module basic_2000_20000_2500_4_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_383,In_1663);
and U1 (N_1,In_1632,In_1299);
nand U2 (N_2,In_1292,In_193);
and U3 (N_3,In_1808,In_1221);
and U4 (N_4,In_1798,In_605);
nor U5 (N_5,In_1262,In_1245);
xor U6 (N_6,In_1651,In_1429);
and U7 (N_7,In_1764,In_1079);
nor U8 (N_8,In_1389,In_361);
or U9 (N_9,In_224,In_228);
nand U10 (N_10,In_1921,In_713);
nand U11 (N_11,In_829,In_1218);
or U12 (N_12,In_32,In_147);
nor U13 (N_13,In_791,In_1633);
xor U14 (N_14,In_660,In_1197);
nor U15 (N_15,In_1065,In_136);
and U16 (N_16,In_1618,In_1029);
or U17 (N_17,In_1511,In_1758);
nand U18 (N_18,In_1031,In_889);
or U19 (N_19,In_1572,In_1027);
or U20 (N_20,In_1432,In_1851);
and U21 (N_21,In_1042,In_1498);
nand U22 (N_22,In_1983,In_1493);
xnor U23 (N_23,In_1509,In_2);
xnor U24 (N_24,In_1222,In_1109);
xor U25 (N_25,In_86,In_1879);
nor U26 (N_26,In_1601,In_807);
and U27 (N_27,In_1490,In_1770);
nor U28 (N_28,In_1642,In_903);
nand U29 (N_29,In_1427,In_1368);
nor U30 (N_30,In_1544,In_1470);
or U31 (N_31,In_644,In_1362);
nor U32 (N_32,In_354,In_1238);
nor U33 (N_33,In_1853,In_684);
and U34 (N_34,In_1112,In_1835);
nand U35 (N_35,In_654,In_1268);
or U36 (N_36,In_1175,In_1820);
nand U37 (N_37,In_1160,In_1384);
nand U38 (N_38,In_1170,In_804);
or U39 (N_39,In_434,In_1837);
or U40 (N_40,In_1423,In_1934);
or U41 (N_41,In_1569,In_1748);
nor U42 (N_42,In_1507,In_194);
or U43 (N_43,In_1884,In_307);
xnor U44 (N_44,In_878,In_1185);
nand U45 (N_45,In_1609,In_1247);
nand U46 (N_46,In_1531,In_1482);
and U47 (N_47,In_1294,In_1319);
xor U48 (N_48,In_497,In_526);
nand U49 (N_49,In_1305,In_152);
nor U50 (N_50,In_853,In_311);
xnor U51 (N_51,In_1785,In_1);
xor U52 (N_52,In_1409,In_864);
nand U53 (N_53,In_1356,In_1577);
xnor U54 (N_54,In_271,In_1426);
nand U55 (N_55,In_337,In_1473);
nand U56 (N_56,In_1043,In_1338);
or U57 (N_57,In_1240,In_603);
or U58 (N_58,In_232,In_388);
nand U59 (N_59,In_1830,In_1462);
nor U60 (N_60,In_783,In_1863);
xor U61 (N_61,In_1888,In_1016);
and U62 (N_62,In_1622,In_1993);
nor U63 (N_63,In_91,In_863);
and U64 (N_64,In_689,In_12);
xor U65 (N_65,In_1745,In_170);
and U66 (N_66,In_20,In_765);
and U67 (N_67,In_1696,In_1492);
nor U68 (N_68,In_1919,In_1720);
xnor U69 (N_69,In_814,In_945);
xnor U70 (N_70,In_1708,In_661);
nor U71 (N_71,In_490,In_49);
nand U72 (N_72,In_191,In_183);
and U73 (N_73,In_1420,In_1290);
and U74 (N_74,In_1495,In_768);
xnor U75 (N_75,In_48,In_1469);
nor U76 (N_76,In_705,In_823);
or U77 (N_77,In_908,In_349);
nor U78 (N_78,In_1710,In_456);
xnor U79 (N_79,In_198,In_930);
nand U80 (N_80,In_1769,In_1539);
nand U81 (N_81,In_1199,In_300);
nand U82 (N_82,In_1334,In_1559);
xnor U83 (N_83,In_769,In_1232);
or U84 (N_84,In_1364,In_1166);
nand U85 (N_85,In_1237,In_229);
and U86 (N_86,In_1717,In_214);
nor U87 (N_87,In_1941,In_1533);
nand U88 (N_88,In_936,In_1840);
nor U89 (N_89,In_1986,In_1719);
or U90 (N_90,In_1760,In_1547);
nand U91 (N_91,In_1737,In_203);
nand U92 (N_92,In_1759,In_1721);
and U93 (N_93,In_18,In_1504);
nand U94 (N_94,In_1455,In_796);
nor U95 (N_95,In_1099,In_1598);
or U96 (N_96,In_1605,In_329);
xor U97 (N_97,In_1126,In_747);
and U98 (N_98,In_698,In_1744);
xor U99 (N_99,In_1591,In_1988);
nor U100 (N_100,In_1475,In_587);
and U101 (N_101,In_101,In_1617);
xnor U102 (N_102,In_1046,In_668);
xor U103 (N_103,In_1214,In_1143);
and U104 (N_104,In_1522,In_1774);
xor U105 (N_105,In_967,In_572);
nand U106 (N_106,In_1589,In_1064);
nand U107 (N_107,In_834,In_1322);
and U108 (N_108,In_1893,In_38);
nor U109 (N_109,In_1897,In_1920);
nor U110 (N_110,In_319,In_1349);
nor U111 (N_111,In_58,In_114);
xnor U112 (N_112,In_536,In_1566);
and U113 (N_113,In_1953,In_272);
nor U114 (N_114,In_14,In_1360);
or U115 (N_115,In_25,In_555);
and U116 (N_116,In_801,In_61);
and U117 (N_117,In_1843,In_31);
nand U118 (N_118,In_797,In_824);
and U119 (N_119,In_657,In_1115);
and U120 (N_120,In_1703,In_1940);
and U121 (N_121,In_714,In_1947);
or U122 (N_122,In_1541,In_1020);
nor U123 (N_123,In_1930,In_391);
nand U124 (N_124,In_1778,In_977);
nand U125 (N_125,In_1107,In_284);
and U126 (N_126,In_1001,In_85);
xnor U127 (N_127,In_763,In_1263);
or U128 (N_128,In_795,In_931);
and U129 (N_129,In_592,In_954);
and U130 (N_130,In_1865,In_1809);
xor U131 (N_131,In_368,In_1603);
nor U132 (N_132,In_1325,In_268);
xnor U133 (N_133,In_1985,In_1416);
or U134 (N_134,In_468,In_1484);
xor U135 (N_135,In_317,In_1480);
nor U136 (N_136,In_827,In_1584);
xnor U137 (N_137,In_932,In_637);
xor U138 (N_138,In_770,In_1549);
xor U139 (N_139,In_1739,In_1053);
and U140 (N_140,In_66,In_1176);
nor U141 (N_141,In_1561,In_169);
and U142 (N_142,In_432,In_586);
nor U143 (N_143,In_1306,In_1188);
nor U144 (N_144,In_1347,In_856);
nand U145 (N_145,In_1844,In_588);
or U146 (N_146,In_543,In_248);
xnor U147 (N_147,In_669,In_47);
nor U148 (N_148,In_1842,In_629);
and U149 (N_149,In_102,In_1873);
xnor U150 (N_150,In_453,In_1724);
nor U151 (N_151,In_1935,In_132);
nor U152 (N_152,In_1510,In_1471);
nand U153 (N_153,In_1520,In_792);
xnor U154 (N_154,In_1406,In_249);
and U155 (N_155,In_609,In_1108);
or U156 (N_156,In_28,In_331);
xor U157 (N_157,In_1731,In_225);
nand U158 (N_158,In_261,In_1984);
nand U159 (N_159,In_1182,In_244);
xor U160 (N_160,In_1151,In_686);
xor U161 (N_161,In_1234,In_794);
and U162 (N_162,In_917,In_1040);
and U163 (N_163,In_1966,In_772);
xnor U164 (N_164,In_607,In_1465);
nor U165 (N_165,In_626,In_699);
xnor U166 (N_166,In_414,In_729);
nand U167 (N_167,In_1678,In_73);
nor U168 (N_168,In_642,In_1265);
xnor U169 (N_169,In_553,In_411);
and U170 (N_170,In_1072,In_700);
nand U171 (N_171,In_335,In_1575);
and U172 (N_172,In_322,In_1912);
and U173 (N_173,In_275,In_480);
or U174 (N_174,In_1258,In_404);
and U175 (N_175,In_1343,In_1383);
nor U176 (N_176,In_315,In_1091);
nand U177 (N_177,In_786,In_719);
nand U178 (N_178,In_995,In_1689);
xor U179 (N_179,In_1171,In_577);
or U180 (N_180,In_761,In_450);
nand U181 (N_181,In_1806,In_1828);
xnor U182 (N_182,In_1574,In_688);
nor U183 (N_183,In_1297,In_905);
nor U184 (N_184,In_1713,In_1230);
and U185 (N_185,In_849,In_1159);
or U186 (N_186,In_133,In_241);
and U187 (N_187,In_323,In_77);
nor U188 (N_188,In_1144,In_882);
or U189 (N_189,In_1316,In_81);
and U190 (N_190,In_1516,In_808);
nand U191 (N_191,In_1960,In_730);
xnor U192 (N_192,In_963,In_172);
or U193 (N_193,In_1179,In_1856);
and U194 (N_194,In_1620,In_1979);
xnor U195 (N_195,In_160,In_1823);
and U196 (N_196,In_993,In_597);
xor U197 (N_197,In_767,In_1335);
nor U198 (N_198,In_1451,In_1747);
nand U199 (N_199,In_563,In_520);
nand U200 (N_200,In_134,In_1148);
and U201 (N_201,In_1336,In_782);
nor U202 (N_202,In_1215,In_491);
and U203 (N_203,In_1363,In_1891);
nand U204 (N_204,In_885,In_234);
or U205 (N_205,In_1366,In_334);
nand U206 (N_206,In_1439,In_659);
xor U207 (N_207,In_466,In_1554);
or U208 (N_208,In_1578,In_1974);
and U209 (N_209,In_1625,In_745);
nor U210 (N_210,In_695,In_98);
and U211 (N_211,In_486,In_940);
xor U212 (N_212,In_70,In_1090);
or U213 (N_213,In_1592,In_624);
or U214 (N_214,In_488,In_619);
nand U215 (N_215,In_1515,In_1468);
or U216 (N_216,In_1180,In_71);
xor U217 (N_217,In_1276,In_1624);
and U218 (N_218,In_1293,In_115);
xnor U219 (N_219,In_645,In_69);
xor U220 (N_220,In_19,In_1525);
and U221 (N_221,In_836,In_1576);
nor U222 (N_222,In_1653,In_1277);
xor U223 (N_223,In_120,In_852);
and U224 (N_224,In_1139,In_1378);
and U225 (N_225,In_515,In_551);
nor U226 (N_226,In_1787,In_1824);
and U227 (N_227,In_1864,In_975);
nor U228 (N_228,In_844,In_1762);
nand U229 (N_229,In_1440,In_922);
and U230 (N_230,In_519,In_816);
xnor U231 (N_231,In_809,In_958);
nor U232 (N_232,In_1519,In_390);
nand U233 (N_233,In_916,In_649);
nor U234 (N_234,In_722,In_848);
and U235 (N_235,In_647,In_387);
nand U236 (N_236,In_1007,In_1838);
and U237 (N_237,In_465,In_288);
nand U238 (N_238,In_646,In_1908);
and U239 (N_239,In_376,In_1892);
nor U240 (N_240,In_1186,In_1801);
or U241 (N_241,In_6,In_446);
or U242 (N_242,In_273,In_1995);
nor U243 (N_243,In_1812,In_1400);
and U244 (N_244,In_1909,In_382);
and U245 (N_245,In_1698,In_327);
nor U246 (N_246,In_1404,In_493);
xor U247 (N_247,In_835,In_535);
and U248 (N_248,In_1975,In_1499);
nand U249 (N_249,In_1560,In_1906);
xnor U250 (N_250,In_4,In_304);
or U251 (N_251,In_1956,In_1877);
nand U252 (N_252,In_1430,In_968);
nand U253 (N_253,In_697,In_1928);
nor U254 (N_254,In_1089,In_1761);
nand U255 (N_255,In_1834,In_1444);
xor U256 (N_256,In_1500,In_1667);
and U257 (N_257,In_727,In_1387);
xor U258 (N_258,In_1847,In_1251);
or U259 (N_259,In_1682,In_1743);
and U260 (N_260,In_427,In_1022);
nand U261 (N_261,In_500,In_1178);
or U262 (N_262,In_417,In_998);
nand U263 (N_263,In_177,In_117);
xor U264 (N_264,In_459,In_1301);
or U265 (N_265,In_1890,In_560);
nand U266 (N_266,In_482,In_29);
nand U267 (N_267,In_1883,In_1303);
and U268 (N_268,In_601,In_986);
or U269 (N_269,In_467,In_1668);
or U270 (N_270,In_630,In_1551);
nand U271 (N_271,In_441,In_328);
nor U272 (N_272,In_620,In_924);
xnor U273 (N_273,In_1055,In_397);
nand U274 (N_274,In_1049,In_1433);
nor U275 (N_275,In_437,In_1540);
or U276 (N_276,In_1716,In_310);
nand U277 (N_277,In_744,In_666);
xor U278 (N_278,In_1639,In_1131);
nor U279 (N_279,In_378,In_556);
nor U280 (N_280,In_359,In_1638);
nand U281 (N_281,In_1375,In_1889);
xor U282 (N_282,In_197,In_1529);
or U283 (N_283,In_1410,In_938);
and U284 (N_284,In_343,In_1715);
nor U285 (N_285,In_1324,In_355);
xor U286 (N_286,In_1248,In_506);
xnor U287 (N_287,In_1196,In_243);
and U288 (N_288,In_1850,In_1125);
nor U289 (N_289,In_919,In_1841);
and U290 (N_290,In_498,In_406);
nor U291 (N_291,In_296,In_281);
nor U292 (N_292,In_352,In_1312);
nand U293 (N_293,In_1777,In_990);
and U294 (N_294,In_1066,In_250);
nand U295 (N_295,In_207,In_693);
and U296 (N_296,In_1944,In_914);
or U297 (N_297,In_1693,In_1738);
or U298 (N_298,In_527,In_8);
and U299 (N_299,In_140,In_939);
and U300 (N_300,In_925,In_1562);
xnor U301 (N_301,In_143,In_217);
nand U302 (N_302,In_943,In_1198);
or U303 (N_303,In_1874,In_186);
xor U304 (N_304,In_1267,In_1355);
and U305 (N_305,In_236,In_1054);
and U306 (N_306,In_580,In_1353);
xor U307 (N_307,In_56,In_1817);
nand U308 (N_308,In_162,In_1780);
xnor U309 (N_309,In_711,In_781);
nand U310 (N_310,In_1580,In_1026);
and U311 (N_311,In_819,In_1573);
nor U312 (N_312,In_1583,In_1431);
nand U313 (N_313,In_156,In_78);
or U314 (N_314,In_1386,In_1189);
and U315 (N_315,In_210,In_596);
and U316 (N_316,In_462,In_308);
nand U317 (N_317,In_704,In_1640);
nand U318 (N_318,In_1311,In_472);
and U319 (N_319,In_350,In_201);
or U320 (N_320,In_706,In_533);
xnor U321 (N_321,In_771,In_868);
nor U322 (N_322,In_737,In_1860);
and U323 (N_323,In_1028,In_1272);
or U324 (N_324,In_692,In_643);
nand U325 (N_325,In_1644,In_176);
nand U326 (N_326,In_84,In_1766);
or U327 (N_327,In_1459,In_982);
xor U328 (N_328,In_1488,In_1942);
nand U329 (N_329,In_1169,In_332);
xor U330 (N_330,In_36,In_1127);
and U331 (N_331,In_1195,In_937);
or U332 (N_332,In_992,In_347);
or U333 (N_333,In_512,In_1287);
nor U334 (N_334,In_608,In_1476);
nand U335 (N_335,In_1217,In_1173);
and U336 (N_336,In_1434,In_1280);
xor U337 (N_337,In_295,In_1628);
xor U338 (N_338,In_1735,In_1463);
xor U339 (N_339,In_1922,In_595);
and U340 (N_340,In_375,In_1978);
or U341 (N_341,In_764,In_1671);
xnor U342 (N_342,In_911,In_530);
nor U343 (N_343,In_57,In_723);
or U344 (N_344,In_1521,In_896);
xnor U345 (N_345,In_534,In_934);
or U346 (N_346,In_1034,In_509);
nand U347 (N_347,In_1315,In_585);
and U348 (N_348,In_1999,In_909);
nor U349 (N_349,In_613,In_72);
xnor U350 (N_350,In_1965,In_1084);
xor U351 (N_351,In_96,In_928);
and U352 (N_352,In_1233,In_145);
or U353 (N_353,In_831,In_1771);
xnor U354 (N_354,In_888,In_1021);
and U355 (N_355,In_658,In_1111);
nand U356 (N_356,In_1997,In_1101);
nand U357 (N_357,In_1105,In_141);
nand U358 (N_358,In_1664,In_1220);
nand U359 (N_359,In_610,In_1792);
nand U360 (N_360,In_1443,In_55);
and U361 (N_361,In_947,In_405);
xor U362 (N_362,In_981,In_178);
or U363 (N_363,In_1943,In_870);
xnor U364 (N_364,In_223,In_3);
nand U365 (N_365,In_436,In_1825);
or U366 (N_366,In_97,In_716);
nand U367 (N_367,In_407,In_1815);
xnor U368 (N_368,In_1226,In_1158);
and U369 (N_369,In_549,In_1381);
and U370 (N_370,In_558,In_805);
and U371 (N_371,In_100,In_87);
or U372 (N_372,In_1514,In_633);
nand U373 (N_373,In_150,In_1636);
nor U374 (N_374,In_1679,In_539);
or U375 (N_375,In_1903,In_1328);
or U376 (N_376,In_113,In_438);
nor U377 (N_377,In_495,In_429);
xor U378 (N_378,In_231,In_1970);
nand U379 (N_379,In_584,In_876);
nand U380 (N_380,In_256,In_664);
nor U381 (N_381,In_672,In_1264);
xor U382 (N_382,In_418,In_205);
xor U383 (N_383,In_392,In_314);
and U384 (N_384,In_1829,In_1948);
nor U385 (N_385,In_1309,In_1058);
nor U386 (N_386,In_1257,In_1795);
nand U387 (N_387,In_615,In_67);
nor U388 (N_388,In_316,In_408);
and U389 (N_389,In_285,In_139);
nor U390 (N_390,In_1550,In_1991);
nor U391 (N_391,In_221,In_1818);
and U392 (N_392,In_972,In_274);
nor U393 (N_393,In_1659,In_1907);
or U394 (N_394,In_1441,In_639);
xnor U395 (N_395,In_1457,In_1448);
or U396 (N_396,In_52,In_421);
nand U397 (N_397,In_1848,In_1813);
or U398 (N_398,In_1969,In_529);
xnor U399 (N_399,In_369,In_13);
nor U400 (N_400,In_1634,In_1933);
nand U401 (N_401,In_1564,In_301);
xnor U402 (N_402,In_1989,In_103);
nand U403 (N_403,In_1587,In_1256);
nor U404 (N_404,In_1749,In_818);
and U405 (N_405,In_1967,In_547);
nor U406 (N_406,In_1085,In_1814);
or U407 (N_407,In_1184,In_865);
and U408 (N_408,In_504,In_676);
nand U409 (N_409,In_1296,In_1610);
and U410 (N_410,In_653,In_1038);
nand U411 (N_411,In_1446,In_460);
xor U412 (N_412,In_1142,In_921);
nor U413 (N_413,In_1757,In_1231);
nor U414 (N_414,In_426,In_1502);
nand U415 (N_415,In_1803,In_1939);
or U416 (N_416,In_1658,In_105);
nor U417 (N_417,In_799,In_531);
nand U418 (N_418,In_1466,In_1726);
xor U419 (N_419,In_173,In_1450);
and U420 (N_420,In_788,In_510);
and U421 (N_421,In_251,In_1900);
and U422 (N_422,In_1076,In_1557);
xor U423 (N_423,In_60,In_253);
or U424 (N_424,In_199,In_395);
nor U425 (N_425,In_1385,In_1790);
xor U426 (N_426,In_528,In_1087);
and U427 (N_427,In_820,In_710);
or U428 (N_428,In_1118,In_1754);
nand U429 (N_429,In_1751,In_1080);
xor U430 (N_430,In_1555,In_1326);
and U431 (N_431,In_1741,In_1819);
xor U432 (N_432,In_1209,In_600);
and U433 (N_433,In_1329,In_1295);
nor U434 (N_434,In_561,In_1260);
xnor U435 (N_435,In_838,In_1310);
nand U436 (N_436,In_302,In_623);
nand U437 (N_437,In_787,In_168);
and U438 (N_438,In_1391,In_1648);
or U439 (N_439,In_444,In_318);
xor U440 (N_440,In_638,In_17);
nor U441 (N_441,In_568,In_1487);
and U442 (N_442,In_1351,In_1223);
xor U443 (N_443,In_1781,In_1119);
or U444 (N_444,In_1902,In_978);
nand U445 (N_445,In_760,In_935);
or U446 (N_446,In_208,In_1784);
nor U447 (N_447,In_442,In_358);
or U448 (N_448,In_1376,In_1302);
nor U449 (N_449,In_184,In_1538);
nor U450 (N_450,In_702,In_1286);
nor U451 (N_451,In_1581,In_1100);
nand U452 (N_452,In_1086,In_479);
and U453 (N_453,In_1200,In_1491);
nor U454 (N_454,In_309,In_1931);
nand U455 (N_455,In_777,In_1661);
nor U456 (N_456,In_1714,In_759);
or U457 (N_457,In_1207,In_1867);
or U458 (N_458,In_743,In_340);
and U459 (N_459,In_1565,In_1097);
nand U460 (N_460,In_1881,In_576);
and U461 (N_461,In_579,In_1202);
xnor U462 (N_462,In_1464,In_1588);
or U463 (N_463,In_1542,In_573);
and U464 (N_464,In_215,In_1036);
nand U465 (N_465,In_1291,In_1567);
or U466 (N_466,In_1646,In_129);
nor U467 (N_467,In_1558,In_1205);
nand U468 (N_468,In_1613,In_1826);
xnor U469 (N_469,In_1008,In_1674);
and U470 (N_470,In_857,In_837);
xnor U471 (N_471,In_1249,In_1904);
or U472 (N_472,In_1796,In_1095);
and U473 (N_473,In_1236,In_1074);
and U474 (N_474,In_1421,In_1155);
xnor U475 (N_475,In_1765,In_641);
and U476 (N_476,In_1137,In_1528);
and U477 (N_477,In_1241,In_109);
xor U478 (N_478,In_1833,In_1616);
nand U479 (N_479,In_953,In_124);
and U480 (N_480,In_1827,In_1120);
xor U481 (N_481,In_82,In_1030);
nor U482 (N_482,In_1050,In_675);
or U483 (N_483,In_123,In_1875);
or U484 (N_484,In_679,In_635);
nand U485 (N_485,In_1138,In_1015);
nor U486 (N_486,In_257,In_738);
xor U487 (N_487,In_196,In_522);
or U488 (N_488,In_800,In_1393);
nor U489 (N_489,In_822,In_627);
xnor U490 (N_490,In_1683,In_1699);
and U491 (N_491,In_1152,In_1686);
nor U492 (N_492,In_701,In_1025);
or U493 (N_493,In_678,In_494);
xor U494 (N_494,In_712,In_1839);
nor U495 (N_495,In_1692,In_1705);
nand U496 (N_496,In_238,In_833);
nand U497 (N_497,In_1987,In_1229);
nor U498 (N_498,In_366,In_190);
nand U499 (N_499,In_1859,In_1783);
and U500 (N_500,In_37,In_1069);
and U501 (N_501,In_1571,In_859);
xor U502 (N_502,In_871,In_1854);
or U503 (N_503,In_433,In_518);
and U504 (N_504,In_1479,In_1358);
xnor U505 (N_505,In_107,In_545);
nor U506 (N_506,In_1243,In_235);
and U507 (N_507,In_267,In_1672);
or U508 (N_508,In_1067,In_1395);
or U509 (N_509,In_1321,In_1377);
and U510 (N_510,In_1361,In_1318);
nand U511 (N_511,In_1782,In_906);
nand U512 (N_512,In_1938,In_1411);
nor U513 (N_513,In_505,In_270);
xnor U514 (N_514,In_381,In_312);
nor U515 (N_515,In_552,In_1298);
nand U516 (N_516,In_1916,In_1009);
nor U517 (N_517,In_696,In_245);
nand U518 (N_518,In_1213,In_557);
and U519 (N_519,In_53,In_1081);
and U520 (N_520,In_46,In_346);
or U521 (N_521,In_326,In_1103);
nand U522 (N_522,In_1534,In_762);
xnor U523 (N_523,In_1611,In_851);
xnor U524 (N_524,In_1821,In_440);
xor U525 (N_525,In_1711,In_1702);
and U526 (N_526,In_1849,In_1971);
nor U527 (N_527,In_35,In_662);
nand U528 (N_528,In_789,In_1918);
and U529 (N_529,In_377,In_632);
nand U530 (N_530,In_1106,In_1637);
xnor U531 (N_531,In_1793,In_1866);
nor U532 (N_532,In_1436,In_1858);
nand U533 (N_533,In_1876,In_1508);
xor U534 (N_534,In_1045,In_1870);
xnor U535 (N_535,In_826,In_1254);
nor U536 (N_536,In_846,In_1503);
or U537 (N_537,In_959,In_1871);
nand U538 (N_538,In_1489,In_736);
nor U539 (N_539,In_1323,In_1786);
and U540 (N_540,In_877,In_734);
or U541 (N_541,In_146,In_1804);
or U542 (N_542,In_1486,In_303);
and U543 (N_543,In_1002,In_1187);
or U544 (N_544,In_1582,In_24);
nor U545 (N_545,In_1006,In_1352);
or U546 (N_546,In_559,In_240);
xnor U547 (N_547,In_341,In_881);
nand U548 (N_548,In_691,In_1271);
and U549 (N_549,In_212,In_474);
nor U550 (N_550,In_866,In_1134);
xnor U551 (N_551,In_324,In_1805);
nor U552 (N_552,In_902,In_900);
or U553 (N_553,In_1852,In_398);
nand U554 (N_554,In_478,In_507);
nand U555 (N_555,In_1946,In_402);
nor U556 (N_556,In_703,In_83);
xor U557 (N_557,In_1212,In_443);
and U558 (N_558,In_1733,In_1163);
and U559 (N_559,In_1371,In_306);
nand U560 (N_560,In_740,In_634);
and U561 (N_561,In_867,In_259);
nor U562 (N_562,In_671,In_246);
xor U563 (N_563,In_1102,In_1915);
xor U564 (N_564,In_1882,In_1802);
or U565 (N_565,In_1597,In_1211);
and U566 (N_566,In_1193,In_904);
and U567 (N_567,In_570,In_1269);
xnor U568 (N_568,In_502,In_969);
nor U569 (N_569,In_1285,In_1905);
or U570 (N_570,In_680,In_987);
or U571 (N_571,In_1590,In_1242);
nand U572 (N_572,In_10,In_1425);
or U573 (N_573,In_127,In_1963);
or U574 (N_574,In_1156,In_1563);
and U575 (N_575,In_631,In_185);
or U576 (N_576,In_65,In_1154);
nor U577 (N_577,In_732,In_891);
or U578 (N_578,In_1730,In_983);
and U579 (N_579,In_915,In_9);
xnor U580 (N_580,In_1373,In_774);
xor U581 (N_581,In_1964,In_989);
or U582 (N_582,In_1895,In_599);
or U583 (N_583,In_283,In_1913);
xor U584 (N_584,In_913,In_1253);
xnor U585 (N_585,In_1899,In_118);
or U586 (N_586,In_521,In_886);
nor U587 (N_587,In_164,In_1958);
and U588 (N_588,In_1901,In_158);
or U589 (N_589,In_575,In_1124);
nor U590 (N_590,In_1308,In_44);
or U591 (N_591,In_99,In_428);
or U592 (N_592,In_1422,In_409);
nand U593 (N_593,In_1691,In_1666);
nor U594 (N_594,In_370,In_22);
and U595 (N_595,In_752,In_1192);
and U596 (N_596,In_1317,In_1401);
nand U597 (N_597,In_1585,In_1024);
or U598 (N_598,In_1756,In_683);
xor U599 (N_599,In_1676,In_30);
and U600 (N_600,In_1768,In_1379);
or U601 (N_601,In_386,In_1394);
nor U602 (N_602,In_1688,In_373);
nor U603 (N_603,In_16,In_1116);
nor U604 (N_604,In_11,In_542);
xor U605 (N_605,In_918,In_458);
or U606 (N_606,In_151,In_1627);
and U607 (N_607,In_640,In_778);
nand U608 (N_608,In_1772,In_1684);
nand U609 (N_609,In_708,In_1657);
nor U610 (N_610,In_277,In_1690);
nand U611 (N_611,In_785,In_1505);
nand U612 (N_612,In_687,In_1130);
and U613 (N_613,In_1478,In_1282);
nand U614 (N_614,In_1135,In_353);
or U615 (N_615,In_1660,In_907);
or U616 (N_616,In_583,In_420);
and U617 (N_617,In_289,In_222);
nor U618 (N_618,In_80,In_1998);
xnor U619 (N_619,In_1675,In_157);
nand U620 (N_620,In_1273,In_298);
and U621 (N_621,In_435,In_230);
nand U622 (N_622,In_999,In_62);
and U623 (N_623,In_1952,In_1797);
and U624 (N_624,In_1374,In_1869);
nor U625 (N_625,In_858,In_735);
or U626 (N_626,In_546,In_1012);
nor U627 (N_627,In_524,In_260);
nand U628 (N_628,In_1773,In_1822);
and U629 (N_629,In_667,In_1145);
xnor U630 (N_630,In_927,In_219);
nor U631 (N_631,In_910,In_1727);
nor U632 (N_632,In_1976,In_548);
nand U633 (N_633,In_1018,In_949);
nor U634 (N_634,In_828,In_707);
and U635 (N_635,In_636,In_1122);
or U636 (N_636,In_1281,In_806);
nand U637 (N_637,In_926,In_1044);
nor U638 (N_638,In_1614,In_1005);
nand U639 (N_639,In_1608,In_1435);
and U640 (N_640,In_34,In_1932);
or U641 (N_641,In_1776,In_401);
and U642 (N_642,In_483,In_255);
nor U643 (N_643,In_110,In_1949);
nand U644 (N_644,In_1167,In_1445);
nand U645 (N_645,In_1398,In_1789);
or U646 (N_646,In_810,In_516);
xnor U647 (N_647,In_299,In_830);
or U648 (N_648,In_424,In_161);
nor U649 (N_649,In_1339,In_278);
nand U650 (N_650,In_1181,In_1161);
or U651 (N_651,In_628,In_276);
xnor U652 (N_652,In_677,In_1062);
nor U653 (N_653,In_1454,In_1593);
nor U654 (N_654,In_1140,In_1685);
and U655 (N_655,In_469,In_1723);
or U656 (N_656,In_1390,In_360);
nor U657 (N_657,In_979,In_192);
xor U658 (N_658,In_1607,In_153);
or U659 (N_659,In_1794,In_1359);
nor U660 (N_660,In_54,In_1252);
and U661 (N_661,In_265,In_455);
and U662 (N_662,In_1996,In_1403);
xnor U663 (N_663,In_717,In_860);
and U664 (N_664,In_1800,In_571);
nor U665 (N_665,In_42,In_1673);
or U666 (N_666,In_503,In_1485);
xor U667 (N_667,In_1951,In_554);
xor U668 (N_668,In_280,In_1862);
nand U669 (N_669,In_1331,In_1235);
or U670 (N_670,In_1397,In_766);
nand U671 (N_671,In_955,In_690);
and U672 (N_672,In_1535,In_652);
and U673 (N_673,In_293,In_475);
and U674 (N_674,In_144,In_1496);
and U675 (N_675,In_1153,In_1619);
nor U676 (N_676,In_188,In_1532);
or U677 (N_677,In_872,In_965);
or U678 (N_678,In_754,In_1010);
and U679 (N_679,In_220,In_1959);
nand U680 (N_680,In_724,In_976);
and U681 (N_681,In_980,In_1057);
and U682 (N_682,In_685,In_1048);
xnor U683 (N_683,In_461,In_1442);
nand U684 (N_684,In_477,In_892);
nand U685 (N_685,In_1052,In_845);
or U686 (N_686,In_452,In_496);
nand U687 (N_687,In_1512,In_1687);
or U688 (N_688,In_362,In_798);
and U689 (N_689,In_1344,In_884);
and U690 (N_690,In_1545,In_108);
or U691 (N_691,In_1011,In_957);
nand U692 (N_692,In_447,In_1340);
and U693 (N_693,In_1071,In_1526);
nand U694 (N_694,In_1073,In_1501);
and U695 (N_695,In_1168,In_746);
and U696 (N_696,In_379,In_1289);
nand U697 (N_697,In_951,In_1936);
nand U698 (N_698,In_1146,In_1437);
nand U699 (N_699,In_840,In_1707);
and U700 (N_700,In_23,In_451);
nand U701 (N_701,In_523,In_1700);
or U702 (N_702,In_264,In_1811);
or U703 (N_703,In_753,In_1228);
or U704 (N_704,In_562,In_758);
xor U705 (N_705,In_879,In_399);
nand U706 (N_706,In_1694,In_650);
nor U707 (N_707,In_1275,In_345);
xnor U708 (N_708,In_365,In_1051);
and U709 (N_709,In_811,In_880);
nor U710 (N_710,In_1586,In_971);
or U711 (N_711,In_991,In_448);
nor U712 (N_712,In_126,In_1506);
nand U713 (N_713,In_1530,In_890);
or U714 (N_714,In_1300,In_540);
or U715 (N_715,In_492,In_39);
or U716 (N_716,In_751,In_725);
nor U717 (N_717,In_1396,In_1579);
xor U718 (N_718,In_122,In_1408);
nor U719 (N_719,In_202,In_457);
or U720 (N_720,In_1078,In_912);
and U721 (N_721,In_1924,In_517);
nand U722 (N_722,In_718,In_393);
xnor U723 (N_723,In_90,In_1227);
or U724 (N_724,In_755,In_422);
or U725 (N_725,In_1740,In_855);
and U726 (N_726,In_1370,In_1606);
nor U727 (N_727,In_1654,In_1481);
nand U728 (N_728,In_602,In_445);
or U729 (N_729,In_893,In_1973);
xnor U730 (N_730,In_944,In_1244);
or U731 (N_731,In_1157,In_1548);
or U732 (N_732,In_742,In_68);
nand U733 (N_733,In_1225,In_330);
xnor U734 (N_734,In_1923,In_51);
nor U735 (N_735,In_1483,In_897);
and U736 (N_736,In_843,In_1494);
and U737 (N_737,In_1746,In_1035);
nand U738 (N_738,In_581,In_1517);
or U739 (N_739,In_484,In_883);
nor U740 (N_740,In_1023,In_682);
xor U741 (N_741,In_1133,In_95);
nor U742 (N_742,In_279,In_1259);
nand U743 (N_743,In_1472,In_1424);
or U744 (N_744,In_1467,In_50);
or U745 (N_745,In_1621,In_1128);
nor U746 (N_746,In_1041,In_104);
nand U747 (N_747,In_513,In_933);
nand U748 (N_748,In_396,In_748);
nor U749 (N_749,In_1599,In_1104);
and U750 (N_750,In_1372,In_1060);
nor U751 (N_751,In_471,In_1350);
xnor U752 (N_752,In_204,In_1246);
nor U753 (N_753,In_1438,In_1070);
nor U754 (N_754,In_1527,In_487);
and U755 (N_755,In_1878,In_1742);
and U756 (N_756,In_290,In_159);
xor U757 (N_757,In_1736,In_1330);
or U758 (N_758,In_813,In_1458);
and U759 (N_759,In_1641,In_593);
xnor U760 (N_760,In_1414,In_1831);
and U761 (N_761,In_812,In_1791);
nor U762 (N_762,In_1077,In_663);
and U763 (N_763,In_1652,In_1898);
and U764 (N_764,In_1655,In_1278);
nor U765 (N_765,In_356,In_282);
xnor U766 (N_766,In_617,In_1556);
xnor U767 (N_767,In_403,In_621);
nand U768 (N_768,In_1183,In_1643);
xnor U769 (N_769,In_1650,In_1357);
xnor U770 (N_770,In_1885,In_1845);
and U771 (N_771,In_749,In_1734);
and U772 (N_772,In_166,In_720);
xor U773 (N_773,In_1210,In_1722);
nand U774 (N_774,In_1524,In_739);
nand U775 (N_775,In_1968,In_694);
or U776 (N_776,In_1855,In_1706);
xnor U777 (N_777,In_415,In_862);
xnor U778 (N_778,In_1039,In_363);
nor U779 (N_779,In_213,In_923);
nor U780 (N_780,In_348,In_394);
xnor U781 (N_781,In_1341,In_262);
nor U782 (N_782,In_1543,In_1239);
xnor U783 (N_783,In_1255,In_1162);
and U784 (N_784,In_15,In_1013);
nor U785 (N_785,In_165,In_1615);
or U786 (N_786,In_1113,In_266);
nor U787 (N_787,In_594,In_1752);
xnor U788 (N_788,In_1354,In_962);
and U789 (N_789,In_413,In_179);
xnor U790 (N_790,In_715,In_1216);
and U791 (N_791,In_131,In_1836);
xnor U792 (N_792,In_112,In_952);
xor U793 (N_793,In_1121,In_1019);
and U794 (N_794,In_1003,In_1098);
nand U795 (N_795,In_591,In_1419);
xor U796 (N_796,In_750,In_1096);
and U797 (N_797,In_832,In_119);
and U798 (N_798,In_1807,In_364);
nand U799 (N_799,In_1190,In_1645);
xnor U800 (N_800,In_1136,In_1763);
and U801 (N_801,In_454,In_167);
nor U802 (N_802,In_532,In_473);
and U803 (N_803,In_508,In_1937);
xnor U804 (N_804,In_726,In_1872);
and U805 (N_805,In_239,In_622);
xor U806 (N_806,In_64,In_1452);
nand U807 (N_807,In_227,In_793);
nand U808 (N_808,In_681,In_875);
xnor U809 (N_809,In_94,In_970);
xnor U810 (N_810,In_1709,In_1894);
nor U811 (N_811,In_294,In_449);
xor U812 (N_812,In_1092,In_1961);
and U813 (N_813,In_389,In_0);
nand U814 (N_814,In_374,In_1447);
xnor U815 (N_815,In_1656,In_1513);
xnor U816 (N_816,In_574,In_1047);
nor U817 (N_817,In_1728,In_898);
nand U818 (N_818,In_138,In_297);
and U819 (N_819,In_357,In_1954);
nor U820 (N_820,In_216,In_1816);
xor U821 (N_821,In_180,In_135);
nand U822 (N_822,In_899,In_489);
nor U823 (N_823,In_1313,In_149);
nand U824 (N_824,In_775,In_63);
xor U825 (N_825,In_861,In_1382);
xnor U826 (N_826,In_1604,In_1333);
nand U827 (N_827,In_1164,In_412);
nand U828 (N_828,In_1596,In_33);
nor U829 (N_829,In_339,In_1224);
nor U830 (N_830,In_1950,In_929);
nand U831 (N_831,In_1695,In_1868);
or U832 (N_832,In_269,In_1061);
or U833 (N_833,In_1453,In_1266);
or U834 (N_834,In_137,In_994);
nand U835 (N_835,In_1456,In_154);
or U836 (N_836,In_1304,In_1346);
nor U837 (N_837,In_1075,In_606);
and U838 (N_838,In_1402,In_385);
nor U839 (N_839,In_566,In_1288);
and U840 (N_840,In_195,In_950);
and U841 (N_841,In_92,In_1083);
or U842 (N_842,In_985,In_733);
xor U843 (N_843,In_1208,In_1004);
and U844 (N_844,In_1981,In_321);
xnor U845 (N_845,In_1880,In_1415);
xnor U846 (N_846,In_1460,In_416);
nand U847 (N_847,In_1332,In_1595);
or U848 (N_848,In_901,In_757);
and U849 (N_849,In_670,In_1203);
and U850 (N_850,In_1788,In_651);
nor U851 (N_851,In_1594,In_1365);
and U852 (N_852,In_839,In_88);
xnor U853 (N_853,In_887,In_589);
nor U854 (N_854,In_1206,In_351);
and U855 (N_855,In_336,In_130);
xnor U856 (N_856,In_1150,In_1732);
nor U857 (N_857,In_1523,In_1068);
and U858 (N_858,In_956,In_1380);
nand U859 (N_859,In_1094,In_286);
or U860 (N_860,In_964,In_1412);
nor U861 (N_861,In_5,In_1925);
or U862 (N_862,In_1388,In_1201);
nor U863 (N_863,In_525,In_1477);
nand U864 (N_864,In_1037,In_292);
and U865 (N_865,In_1093,In_1194);
nand U866 (N_866,In_1250,In_1910);
nand U867 (N_867,In_815,In_1337);
or U868 (N_868,In_233,In_1418);
and U869 (N_869,In_200,In_1629);
or U870 (N_870,In_463,In_1413);
nor U871 (N_871,In_973,In_59);
or U872 (N_872,In_121,In_252);
and U873 (N_873,In_537,In_1342);
or U874 (N_874,In_1407,In_590);
xnor U875 (N_875,In_1320,In_1123);
and U876 (N_876,In_665,In_578);
and U877 (N_877,In_1082,In_1327);
nand U878 (N_878,In_776,In_996);
or U879 (N_879,In_565,In_1141);
xor U880 (N_880,In_1191,In_1177);
xnor U881 (N_881,In_1274,In_1110);
nand U882 (N_882,In_226,In_655);
nor U883 (N_883,In_181,In_1367);
nand U884 (N_884,In_1552,In_1755);
or U885 (N_885,In_784,In_1729);
nand U886 (N_886,In_1977,In_802);
nor U887 (N_887,In_780,In_1857);
nor U888 (N_888,In_419,In_1172);
or U889 (N_889,In_1568,In_174);
or U890 (N_890,In_821,In_325);
nand U891 (N_891,In_263,In_1635);
nor U892 (N_892,In_1307,In_779);
xnor U893 (N_893,In_1063,In_287);
nor U894 (N_894,In_410,In_501);
nand U895 (N_895,In_1000,In_1174);
nand U896 (N_896,In_372,In_320);
xor U897 (N_897,In_1750,In_1701);
or U898 (N_898,In_514,In_1861);
xnor U899 (N_899,In_773,In_342);
nand U900 (N_900,In_1132,In_182);
and U901 (N_901,In_187,In_305);
nor U902 (N_902,In_1926,In_869);
nand U903 (N_903,In_564,In_1270);
xnor U904 (N_904,In_841,In_1314);
nor U905 (N_905,In_1670,In_1896);
nor U906 (N_906,In_1114,In_895);
xor U907 (N_907,In_254,In_1348);
or U908 (N_908,In_1725,In_1810);
nand U909 (N_909,In_431,In_920);
xor U910 (N_910,In_400,In_189);
nor U911 (N_911,In_1990,In_1546);
nand U912 (N_912,In_946,In_430);
xnor U913 (N_913,In_873,In_1056);
or U914 (N_914,In_611,In_481);
nor U915 (N_915,In_1681,In_1626);
or U916 (N_916,In_544,In_45);
nor U917 (N_917,In_464,In_1980);
nand U918 (N_918,In_1704,In_485);
nor U919 (N_919,In_756,In_538);
and U920 (N_920,In_206,In_1887);
nand U921 (N_921,In_1059,In_1886);
nand U922 (N_922,In_1662,In_1630);
xnor U923 (N_923,In_27,In_1449);
or U924 (N_924,In_1767,In_1846);
nand U925 (N_925,In_616,In_211);
or U926 (N_926,In_741,In_380);
nor U927 (N_927,In_1518,In_218);
and U928 (N_928,In_21,In_439);
xnor U929 (N_929,In_338,In_242);
xnor U930 (N_930,In_1405,In_850);
xor U931 (N_931,In_1033,In_76);
and U932 (N_932,In_984,In_1219);
or U933 (N_933,In_1718,In_1392);
or U934 (N_934,In_1117,In_550);
or U935 (N_935,In_1602,In_1345);
nor U936 (N_936,In_1399,In_1911);
xor U937 (N_937,In_89,In_128);
or U938 (N_938,In_476,In_155);
and U939 (N_939,In_825,In_1088);
or U940 (N_940,In_1284,In_1832);
nor U941 (N_941,In_648,In_1129);
nor U942 (N_942,In_1665,In_1497);
nand U943 (N_943,In_1917,In_817);
and U944 (N_944,In_1204,In_709);
nor U945 (N_945,In_948,In_598);
or U946 (N_946,In_40,In_371);
nand U947 (N_947,In_74,In_790);
or U948 (N_948,In_569,In_499);
xnor U949 (N_949,In_1647,In_941);
xor U950 (N_950,In_961,In_1955);
xor U951 (N_951,In_1775,In_344);
nand U952 (N_952,In_974,In_1570);
xor U953 (N_953,In_26,In_313);
xor U954 (N_954,In_43,In_384);
and U955 (N_955,In_163,In_1779);
nor U956 (N_956,In_1631,In_1017);
xor U957 (N_957,In_1537,In_106);
and U958 (N_958,In_291,In_116);
nand U959 (N_959,In_842,In_333);
xnor U960 (N_960,In_1461,In_966);
xor U961 (N_961,In_1914,In_1994);
nand U962 (N_962,In_1945,In_511);
xor U963 (N_963,In_423,In_258);
or U964 (N_964,In_942,In_847);
nand U965 (N_965,In_731,In_854);
nor U966 (N_966,In_1032,In_148);
nor U967 (N_967,In_1279,In_367);
and U968 (N_968,In_142,In_1669);
nor U969 (N_969,In_604,In_470);
and U970 (N_970,In_612,In_567);
nor U971 (N_971,In_1283,In_1014);
or U972 (N_972,In_1261,In_874);
or U973 (N_973,In_1417,In_1957);
xor U974 (N_974,In_960,In_1474);
nor U975 (N_975,In_625,In_1649);
nor U976 (N_976,In_1165,In_79);
and U977 (N_977,In_997,In_1369);
and U978 (N_978,In_7,In_894);
and U979 (N_979,In_1712,In_93);
or U980 (N_980,In_674,In_803);
and U981 (N_981,In_209,In_425);
xnor U982 (N_982,In_673,In_1972);
or U983 (N_983,In_1799,In_111);
xnor U984 (N_984,In_1697,In_728);
and U985 (N_985,In_1680,In_656);
and U986 (N_986,In_1147,In_541);
nor U987 (N_987,In_1982,In_1753);
and U988 (N_988,In_1149,In_1553);
and U989 (N_989,In_1929,In_1962);
nor U990 (N_990,In_1677,In_614);
or U991 (N_991,In_721,In_1428);
nor U992 (N_992,In_171,In_1927);
nand U993 (N_993,In_988,In_1623);
nand U994 (N_994,In_582,In_1600);
and U995 (N_995,In_175,In_247);
or U996 (N_996,In_237,In_618);
nand U997 (N_997,In_125,In_1612);
and U998 (N_998,In_1536,In_41);
nand U999 (N_999,In_1992,In_75);
or U1000 (N_1000,In_555,In_270);
nand U1001 (N_1001,In_457,In_1884);
or U1002 (N_1002,In_882,In_925);
nor U1003 (N_1003,In_1291,In_1367);
xor U1004 (N_1004,In_1740,In_1458);
or U1005 (N_1005,In_138,In_756);
xnor U1006 (N_1006,In_1962,In_1537);
and U1007 (N_1007,In_1922,In_1207);
nor U1008 (N_1008,In_803,In_960);
xnor U1009 (N_1009,In_1904,In_152);
or U1010 (N_1010,In_548,In_1344);
nand U1011 (N_1011,In_904,In_11);
and U1012 (N_1012,In_717,In_844);
nor U1013 (N_1013,In_1450,In_684);
nand U1014 (N_1014,In_1463,In_1286);
or U1015 (N_1015,In_812,In_152);
nand U1016 (N_1016,In_1255,In_998);
xnor U1017 (N_1017,In_417,In_1482);
xor U1018 (N_1018,In_1482,In_806);
nand U1019 (N_1019,In_1179,In_432);
or U1020 (N_1020,In_1220,In_4);
xor U1021 (N_1021,In_1099,In_626);
or U1022 (N_1022,In_1186,In_945);
nor U1023 (N_1023,In_1863,In_1796);
nand U1024 (N_1024,In_992,In_1104);
and U1025 (N_1025,In_401,In_1252);
and U1026 (N_1026,In_1687,In_1556);
nand U1027 (N_1027,In_232,In_856);
and U1028 (N_1028,In_1179,In_141);
or U1029 (N_1029,In_23,In_379);
xnor U1030 (N_1030,In_75,In_1901);
xnor U1031 (N_1031,In_1871,In_1417);
nor U1032 (N_1032,In_1849,In_1144);
or U1033 (N_1033,In_1226,In_1174);
or U1034 (N_1034,In_1362,In_13);
nand U1035 (N_1035,In_1938,In_174);
nor U1036 (N_1036,In_1978,In_1515);
nand U1037 (N_1037,In_1387,In_284);
xor U1038 (N_1038,In_357,In_1531);
xnor U1039 (N_1039,In_914,In_933);
or U1040 (N_1040,In_1028,In_1009);
nor U1041 (N_1041,In_1440,In_1098);
nand U1042 (N_1042,In_1926,In_486);
xor U1043 (N_1043,In_1650,In_1237);
or U1044 (N_1044,In_1392,In_1496);
xor U1045 (N_1045,In_298,In_695);
or U1046 (N_1046,In_96,In_1648);
nand U1047 (N_1047,In_1321,In_538);
and U1048 (N_1048,In_377,In_1113);
nand U1049 (N_1049,In_1009,In_947);
nor U1050 (N_1050,In_1674,In_1557);
and U1051 (N_1051,In_1201,In_919);
xor U1052 (N_1052,In_1457,In_185);
and U1053 (N_1053,In_234,In_1390);
or U1054 (N_1054,In_1817,In_1505);
or U1055 (N_1055,In_260,In_1967);
nand U1056 (N_1056,In_1480,In_1564);
xnor U1057 (N_1057,In_305,In_999);
xor U1058 (N_1058,In_840,In_1315);
and U1059 (N_1059,In_68,In_970);
and U1060 (N_1060,In_280,In_648);
and U1061 (N_1061,In_1251,In_717);
or U1062 (N_1062,In_1883,In_1961);
nor U1063 (N_1063,In_336,In_317);
or U1064 (N_1064,In_1892,In_1366);
nand U1065 (N_1065,In_1356,In_1576);
xor U1066 (N_1066,In_1367,In_786);
or U1067 (N_1067,In_820,In_801);
nand U1068 (N_1068,In_803,In_570);
and U1069 (N_1069,In_435,In_1679);
nor U1070 (N_1070,In_212,In_1844);
nor U1071 (N_1071,In_1642,In_325);
xor U1072 (N_1072,In_1336,In_946);
or U1073 (N_1073,In_278,In_962);
and U1074 (N_1074,In_929,In_1610);
or U1075 (N_1075,In_586,In_624);
xnor U1076 (N_1076,In_1779,In_33);
nor U1077 (N_1077,In_1813,In_1758);
nor U1078 (N_1078,In_447,In_1310);
nand U1079 (N_1079,In_723,In_275);
xor U1080 (N_1080,In_29,In_181);
xnor U1081 (N_1081,In_144,In_435);
and U1082 (N_1082,In_1920,In_1033);
and U1083 (N_1083,In_1932,In_844);
nand U1084 (N_1084,In_1555,In_325);
xnor U1085 (N_1085,In_467,In_793);
xor U1086 (N_1086,In_1203,In_449);
and U1087 (N_1087,In_825,In_1884);
and U1088 (N_1088,In_1972,In_276);
nand U1089 (N_1089,In_523,In_645);
nand U1090 (N_1090,In_1765,In_1354);
and U1091 (N_1091,In_425,In_455);
nor U1092 (N_1092,In_814,In_1375);
and U1093 (N_1093,In_200,In_434);
nor U1094 (N_1094,In_70,In_915);
nand U1095 (N_1095,In_1699,In_1906);
or U1096 (N_1096,In_822,In_1087);
xnor U1097 (N_1097,In_1435,In_1524);
and U1098 (N_1098,In_257,In_586);
and U1099 (N_1099,In_1525,In_151);
or U1100 (N_1100,In_219,In_1992);
or U1101 (N_1101,In_782,In_330);
xnor U1102 (N_1102,In_1306,In_854);
xor U1103 (N_1103,In_198,In_329);
nor U1104 (N_1104,In_1949,In_607);
or U1105 (N_1105,In_1517,In_103);
and U1106 (N_1106,In_796,In_1339);
xnor U1107 (N_1107,In_996,In_394);
or U1108 (N_1108,In_182,In_401);
nand U1109 (N_1109,In_1166,In_1249);
nand U1110 (N_1110,In_1766,In_1545);
nand U1111 (N_1111,In_444,In_1868);
nand U1112 (N_1112,In_1774,In_262);
nor U1113 (N_1113,In_1389,In_838);
or U1114 (N_1114,In_529,In_844);
xor U1115 (N_1115,In_1075,In_1499);
xor U1116 (N_1116,In_402,In_237);
nor U1117 (N_1117,In_1762,In_1150);
nand U1118 (N_1118,In_1712,In_1498);
nand U1119 (N_1119,In_672,In_630);
nand U1120 (N_1120,In_727,In_456);
nor U1121 (N_1121,In_502,In_1295);
nor U1122 (N_1122,In_586,In_1281);
and U1123 (N_1123,In_552,In_509);
or U1124 (N_1124,In_594,In_1859);
and U1125 (N_1125,In_499,In_108);
xor U1126 (N_1126,In_1546,In_1297);
nand U1127 (N_1127,In_435,In_849);
or U1128 (N_1128,In_1759,In_1031);
nand U1129 (N_1129,In_1252,In_1247);
or U1130 (N_1130,In_1742,In_1507);
and U1131 (N_1131,In_53,In_1608);
xnor U1132 (N_1132,In_1735,In_1648);
or U1133 (N_1133,In_1251,In_965);
nor U1134 (N_1134,In_1367,In_798);
and U1135 (N_1135,In_1068,In_1574);
and U1136 (N_1136,In_152,In_17);
nor U1137 (N_1137,In_881,In_1296);
xnor U1138 (N_1138,In_862,In_406);
and U1139 (N_1139,In_1851,In_733);
xnor U1140 (N_1140,In_1922,In_1149);
nor U1141 (N_1141,In_1084,In_1305);
xor U1142 (N_1142,In_927,In_605);
and U1143 (N_1143,In_957,In_310);
nor U1144 (N_1144,In_676,In_712);
xnor U1145 (N_1145,In_1158,In_386);
and U1146 (N_1146,In_1048,In_152);
xor U1147 (N_1147,In_732,In_491);
or U1148 (N_1148,In_1737,In_1462);
xor U1149 (N_1149,In_528,In_308);
and U1150 (N_1150,In_228,In_1416);
xor U1151 (N_1151,In_1061,In_558);
nand U1152 (N_1152,In_867,In_420);
xnor U1153 (N_1153,In_1626,In_1249);
or U1154 (N_1154,In_1430,In_50);
xor U1155 (N_1155,In_1085,In_1795);
or U1156 (N_1156,In_294,In_1517);
and U1157 (N_1157,In_64,In_683);
xor U1158 (N_1158,In_213,In_1247);
xor U1159 (N_1159,In_1208,In_156);
nand U1160 (N_1160,In_167,In_1669);
xnor U1161 (N_1161,In_1789,In_655);
nand U1162 (N_1162,In_47,In_125);
nand U1163 (N_1163,In_1630,In_589);
nor U1164 (N_1164,In_1589,In_1920);
xor U1165 (N_1165,In_343,In_1538);
and U1166 (N_1166,In_1328,In_1579);
or U1167 (N_1167,In_704,In_888);
nand U1168 (N_1168,In_1285,In_1302);
nand U1169 (N_1169,In_1198,In_64);
nand U1170 (N_1170,In_272,In_785);
xnor U1171 (N_1171,In_293,In_980);
nand U1172 (N_1172,In_621,In_1100);
or U1173 (N_1173,In_1667,In_853);
and U1174 (N_1174,In_243,In_1314);
and U1175 (N_1175,In_1429,In_1523);
or U1176 (N_1176,In_359,In_1405);
or U1177 (N_1177,In_1212,In_205);
xnor U1178 (N_1178,In_35,In_113);
nand U1179 (N_1179,In_1217,In_130);
nor U1180 (N_1180,In_573,In_1739);
and U1181 (N_1181,In_624,In_781);
xnor U1182 (N_1182,In_167,In_1301);
or U1183 (N_1183,In_1249,In_1341);
xor U1184 (N_1184,In_543,In_1957);
and U1185 (N_1185,In_809,In_190);
or U1186 (N_1186,In_1037,In_1349);
nand U1187 (N_1187,In_1564,In_380);
nand U1188 (N_1188,In_467,In_1752);
nand U1189 (N_1189,In_719,In_1558);
nor U1190 (N_1190,In_1798,In_760);
and U1191 (N_1191,In_757,In_1816);
and U1192 (N_1192,In_491,In_7);
nand U1193 (N_1193,In_1863,In_388);
nand U1194 (N_1194,In_1091,In_1275);
and U1195 (N_1195,In_1653,In_1608);
nand U1196 (N_1196,In_335,In_1623);
and U1197 (N_1197,In_1187,In_824);
nand U1198 (N_1198,In_885,In_1788);
or U1199 (N_1199,In_386,In_380);
and U1200 (N_1200,In_465,In_471);
nand U1201 (N_1201,In_1454,In_499);
or U1202 (N_1202,In_1885,In_873);
or U1203 (N_1203,In_352,In_1681);
nor U1204 (N_1204,In_1791,In_314);
and U1205 (N_1205,In_609,In_286);
or U1206 (N_1206,In_417,In_1681);
and U1207 (N_1207,In_603,In_894);
xnor U1208 (N_1208,In_1834,In_400);
nand U1209 (N_1209,In_1221,In_1293);
and U1210 (N_1210,In_1891,In_671);
xnor U1211 (N_1211,In_919,In_1199);
or U1212 (N_1212,In_1213,In_1532);
xnor U1213 (N_1213,In_1034,In_1455);
or U1214 (N_1214,In_348,In_897);
or U1215 (N_1215,In_1768,In_916);
xnor U1216 (N_1216,In_56,In_1833);
nand U1217 (N_1217,In_281,In_1665);
nor U1218 (N_1218,In_1239,In_377);
and U1219 (N_1219,In_1319,In_1456);
nand U1220 (N_1220,In_1518,In_719);
and U1221 (N_1221,In_1550,In_437);
xor U1222 (N_1222,In_749,In_1269);
xor U1223 (N_1223,In_837,In_280);
xor U1224 (N_1224,In_1535,In_1886);
nor U1225 (N_1225,In_140,In_1441);
xnor U1226 (N_1226,In_1677,In_152);
and U1227 (N_1227,In_381,In_636);
nand U1228 (N_1228,In_1256,In_114);
xor U1229 (N_1229,In_771,In_548);
and U1230 (N_1230,In_709,In_1896);
and U1231 (N_1231,In_220,In_1315);
nand U1232 (N_1232,In_1670,In_1236);
or U1233 (N_1233,In_1768,In_1894);
xor U1234 (N_1234,In_1508,In_204);
or U1235 (N_1235,In_1304,In_680);
and U1236 (N_1236,In_1831,In_88);
nand U1237 (N_1237,In_1263,In_1069);
nor U1238 (N_1238,In_1398,In_283);
and U1239 (N_1239,In_17,In_75);
nor U1240 (N_1240,In_1308,In_1527);
or U1241 (N_1241,In_1385,In_498);
nor U1242 (N_1242,In_1251,In_657);
or U1243 (N_1243,In_450,In_225);
xnor U1244 (N_1244,In_143,In_1778);
nand U1245 (N_1245,In_1933,In_173);
nor U1246 (N_1246,In_1714,In_452);
nand U1247 (N_1247,In_471,In_249);
xor U1248 (N_1248,In_516,In_450);
nand U1249 (N_1249,In_590,In_1156);
xnor U1250 (N_1250,In_1521,In_184);
xor U1251 (N_1251,In_1862,In_609);
and U1252 (N_1252,In_866,In_1671);
and U1253 (N_1253,In_704,In_1373);
or U1254 (N_1254,In_1740,In_621);
and U1255 (N_1255,In_1739,In_904);
and U1256 (N_1256,In_572,In_343);
xnor U1257 (N_1257,In_442,In_1097);
xor U1258 (N_1258,In_1648,In_1682);
and U1259 (N_1259,In_1465,In_1891);
nand U1260 (N_1260,In_149,In_964);
and U1261 (N_1261,In_1802,In_1028);
nand U1262 (N_1262,In_413,In_1881);
and U1263 (N_1263,In_389,In_1873);
nor U1264 (N_1264,In_14,In_523);
and U1265 (N_1265,In_1566,In_421);
or U1266 (N_1266,In_613,In_1568);
xnor U1267 (N_1267,In_1198,In_1950);
or U1268 (N_1268,In_177,In_690);
xnor U1269 (N_1269,In_1722,In_639);
xor U1270 (N_1270,In_1853,In_12);
xor U1271 (N_1271,In_370,In_131);
xnor U1272 (N_1272,In_670,In_699);
nor U1273 (N_1273,In_1925,In_93);
nor U1274 (N_1274,In_35,In_1119);
nand U1275 (N_1275,In_1731,In_1482);
xor U1276 (N_1276,In_383,In_1703);
xnor U1277 (N_1277,In_262,In_809);
nor U1278 (N_1278,In_622,In_174);
and U1279 (N_1279,In_1028,In_666);
and U1280 (N_1280,In_596,In_198);
and U1281 (N_1281,In_1726,In_713);
nand U1282 (N_1282,In_1025,In_940);
nor U1283 (N_1283,In_269,In_1476);
and U1284 (N_1284,In_982,In_1657);
nand U1285 (N_1285,In_981,In_938);
xnor U1286 (N_1286,In_346,In_595);
or U1287 (N_1287,In_1009,In_1946);
and U1288 (N_1288,In_1309,In_519);
nor U1289 (N_1289,In_540,In_482);
and U1290 (N_1290,In_711,In_289);
nand U1291 (N_1291,In_1843,In_1437);
nor U1292 (N_1292,In_1004,In_288);
and U1293 (N_1293,In_1293,In_1709);
or U1294 (N_1294,In_1714,In_379);
nand U1295 (N_1295,In_304,In_1111);
xor U1296 (N_1296,In_211,In_1975);
nand U1297 (N_1297,In_494,In_327);
nand U1298 (N_1298,In_334,In_44);
and U1299 (N_1299,In_208,In_1005);
nand U1300 (N_1300,In_1365,In_486);
nand U1301 (N_1301,In_414,In_434);
xor U1302 (N_1302,In_1267,In_1387);
nor U1303 (N_1303,In_1549,In_1624);
and U1304 (N_1304,In_1495,In_344);
or U1305 (N_1305,In_1227,In_1634);
and U1306 (N_1306,In_802,In_955);
nor U1307 (N_1307,In_818,In_932);
xor U1308 (N_1308,In_1108,In_790);
nand U1309 (N_1309,In_654,In_422);
or U1310 (N_1310,In_1939,In_499);
nand U1311 (N_1311,In_863,In_1256);
xor U1312 (N_1312,In_878,In_1117);
nand U1313 (N_1313,In_1944,In_405);
and U1314 (N_1314,In_214,In_1625);
and U1315 (N_1315,In_1256,In_1942);
nor U1316 (N_1316,In_1565,In_1247);
and U1317 (N_1317,In_1036,In_1625);
and U1318 (N_1318,In_146,In_1142);
or U1319 (N_1319,In_638,In_692);
nor U1320 (N_1320,In_1148,In_1540);
xnor U1321 (N_1321,In_936,In_795);
nand U1322 (N_1322,In_1479,In_1699);
nand U1323 (N_1323,In_1255,In_1020);
nand U1324 (N_1324,In_1922,In_667);
and U1325 (N_1325,In_1533,In_775);
nor U1326 (N_1326,In_1428,In_779);
or U1327 (N_1327,In_1642,In_821);
xnor U1328 (N_1328,In_32,In_751);
or U1329 (N_1329,In_995,In_1105);
or U1330 (N_1330,In_1365,In_1617);
and U1331 (N_1331,In_1801,In_1837);
xor U1332 (N_1332,In_798,In_811);
nor U1333 (N_1333,In_1420,In_1649);
xor U1334 (N_1334,In_1360,In_742);
xnor U1335 (N_1335,In_1110,In_354);
or U1336 (N_1336,In_1181,In_283);
and U1337 (N_1337,In_1473,In_1200);
and U1338 (N_1338,In_760,In_1515);
or U1339 (N_1339,In_619,In_723);
and U1340 (N_1340,In_1047,In_1938);
or U1341 (N_1341,In_1293,In_804);
or U1342 (N_1342,In_443,In_561);
nand U1343 (N_1343,In_556,In_724);
nand U1344 (N_1344,In_288,In_1075);
or U1345 (N_1345,In_1926,In_1894);
and U1346 (N_1346,In_291,In_815);
nand U1347 (N_1347,In_1386,In_179);
xnor U1348 (N_1348,In_20,In_395);
xor U1349 (N_1349,In_1929,In_78);
or U1350 (N_1350,In_1157,In_1283);
xor U1351 (N_1351,In_387,In_483);
or U1352 (N_1352,In_908,In_1895);
xor U1353 (N_1353,In_1369,In_266);
and U1354 (N_1354,In_1644,In_875);
or U1355 (N_1355,In_1751,In_1381);
or U1356 (N_1356,In_1021,In_650);
or U1357 (N_1357,In_1512,In_1552);
and U1358 (N_1358,In_1810,In_44);
or U1359 (N_1359,In_436,In_1753);
nand U1360 (N_1360,In_348,In_742);
or U1361 (N_1361,In_433,In_1844);
nand U1362 (N_1362,In_1531,In_625);
xor U1363 (N_1363,In_750,In_872);
or U1364 (N_1364,In_240,In_742);
nor U1365 (N_1365,In_1961,In_473);
nand U1366 (N_1366,In_1418,In_1162);
nand U1367 (N_1367,In_885,In_737);
nor U1368 (N_1368,In_1192,In_1443);
nor U1369 (N_1369,In_1262,In_261);
nand U1370 (N_1370,In_506,In_504);
and U1371 (N_1371,In_1659,In_4);
or U1372 (N_1372,In_1052,In_891);
xor U1373 (N_1373,In_1600,In_257);
or U1374 (N_1374,In_888,In_913);
nand U1375 (N_1375,In_424,In_473);
and U1376 (N_1376,In_16,In_1930);
nand U1377 (N_1377,In_1059,In_1237);
xnor U1378 (N_1378,In_611,In_720);
nor U1379 (N_1379,In_244,In_979);
xnor U1380 (N_1380,In_1850,In_1422);
nor U1381 (N_1381,In_1724,In_1968);
and U1382 (N_1382,In_160,In_1194);
or U1383 (N_1383,In_1162,In_421);
nor U1384 (N_1384,In_228,In_1627);
nor U1385 (N_1385,In_1898,In_757);
xor U1386 (N_1386,In_206,In_307);
xor U1387 (N_1387,In_1405,In_910);
xor U1388 (N_1388,In_1203,In_620);
and U1389 (N_1389,In_1200,In_1006);
and U1390 (N_1390,In_624,In_255);
nor U1391 (N_1391,In_1273,In_913);
and U1392 (N_1392,In_734,In_1598);
nor U1393 (N_1393,In_255,In_1188);
or U1394 (N_1394,In_447,In_1905);
xor U1395 (N_1395,In_20,In_1073);
and U1396 (N_1396,In_576,In_1130);
and U1397 (N_1397,In_8,In_1406);
or U1398 (N_1398,In_58,In_686);
or U1399 (N_1399,In_276,In_148);
and U1400 (N_1400,In_1891,In_778);
nor U1401 (N_1401,In_1267,In_1229);
xnor U1402 (N_1402,In_447,In_1821);
nand U1403 (N_1403,In_872,In_631);
or U1404 (N_1404,In_1286,In_96);
and U1405 (N_1405,In_1789,In_462);
xor U1406 (N_1406,In_1502,In_1811);
nand U1407 (N_1407,In_940,In_1225);
or U1408 (N_1408,In_1051,In_1353);
or U1409 (N_1409,In_1308,In_54);
or U1410 (N_1410,In_954,In_875);
or U1411 (N_1411,In_1724,In_1222);
or U1412 (N_1412,In_1856,In_1960);
or U1413 (N_1413,In_1283,In_1116);
xnor U1414 (N_1414,In_1052,In_920);
xor U1415 (N_1415,In_232,In_1153);
xor U1416 (N_1416,In_925,In_1116);
xor U1417 (N_1417,In_1966,In_1678);
and U1418 (N_1418,In_826,In_1979);
nand U1419 (N_1419,In_1690,In_479);
xnor U1420 (N_1420,In_720,In_843);
and U1421 (N_1421,In_1275,In_518);
and U1422 (N_1422,In_223,In_877);
nor U1423 (N_1423,In_787,In_1007);
and U1424 (N_1424,In_1841,In_1696);
and U1425 (N_1425,In_861,In_1244);
and U1426 (N_1426,In_1544,In_1284);
xor U1427 (N_1427,In_1037,In_784);
or U1428 (N_1428,In_1495,In_856);
or U1429 (N_1429,In_629,In_543);
and U1430 (N_1430,In_369,In_628);
and U1431 (N_1431,In_379,In_116);
xnor U1432 (N_1432,In_102,In_4);
nand U1433 (N_1433,In_111,In_763);
nand U1434 (N_1434,In_2,In_1150);
xnor U1435 (N_1435,In_254,In_1469);
xnor U1436 (N_1436,In_1937,In_1886);
and U1437 (N_1437,In_1633,In_1920);
nand U1438 (N_1438,In_1957,In_912);
or U1439 (N_1439,In_871,In_1588);
and U1440 (N_1440,In_112,In_63);
or U1441 (N_1441,In_89,In_1450);
nor U1442 (N_1442,In_1288,In_1952);
nand U1443 (N_1443,In_753,In_489);
nor U1444 (N_1444,In_298,In_1343);
nor U1445 (N_1445,In_515,In_297);
and U1446 (N_1446,In_390,In_1580);
xor U1447 (N_1447,In_1762,In_1924);
or U1448 (N_1448,In_240,In_1970);
or U1449 (N_1449,In_646,In_1556);
nor U1450 (N_1450,In_1802,In_744);
nor U1451 (N_1451,In_1500,In_1249);
nand U1452 (N_1452,In_471,In_1141);
xor U1453 (N_1453,In_1338,In_1080);
nor U1454 (N_1454,In_829,In_184);
nand U1455 (N_1455,In_1002,In_523);
nand U1456 (N_1456,In_1702,In_1983);
xnor U1457 (N_1457,In_84,In_100);
xor U1458 (N_1458,In_1221,In_229);
xnor U1459 (N_1459,In_1165,In_988);
or U1460 (N_1460,In_753,In_1734);
or U1461 (N_1461,In_1123,In_1095);
nand U1462 (N_1462,In_821,In_1280);
nor U1463 (N_1463,In_295,In_47);
nand U1464 (N_1464,In_1752,In_1867);
xor U1465 (N_1465,In_1011,In_557);
nand U1466 (N_1466,In_1822,In_946);
or U1467 (N_1467,In_1993,In_1215);
nand U1468 (N_1468,In_1680,In_1245);
or U1469 (N_1469,In_1602,In_1771);
or U1470 (N_1470,In_1929,In_1317);
nand U1471 (N_1471,In_888,In_1635);
xnor U1472 (N_1472,In_349,In_1936);
or U1473 (N_1473,In_215,In_804);
xnor U1474 (N_1474,In_1383,In_771);
nand U1475 (N_1475,In_87,In_456);
and U1476 (N_1476,In_1490,In_701);
xnor U1477 (N_1477,In_987,In_716);
nor U1478 (N_1478,In_310,In_710);
nor U1479 (N_1479,In_1739,In_1031);
nand U1480 (N_1480,In_369,In_1620);
nor U1481 (N_1481,In_1635,In_190);
nand U1482 (N_1482,In_1041,In_1039);
nand U1483 (N_1483,In_1217,In_1354);
nor U1484 (N_1484,In_1837,In_1162);
xnor U1485 (N_1485,In_1238,In_1494);
nor U1486 (N_1486,In_1558,In_1887);
xnor U1487 (N_1487,In_287,In_1860);
or U1488 (N_1488,In_369,In_14);
and U1489 (N_1489,In_1131,In_751);
or U1490 (N_1490,In_218,In_1516);
nand U1491 (N_1491,In_248,In_792);
xnor U1492 (N_1492,In_345,In_214);
nor U1493 (N_1493,In_808,In_925);
nor U1494 (N_1494,In_582,In_1531);
nor U1495 (N_1495,In_780,In_1394);
or U1496 (N_1496,In_1429,In_1674);
nand U1497 (N_1497,In_829,In_1636);
nor U1498 (N_1498,In_1910,In_682);
or U1499 (N_1499,In_608,In_1530);
nand U1500 (N_1500,In_1496,In_1336);
xnor U1501 (N_1501,In_47,In_1914);
nor U1502 (N_1502,In_549,In_1285);
xnor U1503 (N_1503,In_205,In_643);
nor U1504 (N_1504,In_897,In_938);
nand U1505 (N_1505,In_1816,In_1842);
or U1506 (N_1506,In_1620,In_737);
xor U1507 (N_1507,In_688,In_774);
xnor U1508 (N_1508,In_1401,In_1162);
nor U1509 (N_1509,In_1289,In_1121);
xor U1510 (N_1510,In_1346,In_1119);
and U1511 (N_1511,In_1573,In_1772);
nor U1512 (N_1512,In_1253,In_506);
nand U1513 (N_1513,In_211,In_821);
xor U1514 (N_1514,In_1767,In_1506);
nand U1515 (N_1515,In_53,In_302);
or U1516 (N_1516,In_1754,In_1403);
nand U1517 (N_1517,In_1778,In_1619);
xor U1518 (N_1518,In_1589,In_1880);
nor U1519 (N_1519,In_1355,In_273);
xor U1520 (N_1520,In_1281,In_1844);
nand U1521 (N_1521,In_1279,In_186);
nand U1522 (N_1522,In_107,In_1143);
nand U1523 (N_1523,In_645,In_656);
nand U1524 (N_1524,In_1399,In_1308);
nand U1525 (N_1525,In_1984,In_750);
nand U1526 (N_1526,In_1,In_482);
nor U1527 (N_1527,In_391,In_1266);
nor U1528 (N_1528,In_559,In_1599);
nor U1529 (N_1529,In_56,In_957);
or U1530 (N_1530,In_328,In_854);
xor U1531 (N_1531,In_30,In_241);
xor U1532 (N_1532,In_1207,In_1807);
nor U1533 (N_1533,In_1032,In_394);
or U1534 (N_1534,In_1294,In_1479);
or U1535 (N_1535,In_1356,In_490);
nand U1536 (N_1536,In_467,In_998);
nand U1537 (N_1537,In_1281,In_902);
and U1538 (N_1538,In_1490,In_221);
or U1539 (N_1539,In_1692,In_722);
or U1540 (N_1540,In_134,In_1463);
or U1541 (N_1541,In_11,In_1313);
and U1542 (N_1542,In_1359,In_894);
or U1543 (N_1543,In_1145,In_528);
and U1544 (N_1544,In_405,In_1003);
or U1545 (N_1545,In_959,In_1639);
or U1546 (N_1546,In_38,In_287);
xnor U1547 (N_1547,In_1688,In_249);
or U1548 (N_1548,In_810,In_1332);
nor U1549 (N_1549,In_516,In_1796);
and U1550 (N_1550,In_370,In_1950);
xnor U1551 (N_1551,In_279,In_1455);
nand U1552 (N_1552,In_1451,In_221);
nor U1553 (N_1553,In_902,In_968);
nand U1554 (N_1554,In_1880,In_114);
nor U1555 (N_1555,In_327,In_608);
nor U1556 (N_1556,In_1618,In_340);
xor U1557 (N_1557,In_1886,In_72);
nor U1558 (N_1558,In_1229,In_1199);
and U1559 (N_1559,In_1880,In_1788);
nand U1560 (N_1560,In_727,In_147);
nor U1561 (N_1561,In_1289,In_384);
nor U1562 (N_1562,In_1926,In_1123);
nor U1563 (N_1563,In_302,In_964);
nand U1564 (N_1564,In_670,In_490);
nand U1565 (N_1565,In_144,In_1166);
nand U1566 (N_1566,In_194,In_1232);
nand U1567 (N_1567,In_1065,In_1152);
nand U1568 (N_1568,In_1400,In_780);
or U1569 (N_1569,In_460,In_1802);
and U1570 (N_1570,In_1499,In_1871);
nand U1571 (N_1571,In_1084,In_529);
nand U1572 (N_1572,In_167,In_1199);
xnor U1573 (N_1573,In_1684,In_287);
xnor U1574 (N_1574,In_447,In_437);
xnor U1575 (N_1575,In_1201,In_992);
nor U1576 (N_1576,In_1895,In_150);
or U1577 (N_1577,In_321,In_606);
or U1578 (N_1578,In_1963,In_349);
and U1579 (N_1579,In_1882,In_1952);
nor U1580 (N_1580,In_657,In_1103);
or U1581 (N_1581,In_990,In_1354);
nor U1582 (N_1582,In_231,In_1153);
nand U1583 (N_1583,In_340,In_545);
nand U1584 (N_1584,In_63,In_858);
nand U1585 (N_1585,In_1464,In_1302);
or U1586 (N_1586,In_205,In_1223);
and U1587 (N_1587,In_489,In_1964);
xor U1588 (N_1588,In_738,In_1963);
nand U1589 (N_1589,In_1589,In_1912);
and U1590 (N_1590,In_168,In_1010);
xor U1591 (N_1591,In_1553,In_394);
nor U1592 (N_1592,In_1716,In_1959);
nand U1593 (N_1593,In_345,In_1970);
or U1594 (N_1594,In_1231,In_1663);
and U1595 (N_1595,In_74,In_717);
nand U1596 (N_1596,In_1837,In_401);
or U1597 (N_1597,In_840,In_835);
nor U1598 (N_1598,In_200,In_1267);
xor U1599 (N_1599,In_1664,In_1784);
and U1600 (N_1600,In_1442,In_1888);
nor U1601 (N_1601,In_109,In_1619);
nand U1602 (N_1602,In_1439,In_186);
nand U1603 (N_1603,In_535,In_783);
nor U1604 (N_1604,In_1845,In_1005);
nand U1605 (N_1605,In_483,In_641);
nand U1606 (N_1606,In_163,In_1282);
nor U1607 (N_1607,In_1726,In_476);
or U1608 (N_1608,In_833,In_1353);
and U1609 (N_1609,In_565,In_544);
nand U1610 (N_1610,In_129,In_502);
or U1611 (N_1611,In_281,In_1426);
nand U1612 (N_1612,In_1377,In_632);
nand U1613 (N_1613,In_1724,In_1453);
nand U1614 (N_1614,In_1485,In_308);
nor U1615 (N_1615,In_1894,In_893);
and U1616 (N_1616,In_72,In_619);
nor U1617 (N_1617,In_846,In_1143);
nor U1618 (N_1618,In_842,In_1496);
nor U1619 (N_1619,In_965,In_1996);
nor U1620 (N_1620,In_204,In_320);
xnor U1621 (N_1621,In_600,In_307);
nand U1622 (N_1622,In_1925,In_107);
nor U1623 (N_1623,In_1951,In_251);
or U1624 (N_1624,In_1559,In_92);
nand U1625 (N_1625,In_1418,In_1293);
and U1626 (N_1626,In_820,In_736);
and U1627 (N_1627,In_1242,In_1368);
nand U1628 (N_1628,In_776,In_382);
nand U1629 (N_1629,In_15,In_1596);
and U1630 (N_1630,In_1767,In_33);
and U1631 (N_1631,In_1374,In_178);
or U1632 (N_1632,In_1803,In_1358);
and U1633 (N_1633,In_260,In_1527);
and U1634 (N_1634,In_317,In_86);
xor U1635 (N_1635,In_662,In_376);
and U1636 (N_1636,In_1513,In_1569);
or U1637 (N_1637,In_1891,In_55);
nor U1638 (N_1638,In_1625,In_1264);
or U1639 (N_1639,In_1786,In_64);
and U1640 (N_1640,In_276,In_1977);
or U1641 (N_1641,In_1203,In_1010);
and U1642 (N_1642,In_1356,In_356);
nand U1643 (N_1643,In_1263,In_774);
nor U1644 (N_1644,In_812,In_495);
and U1645 (N_1645,In_460,In_469);
and U1646 (N_1646,In_1879,In_1885);
xor U1647 (N_1647,In_1993,In_30);
nand U1648 (N_1648,In_1166,In_724);
and U1649 (N_1649,In_1786,In_1276);
or U1650 (N_1650,In_837,In_817);
xnor U1651 (N_1651,In_120,In_463);
xnor U1652 (N_1652,In_302,In_315);
nor U1653 (N_1653,In_215,In_972);
nor U1654 (N_1654,In_1084,In_1043);
xor U1655 (N_1655,In_1677,In_1288);
and U1656 (N_1656,In_225,In_1984);
nor U1657 (N_1657,In_684,In_1222);
nand U1658 (N_1658,In_1843,In_634);
nor U1659 (N_1659,In_392,In_291);
and U1660 (N_1660,In_1639,In_215);
xor U1661 (N_1661,In_113,In_1233);
or U1662 (N_1662,In_1754,In_1334);
nand U1663 (N_1663,In_1175,In_1657);
and U1664 (N_1664,In_750,In_781);
and U1665 (N_1665,In_954,In_1923);
and U1666 (N_1666,In_274,In_1636);
or U1667 (N_1667,In_1574,In_1739);
nor U1668 (N_1668,In_1584,In_1315);
nor U1669 (N_1669,In_1067,In_992);
or U1670 (N_1670,In_552,In_173);
nor U1671 (N_1671,In_846,In_723);
or U1672 (N_1672,In_1541,In_233);
nor U1673 (N_1673,In_77,In_1388);
nor U1674 (N_1674,In_1161,In_1798);
xor U1675 (N_1675,In_1617,In_582);
nand U1676 (N_1676,In_719,In_1769);
or U1677 (N_1677,In_1369,In_399);
and U1678 (N_1678,In_324,In_1329);
nand U1679 (N_1679,In_88,In_1231);
or U1680 (N_1680,In_1436,In_1428);
or U1681 (N_1681,In_1481,In_134);
xnor U1682 (N_1682,In_1473,In_407);
or U1683 (N_1683,In_711,In_732);
and U1684 (N_1684,In_1072,In_822);
xor U1685 (N_1685,In_1217,In_270);
and U1686 (N_1686,In_620,In_1624);
xnor U1687 (N_1687,In_770,In_906);
or U1688 (N_1688,In_1858,In_568);
nand U1689 (N_1689,In_1549,In_1971);
xnor U1690 (N_1690,In_1617,In_701);
or U1691 (N_1691,In_31,In_1992);
nand U1692 (N_1692,In_1883,In_1425);
xnor U1693 (N_1693,In_10,In_1189);
or U1694 (N_1694,In_1753,In_1431);
nand U1695 (N_1695,In_426,In_1060);
xnor U1696 (N_1696,In_1228,In_140);
or U1697 (N_1697,In_1221,In_1538);
nand U1698 (N_1698,In_959,In_1694);
xor U1699 (N_1699,In_1293,In_1496);
xor U1700 (N_1700,In_1154,In_75);
and U1701 (N_1701,In_1486,In_357);
xnor U1702 (N_1702,In_319,In_1011);
or U1703 (N_1703,In_1316,In_471);
and U1704 (N_1704,In_230,In_1663);
or U1705 (N_1705,In_683,In_465);
xor U1706 (N_1706,In_1529,In_1615);
or U1707 (N_1707,In_1556,In_1531);
or U1708 (N_1708,In_274,In_280);
nand U1709 (N_1709,In_657,In_344);
and U1710 (N_1710,In_701,In_1043);
nor U1711 (N_1711,In_421,In_707);
xnor U1712 (N_1712,In_1823,In_1173);
and U1713 (N_1713,In_537,In_965);
nand U1714 (N_1714,In_910,In_230);
and U1715 (N_1715,In_1589,In_1294);
nor U1716 (N_1716,In_289,In_1663);
xnor U1717 (N_1717,In_224,In_1879);
xor U1718 (N_1718,In_1860,In_339);
and U1719 (N_1719,In_1928,In_777);
nand U1720 (N_1720,In_74,In_1151);
and U1721 (N_1721,In_1176,In_115);
and U1722 (N_1722,In_261,In_1867);
or U1723 (N_1723,In_941,In_1288);
xor U1724 (N_1724,In_446,In_1771);
nand U1725 (N_1725,In_1645,In_439);
and U1726 (N_1726,In_283,In_818);
and U1727 (N_1727,In_1993,In_824);
nor U1728 (N_1728,In_694,In_120);
nor U1729 (N_1729,In_1432,In_1763);
and U1730 (N_1730,In_1810,In_1834);
or U1731 (N_1731,In_1254,In_443);
and U1732 (N_1732,In_490,In_82);
xnor U1733 (N_1733,In_1893,In_1019);
nor U1734 (N_1734,In_1576,In_1727);
nand U1735 (N_1735,In_1652,In_671);
or U1736 (N_1736,In_1337,In_772);
nand U1737 (N_1737,In_1516,In_1709);
xnor U1738 (N_1738,In_45,In_281);
xnor U1739 (N_1739,In_1533,In_1103);
nor U1740 (N_1740,In_1676,In_875);
or U1741 (N_1741,In_1810,In_1177);
or U1742 (N_1742,In_1342,In_1675);
or U1743 (N_1743,In_538,In_1828);
nor U1744 (N_1744,In_1207,In_685);
and U1745 (N_1745,In_199,In_1989);
nand U1746 (N_1746,In_15,In_803);
nor U1747 (N_1747,In_1522,In_510);
and U1748 (N_1748,In_1267,In_1647);
or U1749 (N_1749,In_383,In_1211);
xnor U1750 (N_1750,In_1491,In_1567);
nand U1751 (N_1751,In_170,In_985);
nor U1752 (N_1752,In_177,In_1151);
or U1753 (N_1753,In_890,In_1687);
nor U1754 (N_1754,In_1365,In_1498);
nor U1755 (N_1755,In_1425,In_1737);
or U1756 (N_1756,In_150,In_965);
nand U1757 (N_1757,In_775,In_340);
xnor U1758 (N_1758,In_1896,In_1546);
nand U1759 (N_1759,In_910,In_1916);
or U1760 (N_1760,In_189,In_1452);
or U1761 (N_1761,In_1635,In_1288);
or U1762 (N_1762,In_1207,In_1469);
or U1763 (N_1763,In_510,In_1810);
nand U1764 (N_1764,In_221,In_808);
xor U1765 (N_1765,In_1299,In_1101);
nor U1766 (N_1766,In_1018,In_1405);
nand U1767 (N_1767,In_409,In_583);
nor U1768 (N_1768,In_58,In_1487);
or U1769 (N_1769,In_1423,In_1898);
nor U1770 (N_1770,In_1980,In_1092);
nor U1771 (N_1771,In_1149,In_1354);
nand U1772 (N_1772,In_422,In_515);
and U1773 (N_1773,In_700,In_1539);
or U1774 (N_1774,In_92,In_759);
nand U1775 (N_1775,In_1070,In_848);
nand U1776 (N_1776,In_1672,In_1417);
nor U1777 (N_1777,In_1508,In_1498);
or U1778 (N_1778,In_948,In_626);
nor U1779 (N_1779,In_1614,In_1013);
and U1780 (N_1780,In_1828,In_1247);
nand U1781 (N_1781,In_1863,In_1569);
xor U1782 (N_1782,In_1278,In_486);
xor U1783 (N_1783,In_320,In_1481);
nand U1784 (N_1784,In_1656,In_1766);
xnor U1785 (N_1785,In_1741,In_1071);
and U1786 (N_1786,In_1106,In_846);
and U1787 (N_1787,In_1523,In_1245);
and U1788 (N_1788,In_1756,In_587);
and U1789 (N_1789,In_1662,In_1831);
and U1790 (N_1790,In_123,In_28);
nor U1791 (N_1791,In_802,In_1941);
and U1792 (N_1792,In_811,In_813);
or U1793 (N_1793,In_1082,In_290);
and U1794 (N_1794,In_1242,In_1889);
or U1795 (N_1795,In_201,In_1536);
and U1796 (N_1796,In_229,In_275);
nand U1797 (N_1797,In_1375,In_872);
nand U1798 (N_1798,In_1404,In_1823);
or U1799 (N_1799,In_463,In_108);
and U1800 (N_1800,In_1115,In_887);
or U1801 (N_1801,In_1965,In_1571);
nor U1802 (N_1802,In_40,In_944);
and U1803 (N_1803,In_640,In_419);
xor U1804 (N_1804,In_463,In_1277);
nor U1805 (N_1805,In_1576,In_155);
xnor U1806 (N_1806,In_1156,In_1158);
nand U1807 (N_1807,In_387,In_111);
xnor U1808 (N_1808,In_1875,In_1102);
nor U1809 (N_1809,In_1550,In_101);
xnor U1810 (N_1810,In_1907,In_1940);
and U1811 (N_1811,In_874,In_589);
and U1812 (N_1812,In_1408,In_487);
xor U1813 (N_1813,In_1616,In_1064);
or U1814 (N_1814,In_942,In_621);
xor U1815 (N_1815,In_700,In_945);
and U1816 (N_1816,In_1117,In_127);
nand U1817 (N_1817,In_1105,In_87);
nor U1818 (N_1818,In_1002,In_1442);
xnor U1819 (N_1819,In_162,In_1108);
nor U1820 (N_1820,In_718,In_1367);
xnor U1821 (N_1821,In_319,In_1481);
xor U1822 (N_1822,In_750,In_15);
nand U1823 (N_1823,In_119,In_421);
nand U1824 (N_1824,In_519,In_1066);
and U1825 (N_1825,In_212,In_748);
and U1826 (N_1826,In_1120,In_1943);
xor U1827 (N_1827,In_1271,In_785);
or U1828 (N_1828,In_1692,In_427);
nor U1829 (N_1829,In_904,In_57);
or U1830 (N_1830,In_109,In_702);
nand U1831 (N_1831,In_1077,In_523);
or U1832 (N_1832,In_144,In_304);
nand U1833 (N_1833,In_1798,In_698);
nand U1834 (N_1834,In_1468,In_427);
or U1835 (N_1835,In_1053,In_1774);
xnor U1836 (N_1836,In_453,In_1891);
or U1837 (N_1837,In_1275,In_1039);
nor U1838 (N_1838,In_1795,In_1624);
xnor U1839 (N_1839,In_1280,In_1687);
nand U1840 (N_1840,In_141,In_1694);
xor U1841 (N_1841,In_1155,In_207);
xor U1842 (N_1842,In_1460,In_1262);
xor U1843 (N_1843,In_542,In_1330);
or U1844 (N_1844,In_1667,In_259);
nand U1845 (N_1845,In_589,In_1101);
nand U1846 (N_1846,In_899,In_694);
nand U1847 (N_1847,In_1556,In_425);
nor U1848 (N_1848,In_428,In_299);
xnor U1849 (N_1849,In_892,In_621);
or U1850 (N_1850,In_1368,In_354);
and U1851 (N_1851,In_596,In_395);
nand U1852 (N_1852,In_1384,In_1377);
nor U1853 (N_1853,In_763,In_635);
nand U1854 (N_1854,In_1235,In_125);
and U1855 (N_1855,In_1826,In_531);
nor U1856 (N_1856,In_821,In_1884);
or U1857 (N_1857,In_1654,In_1847);
and U1858 (N_1858,In_1661,In_1423);
nand U1859 (N_1859,In_1590,In_556);
xor U1860 (N_1860,In_219,In_1115);
or U1861 (N_1861,In_857,In_877);
xor U1862 (N_1862,In_4,In_1796);
or U1863 (N_1863,In_718,In_419);
xnor U1864 (N_1864,In_1334,In_1985);
or U1865 (N_1865,In_1118,In_1207);
xor U1866 (N_1866,In_1043,In_1224);
nand U1867 (N_1867,In_1327,In_1867);
xnor U1868 (N_1868,In_1819,In_1980);
nand U1869 (N_1869,In_1724,In_688);
or U1870 (N_1870,In_666,In_1296);
nand U1871 (N_1871,In_1679,In_1817);
nor U1872 (N_1872,In_1268,In_1611);
or U1873 (N_1873,In_493,In_377);
nand U1874 (N_1874,In_292,In_1710);
xor U1875 (N_1875,In_740,In_489);
xor U1876 (N_1876,In_781,In_497);
or U1877 (N_1877,In_293,In_1512);
and U1878 (N_1878,In_1807,In_1441);
nor U1879 (N_1879,In_125,In_1430);
and U1880 (N_1880,In_1244,In_268);
nor U1881 (N_1881,In_234,In_1100);
xor U1882 (N_1882,In_219,In_378);
nand U1883 (N_1883,In_137,In_1505);
xnor U1884 (N_1884,In_1961,In_770);
and U1885 (N_1885,In_666,In_246);
or U1886 (N_1886,In_963,In_36);
xnor U1887 (N_1887,In_350,In_1927);
xnor U1888 (N_1888,In_794,In_820);
or U1889 (N_1889,In_304,In_415);
nor U1890 (N_1890,In_1555,In_1094);
or U1891 (N_1891,In_13,In_1221);
or U1892 (N_1892,In_1298,In_1773);
and U1893 (N_1893,In_1015,In_59);
xnor U1894 (N_1894,In_1086,In_814);
and U1895 (N_1895,In_762,In_474);
xor U1896 (N_1896,In_1365,In_640);
nor U1897 (N_1897,In_1021,In_133);
or U1898 (N_1898,In_1588,In_1238);
nand U1899 (N_1899,In_917,In_900);
or U1900 (N_1900,In_92,In_749);
xor U1901 (N_1901,In_643,In_1346);
nor U1902 (N_1902,In_356,In_747);
and U1903 (N_1903,In_1625,In_242);
and U1904 (N_1904,In_0,In_1609);
xnor U1905 (N_1905,In_778,In_1344);
xnor U1906 (N_1906,In_184,In_1058);
xor U1907 (N_1907,In_1975,In_514);
and U1908 (N_1908,In_953,In_162);
and U1909 (N_1909,In_1362,In_1260);
and U1910 (N_1910,In_1066,In_1806);
and U1911 (N_1911,In_1997,In_1198);
xor U1912 (N_1912,In_1383,In_1180);
xor U1913 (N_1913,In_7,In_150);
xor U1914 (N_1914,In_1555,In_431);
or U1915 (N_1915,In_1952,In_1060);
nand U1916 (N_1916,In_1643,In_1406);
nand U1917 (N_1917,In_237,In_1118);
and U1918 (N_1918,In_1278,In_1970);
nand U1919 (N_1919,In_1557,In_655);
nand U1920 (N_1920,In_653,In_1889);
and U1921 (N_1921,In_869,In_739);
nand U1922 (N_1922,In_623,In_1288);
or U1923 (N_1923,In_412,In_1078);
or U1924 (N_1924,In_593,In_961);
xor U1925 (N_1925,In_426,In_566);
and U1926 (N_1926,In_1596,In_1262);
nand U1927 (N_1927,In_1626,In_1237);
or U1928 (N_1928,In_562,In_1201);
xnor U1929 (N_1929,In_1499,In_1362);
and U1930 (N_1930,In_1906,In_777);
xnor U1931 (N_1931,In_1191,In_142);
nor U1932 (N_1932,In_1751,In_82);
or U1933 (N_1933,In_1588,In_915);
nor U1934 (N_1934,In_1726,In_1412);
nand U1935 (N_1935,In_1876,In_731);
or U1936 (N_1936,In_948,In_321);
nand U1937 (N_1937,In_1493,In_396);
nor U1938 (N_1938,In_13,In_1887);
xor U1939 (N_1939,In_1796,In_550);
nor U1940 (N_1940,In_593,In_1461);
nor U1941 (N_1941,In_1136,In_510);
or U1942 (N_1942,In_1937,In_1255);
xor U1943 (N_1943,In_793,In_1185);
and U1944 (N_1944,In_300,In_1601);
and U1945 (N_1945,In_1055,In_915);
nand U1946 (N_1946,In_381,In_130);
xnor U1947 (N_1947,In_1453,In_602);
nor U1948 (N_1948,In_708,In_224);
or U1949 (N_1949,In_936,In_1371);
and U1950 (N_1950,In_557,In_44);
and U1951 (N_1951,In_183,In_1020);
and U1952 (N_1952,In_1314,In_708);
and U1953 (N_1953,In_364,In_836);
nand U1954 (N_1954,In_1776,In_1083);
and U1955 (N_1955,In_1716,In_291);
and U1956 (N_1956,In_1275,In_1072);
xor U1957 (N_1957,In_1657,In_1300);
xnor U1958 (N_1958,In_421,In_996);
nor U1959 (N_1959,In_780,In_433);
nand U1960 (N_1960,In_1320,In_979);
nor U1961 (N_1961,In_562,In_343);
nor U1962 (N_1962,In_1804,In_135);
or U1963 (N_1963,In_1108,In_1947);
and U1964 (N_1964,In_173,In_676);
or U1965 (N_1965,In_1850,In_1417);
or U1966 (N_1966,In_1796,In_1591);
nor U1967 (N_1967,In_1934,In_383);
and U1968 (N_1968,In_1003,In_1036);
xnor U1969 (N_1969,In_1877,In_470);
nand U1970 (N_1970,In_1305,In_1938);
nor U1971 (N_1971,In_1136,In_388);
nor U1972 (N_1972,In_33,In_1899);
xor U1973 (N_1973,In_1069,In_737);
and U1974 (N_1974,In_160,In_1802);
or U1975 (N_1975,In_895,In_1079);
and U1976 (N_1976,In_1085,In_861);
xor U1977 (N_1977,In_147,In_194);
and U1978 (N_1978,In_1862,In_281);
or U1979 (N_1979,In_853,In_159);
nor U1980 (N_1980,In_676,In_1046);
xor U1981 (N_1981,In_754,In_560);
and U1982 (N_1982,In_351,In_1979);
or U1983 (N_1983,In_1671,In_157);
and U1984 (N_1984,In_1781,In_1085);
and U1985 (N_1985,In_846,In_1438);
and U1986 (N_1986,In_1702,In_1999);
xor U1987 (N_1987,In_596,In_75);
and U1988 (N_1988,In_1763,In_673);
or U1989 (N_1989,In_1273,In_1753);
or U1990 (N_1990,In_1255,In_1544);
nand U1991 (N_1991,In_65,In_1038);
nor U1992 (N_1992,In_1453,In_1929);
or U1993 (N_1993,In_201,In_1949);
nand U1994 (N_1994,In_791,In_743);
nor U1995 (N_1995,In_733,In_168);
nand U1996 (N_1996,In_789,In_598);
or U1997 (N_1997,In_711,In_150);
and U1998 (N_1998,In_1464,In_1724);
or U1999 (N_1999,In_1022,In_1634);
and U2000 (N_2000,In_1274,In_706);
nor U2001 (N_2001,In_559,In_1293);
and U2002 (N_2002,In_765,In_1096);
or U2003 (N_2003,In_938,In_749);
or U2004 (N_2004,In_1868,In_1624);
nor U2005 (N_2005,In_1497,In_981);
and U2006 (N_2006,In_425,In_1599);
or U2007 (N_2007,In_73,In_1269);
nand U2008 (N_2008,In_1405,In_1572);
and U2009 (N_2009,In_1926,In_318);
and U2010 (N_2010,In_1702,In_1841);
nor U2011 (N_2011,In_17,In_1605);
and U2012 (N_2012,In_1046,In_456);
and U2013 (N_2013,In_1729,In_980);
or U2014 (N_2014,In_61,In_432);
xnor U2015 (N_2015,In_1058,In_1786);
nor U2016 (N_2016,In_608,In_1971);
or U2017 (N_2017,In_1550,In_1596);
nor U2018 (N_2018,In_754,In_1890);
xor U2019 (N_2019,In_298,In_704);
nor U2020 (N_2020,In_1465,In_1223);
nand U2021 (N_2021,In_1778,In_1772);
nand U2022 (N_2022,In_1080,In_291);
xnor U2023 (N_2023,In_543,In_739);
xnor U2024 (N_2024,In_903,In_285);
xor U2025 (N_2025,In_204,In_1052);
nand U2026 (N_2026,In_55,In_1503);
or U2027 (N_2027,In_448,In_107);
or U2028 (N_2028,In_911,In_1197);
xnor U2029 (N_2029,In_826,In_1664);
nor U2030 (N_2030,In_92,In_751);
or U2031 (N_2031,In_1573,In_1405);
nand U2032 (N_2032,In_1655,In_1967);
xnor U2033 (N_2033,In_1701,In_259);
and U2034 (N_2034,In_1266,In_1312);
or U2035 (N_2035,In_699,In_1193);
nor U2036 (N_2036,In_210,In_165);
nand U2037 (N_2037,In_584,In_1050);
xor U2038 (N_2038,In_1404,In_1422);
and U2039 (N_2039,In_1813,In_1280);
or U2040 (N_2040,In_1573,In_1329);
xnor U2041 (N_2041,In_414,In_159);
and U2042 (N_2042,In_617,In_1625);
nor U2043 (N_2043,In_1514,In_34);
or U2044 (N_2044,In_1147,In_1381);
and U2045 (N_2045,In_1359,In_1722);
or U2046 (N_2046,In_1278,In_609);
xnor U2047 (N_2047,In_1104,In_1963);
and U2048 (N_2048,In_465,In_470);
or U2049 (N_2049,In_1827,In_115);
and U2050 (N_2050,In_606,In_1915);
nor U2051 (N_2051,In_1772,In_665);
nor U2052 (N_2052,In_800,In_921);
xor U2053 (N_2053,In_368,In_1229);
nand U2054 (N_2054,In_1418,In_1669);
and U2055 (N_2055,In_1399,In_101);
or U2056 (N_2056,In_723,In_807);
xor U2057 (N_2057,In_1042,In_1211);
and U2058 (N_2058,In_1815,In_1818);
or U2059 (N_2059,In_1464,In_1141);
nand U2060 (N_2060,In_1316,In_1756);
and U2061 (N_2061,In_781,In_1133);
or U2062 (N_2062,In_926,In_586);
or U2063 (N_2063,In_953,In_1778);
and U2064 (N_2064,In_1167,In_841);
nand U2065 (N_2065,In_1778,In_206);
nor U2066 (N_2066,In_882,In_1248);
or U2067 (N_2067,In_1107,In_772);
xor U2068 (N_2068,In_1408,In_105);
nand U2069 (N_2069,In_1878,In_1294);
nor U2070 (N_2070,In_105,In_1636);
or U2071 (N_2071,In_1960,In_121);
and U2072 (N_2072,In_1069,In_706);
nand U2073 (N_2073,In_1387,In_1189);
or U2074 (N_2074,In_1347,In_645);
xnor U2075 (N_2075,In_191,In_1973);
or U2076 (N_2076,In_1212,In_1717);
nor U2077 (N_2077,In_230,In_1529);
nor U2078 (N_2078,In_1840,In_420);
or U2079 (N_2079,In_111,In_1348);
and U2080 (N_2080,In_1702,In_1036);
nor U2081 (N_2081,In_445,In_24);
and U2082 (N_2082,In_1217,In_1703);
xor U2083 (N_2083,In_664,In_546);
nand U2084 (N_2084,In_834,In_89);
and U2085 (N_2085,In_988,In_1981);
xor U2086 (N_2086,In_676,In_1328);
nand U2087 (N_2087,In_316,In_1559);
or U2088 (N_2088,In_1409,In_562);
and U2089 (N_2089,In_514,In_1119);
nor U2090 (N_2090,In_1404,In_191);
and U2091 (N_2091,In_756,In_1840);
and U2092 (N_2092,In_922,In_1628);
nor U2093 (N_2093,In_1754,In_1286);
and U2094 (N_2094,In_159,In_1557);
nand U2095 (N_2095,In_437,In_651);
xor U2096 (N_2096,In_1645,In_586);
nor U2097 (N_2097,In_1161,In_45);
and U2098 (N_2098,In_1178,In_1535);
or U2099 (N_2099,In_156,In_867);
xor U2100 (N_2100,In_1714,In_1247);
and U2101 (N_2101,In_384,In_1285);
xnor U2102 (N_2102,In_1454,In_1582);
nor U2103 (N_2103,In_1262,In_277);
or U2104 (N_2104,In_1684,In_1047);
nand U2105 (N_2105,In_1929,In_1823);
nor U2106 (N_2106,In_335,In_126);
xor U2107 (N_2107,In_1877,In_1521);
nand U2108 (N_2108,In_1041,In_1712);
and U2109 (N_2109,In_1438,In_869);
nor U2110 (N_2110,In_1640,In_920);
nor U2111 (N_2111,In_823,In_1584);
and U2112 (N_2112,In_1660,In_603);
nor U2113 (N_2113,In_1958,In_891);
nor U2114 (N_2114,In_1588,In_596);
or U2115 (N_2115,In_437,In_773);
and U2116 (N_2116,In_751,In_1289);
and U2117 (N_2117,In_1874,In_613);
nor U2118 (N_2118,In_1448,In_793);
xor U2119 (N_2119,In_566,In_1598);
and U2120 (N_2120,In_1594,In_806);
nor U2121 (N_2121,In_56,In_1235);
nand U2122 (N_2122,In_919,In_1084);
nand U2123 (N_2123,In_1641,In_1066);
nand U2124 (N_2124,In_1043,In_1524);
xor U2125 (N_2125,In_1574,In_267);
nor U2126 (N_2126,In_1182,In_3);
nor U2127 (N_2127,In_94,In_71);
nor U2128 (N_2128,In_381,In_314);
and U2129 (N_2129,In_1643,In_1002);
or U2130 (N_2130,In_1660,In_1929);
nand U2131 (N_2131,In_324,In_1791);
xnor U2132 (N_2132,In_485,In_1886);
and U2133 (N_2133,In_183,In_1819);
xor U2134 (N_2134,In_1179,In_1482);
or U2135 (N_2135,In_1051,In_1378);
xnor U2136 (N_2136,In_194,In_629);
and U2137 (N_2137,In_1830,In_1556);
nand U2138 (N_2138,In_104,In_1737);
or U2139 (N_2139,In_1025,In_129);
nand U2140 (N_2140,In_865,In_311);
or U2141 (N_2141,In_542,In_67);
or U2142 (N_2142,In_949,In_130);
xor U2143 (N_2143,In_536,In_497);
and U2144 (N_2144,In_1950,In_1033);
and U2145 (N_2145,In_1641,In_972);
and U2146 (N_2146,In_163,In_790);
and U2147 (N_2147,In_1373,In_705);
xor U2148 (N_2148,In_1459,In_223);
xnor U2149 (N_2149,In_1520,In_20);
nor U2150 (N_2150,In_667,In_248);
xor U2151 (N_2151,In_1858,In_1250);
nand U2152 (N_2152,In_1004,In_789);
nand U2153 (N_2153,In_712,In_1475);
xor U2154 (N_2154,In_1880,In_952);
nand U2155 (N_2155,In_1830,In_580);
and U2156 (N_2156,In_574,In_15);
xor U2157 (N_2157,In_147,In_199);
or U2158 (N_2158,In_397,In_1719);
nand U2159 (N_2159,In_1559,In_1634);
nand U2160 (N_2160,In_1228,In_465);
xor U2161 (N_2161,In_702,In_409);
xnor U2162 (N_2162,In_253,In_1782);
and U2163 (N_2163,In_1982,In_1301);
or U2164 (N_2164,In_427,In_486);
nand U2165 (N_2165,In_1511,In_1291);
and U2166 (N_2166,In_540,In_508);
nor U2167 (N_2167,In_1904,In_740);
or U2168 (N_2168,In_1598,In_957);
and U2169 (N_2169,In_239,In_1541);
or U2170 (N_2170,In_1768,In_884);
nor U2171 (N_2171,In_1931,In_700);
nand U2172 (N_2172,In_610,In_1954);
and U2173 (N_2173,In_1108,In_1021);
nand U2174 (N_2174,In_1985,In_969);
nor U2175 (N_2175,In_1197,In_981);
xor U2176 (N_2176,In_1180,In_692);
or U2177 (N_2177,In_490,In_576);
xor U2178 (N_2178,In_795,In_1642);
nor U2179 (N_2179,In_1630,In_7);
xnor U2180 (N_2180,In_1157,In_597);
nor U2181 (N_2181,In_587,In_1661);
nor U2182 (N_2182,In_185,In_1115);
nand U2183 (N_2183,In_1770,In_701);
xnor U2184 (N_2184,In_979,In_472);
xnor U2185 (N_2185,In_1072,In_1769);
nor U2186 (N_2186,In_488,In_852);
and U2187 (N_2187,In_1278,In_983);
xor U2188 (N_2188,In_1263,In_64);
or U2189 (N_2189,In_1125,In_1815);
nor U2190 (N_2190,In_1738,In_350);
or U2191 (N_2191,In_1134,In_1324);
or U2192 (N_2192,In_1262,In_1461);
nor U2193 (N_2193,In_260,In_153);
nor U2194 (N_2194,In_1426,In_286);
nor U2195 (N_2195,In_400,In_970);
nor U2196 (N_2196,In_149,In_743);
and U2197 (N_2197,In_1779,In_595);
and U2198 (N_2198,In_275,In_993);
or U2199 (N_2199,In_1402,In_460);
or U2200 (N_2200,In_592,In_133);
nand U2201 (N_2201,In_1437,In_1440);
or U2202 (N_2202,In_444,In_1840);
xor U2203 (N_2203,In_221,In_24);
xnor U2204 (N_2204,In_775,In_1086);
xnor U2205 (N_2205,In_729,In_30);
nor U2206 (N_2206,In_1206,In_14);
or U2207 (N_2207,In_1768,In_1995);
nand U2208 (N_2208,In_1502,In_442);
and U2209 (N_2209,In_1005,In_1846);
xor U2210 (N_2210,In_1605,In_1995);
xnor U2211 (N_2211,In_175,In_1885);
or U2212 (N_2212,In_1181,In_1542);
nor U2213 (N_2213,In_346,In_820);
nand U2214 (N_2214,In_1813,In_721);
or U2215 (N_2215,In_414,In_790);
xor U2216 (N_2216,In_900,In_651);
or U2217 (N_2217,In_1243,In_1279);
nand U2218 (N_2218,In_1660,In_475);
and U2219 (N_2219,In_803,In_1601);
nand U2220 (N_2220,In_169,In_559);
or U2221 (N_2221,In_1609,In_407);
nand U2222 (N_2222,In_1021,In_1222);
nor U2223 (N_2223,In_388,In_1709);
nor U2224 (N_2224,In_99,In_1032);
or U2225 (N_2225,In_1112,In_1851);
xor U2226 (N_2226,In_1101,In_1525);
nand U2227 (N_2227,In_54,In_359);
nand U2228 (N_2228,In_633,In_386);
and U2229 (N_2229,In_767,In_173);
or U2230 (N_2230,In_836,In_1483);
or U2231 (N_2231,In_1242,In_659);
xor U2232 (N_2232,In_965,In_770);
xor U2233 (N_2233,In_1589,In_353);
or U2234 (N_2234,In_1715,In_103);
xor U2235 (N_2235,In_1548,In_309);
or U2236 (N_2236,In_1924,In_937);
nand U2237 (N_2237,In_126,In_547);
nand U2238 (N_2238,In_868,In_176);
xor U2239 (N_2239,In_615,In_1100);
nor U2240 (N_2240,In_681,In_575);
or U2241 (N_2241,In_1357,In_434);
and U2242 (N_2242,In_1187,In_24);
xor U2243 (N_2243,In_540,In_1132);
and U2244 (N_2244,In_1033,In_451);
nor U2245 (N_2245,In_1206,In_1794);
nand U2246 (N_2246,In_311,In_995);
nor U2247 (N_2247,In_975,In_1595);
and U2248 (N_2248,In_637,In_1147);
or U2249 (N_2249,In_179,In_1112);
xor U2250 (N_2250,In_129,In_625);
nand U2251 (N_2251,In_232,In_778);
nand U2252 (N_2252,In_1573,In_375);
xnor U2253 (N_2253,In_1660,In_524);
or U2254 (N_2254,In_828,In_1809);
nor U2255 (N_2255,In_78,In_601);
xor U2256 (N_2256,In_1414,In_241);
or U2257 (N_2257,In_515,In_1165);
or U2258 (N_2258,In_369,In_1688);
and U2259 (N_2259,In_1911,In_1709);
or U2260 (N_2260,In_1714,In_91);
and U2261 (N_2261,In_1851,In_1874);
and U2262 (N_2262,In_960,In_710);
and U2263 (N_2263,In_966,In_866);
or U2264 (N_2264,In_71,In_561);
nand U2265 (N_2265,In_1542,In_1978);
or U2266 (N_2266,In_321,In_1720);
nor U2267 (N_2267,In_847,In_1493);
nor U2268 (N_2268,In_1017,In_1236);
xnor U2269 (N_2269,In_1240,In_1223);
or U2270 (N_2270,In_429,In_860);
nor U2271 (N_2271,In_700,In_1698);
and U2272 (N_2272,In_1568,In_1245);
and U2273 (N_2273,In_20,In_1116);
xnor U2274 (N_2274,In_1510,In_1904);
and U2275 (N_2275,In_232,In_723);
nor U2276 (N_2276,In_1764,In_467);
and U2277 (N_2277,In_821,In_666);
or U2278 (N_2278,In_1843,In_1227);
nand U2279 (N_2279,In_184,In_1998);
nor U2280 (N_2280,In_837,In_1228);
and U2281 (N_2281,In_366,In_678);
nor U2282 (N_2282,In_721,In_271);
nand U2283 (N_2283,In_746,In_765);
and U2284 (N_2284,In_992,In_1668);
or U2285 (N_2285,In_433,In_1328);
and U2286 (N_2286,In_1670,In_1041);
nand U2287 (N_2287,In_1782,In_1779);
or U2288 (N_2288,In_277,In_216);
nor U2289 (N_2289,In_620,In_1558);
or U2290 (N_2290,In_1115,In_101);
nor U2291 (N_2291,In_342,In_1829);
xnor U2292 (N_2292,In_1311,In_1060);
nand U2293 (N_2293,In_1193,In_1618);
and U2294 (N_2294,In_1844,In_1142);
or U2295 (N_2295,In_806,In_1416);
or U2296 (N_2296,In_1372,In_450);
and U2297 (N_2297,In_1688,In_1316);
xnor U2298 (N_2298,In_1023,In_1987);
nand U2299 (N_2299,In_1039,In_829);
xnor U2300 (N_2300,In_527,In_125);
nor U2301 (N_2301,In_262,In_564);
and U2302 (N_2302,In_153,In_1599);
or U2303 (N_2303,In_630,In_1134);
xnor U2304 (N_2304,In_1986,In_835);
xor U2305 (N_2305,In_330,In_691);
or U2306 (N_2306,In_1821,In_1034);
or U2307 (N_2307,In_1407,In_367);
xnor U2308 (N_2308,In_1353,In_58);
or U2309 (N_2309,In_871,In_348);
and U2310 (N_2310,In_1883,In_1289);
nor U2311 (N_2311,In_1024,In_214);
or U2312 (N_2312,In_891,In_436);
or U2313 (N_2313,In_1535,In_686);
and U2314 (N_2314,In_336,In_1991);
or U2315 (N_2315,In_848,In_1273);
nand U2316 (N_2316,In_530,In_1336);
and U2317 (N_2317,In_873,In_222);
xor U2318 (N_2318,In_1051,In_671);
or U2319 (N_2319,In_724,In_1006);
nand U2320 (N_2320,In_585,In_1558);
or U2321 (N_2321,In_1813,In_1556);
nor U2322 (N_2322,In_1416,In_1866);
nor U2323 (N_2323,In_1686,In_33);
nand U2324 (N_2324,In_583,In_1913);
nor U2325 (N_2325,In_1091,In_1835);
nor U2326 (N_2326,In_1214,In_1680);
or U2327 (N_2327,In_30,In_1229);
nor U2328 (N_2328,In_376,In_235);
nand U2329 (N_2329,In_886,In_1902);
xor U2330 (N_2330,In_1217,In_1755);
xor U2331 (N_2331,In_129,In_1275);
and U2332 (N_2332,In_186,In_1861);
nand U2333 (N_2333,In_1792,In_940);
nand U2334 (N_2334,In_65,In_289);
xnor U2335 (N_2335,In_984,In_1213);
nand U2336 (N_2336,In_64,In_139);
nor U2337 (N_2337,In_257,In_1000);
nor U2338 (N_2338,In_226,In_1035);
xor U2339 (N_2339,In_157,In_1165);
and U2340 (N_2340,In_672,In_1115);
xnor U2341 (N_2341,In_1186,In_817);
xor U2342 (N_2342,In_1760,In_367);
nor U2343 (N_2343,In_1802,In_347);
xor U2344 (N_2344,In_1417,In_1777);
nand U2345 (N_2345,In_1369,In_1165);
nand U2346 (N_2346,In_1215,In_636);
xnor U2347 (N_2347,In_1082,In_330);
xor U2348 (N_2348,In_1217,In_1608);
nor U2349 (N_2349,In_376,In_1343);
or U2350 (N_2350,In_1960,In_1778);
or U2351 (N_2351,In_1631,In_1651);
nor U2352 (N_2352,In_948,In_551);
nand U2353 (N_2353,In_830,In_1554);
nand U2354 (N_2354,In_340,In_334);
or U2355 (N_2355,In_987,In_735);
nor U2356 (N_2356,In_959,In_1353);
nor U2357 (N_2357,In_1891,In_873);
and U2358 (N_2358,In_1977,In_489);
and U2359 (N_2359,In_1932,In_1445);
and U2360 (N_2360,In_1651,In_327);
nor U2361 (N_2361,In_156,In_618);
nand U2362 (N_2362,In_858,In_783);
or U2363 (N_2363,In_747,In_7);
nor U2364 (N_2364,In_555,In_1317);
nor U2365 (N_2365,In_33,In_815);
xor U2366 (N_2366,In_1026,In_503);
nor U2367 (N_2367,In_1812,In_267);
nand U2368 (N_2368,In_1432,In_364);
xor U2369 (N_2369,In_1424,In_1060);
and U2370 (N_2370,In_910,In_52);
and U2371 (N_2371,In_1078,In_28);
nand U2372 (N_2372,In_1743,In_548);
and U2373 (N_2373,In_1248,In_421);
nand U2374 (N_2374,In_1863,In_682);
xnor U2375 (N_2375,In_1318,In_1916);
nor U2376 (N_2376,In_503,In_745);
nor U2377 (N_2377,In_1109,In_1907);
nor U2378 (N_2378,In_1255,In_1277);
or U2379 (N_2379,In_1904,In_321);
xor U2380 (N_2380,In_441,In_1856);
or U2381 (N_2381,In_1373,In_1956);
or U2382 (N_2382,In_1629,In_247);
and U2383 (N_2383,In_426,In_202);
nor U2384 (N_2384,In_102,In_1052);
xnor U2385 (N_2385,In_148,In_1767);
and U2386 (N_2386,In_649,In_1338);
or U2387 (N_2387,In_1608,In_1650);
or U2388 (N_2388,In_573,In_847);
nand U2389 (N_2389,In_382,In_1000);
or U2390 (N_2390,In_53,In_769);
nand U2391 (N_2391,In_208,In_1235);
nand U2392 (N_2392,In_1002,In_1964);
nand U2393 (N_2393,In_1485,In_1861);
and U2394 (N_2394,In_493,In_1172);
xnor U2395 (N_2395,In_1288,In_1121);
nand U2396 (N_2396,In_1097,In_1713);
or U2397 (N_2397,In_1787,In_750);
xor U2398 (N_2398,In_851,In_614);
or U2399 (N_2399,In_1426,In_1786);
xor U2400 (N_2400,In_711,In_352);
nand U2401 (N_2401,In_883,In_1648);
and U2402 (N_2402,In_1886,In_274);
and U2403 (N_2403,In_917,In_1198);
or U2404 (N_2404,In_1693,In_71);
xor U2405 (N_2405,In_1568,In_1851);
nand U2406 (N_2406,In_647,In_115);
nand U2407 (N_2407,In_1852,In_622);
and U2408 (N_2408,In_669,In_1338);
xor U2409 (N_2409,In_374,In_930);
xor U2410 (N_2410,In_1871,In_536);
and U2411 (N_2411,In_469,In_1889);
nor U2412 (N_2412,In_362,In_628);
nor U2413 (N_2413,In_704,In_1673);
nor U2414 (N_2414,In_123,In_696);
xor U2415 (N_2415,In_1989,In_1114);
xnor U2416 (N_2416,In_1903,In_647);
or U2417 (N_2417,In_134,In_1306);
nor U2418 (N_2418,In_97,In_463);
and U2419 (N_2419,In_1624,In_1110);
nor U2420 (N_2420,In_1952,In_876);
xor U2421 (N_2421,In_1008,In_660);
or U2422 (N_2422,In_625,In_1240);
and U2423 (N_2423,In_860,In_1802);
or U2424 (N_2424,In_1093,In_1737);
nand U2425 (N_2425,In_838,In_1804);
nor U2426 (N_2426,In_1994,In_69);
nor U2427 (N_2427,In_958,In_126);
nor U2428 (N_2428,In_800,In_1820);
nor U2429 (N_2429,In_1097,In_789);
xor U2430 (N_2430,In_1738,In_1908);
xor U2431 (N_2431,In_269,In_145);
nand U2432 (N_2432,In_351,In_86);
and U2433 (N_2433,In_1681,In_219);
xor U2434 (N_2434,In_936,In_1227);
xor U2435 (N_2435,In_1695,In_117);
or U2436 (N_2436,In_418,In_414);
nor U2437 (N_2437,In_1370,In_90);
or U2438 (N_2438,In_1916,In_955);
xnor U2439 (N_2439,In_785,In_847);
nand U2440 (N_2440,In_1544,In_121);
or U2441 (N_2441,In_1956,In_1816);
and U2442 (N_2442,In_1342,In_806);
xor U2443 (N_2443,In_1613,In_1445);
nand U2444 (N_2444,In_674,In_1068);
and U2445 (N_2445,In_553,In_153);
nand U2446 (N_2446,In_583,In_1173);
or U2447 (N_2447,In_1342,In_543);
xor U2448 (N_2448,In_484,In_1763);
nand U2449 (N_2449,In_1328,In_1921);
and U2450 (N_2450,In_1273,In_1971);
or U2451 (N_2451,In_476,In_591);
nand U2452 (N_2452,In_171,In_62);
nand U2453 (N_2453,In_617,In_1206);
or U2454 (N_2454,In_933,In_1406);
nand U2455 (N_2455,In_233,In_264);
and U2456 (N_2456,In_716,In_1297);
nor U2457 (N_2457,In_596,In_1102);
nand U2458 (N_2458,In_119,In_629);
or U2459 (N_2459,In_1548,In_1917);
nand U2460 (N_2460,In_1233,In_288);
or U2461 (N_2461,In_1714,In_803);
nor U2462 (N_2462,In_165,In_684);
and U2463 (N_2463,In_965,In_1801);
xnor U2464 (N_2464,In_1928,In_1464);
nor U2465 (N_2465,In_1102,In_1231);
nor U2466 (N_2466,In_1291,In_390);
and U2467 (N_2467,In_248,In_1305);
or U2468 (N_2468,In_1911,In_1772);
xnor U2469 (N_2469,In_382,In_621);
xnor U2470 (N_2470,In_1442,In_960);
and U2471 (N_2471,In_62,In_430);
nor U2472 (N_2472,In_1187,In_448);
xnor U2473 (N_2473,In_1196,In_1684);
xor U2474 (N_2474,In_250,In_1466);
nor U2475 (N_2475,In_627,In_210);
nand U2476 (N_2476,In_117,In_1856);
or U2477 (N_2477,In_1124,In_1907);
nor U2478 (N_2478,In_784,In_1673);
nand U2479 (N_2479,In_1080,In_476);
nor U2480 (N_2480,In_858,In_1787);
xnor U2481 (N_2481,In_1332,In_918);
nand U2482 (N_2482,In_162,In_939);
nand U2483 (N_2483,In_1202,In_118);
nand U2484 (N_2484,In_1393,In_1695);
or U2485 (N_2485,In_1549,In_842);
and U2486 (N_2486,In_1873,In_1943);
xnor U2487 (N_2487,In_1389,In_510);
nand U2488 (N_2488,In_1513,In_642);
nor U2489 (N_2489,In_583,In_657);
and U2490 (N_2490,In_1088,In_1311);
nand U2491 (N_2491,In_903,In_1838);
nor U2492 (N_2492,In_311,In_494);
or U2493 (N_2493,In_1940,In_1698);
nand U2494 (N_2494,In_1275,In_1159);
and U2495 (N_2495,In_894,In_1423);
nand U2496 (N_2496,In_964,In_1197);
and U2497 (N_2497,In_1401,In_921);
xor U2498 (N_2498,In_1985,In_833);
nand U2499 (N_2499,In_342,In_506);
nand U2500 (N_2500,In_612,In_505);
nor U2501 (N_2501,In_983,In_911);
or U2502 (N_2502,In_951,In_618);
nor U2503 (N_2503,In_904,In_865);
nand U2504 (N_2504,In_1014,In_335);
xnor U2505 (N_2505,In_1332,In_1437);
xnor U2506 (N_2506,In_421,In_207);
nor U2507 (N_2507,In_1973,In_802);
or U2508 (N_2508,In_1364,In_304);
and U2509 (N_2509,In_1921,In_1658);
xor U2510 (N_2510,In_1303,In_905);
or U2511 (N_2511,In_1764,In_644);
nand U2512 (N_2512,In_670,In_1688);
nand U2513 (N_2513,In_33,In_1540);
or U2514 (N_2514,In_1530,In_1139);
nand U2515 (N_2515,In_177,In_1123);
or U2516 (N_2516,In_716,In_836);
xnor U2517 (N_2517,In_761,In_715);
or U2518 (N_2518,In_1076,In_166);
nor U2519 (N_2519,In_1994,In_1960);
and U2520 (N_2520,In_1128,In_689);
or U2521 (N_2521,In_474,In_145);
nand U2522 (N_2522,In_289,In_1355);
nor U2523 (N_2523,In_823,In_1835);
nand U2524 (N_2524,In_903,In_1532);
or U2525 (N_2525,In_265,In_941);
nor U2526 (N_2526,In_641,In_1411);
xor U2527 (N_2527,In_1192,In_1735);
or U2528 (N_2528,In_574,In_1896);
nor U2529 (N_2529,In_1868,In_472);
nor U2530 (N_2530,In_527,In_1427);
xor U2531 (N_2531,In_661,In_1174);
nor U2532 (N_2532,In_1993,In_1787);
and U2533 (N_2533,In_139,In_1801);
and U2534 (N_2534,In_1778,In_1439);
nor U2535 (N_2535,In_1265,In_219);
nor U2536 (N_2536,In_1967,In_279);
nor U2537 (N_2537,In_1249,In_60);
nor U2538 (N_2538,In_1752,In_1354);
xor U2539 (N_2539,In_1608,In_183);
and U2540 (N_2540,In_1462,In_708);
nor U2541 (N_2541,In_1866,In_385);
or U2542 (N_2542,In_145,In_1232);
or U2543 (N_2543,In_322,In_753);
or U2544 (N_2544,In_1370,In_103);
nor U2545 (N_2545,In_1472,In_1666);
nand U2546 (N_2546,In_1792,In_344);
and U2547 (N_2547,In_231,In_1906);
or U2548 (N_2548,In_599,In_1718);
or U2549 (N_2549,In_1308,In_1978);
xnor U2550 (N_2550,In_1052,In_308);
xor U2551 (N_2551,In_1141,In_216);
and U2552 (N_2552,In_211,In_1654);
xor U2553 (N_2553,In_1654,In_170);
and U2554 (N_2554,In_1681,In_1740);
nand U2555 (N_2555,In_53,In_1881);
or U2556 (N_2556,In_1368,In_1967);
nand U2557 (N_2557,In_1208,In_588);
nor U2558 (N_2558,In_529,In_1041);
nand U2559 (N_2559,In_181,In_851);
nand U2560 (N_2560,In_855,In_554);
and U2561 (N_2561,In_897,In_68);
nand U2562 (N_2562,In_1214,In_620);
nor U2563 (N_2563,In_309,In_1326);
xnor U2564 (N_2564,In_294,In_750);
nand U2565 (N_2565,In_4,In_563);
nor U2566 (N_2566,In_1346,In_1139);
nor U2567 (N_2567,In_868,In_324);
and U2568 (N_2568,In_396,In_1762);
and U2569 (N_2569,In_1002,In_1779);
nor U2570 (N_2570,In_153,In_186);
nand U2571 (N_2571,In_975,In_1510);
xor U2572 (N_2572,In_242,In_1946);
nand U2573 (N_2573,In_265,In_196);
nor U2574 (N_2574,In_776,In_1291);
or U2575 (N_2575,In_1188,In_896);
nor U2576 (N_2576,In_1756,In_1745);
and U2577 (N_2577,In_1704,In_13);
nand U2578 (N_2578,In_1670,In_1482);
nand U2579 (N_2579,In_923,In_1670);
and U2580 (N_2580,In_384,In_563);
or U2581 (N_2581,In_91,In_369);
nand U2582 (N_2582,In_1015,In_1819);
or U2583 (N_2583,In_1418,In_702);
nor U2584 (N_2584,In_173,In_1302);
and U2585 (N_2585,In_891,In_1852);
xor U2586 (N_2586,In_1067,In_1952);
nand U2587 (N_2587,In_1882,In_849);
xnor U2588 (N_2588,In_903,In_777);
nand U2589 (N_2589,In_331,In_919);
and U2590 (N_2590,In_1140,In_563);
or U2591 (N_2591,In_1697,In_1573);
or U2592 (N_2592,In_214,In_1796);
nor U2593 (N_2593,In_1589,In_1458);
nand U2594 (N_2594,In_1372,In_685);
nand U2595 (N_2595,In_1061,In_1240);
or U2596 (N_2596,In_1970,In_812);
xnor U2597 (N_2597,In_906,In_127);
xnor U2598 (N_2598,In_845,In_250);
nand U2599 (N_2599,In_553,In_1473);
nor U2600 (N_2600,In_331,In_1982);
nor U2601 (N_2601,In_682,In_278);
and U2602 (N_2602,In_1251,In_25);
and U2603 (N_2603,In_381,In_861);
xor U2604 (N_2604,In_875,In_760);
or U2605 (N_2605,In_482,In_1757);
nor U2606 (N_2606,In_897,In_1315);
or U2607 (N_2607,In_606,In_346);
nand U2608 (N_2608,In_290,In_1401);
xnor U2609 (N_2609,In_563,In_1038);
nand U2610 (N_2610,In_154,In_457);
xor U2611 (N_2611,In_896,In_449);
or U2612 (N_2612,In_349,In_568);
and U2613 (N_2613,In_477,In_870);
xor U2614 (N_2614,In_294,In_949);
or U2615 (N_2615,In_165,In_1809);
and U2616 (N_2616,In_291,In_50);
nor U2617 (N_2617,In_982,In_632);
or U2618 (N_2618,In_979,In_1217);
and U2619 (N_2619,In_1456,In_94);
nor U2620 (N_2620,In_215,In_1168);
xnor U2621 (N_2621,In_326,In_1543);
nor U2622 (N_2622,In_789,In_572);
or U2623 (N_2623,In_118,In_705);
and U2624 (N_2624,In_695,In_676);
nand U2625 (N_2625,In_201,In_456);
xor U2626 (N_2626,In_21,In_933);
nand U2627 (N_2627,In_1249,In_373);
nor U2628 (N_2628,In_1377,In_1681);
nor U2629 (N_2629,In_1027,In_1861);
nand U2630 (N_2630,In_201,In_1822);
or U2631 (N_2631,In_1771,In_840);
xor U2632 (N_2632,In_910,In_1465);
xor U2633 (N_2633,In_613,In_1136);
xnor U2634 (N_2634,In_1054,In_387);
xor U2635 (N_2635,In_421,In_1066);
nor U2636 (N_2636,In_625,In_180);
xnor U2637 (N_2637,In_307,In_1833);
nor U2638 (N_2638,In_141,In_336);
nand U2639 (N_2639,In_726,In_798);
nor U2640 (N_2640,In_1489,In_1881);
nor U2641 (N_2641,In_1324,In_1136);
or U2642 (N_2642,In_1176,In_181);
xnor U2643 (N_2643,In_1224,In_1586);
xor U2644 (N_2644,In_1692,In_76);
or U2645 (N_2645,In_1594,In_334);
xnor U2646 (N_2646,In_58,In_215);
nor U2647 (N_2647,In_1450,In_894);
nand U2648 (N_2648,In_194,In_936);
and U2649 (N_2649,In_1294,In_795);
and U2650 (N_2650,In_1792,In_55);
or U2651 (N_2651,In_1015,In_29);
nand U2652 (N_2652,In_1451,In_1979);
and U2653 (N_2653,In_1733,In_399);
and U2654 (N_2654,In_215,In_855);
or U2655 (N_2655,In_969,In_929);
or U2656 (N_2656,In_366,In_741);
xnor U2657 (N_2657,In_91,In_401);
or U2658 (N_2658,In_1007,In_1779);
or U2659 (N_2659,In_1343,In_662);
and U2660 (N_2660,In_1168,In_490);
nor U2661 (N_2661,In_861,In_825);
and U2662 (N_2662,In_239,In_270);
nor U2663 (N_2663,In_1423,In_699);
nor U2664 (N_2664,In_1530,In_575);
nand U2665 (N_2665,In_374,In_1433);
or U2666 (N_2666,In_256,In_44);
nand U2667 (N_2667,In_1224,In_316);
nand U2668 (N_2668,In_144,In_1718);
xnor U2669 (N_2669,In_1948,In_533);
or U2670 (N_2670,In_953,In_1638);
xor U2671 (N_2671,In_1239,In_1590);
nor U2672 (N_2672,In_1328,In_698);
nor U2673 (N_2673,In_825,In_1431);
or U2674 (N_2674,In_1353,In_191);
and U2675 (N_2675,In_1643,In_30);
and U2676 (N_2676,In_1723,In_912);
or U2677 (N_2677,In_461,In_1795);
or U2678 (N_2678,In_1634,In_1027);
nand U2679 (N_2679,In_668,In_1875);
or U2680 (N_2680,In_369,In_288);
nand U2681 (N_2681,In_1957,In_1597);
nand U2682 (N_2682,In_897,In_1527);
nand U2683 (N_2683,In_939,In_515);
xnor U2684 (N_2684,In_761,In_1302);
nor U2685 (N_2685,In_308,In_698);
or U2686 (N_2686,In_643,In_1353);
xor U2687 (N_2687,In_593,In_152);
nand U2688 (N_2688,In_1144,In_188);
nor U2689 (N_2689,In_598,In_444);
xor U2690 (N_2690,In_1219,In_1212);
xor U2691 (N_2691,In_1943,In_1776);
nor U2692 (N_2692,In_1237,In_1823);
nand U2693 (N_2693,In_33,In_373);
nand U2694 (N_2694,In_1443,In_880);
nor U2695 (N_2695,In_545,In_1652);
nor U2696 (N_2696,In_1552,In_221);
and U2697 (N_2697,In_811,In_1038);
nor U2698 (N_2698,In_825,In_661);
xor U2699 (N_2699,In_82,In_1051);
or U2700 (N_2700,In_391,In_986);
nand U2701 (N_2701,In_32,In_1670);
and U2702 (N_2702,In_1062,In_59);
nor U2703 (N_2703,In_1286,In_593);
nand U2704 (N_2704,In_1273,In_200);
or U2705 (N_2705,In_1178,In_1558);
or U2706 (N_2706,In_571,In_1378);
nand U2707 (N_2707,In_1073,In_1454);
nand U2708 (N_2708,In_1678,In_636);
or U2709 (N_2709,In_756,In_468);
and U2710 (N_2710,In_1362,In_1347);
xnor U2711 (N_2711,In_868,In_1079);
and U2712 (N_2712,In_1038,In_545);
or U2713 (N_2713,In_1009,In_76);
nor U2714 (N_2714,In_437,In_290);
xnor U2715 (N_2715,In_1852,In_1997);
or U2716 (N_2716,In_362,In_601);
nor U2717 (N_2717,In_750,In_1084);
or U2718 (N_2718,In_1963,In_1246);
and U2719 (N_2719,In_764,In_851);
and U2720 (N_2720,In_1543,In_1041);
nor U2721 (N_2721,In_396,In_1710);
or U2722 (N_2722,In_1943,In_320);
xnor U2723 (N_2723,In_534,In_38);
or U2724 (N_2724,In_340,In_1986);
xnor U2725 (N_2725,In_289,In_789);
or U2726 (N_2726,In_1369,In_413);
and U2727 (N_2727,In_689,In_826);
nor U2728 (N_2728,In_970,In_291);
xnor U2729 (N_2729,In_368,In_1961);
or U2730 (N_2730,In_1143,In_1482);
and U2731 (N_2731,In_1373,In_943);
nor U2732 (N_2732,In_1576,In_1839);
nand U2733 (N_2733,In_1079,In_942);
nand U2734 (N_2734,In_541,In_1884);
nand U2735 (N_2735,In_1499,In_1474);
nand U2736 (N_2736,In_968,In_179);
and U2737 (N_2737,In_129,In_672);
nand U2738 (N_2738,In_956,In_867);
nor U2739 (N_2739,In_1431,In_1605);
or U2740 (N_2740,In_19,In_660);
xnor U2741 (N_2741,In_148,In_1853);
or U2742 (N_2742,In_1513,In_1951);
nand U2743 (N_2743,In_0,In_889);
nand U2744 (N_2744,In_661,In_1263);
nor U2745 (N_2745,In_632,In_1085);
or U2746 (N_2746,In_1067,In_996);
and U2747 (N_2747,In_1322,In_818);
nor U2748 (N_2748,In_1148,In_1927);
nor U2749 (N_2749,In_721,In_1064);
and U2750 (N_2750,In_559,In_726);
or U2751 (N_2751,In_264,In_27);
nand U2752 (N_2752,In_1590,In_1838);
nand U2753 (N_2753,In_405,In_1521);
xnor U2754 (N_2754,In_1639,In_384);
and U2755 (N_2755,In_1492,In_136);
or U2756 (N_2756,In_564,In_1645);
nand U2757 (N_2757,In_909,In_147);
nor U2758 (N_2758,In_1256,In_963);
xor U2759 (N_2759,In_1624,In_552);
or U2760 (N_2760,In_1338,In_48);
nand U2761 (N_2761,In_359,In_1524);
or U2762 (N_2762,In_984,In_777);
xnor U2763 (N_2763,In_1379,In_824);
nor U2764 (N_2764,In_1757,In_981);
or U2765 (N_2765,In_715,In_617);
nand U2766 (N_2766,In_1222,In_1678);
nand U2767 (N_2767,In_470,In_1981);
nor U2768 (N_2768,In_1774,In_373);
and U2769 (N_2769,In_344,In_1158);
nor U2770 (N_2770,In_1168,In_901);
or U2771 (N_2771,In_1473,In_1339);
and U2772 (N_2772,In_605,In_313);
nor U2773 (N_2773,In_1213,In_263);
nor U2774 (N_2774,In_1388,In_784);
nand U2775 (N_2775,In_424,In_1621);
and U2776 (N_2776,In_714,In_1728);
nor U2777 (N_2777,In_670,In_1173);
nand U2778 (N_2778,In_1303,In_891);
and U2779 (N_2779,In_893,In_75);
and U2780 (N_2780,In_603,In_1488);
nor U2781 (N_2781,In_1171,In_554);
xor U2782 (N_2782,In_1253,In_923);
and U2783 (N_2783,In_487,In_927);
and U2784 (N_2784,In_552,In_1399);
nand U2785 (N_2785,In_536,In_1236);
xnor U2786 (N_2786,In_243,In_1746);
or U2787 (N_2787,In_881,In_777);
or U2788 (N_2788,In_216,In_823);
or U2789 (N_2789,In_1745,In_813);
or U2790 (N_2790,In_253,In_633);
xnor U2791 (N_2791,In_139,In_1731);
or U2792 (N_2792,In_1095,In_1168);
nor U2793 (N_2793,In_622,In_1026);
nor U2794 (N_2794,In_1476,In_657);
nand U2795 (N_2795,In_118,In_1384);
nor U2796 (N_2796,In_1743,In_415);
nor U2797 (N_2797,In_543,In_91);
and U2798 (N_2798,In_1202,In_808);
xor U2799 (N_2799,In_539,In_1519);
and U2800 (N_2800,In_1062,In_1000);
or U2801 (N_2801,In_141,In_1992);
nand U2802 (N_2802,In_655,In_576);
or U2803 (N_2803,In_1570,In_253);
nor U2804 (N_2804,In_1613,In_1506);
nand U2805 (N_2805,In_1477,In_1030);
or U2806 (N_2806,In_565,In_278);
xor U2807 (N_2807,In_785,In_1856);
or U2808 (N_2808,In_1302,In_1945);
nand U2809 (N_2809,In_1522,In_1154);
and U2810 (N_2810,In_137,In_989);
nand U2811 (N_2811,In_1541,In_247);
xor U2812 (N_2812,In_1944,In_495);
nand U2813 (N_2813,In_1445,In_1694);
xor U2814 (N_2814,In_1436,In_1853);
xor U2815 (N_2815,In_110,In_1497);
xor U2816 (N_2816,In_991,In_49);
nand U2817 (N_2817,In_936,In_1147);
or U2818 (N_2818,In_513,In_435);
nand U2819 (N_2819,In_1958,In_839);
xnor U2820 (N_2820,In_1950,In_213);
or U2821 (N_2821,In_30,In_1951);
and U2822 (N_2822,In_1064,In_1050);
xnor U2823 (N_2823,In_841,In_304);
nand U2824 (N_2824,In_115,In_1818);
or U2825 (N_2825,In_549,In_1582);
nor U2826 (N_2826,In_1403,In_636);
xnor U2827 (N_2827,In_284,In_1694);
and U2828 (N_2828,In_178,In_774);
xnor U2829 (N_2829,In_1436,In_1661);
or U2830 (N_2830,In_1371,In_1782);
xnor U2831 (N_2831,In_1125,In_1066);
nor U2832 (N_2832,In_136,In_1313);
and U2833 (N_2833,In_942,In_1883);
xnor U2834 (N_2834,In_1963,In_1244);
nand U2835 (N_2835,In_632,In_395);
or U2836 (N_2836,In_1518,In_814);
nand U2837 (N_2837,In_789,In_347);
xnor U2838 (N_2838,In_1370,In_1937);
xor U2839 (N_2839,In_534,In_723);
or U2840 (N_2840,In_888,In_127);
xor U2841 (N_2841,In_712,In_1979);
xor U2842 (N_2842,In_643,In_600);
and U2843 (N_2843,In_894,In_677);
xor U2844 (N_2844,In_920,In_587);
xor U2845 (N_2845,In_1611,In_86);
and U2846 (N_2846,In_1584,In_1094);
and U2847 (N_2847,In_1549,In_209);
nand U2848 (N_2848,In_820,In_828);
nor U2849 (N_2849,In_1652,In_1035);
nor U2850 (N_2850,In_1571,In_275);
and U2851 (N_2851,In_944,In_502);
nand U2852 (N_2852,In_852,In_1570);
and U2853 (N_2853,In_980,In_414);
xnor U2854 (N_2854,In_1934,In_1786);
nor U2855 (N_2855,In_425,In_634);
or U2856 (N_2856,In_743,In_1830);
or U2857 (N_2857,In_29,In_75);
and U2858 (N_2858,In_1493,In_1867);
or U2859 (N_2859,In_1406,In_1477);
xor U2860 (N_2860,In_1567,In_326);
nor U2861 (N_2861,In_763,In_1741);
or U2862 (N_2862,In_1904,In_460);
or U2863 (N_2863,In_696,In_1255);
nor U2864 (N_2864,In_1476,In_1355);
or U2865 (N_2865,In_905,In_1353);
or U2866 (N_2866,In_1612,In_958);
xnor U2867 (N_2867,In_304,In_1207);
or U2868 (N_2868,In_568,In_983);
and U2869 (N_2869,In_422,In_1836);
and U2870 (N_2870,In_1667,In_757);
and U2871 (N_2871,In_1519,In_1247);
and U2872 (N_2872,In_1054,In_1333);
and U2873 (N_2873,In_524,In_1398);
nor U2874 (N_2874,In_177,In_1249);
xor U2875 (N_2875,In_408,In_1150);
nor U2876 (N_2876,In_1874,In_1266);
and U2877 (N_2877,In_656,In_905);
nor U2878 (N_2878,In_1207,In_446);
and U2879 (N_2879,In_669,In_987);
nand U2880 (N_2880,In_982,In_276);
nand U2881 (N_2881,In_852,In_888);
and U2882 (N_2882,In_1267,In_715);
nor U2883 (N_2883,In_1562,In_330);
and U2884 (N_2884,In_348,In_425);
and U2885 (N_2885,In_808,In_1966);
xnor U2886 (N_2886,In_618,In_1462);
xor U2887 (N_2887,In_992,In_1759);
nand U2888 (N_2888,In_1117,In_1007);
and U2889 (N_2889,In_46,In_1608);
or U2890 (N_2890,In_259,In_62);
nand U2891 (N_2891,In_922,In_1790);
or U2892 (N_2892,In_1891,In_1775);
xnor U2893 (N_2893,In_612,In_1041);
nor U2894 (N_2894,In_915,In_219);
or U2895 (N_2895,In_747,In_858);
or U2896 (N_2896,In_363,In_1367);
nand U2897 (N_2897,In_1935,In_238);
nand U2898 (N_2898,In_717,In_221);
nand U2899 (N_2899,In_456,In_272);
nand U2900 (N_2900,In_543,In_1296);
xnor U2901 (N_2901,In_906,In_797);
xnor U2902 (N_2902,In_1695,In_1614);
or U2903 (N_2903,In_1809,In_1390);
and U2904 (N_2904,In_1995,In_609);
nand U2905 (N_2905,In_433,In_1638);
nand U2906 (N_2906,In_1425,In_1583);
xor U2907 (N_2907,In_469,In_286);
xor U2908 (N_2908,In_1874,In_638);
nor U2909 (N_2909,In_1125,In_631);
nor U2910 (N_2910,In_1678,In_699);
xnor U2911 (N_2911,In_1782,In_564);
xnor U2912 (N_2912,In_335,In_809);
nand U2913 (N_2913,In_393,In_1018);
nand U2914 (N_2914,In_1827,In_1860);
or U2915 (N_2915,In_466,In_289);
xnor U2916 (N_2916,In_1093,In_1108);
and U2917 (N_2917,In_452,In_502);
or U2918 (N_2918,In_1996,In_1132);
and U2919 (N_2919,In_1930,In_608);
nor U2920 (N_2920,In_1807,In_1971);
nand U2921 (N_2921,In_817,In_1376);
and U2922 (N_2922,In_807,In_1674);
or U2923 (N_2923,In_1459,In_755);
nor U2924 (N_2924,In_973,In_13);
nand U2925 (N_2925,In_607,In_1310);
or U2926 (N_2926,In_1255,In_1676);
or U2927 (N_2927,In_980,In_1986);
xor U2928 (N_2928,In_1284,In_564);
or U2929 (N_2929,In_334,In_266);
xor U2930 (N_2930,In_1959,In_1229);
or U2931 (N_2931,In_540,In_586);
and U2932 (N_2932,In_815,In_693);
nor U2933 (N_2933,In_568,In_1097);
nor U2934 (N_2934,In_380,In_1042);
nand U2935 (N_2935,In_788,In_411);
nand U2936 (N_2936,In_195,In_1364);
nor U2937 (N_2937,In_855,In_793);
and U2938 (N_2938,In_1418,In_903);
or U2939 (N_2939,In_946,In_1455);
or U2940 (N_2940,In_337,In_936);
nor U2941 (N_2941,In_1940,In_1710);
nand U2942 (N_2942,In_1243,In_1117);
and U2943 (N_2943,In_584,In_1707);
nor U2944 (N_2944,In_641,In_1043);
nand U2945 (N_2945,In_1428,In_1356);
nor U2946 (N_2946,In_1444,In_810);
or U2947 (N_2947,In_1436,In_1453);
xnor U2948 (N_2948,In_408,In_1602);
nand U2949 (N_2949,In_417,In_1717);
nor U2950 (N_2950,In_1597,In_1004);
or U2951 (N_2951,In_1905,In_694);
nor U2952 (N_2952,In_1699,In_40);
nor U2953 (N_2953,In_1070,In_422);
nand U2954 (N_2954,In_1936,In_286);
and U2955 (N_2955,In_1516,In_948);
and U2956 (N_2956,In_1831,In_130);
nand U2957 (N_2957,In_1429,In_1143);
nand U2958 (N_2958,In_1898,In_370);
nand U2959 (N_2959,In_208,In_1474);
and U2960 (N_2960,In_973,In_1658);
nor U2961 (N_2961,In_1684,In_150);
or U2962 (N_2962,In_1095,In_1714);
and U2963 (N_2963,In_657,In_541);
nor U2964 (N_2964,In_1798,In_35);
xor U2965 (N_2965,In_1174,In_1939);
nand U2966 (N_2966,In_377,In_539);
nand U2967 (N_2967,In_83,In_326);
or U2968 (N_2968,In_969,In_1408);
xor U2969 (N_2969,In_1466,In_1474);
nand U2970 (N_2970,In_1874,In_840);
nor U2971 (N_2971,In_1008,In_933);
nor U2972 (N_2972,In_1170,In_671);
or U2973 (N_2973,In_1943,In_1573);
and U2974 (N_2974,In_397,In_1560);
nand U2975 (N_2975,In_1199,In_1837);
xor U2976 (N_2976,In_1232,In_1649);
nor U2977 (N_2977,In_1348,In_835);
or U2978 (N_2978,In_1855,In_1886);
or U2979 (N_2979,In_639,In_1087);
xor U2980 (N_2980,In_9,In_483);
and U2981 (N_2981,In_1106,In_1348);
and U2982 (N_2982,In_330,In_254);
nand U2983 (N_2983,In_1294,In_628);
nor U2984 (N_2984,In_1004,In_271);
xor U2985 (N_2985,In_1579,In_905);
nor U2986 (N_2986,In_803,In_889);
and U2987 (N_2987,In_1052,In_1627);
or U2988 (N_2988,In_1017,In_1561);
xor U2989 (N_2989,In_108,In_1819);
nand U2990 (N_2990,In_1438,In_347);
xor U2991 (N_2991,In_269,In_35);
nand U2992 (N_2992,In_224,In_1712);
or U2993 (N_2993,In_1834,In_251);
nand U2994 (N_2994,In_219,In_996);
nand U2995 (N_2995,In_1206,In_1590);
nor U2996 (N_2996,In_1306,In_1643);
and U2997 (N_2997,In_1259,In_1421);
xor U2998 (N_2998,In_601,In_1282);
nand U2999 (N_2999,In_1326,In_1097);
or U3000 (N_3000,In_1013,In_471);
or U3001 (N_3001,In_433,In_1931);
and U3002 (N_3002,In_229,In_132);
xnor U3003 (N_3003,In_514,In_471);
xor U3004 (N_3004,In_4,In_1424);
or U3005 (N_3005,In_1492,In_1159);
and U3006 (N_3006,In_468,In_228);
or U3007 (N_3007,In_1624,In_894);
and U3008 (N_3008,In_1868,In_1998);
or U3009 (N_3009,In_1460,In_873);
and U3010 (N_3010,In_1598,In_1578);
nor U3011 (N_3011,In_1476,In_348);
nand U3012 (N_3012,In_526,In_1721);
nand U3013 (N_3013,In_217,In_378);
and U3014 (N_3014,In_1860,In_1921);
or U3015 (N_3015,In_1897,In_1764);
xnor U3016 (N_3016,In_717,In_1629);
nand U3017 (N_3017,In_1360,In_801);
or U3018 (N_3018,In_1536,In_878);
nor U3019 (N_3019,In_1269,In_1929);
or U3020 (N_3020,In_1563,In_48);
xnor U3021 (N_3021,In_1126,In_1548);
nor U3022 (N_3022,In_1766,In_241);
nand U3023 (N_3023,In_747,In_1843);
and U3024 (N_3024,In_616,In_1527);
and U3025 (N_3025,In_1317,In_472);
and U3026 (N_3026,In_311,In_1301);
and U3027 (N_3027,In_1202,In_876);
xor U3028 (N_3028,In_248,In_1902);
and U3029 (N_3029,In_1407,In_1294);
nor U3030 (N_3030,In_830,In_1021);
nand U3031 (N_3031,In_653,In_1713);
nor U3032 (N_3032,In_1070,In_282);
and U3033 (N_3033,In_964,In_1765);
nand U3034 (N_3034,In_1415,In_926);
and U3035 (N_3035,In_150,In_1628);
nand U3036 (N_3036,In_1793,In_533);
nand U3037 (N_3037,In_907,In_1190);
nand U3038 (N_3038,In_1406,In_1128);
nand U3039 (N_3039,In_725,In_858);
xnor U3040 (N_3040,In_915,In_1024);
or U3041 (N_3041,In_1133,In_1196);
nand U3042 (N_3042,In_189,In_1649);
xor U3043 (N_3043,In_1761,In_616);
xnor U3044 (N_3044,In_1777,In_1200);
nor U3045 (N_3045,In_841,In_1667);
nand U3046 (N_3046,In_1709,In_1153);
nand U3047 (N_3047,In_259,In_1061);
xnor U3048 (N_3048,In_745,In_919);
nor U3049 (N_3049,In_1362,In_1854);
xnor U3050 (N_3050,In_962,In_217);
nor U3051 (N_3051,In_90,In_38);
nor U3052 (N_3052,In_917,In_843);
nand U3053 (N_3053,In_1607,In_653);
or U3054 (N_3054,In_1054,In_136);
xnor U3055 (N_3055,In_355,In_1180);
and U3056 (N_3056,In_1300,In_1007);
nand U3057 (N_3057,In_566,In_45);
xnor U3058 (N_3058,In_1581,In_1974);
nand U3059 (N_3059,In_7,In_1276);
xnor U3060 (N_3060,In_541,In_877);
xor U3061 (N_3061,In_976,In_135);
nor U3062 (N_3062,In_1911,In_1077);
or U3063 (N_3063,In_639,In_475);
and U3064 (N_3064,In_551,In_1695);
nor U3065 (N_3065,In_1337,In_130);
or U3066 (N_3066,In_1602,In_1663);
nor U3067 (N_3067,In_1876,In_1209);
xnor U3068 (N_3068,In_12,In_1165);
and U3069 (N_3069,In_582,In_438);
or U3070 (N_3070,In_925,In_1381);
nand U3071 (N_3071,In_651,In_895);
or U3072 (N_3072,In_1222,In_258);
or U3073 (N_3073,In_1863,In_1074);
xnor U3074 (N_3074,In_643,In_412);
and U3075 (N_3075,In_347,In_1119);
and U3076 (N_3076,In_223,In_741);
xnor U3077 (N_3077,In_14,In_315);
nand U3078 (N_3078,In_1524,In_1938);
nand U3079 (N_3079,In_1869,In_1848);
and U3080 (N_3080,In_1694,In_371);
or U3081 (N_3081,In_494,In_869);
nor U3082 (N_3082,In_35,In_970);
xor U3083 (N_3083,In_183,In_1140);
xnor U3084 (N_3084,In_127,In_1599);
and U3085 (N_3085,In_1319,In_66);
xor U3086 (N_3086,In_1649,In_367);
or U3087 (N_3087,In_1539,In_1690);
nor U3088 (N_3088,In_1471,In_1573);
nor U3089 (N_3089,In_270,In_1204);
or U3090 (N_3090,In_457,In_1955);
and U3091 (N_3091,In_686,In_1598);
nor U3092 (N_3092,In_1457,In_138);
and U3093 (N_3093,In_942,In_239);
or U3094 (N_3094,In_929,In_1252);
or U3095 (N_3095,In_328,In_595);
or U3096 (N_3096,In_731,In_1331);
or U3097 (N_3097,In_208,In_612);
and U3098 (N_3098,In_1468,In_728);
nor U3099 (N_3099,In_1028,In_1001);
xnor U3100 (N_3100,In_1144,In_781);
or U3101 (N_3101,In_1629,In_672);
and U3102 (N_3102,In_965,In_438);
xnor U3103 (N_3103,In_1109,In_700);
or U3104 (N_3104,In_843,In_700);
and U3105 (N_3105,In_170,In_1914);
and U3106 (N_3106,In_960,In_891);
nor U3107 (N_3107,In_996,In_563);
and U3108 (N_3108,In_1809,In_1905);
nand U3109 (N_3109,In_408,In_42);
nor U3110 (N_3110,In_1423,In_197);
nand U3111 (N_3111,In_807,In_772);
and U3112 (N_3112,In_1628,In_1707);
or U3113 (N_3113,In_681,In_1365);
xor U3114 (N_3114,In_63,In_1761);
and U3115 (N_3115,In_793,In_1699);
or U3116 (N_3116,In_1971,In_186);
or U3117 (N_3117,In_365,In_1264);
or U3118 (N_3118,In_225,In_1275);
xnor U3119 (N_3119,In_884,In_1970);
or U3120 (N_3120,In_1733,In_300);
nor U3121 (N_3121,In_396,In_522);
and U3122 (N_3122,In_306,In_1996);
and U3123 (N_3123,In_1158,In_1569);
or U3124 (N_3124,In_680,In_689);
nand U3125 (N_3125,In_1921,In_560);
or U3126 (N_3126,In_731,In_1289);
or U3127 (N_3127,In_1151,In_1814);
xnor U3128 (N_3128,In_956,In_297);
xor U3129 (N_3129,In_967,In_997);
nor U3130 (N_3130,In_1347,In_1796);
nor U3131 (N_3131,In_1261,In_151);
nor U3132 (N_3132,In_1955,In_436);
nand U3133 (N_3133,In_457,In_391);
or U3134 (N_3134,In_1684,In_1650);
and U3135 (N_3135,In_853,In_1299);
xor U3136 (N_3136,In_1693,In_1756);
xor U3137 (N_3137,In_371,In_875);
and U3138 (N_3138,In_37,In_1266);
nor U3139 (N_3139,In_877,In_200);
nor U3140 (N_3140,In_480,In_1936);
or U3141 (N_3141,In_389,In_536);
nor U3142 (N_3142,In_1787,In_412);
xor U3143 (N_3143,In_439,In_742);
nor U3144 (N_3144,In_1659,In_1151);
or U3145 (N_3145,In_376,In_934);
nor U3146 (N_3146,In_1696,In_164);
xnor U3147 (N_3147,In_1301,In_1356);
xnor U3148 (N_3148,In_1629,In_1483);
nor U3149 (N_3149,In_1730,In_1618);
nor U3150 (N_3150,In_955,In_793);
nand U3151 (N_3151,In_1497,In_850);
xnor U3152 (N_3152,In_175,In_239);
and U3153 (N_3153,In_293,In_1940);
or U3154 (N_3154,In_1977,In_389);
and U3155 (N_3155,In_1788,In_281);
or U3156 (N_3156,In_394,In_396);
and U3157 (N_3157,In_146,In_1471);
or U3158 (N_3158,In_840,In_1979);
xor U3159 (N_3159,In_30,In_1479);
or U3160 (N_3160,In_1430,In_791);
xnor U3161 (N_3161,In_1908,In_1443);
and U3162 (N_3162,In_1986,In_984);
nor U3163 (N_3163,In_956,In_227);
xor U3164 (N_3164,In_484,In_916);
and U3165 (N_3165,In_1637,In_1366);
nor U3166 (N_3166,In_703,In_821);
xnor U3167 (N_3167,In_481,In_1987);
and U3168 (N_3168,In_1944,In_1490);
nor U3169 (N_3169,In_1806,In_442);
nor U3170 (N_3170,In_238,In_470);
or U3171 (N_3171,In_573,In_852);
or U3172 (N_3172,In_996,In_676);
nor U3173 (N_3173,In_409,In_496);
nor U3174 (N_3174,In_1376,In_1653);
xnor U3175 (N_3175,In_37,In_173);
or U3176 (N_3176,In_849,In_1587);
or U3177 (N_3177,In_530,In_1453);
xor U3178 (N_3178,In_821,In_95);
or U3179 (N_3179,In_744,In_1058);
nor U3180 (N_3180,In_1024,In_1007);
and U3181 (N_3181,In_127,In_565);
or U3182 (N_3182,In_485,In_361);
xor U3183 (N_3183,In_1290,In_1013);
nand U3184 (N_3184,In_828,In_406);
and U3185 (N_3185,In_1960,In_1128);
nand U3186 (N_3186,In_1613,In_1738);
or U3187 (N_3187,In_1351,In_861);
or U3188 (N_3188,In_243,In_1175);
nor U3189 (N_3189,In_1374,In_209);
xor U3190 (N_3190,In_274,In_697);
or U3191 (N_3191,In_398,In_473);
nor U3192 (N_3192,In_1419,In_1607);
xnor U3193 (N_3193,In_1291,In_1576);
xnor U3194 (N_3194,In_1049,In_1695);
or U3195 (N_3195,In_1002,In_1383);
nand U3196 (N_3196,In_1817,In_244);
nand U3197 (N_3197,In_89,In_963);
xnor U3198 (N_3198,In_27,In_50);
xnor U3199 (N_3199,In_1808,In_924);
xor U3200 (N_3200,In_1294,In_310);
nor U3201 (N_3201,In_1717,In_1873);
nand U3202 (N_3202,In_1025,In_1693);
xor U3203 (N_3203,In_1198,In_935);
xor U3204 (N_3204,In_207,In_30);
nor U3205 (N_3205,In_780,In_1758);
and U3206 (N_3206,In_179,In_1010);
nand U3207 (N_3207,In_280,In_851);
nand U3208 (N_3208,In_487,In_1579);
or U3209 (N_3209,In_1821,In_403);
nor U3210 (N_3210,In_1935,In_743);
or U3211 (N_3211,In_1470,In_419);
xnor U3212 (N_3212,In_538,In_1412);
or U3213 (N_3213,In_1495,In_399);
xor U3214 (N_3214,In_1901,In_803);
nand U3215 (N_3215,In_1216,In_423);
nand U3216 (N_3216,In_992,In_778);
xnor U3217 (N_3217,In_71,In_1505);
xor U3218 (N_3218,In_764,In_1997);
and U3219 (N_3219,In_1726,In_1532);
and U3220 (N_3220,In_396,In_1037);
xor U3221 (N_3221,In_1898,In_461);
nand U3222 (N_3222,In_534,In_1874);
xnor U3223 (N_3223,In_1756,In_377);
xor U3224 (N_3224,In_985,In_988);
nand U3225 (N_3225,In_1690,In_1003);
nand U3226 (N_3226,In_1133,In_1136);
xnor U3227 (N_3227,In_73,In_1541);
nor U3228 (N_3228,In_498,In_1618);
xnor U3229 (N_3229,In_1775,In_1917);
xnor U3230 (N_3230,In_301,In_459);
and U3231 (N_3231,In_905,In_1332);
or U3232 (N_3232,In_55,In_1256);
and U3233 (N_3233,In_393,In_1303);
nand U3234 (N_3234,In_1411,In_989);
and U3235 (N_3235,In_1736,In_695);
nand U3236 (N_3236,In_1916,In_900);
xor U3237 (N_3237,In_1110,In_711);
xor U3238 (N_3238,In_476,In_51);
nor U3239 (N_3239,In_1267,In_1482);
nand U3240 (N_3240,In_1096,In_1132);
xor U3241 (N_3241,In_156,In_312);
or U3242 (N_3242,In_403,In_1666);
nor U3243 (N_3243,In_1435,In_139);
and U3244 (N_3244,In_1761,In_1873);
nor U3245 (N_3245,In_441,In_1765);
and U3246 (N_3246,In_1196,In_1297);
nand U3247 (N_3247,In_1056,In_798);
xor U3248 (N_3248,In_984,In_1807);
nor U3249 (N_3249,In_617,In_281);
nor U3250 (N_3250,In_832,In_1891);
nor U3251 (N_3251,In_895,In_82);
or U3252 (N_3252,In_1944,In_5);
and U3253 (N_3253,In_673,In_1899);
nor U3254 (N_3254,In_642,In_48);
and U3255 (N_3255,In_1256,In_454);
and U3256 (N_3256,In_809,In_1389);
or U3257 (N_3257,In_1689,In_519);
nand U3258 (N_3258,In_1308,In_546);
xnor U3259 (N_3259,In_1203,In_1288);
or U3260 (N_3260,In_871,In_695);
xor U3261 (N_3261,In_896,In_256);
and U3262 (N_3262,In_761,In_1104);
nor U3263 (N_3263,In_1305,In_252);
and U3264 (N_3264,In_759,In_1025);
and U3265 (N_3265,In_1682,In_1909);
nor U3266 (N_3266,In_3,In_1646);
nor U3267 (N_3267,In_39,In_331);
and U3268 (N_3268,In_1646,In_1098);
nor U3269 (N_3269,In_710,In_1867);
xnor U3270 (N_3270,In_245,In_1461);
or U3271 (N_3271,In_1214,In_50);
or U3272 (N_3272,In_586,In_834);
xor U3273 (N_3273,In_1555,In_1376);
or U3274 (N_3274,In_828,In_762);
xnor U3275 (N_3275,In_1415,In_1379);
nand U3276 (N_3276,In_495,In_158);
or U3277 (N_3277,In_1957,In_1780);
or U3278 (N_3278,In_742,In_1133);
nand U3279 (N_3279,In_11,In_917);
nand U3280 (N_3280,In_381,In_1266);
xnor U3281 (N_3281,In_168,In_186);
nor U3282 (N_3282,In_1389,In_205);
nand U3283 (N_3283,In_383,In_306);
nor U3284 (N_3284,In_1681,In_853);
and U3285 (N_3285,In_387,In_604);
and U3286 (N_3286,In_1282,In_1468);
or U3287 (N_3287,In_1753,In_1432);
nand U3288 (N_3288,In_1740,In_781);
nor U3289 (N_3289,In_1510,In_1647);
nor U3290 (N_3290,In_1807,In_1250);
nand U3291 (N_3291,In_1774,In_498);
xor U3292 (N_3292,In_474,In_1236);
xor U3293 (N_3293,In_1273,In_1479);
nand U3294 (N_3294,In_1466,In_668);
nand U3295 (N_3295,In_634,In_732);
or U3296 (N_3296,In_1748,In_224);
and U3297 (N_3297,In_1398,In_1044);
or U3298 (N_3298,In_1541,In_545);
or U3299 (N_3299,In_755,In_1355);
or U3300 (N_3300,In_1633,In_433);
xor U3301 (N_3301,In_983,In_452);
nand U3302 (N_3302,In_281,In_299);
or U3303 (N_3303,In_1805,In_1708);
xor U3304 (N_3304,In_981,In_1980);
and U3305 (N_3305,In_1363,In_1921);
nor U3306 (N_3306,In_38,In_1537);
nor U3307 (N_3307,In_710,In_90);
nor U3308 (N_3308,In_257,In_37);
nor U3309 (N_3309,In_1418,In_1606);
xnor U3310 (N_3310,In_1503,In_1085);
nand U3311 (N_3311,In_304,In_1026);
nand U3312 (N_3312,In_1660,In_736);
nor U3313 (N_3313,In_32,In_99);
nor U3314 (N_3314,In_1809,In_580);
xor U3315 (N_3315,In_1669,In_1647);
or U3316 (N_3316,In_691,In_1526);
xor U3317 (N_3317,In_33,In_636);
nor U3318 (N_3318,In_1232,In_788);
xor U3319 (N_3319,In_1246,In_584);
and U3320 (N_3320,In_712,In_216);
xnor U3321 (N_3321,In_1166,In_1520);
or U3322 (N_3322,In_521,In_522);
and U3323 (N_3323,In_33,In_294);
nor U3324 (N_3324,In_677,In_211);
xnor U3325 (N_3325,In_908,In_655);
xor U3326 (N_3326,In_1515,In_1146);
or U3327 (N_3327,In_1577,In_121);
nand U3328 (N_3328,In_668,In_358);
and U3329 (N_3329,In_1117,In_1918);
nand U3330 (N_3330,In_1626,In_553);
or U3331 (N_3331,In_1648,In_1128);
nand U3332 (N_3332,In_538,In_797);
and U3333 (N_3333,In_1536,In_519);
xnor U3334 (N_3334,In_1127,In_1688);
xor U3335 (N_3335,In_898,In_1576);
and U3336 (N_3336,In_1825,In_895);
nand U3337 (N_3337,In_1169,In_622);
nand U3338 (N_3338,In_35,In_1596);
nor U3339 (N_3339,In_1578,In_998);
and U3340 (N_3340,In_733,In_1931);
xor U3341 (N_3341,In_385,In_386);
xnor U3342 (N_3342,In_1930,In_527);
or U3343 (N_3343,In_1504,In_1797);
xor U3344 (N_3344,In_546,In_113);
nor U3345 (N_3345,In_1646,In_322);
nand U3346 (N_3346,In_204,In_337);
nor U3347 (N_3347,In_386,In_8);
nand U3348 (N_3348,In_1283,In_1860);
nor U3349 (N_3349,In_457,In_1770);
or U3350 (N_3350,In_1873,In_1883);
xor U3351 (N_3351,In_1737,In_391);
nand U3352 (N_3352,In_1252,In_1743);
and U3353 (N_3353,In_1747,In_424);
xor U3354 (N_3354,In_1307,In_1106);
xor U3355 (N_3355,In_1601,In_51);
and U3356 (N_3356,In_1030,In_211);
nand U3357 (N_3357,In_574,In_1547);
or U3358 (N_3358,In_572,In_1653);
xnor U3359 (N_3359,In_360,In_442);
nor U3360 (N_3360,In_661,In_1127);
nor U3361 (N_3361,In_458,In_1890);
and U3362 (N_3362,In_1997,In_793);
nand U3363 (N_3363,In_1884,In_426);
nand U3364 (N_3364,In_1843,In_1879);
or U3365 (N_3365,In_395,In_119);
or U3366 (N_3366,In_50,In_92);
xnor U3367 (N_3367,In_722,In_1409);
or U3368 (N_3368,In_851,In_1814);
xor U3369 (N_3369,In_974,In_1304);
nor U3370 (N_3370,In_246,In_953);
and U3371 (N_3371,In_64,In_973);
xor U3372 (N_3372,In_1734,In_423);
xor U3373 (N_3373,In_180,In_1793);
nand U3374 (N_3374,In_705,In_1215);
and U3375 (N_3375,In_518,In_27);
xnor U3376 (N_3376,In_251,In_494);
nor U3377 (N_3377,In_1159,In_1027);
and U3378 (N_3378,In_813,In_904);
nand U3379 (N_3379,In_1955,In_46);
nor U3380 (N_3380,In_695,In_864);
nor U3381 (N_3381,In_906,In_323);
nor U3382 (N_3382,In_1694,In_1429);
and U3383 (N_3383,In_1741,In_1747);
and U3384 (N_3384,In_1128,In_1285);
nor U3385 (N_3385,In_818,In_1776);
or U3386 (N_3386,In_810,In_1914);
xor U3387 (N_3387,In_863,In_1821);
xnor U3388 (N_3388,In_1233,In_1697);
and U3389 (N_3389,In_333,In_96);
or U3390 (N_3390,In_795,In_1816);
nor U3391 (N_3391,In_1002,In_217);
xor U3392 (N_3392,In_983,In_1223);
nor U3393 (N_3393,In_982,In_1967);
nand U3394 (N_3394,In_1180,In_1534);
nor U3395 (N_3395,In_1798,In_201);
nand U3396 (N_3396,In_1262,In_1635);
nor U3397 (N_3397,In_377,In_1169);
nand U3398 (N_3398,In_1695,In_1301);
or U3399 (N_3399,In_772,In_1700);
and U3400 (N_3400,In_775,In_813);
nand U3401 (N_3401,In_907,In_975);
nor U3402 (N_3402,In_1583,In_1791);
nor U3403 (N_3403,In_1874,In_499);
and U3404 (N_3404,In_162,In_249);
xor U3405 (N_3405,In_548,In_1982);
and U3406 (N_3406,In_773,In_1347);
xor U3407 (N_3407,In_1825,In_1045);
nor U3408 (N_3408,In_1014,In_1292);
or U3409 (N_3409,In_1155,In_669);
or U3410 (N_3410,In_1975,In_1996);
nor U3411 (N_3411,In_244,In_1898);
or U3412 (N_3412,In_474,In_1741);
nand U3413 (N_3413,In_1053,In_144);
and U3414 (N_3414,In_1525,In_1158);
xor U3415 (N_3415,In_1889,In_1486);
and U3416 (N_3416,In_1309,In_634);
nor U3417 (N_3417,In_614,In_1623);
nand U3418 (N_3418,In_1053,In_899);
nor U3419 (N_3419,In_460,In_748);
and U3420 (N_3420,In_1040,In_1158);
nand U3421 (N_3421,In_197,In_750);
or U3422 (N_3422,In_183,In_1599);
nand U3423 (N_3423,In_1110,In_1979);
or U3424 (N_3424,In_1780,In_1146);
or U3425 (N_3425,In_1641,In_611);
xor U3426 (N_3426,In_692,In_1015);
nor U3427 (N_3427,In_1099,In_617);
nand U3428 (N_3428,In_579,In_275);
nand U3429 (N_3429,In_73,In_1187);
and U3430 (N_3430,In_265,In_1913);
nor U3431 (N_3431,In_1845,In_112);
or U3432 (N_3432,In_1560,In_1173);
and U3433 (N_3433,In_1079,In_539);
or U3434 (N_3434,In_1726,In_101);
xnor U3435 (N_3435,In_735,In_1910);
nand U3436 (N_3436,In_884,In_618);
nand U3437 (N_3437,In_1669,In_921);
or U3438 (N_3438,In_1433,In_1184);
nor U3439 (N_3439,In_137,In_512);
or U3440 (N_3440,In_1423,In_1757);
nand U3441 (N_3441,In_1876,In_1810);
nand U3442 (N_3442,In_1147,In_173);
xnor U3443 (N_3443,In_1796,In_1545);
nand U3444 (N_3444,In_1664,In_707);
nor U3445 (N_3445,In_1911,In_256);
and U3446 (N_3446,In_1433,In_1764);
nor U3447 (N_3447,In_513,In_1092);
nor U3448 (N_3448,In_1438,In_713);
nand U3449 (N_3449,In_415,In_1138);
nand U3450 (N_3450,In_276,In_558);
nand U3451 (N_3451,In_1159,In_264);
and U3452 (N_3452,In_1828,In_757);
nor U3453 (N_3453,In_737,In_961);
nand U3454 (N_3454,In_1800,In_1060);
nor U3455 (N_3455,In_43,In_656);
and U3456 (N_3456,In_1673,In_477);
nand U3457 (N_3457,In_97,In_1603);
or U3458 (N_3458,In_442,In_479);
xor U3459 (N_3459,In_586,In_818);
and U3460 (N_3460,In_1289,In_1768);
nand U3461 (N_3461,In_1395,In_821);
nor U3462 (N_3462,In_1177,In_1663);
or U3463 (N_3463,In_1694,In_1203);
nand U3464 (N_3464,In_431,In_1387);
xor U3465 (N_3465,In_1263,In_1507);
nand U3466 (N_3466,In_466,In_1974);
and U3467 (N_3467,In_902,In_1624);
nand U3468 (N_3468,In_145,In_1894);
nand U3469 (N_3469,In_743,In_1151);
nor U3470 (N_3470,In_1259,In_993);
or U3471 (N_3471,In_233,In_1592);
xnor U3472 (N_3472,In_660,In_201);
and U3473 (N_3473,In_841,In_1224);
or U3474 (N_3474,In_431,In_285);
and U3475 (N_3475,In_1391,In_1625);
nor U3476 (N_3476,In_1049,In_823);
nor U3477 (N_3477,In_133,In_51);
or U3478 (N_3478,In_456,In_368);
nand U3479 (N_3479,In_609,In_555);
nor U3480 (N_3480,In_622,In_1948);
and U3481 (N_3481,In_1636,In_1706);
xnor U3482 (N_3482,In_177,In_1697);
and U3483 (N_3483,In_758,In_909);
nor U3484 (N_3484,In_771,In_630);
and U3485 (N_3485,In_1756,In_153);
nand U3486 (N_3486,In_872,In_16);
and U3487 (N_3487,In_916,In_955);
and U3488 (N_3488,In_1483,In_1919);
xor U3489 (N_3489,In_684,In_1490);
and U3490 (N_3490,In_1460,In_409);
or U3491 (N_3491,In_235,In_1295);
or U3492 (N_3492,In_1915,In_498);
nor U3493 (N_3493,In_1297,In_1806);
and U3494 (N_3494,In_1579,In_1378);
or U3495 (N_3495,In_1631,In_1990);
nand U3496 (N_3496,In_538,In_345);
or U3497 (N_3497,In_989,In_1380);
or U3498 (N_3498,In_1862,In_789);
xor U3499 (N_3499,In_1485,In_234);
xor U3500 (N_3500,In_1669,In_187);
and U3501 (N_3501,In_1921,In_460);
xor U3502 (N_3502,In_414,In_998);
nor U3503 (N_3503,In_80,In_305);
or U3504 (N_3504,In_75,In_46);
xor U3505 (N_3505,In_1794,In_753);
nor U3506 (N_3506,In_64,In_397);
or U3507 (N_3507,In_411,In_695);
and U3508 (N_3508,In_922,In_650);
nor U3509 (N_3509,In_830,In_1735);
or U3510 (N_3510,In_1408,In_40);
nor U3511 (N_3511,In_529,In_1347);
nand U3512 (N_3512,In_1053,In_1618);
nand U3513 (N_3513,In_45,In_226);
xor U3514 (N_3514,In_683,In_1202);
and U3515 (N_3515,In_1104,In_692);
nand U3516 (N_3516,In_1403,In_86);
or U3517 (N_3517,In_368,In_217);
and U3518 (N_3518,In_677,In_787);
or U3519 (N_3519,In_184,In_1893);
or U3520 (N_3520,In_1223,In_1834);
nand U3521 (N_3521,In_1518,In_1926);
nor U3522 (N_3522,In_1767,In_1879);
xor U3523 (N_3523,In_1342,In_1915);
and U3524 (N_3524,In_963,In_1130);
xnor U3525 (N_3525,In_641,In_211);
and U3526 (N_3526,In_1717,In_326);
or U3527 (N_3527,In_760,In_1305);
and U3528 (N_3528,In_1759,In_705);
xnor U3529 (N_3529,In_1620,In_694);
xnor U3530 (N_3530,In_266,In_1095);
or U3531 (N_3531,In_527,In_1221);
or U3532 (N_3532,In_1467,In_302);
nand U3533 (N_3533,In_71,In_1887);
xnor U3534 (N_3534,In_1149,In_195);
or U3535 (N_3535,In_39,In_121);
nand U3536 (N_3536,In_807,In_1047);
nor U3537 (N_3537,In_1014,In_428);
nand U3538 (N_3538,In_1481,In_1125);
nand U3539 (N_3539,In_1389,In_745);
nor U3540 (N_3540,In_942,In_619);
nand U3541 (N_3541,In_1362,In_1195);
nand U3542 (N_3542,In_239,In_1800);
xnor U3543 (N_3543,In_247,In_1378);
and U3544 (N_3544,In_176,In_1868);
or U3545 (N_3545,In_72,In_787);
and U3546 (N_3546,In_249,In_1260);
nor U3547 (N_3547,In_1878,In_1730);
nor U3548 (N_3548,In_12,In_252);
and U3549 (N_3549,In_540,In_1174);
xnor U3550 (N_3550,In_1692,In_649);
or U3551 (N_3551,In_1284,In_1239);
or U3552 (N_3552,In_1656,In_200);
nand U3553 (N_3553,In_94,In_632);
or U3554 (N_3554,In_1241,In_1283);
nand U3555 (N_3555,In_552,In_1899);
and U3556 (N_3556,In_1208,In_1141);
and U3557 (N_3557,In_1126,In_1678);
nand U3558 (N_3558,In_1846,In_1975);
nor U3559 (N_3559,In_1409,In_1146);
or U3560 (N_3560,In_1129,In_961);
nor U3561 (N_3561,In_1323,In_833);
nor U3562 (N_3562,In_769,In_1576);
xor U3563 (N_3563,In_189,In_532);
and U3564 (N_3564,In_711,In_967);
and U3565 (N_3565,In_409,In_1448);
xnor U3566 (N_3566,In_86,In_1826);
and U3567 (N_3567,In_649,In_798);
and U3568 (N_3568,In_1291,In_685);
nand U3569 (N_3569,In_639,In_1866);
or U3570 (N_3570,In_1672,In_1613);
and U3571 (N_3571,In_446,In_691);
xnor U3572 (N_3572,In_1897,In_587);
xnor U3573 (N_3573,In_4,In_971);
xor U3574 (N_3574,In_1782,In_1340);
and U3575 (N_3575,In_706,In_1982);
and U3576 (N_3576,In_8,In_1051);
xor U3577 (N_3577,In_1940,In_1572);
or U3578 (N_3578,In_991,In_1658);
or U3579 (N_3579,In_629,In_1659);
xnor U3580 (N_3580,In_32,In_1861);
xor U3581 (N_3581,In_297,In_344);
or U3582 (N_3582,In_674,In_1755);
xnor U3583 (N_3583,In_1739,In_18);
and U3584 (N_3584,In_774,In_1556);
nand U3585 (N_3585,In_828,In_1367);
nor U3586 (N_3586,In_24,In_710);
nand U3587 (N_3587,In_83,In_1536);
nand U3588 (N_3588,In_564,In_96);
and U3589 (N_3589,In_605,In_267);
nor U3590 (N_3590,In_1452,In_858);
nand U3591 (N_3591,In_1616,In_806);
xnor U3592 (N_3592,In_1345,In_325);
xor U3593 (N_3593,In_1238,In_1161);
xnor U3594 (N_3594,In_1704,In_1483);
nor U3595 (N_3595,In_1887,In_1639);
nand U3596 (N_3596,In_140,In_774);
or U3597 (N_3597,In_461,In_597);
or U3598 (N_3598,In_1709,In_1068);
or U3599 (N_3599,In_1841,In_453);
or U3600 (N_3600,In_542,In_1096);
nor U3601 (N_3601,In_154,In_715);
nand U3602 (N_3602,In_1708,In_1406);
nand U3603 (N_3603,In_1326,In_810);
or U3604 (N_3604,In_1714,In_1362);
and U3605 (N_3605,In_961,In_1472);
or U3606 (N_3606,In_1319,In_1485);
and U3607 (N_3607,In_333,In_480);
nand U3608 (N_3608,In_1387,In_1407);
nor U3609 (N_3609,In_947,In_1929);
and U3610 (N_3610,In_381,In_1806);
and U3611 (N_3611,In_130,In_753);
and U3612 (N_3612,In_1366,In_1977);
xor U3613 (N_3613,In_917,In_688);
and U3614 (N_3614,In_1908,In_420);
and U3615 (N_3615,In_1341,In_854);
or U3616 (N_3616,In_128,In_312);
xor U3617 (N_3617,In_1208,In_68);
nor U3618 (N_3618,In_1112,In_455);
or U3619 (N_3619,In_1326,In_1934);
nor U3620 (N_3620,In_47,In_970);
nor U3621 (N_3621,In_1611,In_576);
and U3622 (N_3622,In_696,In_261);
nor U3623 (N_3623,In_692,In_327);
and U3624 (N_3624,In_1100,In_210);
xnor U3625 (N_3625,In_839,In_662);
and U3626 (N_3626,In_992,In_152);
and U3627 (N_3627,In_1411,In_303);
and U3628 (N_3628,In_1738,In_555);
nor U3629 (N_3629,In_902,In_137);
or U3630 (N_3630,In_1790,In_12);
and U3631 (N_3631,In_304,In_1701);
nand U3632 (N_3632,In_1571,In_1239);
or U3633 (N_3633,In_593,In_1042);
nor U3634 (N_3634,In_963,In_1031);
xnor U3635 (N_3635,In_110,In_1097);
or U3636 (N_3636,In_1498,In_1262);
nor U3637 (N_3637,In_984,In_1606);
or U3638 (N_3638,In_954,In_829);
or U3639 (N_3639,In_190,In_1703);
or U3640 (N_3640,In_406,In_1544);
nand U3641 (N_3641,In_1363,In_1578);
nand U3642 (N_3642,In_1248,In_721);
xnor U3643 (N_3643,In_223,In_1004);
nor U3644 (N_3644,In_723,In_1134);
xnor U3645 (N_3645,In_1707,In_1646);
and U3646 (N_3646,In_1693,In_1272);
and U3647 (N_3647,In_747,In_918);
or U3648 (N_3648,In_1113,In_18);
nand U3649 (N_3649,In_1905,In_736);
nor U3650 (N_3650,In_1705,In_417);
or U3651 (N_3651,In_1070,In_739);
nand U3652 (N_3652,In_1191,In_1419);
and U3653 (N_3653,In_1877,In_32);
or U3654 (N_3654,In_432,In_1925);
nand U3655 (N_3655,In_1673,In_256);
nand U3656 (N_3656,In_211,In_526);
or U3657 (N_3657,In_1122,In_305);
nor U3658 (N_3658,In_833,In_995);
or U3659 (N_3659,In_735,In_1362);
nand U3660 (N_3660,In_1010,In_1819);
nand U3661 (N_3661,In_612,In_502);
nor U3662 (N_3662,In_1086,In_1455);
and U3663 (N_3663,In_618,In_786);
xor U3664 (N_3664,In_1539,In_1913);
xor U3665 (N_3665,In_1180,In_774);
or U3666 (N_3666,In_1924,In_789);
nand U3667 (N_3667,In_676,In_607);
nor U3668 (N_3668,In_931,In_922);
nor U3669 (N_3669,In_720,In_1604);
and U3670 (N_3670,In_755,In_1425);
nand U3671 (N_3671,In_352,In_1000);
nor U3672 (N_3672,In_1043,In_393);
nand U3673 (N_3673,In_931,In_1249);
or U3674 (N_3674,In_308,In_1878);
and U3675 (N_3675,In_1466,In_462);
nor U3676 (N_3676,In_1988,In_836);
nor U3677 (N_3677,In_1657,In_208);
or U3678 (N_3678,In_1903,In_1379);
nor U3679 (N_3679,In_354,In_331);
or U3680 (N_3680,In_1357,In_756);
nor U3681 (N_3681,In_1813,In_1643);
and U3682 (N_3682,In_436,In_1306);
xnor U3683 (N_3683,In_187,In_109);
nor U3684 (N_3684,In_1423,In_1149);
xnor U3685 (N_3685,In_1247,In_590);
and U3686 (N_3686,In_1228,In_1004);
or U3687 (N_3687,In_967,In_1916);
or U3688 (N_3688,In_1311,In_1586);
and U3689 (N_3689,In_1844,In_1189);
or U3690 (N_3690,In_1011,In_1992);
or U3691 (N_3691,In_909,In_1473);
xor U3692 (N_3692,In_1873,In_659);
or U3693 (N_3693,In_1603,In_1804);
nand U3694 (N_3694,In_1291,In_768);
and U3695 (N_3695,In_1464,In_1730);
or U3696 (N_3696,In_156,In_799);
nor U3697 (N_3697,In_1010,In_1323);
xor U3698 (N_3698,In_1436,In_800);
or U3699 (N_3699,In_440,In_93);
nand U3700 (N_3700,In_1154,In_970);
nor U3701 (N_3701,In_329,In_1811);
and U3702 (N_3702,In_1623,In_1925);
or U3703 (N_3703,In_1358,In_1461);
nand U3704 (N_3704,In_1417,In_354);
xnor U3705 (N_3705,In_962,In_837);
or U3706 (N_3706,In_638,In_209);
and U3707 (N_3707,In_252,In_982);
or U3708 (N_3708,In_588,In_1126);
nor U3709 (N_3709,In_534,In_241);
and U3710 (N_3710,In_478,In_1176);
nor U3711 (N_3711,In_523,In_1469);
nor U3712 (N_3712,In_381,In_124);
nand U3713 (N_3713,In_1461,In_1341);
xnor U3714 (N_3714,In_1463,In_1866);
or U3715 (N_3715,In_1998,In_248);
xor U3716 (N_3716,In_1116,In_1024);
nand U3717 (N_3717,In_1587,In_791);
or U3718 (N_3718,In_146,In_1720);
xnor U3719 (N_3719,In_223,In_906);
xor U3720 (N_3720,In_1342,In_193);
nor U3721 (N_3721,In_1448,In_1254);
nor U3722 (N_3722,In_1326,In_219);
and U3723 (N_3723,In_1434,In_742);
and U3724 (N_3724,In_571,In_1583);
nand U3725 (N_3725,In_1648,In_1476);
xnor U3726 (N_3726,In_784,In_880);
xnor U3727 (N_3727,In_1465,In_1874);
or U3728 (N_3728,In_398,In_741);
or U3729 (N_3729,In_514,In_409);
and U3730 (N_3730,In_1185,In_1119);
and U3731 (N_3731,In_78,In_819);
nand U3732 (N_3732,In_908,In_1884);
or U3733 (N_3733,In_1022,In_1728);
nor U3734 (N_3734,In_1142,In_1921);
or U3735 (N_3735,In_1519,In_571);
or U3736 (N_3736,In_702,In_1720);
xnor U3737 (N_3737,In_344,In_168);
or U3738 (N_3738,In_1361,In_558);
and U3739 (N_3739,In_1094,In_1380);
xnor U3740 (N_3740,In_1201,In_1391);
or U3741 (N_3741,In_409,In_584);
xor U3742 (N_3742,In_344,In_1751);
xor U3743 (N_3743,In_930,In_1671);
or U3744 (N_3744,In_1555,In_506);
and U3745 (N_3745,In_1740,In_24);
or U3746 (N_3746,In_1483,In_1345);
or U3747 (N_3747,In_736,In_1688);
nand U3748 (N_3748,In_206,In_1165);
xnor U3749 (N_3749,In_1523,In_169);
and U3750 (N_3750,In_715,In_1020);
and U3751 (N_3751,In_40,In_1577);
xor U3752 (N_3752,In_809,In_1595);
nand U3753 (N_3753,In_1621,In_453);
or U3754 (N_3754,In_1301,In_421);
or U3755 (N_3755,In_1194,In_1249);
xnor U3756 (N_3756,In_1046,In_925);
and U3757 (N_3757,In_1555,In_263);
nor U3758 (N_3758,In_60,In_360);
or U3759 (N_3759,In_133,In_214);
or U3760 (N_3760,In_1713,In_1434);
nand U3761 (N_3761,In_675,In_1577);
nand U3762 (N_3762,In_428,In_109);
and U3763 (N_3763,In_387,In_1554);
xor U3764 (N_3764,In_1103,In_210);
nor U3765 (N_3765,In_734,In_1067);
nor U3766 (N_3766,In_1705,In_920);
and U3767 (N_3767,In_1527,In_1757);
or U3768 (N_3768,In_891,In_1679);
xnor U3769 (N_3769,In_1710,In_1074);
nand U3770 (N_3770,In_192,In_1448);
xor U3771 (N_3771,In_1369,In_1837);
nor U3772 (N_3772,In_111,In_1976);
and U3773 (N_3773,In_1808,In_1518);
or U3774 (N_3774,In_1076,In_1669);
xor U3775 (N_3775,In_756,In_156);
xnor U3776 (N_3776,In_482,In_713);
nand U3777 (N_3777,In_382,In_844);
and U3778 (N_3778,In_305,In_1476);
xor U3779 (N_3779,In_564,In_332);
xor U3780 (N_3780,In_4,In_1467);
xnor U3781 (N_3781,In_1291,In_217);
nand U3782 (N_3782,In_1525,In_1399);
and U3783 (N_3783,In_1736,In_534);
and U3784 (N_3784,In_1099,In_1968);
xor U3785 (N_3785,In_1424,In_1347);
or U3786 (N_3786,In_1923,In_1469);
xnor U3787 (N_3787,In_83,In_349);
xor U3788 (N_3788,In_1384,In_1217);
xor U3789 (N_3789,In_1374,In_1606);
or U3790 (N_3790,In_1191,In_1712);
or U3791 (N_3791,In_1648,In_502);
nor U3792 (N_3792,In_1191,In_1135);
or U3793 (N_3793,In_1198,In_1028);
or U3794 (N_3794,In_1743,In_848);
and U3795 (N_3795,In_1554,In_1682);
nor U3796 (N_3796,In_65,In_1194);
and U3797 (N_3797,In_988,In_1872);
or U3798 (N_3798,In_1488,In_1191);
and U3799 (N_3799,In_1936,In_1719);
nand U3800 (N_3800,In_1117,In_1870);
nor U3801 (N_3801,In_1136,In_1012);
nor U3802 (N_3802,In_1757,In_1316);
nor U3803 (N_3803,In_958,In_1788);
xnor U3804 (N_3804,In_463,In_1991);
nand U3805 (N_3805,In_154,In_1704);
or U3806 (N_3806,In_903,In_1982);
nor U3807 (N_3807,In_665,In_965);
xnor U3808 (N_3808,In_357,In_1082);
nand U3809 (N_3809,In_99,In_559);
nand U3810 (N_3810,In_1398,In_1847);
nand U3811 (N_3811,In_1591,In_1676);
and U3812 (N_3812,In_1748,In_1328);
and U3813 (N_3813,In_1245,In_4);
xnor U3814 (N_3814,In_44,In_1527);
or U3815 (N_3815,In_352,In_714);
or U3816 (N_3816,In_803,In_477);
nor U3817 (N_3817,In_936,In_284);
xnor U3818 (N_3818,In_1529,In_926);
xnor U3819 (N_3819,In_935,In_835);
nand U3820 (N_3820,In_951,In_1790);
xnor U3821 (N_3821,In_307,In_163);
nand U3822 (N_3822,In_1351,In_1664);
nor U3823 (N_3823,In_208,In_1107);
nand U3824 (N_3824,In_905,In_1571);
or U3825 (N_3825,In_1850,In_404);
or U3826 (N_3826,In_1492,In_341);
nor U3827 (N_3827,In_1173,In_98);
nor U3828 (N_3828,In_1192,In_1602);
nand U3829 (N_3829,In_417,In_1399);
xnor U3830 (N_3830,In_1586,In_873);
xor U3831 (N_3831,In_636,In_1597);
nor U3832 (N_3832,In_163,In_1054);
nand U3833 (N_3833,In_348,In_480);
nand U3834 (N_3834,In_640,In_1690);
and U3835 (N_3835,In_1166,In_1325);
or U3836 (N_3836,In_1117,In_1720);
and U3837 (N_3837,In_553,In_377);
and U3838 (N_3838,In_1570,In_691);
nand U3839 (N_3839,In_1883,In_427);
nand U3840 (N_3840,In_1946,In_0);
or U3841 (N_3841,In_1793,In_1678);
nor U3842 (N_3842,In_1707,In_1126);
and U3843 (N_3843,In_1169,In_1211);
nor U3844 (N_3844,In_1669,In_785);
and U3845 (N_3845,In_1968,In_1550);
and U3846 (N_3846,In_1654,In_113);
xor U3847 (N_3847,In_1523,In_313);
and U3848 (N_3848,In_225,In_874);
nor U3849 (N_3849,In_42,In_963);
xor U3850 (N_3850,In_796,In_113);
nand U3851 (N_3851,In_80,In_721);
nor U3852 (N_3852,In_907,In_903);
or U3853 (N_3853,In_1297,In_1914);
or U3854 (N_3854,In_166,In_235);
or U3855 (N_3855,In_122,In_1221);
and U3856 (N_3856,In_388,In_607);
nand U3857 (N_3857,In_1113,In_433);
and U3858 (N_3858,In_1891,In_1695);
xnor U3859 (N_3859,In_214,In_577);
nand U3860 (N_3860,In_435,In_1820);
nor U3861 (N_3861,In_585,In_1039);
xor U3862 (N_3862,In_661,In_355);
nand U3863 (N_3863,In_387,In_1501);
nor U3864 (N_3864,In_441,In_1441);
and U3865 (N_3865,In_93,In_624);
and U3866 (N_3866,In_620,In_938);
and U3867 (N_3867,In_173,In_736);
and U3868 (N_3868,In_1531,In_1540);
or U3869 (N_3869,In_1006,In_1836);
and U3870 (N_3870,In_1845,In_670);
xor U3871 (N_3871,In_1844,In_1437);
or U3872 (N_3872,In_510,In_877);
or U3873 (N_3873,In_1250,In_502);
nor U3874 (N_3874,In_1596,In_836);
nand U3875 (N_3875,In_1732,In_1215);
and U3876 (N_3876,In_824,In_614);
xor U3877 (N_3877,In_756,In_544);
nor U3878 (N_3878,In_1851,In_528);
and U3879 (N_3879,In_1173,In_1587);
nand U3880 (N_3880,In_1367,In_1244);
or U3881 (N_3881,In_880,In_1596);
and U3882 (N_3882,In_1314,In_822);
nand U3883 (N_3883,In_1298,In_1915);
and U3884 (N_3884,In_1248,In_772);
xor U3885 (N_3885,In_665,In_1647);
nand U3886 (N_3886,In_834,In_184);
xnor U3887 (N_3887,In_778,In_1163);
and U3888 (N_3888,In_1029,In_1297);
xor U3889 (N_3889,In_1361,In_1312);
xnor U3890 (N_3890,In_312,In_587);
nor U3891 (N_3891,In_986,In_839);
xor U3892 (N_3892,In_245,In_1012);
and U3893 (N_3893,In_402,In_265);
and U3894 (N_3894,In_510,In_944);
or U3895 (N_3895,In_978,In_1980);
or U3896 (N_3896,In_826,In_1444);
nand U3897 (N_3897,In_221,In_1487);
nor U3898 (N_3898,In_1266,In_610);
xor U3899 (N_3899,In_430,In_213);
nor U3900 (N_3900,In_1186,In_687);
or U3901 (N_3901,In_956,In_821);
or U3902 (N_3902,In_1179,In_607);
or U3903 (N_3903,In_765,In_882);
or U3904 (N_3904,In_392,In_1637);
and U3905 (N_3905,In_1212,In_1650);
xnor U3906 (N_3906,In_828,In_1940);
or U3907 (N_3907,In_1776,In_1006);
xor U3908 (N_3908,In_1634,In_716);
or U3909 (N_3909,In_749,In_1012);
or U3910 (N_3910,In_59,In_141);
or U3911 (N_3911,In_1809,In_382);
nand U3912 (N_3912,In_361,In_425);
xnor U3913 (N_3913,In_1785,In_1072);
and U3914 (N_3914,In_1286,In_804);
xor U3915 (N_3915,In_1573,In_1012);
nand U3916 (N_3916,In_1928,In_1111);
nand U3917 (N_3917,In_689,In_160);
nor U3918 (N_3918,In_899,In_931);
and U3919 (N_3919,In_432,In_417);
and U3920 (N_3920,In_496,In_700);
xor U3921 (N_3921,In_1708,In_79);
nand U3922 (N_3922,In_393,In_1780);
nand U3923 (N_3923,In_1642,In_382);
or U3924 (N_3924,In_937,In_68);
nand U3925 (N_3925,In_103,In_263);
and U3926 (N_3926,In_1806,In_940);
nand U3927 (N_3927,In_870,In_148);
and U3928 (N_3928,In_371,In_1167);
xnor U3929 (N_3929,In_524,In_1039);
nor U3930 (N_3930,In_1278,In_497);
nor U3931 (N_3931,In_1455,In_1026);
xor U3932 (N_3932,In_1783,In_151);
nor U3933 (N_3933,In_1286,In_1094);
xor U3934 (N_3934,In_657,In_1165);
and U3935 (N_3935,In_1046,In_1938);
or U3936 (N_3936,In_1525,In_1354);
nand U3937 (N_3937,In_1376,In_1291);
nor U3938 (N_3938,In_1181,In_1756);
nor U3939 (N_3939,In_1688,In_937);
nor U3940 (N_3940,In_1313,In_178);
or U3941 (N_3941,In_1335,In_1110);
nand U3942 (N_3942,In_1313,In_403);
and U3943 (N_3943,In_1086,In_1085);
nor U3944 (N_3944,In_683,In_22);
nand U3945 (N_3945,In_571,In_1260);
and U3946 (N_3946,In_144,In_583);
nor U3947 (N_3947,In_242,In_1741);
xor U3948 (N_3948,In_674,In_1701);
nand U3949 (N_3949,In_255,In_545);
nor U3950 (N_3950,In_1153,In_1464);
or U3951 (N_3951,In_292,In_742);
and U3952 (N_3952,In_840,In_339);
nand U3953 (N_3953,In_1813,In_1635);
nor U3954 (N_3954,In_1376,In_744);
nand U3955 (N_3955,In_210,In_466);
nand U3956 (N_3956,In_256,In_238);
nand U3957 (N_3957,In_1557,In_1378);
nand U3958 (N_3958,In_459,In_626);
nor U3959 (N_3959,In_1352,In_1693);
nor U3960 (N_3960,In_94,In_1038);
or U3961 (N_3961,In_579,In_1254);
nand U3962 (N_3962,In_1648,In_103);
nand U3963 (N_3963,In_1096,In_622);
xnor U3964 (N_3964,In_184,In_1471);
and U3965 (N_3965,In_1724,In_602);
and U3966 (N_3966,In_72,In_813);
nor U3967 (N_3967,In_1730,In_216);
nor U3968 (N_3968,In_311,In_52);
xnor U3969 (N_3969,In_559,In_1980);
nor U3970 (N_3970,In_1697,In_1175);
and U3971 (N_3971,In_695,In_653);
nor U3972 (N_3972,In_1736,In_1498);
xnor U3973 (N_3973,In_1009,In_1068);
xor U3974 (N_3974,In_864,In_915);
or U3975 (N_3975,In_837,In_1698);
and U3976 (N_3976,In_974,In_1718);
xor U3977 (N_3977,In_178,In_755);
xnor U3978 (N_3978,In_187,In_1535);
nand U3979 (N_3979,In_1362,In_780);
or U3980 (N_3980,In_148,In_1231);
nor U3981 (N_3981,In_1467,In_734);
xnor U3982 (N_3982,In_1039,In_590);
and U3983 (N_3983,In_1095,In_1536);
xor U3984 (N_3984,In_989,In_979);
nand U3985 (N_3985,In_1199,In_1379);
xor U3986 (N_3986,In_1439,In_353);
nor U3987 (N_3987,In_499,In_1598);
nand U3988 (N_3988,In_1180,In_1799);
and U3989 (N_3989,In_61,In_453);
and U3990 (N_3990,In_1635,In_664);
xor U3991 (N_3991,In_1148,In_680);
or U3992 (N_3992,In_1302,In_1797);
nor U3993 (N_3993,In_1809,In_644);
and U3994 (N_3994,In_325,In_1303);
or U3995 (N_3995,In_355,In_218);
xnor U3996 (N_3996,In_1673,In_759);
nor U3997 (N_3997,In_1935,In_1787);
nor U3998 (N_3998,In_264,In_1295);
xnor U3999 (N_3999,In_258,In_709);
xnor U4000 (N_4000,In_1596,In_1125);
and U4001 (N_4001,In_472,In_405);
xor U4002 (N_4002,In_645,In_1993);
and U4003 (N_4003,In_958,In_477);
and U4004 (N_4004,In_143,In_1738);
or U4005 (N_4005,In_861,In_1607);
nor U4006 (N_4006,In_461,In_1778);
xnor U4007 (N_4007,In_1335,In_426);
nor U4008 (N_4008,In_1587,In_1821);
nor U4009 (N_4009,In_1633,In_326);
xor U4010 (N_4010,In_606,In_1381);
nor U4011 (N_4011,In_1746,In_961);
and U4012 (N_4012,In_1101,In_805);
nor U4013 (N_4013,In_1901,In_1068);
xnor U4014 (N_4014,In_1706,In_697);
xor U4015 (N_4015,In_1875,In_1753);
nor U4016 (N_4016,In_684,In_1506);
nor U4017 (N_4017,In_219,In_491);
and U4018 (N_4018,In_745,In_1813);
and U4019 (N_4019,In_1412,In_374);
nand U4020 (N_4020,In_317,In_694);
xnor U4021 (N_4021,In_1637,In_231);
or U4022 (N_4022,In_1764,In_326);
nor U4023 (N_4023,In_389,In_1504);
or U4024 (N_4024,In_182,In_1044);
nor U4025 (N_4025,In_996,In_1431);
xnor U4026 (N_4026,In_918,In_145);
xnor U4027 (N_4027,In_621,In_52);
or U4028 (N_4028,In_1323,In_607);
nor U4029 (N_4029,In_1657,In_20);
and U4030 (N_4030,In_1808,In_1793);
nor U4031 (N_4031,In_829,In_226);
xnor U4032 (N_4032,In_1229,In_1176);
nor U4033 (N_4033,In_110,In_1153);
and U4034 (N_4034,In_767,In_912);
xnor U4035 (N_4035,In_628,In_892);
and U4036 (N_4036,In_848,In_998);
nor U4037 (N_4037,In_699,In_996);
nor U4038 (N_4038,In_687,In_1420);
nand U4039 (N_4039,In_623,In_1958);
and U4040 (N_4040,In_600,In_103);
nand U4041 (N_4041,In_908,In_205);
nand U4042 (N_4042,In_1912,In_1725);
and U4043 (N_4043,In_678,In_1124);
or U4044 (N_4044,In_679,In_492);
or U4045 (N_4045,In_1234,In_1073);
or U4046 (N_4046,In_643,In_978);
and U4047 (N_4047,In_78,In_1589);
or U4048 (N_4048,In_1604,In_737);
xor U4049 (N_4049,In_535,In_1485);
xnor U4050 (N_4050,In_1519,In_930);
and U4051 (N_4051,In_402,In_1353);
nand U4052 (N_4052,In_1461,In_1063);
nor U4053 (N_4053,In_989,In_94);
and U4054 (N_4054,In_1312,In_1020);
and U4055 (N_4055,In_681,In_235);
and U4056 (N_4056,In_1037,In_1289);
xor U4057 (N_4057,In_304,In_846);
nor U4058 (N_4058,In_173,In_632);
nand U4059 (N_4059,In_1248,In_389);
and U4060 (N_4060,In_367,In_1694);
nor U4061 (N_4061,In_1977,In_79);
nand U4062 (N_4062,In_1948,In_1836);
nand U4063 (N_4063,In_1720,In_591);
and U4064 (N_4064,In_979,In_408);
nor U4065 (N_4065,In_1054,In_807);
and U4066 (N_4066,In_1429,In_1436);
or U4067 (N_4067,In_1275,In_31);
nand U4068 (N_4068,In_338,In_863);
nor U4069 (N_4069,In_1295,In_435);
xor U4070 (N_4070,In_1677,In_1326);
and U4071 (N_4071,In_1413,In_521);
nand U4072 (N_4072,In_838,In_1562);
nor U4073 (N_4073,In_782,In_147);
nor U4074 (N_4074,In_818,In_831);
nand U4075 (N_4075,In_1071,In_1974);
nand U4076 (N_4076,In_567,In_430);
xnor U4077 (N_4077,In_500,In_512);
nand U4078 (N_4078,In_78,In_1300);
nand U4079 (N_4079,In_1339,In_42);
and U4080 (N_4080,In_1636,In_259);
and U4081 (N_4081,In_325,In_1088);
nand U4082 (N_4082,In_1919,In_1777);
and U4083 (N_4083,In_691,In_546);
or U4084 (N_4084,In_468,In_917);
nor U4085 (N_4085,In_258,In_1822);
nor U4086 (N_4086,In_1294,In_429);
nor U4087 (N_4087,In_52,In_1568);
nor U4088 (N_4088,In_1191,In_1270);
and U4089 (N_4089,In_538,In_668);
nand U4090 (N_4090,In_1905,In_179);
or U4091 (N_4091,In_101,In_419);
or U4092 (N_4092,In_1477,In_1313);
nor U4093 (N_4093,In_968,In_810);
or U4094 (N_4094,In_1973,In_1426);
and U4095 (N_4095,In_1947,In_1477);
xnor U4096 (N_4096,In_1745,In_1657);
or U4097 (N_4097,In_1254,In_1370);
nand U4098 (N_4098,In_1568,In_579);
and U4099 (N_4099,In_143,In_825);
nand U4100 (N_4100,In_1974,In_1723);
and U4101 (N_4101,In_1562,In_400);
xor U4102 (N_4102,In_515,In_1968);
nor U4103 (N_4103,In_1270,In_645);
and U4104 (N_4104,In_739,In_922);
xor U4105 (N_4105,In_1651,In_704);
xnor U4106 (N_4106,In_1734,In_1271);
and U4107 (N_4107,In_1342,In_47);
nand U4108 (N_4108,In_1503,In_1597);
nand U4109 (N_4109,In_776,In_633);
xnor U4110 (N_4110,In_1330,In_1557);
and U4111 (N_4111,In_91,In_909);
nand U4112 (N_4112,In_1728,In_1360);
and U4113 (N_4113,In_1490,In_1557);
nand U4114 (N_4114,In_1498,In_791);
nor U4115 (N_4115,In_1075,In_1331);
nand U4116 (N_4116,In_614,In_1178);
nand U4117 (N_4117,In_1808,In_97);
nor U4118 (N_4118,In_1840,In_1524);
nor U4119 (N_4119,In_706,In_771);
nand U4120 (N_4120,In_1257,In_1348);
and U4121 (N_4121,In_1143,In_231);
nand U4122 (N_4122,In_1805,In_1640);
nor U4123 (N_4123,In_469,In_676);
nand U4124 (N_4124,In_1888,In_1881);
xor U4125 (N_4125,In_827,In_313);
nand U4126 (N_4126,In_25,In_348);
and U4127 (N_4127,In_1030,In_829);
xnor U4128 (N_4128,In_1616,In_627);
or U4129 (N_4129,In_1764,In_1117);
xnor U4130 (N_4130,In_371,In_328);
and U4131 (N_4131,In_1482,In_1117);
xnor U4132 (N_4132,In_1065,In_466);
xor U4133 (N_4133,In_637,In_1770);
or U4134 (N_4134,In_479,In_1623);
nand U4135 (N_4135,In_817,In_440);
and U4136 (N_4136,In_787,In_916);
and U4137 (N_4137,In_576,In_1195);
nor U4138 (N_4138,In_1878,In_1792);
nor U4139 (N_4139,In_517,In_1936);
or U4140 (N_4140,In_1394,In_1537);
or U4141 (N_4141,In_1187,In_1682);
nor U4142 (N_4142,In_795,In_33);
nand U4143 (N_4143,In_1667,In_1456);
nand U4144 (N_4144,In_0,In_276);
nor U4145 (N_4145,In_406,In_503);
and U4146 (N_4146,In_14,In_160);
xor U4147 (N_4147,In_70,In_955);
or U4148 (N_4148,In_1010,In_835);
nor U4149 (N_4149,In_193,In_1722);
and U4150 (N_4150,In_476,In_1431);
nor U4151 (N_4151,In_1936,In_487);
and U4152 (N_4152,In_1867,In_627);
or U4153 (N_4153,In_106,In_705);
xnor U4154 (N_4154,In_253,In_1464);
nor U4155 (N_4155,In_1004,In_412);
or U4156 (N_4156,In_1420,In_44);
nor U4157 (N_4157,In_930,In_952);
xor U4158 (N_4158,In_1150,In_1028);
nor U4159 (N_4159,In_1648,In_1936);
or U4160 (N_4160,In_1221,In_1341);
xnor U4161 (N_4161,In_532,In_1773);
or U4162 (N_4162,In_1987,In_811);
xnor U4163 (N_4163,In_1584,In_1382);
nand U4164 (N_4164,In_1345,In_1239);
nor U4165 (N_4165,In_1444,In_1230);
nor U4166 (N_4166,In_1571,In_497);
nand U4167 (N_4167,In_1389,In_604);
nand U4168 (N_4168,In_1110,In_391);
nand U4169 (N_4169,In_1294,In_1306);
xnor U4170 (N_4170,In_1315,In_956);
and U4171 (N_4171,In_465,In_1609);
nand U4172 (N_4172,In_117,In_1367);
xnor U4173 (N_4173,In_1167,In_1974);
nor U4174 (N_4174,In_135,In_75);
or U4175 (N_4175,In_1410,In_1635);
xnor U4176 (N_4176,In_842,In_550);
or U4177 (N_4177,In_1515,In_1493);
xor U4178 (N_4178,In_1237,In_948);
nand U4179 (N_4179,In_458,In_1076);
nand U4180 (N_4180,In_70,In_608);
nor U4181 (N_4181,In_761,In_1627);
nor U4182 (N_4182,In_914,In_98);
nor U4183 (N_4183,In_1916,In_920);
or U4184 (N_4184,In_304,In_870);
xnor U4185 (N_4185,In_176,In_1754);
xor U4186 (N_4186,In_1465,In_576);
nor U4187 (N_4187,In_1381,In_959);
xnor U4188 (N_4188,In_303,In_1605);
nor U4189 (N_4189,In_1264,In_1633);
xnor U4190 (N_4190,In_1431,In_1467);
nor U4191 (N_4191,In_685,In_1897);
xor U4192 (N_4192,In_1066,In_1569);
and U4193 (N_4193,In_455,In_1377);
nand U4194 (N_4194,In_448,In_1255);
nand U4195 (N_4195,In_328,In_408);
or U4196 (N_4196,In_1155,In_1158);
nor U4197 (N_4197,In_1424,In_464);
and U4198 (N_4198,In_934,In_821);
xnor U4199 (N_4199,In_833,In_1344);
and U4200 (N_4200,In_234,In_496);
xnor U4201 (N_4201,In_53,In_1991);
xor U4202 (N_4202,In_1960,In_1669);
and U4203 (N_4203,In_721,In_123);
or U4204 (N_4204,In_1226,In_75);
and U4205 (N_4205,In_177,In_1808);
nand U4206 (N_4206,In_632,In_956);
nor U4207 (N_4207,In_1576,In_1956);
nor U4208 (N_4208,In_1951,In_1614);
and U4209 (N_4209,In_990,In_1027);
xnor U4210 (N_4210,In_402,In_835);
nand U4211 (N_4211,In_1564,In_1191);
xnor U4212 (N_4212,In_1008,In_740);
nand U4213 (N_4213,In_1146,In_1774);
and U4214 (N_4214,In_882,In_581);
or U4215 (N_4215,In_261,In_1477);
xor U4216 (N_4216,In_431,In_789);
nor U4217 (N_4217,In_982,In_1395);
nor U4218 (N_4218,In_1700,In_1797);
xor U4219 (N_4219,In_1490,In_1347);
and U4220 (N_4220,In_440,In_497);
xnor U4221 (N_4221,In_1793,In_749);
xor U4222 (N_4222,In_951,In_1986);
xnor U4223 (N_4223,In_999,In_376);
xnor U4224 (N_4224,In_1089,In_979);
or U4225 (N_4225,In_990,In_1451);
and U4226 (N_4226,In_1913,In_528);
and U4227 (N_4227,In_1375,In_1717);
nand U4228 (N_4228,In_156,In_893);
nand U4229 (N_4229,In_482,In_16);
and U4230 (N_4230,In_1563,In_197);
xnor U4231 (N_4231,In_905,In_512);
nor U4232 (N_4232,In_1895,In_1614);
nand U4233 (N_4233,In_268,In_550);
xnor U4234 (N_4234,In_56,In_996);
or U4235 (N_4235,In_1474,In_81);
nor U4236 (N_4236,In_175,In_645);
or U4237 (N_4237,In_1864,In_189);
xor U4238 (N_4238,In_554,In_1797);
nor U4239 (N_4239,In_1017,In_1961);
xor U4240 (N_4240,In_1285,In_106);
and U4241 (N_4241,In_1203,In_48);
or U4242 (N_4242,In_813,In_551);
nor U4243 (N_4243,In_808,In_1354);
xnor U4244 (N_4244,In_910,In_1851);
and U4245 (N_4245,In_321,In_574);
and U4246 (N_4246,In_356,In_452);
nand U4247 (N_4247,In_70,In_1430);
nand U4248 (N_4248,In_1277,In_1411);
or U4249 (N_4249,In_1328,In_1116);
nor U4250 (N_4250,In_799,In_1476);
xor U4251 (N_4251,In_1495,In_689);
and U4252 (N_4252,In_1847,In_1342);
nor U4253 (N_4253,In_548,In_615);
nor U4254 (N_4254,In_206,In_857);
nand U4255 (N_4255,In_1297,In_1);
nand U4256 (N_4256,In_1284,In_607);
or U4257 (N_4257,In_1573,In_1015);
nand U4258 (N_4258,In_1046,In_501);
and U4259 (N_4259,In_569,In_691);
nor U4260 (N_4260,In_138,In_27);
and U4261 (N_4261,In_200,In_671);
and U4262 (N_4262,In_405,In_160);
or U4263 (N_4263,In_1268,In_989);
and U4264 (N_4264,In_246,In_1854);
and U4265 (N_4265,In_1266,In_324);
and U4266 (N_4266,In_688,In_1063);
xor U4267 (N_4267,In_1548,In_1269);
xor U4268 (N_4268,In_1018,In_690);
nor U4269 (N_4269,In_801,In_1350);
and U4270 (N_4270,In_1260,In_1689);
and U4271 (N_4271,In_189,In_1878);
nand U4272 (N_4272,In_602,In_429);
nor U4273 (N_4273,In_831,In_1794);
xor U4274 (N_4274,In_109,In_349);
xor U4275 (N_4275,In_1778,In_425);
and U4276 (N_4276,In_848,In_1252);
nand U4277 (N_4277,In_1061,In_843);
nor U4278 (N_4278,In_638,In_6);
nor U4279 (N_4279,In_1551,In_1885);
or U4280 (N_4280,In_1068,In_876);
or U4281 (N_4281,In_157,In_1163);
and U4282 (N_4282,In_1143,In_1810);
xnor U4283 (N_4283,In_906,In_1387);
and U4284 (N_4284,In_1788,In_887);
or U4285 (N_4285,In_584,In_1326);
xor U4286 (N_4286,In_1458,In_208);
or U4287 (N_4287,In_1037,In_193);
xor U4288 (N_4288,In_110,In_1422);
nor U4289 (N_4289,In_1341,In_1248);
xor U4290 (N_4290,In_455,In_1407);
nand U4291 (N_4291,In_1163,In_140);
nor U4292 (N_4292,In_1333,In_509);
nor U4293 (N_4293,In_365,In_1667);
nor U4294 (N_4294,In_767,In_1776);
nor U4295 (N_4295,In_1098,In_1937);
nor U4296 (N_4296,In_1322,In_1182);
and U4297 (N_4297,In_25,In_1943);
nand U4298 (N_4298,In_62,In_1667);
or U4299 (N_4299,In_799,In_1481);
nand U4300 (N_4300,In_1785,In_454);
and U4301 (N_4301,In_768,In_454);
and U4302 (N_4302,In_1120,In_435);
and U4303 (N_4303,In_21,In_1295);
nand U4304 (N_4304,In_24,In_1108);
or U4305 (N_4305,In_263,In_266);
or U4306 (N_4306,In_896,In_386);
xnor U4307 (N_4307,In_1644,In_348);
and U4308 (N_4308,In_464,In_1250);
nand U4309 (N_4309,In_811,In_432);
xor U4310 (N_4310,In_1373,In_121);
nand U4311 (N_4311,In_158,In_996);
nor U4312 (N_4312,In_335,In_539);
or U4313 (N_4313,In_1946,In_971);
or U4314 (N_4314,In_1049,In_1979);
and U4315 (N_4315,In_1257,In_452);
and U4316 (N_4316,In_1267,In_651);
and U4317 (N_4317,In_1230,In_706);
or U4318 (N_4318,In_1564,In_329);
nand U4319 (N_4319,In_1558,In_559);
and U4320 (N_4320,In_836,In_1615);
nand U4321 (N_4321,In_1108,In_748);
nand U4322 (N_4322,In_1519,In_1563);
or U4323 (N_4323,In_1403,In_90);
and U4324 (N_4324,In_976,In_1023);
nand U4325 (N_4325,In_883,In_1023);
nor U4326 (N_4326,In_1638,In_997);
nand U4327 (N_4327,In_152,In_1230);
nand U4328 (N_4328,In_1334,In_702);
nor U4329 (N_4329,In_876,In_1594);
xor U4330 (N_4330,In_462,In_473);
nand U4331 (N_4331,In_941,In_499);
xor U4332 (N_4332,In_531,In_695);
or U4333 (N_4333,In_1981,In_1586);
nand U4334 (N_4334,In_1596,In_174);
nor U4335 (N_4335,In_508,In_905);
or U4336 (N_4336,In_854,In_384);
and U4337 (N_4337,In_165,In_932);
nor U4338 (N_4338,In_1956,In_1933);
and U4339 (N_4339,In_1283,In_1076);
nor U4340 (N_4340,In_430,In_1664);
nor U4341 (N_4341,In_181,In_175);
nand U4342 (N_4342,In_1622,In_1675);
nand U4343 (N_4343,In_214,In_1175);
and U4344 (N_4344,In_212,In_1819);
and U4345 (N_4345,In_1572,In_963);
nand U4346 (N_4346,In_317,In_493);
or U4347 (N_4347,In_570,In_422);
and U4348 (N_4348,In_1327,In_1940);
and U4349 (N_4349,In_740,In_1637);
xor U4350 (N_4350,In_111,In_96);
nand U4351 (N_4351,In_1851,In_1823);
xor U4352 (N_4352,In_297,In_229);
nor U4353 (N_4353,In_889,In_513);
and U4354 (N_4354,In_1582,In_165);
nand U4355 (N_4355,In_1824,In_1326);
xnor U4356 (N_4356,In_1842,In_1125);
nor U4357 (N_4357,In_1434,In_300);
nand U4358 (N_4358,In_1095,In_1387);
nand U4359 (N_4359,In_405,In_408);
nand U4360 (N_4360,In_1864,In_1135);
nor U4361 (N_4361,In_1415,In_1370);
and U4362 (N_4362,In_1986,In_753);
and U4363 (N_4363,In_784,In_1635);
nand U4364 (N_4364,In_606,In_1988);
and U4365 (N_4365,In_577,In_1333);
nor U4366 (N_4366,In_1451,In_1862);
xnor U4367 (N_4367,In_994,In_542);
and U4368 (N_4368,In_549,In_1511);
nor U4369 (N_4369,In_943,In_1108);
nand U4370 (N_4370,In_1344,In_277);
nand U4371 (N_4371,In_1566,In_1401);
nor U4372 (N_4372,In_796,In_1264);
or U4373 (N_4373,In_1535,In_511);
and U4374 (N_4374,In_1912,In_1275);
and U4375 (N_4375,In_121,In_1339);
nand U4376 (N_4376,In_239,In_426);
and U4377 (N_4377,In_1425,In_1680);
nor U4378 (N_4378,In_1590,In_128);
xnor U4379 (N_4379,In_1023,In_677);
and U4380 (N_4380,In_588,In_641);
nor U4381 (N_4381,In_982,In_236);
nand U4382 (N_4382,In_1000,In_1118);
nor U4383 (N_4383,In_593,In_1664);
nor U4384 (N_4384,In_916,In_1159);
or U4385 (N_4385,In_1167,In_640);
nor U4386 (N_4386,In_1516,In_1223);
or U4387 (N_4387,In_1377,In_365);
nand U4388 (N_4388,In_1753,In_1593);
xnor U4389 (N_4389,In_295,In_237);
xor U4390 (N_4390,In_809,In_1832);
nor U4391 (N_4391,In_1814,In_324);
or U4392 (N_4392,In_1480,In_1724);
nor U4393 (N_4393,In_488,In_1158);
nand U4394 (N_4394,In_1221,In_196);
nand U4395 (N_4395,In_504,In_726);
nor U4396 (N_4396,In_942,In_407);
or U4397 (N_4397,In_1481,In_869);
nor U4398 (N_4398,In_1387,In_1484);
nor U4399 (N_4399,In_607,In_1053);
or U4400 (N_4400,In_111,In_1995);
and U4401 (N_4401,In_586,In_1432);
xnor U4402 (N_4402,In_1602,In_715);
nand U4403 (N_4403,In_1192,In_725);
nand U4404 (N_4404,In_917,In_1508);
nand U4405 (N_4405,In_1388,In_1489);
and U4406 (N_4406,In_1379,In_1601);
xnor U4407 (N_4407,In_489,In_1421);
nor U4408 (N_4408,In_1351,In_89);
nand U4409 (N_4409,In_1285,In_1025);
and U4410 (N_4410,In_1078,In_204);
nor U4411 (N_4411,In_124,In_1099);
xor U4412 (N_4412,In_513,In_1813);
nor U4413 (N_4413,In_1675,In_1767);
nor U4414 (N_4414,In_1342,In_1711);
and U4415 (N_4415,In_664,In_780);
nor U4416 (N_4416,In_594,In_306);
nand U4417 (N_4417,In_1324,In_125);
xor U4418 (N_4418,In_1600,In_164);
xor U4419 (N_4419,In_984,In_602);
xnor U4420 (N_4420,In_54,In_520);
nor U4421 (N_4421,In_18,In_1761);
xnor U4422 (N_4422,In_855,In_506);
nand U4423 (N_4423,In_1251,In_1964);
nor U4424 (N_4424,In_1696,In_699);
and U4425 (N_4425,In_486,In_1880);
nand U4426 (N_4426,In_1863,In_1091);
xor U4427 (N_4427,In_823,In_600);
xor U4428 (N_4428,In_921,In_1161);
and U4429 (N_4429,In_391,In_1401);
nand U4430 (N_4430,In_1023,In_1774);
and U4431 (N_4431,In_540,In_1843);
or U4432 (N_4432,In_980,In_261);
nor U4433 (N_4433,In_29,In_1160);
and U4434 (N_4434,In_383,In_1842);
xnor U4435 (N_4435,In_1066,In_1268);
or U4436 (N_4436,In_1848,In_1658);
and U4437 (N_4437,In_531,In_1545);
nor U4438 (N_4438,In_1783,In_281);
nor U4439 (N_4439,In_942,In_507);
xnor U4440 (N_4440,In_1917,In_1621);
xnor U4441 (N_4441,In_1860,In_1425);
nor U4442 (N_4442,In_615,In_1020);
or U4443 (N_4443,In_266,In_1476);
nor U4444 (N_4444,In_1658,In_1494);
and U4445 (N_4445,In_1552,In_876);
or U4446 (N_4446,In_1199,In_1821);
nor U4447 (N_4447,In_332,In_1576);
nor U4448 (N_4448,In_1213,In_1334);
xnor U4449 (N_4449,In_258,In_1771);
nor U4450 (N_4450,In_460,In_1798);
nor U4451 (N_4451,In_1264,In_1660);
or U4452 (N_4452,In_641,In_1721);
xor U4453 (N_4453,In_1433,In_569);
xnor U4454 (N_4454,In_1712,In_393);
xnor U4455 (N_4455,In_1452,In_1377);
and U4456 (N_4456,In_1223,In_461);
and U4457 (N_4457,In_1253,In_607);
nand U4458 (N_4458,In_1796,In_1703);
nand U4459 (N_4459,In_382,In_205);
or U4460 (N_4460,In_715,In_1115);
or U4461 (N_4461,In_650,In_821);
nor U4462 (N_4462,In_510,In_716);
xnor U4463 (N_4463,In_54,In_973);
and U4464 (N_4464,In_123,In_727);
or U4465 (N_4465,In_1655,In_1135);
xor U4466 (N_4466,In_690,In_1160);
and U4467 (N_4467,In_1598,In_298);
xor U4468 (N_4468,In_1815,In_1916);
xnor U4469 (N_4469,In_1330,In_995);
nor U4470 (N_4470,In_566,In_1056);
nor U4471 (N_4471,In_232,In_968);
and U4472 (N_4472,In_1604,In_105);
nor U4473 (N_4473,In_1149,In_1938);
and U4474 (N_4474,In_1574,In_494);
xnor U4475 (N_4475,In_1067,In_1552);
and U4476 (N_4476,In_550,In_1753);
and U4477 (N_4477,In_984,In_1920);
nor U4478 (N_4478,In_235,In_1911);
or U4479 (N_4479,In_1999,In_664);
or U4480 (N_4480,In_91,In_528);
nor U4481 (N_4481,In_526,In_604);
and U4482 (N_4482,In_265,In_503);
nor U4483 (N_4483,In_1058,In_164);
nor U4484 (N_4484,In_1974,In_1769);
or U4485 (N_4485,In_1002,In_214);
nand U4486 (N_4486,In_281,In_205);
and U4487 (N_4487,In_373,In_1878);
xor U4488 (N_4488,In_1751,In_76);
xor U4489 (N_4489,In_895,In_1749);
nor U4490 (N_4490,In_543,In_43);
or U4491 (N_4491,In_1653,In_119);
and U4492 (N_4492,In_1872,In_1067);
nor U4493 (N_4493,In_574,In_1422);
nand U4494 (N_4494,In_1933,In_1360);
nor U4495 (N_4495,In_225,In_1947);
and U4496 (N_4496,In_173,In_1887);
nand U4497 (N_4497,In_1838,In_1310);
and U4498 (N_4498,In_365,In_450);
xor U4499 (N_4499,In_805,In_553);
xor U4500 (N_4500,In_976,In_670);
nand U4501 (N_4501,In_457,In_612);
nor U4502 (N_4502,In_1679,In_1627);
nor U4503 (N_4503,In_160,In_1731);
xor U4504 (N_4504,In_585,In_71);
and U4505 (N_4505,In_952,In_339);
nand U4506 (N_4506,In_730,In_1266);
and U4507 (N_4507,In_214,In_1244);
nand U4508 (N_4508,In_234,In_1046);
xnor U4509 (N_4509,In_1070,In_1772);
nand U4510 (N_4510,In_1371,In_794);
and U4511 (N_4511,In_175,In_1652);
nand U4512 (N_4512,In_956,In_1604);
nand U4513 (N_4513,In_855,In_1801);
nand U4514 (N_4514,In_1307,In_757);
and U4515 (N_4515,In_1510,In_203);
nand U4516 (N_4516,In_1580,In_1790);
or U4517 (N_4517,In_505,In_1563);
and U4518 (N_4518,In_1690,In_1943);
or U4519 (N_4519,In_734,In_132);
nand U4520 (N_4520,In_1317,In_1729);
nor U4521 (N_4521,In_249,In_1142);
and U4522 (N_4522,In_1670,In_432);
or U4523 (N_4523,In_1103,In_626);
and U4524 (N_4524,In_71,In_1923);
or U4525 (N_4525,In_1246,In_532);
nor U4526 (N_4526,In_940,In_477);
nand U4527 (N_4527,In_1957,In_1342);
or U4528 (N_4528,In_1960,In_1484);
and U4529 (N_4529,In_1587,In_1538);
nand U4530 (N_4530,In_1125,In_435);
nand U4531 (N_4531,In_911,In_412);
or U4532 (N_4532,In_1535,In_189);
or U4533 (N_4533,In_1865,In_47);
nand U4534 (N_4534,In_877,In_333);
or U4535 (N_4535,In_596,In_1096);
nor U4536 (N_4536,In_371,In_508);
xor U4537 (N_4537,In_1251,In_649);
or U4538 (N_4538,In_120,In_1986);
nor U4539 (N_4539,In_92,In_674);
nor U4540 (N_4540,In_1384,In_1433);
nand U4541 (N_4541,In_668,In_409);
nor U4542 (N_4542,In_494,In_1017);
nand U4543 (N_4543,In_1634,In_1859);
nor U4544 (N_4544,In_1054,In_1770);
nor U4545 (N_4545,In_1240,In_1511);
nand U4546 (N_4546,In_1956,In_569);
xor U4547 (N_4547,In_481,In_654);
or U4548 (N_4548,In_436,In_1211);
nand U4549 (N_4549,In_676,In_1855);
and U4550 (N_4550,In_1433,In_543);
nor U4551 (N_4551,In_1999,In_61);
nand U4552 (N_4552,In_479,In_1424);
xor U4553 (N_4553,In_687,In_1406);
nor U4554 (N_4554,In_496,In_760);
nor U4555 (N_4555,In_862,In_1006);
nor U4556 (N_4556,In_1082,In_884);
nand U4557 (N_4557,In_148,In_1020);
and U4558 (N_4558,In_1208,In_1415);
nand U4559 (N_4559,In_424,In_31);
nand U4560 (N_4560,In_1561,In_893);
nand U4561 (N_4561,In_541,In_1314);
and U4562 (N_4562,In_429,In_667);
nand U4563 (N_4563,In_1721,In_1078);
nand U4564 (N_4564,In_1925,In_450);
nand U4565 (N_4565,In_927,In_511);
nor U4566 (N_4566,In_1891,In_783);
and U4567 (N_4567,In_195,In_1805);
or U4568 (N_4568,In_1485,In_346);
or U4569 (N_4569,In_1047,In_819);
nor U4570 (N_4570,In_848,In_1174);
nor U4571 (N_4571,In_731,In_1676);
xor U4572 (N_4572,In_1745,In_741);
and U4573 (N_4573,In_5,In_1876);
nand U4574 (N_4574,In_1559,In_793);
nand U4575 (N_4575,In_1438,In_1997);
and U4576 (N_4576,In_1762,In_1101);
nor U4577 (N_4577,In_6,In_1289);
nor U4578 (N_4578,In_157,In_208);
xnor U4579 (N_4579,In_1992,In_1038);
xor U4580 (N_4580,In_1655,In_1883);
and U4581 (N_4581,In_1852,In_700);
nor U4582 (N_4582,In_692,In_313);
or U4583 (N_4583,In_902,In_1350);
or U4584 (N_4584,In_450,In_1427);
nor U4585 (N_4585,In_914,In_1825);
or U4586 (N_4586,In_1350,In_745);
and U4587 (N_4587,In_1783,In_493);
or U4588 (N_4588,In_1802,In_158);
xor U4589 (N_4589,In_1482,In_349);
xnor U4590 (N_4590,In_1537,In_1);
nor U4591 (N_4591,In_1084,In_1418);
or U4592 (N_4592,In_1558,In_807);
or U4593 (N_4593,In_1605,In_1941);
or U4594 (N_4594,In_1290,In_508);
nor U4595 (N_4595,In_921,In_1364);
or U4596 (N_4596,In_552,In_5);
xor U4597 (N_4597,In_189,In_984);
or U4598 (N_4598,In_1820,In_604);
nand U4599 (N_4599,In_220,In_477);
nor U4600 (N_4600,In_1297,In_1641);
xnor U4601 (N_4601,In_1207,In_1534);
or U4602 (N_4602,In_1175,In_849);
nand U4603 (N_4603,In_794,In_1380);
or U4604 (N_4604,In_889,In_1819);
nand U4605 (N_4605,In_196,In_1504);
or U4606 (N_4606,In_503,In_921);
nor U4607 (N_4607,In_800,In_859);
nor U4608 (N_4608,In_1057,In_1601);
and U4609 (N_4609,In_1292,In_670);
nand U4610 (N_4610,In_596,In_367);
nor U4611 (N_4611,In_464,In_1995);
nor U4612 (N_4612,In_1539,In_618);
or U4613 (N_4613,In_808,In_1522);
nand U4614 (N_4614,In_1222,In_885);
nor U4615 (N_4615,In_1600,In_1900);
nor U4616 (N_4616,In_471,In_321);
xor U4617 (N_4617,In_1151,In_1948);
nor U4618 (N_4618,In_1740,In_1078);
nor U4619 (N_4619,In_1758,In_319);
nand U4620 (N_4620,In_649,In_1391);
nor U4621 (N_4621,In_268,In_1824);
and U4622 (N_4622,In_1711,In_401);
and U4623 (N_4623,In_917,In_606);
or U4624 (N_4624,In_905,In_1283);
nand U4625 (N_4625,In_367,In_1382);
xor U4626 (N_4626,In_790,In_1337);
nor U4627 (N_4627,In_96,In_1972);
and U4628 (N_4628,In_1891,In_414);
and U4629 (N_4629,In_665,In_1962);
or U4630 (N_4630,In_1362,In_1402);
nor U4631 (N_4631,In_129,In_749);
nand U4632 (N_4632,In_507,In_765);
or U4633 (N_4633,In_1606,In_1121);
nor U4634 (N_4634,In_934,In_179);
nor U4635 (N_4635,In_126,In_1063);
nor U4636 (N_4636,In_487,In_335);
nor U4637 (N_4637,In_1555,In_1379);
and U4638 (N_4638,In_1447,In_1857);
nand U4639 (N_4639,In_1014,In_1844);
or U4640 (N_4640,In_1330,In_472);
xor U4641 (N_4641,In_1962,In_979);
nor U4642 (N_4642,In_819,In_612);
and U4643 (N_4643,In_1342,In_101);
nand U4644 (N_4644,In_911,In_1754);
nand U4645 (N_4645,In_1666,In_1701);
nor U4646 (N_4646,In_1049,In_474);
nand U4647 (N_4647,In_1118,In_1656);
nor U4648 (N_4648,In_667,In_1062);
or U4649 (N_4649,In_1553,In_1334);
nand U4650 (N_4650,In_792,In_1333);
xor U4651 (N_4651,In_672,In_1715);
or U4652 (N_4652,In_1029,In_740);
xnor U4653 (N_4653,In_432,In_1413);
nor U4654 (N_4654,In_1209,In_733);
nand U4655 (N_4655,In_1452,In_1772);
nor U4656 (N_4656,In_170,In_266);
nand U4657 (N_4657,In_1374,In_684);
and U4658 (N_4658,In_1302,In_1207);
nand U4659 (N_4659,In_1867,In_179);
xor U4660 (N_4660,In_1357,In_25);
nor U4661 (N_4661,In_1732,In_1186);
and U4662 (N_4662,In_1842,In_65);
nor U4663 (N_4663,In_500,In_1337);
nand U4664 (N_4664,In_1350,In_1851);
nor U4665 (N_4665,In_382,In_588);
or U4666 (N_4666,In_1120,In_742);
or U4667 (N_4667,In_316,In_390);
or U4668 (N_4668,In_414,In_1987);
xor U4669 (N_4669,In_672,In_391);
or U4670 (N_4670,In_145,In_103);
and U4671 (N_4671,In_970,In_845);
or U4672 (N_4672,In_1821,In_1080);
xor U4673 (N_4673,In_1183,In_905);
nand U4674 (N_4674,In_384,In_1293);
nor U4675 (N_4675,In_1680,In_1479);
or U4676 (N_4676,In_1221,In_519);
and U4677 (N_4677,In_857,In_1429);
xor U4678 (N_4678,In_987,In_1443);
nor U4679 (N_4679,In_1968,In_565);
and U4680 (N_4680,In_1014,In_843);
xnor U4681 (N_4681,In_1652,In_104);
and U4682 (N_4682,In_1045,In_644);
and U4683 (N_4683,In_1007,In_1131);
and U4684 (N_4684,In_1009,In_450);
nand U4685 (N_4685,In_1093,In_913);
nor U4686 (N_4686,In_1710,In_1238);
and U4687 (N_4687,In_1017,In_1511);
nor U4688 (N_4688,In_1514,In_23);
xor U4689 (N_4689,In_1127,In_902);
or U4690 (N_4690,In_1224,In_398);
nor U4691 (N_4691,In_1833,In_116);
or U4692 (N_4692,In_1117,In_575);
and U4693 (N_4693,In_332,In_1152);
xor U4694 (N_4694,In_970,In_251);
xnor U4695 (N_4695,In_1818,In_466);
xnor U4696 (N_4696,In_75,In_1167);
xnor U4697 (N_4697,In_1733,In_1852);
or U4698 (N_4698,In_1614,In_994);
and U4699 (N_4699,In_1740,In_777);
nor U4700 (N_4700,In_995,In_1598);
or U4701 (N_4701,In_1249,In_954);
nor U4702 (N_4702,In_1609,In_1428);
and U4703 (N_4703,In_1047,In_975);
nand U4704 (N_4704,In_820,In_960);
nor U4705 (N_4705,In_8,In_1063);
nand U4706 (N_4706,In_1787,In_936);
and U4707 (N_4707,In_15,In_1929);
xor U4708 (N_4708,In_1355,In_1614);
and U4709 (N_4709,In_649,In_63);
or U4710 (N_4710,In_1168,In_1908);
nand U4711 (N_4711,In_1216,In_149);
nand U4712 (N_4712,In_392,In_604);
nand U4713 (N_4713,In_1084,In_1747);
or U4714 (N_4714,In_957,In_1458);
nor U4715 (N_4715,In_520,In_388);
nor U4716 (N_4716,In_1588,In_334);
xor U4717 (N_4717,In_1061,In_652);
nor U4718 (N_4718,In_868,In_330);
and U4719 (N_4719,In_1345,In_319);
xnor U4720 (N_4720,In_388,In_1249);
or U4721 (N_4721,In_1870,In_600);
and U4722 (N_4722,In_551,In_1579);
xor U4723 (N_4723,In_1442,In_937);
or U4724 (N_4724,In_737,In_1999);
nor U4725 (N_4725,In_1719,In_410);
nor U4726 (N_4726,In_1282,In_529);
or U4727 (N_4727,In_185,In_255);
or U4728 (N_4728,In_1173,In_1663);
nand U4729 (N_4729,In_631,In_1752);
nor U4730 (N_4730,In_854,In_1831);
and U4731 (N_4731,In_1459,In_1116);
nand U4732 (N_4732,In_1047,In_1426);
nor U4733 (N_4733,In_1140,In_1846);
xor U4734 (N_4734,In_20,In_854);
and U4735 (N_4735,In_1010,In_780);
nand U4736 (N_4736,In_1665,In_1446);
nand U4737 (N_4737,In_481,In_537);
xnor U4738 (N_4738,In_897,In_1445);
xnor U4739 (N_4739,In_1247,In_14);
or U4740 (N_4740,In_940,In_1321);
and U4741 (N_4741,In_916,In_765);
xor U4742 (N_4742,In_1515,In_1806);
nor U4743 (N_4743,In_1325,In_1269);
or U4744 (N_4744,In_807,In_1768);
nor U4745 (N_4745,In_2,In_385);
nand U4746 (N_4746,In_1543,In_1929);
xor U4747 (N_4747,In_1154,In_100);
nand U4748 (N_4748,In_1563,In_657);
and U4749 (N_4749,In_234,In_1821);
nand U4750 (N_4750,In_1033,In_1905);
and U4751 (N_4751,In_1260,In_1660);
nor U4752 (N_4752,In_1461,In_1129);
xor U4753 (N_4753,In_528,In_1143);
xnor U4754 (N_4754,In_1976,In_863);
nor U4755 (N_4755,In_765,In_566);
nand U4756 (N_4756,In_912,In_402);
and U4757 (N_4757,In_391,In_1832);
nand U4758 (N_4758,In_412,In_345);
and U4759 (N_4759,In_188,In_361);
and U4760 (N_4760,In_1932,In_1679);
nor U4761 (N_4761,In_1331,In_344);
nor U4762 (N_4762,In_367,In_1437);
or U4763 (N_4763,In_1585,In_1944);
or U4764 (N_4764,In_212,In_1845);
or U4765 (N_4765,In_789,In_1375);
and U4766 (N_4766,In_1663,In_960);
nor U4767 (N_4767,In_34,In_2);
xnor U4768 (N_4768,In_131,In_1248);
or U4769 (N_4769,In_627,In_767);
nand U4770 (N_4770,In_1798,In_1456);
nor U4771 (N_4771,In_119,In_1966);
or U4772 (N_4772,In_1245,In_956);
xor U4773 (N_4773,In_560,In_218);
nand U4774 (N_4774,In_934,In_361);
nor U4775 (N_4775,In_1680,In_597);
xnor U4776 (N_4776,In_1619,In_1979);
and U4777 (N_4777,In_1804,In_704);
and U4778 (N_4778,In_708,In_296);
and U4779 (N_4779,In_253,In_1941);
xnor U4780 (N_4780,In_1232,In_880);
nor U4781 (N_4781,In_157,In_1896);
nor U4782 (N_4782,In_1659,In_1771);
xor U4783 (N_4783,In_416,In_6);
nand U4784 (N_4784,In_789,In_1641);
nand U4785 (N_4785,In_600,In_1800);
nor U4786 (N_4786,In_889,In_1327);
or U4787 (N_4787,In_415,In_655);
xor U4788 (N_4788,In_1927,In_1946);
xnor U4789 (N_4789,In_1044,In_764);
nor U4790 (N_4790,In_158,In_670);
nand U4791 (N_4791,In_1084,In_1256);
nand U4792 (N_4792,In_888,In_1358);
or U4793 (N_4793,In_1714,In_188);
or U4794 (N_4794,In_1347,In_1827);
and U4795 (N_4795,In_1686,In_671);
and U4796 (N_4796,In_1272,In_1772);
nor U4797 (N_4797,In_1044,In_1425);
xor U4798 (N_4798,In_1530,In_439);
xnor U4799 (N_4799,In_863,In_1307);
nand U4800 (N_4800,In_388,In_1379);
xnor U4801 (N_4801,In_585,In_211);
nand U4802 (N_4802,In_1000,In_1525);
xnor U4803 (N_4803,In_414,In_712);
xor U4804 (N_4804,In_1476,In_1275);
or U4805 (N_4805,In_538,In_20);
and U4806 (N_4806,In_1867,In_449);
nand U4807 (N_4807,In_886,In_1975);
nand U4808 (N_4808,In_1130,In_438);
or U4809 (N_4809,In_870,In_1383);
and U4810 (N_4810,In_555,In_1538);
nand U4811 (N_4811,In_1396,In_275);
nor U4812 (N_4812,In_1539,In_1662);
nor U4813 (N_4813,In_1368,In_1753);
or U4814 (N_4814,In_263,In_1715);
nor U4815 (N_4815,In_962,In_697);
or U4816 (N_4816,In_1623,In_954);
and U4817 (N_4817,In_506,In_872);
nor U4818 (N_4818,In_522,In_610);
and U4819 (N_4819,In_1579,In_1585);
nand U4820 (N_4820,In_1597,In_657);
xnor U4821 (N_4821,In_1822,In_429);
xnor U4822 (N_4822,In_1863,In_316);
nand U4823 (N_4823,In_1718,In_1675);
nand U4824 (N_4824,In_1132,In_385);
nand U4825 (N_4825,In_156,In_839);
xor U4826 (N_4826,In_1314,In_411);
nand U4827 (N_4827,In_1644,In_67);
nor U4828 (N_4828,In_1579,In_1991);
and U4829 (N_4829,In_493,In_1743);
or U4830 (N_4830,In_418,In_157);
or U4831 (N_4831,In_1778,In_1179);
nor U4832 (N_4832,In_1475,In_474);
and U4833 (N_4833,In_395,In_852);
and U4834 (N_4834,In_817,In_897);
and U4835 (N_4835,In_1921,In_251);
and U4836 (N_4836,In_1166,In_406);
nand U4837 (N_4837,In_156,In_1054);
and U4838 (N_4838,In_1717,In_403);
nand U4839 (N_4839,In_539,In_1189);
xnor U4840 (N_4840,In_1222,In_273);
or U4841 (N_4841,In_1159,In_509);
xor U4842 (N_4842,In_428,In_1716);
nor U4843 (N_4843,In_921,In_1052);
nand U4844 (N_4844,In_576,In_192);
nand U4845 (N_4845,In_655,In_1670);
xnor U4846 (N_4846,In_472,In_558);
nor U4847 (N_4847,In_1973,In_1440);
xor U4848 (N_4848,In_171,In_599);
or U4849 (N_4849,In_729,In_747);
xor U4850 (N_4850,In_409,In_114);
or U4851 (N_4851,In_1240,In_534);
nand U4852 (N_4852,In_621,In_1316);
and U4853 (N_4853,In_1164,In_559);
and U4854 (N_4854,In_780,In_1757);
xor U4855 (N_4855,In_365,In_1741);
xor U4856 (N_4856,In_578,In_1056);
xnor U4857 (N_4857,In_825,In_751);
xnor U4858 (N_4858,In_567,In_1520);
nand U4859 (N_4859,In_95,In_1994);
or U4860 (N_4860,In_1058,In_1633);
nor U4861 (N_4861,In_1079,In_1789);
and U4862 (N_4862,In_323,In_1709);
nand U4863 (N_4863,In_370,In_756);
or U4864 (N_4864,In_678,In_1829);
xor U4865 (N_4865,In_450,In_1874);
nor U4866 (N_4866,In_1401,In_1538);
xnor U4867 (N_4867,In_666,In_120);
xnor U4868 (N_4868,In_357,In_1567);
nand U4869 (N_4869,In_863,In_427);
xor U4870 (N_4870,In_14,In_1535);
nand U4871 (N_4871,In_1536,In_513);
xor U4872 (N_4872,In_1285,In_1394);
xor U4873 (N_4873,In_307,In_1687);
and U4874 (N_4874,In_1870,In_937);
nor U4875 (N_4875,In_1486,In_1456);
nand U4876 (N_4876,In_610,In_954);
or U4877 (N_4877,In_1997,In_642);
nand U4878 (N_4878,In_1863,In_1142);
nor U4879 (N_4879,In_303,In_1689);
nand U4880 (N_4880,In_730,In_734);
xor U4881 (N_4881,In_1514,In_509);
nor U4882 (N_4882,In_1752,In_1111);
nand U4883 (N_4883,In_72,In_1903);
nand U4884 (N_4884,In_787,In_1911);
and U4885 (N_4885,In_625,In_1437);
nor U4886 (N_4886,In_1237,In_38);
xnor U4887 (N_4887,In_1109,In_1374);
and U4888 (N_4888,In_1279,In_218);
or U4889 (N_4889,In_181,In_1879);
and U4890 (N_4890,In_944,In_1383);
xor U4891 (N_4891,In_1427,In_1118);
and U4892 (N_4892,In_614,In_341);
nor U4893 (N_4893,In_1381,In_1474);
nor U4894 (N_4894,In_1199,In_1589);
nor U4895 (N_4895,In_1919,In_1115);
nand U4896 (N_4896,In_408,In_217);
or U4897 (N_4897,In_911,In_1766);
or U4898 (N_4898,In_445,In_1492);
nor U4899 (N_4899,In_1586,In_1565);
xor U4900 (N_4900,In_1255,In_526);
nand U4901 (N_4901,In_939,In_945);
and U4902 (N_4902,In_1465,In_1199);
nand U4903 (N_4903,In_125,In_335);
xnor U4904 (N_4904,In_1751,In_1846);
nor U4905 (N_4905,In_249,In_175);
or U4906 (N_4906,In_1504,In_599);
nand U4907 (N_4907,In_1079,In_300);
nor U4908 (N_4908,In_225,In_883);
or U4909 (N_4909,In_763,In_1745);
xnor U4910 (N_4910,In_1228,In_162);
and U4911 (N_4911,In_266,In_430);
or U4912 (N_4912,In_1332,In_817);
xnor U4913 (N_4913,In_1047,In_811);
and U4914 (N_4914,In_709,In_1206);
nor U4915 (N_4915,In_1932,In_1515);
xnor U4916 (N_4916,In_421,In_1007);
xnor U4917 (N_4917,In_232,In_1031);
xnor U4918 (N_4918,In_981,In_159);
nand U4919 (N_4919,In_1672,In_1709);
xor U4920 (N_4920,In_531,In_383);
nand U4921 (N_4921,In_402,In_476);
nand U4922 (N_4922,In_756,In_1168);
nor U4923 (N_4923,In_1993,In_750);
or U4924 (N_4924,In_636,In_1565);
xnor U4925 (N_4925,In_1605,In_601);
nor U4926 (N_4926,In_1695,In_990);
and U4927 (N_4927,In_80,In_1293);
or U4928 (N_4928,In_507,In_542);
and U4929 (N_4929,In_175,In_1997);
nor U4930 (N_4930,In_1929,In_1791);
or U4931 (N_4931,In_40,In_1841);
xor U4932 (N_4932,In_318,In_303);
and U4933 (N_4933,In_696,In_912);
or U4934 (N_4934,In_555,In_304);
xnor U4935 (N_4935,In_1777,In_1515);
or U4936 (N_4936,In_950,In_741);
and U4937 (N_4937,In_661,In_1997);
nor U4938 (N_4938,In_1733,In_298);
and U4939 (N_4939,In_1568,In_673);
and U4940 (N_4940,In_153,In_1183);
nor U4941 (N_4941,In_626,In_1270);
nor U4942 (N_4942,In_1980,In_277);
nand U4943 (N_4943,In_1958,In_1923);
nor U4944 (N_4944,In_1059,In_1801);
or U4945 (N_4945,In_894,In_1760);
nor U4946 (N_4946,In_787,In_1626);
or U4947 (N_4947,In_1550,In_985);
and U4948 (N_4948,In_766,In_626);
nand U4949 (N_4949,In_1507,In_1336);
or U4950 (N_4950,In_1287,In_707);
nor U4951 (N_4951,In_180,In_837);
nor U4952 (N_4952,In_733,In_1300);
xnor U4953 (N_4953,In_770,In_1523);
xnor U4954 (N_4954,In_1541,In_980);
nand U4955 (N_4955,In_1022,In_1176);
nor U4956 (N_4956,In_65,In_673);
xor U4957 (N_4957,In_1137,In_1739);
and U4958 (N_4958,In_850,In_1884);
nor U4959 (N_4959,In_1525,In_1978);
or U4960 (N_4960,In_76,In_655);
nor U4961 (N_4961,In_1847,In_1079);
xnor U4962 (N_4962,In_371,In_0);
nor U4963 (N_4963,In_466,In_172);
xor U4964 (N_4964,In_407,In_361);
and U4965 (N_4965,In_683,In_607);
nand U4966 (N_4966,In_1640,In_811);
xor U4967 (N_4967,In_1244,In_939);
and U4968 (N_4968,In_561,In_376);
or U4969 (N_4969,In_1073,In_1862);
nand U4970 (N_4970,In_508,In_263);
and U4971 (N_4971,In_1950,In_230);
and U4972 (N_4972,In_1266,In_573);
and U4973 (N_4973,In_1395,In_252);
nor U4974 (N_4974,In_936,In_245);
or U4975 (N_4975,In_343,In_305);
or U4976 (N_4976,In_860,In_628);
xnor U4977 (N_4977,In_478,In_19);
or U4978 (N_4978,In_418,In_244);
or U4979 (N_4979,In_1694,In_1320);
nand U4980 (N_4980,In_1435,In_690);
and U4981 (N_4981,In_269,In_106);
nand U4982 (N_4982,In_1305,In_1029);
and U4983 (N_4983,In_1455,In_297);
and U4984 (N_4984,In_1375,In_1942);
xor U4985 (N_4985,In_1140,In_62);
or U4986 (N_4986,In_906,In_1078);
nand U4987 (N_4987,In_1337,In_1831);
and U4988 (N_4988,In_1901,In_398);
or U4989 (N_4989,In_1450,In_691);
and U4990 (N_4990,In_1496,In_1823);
nor U4991 (N_4991,In_987,In_1284);
nand U4992 (N_4992,In_1408,In_1981);
nor U4993 (N_4993,In_1815,In_985);
or U4994 (N_4994,In_1655,In_443);
and U4995 (N_4995,In_1970,In_1875);
and U4996 (N_4996,In_1450,In_491);
nand U4997 (N_4997,In_860,In_1020);
nor U4998 (N_4998,In_1021,In_875);
nand U4999 (N_4999,In_1814,In_1570);
or U5000 (N_5000,N_4170,N_431);
nor U5001 (N_5001,N_3497,N_1079);
nor U5002 (N_5002,N_2978,N_2321);
nand U5003 (N_5003,N_3225,N_1092);
or U5004 (N_5004,N_442,N_2749);
nand U5005 (N_5005,N_4969,N_530);
nand U5006 (N_5006,N_3244,N_2435);
and U5007 (N_5007,N_4756,N_10);
nor U5008 (N_5008,N_1971,N_3793);
nand U5009 (N_5009,N_1852,N_856);
or U5010 (N_5010,N_1800,N_4165);
and U5011 (N_5011,N_1633,N_1065);
and U5012 (N_5012,N_4568,N_4493);
nor U5013 (N_5013,N_3481,N_443);
xnor U5014 (N_5014,N_4611,N_4628);
nor U5015 (N_5015,N_1774,N_4403);
nand U5016 (N_5016,N_4179,N_1562);
nand U5017 (N_5017,N_2482,N_733);
xor U5018 (N_5018,N_4952,N_191);
nand U5019 (N_5019,N_3183,N_2948);
and U5020 (N_5020,N_3102,N_368);
xnor U5021 (N_5021,N_2272,N_727);
nor U5022 (N_5022,N_2357,N_4050);
nor U5023 (N_5023,N_2368,N_2082);
and U5024 (N_5024,N_1843,N_627);
nor U5025 (N_5025,N_2198,N_1297);
or U5026 (N_5026,N_3799,N_3174);
and U5027 (N_5027,N_4779,N_3919);
xnor U5028 (N_5028,N_2625,N_285);
nand U5029 (N_5029,N_3095,N_2028);
nand U5030 (N_5030,N_3062,N_3554);
and U5031 (N_5031,N_2349,N_444);
xor U5032 (N_5032,N_3956,N_470);
and U5033 (N_5033,N_228,N_1049);
or U5034 (N_5034,N_3840,N_1306);
nand U5035 (N_5035,N_4956,N_2493);
nor U5036 (N_5036,N_4178,N_1036);
xor U5037 (N_5037,N_2745,N_1788);
or U5038 (N_5038,N_3710,N_3614);
nand U5039 (N_5039,N_4004,N_1647);
or U5040 (N_5040,N_4277,N_4026);
nand U5041 (N_5041,N_4434,N_2145);
and U5042 (N_5042,N_935,N_2791);
nand U5043 (N_5043,N_4477,N_4584);
nor U5044 (N_5044,N_2170,N_1072);
or U5045 (N_5045,N_4819,N_1508);
nand U5046 (N_5046,N_3309,N_887);
xnor U5047 (N_5047,N_3534,N_3717);
or U5048 (N_5048,N_4496,N_421);
or U5049 (N_5049,N_3882,N_2589);
and U5050 (N_5050,N_184,N_2585);
or U5051 (N_5051,N_3046,N_124);
xor U5052 (N_5052,N_79,N_3274);
nand U5053 (N_5053,N_2016,N_2548);
and U5054 (N_5054,N_1658,N_1874);
nand U5055 (N_5055,N_948,N_3934);
xor U5056 (N_5056,N_1364,N_1479);
and U5057 (N_5057,N_3590,N_3817);
and U5058 (N_5058,N_911,N_4290);
or U5059 (N_5059,N_972,N_2292);
xor U5060 (N_5060,N_1740,N_143);
nor U5061 (N_5061,N_2070,N_2180);
or U5062 (N_5062,N_4617,N_3511);
nor U5063 (N_5063,N_284,N_1210);
and U5064 (N_5064,N_297,N_3350);
nand U5065 (N_5065,N_594,N_345);
or U5066 (N_5066,N_3591,N_2830);
xor U5067 (N_5067,N_3490,N_266);
nand U5068 (N_5068,N_3258,N_4608);
xor U5069 (N_5069,N_4317,N_608);
xnor U5070 (N_5070,N_1075,N_213);
xnor U5071 (N_5071,N_4389,N_2736);
and U5072 (N_5072,N_3502,N_489);
nand U5073 (N_5073,N_2283,N_4738);
nand U5074 (N_5074,N_3958,N_62);
xnor U5075 (N_5075,N_3159,N_2442);
xor U5076 (N_5076,N_3561,N_3415);
nand U5077 (N_5077,N_1683,N_3881);
nor U5078 (N_5078,N_4375,N_2428);
or U5079 (N_5079,N_1295,N_1201);
xnor U5080 (N_5080,N_688,N_1219);
nor U5081 (N_5081,N_3085,N_2060);
and U5082 (N_5082,N_3571,N_2924);
nand U5083 (N_5083,N_2196,N_3050);
and U5084 (N_5084,N_3250,N_3163);
xor U5085 (N_5085,N_2557,N_693);
or U5086 (N_5086,N_255,N_1898);
xor U5087 (N_5087,N_2708,N_739);
nor U5088 (N_5088,N_4356,N_4286);
xor U5089 (N_5089,N_1496,N_4367);
nand U5090 (N_5090,N_957,N_2371);
nor U5091 (N_5091,N_3482,N_1518);
nor U5092 (N_5092,N_188,N_1048);
nand U5093 (N_5093,N_3873,N_3726);
xor U5094 (N_5094,N_3595,N_836);
nor U5095 (N_5095,N_3669,N_84);
xnor U5096 (N_5096,N_1361,N_1165);
and U5097 (N_5097,N_3655,N_3418);
and U5098 (N_5098,N_630,N_4084);
xnor U5099 (N_5099,N_586,N_331);
xor U5100 (N_5100,N_102,N_2591);
or U5101 (N_5101,N_2176,N_455);
nor U5102 (N_5102,N_1288,N_2496);
and U5103 (N_5103,N_488,N_3063);
nor U5104 (N_5104,N_4152,N_3307);
xnor U5105 (N_5105,N_1356,N_1523);
nand U5106 (N_5106,N_709,N_2339);
or U5107 (N_5107,N_4717,N_2414);
and U5108 (N_5108,N_1817,N_3601);
xor U5109 (N_5109,N_1816,N_3104);
and U5110 (N_5110,N_875,N_4809);
or U5111 (N_5111,N_1875,N_1908);
nand U5112 (N_5112,N_3787,N_1249);
nor U5113 (N_5113,N_2113,N_3851);
or U5114 (N_5114,N_4897,N_2432);
xnor U5115 (N_5115,N_1582,N_2689);
or U5116 (N_5116,N_1552,N_3346);
xnor U5117 (N_5117,N_908,N_3051);
nand U5118 (N_5118,N_4736,N_163);
xnor U5119 (N_5119,N_3690,N_4961);
or U5120 (N_5120,N_4220,N_1812);
nor U5121 (N_5121,N_3245,N_4275);
and U5122 (N_5122,N_2782,N_1478);
or U5123 (N_5123,N_3485,N_2798);
and U5124 (N_5124,N_217,N_1471);
nor U5125 (N_5125,N_1197,N_1712);
and U5126 (N_5126,N_896,N_3359);
and U5127 (N_5127,N_4250,N_2687);
nand U5128 (N_5128,N_71,N_999);
and U5129 (N_5129,N_2223,N_95);
xor U5130 (N_5130,N_4690,N_4746);
nor U5131 (N_5131,N_985,N_498);
and U5132 (N_5132,N_1969,N_4933);
and U5133 (N_5133,N_1230,N_1416);
xor U5134 (N_5134,N_2148,N_2597);
nor U5135 (N_5135,N_3640,N_424);
xnor U5136 (N_5136,N_3798,N_136);
xnor U5137 (N_5137,N_773,N_4301);
xor U5138 (N_5138,N_2893,N_2177);
nand U5139 (N_5139,N_1727,N_4457);
and U5140 (N_5140,N_1586,N_1791);
or U5141 (N_5141,N_492,N_933);
nor U5142 (N_5142,N_3917,N_1531);
or U5143 (N_5143,N_4240,N_3608);
xor U5144 (N_5144,N_4844,N_4550);
nor U5145 (N_5145,N_937,N_3984);
nand U5146 (N_5146,N_4305,N_2005);
nand U5147 (N_5147,N_2726,N_2074);
nand U5148 (N_5148,N_4806,N_2296);
or U5149 (N_5149,N_3354,N_1266);
and U5150 (N_5150,N_2878,N_2273);
xnor U5151 (N_5151,N_2734,N_3935);
nand U5152 (N_5152,N_2233,N_1179);
nor U5153 (N_5153,N_4689,N_3732);
and U5154 (N_5154,N_3734,N_1619);
xnor U5155 (N_5155,N_2741,N_2899);
or U5156 (N_5156,N_3321,N_2568);
and U5157 (N_5157,N_1878,N_3878);
nor U5158 (N_5158,N_1003,N_2385);
xor U5159 (N_5159,N_4521,N_3904);
or U5160 (N_5160,N_1806,N_4221);
nor U5161 (N_5161,N_116,N_992);
nor U5162 (N_5162,N_4721,N_2376);
and U5163 (N_5163,N_500,N_954);
nand U5164 (N_5164,N_1370,N_942);
and U5165 (N_5165,N_3686,N_4635);
nand U5166 (N_5166,N_173,N_1465);
and U5167 (N_5167,N_3234,N_3045);
and U5168 (N_5168,N_2555,N_1198);
nor U5169 (N_5169,N_473,N_4231);
xnor U5170 (N_5170,N_383,N_3315);
xor U5171 (N_5171,N_4527,N_3061);
or U5172 (N_5172,N_1128,N_1746);
nor U5173 (N_5173,N_2367,N_1019);
nor U5174 (N_5174,N_4684,N_1227);
xor U5175 (N_5175,N_1259,N_2529);
nor U5176 (N_5176,N_2290,N_2593);
or U5177 (N_5177,N_4394,N_3989);
nor U5178 (N_5178,N_4781,N_1701);
nand U5179 (N_5179,N_748,N_3200);
and U5180 (N_5180,N_4419,N_2799);
or U5181 (N_5181,N_4884,N_2576);
nor U5182 (N_5182,N_4842,N_3041);
nand U5183 (N_5183,N_1520,N_1233);
nor U5184 (N_5184,N_348,N_4683);
and U5185 (N_5185,N_3764,N_565);
xnor U5186 (N_5186,N_794,N_3083);
nor U5187 (N_5187,N_215,N_1);
xor U5188 (N_5188,N_3407,N_4891);
nand U5189 (N_5189,N_4510,N_598);
nand U5190 (N_5190,N_3982,N_1311);
nor U5191 (N_5191,N_1105,N_3235);
nor U5192 (N_5192,N_304,N_3507);
or U5193 (N_5193,N_1481,N_566);
or U5194 (N_5194,N_2249,N_4184);
nand U5195 (N_5195,N_3205,N_2173);
xor U5196 (N_5196,N_4208,N_4960);
nand U5197 (N_5197,N_320,N_2166);
or U5198 (N_5198,N_357,N_379);
nor U5199 (N_5199,N_1322,N_2842);
xor U5200 (N_5200,N_1603,N_4898);
and U5201 (N_5201,N_3358,N_2390);
xnor U5202 (N_5202,N_4150,N_1568);
nand U5203 (N_5203,N_1509,N_4255);
nand U5204 (N_5204,N_3644,N_3816);
or U5205 (N_5205,N_4765,N_4156);
or U5206 (N_5206,N_81,N_4894);
or U5207 (N_5207,N_705,N_4976);
xor U5208 (N_5208,N_4970,N_1422);
nand U5209 (N_5209,N_367,N_1173);
or U5210 (N_5210,N_2991,N_2881);
and U5211 (N_5211,N_2029,N_1467);
and U5212 (N_5212,N_7,N_2527);
nor U5213 (N_5213,N_4292,N_812);
nor U5214 (N_5214,N_2772,N_1133);
xor U5215 (N_5215,N_1669,N_861);
xor U5216 (N_5216,N_3789,N_3813);
or U5217 (N_5217,N_1590,N_2654);
or U5218 (N_5218,N_1793,N_2473);
and U5219 (N_5219,N_3483,N_728);
and U5220 (N_5220,N_4118,N_1783);
xor U5221 (N_5221,N_1138,N_469);
or U5222 (N_5222,N_1591,N_4117);
or U5223 (N_5223,N_4869,N_1790);
nand U5224 (N_5224,N_2641,N_2002);
nor U5225 (N_5225,N_1171,N_2182);
and U5226 (N_5226,N_4251,N_4872);
and U5227 (N_5227,N_1102,N_1070);
xnor U5228 (N_5228,N_703,N_3795);
nand U5229 (N_5229,N_3284,N_1994);
and U5230 (N_5230,N_1545,N_1177);
nand U5231 (N_5231,N_4731,N_4786);
and U5232 (N_5232,N_1713,N_128);
nor U5233 (N_5233,N_3199,N_397);
or U5234 (N_5234,N_2844,N_2342);
nand U5235 (N_5235,N_4259,N_3096);
nand U5236 (N_5236,N_2590,N_1444);
xor U5237 (N_5237,N_4176,N_3010);
or U5238 (N_5238,N_3172,N_113);
and U5239 (N_5239,N_3265,N_3969);
nor U5240 (N_5240,N_1267,N_2216);
nand U5241 (N_5241,N_3857,N_4161);
or U5242 (N_5242,N_3499,N_4113);
or U5243 (N_5243,N_2603,N_422);
nand U5244 (N_5244,N_551,N_2089);
xor U5245 (N_5245,N_399,N_257);
nor U5246 (N_5246,N_3876,N_4196);
xnor U5247 (N_5247,N_4927,N_2618);
nor U5248 (N_5248,N_3428,N_4469);
or U5249 (N_5249,N_2602,N_1599);
and U5250 (N_5250,N_3874,N_3246);
xnor U5251 (N_5251,N_4461,N_3466);
xor U5252 (N_5252,N_1947,N_4955);
xnor U5253 (N_5253,N_1091,N_2946);
and U5254 (N_5254,N_4463,N_3832);
nor U5255 (N_5255,N_2136,N_4405);
nor U5256 (N_5256,N_2503,N_3004);
nand U5257 (N_5257,N_335,N_1909);
xnor U5258 (N_5258,N_4514,N_4718);
xnor U5259 (N_5259,N_1551,N_181);
xor U5260 (N_5260,N_1796,N_4748);
nor U5261 (N_5261,N_4458,N_4349);
and U5262 (N_5262,N_2259,N_240);
or U5263 (N_5263,N_2270,N_2756);
or U5264 (N_5264,N_323,N_1985);
nor U5265 (N_5265,N_2688,N_2938);
or U5266 (N_5266,N_4895,N_6);
xor U5267 (N_5267,N_717,N_3572);
and U5268 (N_5268,N_2149,N_2594);
nor U5269 (N_5269,N_1871,N_2957);
xor U5270 (N_5270,N_4102,N_4293);
and U5271 (N_5271,N_1248,N_716);
nor U5272 (N_5272,N_2477,N_1116);
nor U5273 (N_5273,N_509,N_1462);
nor U5274 (N_5274,N_4359,N_3241);
or U5275 (N_5275,N_3128,N_197);
and U5276 (N_5276,N_811,N_396);
nor U5277 (N_5277,N_2099,N_1274);
nor U5278 (N_5278,N_3773,N_2402);
or U5279 (N_5279,N_1455,N_3098);
nand U5280 (N_5280,N_2240,N_1225);
and U5281 (N_5281,N_225,N_1394);
nor U5282 (N_5282,N_2506,N_464);
xor U5283 (N_5283,N_356,N_1384);
and U5284 (N_5284,N_1348,N_1906);
or U5285 (N_5285,N_4217,N_3395);
nor U5286 (N_5286,N_3526,N_3416);
nor U5287 (N_5287,N_1572,N_4515);
nand U5288 (N_5288,N_3509,N_1176);
and U5289 (N_5289,N_865,N_3130);
or U5290 (N_5290,N_713,N_692);
and U5291 (N_5291,N_2710,N_2989);
xor U5292 (N_5292,N_2124,N_1369);
nor U5293 (N_5293,N_825,N_4606);
and U5294 (N_5294,N_2316,N_2459);
xnor U5295 (N_5295,N_1205,N_3025);
nor U5296 (N_5296,N_1628,N_4144);
nand U5297 (N_5297,N_3498,N_1272);
nor U5298 (N_5298,N_2142,N_1721);
nand U5299 (N_5299,N_1134,N_2627);
or U5300 (N_5300,N_3627,N_3562);
nand U5301 (N_5301,N_1846,N_3656);
or U5302 (N_5302,N_1841,N_3445);
xor U5303 (N_5303,N_2920,N_3654);
nand U5304 (N_5304,N_2372,N_351);
and U5305 (N_5305,N_4471,N_1211);
or U5306 (N_5306,N_823,N_4040);
nand U5307 (N_5307,N_2701,N_1950);
and U5308 (N_5308,N_4261,N_3008);
xnor U5309 (N_5309,N_1103,N_2247);
nor U5310 (N_5310,N_4658,N_990);
or U5311 (N_5311,N_233,N_1938);
xor U5312 (N_5312,N_2199,N_1007);
or U5313 (N_5313,N_4913,N_3283);
nand U5314 (N_5314,N_4484,N_661);
nor U5315 (N_5315,N_1454,N_4790);
or U5316 (N_5316,N_2391,N_1778);
nor U5317 (N_5317,N_583,N_842);
xor U5318 (N_5318,N_3493,N_1026);
nor U5319 (N_5319,N_3101,N_1094);
or U5320 (N_5320,N_2595,N_1792);
xor U5321 (N_5321,N_1411,N_2866);
nand U5322 (N_5322,N_2320,N_3370);
nor U5323 (N_5323,N_1285,N_1063);
or U5324 (N_5324,N_4041,N_4291);
and U5325 (N_5325,N_1192,N_4086);
or U5326 (N_5326,N_1193,N_3268);
nand U5327 (N_5327,N_2852,N_360);
xnor U5328 (N_5328,N_3181,N_2998);
and U5329 (N_5329,N_4412,N_2486);
nor U5330 (N_5330,N_1321,N_1769);
and U5331 (N_5331,N_1434,N_1818);
or U5332 (N_5332,N_73,N_3639);
nand U5333 (N_5333,N_3386,N_2039);
nand U5334 (N_5334,N_4735,N_4932);
or U5335 (N_5335,N_4307,N_4051);
and U5336 (N_5336,N_4954,N_3550);
nor U5337 (N_5337,N_2347,N_86);
nand U5338 (N_5338,N_989,N_190);
nand U5339 (N_5339,N_146,N_3016);
or U5340 (N_5340,N_2648,N_3923);
nor U5341 (N_5341,N_806,N_3913);
nor U5342 (N_5342,N_1897,N_301);
xor U5343 (N_5343,N_629,N_3675);
or U5344 (N_5344,N_3427,N_2355);
or U5345 (N_5345,N_2757,N_3811);
xnor U5346 (N_5346,N_3220,N_4916);
or U5347 (N_5347,N_3461,N_3463);
nand U5348 (N_5348,N_1954,N_75);
xnor U5349 (N_5349,N_1352,N_3115);
nor U5350 (N_5350,N_1542,N_2340);
xnor U5351 (N_5351,N_4337,N_4402);
nand U5352 (N_5352,N_1538,N_3082);
and U5353 (N_5353,N_1579,N_510);
or U5354 (N_5354,N_4130,N_4476);
xnor U5355 (N_5355,N_1087,N_1125);
or U5356 (N_5356,N_912,N_2601);
or U5357 (N_5357,N_3327,N_1338);
and U5358 (N_5358,N_2307,N_4447);
nor U5359 (N_5359,N_2636,N_4168);
nand U5360 (N_5360,N_1180,N_1707);
nand U5361 (N_5361,N_4232,N_2152);
nand U5362 (N_5362,N_1890,N_1671);
or U5363 (N_5363,N_2883,N_4234);
or U5364 (N_5364,N_4627,N_802);
and U5365 (N_5365,N_1190,N_3039);
or U5366 (N_5366,N_2208,N_1519);
xor U5367 (N_5367,N_4726,N_1608);
xor U5368 (N_5368,N_4889,N_3535);
or U5369 (N_5369,N_111,N_3472);
or U5370 (N_5370,N_3753,N_4468);
or U5371 (N_5371,N_1589,N_377);
or U5372 (N_5372,N_2287,N_3492);
nand U5373 (N_5373,N_1926,N_1992);
xor U5374 (N_5374,N_3606,N_2035);
nand U5375 (N_5375,N_2912,N_4909);
or U5376 (N_5376,N_2611,N_359);
and U5377 (N_5377,N_3353,N_405);
nor U5378 (N_5378,N_2553,N_1879);
and U5379 (N_5379,N_4920,N_324);
nand U5380 (N_5380,N_3630,N_557);
and U5381 (N_5381,N_3340,N_261);
or U5382 (N_5382,N_2324,N_1595);
nand U5383 (N_5383,N_110,N_889);
nand U5384 (N_5384,N_2843,N_4128);
nand U5385 (N_5385,N_4465,N_1062);
and U5386 (N_5386,N_560,N_2450);
and U5387 (N_5387,N_2183,N_57);
or U5388 (N_5388,N_2927,N_441);
and U5389 (N_5389,N_3619,N_736);
nand U5390 (N_5390,N_4829,N_2365);
or U5391 (N_5391,N_2478,N_2081);
and U5392 (N_5392,N_650,N_3993);
and U5393 (N_5393,N_4252,N_700);
xor U5394 (N_5394,N_1876,N_3763);
or U5395 (N_5395,N_4973,N_3759);
nor U5396 (N_5396,N_2079,N_1080);
xor U5397 (N_5397,N_2026,N_3688);
xor U5398 (N_5398,N_4393,N_4655);
nor U5399 (N_5399,N_30,N_3064);
nor U5400 (N_5400,N_131,N_3990);
nand U5401 (N_5401,N_579,N_839);
xnor U5402 (N_5402,N_2076,N_2889);
nor U5403 (N_5403,N_3515,N_201);
and U5404 (N_5404,N_750,N_2024);
xor U5405 (N_5405,N_1964,N_639);
xnor U5406 (N_5406,N_4028,N_333);
xor U5407 (N_5407,N_4800,N_3943);
xnor U5408 (N_5408,N_2807,N_446);
nor U5409 (N_5409,N_3260,N_3184);
nor U5410 (N_5410,N_4485,N_2633);
and U5411 (N_5411,N_2147,N_2257);
xor U5412 (N_5412,N_1825,N_563);
and U5413 (N_5413,N_4436,N_4867);
nor U5414 (N_5414,N_2386,N_1040);
nand U5415 (N_5415,N_2091,N_1312);
and U5416 (N_5416,N_3449,N_1157);
and U5417 (N_5417,N_922,N_1680);
and U5418 (N_5418,N_3603,N_1044);
or U5419 (N_5419,N_721,N_3188);
and U5420 (N_5420,N_602,N_2979);
xnor U5421 (N_5421,N_2723,N_4697);
xor U5422 (N_5422,N_2859,N_4000);
or U5423 (N_5423,N_2515,N_1118);
and U5424 (N_5424,N_701,N_4620);
nand U5425 (N_5425,N_3319,N_699);
xnor U5426 (N_5426,N_4524,N_370);
xnor U5427 (N_5427,N_3451,N_2523);
xnor U5428 (N_5428,N_928,N_2670);
nand U5429 (N_5429,N_2241,N_1486);
or U5430 (N_5430,N_2921,N_2119);
nor U5431 (N_5431,N_3942,N_1298);
and U5432 (N_5432,N_3902,N_1941);
nand U5433 (N_5433,N_1715,N_2655);
nand U5434 (N_5434,N_2381,N_3859);
xor U5435 (N_5435,N_4139,N_274);
and U5436 (N_5436,N_1135,N_3842);
nand U5437 (N_5437,N_4302,N_743);
xor U5438 (N_5438,N_2416,N_3322);
xor U5439 (N_5439,N_3460,N_65);
xor U5440 (N_5440,N_3145,N_365);
nor U5441 (N_5441,N_3865,N_2086);
or U5442 (N_5442,N_4985,N_3826);
xnor U5443 (N_5443,N_1611,N_130);
or U5444 (N_5444,N_4294,N_4940);
nand U5445 (N_5445,N_3171,N_4075);
or U5446 (N_5446,N_1625,N_3531);
nor U5447 (N_5447,N_3801,N_4581);
xor U5448 (N_5448,N_2139,N_2276);
or U5449 (N_5449,N_892,N_1940);
nor U5450 (N_5450,N_799,N_4667);
xnor U5451 (N_5451,N_2470,N_1146);
nor U5452 (N_5452,N_2218,N_4147);
nand U5453 (N_5453,N_1469,N_3363);
and U5454 (N_5454,N_763,N_529);
or U5455 (N_5455,N_3406,N_4647);
nor U5456 (N_5456,N_547,N_499);
or U5457 (N_5457,N_90,N_3077);
nor U5458 (N_5458,N_2134,N_4383);
xor U5459 (N_5459,N_38,N_4571);
or U5460 (N_5460,N_2776,N_941);
or U5461 (N_5461,N_1440,N_3387);
nand U5462 (N_5462,N_2192,N_884);
nand U5463 (N_5463,N_4661,N_4135);
or U5464 (N_5464,N_3477,N_653);
nor U5465 (N_5465,N_4400,N_3578);
or U5466 (N_5466,N_156,N_2574);
or U5467 (N_5467,N_4615,N_4444);
nor U5468 (N_5468,N_4556,N_4490);
or U5469 (N_5469,N_2392,N_1152);
nand U5470 (N_5470,N_829,N_2337);
or U5471 (N_5471,N_1645,N_1853);
nor U5472 (N_5472,N_2704,N_3182);
nor U5473 (N_5473,N_3527,N_793);
and U5474 (N_5474,N_1166,N_1539);
nand U5475 (N_5475,N_3324,N_3446);
nor U5476 (N_5476,N_1869,N_1862);
or U5477 (N_5477,N_2411,N_34);
and U5478 (N_5478,N_2452,N_49);
nand U5479 (N_5479,N_2505,N_54);
xor U5480 (N_5480,N_3837,N_689);
xnor U5481 (N_5481,N_1488,N_2649);
and U5482 (N_5482,N_897,N_4066);
or U5483 (N_5483,N_1163,N_392);
and U5484 (N_5484,N_1514,N_2742);
or U5485 (N_5485,N_1310,N_1826);
nor U5486 (N_5486,N_502,N_4095);
and U5487 (N_5487,N_4306,N_475);
and U5488 (N_5488,N_2657,N_445);
and U5489 (N_5489,N_3365,N_408);
nand U5490 (N_5490,N_522,N_1987);
or U5491 (N_5491,N_4088,N_1718);
nand U5492 (N_5492,N_3808,N_1324);
nand U5493 (N_5493,N_2388,N_3218);
and U5494 (N_5494,N_3844,N_135);
xor U5495 (N_5495,N_4557,N_3412);
or U5496 (N_5496,N_278,N_4052);
or U5497 (N_5497,N_2753,N_3287);
nand U5498 (N_5498,N_4760,N_1574);
nor U5499 (N_5499,N_2858,N_4410);
xnor U5500 (N_5500,N_826,N_47);
and U5501 (N_5501,N_4474,N_24);
and U5502 (N_5502,N_4904,N_3584);
and U5503 (N_5503,N_3592,N_3149);
nor U5504 (N_5504,N_4249,N_879);
and U5505 (N_5505,N_2538,N_2087);
nor U5506 (N_5506,N_4877,N_589);
nor U5507 (N_5507,N_1438,N_1217);
or U5508 (N_5508,N_4958,N_2986);
nand U5509 (N_5509,N_4243,N_3741);
nand U5510 (N_5510,N_133,N_1123);
nand U5511 (N_5511,N_4988,N_4060);
xnor U5512 (N_5512,N_4422,N_3756);
or U5513 (N_5513,N_4965,N_1122);
nand U5514 (N_5514,N_2278,N_527);
nor U5515 (N_5515,N_4081,N_3379);
xnor U5516 (N_5516,N_4201,N_4539);
and U5517 (N_5517,N_4132,N_4820);
or U5518 (N_5518,N_479,N_3564);
nor U5519 (N_5519,N_1013,N_460);
or U5520 (N_5520,N_4046,N_1887);
nand U5521 (N_5521,N_1977,N_1614);
or U5522 (N_5522,N_2100,N_4686);
nor U5523 (N_5523,N_2158,N_533);
nand U5524 (N_5524,N_841,N_4423);
or U5525 (N_5525,N_1613,N_4749);
nand U5526 (N_5526,N_2446,N_1917);
nor U5527 (N_5527,N_4421,N_1607);
and U5528 (N_5528,N_4705,N_1101);
xor U5529 (N_5529,N_786,N_3022);
nand U5530 (N_5530,N_4219,N_2980);
or U5531 (N_5531,N_1942,N_973);
or U5532 (N_5532,N_1881,N_4357);
or U5533 (N_5533,N_12,N_1970);
nor U5534 (N_5534,N_3960,N_4483);
nand U5535 (N_5535,N_4511,N_1723);
nand U5536 (N_5536,N_1474,N_4347);
or U5537 (N_5537,N_3750,N_3021);
nand U5538 (N_5538,N_1612,N_1051);
and U5539 (N_5539,N_1692,N_898);
and U5540 (N_5540,N_2997,N_3855);
nand U5541 (N_5541,N_1333,N_4574);
or U5542 (N_5542,N_4372,N_4883);
nand U5543 (N_5543,N_3232,N_4078);
nor U5544 (N_5544,N_2484,N_1390);
or U5545 (N_5545,N_4720,N_3945);
and U5546 (N_5546,N_3853,N_1358);
xnor U5547 (N_5547,N_984,N_3786);
xor U5548 (N_5548,N_1905,N_4454);
nor U5549 (N_5549,N_3693,N_3683);
and U5550 (N_5550,N_450,N_1360);
xor U5551 (N_5551,N_516,N_4941);
xor U5552 (N_5552,N_4257,N_3056);
xor U5553 (N_5553,N_4971,N_645);
nor U5554 (N_5554,N_1414,N_3312);
nor U5555 (N_5555,N_1403,N_2885);
or U5556 (N_5556,N_4769,N_109);
or U5557 (N_5557,N_4665,N_2015);
xnor U5558 (N_5558,N_4535,N_2094);
nor U5559 (N_5559,N_1181,N_1336);
xnor U5560 (N_5560,N_2966,N_4876);
and U5561 (N_5561,N_3156,N_273);
and U5562 (N_5562,N_710,N_3761);
nor U5563 (N_5563,N_2915,N_3473);
nand U5564 (N_5564,N_1667,N_1453);
or U5565 (N_5565,N_3320,N_67);
nand U5566 (N_5566,N_1216,N_3144);
and U5567 (N_5567,N_3032,N_1609);
and U5568 (N_5568,N_162,N_3946);
nand U5569 (N_5569,N_3388,N_77);
xnor U5570 (N_5570,N_611,N_3369);
nand U5571 (N_5571,N_2126,N_2111);
nand U5572 (N_5572,N_3800,N_1155);
or U5573 (N_5573,N_4241,N_501);
or U5574 (N_5574,N_883,N_1668);
xnor U5575 (N_5575,N_816,N_4377);
nor U5576 (N_5576,N_2874,N_1714);
and U5577 (N_5577,N_4734,N_2488);
nor U5578 (N_5578,N_2934,N_2917);
xnor U5579 (N_5579,N_4803,N_3272);
xnor U5580 (N_5580,N_4924,N_3456);
xnor U5581 (N_5581,N_657,N_4917);
and U5582 (N_5582,N_4676,N_1189);
xor U5583 (N_5583,N_3624,N_1314);
nand U5584 (N_5584,N_809,N_3439);
nand U5585 (N_5585,N_1154,N_2519);
nand U5586 (N_5586,N_3587,N_910);
nor U5587 (N_5587,N_1553,N_3317);
nand U5588 (N_5588,N_1910,N_3212);
xor U5589 (N_5589,N_3632,N_4227);
and U5590 (N_5590,N_4169,N_3294);
nand U5591 (N_5591,N_1742,N_337);
xor U5592 (N_5592,N_1708,N_37);
or U5593 (N_5593,N_4214,N_4287);
or U5594 (N_5594,N_1099,N_2253);
xnor U5595 (N_5595,N_2763,N_3658);
or U5596 (N_5596,N_714,N_4801);
or U5597 (N_5597,N_494,N_154);
or U5598 (N_5598,N_4537,N_2164);
nor U5599 (N_5599,N_1732,N_1045);
or U5600 (N_5600,N_2847,N_4695);
and U5601 (N_5601,N_2898,N_3106);
xor U5602 (N_5602,N_1482,N_646);
nor U5603 (N_5603,N_4816,N_2672);
nor U5604 (N_5604,N_1760,N_4758);
and U5605 (N_5605,N_2905,N_1242);
and U5606 (N_5606,N_503,N_1451);
and U5607 (N_5607,N_4699,N_375);
xor U5608 (N_5608,N_76,N_2031);
nand U5609 (N_5609,N_1581,N_4875);
or U5610 (N_5610,N_4613,N_3516);
nor U5611 (N_5611,N_139,N_4205);
and U5612 (N_5612,N_2724,N_3402);
and U5613 (N_5613,N_3471,N_876);
nand U5614 (N_5614,N_2059,N_457);
or U5615 (N_5615,N_4215,N_3866);
nand U5616 (N_5616,N_4131,N_4902);
nor U5617 (N_5617,N_1844,N_3109);
and U5618 (N_5618,N_3594,N_4133);
nor U5619 (N_5619,N_89,N_1150);
xor U5620 (N_5620,N_1126,N_2498);
xnor U5621 (N_5621,N_1744,N_4767);
nand U5622 (N_5622,N_289,N_1930);
nor U5623 (N_5623,N_3995,N_2839);
nor U5624 (N_5624,N_1280,N_4213);
nor U5625 (N_5625,N_1693,N_918);
xor U5626 (N_5626,N_3997,N_668);
or U5627 (N_5627,N_4885,N_4203);
and U5628 (N_5628,N_1684,N_1430);
nor U5629 (N_5629,N_2159,N_1731);
nor U5630 (N_5630,N_2098,N_92);
xnor U5631 (N_5631,N_2717,N_4439);
nor U5632 (N_5632,N_2150,N_1412);
xor U5633 (N_5633,N_4773,N_2615);
or U5634 (N_5634,N_874,N_1335);
nand U5635 (N_5635,N_765,N_4263);
xor U5636 (N_5636,N_4754,N_575);
or U5637 (N_5637,N_1617,N_934);
nor U5638 (N_5638,N_1386,N_4659);
nor U5639 (N_5639,N_776,N_4044);
or U5640 (N_5640,N_2959,N_2495);
and U5641 (N_5641,N_4420,N_1832);
nor U5642 (N_5642,N_183,N_1724);
nand U5643 (N_5643,N_4810,N_4310);
and U5644 (N_5644,N_1789,N_3178);
xnor U5645 (N_5645,N_891,N_3555);
xor U5646 (N_5646,N_4225,N_2255);
xor U5647 (N_5647,N_4675,N_684);
or U5648 (N_5648,N_873,N_4944);
or U5649 (N_5649,N_4549,N_4006);
xnor U5650 (N_5650,N_747,N_4516);
nor U5651 (N_5651,N_2128,N_276);
xor U5652 (N_5652,N_2434,N_2215);
nor U5653 (N_5653,N_2410,N_2429);
or U5654 (N_5654,N_4473,N_3271);
and U5655 (N_5655,N_1220,N_3299);
xor U5656 (N_5656,N_3748,N_161);
nor U5657 (N_5657,N_3058,N_3110);
nand U5658 (N_5658,N_2764,N_4418);
nand U5659 (N_5659,N_3478,N_1160);
and U5660 (N_5660,N_4791,N_2682);
or U5661 (N_5661,N_4183,N_2237);
nor U5662 (N_5662,N_1802,N_2607);
xor U5663 (N_5663,N_2812,N_2405);
xnor U5664 (N_5664,N_3280,N_2988);
xor U5665 (N_5665,N_4233,N_4398);
xor U5666 (N_5666,N_2280,N_1294);
or U5667 (N_5667,N_4823,N_1372);
and U5668 (N_5668,N_461,N_1287);
and U5669 (N_5669,N_3,N_2962);
and U5670 (N_5670,N_4019,N_900);
xor U5671 (N_5671,N_2825,N_4761);
nand U5672 (N_5672,N_1660,N_2463);
or U5673 (N_5673,N_558,N_2187);
nor U5674 (N_5674,N_779,N_3355);
xnor U5675 (N_5675,N_3625,N_2341);
xnor U5676 (N_5676,N_4506,N_3505);
nor U5677 (N_5677,N_535,N_4448);
and U5678 (N_5678,N_2279,N_2851);
nor U5679 (N_5679,N_2972,N_3454);
nor U5680 (N_5680,N_4332,N_1631);
or U5681 (N_5681,N_3920,N_3403);
nor U5682 (N_5682,N_1745,N_1247);
and U5683 (N_5683,N_3108,N_4497);
or U5684 (N_5684,N_3847,N_1799);
and U5685 (N_5685,N_2120,N_2513);
or U5686 (N_5686,N_4406,N_296);
and U5687 (N_5687,N_2476,N_3027);
and U5688 (N_5688,N_4452,N_328);
nand U5689 (N_5689,N_554,N_1273);
xor U5690 (N_5690,N_916,N_1289);
nor U5691 (N_5691,N_4915,N_1034);
xor U5692 (N_5692,N_1847,N_3476);
nand U5693 (N_5693,N_3557,N_114);
or U5694 (N_5694,N_4224,N_209);
and U5695 (N_5695,N_4326,N_690);
xnor U5696 (N_5696,N_2630,N_1477);
nor U5697 (N_5697,N_3206,N_3972);
nand U5698 (N_5698,N_2650,N_3701);
or U5699 (N_5699,N_27,N_1162);
xor U5700 (N_5700,N_3393,N_3558);
xor U5701 (N_5701,N_2642,N_2384);
nand U5702 (N_5702,N_1191,N_581);
xnor U5703 (N_5703,N_920,N_797);
or U5704 (N_5704,N_180,N_2577);
and U5705 (N_5705,N_1346,N_2828);
xnor U5706 (N_5706,N_2976,N_3903);
and U5707 (N_5707,N_4413,N_1821);
or U5708 (N_5708,N_3352,N_800);
xor U5709 (N_5709,N_744,N_867);
or U5710 (N_5710,N_1131,N_1524);
nor U5711 (N_5711,N_1387,N_3974);
nor U5712 (N_5712,N_4464,N_3450);
nand U5713 (N_5713,N_1140,N_2674);
xnor U5714 (N_5714,N_930,N_299);
nand U5715 (N_5715,N_435,N_4653);
and U5716 (N_5716,N_1124,N_21);
nand U5717 (N_5717,N_781,N_427);
nor U5718 (N_5718,N_2256,N_3400);
and U5719 (N_5719,N_963,N_2969);
xnor U5720 (N_5720,N_4937,N_3987);
or U5721 (N_5721,N_628,N_4472);
nor U5722 (N_5722,N_3819,N_3377);
nor U5723 (N_5723,N_4351,N_582);
or U5724 (N_5724,N_572,N_4501);
xnor U5725 (N_5725,N_2534,N_4874);
and U5726 (N_5726,N_2658,N_4901);
xor U5727 (N_5727,N_2317,N_3443);
or U5728 (N_5728,N_3908,N_158);
and U5729 (N_5729,N_1529,N_672);
or U5730 (N_5730,N_4120,N_231);
xnor U5731 (N_5731,N_1738,N_3092);
or U5732 (N_5732,N_2112,N_4762);
nor U5733 (N_5733,N_526,N_1093);
nand U5734 (N_5734,N_2333,N_2037);
xor U5735 (N_5735,N_2542,N_417);
xor U5736 (N_5736,N_186,N_1653);
nor U5737 (N_5737,N_2779,N_1466);
or U5738 (N_5738,N_4614,N_2624);
and U5739 (N_5739,N_1848,N_3560);
or U5740 (N_5740,N_2071,N_411);
nand U5741 (N_5741,N_1064,N_3437);
nand U5742 (N_5742,N_1028,N_31);
and U5743 (N_5743,N_3155,N_3755);
and U5744 (N_5744,N_4657,N_4818);
or U5745 (N_5745,N_2213,N_2301);
nand U5746 (N_5746,N_1860,N_2133);
xnor U5747 (N_5747,N_2932,N_2600);
nand U5748 (N_5748,N_1255,N_3699);
and U5749 (N_5749,N_2507,N_3348);
nor U5750 (N_5750,N_1264,N_632);
nor U5751 (N_5751,N_3950,N_3953);
xnor U5752 (N_5752,N_145,N_543);
and U5753 (N_5753,N_98,N_4371);
xnor U5754 (N_5754,N_2831,N_635);
and U5755 (N_5755,N_4442,N_2747);
and U5756 (N_5756,N_3841,N_4805);
nand U5757 (N_5757,N_4630,N_2036);
xnor U5758 (N_5758,N_573,N_3433);
nor U5759 (N_5759,N_4799,N_2775);
or U5760 (N_5760,N_3991,N_2795);
or U5761 (N_5761,N_631,N_4945);
or U5762 (N_5762,N_402,N_4929);
nor U5763 (N_5763,N_1436,N_1137);
or U5764 (N_5764,N_2359,N_2855);
nand U5765 (N_5765,N_766,N_666);
nor U5766 (N_5766,N_4148,N_462);
nor U5767 (N_5767,N_1279,N_4663);
nor U5768 (N_5768,N_474,N_2397);
nor U5769 (N_5769,N_85,N_1652);
xor U5770 (N_5770,N_1894,N_4185);
nor U5771 (N_5771,N_3519,N_2911);
nand U5772 (N_5772,N_4235,N_3442);
nand U5773 (N_5773,N_1407,N_3276);
xnor U5774 (N_5774,N_3898,N_4466);
xnor U5775 (N_5775,N_1304,N_2345);
nor U5776 (N_5776,N_3660,N_3086);
or U5777 (N_5777,N_1317,N_3221);
nand U5778 (N_5778,N_2325,N_3316);
nand U5779 (N_5779,N_1811,N_3687);
nor U5780 (N_5780,N_2204,N_4604);
nor U5781 (N_5781,N_4975,N_4662);
nand U5782 (N_5782,N_3131,N_4845);
or U5783 (N_5783,N_2908,N_792);
and U5784 (N_5784,N_4207,N_711);
nand U5785 (N_5785,N_2041,N_3076);
and U5786 (N_5786,N_185,N_436);
or U5787 (N_5787,N_3822,N_3279);
and U5788 (N_5788,N_3223,N_295);
nand U5789 (N_5789,N_2916,N_3698);
nor U5790 (N_5790,N_4171,N_1098);
xor U5791 (N_5791,N_850,N_3867);
nor U5792 (N_5792,N_2191,N_4780);
nor U5793 (N_5793,N_1493,N_2203);
xor U5794 (N_5794,N_127,N_2066);
or U5795 (N_5795,N_552,N_3243);
nor U5796 (N_5796,N_3209,N_931);
nor U5797 (N_5797,N_4893,N_539);
nor U5798 (N_5798,N_959,N_2138);
or U5799 (N_5799,N_2549,N_1426);
nand U5800 (N_5800,N_2592,N_4396);
nand U5801 (N_5801,N_1765,N_3467);
nand U5802 (N_5802,N_1918,N_412);
or U5803 (N_5803,N_1548,N_4737);
nor U5804 (N_5804,N_1859,N_4743);
and U5805 (N_5805,N_3702,N_983);
nand U5806 (N_5806,N_4906,N_395);
nor U5807 (N_5807,N_4374,N_1473);
or U5808 (N_5808,N_3662,N_2067);
or U5809 (N_5809,N_3005,N_2288);
xor U5810 (N_5810,N_1867,N_2935);
nand U5811 (N_5811,N_3520,N_2752);
nand U5812 (N_5812,N_995,N_4859);
nor U5813 (N_5813,N_3335,N_2500);
nand U5814 (N_5814,N_310,N_3742);
or U5815 (N_5815,N_3087,N_2396);
or U5816 (N_5816,N_2030,N_604);
xor U5817 (N_5817,N_4919,N_1834);
or U5818 (N_5818,N_4590,N_437);
xor U5819 (N_5819,N_3780,N_4063);
and U5820 (N_5820,N_3807,N_3382);
nand U5821 (N_5821,N_3914,N_3648);
and U5822 (N_5822,N_4994,N_4338);
nand U5823 (N_5823,N_1656,N_3001);
or U5824 (N_5824,N_3068,N_2914);
xnor U5825 (N_5825,N_4195,N_327);
xor U5826 (N_5826,N_3230,N_3673);
xor U5827 (N_5827,N_2771,N_1344);
and U5828 (N_5828,N_279,N_3593);
nor U5829 (N_5829,N_3431,N_3411);
nand U5830 (N_5830,N_2569,N_2127);
nor U5831 (N_5831,N_2684,N_760);
xnor U5832 (N_5832,N_3924,N_1206);
xor U5833 (N_5833,N_4187,N_3362);
nand U5834 (N_5834,N_4708,N_769);
or U5835 (N_5835,N_2338,N_3055);
and U5836 (N_5836,N_4959,N_425);
and U5837 (N_5837,N_478,N_410);
nor U5838 (N_5838,N_4416,N_2755);
xor U5839 (N_5839,N_3986,N_4950);
xnor U5840 (N_5840,N_4014,N_1963);
xor U5841 (N_5841,N_1503,N_2132);
xnor U5842 (N_5842,N_685,N_3818);
and U5843 (N_5843,N_979,N_2460);
and U5844 (N_5844,N_1831,N_2370);
xnor U5845 (N_5845,N_346,N_137);
and U5846 (N_5846,N_4724,N_734);
xnor U5847 (N_5847,N_1148,N_4863);
and U5848 (N_5848,N_1828,N_3425);
or U5849 (N_5849,N_2222,N_1275);
and U5850 (N_5850,N_1814,N_868);
nor U5851 (N_5851,N_1900,N_4888);
and U5852 (N_5852,N_3574,N_506);
or U5853 (N_5853,N_4595,N_2034);
nand U5854 (N_5854,N_3887,N_2913);
and U5855 (N_5855,N_4784,N_2543);
xor U5856 (N_5856,N_493,N_1497);
xnor U5857 (N_5857,N_1300,N_1929);
or U5858 (N_5858,N_3907,N_2873);
nor U5859 (N_5859,N_4429,N_665);
xnor U5860 (N_5860,N_1262,N_222);
nor U5861 (N_5861,N_4193,N_872);
xor U5862 (N_5862,N_1084,N_2535);
nor U5863 (N_5863,N_2993,N_2692);
and U5864 (N_5864,N_4968,N_3253);
xor U5865 (N_5865,N_3556,N_4727);
nor U5866 (N_5866,N_244,N_325);
nor U5867 (N_5867,N_2744,N_3704);
and U5868 (N_5868,N_1169,N_3292);
or U5869 (N_5869,N_3757,N_3988);
nand U5870 (N_5870,N_2879,N_2850);
nand U5871 (N_5871,N_1694,N_1733);
or U5872 (N_5872,N_3278,N_4752);
or U5873 (N_5873,N_3537,N_1351);
xor U5874 (N_5874,N_35,N_1536);
nand U5875 (N_5875,N_1883,N_4157);
nand U5876 (N_5876,N_2897,N_4980);
nor U5877 (N_5877,N_2464,N_2796);
or U5878 (N_5878,N_1670,N_2078);
nor U5879 (N_5879,N_2418,N_82);
and U5880 (N_5880,N_3289,N_3011);
xnor U5881 (N_5881,N_43,N_3420);
xor U5882 (N_5882,N_1686,N_1033);
nand U5883 (N_5883,N_3029,N_754);
nand U5884 (N_5884,N_2228,N_4324);
nor U5885 (N_5885,N_2072,N_2200);
or U5886 (N_5886,N_4771,N_4685);
or U5887 (N_5887,N_3724,N_622);
xnor U5888 (N_5888,N_2186,N_977);
and U5889 (N_5889,N_1710,N_256);
or U5890 (N_5890,N_3932,N_4115);
nand U5891 (N_5891,N_4691,N_3911);
nor U5892 (N_5892,N_2264,N_2356);
and U5893 (N_5893,N_4172,N_2669);
xor U5894 (N_5894,N_1835,N_3524);
or U5895 (N_5895,N_755,N_4089);
xnor U5896 (N_5896,N_3117,N_778);
xnor U5897 (N_5897,N_3080,N_3664);
xnor U5898 (N_5898,N_702,N_3745);
nor U5899 (N_5899,N_1420,N_2050);
or U5900 (N_5900,N_270,N_1962);
nor U5901 (N_5901,N_590,N_2054);
xnor U5902 (N_5902,N_1229,N_2064);
and U5903 (N_5903,N_1838,N_3464);
nand U5904 (N_5904,N_1505,N_4308);
or U5905 (N_5905,N_3544,N_3829);
nand U5906 (N_5906,N_3752,N_3384);
nand U5907 (N_5907,N_2640,N_1698);
or U5908 (N_5908,N_2281,N_1445);
and U5909 (N_5909,N_1923,N_697);
or U5910 (N_5910,N_2846,N_3886);
xor U5911 (N_5911,N_4942,N_1772);
nor U5912 (N_5912,N_2616,N_3651);
nand U5913 (N_5913,N_3465,N_227);
xnor U5914 (N_5914,N_4271,N_4058);
xor U5915 (N_5915,N_2675,N_3992);
xor U5916 (N_5916,N_2826,N_1349);
or U5917 (N_5917,N_1955,N_4951);
xnor U5918 (N_5918,N_1195,N_3462);
xor U5919 (N_5919,N_3721,N_3093);
xnor U5920 (N_5920,N_2421,N_387);
nand U5921 (N_5921,N_2579,N_4407);
nor U5922 (N_5922,N_2941,N_4318);
nand U5923 (N_5923,N_3569,N_3113);
or U5924 (N_5924,N_3746,N_1728);
or U5925 (N_5925,N_2609,N_2759);
xor U5926 (N_5926,N_3187,N_2784);
and U5927 (N_5927,N_4978,N_4837);
xor U5928 (N_5928,N_1877,N_4609);
and U5929 (N_5929,N_966,N_3877);
and U5930 (N_5930,N_2720,N_3007);
nand U5931 (N_5931,N_4177,N_4072);
or U5932 (N_5932,N_2656,N_3731);
and U5933 (N_5933,N_2271,N_1114);
or U5934 (N_5934,N_4719,N_3565);
or U5935 (N_5935,N_2104,N_3288);
or U5936 (N_5936,N_2731,N_3668);
nor U5937 (N_5937,N_1060,N_1241);
nor U5938 (N_5938,N_596,N_3432);
or U5939 (N_5939,N_2875,N_1330);
xnor U5940 (N_5940,N_3933,N_1775);
nand U5941 (N_5941,N_3023,N_2293);
xnor U5942 (N_5942,N_2424,N_3344);
xnor U5943 (N_5943,N_3336,N_2348);
nor U5944 (N_5944,N_4824,N_3148);
or U5945 (N_5945,N_4700,N_3863);
xor U5946 (N_5946,N_1458,N_4828);
nand U5947 (N_5947,N_2718,N_2748);
nor U5948 (N_5948,N_4210,N_603);
and U5949 (N_5949,N_3457,N_3769);
nor U5950 (N_5950,N_3227,N_3508);
or U5951 (N_5951,N_3474,N_2818);
nand U5952 (N_5952,N_3210,N_4142);
and U5953 (N_5953,N_3231,N_4368);
nand U5954 (N_5954,N_307,N_4427);
or U5955 (N_5955,N_3910,N_683);
or U5956 (N_5956,N_430,N_2319);
nand U5957 (N_5957,N_3622,N_1813);
nor U5958 (N_5958,N_4329,N_3567);
or U5959 (N_5959,N_967,N_4199);
xor U5960 (N_5960,N_2004,N_403);
xnor U5961 (N_5961,N_2606,N_2895);
nand U5962 (N_5962,N_4011,N_2299);
nand U5963 (N_5963,N_3448,N_1226);
nor U5964 (N_5964,N_2379,N_706);
or U5965 (N_5965,N_2740,N_205);
or U5966 (N_5966,N_607,N_3858);
and U5967 (N_5967,N_2762,N_1931);
nand U5968 (N_5968,N_4289,N_1798);
and U5969 (N_5969,N_221,N_2696);
and U5970 (N_5970,N_2027,N_303);
and U5971 (N_5971,N_280,N_1326);
nor U5972 (N_5972,N_1246,N_4355);
nor U5973 (N_5973,N_2760,N_3785);
nand U5974 (N_5974,N_4666,N_120);
xnor U5975 (N_5975,N_3186,N_1573);
nand U5976 (N_5976,N_4494,N_3170);
nor U5977 (N_5977,N_2896,N_1223);
nand U5978 (N_5978,N_3650,N_2690);
and U5979 (N_5979,N_3489,N_1978);
xor U5980 (N_5980,N_1768,N_432);
nor U5981 (N_5981,N_3259,N_3862);
nand U5982 (N_5982,N_1866,N_291);
and U5983 (N_5983,N_2900,N_3597);
xor U5984 (N_5984,N_336,N_4854);
xnor U5985 (N_5985,N_4364,N_768);
or U5986 (N_5986,N_1919,N_3254);
xnor U5987 (N_5987,N_4270,N_2175);
nand U5988 (N_5988,N_2707,N_4601);
xnor U5989 (N_5989,N_4553,N_3633);
and U5990 (N_5990,N_2702,N_2400);
nor U5991 (N_5991,N_2383,N_1261);
xnor U5992 (N_5992,N_2635,N_2012);
nor U5993 (N_5993,N_1271,N_4236);
and U5994 (N_5994,N_4146,N_100);
nand U5995 (N_5995,N_3060,N_1602);
nand U5996 (N_5996,N_354,N_813);
nor U5997 (N_5997,N_4415,N_1130);
nor U5998 (N_5998,N_361,N_4512);
or U5999 (N_5999,N_4440,N_4487);
nor U6000 (N_6000,N_3360,N_3838);
nor U6001 (N_6001,N_2190,N_1151);
and U6002 (N_6002,N_4276,N_1388);
xor U6003 (N_6003,N_3173,N_1634);
and U6004 (N_6004,N_4745,N_1046);
and U6005 (N_6005,N_1880,N_3065);
and U6006 (N_6006,N_3125,N_2205);
or U6007 (N_6007,N_4038,N_1737);
nor U6008 (N_6008,N_2472,N_4426);
nor U6009 (N_6009,N_616,N_1398);
nand U6010 (N_6010,N_4079,N_2235);
and U6011 (N_6011,N_3111,N_4409);
nor U6012 (N_6012,N_2243,N_4817);
nand U6013 (N_6013,N_3778,N_3468);
nor U6014 (N_6014,N_4660,N_651);
and U6015 (N_6015,N_1022,N_708);
and U6016 (N_6016,N_164,N_140);
and U6017 (N_6017,N_2395,N_1868);
nor U6018 (N_6018,N_4009,N_925);
nand U6019 (N_6019,N_2801,N_1435);
nand U6020 (N_6020,N_4651,N_1952);
and U6021 (N_6021,N_2231,N_2721);
xor U6022 (N_6022,N_3261,N_3927);
and U6023 (N_6023,N_53,N_4446);
or U6024 (N_6024,N_3248,N_4751);
xor U6025 (N_6025,N_4340,N_3003);
nor U6026 (N_6026,N_1526,N_3909);
nor U6027 (N_6027,N_988,N_3240);
xor U6028 (N_6028,N_2697,N_3193);
nand U6029 (N_6029,N_864,N_1924);
nor U6030 (N_6030,N_2045,N_4114);
xor U6031 (N_6031,N_1069,N_3399);
nor U6032 (N_6032,N_4411,N_4365);
and U6033 (N_6033,N_4505,N_3014);
and U6034 (N_6034,N_141,N_1218);
nand U6035 (N_6035,N_4592,N_1709);
and U6036 (N_6036,N_927,N_538);
xor U6037 (N_6037,N_4814,N_3626);
nor U6038 (N_6038,N_3770,N_998);
xnor U6039 (N_6039,N_4460,N_4);
xor U6040 (N_6040,N_391,N_152);
nand U6041 (N_6041,N_1601,N_4839);
or U6042 (N_6042,N_3119,N_4182);
xnor U6043 (N_6043,N_4322,N_2891);
and U6044 (N_6044,N_4578,N_486);
and U6045 (N_6045,N_1437,N_3653);
or U6046 (N_6046,N_2722,N_2363);
nor U6047 (N_6047,N_758,N_4087);
nor U6048 (N_6048,N_4158,N_3539);
and U6049 (N_6049,N_2105,N_2315);
or U6050 (N_6050,N_513,N_4858);
nor U6051 (N_6051,N_1380,N_1646);
xnor U6052 (N_6052,N_4634,N_2770);
or U6053 (N_6053,N_4860,N_675);
and U6054 (N_6054,N_1343,N_2581);
nand U6055 (N_6055,N_1404,N_3782);
xor U6056 (N_6056,N_4709,N_1563);
or U6057 (N_6057,N_2711,N_245);
or U6058 (N_6058,N_3579,N_849);
and U6059 (N_6059,N_380,N_1301);
and U6060 (N_6060,N_1622,N_4949);
or U6061 (N_6061,N_2961,N_2246);
nor U6062 (N_6062,N_1615,N_2698);
nand U6063 (N_6063,N_3332,N_1302);
nand U6064 (N_6064,N_259,N_4071);
and U6065 (N_6065,N_2289,N_1234);
nor U6066 (N_6066,N_1755,N_4740);
nand U6067 (N_6067,N_1354,N_3869);
or U6068 (N_6068,N_3677,N_3647);
xnor U6069 (N_6069,N_636,N_2422);
or U6070 (N_6070,N_4880,N_384);
nor U6071 (N_6071,N_39,N_620);
xnor U6072 (N_6072,N_159,N_4034);
and U6073 (N_6073,N_1851,N_2737);
xnor U6074 (N_6074,N_2038,N_2571);
xnor U6075 (N_6075,N_316,N_287);
nand U6076 (N_6076,N_1982,N_3559);
xnor U6077 (N_6077,N_3809,N_3424);
xnor U6078 (N_6078,N_1056,N_1359);
or U6079 (N_6079,N_2870,N_2971);
nand U6080 (N_6080,N_4963,N_805);
or U6081 (N_6081,N_4206,N_3503);
nor U6082 (N_6082,N_3072,N_3296);
nand U6083 (N_6083,N_1015,N_528);
nor U6084 (N_6084,N_2462,N_4864);
xor U6085 (N_6085,N_1213,N_4237);
nor U6086 (N_6086,N_4648,N_4192);
or U6087 (N_6087,N_3504,N_1717);
nor U6088 (N_6088,N_3242,N_1566);
nand U6089 (N_6089,N_458,N_4266);
and U6090 (N_6090,N_612,N_3410);
nor U6091 (N_6091,N_1097,N_4934);
xnor U6092 (N_6092,N_4491,N_2361);
or U6093 (N_6093,N_4390,N_118);
nor U6094 (N_6094,N_938,N_3408);
xnor U6095 (N_6095,N_290,N_1450);
or U6096 (N_6096,N_4957,N_4703);
xnor U6097 (N_6097,N_2789,N_1696);
or U6098 (N_6098,N_2117,N_3002);
or U6099 (N_6099,N_1885,N_3367);
and U6100 (N_6100,N_329,N_1377);
or U6101 (N_6101,N_2939,N_3202);
nor U6102 (N_6102,N_138,N_3067);
nor U6103 (N_6103,N_2563,N_2244);
nand U6104 (N_6104,N_570,N_649);
nand U6105 (N_6105,N_4529,N_4792);
nor U6106 (N_6106,N_283,N_4417);
or U6107 (N_6107,N_4668,N_718);
nor U6108 (N_6108,N_2141,N_853);
and U6109 (N_6109,N_4064,N_1522);
nor U6110 (N_6110,N_1886,N_1682);
nor U6111 (N_6111,N_2302,N_4300);
or U6112 (N_6112,N_3957,N_1935);
nor U6113 (N_6113,N_3054,N_2011);
and U6114 (N_6114,N_2876,N_1032);
xor U6115 (N_6115,N_854,N_1674);
and U6116 (N_6116,N_1023,N_32);
nor U6117 (N_6117,N_169,N_4280);
xor U6118 (N_6118,N_3139,N_2565);
or U6119 (N_6119,N_1425,N_633);
and U6120 (N_6120,N_1037,N_272);
and U6121 (N_6121,N_1320,N_4990);
nand U6122 (N_6122,N_4998,N_2910);
or U6123 (N_6123,N_3197,N_2531);
nor U6124 (N_6124,N_1546,N_2699);
nor U6125 (N_6125,N_4930,N_4129);
nand U6126 (N_6126,N_4499,N_761);
or U6127 (N_6127,N_484,N_924);
and U6128 (N_6128,N_3670,N_4397);
nand U6129 (N_6129,N_4024,N_3330);
and U6130 (N_6130,N_2582,N_723);
nor U6131 (N_6131,N_3767,N_3600);
nor U6132 (N_6132,N_2137,N_4083);
nor U6133 (N_6133,N_1903,N_3338);
nor U6134 (N_6134,N_4399,N_4599);
nand U6135 (N_6135,N_3530,N_2845);
nand U6136 (N_6136,N_4570,N_1258);
nand U6137 (N_6137,N_2929,N_3385);
and U6138 (N_6138,N_548,N_1576);
xnor U6139 (N_6139,N_4856,N_1512);
nand U6140 (N_6140,N_648,N_3628);
nand U6141 (N_6141,N_696,N_350);
and U6142 (N_6142,N_2189,N_2766);
or U6143 (N_6143,N_3251,N_167);
and U6144 (N_6144,N_4573,N_144);
nand U6145 (N_6145,N_1144,N_60);
nand U6146 (N_6146,N_585,N_511);
nor U6147 (N_6147,N_2336,N_2457);
or U6148 (N_6148,N_3602,N_4348);
nor U6149 (N_6149,N_216,N_451);
and U6150 (N_6150,N_3617,N_1833);
nand U6151 (N_6151,N_2551,N_3861);
nor U6152 (N_6152,N_1010,N_3522);
nand U6153 (N_6153,N_19,N_3089);
or U6154 (N_6154,N_2931,N_4154);
xor U6155 (N_6155,N_4202,N_2841);
nor U6156 (N_6156,N_3452,N_305);
xor U6157 (N_6157,N_4914,N_1252);
nand U6158 (N_6158,N_2399,N_433);
and U6159 (N_6159,N_726,N_4376);
and U6160 (N_6160,N_2439,N_242);
nor U6161 (N_6161,N_4288,N_2118);
nand U6162 (N_6162,N_3389,N_1374);
or U6163 (N_6163,N_1777,N_600);
xnor U6164 (N_6164,N_326,N_3099);
xnor U6165 (N_6165,N_4725,N_2793);
or U6166 (N_6166,N_4122,N_753);
nand U6167 (N_6167,N_2161,N_2637);
xor U6168 (N_6168,N_4807,N_3718);
nor U6169 (N_6169,N_1399,N_2262);
nor U6170 (N_6170,N_1418,N_870);
nand U6171 (N_6171,N_1292,N_4596);
xor U6172 (N_6172,N_4523,N_4036);
nand U6173 (N_6173,N_265,N_1096);
nand U6174 (N_6174,N_2010,N_4575);
xor U6175 (N_6175,N_2122,N_64);
or U6176 (N_6176,N_3774,N_4564);
or U6177 (N_6177,N_817,N_2714);
or U6178 (N_6178,N_1734,N_4111);
or U6179 (N_6179,N_2524,N_1530);
nand U6180 (N_6180,N_1842,N_921);
nor U6181 (N_6181,N_1750,N_223);
xnor U6182 (N_6182,N_4964,N_971);
and U6183 (N_6183,N_1004,N_2268);
or U6184 (N_6184,N_2562,N_2043);
nor U6185 (N_6185,N_2360,N_4107);
nor U6186 (N_6186,N_2354,N_3973);
or U6187 (N_6187,N_2171,N_3040);
nor U6188 (N_6188,N_4059,N_2479);
or U6189 (N_6189,N_4430,N_730);
or U6190 (N_6190,N_807,N_1182);
nand U6191 (N_6191,N_2265,N_2613);
nor U6192 (N_6192,N_4282,N_2541);
nand U6193 (N_6193,N_2942,N_3357);
nor U6194 (N_6194,N_68,N_58);
nand U6195 (N_6195,N_4106,N_1328);
or U6196 (N_6196,N_243,N_3541);
nor U6197 (N_6197,N_3678,N_1232);
nor U6198 (N_6198,N_3792,N_268);
or U6199 (N_6199,N_3596,N_142);
or U6200 (N_6200,N_1319,N_2263);
nor U6201 (N_6201,N_1650,N_3129);
and U6202 (N_6202,N_4229,N_2886);
and U6203 (N_6203,N_1822,N_4517);
xor U6204 (N_6204,N_248,N_4759);
nor U6205 (N_6205,N_3079,N_1845);
and U6206 (N_6206,N_3328,N_2769);
xor U6207 (N_6207,N_2671,N_946);
nor U6208 (N_6208,N_3570,N_29);
or U6209 (N_6209,N_742,N_4865);
and U6210 (N_6210,N_775,N_4641);
and U6211 (N_6211,N_3896,N_477);
nor U6212 (N_6212,N_3605,N_1307);
xor U6213 (N_6213,N_3839,N_3901);
xor U6214 (N_6214,N_4180,N_3615);
and U6215 (N_6215,N_4522,N_1915);
nor U6216 (N_6216,N_2638,N_1119);
nand U6217 (N_6217,N_877,N_3725);
and U6218 (N_6218,N_2022,N_3136);
nor U6219 (N_6219,N_1672,N_4619);
and U6220 (N_6220,N_863,N_4561);
and U6221 (N_6221,N_1447,N_2211);
and U6222 (N_6222,N_4997,N_1347);
and U6223 (N_6223,N_2853,N_1100);
nand U6224 (N_6224,N_3875,N_647);
nor U6225 (N_6225,N_1507,N_1433);
nor U6226 (N_6226,N_2787,N_2436);
nor U6227 (N_6227,N_3937,N_1999);
nor U6228 (N_6228,N_3044,N_1934);
nor U6229 (N_6229,N_1747,N_4835);
nor U6230 (N_6230,N_978,N_97);
xnor U6231 (N_6231,N_4851,N_2953);
and U6232 (N_6232,N_843,N_4887);
and U6233 (N_6233,N_3548,N_4548);
nor U6234 (N_6234,N_2960,N_3169);
and U6235 (N_6235,N_4414,N_3052);
nand U6236 (N_6236,N_2207,N_3323);
nand U6237 (N_6237,N_614,N_4498);
and U6238 (N_6238,N_1331,N_4373);
or U6239 (N_6239,N_1415,N_4774);
and U6240 (N_6240,N_4126,N_322);
nand U6241 (N_6241,N_1504,N_4151);
nand U6242 (N_6242,N_4532,N_2440);
or U6243 (N_6243,N_756,N_2326);
nand U6244 (N_6244,N_1086,N_3949);
xnor U6245 (N_6245,N_4037,N_729);
and U6246 (N_6246,N_2485,N_4082);
nand U6247 (N_6247,N_374,N_3401);
and U6248 (N_6248,N_848,N_1472);
nor U6249 (N_6249,N_1857,N_964);
nor U6250 (N_6250,N_3931,N_1946);
nand U6251 (N_6251,N_2544,N_4488);
xor U6252 (N_6252,N_4701,N_523);
xnor U6253 (N_6253,N_1284,N_219);
and U6254 (N_6254,N_2090,N_2362);
nand U6255 (N_6255,N_3849,N_707);
nor U6256 (N_6256,N_759,N_496);
xor U6257 (N_6257,N_4543,N_4031);
or U6258 (N_6258,N_429,N_952);
and U6259 (N_6259,N_313,N_2981);
or U6260 (N_6260,N_2788,N_3944);
nor U6261 (N_6261,N_3378,N_982);
or U6262 (N_6262,N_1925,N_2021);
or U6263 (N_6263,N_1555,N_66);
nor U6264 (N_6264,N_1927,N_1286);
or U6265 (N_6265,N_5,N_4077);
or U6266 (N_6266,N_1168,N_601);
nor U6267 (N_6267,N_674,N_3168);
nor U6268 (N_6268,N_2096,N_1127);
and U6269 (N_6269,N_991,N_2863);
and U6270 (N_6270,N_2068,N_3213);
and U6271 (N_6271,N_1199,N_3486);
nor U6272 (N_6272,N_4110,N_2214);
nor U6273 (N_6273,N_680,N_1558);
or U6274 (N_6274,N_618,N_3954);
nand U6275 (N_6275,N_881,N_3447);
xnor U6276 (N_6276,N_4783,N_3331);
and U6277 (N_6277,N_1035,N_401);
or U6278 (N_6278,N_2121,N_4544);
nand U6279 (N_6279,N_2967,N_525);
or U6280 (N_6280,N_2398,N_3830);
nand U6281 (N_6281,N_3237,N_3598);
nand U6282 (N_6282,N_1786,N_2);
and U6283 (N_6283,N_3053,N_3306);
nor U6284 (N_6284,N_1781,N_4103);
nand U6285 (N_6285,N_4323,N_4149);
nand U6286 (N_6286,N_4175,N_3696);
or U6287 (N_6287,N_1639,N_1158);
nand U6288 (N_6288,N_2154,N_4096);
xnor U6289 (N_6289,N_670,N_11);
nor U6290 (N_6290,N_542,N_673);
xnor U6291 (N_6291,N_827,N_119);
and U6292 (N_6292,N_3981,N_1870);
nor U6293 (N_6293,N_448,N_105);
nor U6294 (N_6294,N_1640,N_1991);
and U6295 (N_6295,N_1281,N_252);
nand U6296 (N_6296,N_3846,N_306);
nor U6297 (N_6297,N_2334,N_2974);
and U6298 (N_6298,N_731,N_3134);
xor U6299 (N_6299,N_4495,N_2728);
or U6300 (N_6300,N_302,N_655);
nand U6301 (N_6301,N_4530,N_4742);
and U6302 (N_6302,N_3970,N_3264);
and U6303 (N_6303,N_4670,N_1785);
or U6304 (N_6304,N_660,N_3088);
xor U6305 (N_6305,N_1719,N_2705);
or U6306 (N_6306,N_36,N_4794);
and U6307 (N_6307,N_1998,N_1381);
nand U6308 (N_6308,N_2417,N_1782);
xnor U6309 (N_6309,N_1222,N_3123);
and U6310 (N_6310,N_2322,N_2080);
xor U6311 (N_6311,N_250,N_2329);
and U6312 (N_6312,N_2586,N_4850);
and U6313 (N_6313,N_1920,N_2108);
xnor U6314 (N_6314,N_2552,N_4445);
xnor U6315 (N_6315,N_1748,N_745);
and U6316 (N_6316,N_4565,N_3884);
or U6317 (N_6317,N_3743,N_671);
nand U6318 (N_6318,N_4017,N_687);
xnor U6319 (N_6319,N_4992,N_3167);
xnor U6320 (N_6320,N_837,N_0);
nand U6321 (N_6321,N_3772,N_550);
nand U6322 (N_6322,N_4621,N_3959);
xor U6323 (N_6323,N_2295,N_4886);
xor U6324 (N_6324,N_3758,N_4903);
or U6325 (N_6325,N_1839,N_319);
xor U6326 (N_6326,N_3843,N_1145);
nor U6327 (N_6327,N_1293,N_1277);
and U6328 (N_6328,N_4381,N_3680);
or U6329 (N_6329,N_969,N_4993);
nand U6330 (N_6330,N_1980,N_343);
nand U6331 (N_6331,N_91,N_275);
nand U6332 (N_6332,N_4480,N_312);
xor U6333 (N_6333,N_4729,N_951);
or U6334 (N_6334,N_4459,N_835);
and U6335 (N_6335,N_3512,N_1627);
xor U6336 (N_6336,N_1030,N_4054);
or U6337 (N_6337,N_3140,N_3494);
and U6338 (N_6338,N_3870,N_1972);
xnor U6339 (N_6339,N_3195,N_258);
and U6340 (N_6340,N_4001,N_641);
or U6341 (N_6341,N_3722,N_2918);
xor U6342 (N_6342,N_1088,N_2628);
or U6343 (N_6343,N_752,N_913);
xnor U6344 (N_6344,N_1921,N_1464);
or U6345 (N_6345,N_3888,N_74);
or U6346 (N_6346,N_2834,N_4304);
nor U6347 (N_6347,N_3013,N_23);
nor U6348 (N_6348,N_1637,N_2404);
xnor U6349 (N_6349,N_2297,N_3020);
or U6350 (N_6350,N_3203,N_3018);
nand U6351 (N_6351,N_724,N_1685);
xnor U6352 (N_6352,N_2676,N_3137);
nand U6353 (N_6353,N_3037,N_1739);
xnor U6354 (N_6354,N_2508,N_960);
nand U6355 (N_6355,N_846,N_1365);
nand U6356 (N_6356,N_1605,N_2644);
nand U6357 (N_6357,N_3961,N_1367);
nor U6358 (N_6358,N_1606,N_1141);
nor U6359 (N_6359,N_4741,N_3738);
xor U6360 (N_6360,N_389,N_4625);
nand U6361 (N_6361,N_3417,N_3540);
xor U6362 (N_6362,N_4722,N_4267);
nand U6363 (N_6363,N_3916,N_4853);
and U6364 (N_6364,N_465,N_1665);
and U6365 (N_6365,N_3712,N_4167);
xnor U6366 (N_6366,N_94,N_1939);
or U6367 (N_6367,N_1021,N_369);
nand U6368 (N_6368,N_2530,N_347);
or U6369 (N_6369,N_4188,N_587);
nor U6370 (N_6370,N_1231,N_1318);
xnor U6371 (N_6371,N_4333,N_4962);
nand U6372 (N_6372,N_4453,N_3794);
xnor U6373 (N_6373,N_4673,N_2178);
nor U6374 (N_6374,N_1042,N_1743);
or U6375 (N_6375,N_4070,N_955);
nand U6376 (N_6376,N_4030,N_1057);
nor U6377 (N_6377,N_4787,N_564);
xor U6378 (N_6378,N_4775,N_1129);
xor U6379 (N_6379,N_1270,N_2733);
xnor U6380 (N_6380,N_1187,N_4643);
xnor U6381 (N_6381,N_298,N_487);
xnor U6382 (N_6382,N_3513,N_4796);
or U6383 (N_6383,N_78,N_2572);
or U6384 (N_6384,N_309,N_4256);
and U6385 (N_6385,N_1209,N_3383);
and U6386 (N_6386,N_4025,N_3883);
or U6387 (N_6387,N_3151,N_860);
or U6388 (N_6388,N_3906,N_2522);
nor U6389 (N_6389,N_2504,N_3709);
nand U6390 (N_6390,N_388,N_471);
and U6391 (N_6391,N_1893,N_208);
and U6392 (N_6392,N_407,N_1888);
nor U6393 (N_6393,N_202,N_3154);
or U6394 (N_6394,N_1332,N_2520);
xor U6395 (N_6395,N_3318,N_3697);
nand U6396 (N_6396,N_2928,N_378);
xor U6397 (N_6397,N_2413,N_3533);
or U6398 (N_6398,N_2836,N_3310);
xnor U6399 (N_6399,N_4100,N_2125);
xor U6400 (N_6400,N_1456,N_1741);
nor U6401 (N_6401,N_1953,N_2871);
and U6402 (N_6402,N_4825,N_2992);
nand U6403 (N_6403,N_3375,N_262);
or U6404 (N_6404,N_3661,N_4504);
nand U6405 (N_6405,N_2890,N_4943);
or U6406 (N_6406,N_4770,N_3142);
or U6407 (N_6407,N_2680,N_80);
nor U6408 (N_6408,N_1117,N_2617);
or U6409 (N_6409,N_534,N_2433);
nand U6410 (N_6410,N_4554,N_591);
and U6411 (N_6411,N_2631,N_2444);
nand U6412 (N_6412,N_4899,N_945);
xor U6413 (N_6413,N_115,N_2950);
xor U6414 (N_6414,N_4622,N_3868);
or U6415 (N_6415,N_1973,N_3977);
nand U6416 (N_6416,N_3936,N_4905);
xnor U6417 (N_6417,N_3506,N_4016);
nor U6418 (N_6418,N_1269,N_452);
or U6419 (N_6419,N_2792,N_2608);
and U6420 (N_6420,N_4432,N_777);
xor U6421 (N_6421,N_1583,N_2963);
and U6422 (N_6422,N_2817,N_4508);
xor U6423 (N_6423,N_2761,N_3372);
or U6424 (N_6424,N_1397,N_3177);
xor U6425 (N_6425,N_1449,N_3006);
nor U6426 (N_6426,N_2936,N_1810);
nor U6427 (N_6427,N_2949,N_4536);
nor U6428 (N_6428,N_504,N_1260);
xor U6429 (N_6429,N_2629,N_2151);
xnor U6430 (N_6430,N_3733,N_4339);
and U6431 (N_6431,N_2008,N_4273);
or U6432 (N_6432,N_1528,N_4640);
xnor U6433 (N_6433,N_4283,N_4802);
xor U6434 (N_6434,N_3543,N_2252);
nand U6435 (N_6435,N_3308,N_2709);
and U6436 (N_6436,N_4279,N_3599);
or U6437 (N_6437,N_885,N_694);
xnor U6438 (N_6438,N_819,N_4910);
or U6439 (N_6439,N_1616,N_1395);
nand U6440 (N_6440,N_606,N_251);
nand U6441 (N_6441,N_4711,N_3469);
and U6442 (N_6442,N_419,N_1928);
or U6443 (N_6443,N_2069,N_830);
nor U6444 (N_6444,N_8,N_3024);
or U6445 (N_6445,N_55,N_4928);
nor U6446 (N_6446,N_578,N_13);
nor U6447 (N_6447,N_4053,N_2958);
nand U6448 (N_6448,N_1827,N_1442);
or U6449 (N_6449,N_2605,N_1061);
and U6450 (N_6450,N_3879,N_3629);
xor U6451 (N_6451,N_2062,N_1965);
xor U6452 (N_6452,N_2049,N_2888);
and U6453 (N_6453,N_4341,N_3351);
or U6454 (N_6454,N_609,N_4043);
or U6455 (N_6455,N_1533,N_2518);
xor U6456 (N_6456,N_4597,N_767);
xor U6457 (N_6457,N_172,N_2827);
xor U6458 (N_6458,N_2065,N_2197);
nor U6459 (N_6459,N_2560,N_4141);
nand U6460 (N_6460,N_2453,N_866);
nand U6461 (N_6461,N_2892,N_3976);
or U6462 (N_6462,N_2820,N_2044);
and U6463 (N_6463,N_2691,N_2903);
xnor U6464 (N_6464,N_4404,N_393);
and U6465 (N_6465,N_2040,N_3810);
and U6466 (N_6466,N_2786,N_4600);
and U6467 (N_6467,N_4080,N_1706);
xor U6468 (N_6468,N_3646,N_4518);
xnor U6469 (N_6469,N_3791,N_4572);
and U6470 (N_6470,N_919,N_2877);
or U6471 (N_6471,N_263,N_2811);
xnor U6472 (N_6472,N_2837,N_857);
or U6473 (N_6473,N_720,N_1556);
nand U6474 (N_6474,N_1974,N_4303);
nor U6475 (N_6475,N_980,N_3015);
or U6476 (N_6476,N_4808,N_1988);
nor U6477 (N_6477,N_2539,N_4345);
or U6478 (N_6478,N_4840,N_3153);
and U6479 (N_6479,N_801,N_1630);
or U6480 (N_6480,N_4922,N_3912);
and U6481 (N_6481,N_4987,N_2291);
or U6482 (N_6482,N_4428,N_4450);
and U6483 (N_6483,N_4481,N_4391);
nand U6484 (N_6484,N_1525,N_1618);
or U6485 (N_6485,N_532,N_3781);
xor U6486 (N_6486,N_2983,N_456);
and U6487 (N_6487,N_2765,N_3679);
xnor U6488 (N_6488,N_704,N_1854);
nand U6489 (N_6489,N_1968,N_774);
nor U6490 (N_6490,N_1487,N_4520);
nor U6491 (N_6491,N_2306,N_2425);
and U6492 (N_6492,N_2985,N_3208);
xor U6493 (N_6493,N_878,N_2621);
and U6494 (N_6494,N_4098,N_1787);
and U6495 (N_6495,N_852,N_4153);
and U6496 (N_6496,N_1648,N_4191);
nor U6497 (N_6497,N_3546,N_2823);
and U6498 (N_6498,N_2318,N_3586);
nor U6499 (N_6499,N_4502,N_4654);
nor U6500 (N_6500,N_104,N_3703);
xor U6501 (N_6501,N_4739,N_4785);
and U6502 (N_6502,N_4361,N_1803);
nor U6503 (N_6503,N_2864,N_2933);
or U6504 (N_6504,N_2298,N_1510);
nand U6505 (N_6505,N_1170,N_3229);
nor U6506 (N_6506,N_2032,N_2975);
nor U6507 (N_6507,N_3185,N_2956);
nand U6508 (N_6508,N_1588,N_2331);
nor U6509 (N_6509,N_4646,N_3329);
or U6510 (N_6510,N_4873,N_2229);
nand U6511 (N_6511,N_1621,N_3952);
or U6512 (N_6512,N_4972,N_1770);
nand U6513 (N_6513,N_2944,N_2469);
xnor U6514 (N_6514,N_3075,N_2483);
xnor U6515 (N_6515,N_2940,N_1807);
xor U6516 (N_6516,N_200,N_4710);
nor U6517 (N_6517,N_540,N_1976);
nor U6518 (N_6518,N_780,N_4707);
and U6519 (N_6519,N_1296,N_1864);
and U6520 (N_6520,N_4545,N_2677);
and U6521 (N_6521,N_4105,N_4908);
and U6522 (N_6522,N_2785,N_2351);
or U6523 (N_6523,N_2819,N_1600);
nor U6524 (N_6524,N_828,N_1167);
nand U6525 (N_6525,N_2461,N_2389);
nor U6526 (N_6526,N_476,N_3790);
nand U6527 (N_6527,N_4343,N_123);
nand U6528 (N_6528,N_2754,N_1687);
and U6529 (N_6529,N_3364,N_3207);
xnor U6530 (N_6530,N_1823,N_3532);
or U6531 (N_6531,N_409,N_725);
or U6532 (N_6532,N_2184,N_2533);
nor U6533 (N_6533,N_3659,N_1184);
or U6534 (N_6534,N_4642,N_1204);
nor U6535 (N_6535,N_785,N_1389);
and U6536 (N_6536,N_4755,N_4136);
nor U6537 (N_6537,N_4325,N_2491);
nor U6538 (N_6538,N_3204,N_155);
or U6539 (N_6539,N_4335,N_3893);
or U6540 (N_6540,N_2612,N_1795);
and U6541 (N_6541,N_1203,N_2047);
nor U6542 (N_6542,N_1517,N_1342);
xnor U6543 (N_6543,N_1751,N_4045);
or U6544 (N_6544,N_4328,N_1662);
nor U6545 (N_6545,N_4392,N_1889);
nor U6546 (N_6546,N_1194,N_1895);
xnor U6547 (N_6547,N_654,N_544);
xnor U6548 (N_6548,N_1413,N_3069);
nor U6549 (N_6549,N_2780,N_1104);
xnor U6550 (N_6550,N_3160,N_1676);
and U6551 (N_6551,N_782,N_1596);
nand U6552 (N_6552,N_3257,N_531);
nand U6553 (N_6553,N_2063,N_2494);
or U6554 (N_6554,N_4190,N_1159);
and U6555 (N_6555,N_4268,N_4605);
nand U6556 (N_6556,N_2480,N_2403);
or U6557 (N_6557,N_3175,N_4849);
nand U6558 (N_6558,N_4076,N_1697);
xnor U6559 (N_6559,N_3191,N_915);
and U6560 (N_6560,N_2344,N_3368);
nand U6561 (N_6561,N_1215,N_4047);
and U6562 (N_6562,N_4032,N_588);
or U6563 (N_6563,N_376,N_4297);
or U6564 (N_6564,N_2925,N_2599);
and U6565 (N_6565,N_182,N_344);
nor U6566 (N_6566,N_4284,N_2790);
xor U6567 (N_6567,N_2378,N_996);
xnor U6568 (N_6568,N_4108,N_613);
xor U6569 (N_6569,N_3285,N_3689);
xnor U6570 (N_6570,N_3835,N_2455);
nor U6571 (N_6571,N_3216,N_4470);
nand U6572 (N_6572,N_4216,N_2497);
and U6573 (N_6573,N_2057,N_3122);
or U6574 (N_6574,N_3637,N_2502);
or U6575 (N_6575,N_4162,N_3620);
nor U6576 (N_6576,N_2501,N_3295);
or U6577 (N_6577,N_463,N_3436);
nor U6578 (N_6578,N_2055,N_1038);
and U6579 (N_6579,N_4228,N_1409);
nand U6580 (N_6580,N_1457,N_3749);
nor U6581 (N_6581,N_698,N_4857);
or U6582 (N_6582,N_712,N_3915);
nand U6583 (N_6583,N_453,N_643);
nor U6584 (N_6584,N_4793,N_112);
and U6585 (N_6585,N_1735,N_4714);
or U6586 (N_6586,N_1236,N_2454);
xnor U6587 (N_6587,N_1604,N_2738);
or U6588 (N_6588,N_3736,N_4984);
nor U6589 (N_6589,N_2803,N_1200);
or U6590 (N_6590,N_468,N_1183);
xnor U6591 (N_6591,N_2528,N_858);
and U6592 (N_6592,N_2685,N_789);
nand U6593 (N_6593,N_2882,N_4462);
or U6594 (N_6594,N_1383,N_1174);
xor U6595 (N_6595,N_4015,N_2407);
nor U6596 (N_6596,N_3070,N_3249);
nand U6597 (N_6597,N_134,N_3706);
nand U6598 (N_6598,N_1077,N_160);
or U6599 (N_6599,N_3607,N_3684);
nor U6600 (N_6600,N_3918,N_2526);
xnor U6601 (N_6601,N_4623,N_3263);
or U6602 (N_6602,N_4533,N_125);
or U6603 (N_6603,N_4492,N_2719);
nor U6604 (N_6604,N_4882,N_2647);
or U6605 (N_6605,N_2181,N_1008);
xnor U6606 (N_6606,N_3939,N_791);
nor U6607 (N_6607,N_4938,N_4198);
or U6608 (N_6608,N_467,N_1083);
xor U6609 (N_6609,N_4946,N_1147);
xnor U6610 (N_6610,N_1797,N_1001);
nand U6611 (N_6611,N_3349,N_3729);
nor U6612 (N_6612,N_4664,N_2947);
nand U6613 (N_6613,N_2358,N_1484);
xnor U6614 (N_6614,N_757,N_3760);
xnor U6615 (N_6615,N_1959,N_254);
nor U6616 (N_6616,N_1989,N_3719);
and U6617 (N_6617,N_2923,N_4029);
or U6618 (N_6618,N_236,N_4295);
nand U6619 (N_6619,N_2694,N_153);
nand U6620 (N_6620,N_905,N_4320);
or U6621 (N_6621,N_1238,N_2456);
or U6622 (N_6622,N_4798,N_1305);
nand U6623 (N_6623,N_3609,N_3042);
or U6624 (N_6624,N_2751,N_619);
and U6625 (N_6625,N_3744,N_4378);
or U6626 (N_6626,N_4449,N_1350);
or U6627 (N_6627,N_472,N_536);
or U6628 (N_6628,N_2990,N_3495);
and U6629 (N_6629,N_2020,N_193);
or U6630 (N_6630,N_798,N_267);
and U6631 (N_6631,N_555,N_2239);
and U6632 (N_6632,N_2584,N_4836);
nor U6633 (N_6633,N_4163,N_2408);
xor U6634 (N_6634,N_4226,N_1373);
nor U6635 (N_6635,N_719,N_1636);
nand U6636 (N_6636,N_3922,N_3126);
nor U6637 (N_6637,N_4861,N_4379);
xor U6638 (N_6638,N_2053,N_4467);
and U6639 (N_6639,N_4587,N_2729);
nor U6640 (N_6640,N_2106,N_416);
or U6641 (N_6641,N_2130,N_2824);
and U6642 (N_6642,N_311,N_3341);
or U6643 (N_6643,N_3685,N_1053);
or U6644 (N_6644,N_3380,N_4588);
or U6645 (N_6645,N_3739,N_203);
nand U6646 (N_6646,N_1120,N_1703);
and U6647 (N_6647,N_88,N_4312);
and U6648 (N_6648,N_2423,N_4593);
and U6649 (N_6649,N_373,N_2048);
or U6650 (N_6650,N_2833,N_4482);
nor U6651 (N_6651,N_4692,N_2773);
xnor U6652 (N_6652,N_2715,N_1975);
nand U6653 (N_6653,N_3500,N_2202);
xnor U6654 (N_6654,N_678,N_1577);
xnor U6655 (N_6655,N_3286,N_4541);
and U6656 (N_6656,N_4715,N_3925);
nor U6657 (N_6657,N_355,N_3496);
nand U6658 (N_6658,N_106,N_1836);
nor U6659 (N_6659,N_1499,N_3028);
or U6660 (N_6660,N_4624,N_1700);
or U6661 (N_6661,N_3236,N_3161);
nand U6662 (N_6662,N_1679,N_2904);
nand U6663 (N_6663,N_956,N_288);
or U6664 (N_6664,N_2777,N_4528);
xor U6665 (N_6665,N_3150,N_4974);
xor U6666 (N_6666,N_3928,N_3968);
and U6667 (N_6667,N_4116,N_1567);
and U6668 (N_6668,N_1268,N_4321);
nor U6669 (N_6669,N_3676,N_2238);
or U6670 (N_6670,N_4380,N_3048);
or U6671 (N_6671,N_308,N_2394);
or U6672 (N_6672,N_1303,N_1256);
xnor U6673 (N_6673,N_1353,N_3059);
nand U6674 (N_6674,N_2499,N_4826);
or U6675 (N_6675,N_541,N_4073);
and U6676 (N_6676,N_1039,N_3078);
and U6677 (N_6677,N_3097,N_840);
and U6678 (N_6678,N_2303,N_4090);
nor U6679 (N_6679,N_1228,N_3674);
or U6680 (N_6680,N_482,N_4401);
or U6681 (N_6681,N_3582,N_2210);
xnor U6682 (N_6682,N_4353,N_4546);
xor U6683 (N_6683,N_993,N_901);
or U6684 (N_6684,N_926,N_423);
or U6685 (N_6685,N_2313,N_2492);
nand U6686 (N_6686,N_2412,N_1638);
and U6687 (N_6687,N_2236,N_96);
or U6688 (N_6688,N_2965,N_1623);
nand U6689 (N_6689,N_4274,N_1933);
nor U6690 (N_6690,N_438,N_4682);
nand U6691 (N_6691,N_634,N_834);
nor U6692 (N_6692,N_2375,N_1699);
or U6693 (N_6693,N_1570,N_3784);
and U6694 (N_6694,N_4677,N_3124);
and U6695 (N_6695,N_944,N_4681);
nand U6696 (N_6696,N_3623,N_4258);
and U6697 (N_6697,N_2088,N_1829);
nor U6698 (N_6698,N_3845,N_1251);
or U6699 (N_6699,N_1055,N_3978);
nor U6700 (N_6700,N_3890,N_2073);
nand U6701 (N_6701,N_4870,N_1559);
xor U6702 (N_6702,N_4478,N_3657);
xnor U6703 (N_6703,N_3994,N_3951);
xor U6704 (N_6704,N_1837,N_2101);
nand U6705 (N_6705,N_4772,N_2441);
xor U6706 (N_6706,N_2058,N_3831);
and U6707 (N_6707,N_3293,N_3470);
xnor U6708 (N_6708,N_364,N_2596);
nand U6709 (N_6709,N_4507,N_4812);
xor U6710 (N_6710,N_2767,N_1068);
nand U6711 (N_6711,N_192,N_3026);
and U6712 (N_6712,N_2294,N_4674);
nand U6713 (N_6713,N_3090,N_1424);
xnor U6714 (N_6714,N_3588,N_652);
or U6715 (N_6715,N_3017,N_332);
or U6716 (N_6716,N_1111,N_4035);
and U6717 (N_6717,N_4386,N_2580);
or U6718 (N_6718,N_2143,N_2468);
and U6719 (N_6719,N_2532,N_3806);
xor U6720 (N_6720,N_3899,N_1902);
nor U6721 (N_6721,N_4750,N_882);
and U6722 (N_6722,N_974,N_1429);
xnor U6723 (N_6723,N_2377,N_189);
and U6724 (N_6724,N_4979,N_965);
xnor U6725 (N_6725,N_1378,N_2951);
nand U6726 (N_6726,N_4558,N_4999);
or U6727 (N_6727,N_1932,N_269);
and U6728 (N_6728,N_4923,N_4239);
or U6729 (N_6729,N_2103,N_385);
nand U6730 (N_6730,N_1323,N_4443);
xnor U6731 (N_6731,N_626,N_3381);
nor U6732 (N_6732,N_3723,N_4912);
or U6733 (N_6733,N_3610,N_2201);
or U6734 (N_6734,N_2982,N_226);
nand U6735 (N_6735,N_449,N_4782);
xnor U6736 (N_6736,N_1585,N_2114);
xnor U6737 (N_6737,N_1156,N_2570);
or U6738 (N_6738,N_4953,N_623);
and U6739 (N_6739,N_4645,N_1014);
nor U6740 (N_6740,N_1178,N_2415);
and U6741 (N_6741,N_1805,N_4947);
xor U6742 (N_6742,N_1254,N_3409);
or U6743 (N_6743,N_33,N_2330);
and U6744 (N_6744,N_4855,N_2144);
xor U6745 (N_6745,N_2822,N_936);
nand U6746 (N_6746,N_1720,N_4435);
nor U6747 (N_6747,N_2730,N_1334);
nor U6748 (N_6748,N_4602,N_1392);
and U6749 (N_6749,N_820,N_3549);
nor U6750 (N_6750,N_4967,N_3563);
or U6751 (N_6751,N_4155,N_3833);
xor U6752 (N_6752,N_2274,N_3303);
xnor U6753 (N_6753,N_229,N_4892);
nand U6754 (N_6754,N_986,N_3854);
xor U6755 (N_6755,N_198,N_1643);
or U6756 (N_6756,N_679,N_480);
xor U6757 (N_6757,N_25,N_810);
xor U6758 (N_6758,N_3414,N_1716);
or U6759 (N_6759,N_1308,N_1704);
and U6760 (N_6760,N_4862,N_917);
and U6761 (N_6761,N_1762,N_1865);
and U6762 (N_6762,N_624,N_2487);
and U6763 (N_6763,N_976,N_2232);
or U6764 (N_6764,N_3107,N_4629);
and U6765 (N_6765,N_1779,N_1115);
nor U6766 (N_6766,N_122,N_1575);
nand U6767 (N_6767,N_4186,N_418);
nor U6768 (N_6768,N_264,N_1073);
xor U6769 (N_6769,N_4831,N_2716);
or U6770 (N_6770,N_605,N_4551);
and U6771 (N_6771,N_3290,N_2620);
or U6772 (N_6772,N_1290,N_2097);
and U6773 (N_6773,N_784,N_667);
nand U6774 (N_6774,N_260,N_2212);
xor U6775 (N_6775,N_1212,N_3814);
nand U6776 (N_6776,N_929,N_795);
xor U6777 (N_6777,N_642,N_2305);
nor U6778 (N_6778,N_2277,N_2465);
and U6779 (N_6779,N_4513,N_4366);
and U6780 (N_6780,N_2353,N_358);
nand U6781 (N_6781,N_1984,N_4687);
xor U6782 (N_6782,N_3681,N_1635);
and U6783 (N_6783,N_4696,N_3396);
nor U6784 (N_6784,N_4360,N_1993);
xor U6785 (N_6785,N_1071,N_1058);
and U6786 (N_6786,N_1549,N_663);
and U6787 (N_6787,N_1329,N_770);
or U6788 (N_6788,N_3282,N_2431);
xnor U6789 (N_6789,N_1491,N_2610);
nor U6790 (N_6790,N_1560,N_334);
nand U6791 (N_6791,N_199,N_833);
or U6792 (N_6792,N_4209,N_4616);
or U6793 (N_6793,N_495,N_1112);
or U6794 (N_6794,N_2409,N_3214);
or U6795 (N_6795,N_166,N_1052);
or U6796 (N_6796,N_386,N_808);
and U6797 (N_6797,N_196,N_3796);
or U6798 (N_6798,N_3118,N_1113);
and U6799 (N_6799,N_871,N_4989);
and U6800 (N_6800,N_4104,N_1511);
nor U6801 (N_6801,N_2805,N_1691);
or U6802 (N_6802,N_880,N_4563);
nand U6803 (N_6803,N_1995,N_4580);
nand U6804 (N_6804,N_4626,N_1095);
nand U6805 (N_6805,N_1110,N_2346);
nor U6806 (N_6806,N_3765,N_3583);
and U6807 (N_6807,N_2077,N_3480);
nand U6808 (N_6808,N_3100,N_2829);
or U6809 (N_6809,N_3529,N_1376);
or U6810 (N_6810,N_3836,N_3536);
xnor U6811 (N_6811,N_1489,N_179);
xnor U6812 (N_6812,N_3905,N_1756);
xor U6813 (N_6813,N_1752,N_844);
or U6814 (N_6814,N_3737,N_1561);
nor U6815 (N_6815,N_4039,N_1250);
xor U6816 (N_6816,N_4526,N_1554);
xor U6817 (N_6817,N_3291,N_1313);
and U6818 (N_6818,N_3133,N_4486);
xor U6819 (N_6819,N_3852,N_1711);
xnor U6820 (N_6820,N_4931,N_4815);
or U6821 (N_6821,N_3057,N_4455);
nor U6822 (N_6822,N_4728,N_3860);
or U6823 (N_6823,N_997,N_1557);
and U6824 (N_6824,N_2652,N_3273);
or U6825 (N_6825,N_3356,N_4688);
and U6826 (N_6826,N_3475,N_3577);
or U6827 (N_6827,N_1027,N_4092);
nand U6828 (N_6828,N_2387,N_659);
xnor U6829 (N_6829,N_1090,N_2234);
xor U6830 (N_6830,N_371,N_4010);
and U6831 (N_6831,N_669,N_121);
nand U6832 (N_6832,N_2869,N_2517);
nand U6833 (N_6833,N_1904,N_1654);
xor U6834 (N_6834,N_1316,N_1452);
nand U6835 (N_6835,N_2619,N_2311);
nand U6836 (N_6836,N_390,N_1355);
xnor U6837 (N_6837,N_4382,N_4712);
or U6838 (N_6838,N_3094,N_2323);
xor U6839 (N_6839,N_2977,N_63);
nand U6840 (N_6840,N_3347,N_4145);
nor U6841 (N_6841,N_1263,N_101);
xnor U6842 (N_6842,N_1690,N_1960);
and U6843 (N_6843,N_3517,N_4181);
nand U6844 (N_6844,N_2165,N_895);
nor U6845 (N_6845,N_2194,N_822);
and U6846 (N_6846,N_3373,N_2735);
nand U6847 (N_6847,N_4245,N_1642);
and U6848 (N_6848,N_2310,N_1677);
nor U6849 (N_6849,N_2018,N_381);
nor U6850 (N_6850,N_3423,N_4603);
or U6851 (N_6851,N_1327,N_4926);
or U6852 (N_6852,N_3938,N_3333);
nand U6853 (N_6853,N_1475,N_1763);
xor U6854 (N_6854,N_2286,N_1315);
nor U6855 (N_6855,N_341,N_4569);
xor U6856 (N_6856,N_1441,N_958);
nand U6857 (N_6857,N_2332,N_4534);
nand U6858 (N_6858,N_87,N_664);
or U6859 (N_6859,N_2309,N_722);
or U6860 (N_6860,N_3298,N_3971);
nor U6861 (N_6861,N_3802,N_4878);
nand U6862 (N_6862,N_3434,N_4866);
nand U6863 (N_6863,N_1265,N_4848);
nor U6864 (N_6864,N_4594,N_3224);
xor U6865 (N_6865,N_2206,N_4846);
or U6866 (N_6866,N_2794,N_2335);
or U6867 (N_6867,N_1957,N_2242);
nand U6868 (N_6868,N_4159,N_592);
or U6869 (N_6869,N_4362,N_1620);
nand U6870 (N_6870,N_4811,N_1722);
nor U6871 (N_6871,N_2123,N_4313);
nand U6872 (N_6872,N_845,N_1749);
or U6873 (N_6873,N_1002,N_382);
or U6874 (N_6874,N_4124,N_1983);
nor U6875 (N_6875,N_2659,N_1495);
and U6876 (N_6876,N_1598,N_4766);
nor U6877 (N_6877,N_1443,N_961);
nor U6878 (N_6878,N_656,N_869);
and U6879 (N_6879,N_170,N_814);
nor U6880 (N_6880,N_3547,N_2800);
nor U6881 (N_6881,N_3940,N_3157);
or U6882 (N_6882,N_3671,N_3217);
and U6883 (N_6883,N_2964,N_2438);
nand U6884 (N_6884,N_2813,N_214);
or U6885 (N_6885,N_1597,N_1253);
xnor U6886 (N_6886,N_518,N_4649);
nand U6887 (N_6887,N_695,N_1824);
nand U6888 (N_6888,N_1922,N_3889);
or U6889 (N_6889,N_615,N_2999);
xor U6890 (N_6890,N_3754,N_574);
nand U6891 (N_6891,N_4560,N_1054);
nor U6892 (N_6892,N_1882,N_4813);
nand U6893 (N_6893,N_3071,N_1470);
xnor U6894 (N_6894,N_4598,N_3566);
nor U6895 (N_6895,N_764,N_340);
or U6896 (N_6896,N_3479,N_1000);
and U6897 (N_6897,N_521,N_237);
and U6898 (N_6898,N_2419,N_4778);
xnor U6899 (N_6899,N_1490,N_4137);
nand U6900 (N_6900,N_3394,N_1224);
and U6901 (N_6901,N_481,N_317);
and U6902 (N_6902,N_1009,N_4744);
or U6903 (N_6903,N_3135,N_1371);
nand U6904 (N_6904,N_3038,N_559);
and U6905 (N_6905,N_4764,N_4023);
or U6906 (N_6906,N_2420,N_3666);
nor U6907 (N_6907,N_108,N_2695);
and U6908 (N_6908,N_1468,N_1410);
or U6909 (N_6909,N_1655,N_439);
nor U6910 (N_6910,N_2374,N_3714);
nand U6911 (N_6911,N_577,N_3233);
nand U6912 (N_6912,N_686,N_1949);
xor U6913 (N_6913,N_1483,N_3019);
and U6914 (N_6914,N_2758,N_4285);
nor U6915 (N_6915,N_4065,N_4007);
or U6916 (N_6916,N_981,N_4262);
xor U6917 (N_6917,N_1143,N_2919);
nand U6918 (N_6918,N_3269,N_1695);
and U6919 (N_6919,N_4296,N_681);
and U6920 (N_6920,N_2046,N_1771);
xnor U6921 (N_6921,N_2510,N_3194);
or U6922 (N_6922,N_1997,N_1448);
or U6923 (N_6923,N_2109,N_1849);
xor U6924 (N_6924,N_3663,N_537);
and U6925 (N_6925,N_2536,N_2750);
nand U6926 (N_6926,N_4475,N_4018);
and U6927 (N_6927,N_4299,N_4033);
and U6928 (N_6928,N_1689,N_1340);
xor U6929 (N_6929,N_426,N_4218);
and U6930 (N_6930,N_3334,N_899);
nor U6931 (N_6931,N_2540,N_176);
nand U6932 (N_6932,N_2550,N_3440);
nand U6933 (N_6933,N_1550,N_3219);
or U6934 (N_6934,N_1990,N_3484);
nor U6935 (N_6935,N_3631,N_3576);
or U6936 (N_6936,N_2033,N_4503);
and U6937 (N_6937,N_4669,N_3152);
nor U6938 (N_6938,N_9,N_4896);
nor U6939 (N_6939,N_3366,N_3180);
nor U6940 (N_6940,N_3700,N_187);
and U6941 (N_6941,N_42,N_3033);
nand U6942 (N_6942,N_4637,N_1382);
and U6943 (N_6943,N_2023,N_2725);
xor U6944 (N_6944,N_2135,N_4702);
and U6945 (N_6945,N_2727,N_2848);
nand U6946 (N_6946,N_3551,N_893);
nor U6947 (N_6947,N_2804,N_434);
xor U6948 (N_6948,N_3132,N_2174);
xnor U6949 (N_6949,N_1651,N_2651);
nand U6950 (N_6950,N_2588,N_2443);
and U6951 (N_6951,N_902,N_150);
and U6952 (N_6952,N_2110,N_1629);
or U6953 (N_6953,N_545,N_353);
xor U6954 (N_6954,N_4431,N_2995);
xnor U6955 (N_6955,N_2575,N_4342);
xnor U6956 (N_6956,N_4125,N_621);
nand U6957 (N_6957,N_1494,N_3613);
nor U6958 (N_6958,N_2815,N_497);
and U6959 (N_6959,N_4678,N_2634);
or U6960 (N_6960,N_1050,N_3066);
nand U6961 (N_6961,N_1240,N_4525);
and U6962 (N_6962,N_178,N_3975);
and U6963 (N_6963,N_1153,N_3672);
nor U6964 (N_6964,N_3201,N_3828);
or U6965 (N_6965,N_2185,N_3589);
xnor U6966 (N_6966,N_1515,N_4344);
nand U6967 (N_6967,N_4230,N_1363);
and U6968 (N_6968,N_4871,N_4519);
xor U6969 (N_6969,N_318,N_947);
or U6970 (N_6970,N_2662,N_3114);
nor U6971 (N_6971,N_1405,N_3459);
nor U6972 (N_6972,N_1427,N_3455);
xnor U6973 (N_6973,N_3880,N_3262);
xor U6974 (N_6974,N_4091,N_2083);
nor U6975 (N_6975,N_174,N_4123);
nand U6976 (N_6976,N_2922,N_404);
xor U6977 (N_6977,N_851,N_2673);
xnor U6978 (N_6978,N_3708,N_4264);
and U6979 (N_6979,N_3815,N_2489);
nor U6980 (N_6980,N_1936,N_855);
xor U6981 (N_6981,N_230,N_2282);
and U6982 (N_6982,N_3215,N_40);
or U6983 (N_6983,N_1031,N_3891);
or U6984 (N_6984,N_2937,N_293);
xnor U6985 (N_6985,N_3948,N_2683);
nor U6986 (N_6986,N_2678,N_4804);
xnor U6987 (N_6987,N_175,N_1784);
nor U6988 (N_6988,N_4479,N_2025);
xor U6989 (N_6989,N_4995,N_4852);
nor U6990 (N_6990,N_2327,N_3636);
nor U6991 (N_6991,N_4384,N_4822);
and U6992 (N_6992,N_2102,N_147);
xor U6993 (N_6993,N_3812,N_4763);
nand U6994 (N_6994,N_1278,N_1872);
xnor U6995 (N_6995,N_1337,N_4547);
or U6996 (N_6996,N_4003,N_2573);
nor U6997 (N_6997,N_1172,N_4925);
xor U6998 (N_6998,N_546,N_1914);
or U6999 (N_6999,N_1282,N_398);
nor U7000 (N_7000,N_1132,N_3635);
nor U7001 (N_7001,N_3941,N_349);
and U7002 (N_7002,N_3604,N_1705);
and U7003 (N_7003,N_1776,N_4618);
nand U7004 (N_7004,N_1981,N_923);
or U7005 (N_7005,N_4966,N_490);
xnor U7006 (N_7006,N_1956,N_3000);
nor U7007 (N_7007,N_599,N_4008);
nand U7008 (N_7008,N_2884,N_4644);
or U7009 (N_7009,N_3930,N_2061);
or U7010 (N_7010,N_2251,N_224);
or U7011 (N_7011,N_4713,N_4260);
xor U7012 (N_7012,N_903,N_2092);
nand U7013 (N_7013,N_3612,N_14);
nand U7014 (N_7014,N_3805,N_4693);
nor U7015 (N_7015,N_2632,N_796);
nor U7016 (N_7016,N_1543,N_1544);
nor U7017 (N_7017,N_3834,N_4868);
nor U7018 (N_7018,N_4140,N_1025);
nand U7019 (N_7019,N_4918,N_3983);
nor U7020 (N_7020,N_4048,N_2623);
nor U7021 (N_7021,N_4983,N_950);
xor U7022 (N_7022,N_4062,N_4352);
xnor U7023 (N_7023,N_1641,N_1149);
or U7024 (N_7024,N_1081,N_2567);
xnor U7025 (N_7025,N_2116,N_1659);
xor U7026 (N_7026,N_4248,N_715);
xnor U7027 (N_7027,N_676,N_454);
or U7028 (N_7028,N_732,N_466);
and U7029 (N_7029,N_2000,N_3803);
nor U7030 (N_7030,N_2732,N_2006);
or U7031 (N_7031,N_2430,N_1736);
and U7032 (N_7032,N_2668,N_1396);
and U7033 (N_7033,N_2872,N_149);
or U7034 (N_7034,N_1136,N_597);
and U7035 (N_7035,N_4509,N_1109);
and U7036 (N_7036,N_2945,N_914);
and U7037 (N_7037,N_1006,N_2816);
xnor U7038 (N_7038,N_2901,N_1085);
nor U7039 (N_7039,N_2598,N_4732);
or U7040 (N_7040,N_1502,N_975);
and U7041 (N_7041,N_569,N_3979);
nand U7042 (N_7042,N_1339,N_314);
or U7043 (N_7043,N_195,N_1506);
and U7044 (N_7044,N_148,N_787);
xor U7045 (N_7045,N_2300,N_4559);
or U7046 (N_7046,N_1547,N_3824);
and U7047 (N_7047,N_1391,N_1986);
and U7048 (N_7048,N_4706,N_3300);
nand U7049 (N_7049,N_4562,N_4939);
nor U7050 (N_7050,N_3523,N_2449);
nand U7051 (N_7051,N_2952,N_2887);
xnor U7052 (N_7052,N_3643,N_2471);
nor U7053 (N_7053,N_571,N_507);
xnor U7054 (N_7054,N_4694,N_3127);
or U7055 (N_7055,N_2017,N_4456);
or U7056 (N_7056,N_2537,N_3980);
or U7057 (N_7057,N_1861,N_2285);
xnor U7058 (N_7058,N_1366,N_1309);
xor U7059 (N_7059,N_2547,N_1801);
or U7060 (N_7060,N_2269,N_4049);
and U7061 (N_7061,N_2906,N_459);
xnor U7062 (N_7062,N_4753,N_1082);
nand U7063 (N_7063,N_1188,N_2679);
or U7064 (N_7064,N_1945,N_4350);
or U7065 (N_7065,N_2448,N_2516);
or U7066 (N_7066,N_2312,N_1106);
or U7067 (N_7067,N_4022,N_519);
or U7068 (N_7068,N_803,N_783);
nor U7069 (N_7069,N_4358,N_4109);
nand U7070 (N_7070,N_362,N_238);
nand U7071 (N_7071,N_2525,N_1855);
xnor U7072 (N_7072,N_4704,N_2703);
or U7073 (N_7073,N_2350,N_440);
nor U7074 (N_7074,N_2646,N_4388);
nor U7075 (N_7075,N_968,N_4067);
and U7076 (N_7076,N_1951,N_1593);
and U7077 (N_7077,N_2686,N_1537);
and U7078 (N_7078,N_2284,N_1565);
and U7079 (N_7079,N_987,N_3313);
nor U7080 (N_7080,N_3391,N_1592);
and U7081 (N_7081,N_3528,N_512);
or U7082 (N_7082,N_2366,N_4246);
nand U7083 (N_7083,N_4012,N_1500);
xor U7084 (N_7084,N_2115,N_2968);
nand U7085 (N_7085,N_3575,N_1362);
nand U7086 (N_7086,N_2626,N_3966);
or U7087 (N_7087,N_3103,N_1431);
or U7088 (N_7088,N_51,N_2706);
nor U7089 (N_7089,N_4639,N_3275);
nand U7090 (N_7090,N_2095,N_1186);
or U7091 (N_7091,N_2865,N_3998);
nor U7092 (N_7092,N_949,N_832);
xnor U7093 (N_7093,N_2814,N_3390);
xor U7094 (N_7094,N_4027,N_994);
xnor U7095 (N_7095,N_2564,N_508);
nor U7096 (N_7096,N_4577,N_4265);
xnor U7097 (N_7097,N_4680,N_3397);
nand U7098 (N_7098,N_3034,N_394);
nand U7099 (N_7099,N_247,N_3266);
or U7100 (N_7100,N_1863,N_2835);
or U7101 (N_7101,N_1476,N_2867);
xnor U7102 (N_7102,N_2810,N_1012);
and U7103 (N_7103,N_103,N_372);
or U7104 (N_7104,N_4991,N_2994);
nand U7105 (N_7105,N_1678,N_1345);
or U7106 (N_7106,N_3501,N_3314);
nor U7107 (N_7107,N_1202,N_211);
nand U7108 (N_7108,N_3871,N_2806);
xor U7109 (N_7109,N_970,N_282);
nor U7110 (N_7110,N_1780,N_1214);
or U7111 (N_7111,N_3965,N_1423);
or U7112 (N_7112,N_4238,N_3611);
and U7113 (N_7113,N_2926,N_3176);
or U7114 (N_7114,N_4244,N_1858);
nand U7115 (N_7115,N_2768,N_3165);
or U7116 (N_7116,N_562,N_4336);
xor U7117 (N_7117,N_4977,N_1624);
or U7118 (N_7118,N_1564,N_1912);
nor U7119 (N_7119,N_821,N_1916);
or U7120 (N_7120,N_1142,N_1459);
nand U7121 (N_7121,N_1891,N_3488);
and U7122 (N_7122,N_3985,N_3967);
xor U7123 (N_7123,N_2260,N_815);
nand U7124 (N_7124,N_1357,N_3788);
xnor U7125 (N_7125,N_593,N_3823);
and U7126 (N_7126,N_1996,N_485);
or U7127 (N_7127,N_749,N_738);
and U7128 (N_7128,N_1753,N_406);
nand U7129 (N_7129,N_1419,N_168);
nor U7130 (N_7130,N_4451,N_4085);
nand U7131 (N_7131,N_962,N_4776);
xor U7132 (N_7132,N_1578,N_2373);
xnor U7133 (N_7133,N_2653,N_3116);
nor U7134 (N_7134,N_3222,N_2643);
nor U7135 (N_7135,N_2514,N_2107);
nor U7136 (N_7136,N_3652,N_1368);
or U7137 (N_7137,N_1185,N_2364);
xnor U7138 (N_7138,N_3190,N_515);
xor U7139 (N_7139,N_790,N_3542);
nand U7140 (N_7140,N_1243,N_2314);
xnor U7141 (N_7141,N_1729,N_3525);
nand U7142 (N_7142,N_1513,N_4242);
and U7143 (N_7143,N_3398,N_640);
xnor U7144 (N_7144,N_1979,N_1808);
or U7145 (N_7145,N_483,N_2393);
or U7146 (N_7146,N_50,N_3301);
nor U7147 (N_7147,N_2868,N_1958);
and U7148 (N_7148,N_762,N_4194);
nand U7149 (N_7149,N_3091,N_1754);
nand U7150 (N_7150,N_1759,N_2458);
xnor U7151 (N_7151,N_2146,N_658);
nor U7152 (N_7152,N_1761,N_505);
nor U7153 (N_7153,N_888,N_524);
xor U7154 (N_7154,N_4797,N_330);
nand U7155 (N_7155,N_4582,N_4425);
nand U7156 (N_7156,N_4757,N_4346);
nand U7157 (N_7157,N_1498,N_414);
nor U7158 (N_7158,N_4438,N_3404);
or U7159 (N_7159,N_1417,N_4099);
or U7160 (N_7160,N_3311,N_45);
or U7161 (N_7161,N_4143,N_413);
or U7162 (N_7162,N_4101,N_862);
xor U7163 (N_7163,N_1766,N_3179);
and U7164 (N_7164,N_4489,N_2153);
or U7165 (N_7165,N_4538,N_17);
nand U7166 (N_7166,N_4042,N_177);
and U7167 (N_7167,N_1043,N_3747);
or U7168 (N_7168,N_1020,N_3820);
nor U7169 (N_7169,N_4586,N_4254);
nor U7170 (N_7170,N_1943,N_4982);
nand U7171 (N_7171,N_771,N_4269);
xnor U7172 (N_7172,N_1587,N_737);
xor U7173 (N_7173,N_69,N_4074);
nand U7174 (N_7174,N_2955,N_4631);
nand U7175 (N_7175,N_2227,N_1850);
or U7176 (N_7176,N_1830,N_909);
and U7177 (N_7177,N_2943,N_520);
xor U7178 (N_7178,N_1257,N_4500);
nand U7179 (N_7179,N_26,N_1406);
and U7180 (N_7180,N_4841,N_3112);
xor U7181 (N_7181,N_1237,N_567);
nand U7182 (N_7182,N_1244,N_3705);
and U7183 (N_7183,N_204,N_15);
or U7184 (N_7184,N_1661,N_46);
nor U7185 (N_7185,N_3962,N_3302);
and U7186 (N_7186,N_3419,N_3921);
nand U7187 (N_7187,N_1074,N_70);
xor U7188 (N_7188,N_3634,N_4316);
nand U7189 (N_7189,N_3553,N_41);
nand U7190 (N_7190,N_2713,N_1164);
nor U7191 (N_7191,N_1773,N_3568);
nand U7192 (N_7192,N_241,N_804);
and U7193 (N_7193,N_3012,N_904);
and U7194 (N_7194,N_1041,N_4331);
nand U7195 (N_7195,N_3894,N_2179);
or U7196 (N_7196,N_1221,N_3510);
nor U7197 (N_7197,N_3392,N_2665);
nor U7198 (N_7198,N_3281,N_3376);
and U7199 (N_7199,N_2129,N_1245);
nor U7200 (N_7200,N_549,N_2167);
nand U7201 (N_7201,N_3711,N_4723);
xor U7202 (N_7202,N_4315,N_1078);
nor U7203 (N_7203,N_1408,N_1196);
nand U7204 (N_7204,N_1644,N_3585);
or U7205 (N_7205,N_415,N_4370);
and U7206 (N_7206,N_4068,N_2056);
and U7207 (N_7207,N_2861,N_1688);
nor U7208 (N_7208,N_4121,N_1884);
or U7209 (N_7209,N_1207,N_44);
or U7210 (N_7210,N_4311,N_2140);
or U7211 (N_7211,N_1794,N_3740);
nor U7212 (N_7212,N_4531,N_3779);
or U7213 (N_7213,N_3872,N_3735);
and U7214 (N_7214,N_691,N_3361);
xnor U7215 (N_7215,N_48,N_4716);
and U7216 (N_7216,N_3856,N_1819);
nor U7217 (N_7217,N_4838,N_3192);
and U7218 (N_7218,N_2225,N_2245);
and U7219 (N_7219,N_218,N_1501);
or U7220 (N_7220,N_953,N_363);
or U7221 (N_7221,N_4552,N_2930);
or U7222 (N_7222,N_4222,N_2042);
xnor U7223 (N_7223,N_3413,N_2467);
and U7224 (N_7224,N_1820,N_4981);
and U7225 (N_7225,N_3514,N_4056);
nand U7226 (N_7226,N_890,N_4020);
nor U7227 (N_7227,N_2352,N_3162);
xor U7228 (N_7228,N_3730,N_4173);
nand U7229 (N_7229,N_281,N_2481);
and U7230 (N_7230,N_2160,N_2261);
xnor U7231 (N_7231,N_3751,N_2451);
and U7232 (N_7232,N_1017,N_2614);
nand U7233 (N_7233,N_1944,N_4437);
xnor U7234 (N_7234,N_2304,N_932);
nor U7235 (N_7235,N_1702,N_420);
xor U7236 (N_7236,N_4827,N_4119);
or U7237 (N_7237,N_1516,N_2490);
or U7238 (N_7238,N_4334,N_746);
or U7239 (N_7239,N_2854,N_625);
nand U7240 (N_7240,N_859,N_4833);
and U7241 (N_7241,N_3009,N_3138);
nand U7242 (N_7242,N_2209,N_3267);
or U7243 (N_7243,N_3430,N_4788);
nand U7244 (N_7244,N_838,N_1675);
xnor U7245 (N_7245,N_2783,N_2019);
xnor U7246 (N_7246,N_4330,N_300);
nor U7247 (N_7247,N_2996,N_2369);
xnor U7248 (N_7248,N_1385,N_1725);
nor U7249 (N_7249,N_2447,N_3047);
nand U7250 (N_7250,N_2566,N_2193);
or U7251 (N_7251,N_2188,N_735);
and U7252 (N_7252,N_2275,N_3538);
nor U7253 (N_7253,N_3641,N_2437);
nand U7254 (N_7254,N_2712,N_3645);
xnor U7255 (N_7255,N_1569,N_2155);
or U7256 (N_7256,N_232,N_4540);
xnor U7257 (N_7257,N_338,N_1527);
xnor U7258 (N_7258,N_2224,N_4197);
nand U7259 (N_7259,N_1571,N_2426);
or U7260 (N_7260,N_637,N_3580);
nor U7261 (N_7261,N_2802,N_1764);
or U7262 (N_7262,N_2254,N_638);
or U7263 (N_7263,N_207,N_3325);
and U7264 (N_7264,N_1067,N_93);
or U7265 (N_7265,N_4363,N_3049);
nor U7266 (N_7266,N_4002,N_4134);
nand U7267 (N_7267,N_1428,N_4223);
nand U7268 (N_7268,N_595,N_2131);
xnor U7269 (N_7269,N_2009,N_2902);
or U7270 (N_7270,N_2693,N_3158);
and U7271 (N_7271,N_1726,N_3692);
nor U7272 (N_7272,N_2604,N_943);
or U7273 (N_7273,N_1239,N_3252);
and U7274 (N_7274,N_4936,N_3713);
xor U7275 (N_7275,N_3797,N_1375);
xor U7276 (N_7276,N_644,N_3616);
xor U7277 (N_7277,N_3996,N_2511);
or U7278 (N_7278,N_2554,N_2267);
xnor U7279 (N_7279,N_1840,N_4607);
and U7280 (N_7280,N_4395,N_4253);
or U7281 (N_7281,N_2832,N_2075);
xor U7282 (N_7282,N_1341,N_4567);
and U7283 (N_7283,N_3716,N_2217);
nand U7284 (N_7284,N_3682,N_3848);
and U7285 (N_7285,N_4612,N_1029);
and U7286 (N_7286,N_4272,N_2774);
nand U7287 (N_7287,N_4789,N_3827);
nand U7288 (N_7288,N_1961,N_3228);
xnor U7289 (N_7289,N_788,N_2157);
nand U7290 (N_7290,N_4204,N_576);
nand U7291 (N_7291,N_339,N_4319);
nand U7292 (N_7292,N_1594,N_4881);
and U7293 (N_7293,N_2308,N_1892);
nand U7294 (N_7294,N_3247,N_4408);
or U7295 (N_7295,N_1175,N_1446);
and U7296 (N_7296,N_4566,N_4127);
nand U7297 (N_7297,N_2778,N_4834);
and U7298 (N_7298,N_56,N_2051);
and U7299 (N_7299,N_3405,N_2583);
xor U7300 (N_7300,N_2739,N_2093);
or U7301 (N_7301,N_1047,N_1325);
nor U7302 (N_7302,N_3707,N_2838);
or U7303 (N_7303,N_831,N_2007);
nor U7304 (N_7304,N_4069,N_1401);
and U7305 (N_7305,N_2821,N_2970);
nand U7306 (N_7306,N_2168,N_3345);
xor U7307 (N_7307,N_2427,N_165);
or U7308 (N_7308,N_1856,N_3422);
and U7309 (N_7309,N_1901,N_1580);
xnor U7310 (N_7310,N_2558,N_4166);
xnor U7311 (N_7311,N_249,N_1664);
nor U7312 (N_7312,N_117,N_4174);
or U7313 (N_7313,N_1758,N_4650);
nand U7314 (N_7314,N_2856,N_151);
and U7315 (N_7315,N_1402,N_3030);
or U7316 (N_7316,N_3964,N_3198);
xor U7317 (N_7317,N_3777,N_580);
nor U7318 (N_7318,N_3277,N_3775);
xor U7319 (N_7319,N_886,N_584);
nor U7320 (N_7320,N_4013,N_428);
or U7321 (N_7321,N_3226,N_4585);
nand U7322 (N_7322,N_292,N_4843);
xnor U7323 (N_7323,N_52,N_3955);
xnor U7324 (N_7324,N_906,N_2085);
nand U7325 (N_7325,N_2849,N_3043);
and U7326 (N_7326,N_4986,N_61);
nor U7327 (N_7327,N_1108,N_1379);
nand U7328 (N_7328,N_3141,N_3766);
nor U7329 (N_7329,N_3374,N_1657);
and U7330 (N_7330,N_1018,N_239);
xor U7331 (N_7331,N_2622,N_2909);
nand U7332 (N_7332,N_2248,N_4061);
nand U7333 (N_7333,N_2894,N_847);
nor U7334 (N_7334,N_2797,N_3897);
xor U7335 (N_7335,N_3339,N_682);
xor U7336 (N_7336,N_553,N_3342);
nor U7337 (N_7337,N_2666,N_1632);
nand U7338 (N_7338,N_2561,N_1815);
xnor U7339 (N_7339,N_1421,N_2003);
and U7340 (N_7340,N_3146,N_610);
and U7341 (N_7341,N_1089,N_3691);
nand U7342 (N_7342,N_4795,N_157);
nand U7343 (N_7343,N_3864,N_561);
nor U7344 (N_7344,N_2084,N_3642);
and U7345 (N_7345,N_3621,N_3084);
nand U7346 (N_7346,N_3926,N_3762);
nand U7347 (N_7347,N_3035,N_677);
xor U7348 (N_7348,N_2445,N_3720);
nand U7349 (N_7349,N_1681,N_894);
or U7350 (N_7350,N_3256,N_2880);
xnor U7351 (N_7351,N_2809,N_514);
or U7352 (N_7352,N_4733,N_4672);
xor U7353 (N_7353,N_4112,N_3581);
or U7354 (N_7354,N_568,N_1532);
xnor U7355 (N_7355,N_2667,N_3421);
xnor U7356 (N_7356,N_3438,N_1492);
or U7357 (N_7357,N_3821,N_4832);
and U7358 (N_7358,N_2156,N_2907);
nand U7359 (N_7359,N_2195,N_1283);
xor U7360 (N_7360,N_2474,N_1016);
or U7361 (N_7361,N_4610,N_2556);
or U7362 (N_7362,N_1907,N_3196);
xnor U7363 (N_7363,N_3120,N_3121);
nor U7364 (N_7364,N_4656,N_2512);
or U7365 (N_7365,N_2466,N_126);
xor U7366 (N_7366,N_352,N_1461);
xor U7367 (N_7367,N_1066,N_3695);
and U7368 (N_7368,N_939,N_2781);
nor U7369 (N_7369,N_2987,N_4281);
and U7370 (N_7370,N_2840,N_4247);
xor U7371 (N_7371,N_342,N_556);
nor U7372 (N_7372,N_4309,N_4576);
xnor U7373 (N_7373,N_3768,N_4369);
or U7374 (N_7374,N_3895,N_2052);
and U7375 (N_7375,N_3255,N_4212);
and U7376 (N_7376,N_3343,N_1666);
nor U7377 (N_7377,N_321,N_3211);
nand U7378 (N_7378,N_3435,N_2169);
or U7379 (N_7379,N_3441,N_2857);
nor U7380 (N_7380,N_4921,N_4907);
or U7381 (N_7381,N_2521,N_3305);
nor U7382 (N_7382,N_400,N_3491);
nor U7383 (N_7383,N_3999,N_4996);
or U7384 (N_7384,N_4821,N_3728);
or U7385 (N_7385,N_171,N_2380);
nand U7386 (N_7386,N_2401,N_2172);
or U7387 (N_7387,N_4424,N_107);
nand U7388 (N_7388,N_3270,N_3073);
nand U7389 (N_7389,N_940,N_3031);
xnor U7390 (N_7390,N_3189,N_3573);
nor U7391 (N_7391,N_2973,N_4433);
or U7392 (N_7392,N_4097,N_1663);
nand U7393 (N_7393,N_22,N_3518);
or U7394 (N_7394,N_1011,N_4542);
nor U7395 (N_7395,N_4314,N_2226);
xor U7396 (N_7396,N_1649,N_4730);
xor U7397 (N_7397,N_4057,N_2645);
and U7398 (N_7398,N_3850,N_1913);
xor U7399 (N_7399,N_3487,N_3900);
nor U7400 (N_7400,N_2001,N_1005);
xnor U7401 (N_7401,N_4211,N_3892);
or U7402 (N_7402,N_3147,N_617);
and U7403 (N_7403,N_253,N_662);
xnor U7404 (N_7404,N_4160,N_1299);
and U7405 (N_7405,N_4747,N_234);
xor U7406 (N_7406,N_3074,N_1439);
and U7407 (N_7407,N_2014,N_4298);
and U7408 (N_7408,N_4021,N_1121);
nand U7409 (N_7409,N_294,N_4189);
nor U7410 (N_7410,N_1911,N_4385);
xnor U7411 (N_7411,N_1534,N_1393);
and U7412 (N_7412,N_3458,N_1400);
nand U7413 (N_7413,N_16,N_4200);
or U7414 (N_7414,N_3297,N_3947);
xor U7415 (N_7415,N_3426,N_3166);
and U7416 (N_7416,N_3783,N_2862);
and U7417 (N_7417,N_2382,N_3667);
and U7418 (N_7418,N_2230,N_3727);
nand U7419 (N_7419,N_1161,N_741);
xor U7420 (N_7420,N_3444,N_1757);
xnor U7421 (N_7421,N_1873,N_1291);
nand U7422 (N_7422,N_4636,N_1967);
nor U7423 (N_7423,N_3649,N_3552);
xor U7424 (N_7424,N_4671,N_447);
xnor U7425 (N_7425,N_4830,N_3804);
nand U7426 (N_7426,N_4387,N_3825);
nor U7427 (N_7427,N_3618,N_4698);
nor U7428 (N_7428,N_740,N_4638);
nor U7429 (N_7429,N_4900,N_4138);
or U7430 (N_7430,N_1480,N_1626);
nand U7431 (N_7431,N_4094,N_2743);
xnor U7432 (N_7432,N_4055,N_4354);
xnor U7433 (N_7433,N_2559,N_3715);
or U7434 (N_7434,N_1024,N_1521);
or U7435 (N_7435,N_4847,N_3326);
nand U7436 (N_7436,N_751,N_1804);
or U7437 (N_7437,N_907,N_2162);
xor U7438 (N_7438,N_206,N_2546);
and U7439 (N_7439,N_1059,N_1139);
xnor U7440 (N_7440,N_2746,N_2681);
nor U7441 (N_7441,N_1966,N_1076);
nand U7442 (N_7442,N_271,N_3105);
or U7443 (N_7443,N_129,N_4948);
nand U7444 (N_7444,N_4632,N_2808);
or U7445 (N_7445,N_2328,N_2954);
nor U7446 (N_7446,N_4679,N_1610);
nand U7447 (N_7447,N_286,N_4652);
xor U7448 (N_7448,N_3081,N_1107);
or U7449 (N_7449,N_1673,N_3337);
or U7450 (N_7450,N_2475,N_2013);
and U7451 (N_7451,N_1937,N_72);
or U7452 (N_7452,N_3638,N_3304);
nand U7453 (N_7453,N_20,N_4591);
and U7454 (N_7454,N_2545,N_4164);
xor U7455 (N_7455,N_99,N_2661);
and U7456 (N_7456,N_4278,N_220);
and U7457 (N_7457,N_2860,N_4327);
xor U7458 (N_7458,N_2258,N_1276);
or U7459 (N_7459,N_3885,N_212);
xor U7460 (N_7460,N_315,N_3429);
xor U7461 (N_7461,N_210,N_132);
and U7462 (N_7462,N_2984,N_4768);
or U7463 (N_7463,N_2343,N_4935);
nand U7464 (N_7464,N_1896,N_4911);
nand U7465 (N_7465,N_2219,N_1541);
or U7466 (N_7466,N_1463,N_3694);
or U7467 (N_7467,N_2660,N_4589);
xnor U7468 (N_7468,N_2700,N_1899);
xor U7469 (N_7469,N_1235,N_4777);
nor U7470 (N_7470,N_1809,N_3929);
nand U7471 (N_7471,N_772,N_2220);
nor U7472 (N_7472,N_1730,N_4890);
nand U7473 (N_7473,N_28,N_1485);
or U7474 (N_7474,N_491,N_2639);
xnor U7475 (N_7475,N_4583,N_2266);
and U7476 (N_7476,N_194,N_1767);
or U7477 (N_7477,N_2587,N_3665);
and U7478 (N_7478,N_18,N_277);
and U7479 (N_7479,N_4579,N_824);
nor U7480 (N_7480,N_3238,N_2250);
or U7481 (N_7481,N_3771,N_3963);
nor U7482 (N_7482,N_366,N_59);
and U7483 (N_7483,N_3143,N_4093);
nand U7484 (N_7484,N_1460,N_4441);
nand U7485 (N_7485,N_4879,N_2578);
and U7486 (N_7486,N_2509,N_3453);
nor U7487 (N_7487,N_2221,N_818);
nand U7488 (N_7488,N_3545,N_4005);
and U7489 (N_7489,N_1208,N_2664);
nor U7490 (N_7490,N_4633,N_3776);
or U7491 (N_7491,N_2163,N_83);
or U7492 (N_7492,N_517,N_1540);
nor U7493 (N_7493,N_1584,N_1948);
nand U7494 (N_7494,N_3239,N_3036);
nor U7495 (N_7495,N_246,N_3164);
or U7496 (N_7496,N_2663,N_1535);
nor U7497 (N_7497,N_3521,N_1432);
or U7498 (N_7498,N_3371,N_4555);
xor U7499 (N_7499,N_235,N_2406);
xnor U7500 (N_7500,N_3426,N_3551);
or U7501 (N_7501,N_1434,N_2936);
xnor U7502 (N_7502,N_2773,N_276);
or U7503 (N_7503,N_2328,N_2087);
xnor U7504 (N_7504,N_94,N_504);
nand U7505 (N_7505,N_1122,N_642);
nand U7506 (N_7506,N_1047,N_4177);
xor U7507 (N_7507,N_1860,N_3006);
nand U7508 (N_7508,N_868,N_89);
xor U7509 (N_7509,N_1657,N_1983);
nand U7510 (N_7510,N_638,N_2946);
nand U7511 (N_7511,N_1853,N_3174);
nand U7512 (N_7512,N_1380,N_2386);
nor U7513 (N_7513,N_706,N_1829);
nor U7514 (N_7514,N_1664,N_1558);
nor U7515 (N_7515,N_4257,N_4726);
xor U7516 (N_7516,N_288,N_4970);
nor U7517 (N_7517,N_4343,N_172);
nand U7518 (N_7518,N_2399,N_2299);
nor U7519 (N_7519,N_1577,N_4650);
xnor U7520 (N_7520,N_2145,N_200);
or U7521 (N_7521,N_3308,N_2610);
nand U7522 (N_7522,N_1464,N_32);
or U7523 (N_7523,N_4994,N_1492);
or U7524 (N_7524,N_1271,N_1665);
or U7525 (N_7525,N_3947,N_1783);
nand U7526 (N_7526,N_4087,N_1193);
and U7527 (N_7527,N_4615,N_541);
and U7528 (N_7528,N_106,N_537);
xnor U7529 (N_7529,N_1127,N_1435);
nor U7530 (N_7530,N_1111,N_4084);
or U7531 (N_7531,N_2833,N_4357);
and U7532 (N_7532,N_119,N_3006);
nand U7533 (N_7533,N_4146,N_1511);
nand U7534 (N_7534,N_1256,N_4381);
nor U7535 (N_7535,N_150,N_3081);
and U7536 (N_7536,N_1591,N_1741);
nor U7537 (N_7537,N_4493,N_4081);
and U7538 (N_7538,N_1144,N_3921);
xor U7539 (N_7539,N_1711,N_1877);
or U7540 (N_7540,N_733,N_392);
nand U7541 (N_7541,N_783,N_3290);
xnor U7542 (N_7542,N_2582,N_4655);
nor U7543 (N_7543,N_3373,N_3403);
xor U7544 (N_7544,N_541,N_4406);
nand U7545 (N_7545,N_4674,N_4828);
xnor U7546 (N_7546,N_2962,N_2611);
xnor U7547 (N_7547,N_3466,N_4142);
nor U7548 (N_7548,N_266,N_286);
nor U7549 (N_7549,N_4944,N_4836);
nor U7550 (N_7550,N_2933,N_2106);
nand U7551 (N_7551,N_386,N_1906);
nand U7552 (N_7552,N_1363,N_3935);
nand U7553 (N_7553,N_1033,N_4635);
nor U7554 (N_7554,N_2677,N_3164);
xnor U7555 (N_7555,N_1679,N_4050);
xnor U7556 (N_7556,N_4330,N_298);
and U7557 (N_7557,N_4951,N_1335);
nand U7558 (N_7558,N_4261,N_2737);
nor U7559 (N_7559,N_3222,N_4418);
nand U7560 (N_7560,N_3837,N_352);
and U7561 (N_7561,N_3755,N_117);
and U7562 (N_7562,N_4237,N_3168);
or U7563 (N_7563,N_4116,N_4168);
or U7564 (N_7564,N_3640,N_4207);
or U7565 (N_7565,N_4651,N_2029);
nor U7566 (N_7566,N_2292,N_845);
and U7567 (N_7567,N_4392,N_4959);
and U7568 (N_7568,N_2771,N_4736);
and U7569 (N_7569,N_2488,N_1647);
xnor U7570 (N_7570,N_2828,N_4502);
nor U7571 (N_7571,N_601,N_2564);
nor U7572 (N_7572,N_965,N_1622);
nor U7573 (N_7573,N_3051,N_297);
or U7574 (N_7574,N_4718,N_4091);
and U7575 (N_7575,N_2887,N_280);
nor U7576 (N_7576,N_3415,N_4945);
nand U7577 (N_7577,N_2795,N_491);
xor U7578 (N_7578,N_3277,N_896);
and U7579 (N_7579,N_2818,N_2919);
xnor U7580 (N_7580,N_4154,N_634);
nand U7581 (N_7581,N_3083,N_4045);
or U7582 (N_7582,N_1611,N_3773);
or U7583 (N_7583,N_966,N_1848);
nand U7584 (N_7584,N_3387,N_3539);
nand U7585 (N_7585,N_725,N_2435);
and U7586 (N_7586,N_4310,N_2186);
nand U7587 (N_7587,N_1452,N_4033);
or U7588 (N_7588,N_4764,N_3068);
xor U7589 (N_7589,N_537,N_912);
nand U7590 (N_7590,N_3385,N_1970);
nor U7591 (N_7591,N_3596,N_3589);
and U7592 (N_7592,N_537,N_1679);
nor U7593 (N_7593,N_448,N_217);
xnor U7594 (N_7594,N_2341,N_115);
nand U7595 (N_7595,N_1992,N_138);
xnor U7596 (N_7596,N_2855,N_2154);
nor U7597 (N_7597,N_3258,N_106);
and U7598 (N_7598,N_72,N_1380);
nand U7599 (N_7599,N_2477,N_2685);
xnor U7600 (N_7600,N_2787,N_4945);
xnor U7601 (N_7601,N_3074,N_1499);
or U7602 (N_7602,N_1153,N_1303);
xor U7603 (N_7603,N_3107,N_2532);
or U7604 (N_7604,N_2353,N_4475);
and U7605 (N_7605,N_2611,N_1842);
nand U7606 (N_7606,N_839,N_1753);
and U7607 (N_7607,N_2696,N_3839);
xnor U7608 (N_7608,N_2274,N_1140);
nor U7609 (N_7609,N_3623,N_214);
xnor U7610 (N_7610,N_1922,N_1953);
and U7611 (N_7611,N_4757,N_868);
xor U7612 (N_7612,N_2764,N_3358);
nand U7613 (N_7613,N_326,N_4175);
and U7614 (N_7614,N_655,N_4374);
and U7615 (N_7615,N_3693,N_2016);
nor U7616 (N_7616,N_4792,N_3735);
nor U7617 (N_7617,N_4143,N_3473);
nor U7618 (N_7618,N_2259,N_4772);
nor U7619 (N_7619,N_71,N_2145);
nor U7620 (N_7620,N_3981,N_106);
or U7621 (N_7621,N_3295,N_1917);
nand U7622 (N_7622,N_1481,N_2774);
nand U7623 (N_7623,N_3222,N_2353);
xnor U7624 (N_7624,N_3724,N_1156);
or U7625 (N_7625,N_2908,N_847);
or U7626 (N_7626,N_4395,N_937);
and U7627 (N_7627,N_1799,N_4205);
nand U7628 (N_7628,N_1639,N_1171);
xor U7629 (N_7629,N_3364,N_4311);
xor U7630 (N_7630,N_1147,N_794);
and U7631 (N_7631,N_4256,N_1009);
nor U7632 (N_7632,N_1893,N_4607);
nand U7633 (N_7633,N_3639,N_4809);
nand U7634 (N_7634,N_2572,N_214);
xnor U7635 (N_7635,N_1477,N_4311);
xnor U7636 (N_7636,N_1798,N_2928);
nand U7637 (N_7637,N_4126,N_1888);
xnor U7638 (N_7638,N_40,N_792);
and U7639 (N_7639,N_3479,N_905);
xor U7640 (N_7640,N_892,N_769);
and U7641 (N_7641,N_2134,N_1498);
nand U7642 (N_7642,N_3229,N_2821);
xnor U7643 (N_7643,N_420,N_3263);
nand U7644 (N_7644,N_1539,N_499);
nand U7645 (N_7645,N_760,N_39);
nor U7646 (N_7646,N_721,N_1449);
or U7647 (N_7647,N_780,N_3330);
nand U7648 (N_7648,N_2827,N_3175);
nor U7649 (N_7649,N_3425,N_128);
and U7650 (N_7650,N_4803,N_1622);
or U7651 (N_7651,N_2469,N_4092);
or U7652 (N_7652,N_1761,N_4811);
nor U7653 (N_7653,N_4508,N_3719);
nand U7654 (N_7654,N_3895,N_3904);
and U7655 (N_7655,N_2990,N_127);
or U7656 (N_7656,N_757,N_916);
nor U7657 (N_7657,N_814,N_713);
nor U7658 (N_7658,N_506,N_1765);
nor U7659 (N_7659,N_3926,N_888);
or U7660 (N_7660,N_1780,N_4946);
or U7661 (N_7661,N_1351,N_3913);
or U7662 (N_7662,N_4981,N_4588);
nand U7663 (N_7663,N_1239,N_585);
nor U7664 (N_7664,N_2677,N_581);
and U7665 (N_7665,N_1396,N_138);
nand U7666 (N_7666,N_3573,N_2278);
xnor U7667 (N_7667,N_2021,N_3208);
and U7668 (N_7668,N_2149,N_3683);
or U7669 (N_7669,N_2924,N_1394);
nand U7670 (N_7670,N_1654,N_313);
xor U7671 (N_7671,N_321,N_1687);
nand U7672 (N_7672,N_4910,N_4103);
or U7673 (N_7673,N_4943,N_4855);
or U7674 (N_7674,N_4767,N_1337);
and U7675 (N_7675,N_251,N_4173);
nor U7676 (N_7676,N_2739,N_2995);
and U7677 (N_7677,N_2022,N_1399);
and U7678 (N_7678,N_373,N_1694);
xor U7679 (N_7679,N_4096,N_4207);
or U7680 (N_7680,N_2274,N_348);
or U7681 (N_7681,N_1599,N_1765);
xnor U7682 (N_7682,N_998,N_4491);
or U7683 (N_7683,N_361,N_918);
nor U7684 (N_7684,N_819,N_718);
xor U7685 (N_7685,N_411,N_4896);
or U7686 (N_7686,N_1339,N_2597);
xor U7687 (N_7687,N_4408,N_2949);
xor U7688 (N_7688,N_4247,N_4302);
xnor U7689 (N_7689,N_1128,N_800);
nor U7690 (N_7690,N_609,N_1025);
xor U7691 (N_7691,N_4280,N_520);
or U7692 (N_7692,N_2885,N_2400);
and U7693 (N_7693,N_737,N_2415);
or U7694 (N_7694,N_2987,N_3267);
or U7695 (N_7695,N_3611,N_3754);
nor U7696 (N_7696,N_3827,N_3530);
nand U7697 (N_7697,N_3747,N_52);
nand U7698 (N_7698,N_1833,N_1122);
and U7699 (N_7699,N_390,N_4954);
xor U7700 (N_7700,N_233,N_2021);
nor U7701 (N_7701,N_4683,N_1596);
nor U7702 (N_7702,N_4926,N_1548);
and U7703 (N_7703,N_999,N_2476);
nor U7704 (N_7704,N_1342,N_471);
nand U7705 (N_7705,N_4330,N_995);
or U7706 (N_7706,N_585,N_1562);
or U7707 (N_7707,N_1505,N_2158);
nand U7708 (N_7708,N_281,N_1957);
and U7709 (N_7709,N_2690,N_786);
nand U7710 (N_7710,N_3539,N_4540);
xor U7711 (N_7711,N_4755,N_2409);
and U7712 (N_7712,N_1387,N_1718);
nor U7713 (N_7713,N_2779,N_725);
nand U7714 (N_7714,N_1610,N_1728);
or U7715 (N_7715,N_4494,N_1357);
or U7716 (N_7716,N_2975,N_2807);
and U7717 (N_7717,N_1881,N_1937);
nor U7718 (N_7718,N_290,N_2301);
nand U7719 (N_7719,N_1981,N_1914);
nand U7720 (N_7720,N_4153,N_3242);
or U7721 (N_7721,N_3568,N_2147);
nand U7722 (N_7722,N_771,N_2920);
or U7723 (N_7723,N_554,N_4450);
nor U7724 (N_7724,N_207,N_4556);
xor U7725 (N_7725,N_3617,N_3278);
nand U7726 (N_7726,N_4657,N_203);
nand U7727 (N_7727,N_4600,N_1033);
xor U7728 (N_7728,N_1970,N_3308);
or U7729 (N_7729,N_3710,N_3823);
or U7730 (N_7730,N_1605,N_1764);
xnor U7731 (N_7731,N_4649,N_1502);
xnor U7732 (N_7732,N_896,N_4891);
xnor U7733 (N_7733,N_3690,N_416);
and U7734 (N_7734,N_4069,N_1795);
nor U7735 (N_7735,N_112,N_2782);
or U7736 (N_7736,N_4324,N_746);
or U7737 (N_7737,N_1014,N_3038);
xor U7738 (N_7738,N_1051,N_1592);
nand U7739 (N_7739,N_1637,N_4816);
or U7740 (N_7740,N_3236,N_4211);
nand U7741 (N_7741,N_852,N_2131);
nand U7742 (N_7742,N_2553,N_460);
nand U7743 (N_7743,N_1589,N_3202);
xor U7744 (N_7744,N_3718,N_2706);
and U7745 (N_7745,N_2563,N_3966);
nor U7746 (N_7746,N_4459,N_517);
xnor U7747 (N_7747,N_2613,N_269);
nand U7748 (N_7748,N_1480,N_2978);
nor U7749 (N_7749,N_1137,N_1183);
nor U7750 (N_7750,N_1435,N_3501);
nand U7751 (N_7751,N_2308,N_3136);
nand U7752 (N_7752,N_3743,N_1474);
xnor U7753 (N_7753,N_1409,N_2589);
xor U7754 (N_7754,N_4878,N_4954);
nand U7755 (N_7755,N_3481,N_2976);
and U7756 (N_7756,N_3687,N_2739);
or U7757 (N_7757,N_2435,N_3706);
xnor U7758 (N_7758,N_1234,N_4796);
and U7759 (N_7759,N_3073,N_1225);
or U7760 (N_7760,N_3979,N_2763);
xnor U7761 (N_7761,N_3633,N_1972);
and U7762 (N_7762,N_1275,N_1554);
and U7763 (N_7763,N_3725,N_3187);
or U7764 (N_7764,N_1918,N_2952);
nor U7765 (N_7765,N_2942,N_2867);
nor U7766 (N_7766,N_1817,N_723);
xnor U7767 (N_7767,N_2891,N_2712);
or U7768 (N_7768,N_4012,N_3728);
and U7769 (N_7769,N_4100,N_617);
xor U7770 (N_7770,N_2124,N_1539);
nand U7771 (N_7771,N_3114,N_710);
and U7772 (N_7772,N_3739,N_4654);
nor U7773 (N_7773,N_2595,N_100);
xnor U7774 (N_7774,N_3390,N_2949);
xor U7775 (N_7775,N_3328,N_1498);
nand U7776 (N_7776,N_1124,N_4174);
nand U7777 (N_7777,N_4413,N_4735);
or U7778 (N_7778,N_3897,N_748);
and U7779 (N_7779,N_3252,N_315);
xor U7780 (N_7780,N_3882,N_4305);
nor U7781 (N_7781,N_40,N_1001);
or U7782 (N_7782,N_851,N_1826);
nand U7783 (N_7783,N_2146,N_3926);
nand U7784 (N_7784,N_4151,N_4777);
and U7785 (N_7785,N_2384,N_3849);
or U7786 (N_7786,N_1865,N_1358);
nand U7787 (N_7787,N_3051,N_685);
or U7788 (N_7788,N_1463,N_4285);
nand U7789 (N_7789,N_2168,N_3624);
and U7790 (N_7790,N_3529,N_4042);
and U7791 (N_7791,N_3160,N_1976);
nor U7792 (N_7792,N_4714,N_1525);
xnor U7793 (N_7793,N_4577,N_4817);
nor U7794 (N_7794,N_1996,N_2463);
nand U7795 (N_7795,N_1347,N_501);
nor U7796 (N_7796,N_1603,N_277);
nor U7797 (N_7797,N_179,N_1034);
nand U7798 (N_7798,N_2193,N_4085);
or U7799 (N_7799,N_2200,N_4992);
and U7800 (N_7800,N_3473,N_1063);
or U7801 (N_7801,N_2060,N_529);
xnor U7802 (N_7802,N_4751,N_3908);
nor U7803 (N_7803,N_2260,N_1488);
nor U7804 (N_7804,N_469,N_1955);
or U7805 (N_7805,N_4449,N_1171);
nand U7806 (N_7806,N_2648,N_4505);
and U7807 (N_7807,N_4302,N_135);
nor U7808 (N_7808,N_3193,N_3337);
nor U7809 (N_7809,N_2809,N_4304);
nor U7810 (N_7810,N_3742,N_4436);
or U7811 (N_7811,N_111,N_932);
xnor U7812 (N_7812,N_1376,N_300);
nor U7813 (N_7813,N_2173,N_170);
nor U7814 (N_7814,N_1156,N_465);
or U7815 (N_7815,N_156,N_865);
xor U7816 (N_7816,N_3519,N_2070);
and U7817 (N_7817,N_3070,N_3525);
xnor U7818 (N_7818,N_3091,N_1372);
nand U7819 (N_7819,N_1772,N_574);
nor U7820 (N_7820,N_1474,N_1362);
and U7821 (N_7821,N_3139,N_652);
xor U7822 (N_7822,N_603,N_450);
nand U7823 (N_7823,N_1966,N_82);
nor U7824 (N_7824,N_988,N_4724);
and U7825 (N_7825,N_1052,N_3673);
xor U7826 (N_7826,N_626,N_3209);
nand U7827 (N_7827,N_215,N_4749);
xor U7828 (N_7828,N_1932,N_949);
xnor U7829 (N_7829,N_4417,N_1832);
or U7830 (N_7830,N_3990,N_727);
and U7831 (N_7831,N_1396,N_3621);
and U7832 (N_7832,N_4176,N_4316);
nor U7833 (N_7833,N_3393,N_374);
nor U7834 (N_7834,N_4570,N_4441);
nor U7835 (N_7835,N_800,N_4051);
nand U7836 (N_7836,N_2947,N_993);
xnor U7837 (N_7837,N_192,N_2809);
or U7838 (N_7838,N_4786,N_574);
nor U7839 (N_7839,N_348,N_340);
nand U7840 (N_7840,N_2850,N_3645);
nor U7841 (N_7841,N_573,N_2143);
or U7842 (N_7842,N_673,N_632);
nor U7843 (N_7843,N_1889,N_1576);
nand U7844 (N_7844,N_1214,N_1425);
or U7845 (N_7845,N_324,N_490);
xnor U7846 (N_7846,N_1853,N_359);
or U7847 (N_7847,N_4811,N_409);
nand U7848 (N_7848,N_1697,N_942);
and U7849 (N_7849,N_2556,N_2106);
nand U7850 (N_7850,N_2183,N_3800);
xnor U7851 (N_7851,N_191,N_2810);
or U7852 (N_7852,N_2195,N_1030);
nand U7853 (N_7853,N_4352,N_2641);
or U7854 (N_7854,N_2870,N_1104);
nand U7855 (N_7855,N_4980,N_3047);
nand U7856 (N_7856,N_327,N_1003);
nor U7857 (N_7857,N_4032,N_3709);
nor U7858 (N_7858,N_464,N_2341);
and U7859 (N_7859,N_1028,N_4478);
and U7860 (N_7860,N_7,N_4237);
and U7861 (N_7861,N_557,N_3556);
xnor U7862 (N_7862,N_4320,N_3947);
nand U7863 (N_7863,N_3187,N_218);
xor U7864 (N_7864,N_1496,N_1136);
nand U7865 (N_7865,N_1076,N_3905);
xnor U7866 (N_7866,N_3724,N_1388);
nand U7867 (N_7867,N_1879,N_4255);
nand U7868 (N_7868,N_1783,N_4474);
or U7869 (N_7869,N_4235,N_1245);
and U7870 (N_7870,N_1989,N_2534);
and U7871 (N_7871,N_3922,N_2435);
and U7872 (N_7872,N_1601,N_4167);
or U7873 (N_7873,N_710,N_1296);
nand U7874 (N_7874,N_3611,N_2833);
xor U7875 (N_7875,N_4042,N_3549);
nand U7876 (N_7876,N_4886,N_4352);
and U7877 (N_7877,N_2973,N_1122);
and U7878 (N_7878,N_4511,N_390);
xnor U7879 (N_7879,N_4347,N_1518);
nand U7880 (N_7880,N_1473,N_2240);
xnor U7881 (N_7881,N_533,N_1357);
xnor U7882 (N_7882,N_3874,N_4929);
nor U7883 (N_7883,N_2420,N_4690);
or U7884 (N_7884,N_2109,N_2736);
and U7885 (N_7885,N_1967,N_3660);
nor U7886 (N_7886,N_1691,N_1391);
and U7887 (N_7887,N_3499,N_2669);
xor U7888 (N_7888,N_2581,N_1886);
nand U7889 (N_7889,N_3637,N_3156);
nand U7890 (N_7890,N_167,N_993);
and U7891 (N_7891,N_3977,N_907);
nand U7892 (N_7892,N_1967,N_3082);
nand U7893 (N_7893,N_103,N_2581);
nor U7894 (N_7894,N_125,N_2682);
nor U7895 (N_7895,N_4422,N_615);
and U7896 (N_7896,N_1496,N_937);
or U7897 (N_7897,N_511,N_4692);
nand U7898 (N_7898,N_285,N_765);
xnor U7899 (N_7899,N_302,N_1210);
and U7900 (N_7900,N_2598,N_2043);
and U7901 (N_7901,N_4780,N_3765);
or U7902 (N_7902,N_3603,N_1229);
xnor U7903 (N_7903,N_134,N_4415);
xnor U7904 (N_7904,N_444,N_1768);
nor U7905 (N_7905,N_2631,N_4469);
and U7906 (N_7906,N_62,N_1131);
or U7907 (N_7907,N_551,N_4273);
nand U7908 (N_7908,N_323,N_4210);
xor U7909 (N_7909,N_4525,N_1915);
xor U7910 (N_7910,N_747,N_2022);
nor U7911 (N_7911,N_1116,N_2522);
or U7912 (N_7912,N_4064,N_2610);
or U7913 (N_7913,N_3682,N_2660);
xnor U7914 (N_7914,N_1972,N_3912);
and U7915 (N_7915,N_3378,N_2226);
nand U7916 (N_7916,N_574,N_1264);
xor U7917 (N_7917,N_2745,N_3769);
and U7918 (N_7918,N_1271,N_600);
nand U7919 (N_7919,N_4930,N_4897);
xor U7920 (N_7920,N_4546,N_3683);
or U7921 (N_7921,N_848,N_343);
or U7922 (N_7922,N_472,N_765);
nand U7923 (N_7923,N_4184,N_4811);
or U7924 (N_7924,N_2727,N_3076);
nand U7925 (N_7925,N_1333,N_2985);
or U7926 (N_7926,N_692,N_4237);
nand U7927 (N_7927,N_2839,N_4118);
nor U7928 (N_7928,N_1178,N_2516);
and U7929 (N_7929,N_3444,N_563);
nor U7930 (N_7930,N_3713,N_4436);
and U7931 (N_7931,N_835,N_2314);
or U7932 (N_7932,N_4165,N_197);
or U7933 (N_7933,N_3565,N_4143);
nor U7934 (N_7934,N_1028,N_2604);
nand U7935 (N_7935,N_2051,N_4935);
xor U7936 (N_7936,N_4170,N_3525);
nand U7937 (N_7937,N_132,N_3322);
nor U7938 (N_7938,N_4203,N_2837);
or U7939 (N_7939,N_2399,N_3871);
nand U7940 (N_7940,N_338,N_989);
nor U7941 (N_7941,N_493,N_2444);
and U7942 (N_7942,N_4858,N_4874);
or U7943 (N_7943,N_2558,N_211);
and U7944 (N_7944,N_3015,N_2638);
nor U7945 (N_7945,N_1846,N_4752);
or U7946 (N_7946,N_2229,N_430);
and U7947 (N_7947,N_1782,N_1997);
xor U7948 (N_7948,N_3946,N_4874);
nor U7949 (N_7949,N_193,N_4431);
and U7950 (N_7950,N_1030,N_3564);
nand U7951 (N_7951,N_3950,N_1256);
and U7952 (N_7952,N_3269,N_1549);
or U7953 (N_7953,N_4168,N_3927);
nor U7954 (N_7954,N_3943,N_2177);
nor U7955 (N_7955,N_1449,N_1184);
xnor U7956 (N_7956,N_2910,N_4567);
and U7957 (N_7957,N_3245,N_3822);
nand U7958 (N_7958,N_1562,N_4018);
or U7959 (N_7959,N_3643,N_4689);
and U7960 (N_7960,N_491,N_4411);
nand U7961 (N_7961,N_264,N_1246);
nand U7962 (N_7962,N_3909,N_4409);
or U7963 (N_7963,N_2074,N_2811);
or U7964 (N_7964,N_3044,N_3359);
or U7965 (N_7965,N_1564,N_2319);
nand U7966 (N_7966,N_243,N_2387);
and U7967 (N_7967,N_335,N_3644);
nor U7968 (N_7968,N_498,N_1795);
and U7969 (N_7969,N_3595,N_3304);
or U7970 (N_7970,N_303,N_2234);
xnor U7971 (N_7971,N_611,N_1596);
nor U7972 (N_7972,N_1269,N_3816);
or U7973 (N_7973,N_3603,N_1930);
or U7974 (N_7974,N_4905,N_921);
nor U7975 (N_7975,N_3488,N_4822);
nand U7976 (N_7976,N_459,N_4876);
nor U7977 (N_7977,N_557,N_2841);
and U7978 (N_7978,N_4417,N_1935);
or U7979 (N_7979,N_2000,N_1519);
nand U7980 (N_7980,N_4354,N_1741);
xnor U7981 (N_7981,N_2616,N_2416);
nand U7982 (N_7982,N_4459,N_1627);
nor U7983 (N_7983,N_1600,N_3388);
nand U7984 (N_7984,N_2324,N_305);
and U7985 (N_7985,N_932,N_2610);
and U7986 (N_7986,N_3855,N_4417);
nand U7987 (N_7987,N_3807,N_4530);
xor U7988 (N_7988,N_2713,N_2949);
nor U7989 (N_7989,N_893,N_235);
nor U7990 (N_7990,N_2,N_1752);
or U7991 (N_7991,N_2026,N_4628);
nor U7992 (N_7992,N_3652,N_1050);
and U7993 (N_7993,N_144,N_4109);
xor U7994 (N_7994,N_2522,N_592);
xor U7995 (N_7995,N_3504,N_867);
nand U7996 (N_7996,N_2515,N_2124);
xor U7997 (N_7997,N_754,N_1417);
xor U7998 (N_7998,N_2731,N_1149);
xor U7999 (N_7999,N_1266,N_2417);
xor U8000 (N_8000,N_1550,N_4942);
and U8001 (N_8001,N_3255,N_2568);
nand U8002 (N_8002,N_1057,N_2142);
xnor U8003 (N_8003,N_682,N_3843);
nand U8004 (N_8004,N_612,N_1900);
nand U8005 (N_8005,N_4098,N_4225);
or U8006 (N_8006,N_4241,N_2466);
nor U8007 (N_8007,N_3572,N_3142);
and U8008 (N_8008,N_4532,N_4508);
xor U8009 (N_8009,N_1114,N_2566);
nand U8010 (N_8010,N_3372,N_9);
nor U8011 (N_8011,N_2905,N_3978);
nor U8012 (N_8012,N_3463,N_3302);
nor U8013 (N_8013,N_1024,N_4630);
nor U8014 (N_8014,N_1299,N_530);
or U8015 (N_8015,N_2415,N_2345);
nor U8016 (N_8016,N_1627,N_4429);
or U8017 (N_8017,N_4714,N_529);
or U8018 (N_8018,N_3490,N_1873);
and U8019 (N_8019,N_1857,N_4702);
or U8020 (N_8020,N_2544,N_1887);
nor U8021 (N_8021,N_2610,N_2334);
nor U8022 (N_8022,N_1662,N_3717);
or U8023 (N_8023,N_2889,N_720);
and U8024 (N_8024,N_1278,N_3743);
xor U8025 (N_8025,N_1787,N_208);
nand U8026 (N_8026,N_4011,N_2319);
and U8027 (N_8027,N_4996,N_188);
and U8028 (N_8028,N_1565,N_2156);
and U8029 (N_8029,N_4918,N_4531);
nand U8030 (N_8030,N_1896,N_1015);
nor U8031 (N_8031,N_15,N_3805);
xnor U8032 (N_8032,N_1025,N_3672);
and U8033 (N_8033,N_4665,N_2184);
nor U8034 (N_8034,N_2874,N_1772);
nor U8035 (N_8035,N_696,N_3427);
nand U8036 (N_8036,N_483,N_1734);
nor U8037 (N_8037,N_4342,N_3610);
or U8038 (N_8038,N_19,N_2196);
or U8039 (N_8039,N_1780,N_2536);
or U8040 (N_8040,N_1228,N_110);
or U8041 (N_8041,N_3588,N_1255);
and U8042 (N_8042,N_2972,N_2271);
nor U8043 (N_8043,N_1892,N_3173);
xor U8044 (N_8044,N_3238,N_4714);
xnor U8045 (N_8045,N_465,N_2765);
xnor U8046 (N_8046,N_1643,N_1936);
or U8047 (N_8047,N_147,N_3513);
or U8048 (N_8048,N_670,N_2455);
nand U8049 (N_8049,N_1062,N_1460);
and U8050 (N_8050,N_3088,N_4237);
and U8051 (N_8051,N_4757,N_197);
and U8052 (N_8052,N_4070,N_1143);
or U8053 (N_8053,N_4399,N_2378);
nor U8054 (N_8054,N_1330,N_4732);
or U8055 (N_8055,N_4947,N_756);
nand U8056 (N_8056,N_287,N_1418);
xnor U8057 (N_8057,N_1498,N_3400);
nand U8058 (N_8058,N_1107,N_3539);
nand U8059 (N_8059,N_4379,N_452);
nor U8060 (N_8060,N_992,N_3532);
and U8061 (N_8061,N_4046,N_3845);
or U8062 (N_8062,N_525,N_4533);
and U8063 (N_8063,N_3570,N_1863);
or U8064 (N_8064,N_2066,N_505);
nand U8065 (N_8065,N_4587,N_2156);
xnor U8066 (N_8066,N_181,N_2989);
nand U8067 (N_8067,N_2290,N_4751);
xnor U8068 (N_8068,N_4705,N_4880);
and U8069 (N_8069,N_4803,N_424);
or U8070 (N_8070,N_4754,N_2901);
and U8071 (N_8071,N_4760,N_4180);
nor U8072 (N_8072,N_4422,N_4216);
nand U8073 (N_8073,N_4714,N_3096);
nand U8074 (N_8074,N_3913,N_2832);
and U8075 (N_8075,N_1924,N_4918);
nand U8076 (N_8076,N_2470,N_1227);
xor U8077 (N_8077,N_1266,N_3757);
nand U8078 (N_8078,N_2231,N_4358);
xor U8079 (N_8079,N_3305,N_1510);
or U8080 (N_8080,N_458,N_1213);
xor U8081 (N_8081,N_3009,N_2797);
nand U8082 (N_8082,N_2611,N_1997);
xnor U8083 (N_8083,N_4185,N_3903);
and U8084 (N_8084,N_3284,N_2929);
or U8085 (N_8085,N_229,N_2190);
or U8086 (N_8086,N_2834,N_411);
xor U8087 (N_8087,N_4437,N_4044);
xnor U8088 (N_8088,N_1433,N_4238);
and U8089 (N_8089,N_1940,N_2086);
or U8090 (N_8090,N_289,N_2302);
nor U8091 (N_8091,N_1787,N_3247);
nand U8092 (N_8092,N_2587,N_1449);
xnor U8093 (N_8093,N_4339,N_3839);
or U8094 (N_8094,N_4420,N_655);
and U8095 (N_8095,N_2772,N_3158);
nor U8096 (N_8096,N_2951,N_2825);
and U8097 (N_8097,N_4291,N_3989);
nor U8098 (N_8098,N_40,N_1624);
xnor U8099 (N_8099,N_1463,N_1956);
and U8100 (N_8100,N_643,N_1995);
and U8101 (N_8101,N_2581,N_162);
or U8102 (N_8102,N_2589,N_4029);
and U8103 (N_8103,N_547,N_2238);
nor U8104 (N_8104,N_967,N_2137);
nor U8105 (N_8105,N_1876,N_3961);
and U8106 (N_8106,N_203,N_4279);
nor U8107 (N_8107,N_3632,N_4458);
nand U8108 (N_8108,N_4780,N_1052);
nand U8109 (N_8109,N_2839,N_1780);
and U8110 (N_8110,N_3677,N_945);
and U8111 (N_8111,N_830,N_2427);
and U8112 (N_8112,N_3418,N_4987);
and U8113 (N_8113,N_4860,N_1158);
nor U8114 (N_8114,N_3569,N_1661);
and U8115 (N_8115,N_3746,N_3223);
xnor U8116 (N_8116,N_1719,N_3969);
nand U8117 (N_8117,N_2058,N_2253);
nand U8118 (N_8118,N_3378,N_369);
or U8119 (N_8119,N_3622,N_597);
xnor U8120 (N_8120,N_4732,N_309);
nor U8121 (N_8121,N_3067,N_1008);
nand U8122 (N_8122,N_940,N_3441);
and U8123 (N_8123,N_2703,N_2662);
or U8124 (N_8124,N_4077,N_835);
or U8125 (N_8125,N_3088,N_3286);
and U8126 (N_8126,N_1720,N_391);
nand U8127 (N_8127,N_4064,N_399);
nand U8128 (N_8128,N_2135,N_2225);
or U8129 (N_8129,N_1514,N_1241);
xnor U8130 (N_8130,N_3063,N_2967);
and U8131 (N_8131,N_4686,N_926);
nor U8132 (N_8132,N_3840,N_276);
and U8133 (N_8133,N_670,N_637);
or U8134 (N_8134,N_4954,N_1446);
nor U8135 (N_8135,N_110,N_1083);
or U8136 (N_8136,N_1053,N_4432);
xnor U8137 (N_8137,N_4669,N_3317);
nor U8138 (N_8138,N_4340,N_323);
and U8139 (N_8139,N_1981,N_1851);
and U8140 (N_8140,N_2207,N_770);
or U8141 (N_8141,N_4322,N_2507);
nor U8142 (N_8142,N_664,N_2029);
nor U8143 (N_8143,N_2837,N_1069);
nand U8144 (N_8144,N_26,N_1321);
nand U8145 (N_8145,N_4231,N_4527);
xnor U8146 (N_8146,N_1095,N_4042);
or U8147 (N_8147,N_1747,N_372);
and U8148 (N_8148,N_1596,N_4029);
nand U8149 (N_8149,N_1576,N_1007);
nor U8150 (N_8150,N_7,N_2217);
nand U8151 (N_8151,N_250,N_3364);
or U8152 (N_8152,N_59,N_1809);
or U8153 (N_8153,N_3546,N_4148);
or U8154 (N_8154,N_405,N_76);
nor U8155 (N_8155,N_2144,N_3644);
xnor U8156 (N_8156,N_2627,N_3870);
xor U8157 (N_8157,N_2267,N_365);
nand U8158 (N_8158,N_2308,N_2309);
nor U8159 (N_8159,N_1810,N_2610);
and U8160 (N_8160,N_3452,N_2559);
or U8161 (N_8161,N_3286,N_4919);
or U8162 (N_8162,N_3470,N_49);
nor U8163 (N_8163,N_3818,N_1542);
and U8164 (N_8164,N_1688,N_4393);
nor U8165 (N_8165,N_4850,N_1650);
nor U8166 (N_8166,N_2470,N_4472);
nand U8167 (N_8167,N_2470,N_4604);
nor U8168 (N_8168,N_2222,N_3973);
xnor U8169 (N_8169,N_4300,N_4996);
and U8170 (N_8170,N_1716,N_3391);
nor U8171 (N_8171,N_1323,N_1696);
nor U8172 (N_8172,N_4528,N_2420);
and U8173 (N_8173,N_2087,N_178);
xnor U8174 (N_8174,N_2354,N_1524);
nor U8175 (N_8175,N_2138,N_3128);
nor U8176 (N_8176,N_136,N_2239);
xnor U8177 (N_8177,N_772,N_3555);
or U8178 (N_8178,N_4909,N_2362);
or U8179 (N_8179,N_3433,N_2826);
or U8180 (N_8180,N_1206,N_3393);
nand U8181 (N_8181,N_2613,N_1681);
and U8182 (N_8182,N_2493,N_1270);
nor U8183 (N_8183,N_2661,N_4730);
xnor U8184 (N_8184,N_1076,N_1659);
nand U8185 (N_8185,N_3514,N_2728);
nand U8186 (N_8186,N_1809,N_1978);
xor U8187 (N_8187,N_4114,N_4260);
xor U8188 (N_8188,N_3585,N_585);
nand U8189 (N_8189,N_3345,N_2205);
or U8190 (N_8190,N_2205,N_4338);
nand U8191 (N_8191,N_4911,N_3245);
nand U8192 (N_8192,N_3448,N_666);
and U8193 (N_8193,N_2247,N_2948);
nand U8194 (N_8194,N_635,N_963);
or U8195 (N_8195,N_4071,N_211);
xnor U8196 (N_8196,N_3250,N_2475);
nor U8197 (N_8197,N_1167,N_2575);
xnor U8198 (N_8198,N_4836,N_3021);
nand U8199 (N_8199,N_4451,N_595);
nand U8200 (N_8200,N_2794,N_652);
xnor U8201 (N_8201,N_1913,N_808);
and U8202 (N_8202,N_2685,N_586);
nor U8203 (N_8203,N_4646,N_2250);
nand U8204 (N_8204,N_1859,N_1831);
or U8205 (N_8205,N_2050,N_4162);
and U8206 (N_8206,N_1932,N_485);
nor U8207 (N_8207,N_809,N_4975);
nor U8208 (N_8208,N_3284,N_2573);
xor U8209 (N_8209,N_4094,N_538);
nor U8210 (N_8210,N_3012,N_664);
nor U8211 (N_8211,N_278,N_2818);
nor U8212 (N_8212,N_3845,N_819);
or U8213 (N_8213,N_4690,N_3918);
or U8214 (N_8214,N_4876,N_4984);
xnor U8215 (N_8215,N_1529,N_3667);
nor U8216 (N_8216,N_4042,N_3265);
and U8217 (N_8217,N_4168,N_2083);
and U8218 (N_8218,N_2191,N_1659);
xnor U8219 (N_8219,N_792,N_2540);
and U8220 (N_8220,N_54,N_4892);
nor U8221 (N_8221,N_4185,N_945);
nor U8222 (N_8222,N_3558,N_3913);
or U8223 (N_8223,N_176,N_11);
or U8224 (N_8224,N_1825,N_4662);
xnor U8225 (N_8225,N_1726,N_1978);
xnor U8226 (N_8226,N_4052,N_4225);
nor U8227 (N_8227,N_4539,N_1534);
and U8228 (N_8228,N_1553,N_3831);
nand U8229 (N_8229,N_3407,N_857);
xor U8230 (N_8230,N_870,N_4448);
nand U8231 (N_8231,N_4648,N_3283);
and U8232 (N_8232,N_2647,N_2418);
or U8233 (N_8233,N_4074,N_1135);
and U8234 (N_8234,N_438,N_2539);
xnor U8235 (N_8235,N_4874,N_1025);
nand U8236 (N_8236,N_4767,N_1348);
xor U8237 (N_8237,N_2976,N_30);
or U8238 (N_8238,N_3391,N_4692);
or U8239 (N_8239,N_1282,N_3725);
and U8240 (N_8240,N_2339,N_4691);
or U8241 (N_8241,N_3680,N_1610);
or U8242 (N_8242,N_4284,N_4874);
and U8243 (N_8243,N_4294,N_2728);
nand U8244 (N_8244,N_3062,N_4784);
and U8245 (N_8245,N_4924,N_2337);
nor U8246 (N_8246,N_121,N_130);
nand U8247 (N_8247,N_1124,N_4420);
or U8248 (N_8248,N_2334,N_2190);
and U8249 (N_8249,N_1352,N_1773);
nand U8250 (N_8250,N_4336,N_4020);
and U8251 (N_8251,N_2111,N_4436);
and U8252 (N_8252,N_531,N_770);
nor U8253 (N_8253,N_4257,N_128);
and U8254 (N_8254,N_3213,N_2800);
or U8255 (N_8255,N_1832,N_142);
nand U8256 (N_8256,N_1080,N_1854);
nand U8257 (N_8257,N_4552,N_4938);
nor U8258 (N_8258,N_2699,N_3304);
and U8259 (N_8259,N_2076,N_4230);
xnor U8260 (N_8260,N_3475,N_2658);
or U8261 (N_8261,N_3901,N_4692);
or U8262 (N_8262,N_4606,N_2565);
xor U8263 (N_8263,N_4915,N_3558);
nand U8264 (N_8264,N_320,N_2470);
and U8265 (N_8265,N_3432,N_587);
nor U8266 (N_8266,N_177,N_4043);
nand U8267 (N_8267,N_759,N_1012);
nand U8268 (N_8268,N_3735,N_1318);
and U8269 (N_8269,N_447,N_422);
nor U8270 (N_8270,N_4965,N_2355);
or U8271 (N_8271,N_807,N_1137);
nand U8272 (N_8272,N_169,N_66);
nand U8273 (N_8273,N_2400,N_3943);
and U8274 (N_8274,N_1116,N_3940);
nand U8275 (N_8275,N_3267,N_3322);
xnor U8276 (N_8276,N_3573,N_2390);
nor U8277 (N_8277,N_1770,N_3684);
xor U8278 (N_8278,N_711,N_272);
and U8279 (N_8279,N_4358,N_1213);
or U8280 (N_8280,N_448,N_4468);
nand U8281 (N_8281,N_1310,N_4722);
nand U8282 (N_8282,N_3115,N_969);
or U8283 (N_8283,N_4374,N_3618);
and U8284 (N_8284,N_372,N_3499);
or U8285 (N_8285,N_878,N_3740);
nand U8286 (N_8286,N_3139,N_3949);
nor U8287 (N_8287,N_3391,N_4978);
xor U8288 (N_8288,N_4418,N_96);
or U8289 (N_8289,N_3638,N_2155);
and U8290 (N_8290,N_2805,N_3165);
or U8291 (N_8291,N_2254,N_1996);
and U8292 (N_8292,N_2286,N_1600);
nor U8293 (N_8293,N_1899,N_3172);
xnor U8294 (N_8294,N_429,N_266);
and U8295 (N_8295,N_4848,N_4466);
nand U8296 (N_8296,N_219,N_3948);
or U8297 (N_8297,N_2446,N_4113);
nor U8298 (N_8298,N_2750,N_3009);
and U8299 (N_8299,N_3331,N_1899);
nand U8300 (N_8300,N_531,N_4649);
nand U8301 (N_8301,N_3270,N_2052);
or U8302 (N_8302,N_3530,N_1084);
xor U8303 (N_8303,N_3543,N_1935);
and U8304 (N_8304,N_421,N_1960);
nand U8305 (N_8305,N_3397,N_4374);
nand U8306 (N_8306,N_1954,N_1436);
and U8307 (N_8307,N_4352,N_1665);
nor U8308 (N_8308,N_258,N_4903);
nor U8309 (N_8309,N_3455,N_3306);
or U8310 (N_8310,N_588,N_973);
nand U8311 (N_8311,N_2057,N_3874);
nand U8312 (N_8312,N_4412,N_2511);
nor U8313 (N_8313,N_2925,N_690);
xor U8314 (N_8314,N_4501,N_2709);
or U8315 (N_8315,N_3039,N_2855);
xor U8316 (N_8316,N_1820,N_4474);
xor U8317 (N_8317,N_643,N_566);
nor U8318 (N_8318,N_4870,N_2615);
nor U8319 (N_8319,N_1880,N_1818);
xor U8320 (N_8320,N_4378,N_3405);
nor U8321 (N_8321,N_2531,N_1517);
nand U8322 (N_8322,N_2824,N_2847);
xnor U8323 (N_8323,N_411,N_940);
nor U8324 (N_8324,N_966,N_4247);
and U8325 (N_8325,N_2736,N_3430);
nor U8326 (N_8326,N_4421,N_1945);
nand U8327 (N_8327,N_4241,N_4682);
xor U8328 (N_8328,N_82,N_2563);
xor U8329 (N_8329,N_3803,N_695);
and U8330 (N_8330,N_3863,N_2489);
xnor U8331 (N_8331,N_672,N_2980);
nand U8332 (N_8332,N_2221,N_4362);
xnor U8333 (N_8333,N_2108,N_1789);
nor U8334 (N_8334,N_1624,N_1061);
xor U8335 (N_8335,N_1015,N_2001);
and U8336 (N_8336,N_3125,N_2170);
xnor U8337 (N_8337,N_3133,N_2785);
nand U8338 (N_8338,N_2860,N_2234);
nor U8339 (N_8339,N_2978,N_944);
or U8340 (N_8340,N_727,N_440);
nand U8341 (N_8341,N_4609,N_1963);
xnor U8342 (N_8342,N_3103,N_2142);
xnor U8343 (N_8343,N_1726,N_887);
xor U8344 (N_8344,N_2097,N_1427);
or U8345 (N_8345,N_1705,N_2202);
xor U8346 (N_8346,N_4675,N_4246);
and U8347 (N_8347,N_1613,N_174);
nand U8348 (N_8348,N_1968,N_3030);
or U8349 (N_8349,N_4670,N_1145);
and U8350 (N_8350,N_4436,N_792);
xnor U8351 (N_8351,N_2110,N_4220);
nor U8352 (N_8352,N_4044,N_2789);
or U8353 (N_8353,N_2734,N_182);
nor U8354 (N_8354,N_1971,N_527);
nand U8355 (N_8355,N_3210,N_3090);
and U8356 (N_8356,N_2909,N_820);
xor U8357 (N_8357,N_2190,N_2622);
nand U8358 (N_8358,N_2207,N_3968);
and U8359 (N_8359,N_4510,N_3712);
nor U8360 (N_8360,N_4892,N_3719);
or U8361 (N_8361,N_1783,N_708);
nand U8362 (N_8362,N_2692,N_419);
and U8363 (N_8363,N_978,N_493);
or U8364 (N_8364,N_3128,N_4157);
or U8365 (N_8365,N_4649,N_4308);
and U8366 (N_8366,N_852,N_3018);
and U8367 (N_8367,N_3884,N_4559);
xor U8368 (N_8368,N_4808,N_3483);
nand U8369 (N_8369,N_4706,N_2194);
or U8370 (N_8370,N_3680,N_4144);
or U8371 (N_8371,N_3225,N_4030);
or U8372 (N_8372,N_720,N_3871);
nand U8373 (N_8373,N_3102,N_3844);
nand U8374 (N_8374,N_1694,N_110);
nor U8375 (N_8375,N_2521,N_821);
nand U8376 (N_8376,N_4249,N_592);
xor U8377 (N_8377,N_4755,N_2147);
nor U8378 (N_8378,N_4279,N_827);
nand U8379 (N_8379,N_4880,N_143);
xor U8380 (N_8380,N_4495,N_4313);
and U8381 (N_8381,N_2976,N_1417);
and U8382 (N_8382,N_1320,N_3785);
or U8383 (N_8383,N_2902,N_1302);
xor U8384 (N_8384,N_4655,N_1959);
and U8385 (N_8385,N_424,N_4016);
xnor U8386 (N_8386,N_1452,N_1612);
nor U8387 (N_8387,N_548,N_2079);
xor U8388 (N_8388,N_3906,N_4755);
and U8389 (N_8389,N_902,N_1193);
xor U8390 (N_8390,N_161,N_3019);
or U8391 (N_8391,N_775,N_1997);
nand U8392 (N_8392,N_94,N_2814);
and U8393 (N_8393,N_1752,N_1121);
xor U8394 (N_8394,N_2808,N_3552);
or U8395 (N_8395,N_3254,N_2494);
or U8396 (N_8396,N_3937,N_2457);
or U8397 (N_8397,N_354,N_933);
or U8398 (N_8398,N_536,N_1160);
nor U8399 (N_8399,N_3664,N_3506);
and U8400 (N_8400,N_2126,N_3937);
nand U8401 (N_8401,N_1729,N_2569);
and U8402 (N_8402,N_291,N_4823);
nor U8403 (N_8403,N_3015,N_2385);
xor U8404 (N_8404,N_1014,N_3735);
nor U8405 (N_8405,N_4500,N_561);
nand U8406 (N_8406,N_2746,N_4460);
nor U8407 (N_8407,N_2537,N_4554);
nor U8408 (N_8408,N_4236,N_4047);
or U8409 (N_8409,N_2408,N_4458);
nor U8410 (N_8410,N_3184,N_1049);
nand U8411 (N_8411,N_4570,N_535);
nor U8412 (N_8412,N_3950,N_3600);
and U8413 (N_8413,N_593,N_1832);
or U8414 (N_8414,N_2713,N_439);
and U8415 (N_8415,N_1598,N_3492);
nand U8416 (N_8416,N_518,N_4364);
or U8417 (N_8417,N_2810,N_4674);
or U8418 (N_8418,N_2128,N_3793);
nand U8419 (N_8419,N_4691,N_4703);
nor U8420 (N_8420,N_363,N_4662);
and U8421 (N_8421,N_1847,N_1976);
nand U8422 (N_8422,N_1291,N_4836);
nand U8423 (N_8423,N_1235,N_2101);
or U8424 (N_8424,N_3850,N_3593);
nor U8425 (N_8425,N_4343,N_1760);
nor U8426 (N_8426,N_1369,N_3640);
nand U8427 (N_8427,N_73,N_367);
and U8428 (N_8428,N_664,N_1242);
or U8429 (N_8429,N_2705,N_3564);
and U8430 (N_8430,N_1750,N_1340);
nand U8431 (N_8431,N_1567,N_4932);
or U8432 (N_8432,N_3109,N_688);
and U8433 (N_8433,N_3195,N_2944);
xnor U8434 (N_8434,N_1069,N_4119);
and U8435 (N_8435,N_4679,N_965);
or U8436 (N_8436,N_2643,N_4465);
nand U8437 (N_8437,N_4418,N_3231);
and U8438 (N_8438,N_3991,N_2513);
or U8439 (N_8439,N_4445,N_2543);
xnor U8440 (N_8440,N_3577,N_2492);
nand U8441 (N_8441,N_4892,N_2553);
xor U8442 (N_8442,N_4117,N_3545);
xor U8443 (N_8443,N_3857,N_1310);
and U8444 (N_8444,N_3001,N_1507);
xnor U8445 (N_8445,N_2393,N_4705);
nand U8446 (N_8446,N_1883,N_1);
and U8447 (N_8447,N_1032,N_2196);
and U8448 (N_8448,N_2347,N_4724);
xor U8449 (N_8449,N_4402,N_3860);
and U8450 (N_8450,N_923,N_553);
nor U8451 (N_8451,N_1365,N_2699);
xor U8452 (N_8452,N_3773,N_1232);
and U8453 (N_8453,N_2685,N_1292);
and U8454 (N_8454,N_2104,N_1887);
and U8455 (N_8455,N_2902,N_1576);
nor U8456 (N_8456,N_3567,N_1356);
nor U8457 (N_8457,N_3492,N_2011);
nor U8458 (N_8458,N_34,N_4949);
or U8459 (N_8459,N_878,N_4898);
and U8460 (N_8460,N_3590,N_1344);
xor U8461 (N_8461,N_4298,N_4359);
nor U8462 (N_8462,N_1146,N_1349);
nor U8463 (N_8463,N_252,N_3553);
nand U8464 (N_8464,N_683,N_3351);
xor U8465 (N_8465,N_2639,N_328);
or U8466 (N_8466,N_4775,N_2851);
xnor U8467 (N_8467,N_2041,N_2591);
nor U8468 (N_8468,N_2508,N_706);
and U8469 (N_8469,N_3118,N_2103);
and U8470 (N_8470,N_865,N_1089);
nor U8471 (N_8471,N_1112,N_1162);
xnor U8472 (N_8472,N_73,N_1253);
nand U8473 (N_8473,N_3596,N_4879);
nor U8474 (N_8474,N_2830,N_3974);
and U8475 (N_8475,N_61,N_762);
nor U8476 (N_8476,N_1444,N_4967);
nand U8477 (N_8477,N_2565,N_2842);
nor U8478 (N_8478,N_1702,N_2999);
and U8479 (N_8479,N_2119,N_78);
xor U8480 (N_8480,N_980,N_1353);
xor U8481 (N_8481,N_3129,N_3040);
xnor U8482 (N_8482,N_3500,N_840);
xor U8483 (N_8483,N_111,N_1415);
nor U8484 (N_8484,N_73,N_683);
xor U8485 (N_8485,N_3647,N_4741);
nand U8486 (N_8486,N_24,N_1693);
nor U8487 (N_8487,N_3709,N_1834);
and U8488 (N_8488,N_3689,N_2738);
nor U8489 (N_8489,N_3632,N_4495);
and U8490 (N_8490,N_43,N_248);
nor U8491 (N_8491,N_4205,N_3827);
or U8492 (N_8492,N_2419,N_1167);
xor U8493 (N_8493,N_4912,N_3844);
nor U8494 (N_8494,N_681,N_2529);
xnor U8495 (N_8495,N_2412,N_4515);
xnor U8496 (N_8496,N_3047,N_4838);
nand U8497 (N_8497,N_2836,N_3307);
nor U8498 (N_8498,N_4929,N_1272);
xnor U8499 (N_8499,N_629,N_3217);
nor U8500 (N_8500,N_710,N_326);
nor U8501 (N_8501,N_944,N_369);
or U8502 (N_8502,N_3153,N_3224);
nor U8503 (N_8503,N_4600,N_1053);
and U8504 (N_8504,N_659,N_1803);
xor U8505 (N_8505,N_2138,N_1597);
nor U8506 (N_8506,N_2984,N_5);
or U8507 (N_8507,N_4991,N_1992);
xor U8508 (N_8508,N_3768,N_1671);
xor U8509 (N_8509,N_2925,N_1359);
xnor U8510 (N_8510,N_3649,N_1182);
nand U8511 (N_8511,N_426,N_389);
nor U8512 (N_8512,N_160,N_806);
xor U8513 (N_8513,N_1615,N_1796);
nor U8514 (N_8514,N_421,N_601);
nor U8515 (N_8515,N_1875,N_1782);
or U8516 (N_8516,N_2248,N_1832);
or U8517 (N_8517,N_1017,N_646);
and U8518 (N_8518,N_4343,N_2770);
and U8519 (N_8519,N_4710,N_1679);
or U8520 (N_8520,N_3584,N_4468);
xnor U8521 (N_8521,N_1200,N_2821);
or U8522 (N_8522,N_3790,N_3944);
nand U8523 (N_8523,N_669,N_4472);
xor U8524 (N_8524,N_1309,N_3914);
nand U8525 (N_8525,N_3347,N_2702);
nand U8526 (N_8526,N_232,N_1608);
or U8527 (N_8527,N_2598,N_4413);
or U8528 (N_8528,N_4744,N_4134);
nor U8529 (N_8529,N_654,N_4261);
xor U8530 (N_8530,N_4500,N_1963);
xor U8531 (N_8531,N_2770,N_3782);
nor U8532 (N_8532,N_3513,N_4851);
nand U8533 (N_8533,N_3262,N_997);
and U8534 (N_8534,N_4618,N_478);
xnor U8535 (N_8535,N_717,N_1949);
or U8536 (N_8536,N_4018,N_3344);
nand U8537 (N_8537,N_1581,N_3560);
and U8538 (N_8538,N_3883,N_1370);
nor U8539 (N_8539,N_201,N_4244);
nor U8540 (N_8540,N_1967,N_1610);
nand U8541 (N_8541,N_4052,N_3246);
xor U8542 (N_8542,N_1593,N_4658);
nor U8543 (N_8543,N_1565,N_1165);
nand U8544 (N_8544,N_2043,N_1893);
xnor U8545 (N_8545,N_945,N_3142);
or U8546 (N_8546,N_2141,N_2720);
xnor U8547 (N_8547,N_668,N_1660);
nor U8548 (N_8548,N_685,N_671);
nand U8549 (N_8549,N_4330,N_622);
or U8550 (N_8550,N_2972,N_2737);
nor U8551 (N_8551,N_1205,N_1309);
or U8552 (N_8552,N_3680,N_480);
nor U8553 (N_8553,N_756,N_174);
xor U8554 (N_8554,N_720,N_4427);
nand U8555 (N_8555,N_4102,N_1723);
nor U8556 (N_8556,N_862,N_2844);
nor U8557 (N_8557,N_962,N_1614);
and U8558 (N_8558,N_1050,N_2558);
and U8559 (N_8559,N_2033,N_1896);
nand U8560 (N_8560,N_2526,N_2705);
nand U8561 (N_8561,N_65,N_3085);
nand U8562 (N_8562,N_817,N_529);
and U8563 (N_8563,N_2132,N_2493);
or U8564 (N_8564,N_1632,N_710);
xor U8565 (N_8565,N_4356,N_2605);
nor U8566 (N_8566,N_4682,N_2387);
xor U8567 (N_8567,N_4225,N_3468);
or U8568 (N_8568,N_1679,N_3657);
and U8569 (N_8569,N_3055,N_711);
nor U8570 (N_8570,N_1122,N_840);
xnor U8571 (N_8571,N_3390,N_2110);
and U8572 (N_8572,N_4212,N_4613);
nand U8573 (N_8573,N_2212,N_4390);
nor U8574 (N_8574,N_1235,N_3583);
xor U8575 (N_8575,N_4646,N_2667);
xnor U8576 (N_8576,N_2749,N_3475);
nor U8577 (N_8577,N_565,N_4882);
nor U8578 (N_8578,N_2881,N_2742);
or U8579 (N_8579,N_1838,N_609);
nor U8580 (N_8580,N_4736,N_3315);
or U8581 (N_8581,N_3837,N_2565);
and U8582 (N_8582,N_3001,N_3749);
nor U8583 (N_8583,N_2531,N_3993);
or U8584 (N_8584,N_1791,N_164);
or U8585 (N_8585,N_1533,N_2604);
and U8586 (N_8586,N_1185,N_4913);
and U8587 (N_8587,N_3603,N_3308);
or U8588 (N_8588,N_2493,N_1151);
nand U8589 (N_8589,N_4495,N_264);
or U8590 (N_8590,N_358,N_3229);
and U8591 (N_8591,N_1850,N_1912);
xor U8592 (N_8592,N_3372,N_2361);
nor U8593 (N_8593,N_1611,N_622);
nand U8594 (N_8594,N_680,N_1949);
nand U8595 (N_8595,N_4431,N_1496);
nor U8596 (N_8596,N_4487,N_3821);
nor U8597 (N_8597,N_4011,N_3406);
nor U8598 (N_8598,N_3176,N_1956);
nand U8599 (N_8599,N_3652,N_1082);
or U8600 (N_8600,N_2991,N_2194);
or U8601 (N_8601,N_411,N_4336);
nand U8602 (N_8602,N_2483,N_3442);
xnor U8603 (N_8603,N_414,N_2768);
or U8604 (N_8604,N_3482,N_4370);
nor U8605 (N_8605,N_1791,N_4391);
nor U8606 (N_8606,N_1081,N_1173);
nand U8607 (N_8607,N_3125,N_2985);
and U8608 (N_8608,N_889,N_1389);
and U8609 (N_8609,N_2596,N_4358);
and U8610 (N_8610,N_781,N_3353);
nor U8611 (N_8611,N_4590,N_3061);
xor U8612 (N_8612,N_761,N_3624);
or U8613 (N_8613,N_2007,N_2916);
or U8614 (N_8614,N_417,N_2164);
nand U8615 (N_8615,N_1984,N_768);
nor U8616 (N_8616,N_4618,N_29);
nand U8617 (N_8617,N_1689,N_4252);
or U8618 (N_8618,N_3988,N_4793);
and U8619 (N_8619,N_1298,N_4817);
xor U8620 (N_8620,N_4250,N_501);
and U8621 (N_8621,N_2354,N_3950);
xor U8622 (N_8622,N_1435,N_508);
nand U8623 (N_8623,N_121,N_4007);
and U8624 (N_8624,N_2696,N_4090);
nand U8625 (N_8625,N_1320,N_2693);
and U8626 (N_8626,N_699,N_4508);
and U8627 (N_8627,N_277,N_3779);
nor U8628 (N_8628,N_993,N_135);
nand U8629 (N_8629,N_2647,N_974);
nor U8630 (N_8630,N_1860,N_3249);
nand U8631 (N_8631,N_1326,N_1504);
and U8632 (N_8632,N_4551,N_1983);
nor U8633 (N_8633,N_2063,N_3077);
nand U8634 (N_8634,N_2103,N_2975);
nand U8635 (N_8635,N_4029,N_4037);
nor U8636 (N_8636,N_2184,N_2099);
xnor U8637 (N_8637,N_1357,N_2862);
and U8638 (N_8638,N_3547,N_1462);
xor U8639 (N_8639,N_4830,N_293);
nand U8640 (N_8640,N_2732,N_3940);
or U8641 (N_8641,N_838,N_3376);
or U8642 (N_8642,N_3167,N_96);
and U8643 (N_8643,N_4926,N_3238);
or U8644 (N_8644,N_3863,N_935);
nor U8645 (N_8645,N_718,N_2517);
xor U8646 (N_8646,N_4894,N_1443);
nor U8647 (N_8647,N_1270,N_819);
xor U8648 (N_8648,N_724,N_394);
and U8649 (N_8649,N_2010,N_2131);
or U8650 (N_8650,N_2619,N_1375);
or U8651 (N_8651,N_1588,N_1286);
nand U8652 (N_8652,N_4632,N_333);
and U8653 (N_8653,N_3297,N_4081);
nand U8654 (N_8654,N_4710,N_3762);
nor U8655 (N_8655,N_4062,N_2522);
xor U8656 (N_8656,N_684,N_51);
and U8657 (N_8657,N_1132,N_674);
and U8658 (N_8658,N_548,N_3898);
xnor U8659 (N_8659,N_1445,N_2228);
nor U8660 (N_8660,N_4122,N_2499);
xor U8661 (N_8661,N_4782,N_927);
nand U8662 (N_8662,N_2475,N_1972);
nand U8663 (N_8663,N_1302,N_4511);
nor U8664 (N_8664,N_3327,N_216);
nand U8665 (N_8665,N_2449,N_2350);
xnor U8666 (N_8666,N_233,N_4488);
nand U8667 (N_8667,N_602,N_3951);
or U8668 (N_8668,N_3091,N_2307);
and U8669 (N_8669,N_3998,N_2886);
or U8670 (N_8670,N_4125,N_3105);
and U8671 (N_8671,N_1169,N_62);
nor U8672 (N_8672,N_2553,N_401);
nand U8673 (N_8673,N_1282,N_1599);
and U8674 (N_8674,N_3900,N_1193);
nand U8675 (N_8675,N_3404,N_4651);
and U8676 (N_8676,N_4373,N_1483);
or U8677 (N_8677,N_210,N_4504);
and U8678 (N_8678,N_2322,N_515);
nand U8679 (N_8679,N_1628,N_3081);
or U8680 (N_8680,N_4218,N_2572);
and U8681 (N_8681,N_2489,N_3306);
or U8682 (N_8682,N_3801,N_4498);
nand U8683 (N_8683,N_3996,N_2031);
nor U8684 (N_8684,N_4520,N_4030);
or U8685 (N_8685,N_1111,N_3938);
and U8686 (N_8686,N_3887,N_2630);
nor U8687 (N_8687,N_1745,N_3464);
nor U8688 (N_8688,N_4474,N_4107);
nand U8689 (N_8689,N_2951,N_3521);
and U8690 (N_8690,N_3629,N_3728);
nand U8691 (N_8691,N_2223,N_2518);
xnor U8692 (N_8692,N_2564,N_523);
xor U8693 (N_8693,N_4610,N_3729);
and U8694 (N_8694,N_2548,N_368);
or U8695 (N_8695,N_2138,N_3438);
nor U8696 (N_8696,N_298,N_4713);
or U8697 (N_8697,N_2834,N_2287);
or U8698 (N_8698,N_45,N_3930);
or U8699 (N_8699,N_3258,N_815);
or U8700 (N_8700,N_2296,N_551);
or U8701 (N_8701,N_3872,N_1496);
nand U8702 (N_8702,N_3648,N_1590);
xnor U8703 (N_8703,N_4175,N_1587);
nand U8704 (N_8704,N_4,N_4486);
xor U8705 (N_8705,N_578,N_4851);
nor U8706 (N_8706,N_4190,N_558);
nand U8707 (N_8707,N_418,N_1543);
nand U8708 (N_8708,N_1244,N_1279);
nor U8709 (N_8709,N_693,N_3032);
and U8710 (N_8710,N_291,N_4793);
or U8711 (N_8711,N_3864,N_4402);
nand U8712 (N_8712,N_4886,N_1817);
and U8713 (N_8713,N_3592,N_2287);
nor U8714 (N_8714,N_529,N_4657);
nand U8715 (N_8715,N_4736,N_4797);
or U8716 (N_8716,N_1201,N_3068);
or U8717 (N_8717,N_390,N_2973);
or U8718 (N_8718,N_4764,N_2847);
and U8719 (N_8719,N_2035,N_3093);
and U8720 (N_8720,N_3093,N_1163);
or U8721 (N_8721,N_2194,N_2834);
and U8722 (N_8722,N_4821,N_3352);
nand U8723 (N_8723,N_4141,N_791);
xnor U8724 (N_8724,N_535,N_618);
and U8725 (N_8725,N_4936,N_2953);
or U8726 (N_8726,N_4643,N_3595);
nand U8727 (N_8727,N_585,N_3019);
xor U8728 (N_8728,N_4238,N_2098);
nor U8729 (N_8729,N_4827,N_4116);
nor U8730 (N_8730,N_1907,N_1099);
or U8731 (N_8731,N_4639,N_1212);
nor U8732 (N_8732,N_474,N_1432);
nand U8733 (N_8733,N_786,N_572);
or U8734 (N_8734,N_1925,N_2179);
or U8735 (N_8735,N_2951,N_2263);
and U8736 (N_8736,N_1872,N_2948);
xor U8737 (N_8737,N_663,N_694);
and U8738 (N_8738,N_4354,N_2054);
and U8739 (N_8739,N_2495,N_430);
xor U8740 (N_8740,N_4266,N_4223);
or U8741 (N_8741,N_4024,N_883);
and U8742 (N_8742,N_4306,N_1819);
or U8743 (N_8743,N_813,N_4945);
or U8744 (N_8744,N_358,N_4364);
nand U8745 (N_8745,N_556,N_2433);
or U8746 (N_8746,N_1379,N_3591);
nor U8747 (N_8747,N_4551,N_4581);
nor U8748 (N_8748,N_4513,N_1283);
nand U8749 (N_8749,N_2969,N_2607);
or U8750 (N_8750,N_839,N_3908);
nand U8751 (N_8751,N_3423,N_4437);
xor U8752 (N_8752,N_4778,N_4535);
xnor U8753 (N_8753,N_2655,N_3940);
or U8754 (N_8754,N_1762,N_3015);
xnor U8755 (N_8755,N_3169,N_3033);
xnor U8756 (N_8756,N_69,N_399);
or U8757 (N_8757,N_4400,N_1564);
or U8758 (N_8758,N_1548,N_207);
xor U8759 (N_8759,N_515,N_3536);
and U8760 (N_8760,N_3249,N_2826);
nand U8761 (N_8761,N_294,N_2794);
nand U8762 (N_8762,N_4604,N_104);
and U8763 (N_8763,N_605,N_2522);
nand U8764 (N_8764,N_2037,N_4191);
and U8765 (N_8765,N_3840,N_4531);
or U8766 (N_8766,N_2328,N_926);
or U8767 (N_8767,N_220,N_1276);
and U8768 (N_8768,N_541,N_2850);
nor U8769 (N_8769,N_1047,N_3625);
nor U8770 (N_8770,N_2664,N_879);
and U8771 (N_8771,N_4141,N_4236);
xnor U8772 (N_8772,N_4761,N_480);
or U8773 (N_8773,N_2938,N_716);
and U8774 (N_8774,N_614,N_2894);
or U8775 (N_8775,N_3934,N_754);
or U8776 (N_8776,N_4131,N_1410);
or U8777 (N_8777,N_3893,N_2020);
and U8778 (N_8778,N_4462,N_2811);
nor U8779 (N_8779,N_4839,N_4255);
nor U8780 (N_8780,N_3601,N_1019);
or U8781 (N_8781,N_889,N_4659);
nand U8782 (N_8782,N_4791,N_1027);
xnor U8783 (N_8783,N_4317,N_2776);
and U8784 (N_8784,N_3609,N_1299);
and U8785 (N_8785,N_3007,N_3679);
nor U8786 (N_8786,N_3697,N_4721);
or U8787 (N_8787,N_3870,N_4777);
and U8788 (N_8788,N_4224,N_1282);
or U8789 (N_8789,N_2020,N_4866);
and U8790 (N_8790,N_4742,N_2012);
xnor U8791 (N_8791,N_1813,N_3900);
nand U8792 (N_8792,N_255,N_1148);
nand U8793 (N_8793,N_3355,N_856);
xnor U8794 (N_8794,N_434,N_3033);
nand U8795 (N_8795,N_3115,N_1948);
or U8796 (N_8796,N_129,N_2868);
or U8797 (N_8797,N_225,N_1130);
or U8798 (N_8798,N_1828,N_325);
xor U8799 (N_8799,N_2262,N_3590);
nand U8800 (N_8800,N_4564,N_1823);
and U8801 (N_8801,N_592,N_2533);
or U8802 (N_8802,N_2022,N_1094);
xnor U8803 (N_8803,N_1844,N_423);
or U8804 (N_8804,N_1641,N_235);
nor U8805 (N_8805,N_4469,N_1384);
nor U8806 (N_8806,N_2388,N_1812);
nand U8807 (N_8807,N_111,N_3244);
or U8808 (N_8808,N_3050,N_3974);
and U8809 (N_8809,N_376,N_534);
nand U8810 (N_8810,N_2719,N_504);
xor U8811 (N_8811,N_462,N_3387);
and U8812 (N_8812,N_1915,N_748);
nand U8813 (N_8813,N_328,N_2342);
nand U8814 (N_8814,N_1891,N_3911);
and U8815 (N_8815,N_277,N_203);
and U8816 (N_8816,N_703,N_4738);
xor U8817 (N_8817,N_2428,N_2928);
nor U8818 (N_8818,N_3696,N_1769);
or U8819 (N_8819,N_3033,N_1722);
nand U8820 (N_8820,N_103,N_2712);
and U8821 (N_8821,N_2761,N_414);
or U8822 (N_8822,N_2366,N_1313);
nand U8823 (N_8823,N_3201,N_2338);
xor U8824 (N_8824,N_576,N_3016);
nor U8825 (N_8825,N_2043,N_4160);
and U8826 (N_8826,N_3873,N_2737);
or U8827 (N_8827,N_4341,N_540);
nand U8828 (N_8828,N_71,N_1556);
nand U8829 (N_8829,N_3139,N_340);
nand U8830 (N_8830,N_3479,N_4870);
xor U8831 (N_8831,N_1799,N_3524);
and U8832 (N_8832,N_1647,N_1071);
nand U8833 (N_8833,N_1124,N_3077);
xnor U8834 (N_8834,N_2124,N_3670);
nor U8835 (N_8835,N_638,N_961);
xnor U8836 (N_8836,N_1419,N_1362);
nand U8837 (N_8837,N_2267,N_4415);
or U8838 (N_8838,N_2976,N_1585);
nand U8839 (N_8839,N_3710,N_1911);
nand U8840 (N_8840,N_4327,N_554);
or U8841 (N_8841,N_3572,N_847);
and U8842 (N_8842,N_1175,N_4662);
and U8843 (N_8843,N_1465,N_3419);
xor U8844 (N_8844,N_1839,N_2290);
nand U8845 (N_8845,N_2599,N_3002);
and U8846 (N_8846,N_4588,N_3641);
or U8847 (N_8847,N_1208,N_4344);
nand U8848 (N_8848,N_1925,N_2458);
nand U8849 (N_8849,N_966,N_3680);
or U8850 (N_8850,N_562,N_213);
or U8851 (N_8851,N_2149,N_2230);
or U8852 (N_8852,N_2245,N_1406);
or U8853 (N_8853,N_4450,N_3429);
xor U8854 (N_8854,N_4358,N_3281);
and U8855 (N_8855,N_3653,N_1857);
nand U8856 (N_8856,N_2377,N_4242);
nor U8857 (N_8857,N_1123,N_519);
and U8858 (N_8858,N_2076,N_2654);
nand U8859 (N_8859,N_2186,N_4691);
or U8860 (N_8860,N_3160,N_1632);
nor U8861 (N_8861,N_504,N_2110);
or U8862 (N_8862,N_3801,N_1151);
nor U8863 (N_8863,N_309,N_2948);
xnor U8864 (N_8864,N_849,N_283);
or U8865 (N_8865,N_3035,N_3970);
or U8866 (N_8866,N_3736,N_2958);
or U8867 (N_8867,N_1524,N_588);
and U8868 (N_8868,N_3170,N_1160);
and U8869 (N_8869,N_4793,N_1112);
xnor U8870 (N_8870,N_4711,N_1487);
xnor U8871 (N_8871,N_1434,N_3721);
nor U8872 (N_8872,N_4648,N_16);
xor U8873 (N_8873,N_2754,N_3282);
nor U8874 (N_8874,N_1211,N_4682);
nand U8875 (N_8875,N_3354,N_4402);
or U8876 (N_8876,N_3388,N_1880);
xnor U8877 (N_8877,N_2208,N_1147);
and U8878 (N_8878,N_4695,N_733);
nand U8879 (N_8879,N_2423,N_546);
nand U8880 (N_8880,N_3827,N_422);
nand U8881 (N_8881,N_3398,N_3231);
xnor U8882 (N_8882,N_4931,N_694);
or U8883 (N_8883,N_1401,N_1731);
xnor U8884 (N_8884,N_807,N_1960);
nor U8885 (N_8885,N_2954,N_2516);
nor U8886 (N_8886,N_3758,N_883);
nand U8887 (N_8887,N_4626,N_1367);
nand U8888 (N_8888,N_517,N_1485);
or U8889 (N_8889,N_4169,N_642);
nand U8890 (N_8890,N_3132,N_2044);
or U8891 (N_8891,N_1527,N_2119);
xnor U8892 (N_8892,N_4086,N_221);
or U8893 (N_8893,N_4992,N_1335);
nor U8894 (N_8894,N_2865,N_3115);
or U8895 (N_8895,N_3718,N_484);
or U8896 (N_8896,N_1974,N_4706);
nor U8897 (N_8897,N_3513,N_2135);
or U8898 (N_8898,N_4818,N_148);
nor U8899 (N_8899,N_1784,N_4001);
nor U8900 (N_8900,N_3459,N_1266);
nand U8901 (N_8901,N_4624,N_3646);
or U8902 (N_8902,N_2776,N_3488);
xnor U8903 (N_8903,N_2900,N_3478);
and U8904 (N_8904,N_1340,N_4429);
and U8905 (N_8905,N_348,N_2671);
and U8906 (N_8906,N_2110,N_417);
nor U8907 (N_8907,N_2278,N_4796);
or U8908 (N_8908,N_3010,N_3081);
and U8909 (N_8909,N_3575,N_3721);
nor U8910 (N_8910,N_1853,N_3878);
nand U8911 (N_8911,N_824,N_4025);
and U8912 (N_8912,N_4496,N_2574);
nand U8913 (N_8913,N_2586,N_1947);
nor U8914 (N_8914,N_21,N_4328);
or U8915 (N_8915,N_4527,N_1099);
nand U8916 (N_8916,N_3146,N_4657);
xor U8917 (N_8917,N_2014,N_173);
and U8918 (N_8918,N_94,N_1909);
nand U8919 (N_8919,N_4906,N_3297);
nand U8920 (N_8920,N_594,N_978);
and U8921 (N_8921,N_4551,N_1091);
nor U8922 (N_8922,N_2912,N_3032);
or U8923 (N_8923,N_339,N_4146);
nor U8924 (N_8924,N_3823,N_1018);
xnor U8925 (N_8925,N_2549,N_3973);
nor U8926 (N_8926,N_2474,N_2136);
or U8927 (N_8927,N_47,N_920);
and U8928 (N_8928,N_1336,N_1045);
and U8929 (N_8929,N_4,N_2268);
nand U8930 (N_8930,N_1587,N_4615);
xnor U8931 (N_8931,N_3322,N_2279);
nor U8932 (N_8932,N_2449,N_2616);
or U8933 (N_8933,N_3818,N_986);
nand U8934 (N_8934,N_3133,N_4607);
and U8935 (N_8935,N_2548,N_1685);
xor U8936 (N_8936,N_56,N_132);
and U8937 (N_8937,N_2215,N_2187);
xnor U8938 (N_8938,N_2474,N_3307);
nand U8939 (N_8939,N_715,N_102);
nand U8940 (N_8940,N_3064,N_4917);
and U8941 (N_8941,N_4679,N_4359);
nor U8942 (N_8942,N_2544,N_356);
and U8943 (N_8943,N_1097,N_626);
nand U8944 (N_8944,N_2574,N_2640);
nor U8945 (N_8945,N_3967,N_3506);
nor U8946 (N_8946,N_2294,N_2690);
nand U8947 (N_8947,N_915,N_34);
nor U8948 (N_8948,N_1768,N_3505);
and U8949 (N_8949,N_213,N_3910);
and U8950 (N_8950,N_2490,N_3309);
nor U8951 (N_8951,N_3362,N_4069);
nor U8952 (N_8952,N_1822,N_180);
or U8953 (N_8953,N_1539,N_3204);
and U8954 (N_8954,N_3748,N_1516);
and U8955 (N_8955,N_1067,N_635);
or U8956 (N_8956,N_4079,N_4897);
and U8957 (N_8957,N_4659,N_2553);
xor U8958 (N_8958,N_3410,N_589);
xor U8959 (N_8959,N_770,N_1651);
and U8960 (N_8960,N_967,N_1662);
nand U8961 (N_8961,N_507,N_2075);
and U8962 (N_8962,N_143,N_441);
xor U8963 (N_8963,N_4383,N_2677);
xor U8964 (N_8964,N_4770,N_2876);
and U8965 (N_8965,N_4174,N_4766);
nor U8966 (N_8966,N_326,N_2124);
and U8967 (N_8967,N_2845,N_2923);
nor U8968 (N_8968,N_576,N_2283);
and U8969 (N_8969,N_734,N_332);
nand U8970 (N_8970,N_1901,N_1225);
nor U8971 (N_8971,N_4098,N_2620);
xnor U8972 (N_8972,N_576,N_3178);
nor U8973 (N_8973,N_1592,N_2497);
nor U8974 (N_8974,N_4189,N_3577);
nor U8975 (N_8975,N_4129,N_306);
xnor U8976 (N_8976,N_88,N_1704);
and U8977 (N_8977,N_3799,N_3613);
or U8978 (N_8978,N_1167,N_3789);
or U8979 (N_8979,N_2739,N_1854);
xnor U8980 (N_8980,N_406,N_1231);
and U8981 (N_8981,N_3665,N_3764);
nand U8982 (N_8982,N_3288,N_629);
nor U8983 (N_8983,N_3467,N_3343);
and U8984 (N_8984,N_38,N_2455);
xor U8985 (N_8985,N_4058,N_1133);
nand U8986 (N_8986,N_27,N_2954);
nand U8987 (N_8987,N_3056,N_2302);
nor U8988 (N_8988,N_2401,N_4784);
or U8989 (N_8989,N_1027,N_2171);
or U8990 (N_8990,N_1013,N_2753);
and U8991 (N_8991,N_2146,N_3625);
and U8992 (N_8992,N_1077,N_782);
xor U8993 (N_8993,N_1997,N_2732);
xor U8994 (N_8994,N_4250,N_1614);
or U8995 (N_8995,N_957,N_2289);
nor U8996 (N_8996,N_4679,N_2112);
nor U8997 (N_8997,N_1451,N_710);
xor U8998 (N_8998,N_2215,N_4650);
and U8999 (N_8999,N_3686,N_3134);
nor U9000 (N_9000,N_2746,N_1798);
or U9001 (N_9001,N_1763,N_3321);
or U9002 (N_9002,N_4892,N_3713);
or U9003 (N_9003,N_361,N_3024);
xnor U9004 (N_9004,N_1494,N_4747);
or U9005 (N_9005,N_3521,N_2358);
xnor U9006 (N_9006,N_4291,N_24);
and U9007 (N_9007,N_1801,N_756);
xnor U9008 (N_9008,N_2510,N_812);
xnor U9009 (N_9009,N_2019,N_4147);
nand U9010 (N_9010,N_4849,N_1185);
nor U9011 (N_9011,N_3029,N_4870);
and U9012 (N_9012,N_2933,N_3493);
and U9013 (N_9013,N_990,N_2945);
or U9014 (N_9014,N_2333,N_3430);
nand U9015 (N_9015,N_4258,N_2531);
and U9016 (N_9016,N_3700,N_407);
nor U9017 (N_9017,N_1052,N_4709);
or U9018 (N_9018,N_2649,N_1145);
nand U9019 (N_9019,N_1446,N_1646);
nor U9020 (N_9020,N_253,N_506);
xor U9021 (N_9021,N_4201,N_2266);
and U9022 (N_9022,N_209,N_215);
nand U9023 (N_9023,N_3404,N_3987);
or U9024 (N_9024,N_3461,N_392);
or U9025 (N_9025,N_1452,N_1003);
and U9026 (N_9026,N_2758,N_1668);
and U9027 (N_9027,N_4448,N_1092);
or U9028 (N_9028,N_2394,N_4742);
xnor U9029 (N_9029,N_4743,N_1975);
and U9030 (N_9030,N_1432,N_13);
nor U9031 (N_9031,N_1982,N_3375);
or U9032 (N_9032,N_2398,N_3754);
xnor U9033 (N_9033,N_4090,N_1711);
and U9034 (N_9034,N_359,N_1300);
or U9035 (N_9035,N_1251,N_4567);
and U9036 (N_9036,N_1302,N_4447);
xnor U9037 (N_9037,N_624,N_1721);
or U9038 (N_9038,N_330,N_2042);
xnor U9039 (N_9039,N_1274,N_252);
or U9040 (N_9040,N_2469,N_2113);
or U9041 (N_9041,N_2227,N_1394);
or U9042 (N_9042,N_1264,N_1095);
or U9043 (N_9043,N_1002,N_2286);
and U9044 (N_9044,N_4414,N_4604);
or U9045 (N_9045,N_3030,N_1031);
and U9046 (N_9046,N_2972,N_3039);
or U9047 (N_9047,N_1790,N_292);
xor U9048 (N_9048,N_794,N_1784);
nand U9049 (N_9049,N_4505,N_1166);
or U9050 (N_9050,N_545,N_4188);
or U9051 (N_9051,N_4293,N_933);
nor U9052 (N_9052,N_2713,N_674);
nor U9053 (N_9053,N_1621,N_2337);
xor U9054 (N_9054,N_1263,N_2689);
nand U9055 (N_9055,N_1484,N_309);
and U9056 (N_9056,N_1174,N_4703);
nand U9057 (N_9057,N_90,N_1232);
nor U9058 (N_9058,N_2176,N_63);
nor U9059 (N_9059,N_1942,N_3159);
or U9060 (N_9060,N_1453,N_1808);
nand U9061 (N_9061,N_2549,N_4354);
xnor U9062 (N_9062,N_3461,N_3896);
xor U9063 (N_9063,N_4302,N_1853);
nand U9064 (N_9064,N_4706,N_731);
nor U9065 (N_9065,N_395,N_4560);
xor U9066 (N_9066,N_1564,N_3576);
nand U9067 (N_9067,N_2531,N_2795);
nand U9068 (N_9068,N_1312,N_2296);
nand U9069 (N_9069,N_4504,N_4665);
xnor U9070 (N_9070,N_779,N_2124);
nand U9071 (N_9071,N_3535,N_2326);
xnor U9072 (N_9072,N_3343,N_2370);
or U9073 (N_9073,N_4078,N_2552);
nand U9074 (N_9074,N_4757,N_829);
and U9075 (N_9075,N_3446,N_3410);
and U9076 (N_9076,N_3532,N_3552);
and U9077 (N_9077,N_2488,N_1055);
nand U9078 (N_9078,N_4520,N_1384);
nand U9079 (N_9079,N_4655,N_3112);
nor U9080 (N_9080,N_2669,N_1143);
or U9081 (N_9081,N_2629,N_2717);
nor U9082 (N_9082,N_3970,N_2247);
nor U9083 (N_9083,N_275,N_4038);
and U9084 (N_9084,N_3052,N_4742);
or U9085 (N_9085,N_4355,N_1128);
xor U9086 (N_9086,N_431,N_4062);
nand U9087 (N_9087,N_4895,N_3809);
or U9088 (N_9088,N_4918,N_2020);
nor U9089 (N_9089,N_1773,N_4452);
and U9090 (N_9090,N_2788,N_142);
and U9091 (N_9091,N_724,N_3775);
nor U9092 (N_9092,N_327,N_589);
nor U9093 (N_9093,N_2667,N_4804);
and U9094 (N_9094,N_534,N_2255);
and U9095 (N_9095,N_2695,N_2807);
nor U9096 (N_9096,N_1507,N_3666);
xnor U9097 (N_9097,N_4540,N_3298);
or U9098 (N_9098,N_2107,N_3537);
and U9099 (N_9099,N_3691,N_876);
or U9100 (N_9100,N_2815,N_1430);
nor U9101 (N_9101,N_2830,N_2344);
nand U9102 (N_9102,N_4999,N_966);
xor U9103 (N_9103,N_581,N_672);
xor U9104 (N_9104,N_3945,N_3194);
nand U9105 (N_9105,N_576,N_71);
nand U9106 (N_9106,N_4701,N_304);
or U9107 (N_9107,N_4234,N_1873);
xor U9108 (N_9108,N_3703,N_4659);
xor U9109 (N_9109,N_280,N_1599);
xnor U9110 (N_9110,N_3286,N_137);
nand U9111 (N_9111,N_3761,N_3187);
or U9112 (N_9112,N_842,N_3125);
nor U9113 (N_9113,N_2947,N_2688);
nor U9114 (N_9114,N_806,N_2412);
nand U9115 (N_9115,N_955,N_4436);
nor U9116 (N_9116,N_226,N_3626);
xor U9117 (N_9117,N_4303,N_2109);
and U9118 (N_9118,N_2960,N_1328);
xnor U9119 (N_9119,N_4613,N_4199);
and U9120 (N_9120,N_6,N_3460);
nand U9121 (N_9121,N_3546,N_699);
xor U9122 (N_9122,N_2819,N_2780);
nor U9123 (N_9123,N_4018,N_325);
and U9124 (N_9124,N_4876,N_3167);
nor U9125 (N_9125,N_305,N_2391);
nor U9126 (N_9126,N_4175,N_1393);
or U9127 (N_9127,N_2815,N_3127);
nand U9128 (N_9128,N_4547,N_1430);
and U9129 (N_9129,N_4292,N_4053);
and U9130 (N_9130,N_3749,N_640);
and U9131 (N_9131,N_1991,N_3884);
and U9132 (N_9132,N_4322,N_4949);
nand U9133 (N_9133,N_3431,N_4370);
xor U9134 (N_9134,N_1469,N_2839);
or U9135 (N_9135,N_3326,N_241);
nand U9136 (N_9136,N_2039,N_2028);
nand U9137 (N_9137,N_4208,N_2439);
nor U9138 (N_9138,N_4228,N_107);
xnor U9139 (N_9139,N_4833,N_3709);
nor U9140 (N_9140,N_1255,N_385);
nand U9141 (N_9141,N_3892,N_1281);
and U9142 (N_9142,N_3147,N_4518);
nor U9143 (N_9143,N_271,N_1023);
xor U9144 (N_9144,N_1190,N_1299);
xnor U9145 (N_9145,N_1836,N_1677);
nand U9146 (N_9146,N_2801,N_2405);
xnor U9147 (N_9147,N_3614,N_1546);
nor U9148 (N_9148,N_1713,N_2478);
nor U9149 (N_9149,N_2621,N_2205);
nand U9150 (N_9150,N_348,N_2902);
xnor U9151 (N_9151,N_204,N_1598);
xnor U9152 (N_9152,N_4570,N_3191);
xnor U9153 (N_9153,N_2370,N_421);
nand U9154 (N_9154,N_3999,N_3726);
nand U9155 (N_9155,N_3775,N_58);
xnor U9156 (N_9156,N_921,N_1900);
or U9157 (N_9157,N_3479,N_2538);
and U9158 (N_9158,N_4416,N_3405);
nand U9159 (N_9159,N_573,N_1283);
and U9160 (N_9160,N_927,N_1466);
and U9161 (N_9161,N_1710,N_1);
xnor U9162 (N_9162,N_3181,N_1423);
and U9163 (N_9163,N_1701,N_3425);
and U9164 (N_9164,N_1578,N_539);
nor U9165 (N_9165,N_3758,N_2724);
or U9166 (N_9166,N_3687,N_2141);
nor U9167 (N_9167,N_615,N_202);
xnor U9168 (N_9168,N_3885,N_4223);
nor U9169 (N_9169,N_708,N_2249);
nand U9170 (N_9170,N_2929,N_2756);
and U9171 (N_9171,N_532,N_3872);
or U9172 (N_9172,N_3380,N_4605);
and U9173 (N_9173,N_1509,N_3938);
nand U9174 (N_9174,N_3209,N_4102);
xnor U9175 (N_9175,N_3283,N_817);
and U9176 (N_9176,N_1594,N_3707);
xnor U9177 (N_9177,N_1566,N_2761);
xnor U9178 (N_9178,N_3365,N_4437);
nor U9179 (N_9179,N_3586,N_1401);
xor U9180 (N_9180,N_4507,N_929);
and U9181 (N_9181,N_4845,N_154);
or U9182 (N_9182,N_436,N_63);
nor U9183 (N_9183,N_1796,N_4998);
or U9184 (N_9184,N_3680,N_703);
and U9185 (N_9185,N_1041,N_2842);
or U9186 (N_9186,N_3651,N_4879);
xor U9187 (N_9187,N_1163,N_3274);
nor U9188 (N_9188,N_2257,N_2055);
xnor U9189 (N_9189,N_476,N_1599);
xor U9190 (N_9190,N_350,N_4532);
nand U9191 (N_9191,N_1341,N_1749);
or U9192 (N_9192,N_2325,N_4558);
nor U9193 (N_9193,N_2604,N_366);
xor U9194 (N_9194,N_3124,N_2282);
xnor U9195 (N_9195,N_4496,N_4104);
xor U9196 (N_9196,N_3063,N_1247);
nand U9197 (N_9197,N_409,N_3141);
or U9198 (N_9198,N_3208,N_3230);
xnor U9199 (N_9199,N_2289,N_2705);
xnor U9200 (N_9200,N_3137,N_4327);
xnor U9201 (N_9201,N_4174,N_3884);
nand U9202 (N_9202,N_891,N_3220);
nor U9203 (N_9203,N_5,N_1871);
or U9204 (N_9204,N_4968,N_1186);
nand U9205 (N_9205,N_3848,N_3777);
nor U9206 (N_9206,N_767,N_1855);
nand U9207 (N_9207,N_4863,N_1259);
and U9208 (N_9208,N_832,N_3461);
xor U9209 (N_9209,N_2701,N_2009);
nand U9210 (N_9210,N_262,N_3823);
xor U9211 (N_9211,N_3410,N_2704);
or U9212 (N_9212,N_4014,N_1154);
or U9213 (N_9213,N_2835,N_466);
and U9214 (N_9214,N_3169,N_1242);
nand U9215 (N_9215,N_221,N_10);
xnor U9216 (N_9216,N_2866,N_3706);
and U9217 (N_9217,N_4894,N_1403);
xnor U9218 (N_9218,N_422,N_2886);
nor U9219 (N_9219,N_1600,N_286);
xnor U9220 (N_9220,N_78,N_4239);
or U9221 (N_9221,N_4258,N_2319);
or U9222 (N_9222,N_4126,N_45);
and U9223 (N_9223,N_110,N_374);
xnor U9224 (N_9224,N_3956,N_2558);
xor U9225 (N_9225,N_3601,N_2124);
nand U9226 (N_9226,N_1922,N_1736);
or U9227 (N_9227,N_2780,N_2106);
nand U9228 (N_9228,N_728,N_915);
or U9229 (N_9229,N_4943,N_3024);
nand U9230 (N_9230,N_127,N_2560);
nor U9231 (N_9231,N_1228,N_328);
or U9232 (N_9232,N_3667,N_328);
xor U9233 (N_9233,N_1207,N_1467);
and U9234 (N_9234,N_2642,N_101);
nor U9235 (N_9235,N_4163,N_4827);
and U9236 (N_9236,N_1817,N_1604);
and U9237 (N_9237,N_4975,N_819);
nand U9238 (N_9238,N_4700,N_1750);
or U9239 (N_9239,N_3214,N_299);
or U9240 (N_9240,N_3695,N_1934);
or U9241 (N_9241,N_1175,N_3765);
xor U9242 (N_9242,N_4095,N_785);
nand U9243 (N_9243,N_3806,N_1785);
or U9244 (N_9244,N_2675,N_2674);
and U9245 (N_9245,N_1945,N_3355);
xor U9246 (N_9246,N_4567,N_2128);
xor U9247 (N_9247,N_1551,N_3667);
and U9248 (N_9248,N_4567,N_452);
nor U9249 (N_9249,N_913,N_59);
nor U9250 (N_9250,N_4502,N_3394);
and U9251 (N_9251,N_3561,N_4568);
nor U9252 (N_9252,N_1980,N_4380);
nor U9253 (N_9253,N_3564,N_3083);
nand U9254 (N_9254,N_3074,N_3723);
xnor U9255 (N_9255,N_982,N_1907);
nand U9256 (N_9256,N_4725,N_4071);
nand U9257 (N_9257,N_1431,N_2650);
and U9258 (N_9258,N_1304,N_4581);
or U9259 (N_9259,N_529,N_4192);
xnor U9260 (N_9260,N_350,N_755);
or U9261 (N_9261,N_3538,N_3712);
and U9262 (N_9262,N_2341,N_381);
xnor U9263 (N_9263,N_4403,N_2875);
xnor U9264 (N_9264,N_1162,N_1350);
and U9265 (N_9265,N_142,N_3928);
xnor U9266 (N_9266,N_1321,N_4450);
xnor U9267 (N_9267,N_3247,N_3647);
nor U9268 (N_9268,N_3280,N_2450);
nor U9269 (N_9269,N_3975,N_3581);
xor U9270 (N_9270,N_1564,N_1486);
and U9271 (N_9271,N_2865,N_1266);
xor U9272 (N_9272,N_482,N_2407);
and U9273 (N_9273,N_1428,N_1901);
xor U9274 (N_9274,N_3368,N_1033);
nor U9275 (N_9275,N_1630,N_3681);
and U9276 (N_9276,N_2909,N_1387);
nor U9277 (N_9277,N_539,N_955);
or U9278 (N_9278,N_3215,N_78);
nor U9279 (N_9279,N_2961,N_1413);
or U9280 (N_9280,N_3896,N_405);
nor U9281 (N_9281,N_66,N_2222);
nor U9282 (N_9282,N_4691,N_1694);
and U9283 (N_9283,N_1716,N_3510);
xor U9284 (N_9284,N_3133,N_946);
xnor U9285 (N_9285,N_2701,N_4698);
and U9286 (N_9286,N_1552,N_3957);
and U9287 (N_9287,N_2163,N_4738);
xnor U9288 (N_9288,N_1966,N_1250);
nor U9289 (N_9289,N_1974,N_2838);
nor U9290 (N_9290,N_4476,N_603);
nand U9291 (N_9291,N_216,N_3800);
and U9292 (N_9292,N_4288,N_2523);
nor U9293 (N_9293,N_4666,N_2058);
nor U9294 (N_9294,N_1896,N_677);
and U9295 (N_9295,N_3519,N_1024);
xor U9296 (N_9296,N_3093,N_4805);
and U9297 (N_9297,N_2975,N_208);
nand U9298 (N_9298,N_1749,N_4229);
or U9299 (N_9299,N_4319,N_4244);
nor U9300 (N_9300,N_2136,N_2616);
nand U9301 (N_9301,N_1858,N_4259);
nand U9302 (N_9302,N_1562,N_3208);
xnor U9303 (N_9303,N_3991,N_2067);
and U9304 (N_9304,N_2619,N_4120);
xor U9305 (N_9305,N_1913,N_801);
nand U9306 (N_9306,N_340,N_2272);
xnor U9307 (N_9307,N_4678,N_4378);
nand U9308 (N_9308,N_2239,N_2257);
and U9309 (N_9309,N_119,N_35);
nand U9310 (N_9310,N_1691,N_774);
and U9311 (N_9311,N_1856,N_1538);
and U9312 (N_9312,N_3056,N_4324);
and U9313 (N_9313,N_1776,N_2516);
nand U9314 (N_9314,N_2828,N_1052);
nand U9315 (N_9315,N_30,N_3968);
nor U9316 (N_9316,N_2440,N_2400);
nand U9317 (N_9317,N_3868,N_462);
or U9318 (N_9318,N_824,N_2357);
nand U9319 (N_9319,N_1634,N_2113);
nor U9320 (N_9320,N_2094,N_354);
nand U9321 (N_9321,N_2702,N_4248);
xor U9322 (N_9322,N_3199,N_806);
or U9323 (N_9323,N_3748,N_3152);
xnor U9324 (N_9324,N_1628,N_4477);
nor U9325 (N_9325,N_1442,N_2706);
or U9326 (N_9326,N_3058,N_3133);
nand U9327 (N_9327,N_398,N_412);
or U9328 (N_9328,N_4941,N_70);
and U9329 (N_9329,N_651,N_4204);
nand U9330 (N_9330,N_977,N_1020);
or U9331 (N_9331,N_2623,N_3602);
or U9332 (N_9332,N_151,N_859);
nor U9333 (N_9333,N_644,N_1773);
nor U9334 (N_9334,N_2196,N_2430);
xor U9335 (N_9335,N_4797,N_4219);
and U9336 (N_9336,N_3064,N_1040);
nor U9337 (N_9337,N_2405,N_124);
nor U9338 (N_9338,N_2189,N_693);
and U9339 (N_9339,N_4713,N_1763);
nand U9340 (N_9340,N_1864,N_2860);
or U9341 (N_9341,N_4239,N_2401);
or U9342 (N_9342,N_2404,N_739);
and U9343 (N_9343,N_3585,N_158);
xnor U9344 (N_9344,N_1943,N_3536);
and U9345 (N_9345,N_4288,N_4046);
or U9346 (N_9346,N_72,N_3701);
or U9347 (N_9347,N_1604,N_1363);
or U9348 (N_9348,N_3271,N_1328);
and U9349 (N_9349,N_2045,N_2492);
nand U9350 (N_9350,N_1032,N_1994);
nor U9351 (N_9351,N_3503,N_2465);
nor U9352 (N_9352,N_2709,N_3033);
nand U9353 (N_9353,N_2558,N_3555);
or U9354 (N_9354,N_118,N_1833);
xnor U9355 (N_9355,N_1463,N_1982);
nand U9356 (N_9356,N_670,N_3509);
xor U9357 (N_9357,N_1122,N_30);
nand U9358 (N_9358,N_3042,N_655);
nor U9359 (N_9359,N_4415,N_3577);
nand U9360 (N_9360,N_3660,N_3097);
nor U9361 (N_9361,N_507,N_2024);
and U9362 (N_9362,N_3329,N_3822);
nand U9363 (N_9363,N_431,N_3427);
xor U9364 (N_9364,N_535,N_1576);
nand U9365 (N_9365,N_3378,N_4987);
nor U9366 (N_9366,N_1614,N_4717);
nor U9367 (N_9367,N_1757,N_4349);
or U9368 (N_9368,N_2404,N_4665);
or U9369 (N_9369,N_4333,N_3277);
nor U9370 (N_9370,N_1150,N_3102);
nor U9371 (N_9371,N_1292,N_2564);
nor U9372 (N_9372,N_1936,N_4780);
or U9373 (N_9373,N_1350,N_4101);
nor U9374 (N_9374,N_2003,N_3465);
xor U9375 (N_9375,N_152,N_371);
nor U9376 (N_9376,N_4130,N_685);
nor U9377 (N_9377,N_4901,N_1686);
nand U9378 (N_9378,N_159,N_605);
xor U9379 (N_9379,N_4895,N_2394);
nand U9380 (N_9380,N_270,N_3521);
nand U9381 (N_9381,N_3617,N_1912);
or U9382 (N_9382,N_608,N_4950);
nor U9383 (N_9383,N_1489,N_2646);
xnor U9384 (N_9384,N_2537,N_1600);
xor U9385 (N_9385,N_2838,N_2279);
xor U9386 (N_9386,N_2850,N_3146);
nand U9387 (N_9387,N_849,N_3987);
or U9388 (N_9388,N_4161,N_4412);
or U9389 (N_9389,N_2334,N_4720);
nand U9390 (N_9390,N_4718,N_1019);
nor U9391 (N_9391,N_3483,N_715);
nor U9392 (N_9392,N_813,N_4848);
nor U9393 (N_9393,N_4388,N_1057);
nor U9394 (N_9394,N_975,N_684);
nand U9395 (N_9395,N_1933,N_2203);
nor U9396 (N_9396,N_4270,N_1136);
nand U9397 (N_9397,N_2045,N_1956);
xnor U9398 (N_9398,N_4113,N_2798);
nand U9399 (N_9399,N_1914,N_857);
or U9400 (N_9400,N_1474,N_3930);
and U9401 (N_9401,N_1331,N_3460);
xor U9402 (N_9402,N_2297,N_664);
nor U9403 (N_9403,N_1797,N_4983);
xor U9404 (N_9404,N_3885,N_4875);
nor U9405 (N_9405,N_2268,N_1476);
nor U9406 (N_9406,N_2475,N_114);
or U9407 (N_9407,N_4370,N_2237);
nand U9408 (N_9408,N_383,N_3351);
nor U9409 (N_9409,N_2251,N_4574);
or U9410 (N_9410,N_3180,N_2136);
xnor U9411 (N_9411,N_611,N_3007);
and U9412 (N_9412,N_3126,N_2021);
nand U9413 (N_9413,N_1137,N_3104);
nand U9414 (N_9414,N_4977,N_2010);
nand U9415 (N_9415,N_4516,N_482);
nand U9416 (N_9416,N_2528,N_2005);
or U9417 (N_9417,N_1783,N_366);
nand U9418 (N_9418,N_4198,N_4723);
nor U9419 (N_9419,N_266,N_1786);
nor U9420 (N_9420,N_96,N_4268);
nand U9421 (N_9421,N_2393,N_1485);
nand U9422 (N_9422,N_4617,N_3315);
nand U9423 (N_9423,N_553,N_3200);
nand U9424 (N_9424,N_1280,N_2886);
nand U9425 (N_9425,N_3649,N_4478);
or U9426 (N_9426,N_2273,N_133);
nand U9427 (N_9427,N_3287,N_2743);
xnor U9428 (N_9428,N_2050,N_2067);
xor U9429 (N_9429,N_4768,N_1236);
and U9430 (N_9430,N_1810,N_1521);
nor U9431 (N_9431,N_4196,N_994);
or U9432 (N_9432,N_1745,N_870);
and U9433 (N_9433,N_1063,N_3035);
or U9434 (N_9434,N_3714,N_918);
xor U9435 (N_9435,N_1390,N_3974);
xor U9436 (N_9436,N_1120,N_3991);
nor U9437 (N_9437,N_1325,N_3035);
nand U9438 (N_9438,N_4418,N_1116);
or U9439 (N_9439,N_4088,N_1627);
and U9440 (N_9440,N_3543,N_4204);
or U9441 (N_9441,N_3173,N_3151);
and U9442 (N_9442,N_3019,N_4141);
or U9443 (N_9443,N_3227,N_4008);
or U9444 (N_9444,N_2715,N_334);
and U9445 (N_9445,N_3642,N_4970);
xnor U9446 (N_9446,N_161,N_4294);
xor U9447 (N_9447,N_3929,N_1562);
xnor U9448 (N_9448,N_992,N_2052);
and U9449 (N_9449,N_4886,N_2816);
xor U9450 (N_9450,N_1599,N_1483);
nand U9451 (N_9451,N_557,N_731);
xor U9452 (N_9452,N_3557,N_2228);
nand U9453 (N_9453,N_4370,N_4541);
and U9454 (N_9454,N_4677,N_4694);
xnor U9455 (N_9455,N_259,N_4929);
nor U9456 (N_9456,N_1806,N_4668);
or U9457 (N_9457,N_535,N_367);
nor U9458 (N_9458,N_4225,N_494);
nand U9459 (N_9459,N_1068,N_595);
nor U9460 (N_9460,N_4814,N_1699);
and U9461 (N_9461,N_2010,N_4470);
nand U9462 (N_9462,N_4467,N_3850);
xnor U9463 (N_9463,N_503,N_3026);
xnor U9464 (N_9464,N_2977,N_533);
nand U9465 (N_9465,N_2868,N_1129);
nand U9466 (N_9466,N_3086,N_2465);
and U9467 (N_9467,N_1951,N_1077);
and U9468 (N_9468,N_4185,N_3285);
or U9469 (N_9469,N_2221,N_2590);
and U9470 (N_9470,N_4976,N_524);
nor U9471 (N_9471,N_374,N_492);
or U9472 (N_9472,N_4811,N_379);
nand U9473 (N_9473,N_2245,N_2230);
or U9474 (N_9474,N_2772,N_2982);
nand U9475 (N_9475,N_1121,N_3399);
or U9476 (N_9476,N_4546,N_4250);
and U9477 (N_9477,N_1449,N_2549);
or U9478 (N_9478,N_330,N_141);
nand U9479 (N_9479,N_730,N_287);
xnor U9480 (N_9480,N_17,N_4366);
nor U9481 (N_9481,N_1576,N_1936);
xor U9482 (N_9482,N_403,N_830);
and U9483 (N_9483,N_1183,N_1872);
and U9484 (N_9484,N_4861,N_3949);
or U9485 (N_9485,N_1830,N_1877);
and U9486 (N_9486,N_4599,N_239);
and U9487 (N_9487,N_645,N_1007);
and U9488 (N_9488,N_2582,N_2983);
or U9489 (N_9489,N_2202,N_1137);
or U9490 (N_9490,N_177,N_2708);
nand U9491 (N_9491,N_4285,N_2585);
nor U9492 (N_9492,N_2215,N_2260);
and U9493 (N_9493,N_716,N_1343);
nand U9494 (N_9494,N_1812,N_3934);
and U9495 (N_9495,N_4043,N_2562);
nand U9496 (N_9496,N_2935,N_287);
or U9497 (N_9497,N_1828,N_2575);
nand U9498 (N_9498,N_4351,N_2697);
xor U9499 (N_9499,N_4364,N_3151);
or U9500 (N_9500,N_4649,N_4450);
xnor U9501 (N_9501,N_1153,N_2097);
nand U9502 (N_9502,N_1698,N_1296);
or U9503 (N_9503,N_4786,N_551);
and U9504 (N_9504,N_1719,N_1601);
and U9505 (N_9505,N_800,N_4115);
nand U9506 (N_9506,N_1303,N_1125);
or U9507 (N_9507,N_622,N_2407);
nor U9508 (N_9508,N_4563,N_3600);
xor U9509 (N_9509,N_822,N_3021);
xor U9510 (N_9510,N_999,N_3708);
xor U9511 (N_9511,N_4547,N_4136);
and U9512 (N_9512,N_4513,N_1193);
nor U9513 (N_9513,N_2658,N_626);
xor U9514 (N_9514,N_4480,N_3791);
xnor U9515 (N_9515,N_2479,N_4125);
nand U9516 (N_9516,N_2643,N_2397);
nor U9517 (N_9517,N_4924,N_3814);
xnor U9518 (N_9518,N_858,N_3537);
nor U9519 (N_9519,N_1650,N_443);
nor U9520 (N_9520,N_1950,N_355);
nor U9521 (N_9521,N_3816,N_679);
xor U9522 (N_9522,N_2741,N_3035);
or U9523 (N_9523,N_3400,N_1504);
and U9524 (N_9524,N_607,N_2249);
or U9525 (N_9525,N_396,N_1041);
xor U9526 (N_9526,N_252,N_883);
nor U9527 (N_9527,N_4301,N_1269);
or U9528 (N_9528,N_2329,N_2044);
and U9529 (N_9529,N_2987,N_1504);
nor U9530 (N_9530,N_3209,N_1188);
xnor U9531 (N_9531,N_3360,N_4602);
and U9532 (N_9532,N_4964,N_3296);
and U9533 (N_9533,N_2293,N_2514);
xnor U9534 (N_9534,N_2601,N_567);
nor U9535 (N_9535,N_1268,N_892);
nand U9536 (N_9536,N_1015,N_2373);
nor U9537 (N_9537,N_2715,N_1402);
or U9538 (N_9538,N_2472,N_1333);
nand U9539 (N_9539,N_2128,N_3917);
nand U9540 (N_9540,N_987,N_1010);
or U9541 (N_9541,N_4576,N_1048);
and U9542 (N_9542,N_2348,N_2616);
xor U9543 (N_9543,N_1909,N_2590);
and U9544 (N_9544,N_1560,N_804);
nand U9545 (N_9545,N_1764,N_1547);
xnor U9546 (N_9546,N_1640,N_877);
xor U9547 (N_9547,N_329,N_708);
nor U9548 (N_9548,N_2461,N_2310);
and U9549 (N_9549,N_745,N_4316);
xnor U9550 (N_9550,N_3229,N_655);
xor U9551 (N_9551,N_3448,N_3257);
or U9552 (N_9552,N_2242,N_4195);
nor U9553 (N_9553,N_2693,N_4525);
and U9554 (N_9554,N_2521,N_2267);
xnor U9555 (N_9555,N_2414,N_329);
nand U9556 (N_9556,N_2242,N_1502);
and U9557 (N_9557,N_1389,N_2363);
or U9558 (N_9558,N_878,N_3181);
nor U9559 (N_9559,N_1533,N_4654);
and U9560 (N_9560,N_2512,N_1482);
and U9561 (N_9561,N_519,N_1767);
nand U9562 (N_9562,N_2512,N_3200);
nand U9563 (N_9563,N_2573,N_1177);
nor U9564 (N_9564,N_665,N_630);
and U9565 (N_9565,N_3684,N_2943);
or U9566 (N_9566,N_2664,N_2352);
xor U9567 (N_9567,N_1462,N_1482);
xnor U9568 (N_9568,N_4474,N_2323);
or U9569 (N_9569,N_3221,N_1807);
xor U9570 (N_9570,N_3868,N_1361);
and U9571 (N_9571,N_2998,N_3470);
nor U9572 (N_9572,N_2686,N_927);
xor U9573 (N_9573,N_184,N_14);
nor U9574 (N_9574,N_1827,N_772);
nand U9575 (N_9575,N_3545,N_4208);
nor U9576 (N_9576,N_1948,N_2960);
nor U9577 (N_9577,N_3809,N_2567);
nand U9578 (N_9578,N_3034,N_2042);
or U9579 (N_9579,N_3494,N_1045);
xnor U9580 (N_9580,N_3820,N_1500);
xnor U9581 (N_9581,N_1090,N_2788);
and U9582 (N_9582,N_1776,N_1882);
nor U9583 (N_9583,N_4773,N_406);
or U9584 (N_9584,N_3502,N_1146);
nor U9585 (N_9585,N_1068,N_263);
or U9586 (N_9586,N_2857,N_2580);
nand U9587 (N_9587,N_2527,N_2418);
and U9588 (N_9588,N_1865,N_4639);
or U9589 (N_9589,N_4248,N_3560);
nand U9590 (N_9590,N_2395,N_1154);
or U9591 (N_9591,N_1047,N_1178);
nand U9592 (N_9592,N_1264,N_4894);
or U9593 (N_9593,N_402,N_3298);
nor U9594 (N_9594,N_549,N_1174);
xnor U9595 (N_9595,N_523,N_3389);
xnor U9596 (N_9596,N_4652,N_4138);
or U9597 (N_9597,N_704,N_1736);
nor U9598 (N_9598,N_3287,N_2781);
or U9599 (N_9599,N_59,N_4349);
xor U9600 (N_9600,N_913,N_2351);
nor U9601 (N_9601,N_1814,N_2337);
nand U9602 (N_9602,N_3321,N_1162);
xnor U9603 (N_9603,N_917,N_4204);
xnor U9604 (N_9604,N_608,N_4468);
or U9605 (N_9605,N_998,N_4332);
or U9606 (N_9606,N_3832,N_4853);
xor U9607 (N_9607,N_1085,N_3165);
nor U9608 (N_9608,N_908,N_1315);
or U9609 (N_9609,N_2913,N_3719);
xor U9610 (N_9610,N_423,N_3907);
nor U9611 (N_9611,N_2636,N_690);
nor U9612 (N_9612,N_1559,N_3140);
and U9613 (N_9613,N_1773,N_1486);
nor U9614 (N_9614,N_1514,N_3594);
nor U9615 (N_9615,N_32,N_3950);
xor U9616 (N_9616,N_2517,N_4445);
xor U9617 (N_9617,N_3934,N_2242);
nor U9618 (N_9618,N_804,N_3586);
nor U9619 (N_9619,N_3801,N_295);
and U9620 (N_9620,N_2789,N_4167);
or U9621 (N_9621,N_3736,N_3258);
and U9622 (N_9622,N_3283,N_1916);
nor U9623 (N_9623,N_4529,N_3723);
or U9624 (N_9624,N_4035,N_4977);
or U9625 (N_9625,N_3279,N_2526);
nor U9626 (N_9626,N_4823,N_2991);
nand U9627 (N_9627,N_2471,N_429);
xnor U9628 (N_9628,N_3876,N_4052);
nor U9629 (N_9629,N_4927,N_553);
or U9630 (N_9630,N_4385,N_3096);
and U9631 (N_9631,N_1270,N_2243);
or U9632 (N_9632,N_3206,N_875);
and U9633 (N_9633,N_1647,N_2835);
nand U9634 (N_9634,N_3476,N_2114);
nand U9635 (N_9635,N_4282,N_4637);
and U9636 (N_9636,N_3048,N_4910);
xnor U9637 (N_9637,N_222,N_1838);
nor U9638 (N_9638,N_4725,N_1728);
nand U9639 (N_9639,N_3900,N_2835);
xor U9640 (N_9640,N_824,N_4835);
nand U9641 (N_9641,N_4820,N_94);
nor U9642 (N_9642,N_1055,N_2972);
and U9643 (N_9643,N_4359,N_4023);
nand U9644 (N_9644,N_682,N_1787);
nor U9645 (N_9645,N_295,N_3602);
nor U9646 (N_9646,N_2694,N_2389);
nor U9647 (N_9647,N_2610,N_441);
nor U9648 (N_9648,N_3228,N_2042);
or U9649 (N_9649,N_465,N_1727);
or U9650 (N_9650,N_3697,N_2871);
or U9651 (N_9651,N_4421,N_853);
nand U9652 (N_9652,N_3892,N_3425);
nand U9653 (N_9653,N_3804,N_4506);
nor U9654 (N_9654,N_420,N_249);
xor U9655 (N_9655,N_2842,N_3128);
nand U9656 (N_9656,N_3287,N_4342);
nor U9657 (N_9657,N_2886,N_1574);
or U9658 (N_9658,N_264,N_2849);
and U9659 (N_9659,N_4745,N_1558);
nand U9660 (N_9660,N_620,N_1196);
nor U9661 (N_9661,N_732,N_1071);
nor U9662 (N_9662,N_4398,N_4301);
nor U9663 (N_9663,N_1525,N_4709);
nor U9664 (N_9664,N_1333,N_1756);
and U9665 (N_9665,N_4007,N_423);
nor U9666 (N_9666,N_3872,N_1817);
or U9667 (N_9667,N_958,N_2682);
nand U9668 (N_9668,N_1724,N_937);
nor U9669 (N_9669,N_4579,N_3589);
or U9670 (N_9670,N_1415,N_4715);
nand U9671 (N_9671,N_2476,N_2449);
nand U9672 (N_9672,N_3855,N_1182);
nor U9673 (N_9673,N_1114,N_3024);
xor U9674 (N_9674,N_3010,N_4667);
and U9675 (N_9675,N_4948,N_2011);
nor U9676 (N_9676,N_1375,N_673);
nor U9677 (N_9677,N_3602,N_367);
or U9678 (N_9678,N_677,N_1436);
and U9679 (N_9679,N_1433,N_3539);
nand U9680 (N_9680,N_1180,N_4870);
and U9681 (N_9681,N_2436,N_4768);
or U9682 (N_9682,N_2655,N_1099);
xor U9683 (N_9683,N_906,N_4014);
and U9684 (N_9684,N_3967,N_1472);
xnor U9685 (N_9685,N_1379,N_3905);
and U9686 (N_9686,N_1409,N_3763);
and U9687 (N_9687,N_1879,N_1124);
nor U9688 (N_9688,N_4868,N_2087);
nand U9689 (N_9689,N_3946,N_676);
and U9690 (N_9690,N_2048,N_3895);
nand U9691 (N_9691,N_3899,N_512);
nand U9692 (N_9692,N_448,N_2960);
nor U9693 (N_9693,N_4195,N_1119);
xor U9694 (N_9694,N_4112,N_1056);
nor U9695 (N_9695,N_1511,N_2714);
and U9696 (N_9696,N_3891,N_1417);
nor U9697 (N_9697,N_297,N_4292);
or U9698 (N_9698,N_4681,N_701);
xor U9699 (N_9699,N_3297,N_789);
nand U9700 (N_9700,N_4975,N_3827);
xor U9701 (N_9701,N_539,N_1819);
nand U9702 (N_9702,N_1716,N_1776);
or U9703 (N_9703,N_1900,N_1761);
nor U9704 (N_9704,N_4358,N_1353);
nor U9705 (N_9705,N_1374,N_1711);
nand U9706 (N_9706,N_237,N_2462);
and U9707 (N_9707,N_627,N_2533);
nand U9708 (N_9708,N_836,N_1723);
xnor U9709 (N_9709,N_1658,N_4438);
and U9710 (N_9710,N_4969,N_3545);
nor U9711 (N_9711,N_1112,N_3872);
nor U9712 (N_9712,N_1242,N_1837);
xnor U9713 (N_9713,N_3794,N_519);
xnor U9714 (N_9714,N_2002,N_2013);
and U9715 (N_9715,N_3178,N_2827);
or U9716 (N_9716,N_1714,N_1356);
nand U9717 (N_9717,N_1594,N_1720);
and U9718 (N_9718,N_2497,N_2166);
and U9719 (N_9719,N_2638,N_4796);
and U9720 (N_9720,N_2928,N_3954);
xnor U9721 (N_9721,N_3169,N_4020);
nand U9722 (N_9722,N_2370,N_4942);
or U9723 (N_9723,N_2318,N_2093);
and U9724 (N_9724,N_2887,N_311);
nor U9725 (N_9725,N_77,N_3323);
or U9726 (N_9726,N_305,N_2060);
xor U9727 (N_9727,N_142,N_3076);
and U9728 (N_9728,N_4906,N_31);
and U9729 (N_9729,N_3620,N_3374);
or U9730 (N_9730,N_4136,N_2301);
nor U9731 (N_9731,N_1870,N_3886);
or U9732 (N_9732,N_1522,N_3624);
and U9733 (N_9733,N_3811,N_4722);
nand U9734 (N_9734,N_1344,N_2351);
xor U9735 (N_9735,N_4700,N_4565);
xor U9736 (N_9736,N_1854,N_3798);
nand U9737 (N_9737,N_1720,N_4783);
and U9738 (N_9738,N_2490,N_1073);
or U9739 (N_9739,N_773,N_2094);
or U9740 (N_9740,N_2932,N_742);
xnor U9741 (N_9741,N_3806,N_4090);
nor U9742 (N_9742,N_577,N_2759);
nand U9743 (N_9743,N_2589,N_1372);
nor U9744 (N_9744,N_3569,N_4212);
xnor U9745 (N_9745,N_4730,N_246);
nor U9746 (N_9746,N_2521,N_2764);
xor U9747 (N_9747,N_2929,N_1283);
xnor U9748 (N_9748,N_3714,N_2033);
or U9749 (N_9749,N_4116,N_2020);
or U9750 (N_9750,N_4782,N_2582);
nand U9751 (N_9751,N_146,N_3240);
xnor U9752 (N_9752,N_2236,N_4515);
and U9753 (N_9753,N_4065,N_1082);
or U9754 (N_9754,N_4413,N_4482);
nor U9755 (N_9755,N_2914,N_291);
and U9756 (N_9756,N_3964,N_404);
or U9757 (N_9757,N_1861,N_2742);
and U9758 (N_9758,N_4333,N_34);
xor U9759 (N_9759,N_4393,N_89);
and U9760 (N_9760,N_1073,N_1288);
and U9761 (N_9761,N_3783,N_1355);
nand U9762 (N_9762,N_3248,N_808);
nand U9763 (N_9763,N_2456,N_2747);
nor U9764 (N_9764,N_3062,N_2731);
nor U9765 (N_9765,N_4017,N_1398);
nor U9766 (N_9766,N_896,N_3078);
xor U9767 (N_9767,N_4333,N_4717);
nor U9768 (N_9768,N_1404,N_430);
nand U9769 (N_9769,N_3792,N_1136);
nor U9770 (N_9770,N_652,N_1204);
xnor U9771 (N_9771,N_2279,N_2855);
and U9772 (N_9772,N_3477,N_2535);
xnor U9773 (N_9773,N_1880,N_3904);
nor U9774 (N_9774,N_3579,N_1398);
or U9775 (N_9775,N_799,N_2142);
nor U9776 (N_9776,N_4917,N_4051);
nor U9777 (N_9777,N_754,N_54);
and U9778 (N_9778,N_2089,N_1200);
and U9779 (N_9779,N_2317,N_3358);
nor U9780 (N_9780,N_1067,N_638);
xor U9781 (N_9781,N_3051,N_4506);
nand U9782 (N_9782,N_1166,N_1599);
nor U9783 (N_9783,N_197,N_3379);
or U9784 (N_9784,N_2947,N_122);
and U9785 (N_9785,N_1621,N_4679);
nor U9786 (N_9786,N_2896,N_4879);
or U9787 (N_9787,N_2519,N_906);
or U9788 (N_9788,N_4242,N_1546);
nand U9789 (N_9789,N_3072,N_887);
nand U9790 (N_9790,N_2228,N_2521);
xor U9791 (N_9791,N_4466,N_2366);
nand U9792 (N_9792,N_1718,N_1318);
nand U9793 (N_9793,N_539,N_2181);
nand U9794 (N_9794,N_1025,N_4122);
and U9795 (N_9795,N_1345,N_665);
xnor U9796 (N_9796,N_224,N_2684);
xnor U9797 (N_9797,N_762,N_468);
nor U9798 (N_9798,N_1366,N_4);
or U9799 (N_9799,N_57,N_2884);
nand U9800 (N_9800,N_2867,N_299);
and U9801 (N_9801,N_1233,N_469);
nand U9802 (N_9802,N_3015,N_3793);
and U9803 (N_9803,N_3981,N_2987);
and U9804 (N_9804,N_3453,N_2865);
xor U9805 (N_9805,N_2433,N_1323);
nand U9806 (N_9806,N_3104,N_1724);
nor U9807 (N_9807,N_3596,N_2378);
nand U9808 (N_9808,N_9,N_1383);
and U9809 (N_9809,N_1950,N_1131);
or U9810 (N_9810,N_2212,N_1547);
and U9811 (N_9811,N_1483,N_2458);
and U9812 (N_9812,N_930,N_1061);
or U9813 (N_9813,N_4610,N_563);
or U9814 (N_9814,N_2448,N_1077);
nor U9815 (N_9815,N_4391,N_2639);
xnor U9816 (N_9816,N_4039,N_2938);
and U9817 (N_9817,N_3605,N_4506);
and U9818 (N_9818,N_2649,N_3411);
or U9819 (N_9819,N_1222,N_3302);
nand U9820 (N_9820,N_4341,N_4464);
nor U9821 (N_9821,N_4771,N_549);
or U9822 (N_9822,N_822,N_3672);
or U9823 (N_9823,N_728,N_2014);
xor U9824 (N_9824,N_1003,N_311);
nor U9825 (N_9825,N_2759,N_2794);
nand U9826 (N_9826,N_960,N_3216);
xnor U9827 (N_9827,N_1234,N_1120);
nor U9828 (N_9828,N_3249,N_381);
nor U9829 (N_9829,N_4211,N_1147);
and U9830 (N_9830,N_3400,N_1486);
nor U9831 (N_9831,N_1693,N_4430);
xnor U9832 (N_9832,N_2458,N_4123);
nor U9833 (N_9833,N_1268,N_211);
nand U9834 (N_9834,N_196,N_4207);
or U9835 (N_9835,N_4887,N_3457);
and U9836 (N_9836,N_3641,N_4127);
and U9837 (N_9837,N_1306,N_4368);
nor U9838 (N_9838,N_4122,N_4275);
and U9839 (N_9839,N_4878,N_3274);
or U9840 (N_9840,N_123,N_1164);
and U9841 (N_9841,N_3806,N_3345);
and U9842 (N_9842,N_4789,N_4507);
or U9843 (N_9843,N_4831,N_2799);
nand U9844 (N_9844,N_3799,N_4367);
xnor U9845 (N_9845,N_3774,N_2841);
xnor U9846 (N_9846,N_1098,N_3511);
nor U9847 (N_9847,N_3244,N_3574);
xnor U9848 (N_9848,N_1999,N_671);
nor U9849 (N_9849,N_2791,N_3313);
xnor U9850 (N_9850,N_1642,N_4628);
xor U9851 (N_9851,N_3946,N_3616);
and U9852 (N_9852,N_4237,N_1011);
xor U9853 (N_9853,N_4076,N_1398);
xor U9854 (N_9854,N_848,N_3209);
nor U9855 (N_9855,N_4069,N_1634);
nand U9856 (N_9856,N_3705,N_1271);
nand U9857 (N_9857,N_1153,N_3713);
nand U9858 (N_9858,N_953,N_1538);
and U9859 (N_9859,N_3156,N_86);
and U9860 (N_9860,N_1263,N_2361);
nand U9861 (N_9861,N_4277,N_4230);
nor U9862 (N_9862,N_4930,N_4118);
xor U9863 (N_9863,N_4146,N_3012);
nand U9864 (N_9864,N_2712,N_3232);
xnor U9865 (N_9865,N_2037,N_619);
nand U9866 (N_9866,N_331,N_3873);
and U9867 (N_9867,N_2310,N_1182);
nand U9868 (N_9868,N_143,N_4782);
xnor U9869 (N_9869,N_1508,N_2814);
xor U9870 (N_9870,N_4625,N_1323);
xnor U9871 (N_9871,N_3772,N_1395);
or U9872 (N_9872,N_4231,N_4190);
nand U9873 (N_9873,N_1373,N_1681);
xor U9874 (N_9874,N_1520,N_513);
and U9875 (N_9875,N_1428,N_234);
nand U9876 (N_9876,N_836,N_1323);
or U9877 (N_9877,N_348,N_1610);
and U9878 (N_9878,N_2314,N_4721);
or U9879 (N_9879,N_1812,N_989);
nor U9880 (N_9880,N_3902,N_3928);
xnor U9881 (N_9881,N_2185,N_2081);
or U9882 (N_9882,N_887,N_2169);
and U9883 (N_9883,N_2001,N_3036);
nor U9884 (N_9884,N_435,N_4866);
and U9885 (N_9885,N_529,N_1391);
nor U9886 (N_9886,N_2375,N_726);
xnor U9887 (N_9887,N_4330,N_3344);
and U9888 (N_9888,N_4743,N_2409);
or U9889 (N_9889,N_3604,N_130);
xnor U9890 (N_9890,N_4464,N_2720);
and U9891 (N_9891,N_3397,N_1392);
nor U9892 (N_9892,N_1077,N_1977);
and U9893 (N_9893,N_3752,N_937);
nand U9894 (N_9894,N_3777,N_1713);
xnor U9895 (N_9895,N_2509,N_2621);
and U9896 (N_9896,N_1081,N_661);
and U9897 (N_9897,N_1696,N_3080);
or U9898 (N_9898,N_3870,N_2402);
nor U9899 (N_9899,N_2897,N_4500);
or U9900 (N_9900,N_2277,N_1264);
or U9901 (N_9901,N_3590,N_1398);
xor U9902 (N_9902,N_3614,N_1933);
and U9903 (N_9903,N_2000,N_3847);
xnor U9904 (N_9904,N_1301,N_1201);
nand U9905 (N_9905,N_2856,N_921);
nand U9906 (N_9906,N_2679,N_2866);
nand U9907 (N_9907,N_304,N_187);
xnor U9908 (N_9908,N_1051,N_2451);
nand U9909 (N_9909,N_566,N_1857);
xor U9910 (N_9910,N_1689,N_3107);
nand U9911 (N_9911,N_1754,N_1464);
xnor U9912 (N_9912,N_1672,N_3554);
and U9913 (N_9913,N_915,N_2518);
nor U9914 (N_9914,N_141,N_4490);
nand U9915 (N_9915,N_1504,N_1380);
and U9916 (N_9916,N_4827,N_894);
and U9917 (N_9917,N_3993,N_4160);
xor U9918 (N_9918,N_4700,N_1854);
and U9919 (N_9919,N_4337,N_1659);
and U9920 (N_9920,N_552,N_1039);
and U9921 (N_9921,N_757,N_3527);
or U9922 (N_9922,N_2579,N_1658);
nor U9923 (N_9923,N_694,N_2522);
or U9924 (N_9924,N_4254,N_3272);
nor U9925 (N_9925,N_2482,N_882);
or U9926 (N_9926,N_3363,N_1702);
nand U9927 (N_9927,N_342,N_3633);
and U9928 (N_9928,N_3004,N_3862);
xnor U9929 (N_9929,N_1753,N_67);
nor U9930 (N_9930,N_2413,N_114);
or U9931 (N_9931,N_2764,N_1856);
nor U9932 (N_9932,N_1660,N_4381);
xor U9933 (N_9933,N_4755,N_2650);
or U9934 (N_9934,N_3122,N_1757);
xor U9935 (N_9935,N_1225,N_1443);
nand U9936 (N_9936,N_49,N_3024);
and U9937 (N_9937,N_2407,N_3821);
or U9938 (N_9938,N_667,N_655);
nor U9939 (N_9939,N_4543,N_2367);
nand U9940 (N_9940,N_2991,N_1736);
xnor U9941 (N_9941,N_1522,N_2068);
nand U9942 (N_9942,N_783,N_3764);
and U9943 (N_9943,N_2327,N_1918);
xor U9944 (N_9944,N_653,N_2263);
or U9945 (N_9945,N_2284,N_3332);
xor U9946 (N_9946,N_3445,N_337);
nor U9947 (N_9947,N_2410,N_1020);
or U9948 (N_9948,N_3640,N_790);
and U9949 (N_9949,N_3835,N_4080);
or U9950 (N_9950,N_228,N_1985);
nor U9951 (N_9951,N_1915,N_2179);
nor U9952 (N_9952,N_52,N_3449);
nor U9953 (N_9953,N_728,N_3834);
nand U9954 (N_9954,N_125,N_4218);
nor U9955 (N_9955,N_4368,N_462);
xor U9956 (N_9956,N_313,N_4718);
xor U9957 (N_9957,N_4111,N_4431);
nor U9958 (N_9958,N_2831,N_3421);
nand U9959 (N_9959,N_4510,N_4492);
nor U9960 (N_9960,N_405,N_3926);
nand U9961 (N_9961,N_177,N_33);
and U9962 (N_9962,N_3015,N_413);
nand U9963 (N_9963,N_1016,N_4327);
nor U9964 (N_9964,N_2396,N_4655);
nor U9965 (N_9965,N_3196,N_1459);
or U9966 (N_9966,N_422,N_881);
nand U9967 (N_9967,N_582,N_1533);
nand U9968 (N_9968,N_11,N_431);
nor U9969 (N_9969,N_4099,N_294);
xnor U9970 (N_9970,N_894,N_2785);
or U9971 (N_9971,N_4768,N_87);
or U9972 (N_9972,N_767,N_425);
and U9973 (N_9973,N_731,N_1263);
and U9974 (N_9974,N_2732,N_877);
nand U9975 (N_9975,N_1032,N_1723);
nand U9976 (N_9976,N_2383,N_2369);
nand U9977 (N_9977,N_723,N_3300);
xor U9978 (N_9978,N_1331,N_1837);
or U9979 (N_9979,N_4793,N_3485);
or U9980 (N_9980,N_1422,N_1395);
xor U9981 (N_9981,N_3231,N_1443);
nand U9982 (N_9982,N_2222,N_3593);
nand U9983 (N_9983,N_499,N_2135);
nor U9984 (N_9984,N_1519,N_373);
nand U9985 (N_9985,N_3916,N_1957);
nand U9986 (N_9986,N_3413,N_238);
xor U9987 (N_9987,N_2519,N_2253);
or U9988 (N_9988,N_1883,N_3511);
or U9989 (N_9989,N_3322,N_2127);
and U9990 (N_9990,N_3666,N_4268);
nor U9991 (N_9991,N_4211,N_826);
xnor U9992 (N_9992,N_129,N_977);
xnor U9993 (N_9993,N_3872,N_1551);
xnor U9994 (N_9994,N_2125,N_4580);
and U9995 (N_9995,N_4172,N_969);
nand U9996 (N_9996,N_3353,N_3512);
and U9997 (N_9997,N_3525,N_4864);
nor U9998 (N_9998,N_2250,N_4580);
nand U9999 (N_9999,N_2354,N_367);
or U10000 (N_10000,N_6217,N_5886);
xnor U10001 (N_10001,N_5664,N_5024);
nand U10002 (N_10002,N_6152,N_8595);
nor U10003 (N_10003,N_7808,N_8708);
nor U10004 (N_10004,N_9253,N_7506);
and U10005 (N_10005,N_6768,N_8117);
xor U10006 (N_10006,N_6443,N_6434);
xnor U10007 (N_10007,N_6765,N_5410);
and U10008 (N_10008,N_8724,N_9610);
and U10009 (N_10009,N_8444,N_7796);
or U10010 (N_10010,N_7565,N_5123);
and U10011 (N_10011,N_9095,N_6780);
and U10012 (N_10012,N_6947,N_7539);
nor U10013 (N_10013,N_6690,N_5184);
and U10014 (N_10014,N_7508,N_6719);
nand U10015 (N_10015,N_5057,N_6772);
nand U10016 (N_10016,N_9763,N_7676);
nand U10017 (N_10017,N_6148,N_7838);
or U10018 (N_10018,N_6923,N_7147);
or U10019 (N_10019,N_5264,N_8493);
xnor U10020 (N_10020,N_9984,N_6352);
and U10021 (N_10021,N_6831,N_5370);
nand U10022 (N_10022,N_7721,N_5812);
nand U10023 (N_10023,N_8120,N_9276);
or U10024 (N_10024,N_7278,N_6094);
nor U10025 (N_10025,N_7964,N_8409);
and U10026 (N_10026,N_8950,N_8695);
nand U10027 (N_10027,N_9089,N_5549);
nor U10028 (N_10028,N_9171,N_8810);
and U10029 (N_10029,N_8463,N_5963);
nor U10030 (N_10030,N_6431,N_5400);
nor U10031 (N_10031,N_6079,N_6065);
and U10032 (N_10032,N_6536,N_8496);
and U10033 (N_10033,N_6648,N_5780);
or U10034 (N_10034,N_9373,N_7321);
and U10035 (N_10035,N_8947,N_7834);
xnor U10036 (N_10036,N_7849,N_9492);
nor U10037 (N_10037,N_6547,N_7000);
nor U10038 (N_10038,N_8566,N_9819);
xor U10039 (N_10039,N_5778,N_7449);
and U10040 (N_10040,N_6789,N_9474);
and U10041 (N_10041,N_9219,N_8282);
and U10042 (N_10042,N_5904,N_8725);
nor U10043 (N_10043,N_5501,N_5276);
and U10044 (N_10044,N_7988,N_8435);
or U10045 (N_10045,N_5872,N_5883);
xnor U10046 (N_10046,N_6658,N_5471);
xnor U10047 (N_10047,N_5649,N_5205);
nand U10048 (N_10048,N_7741,N_6977);
nor U10049 (N_10049,N_6940,N_7687);
nand U10050 (N_10050,N_5039,N_6819);
xor U10051 (N_10051,N_9488,N_9187);
nor U10052 (N_10052,N_7400,N_5532);
nand U10053 (N_10053,N_5573,N_5455);
or U10054 (N_10054,N_7525,N_7653);
nor U10055 (N_10055,N_7727,N_7107);
xnor U10056 (N_10056,N_6852,N_8430);
or U10057 (N_10057,N_8327,N_5157);
and U10058 (N_10058,N_9047,N_5199);
xor U10059 (N_10059,N_5879,N_7415);
nand U10060 (N_10060,N_8143,N_8255);
xor U10061 (N_10061,N_8349,N_7809);
xnor U10062 (N_10062,N_8307,N_9658);
xor U10063 (N_10063,N_9490,N_5959);
nand U10064 (N_10064,N_5472,N_9486);
nand U10065 (N_10065,N_6861,N_9558);
nor U10066 (N_10066,N_6716,N_7077);
nor U10067 (N_10067,N_9156,N_8302);
or U10068 (N_10068,N_5875,N_8765);
and U10069 (N_10069,N_7122,N_5957);
nor U10070 (N_10070,N_5418,N_6311);
xnor U10071 (N_10071,N_5226,N_7357);
nand U10072 (N_10072,N_6890,N_7833);
or U10073 (N_10073,N_6614,N_5245);
and U10074 (N_10074,N_6145,N_7324);
nor U10075 (N_10075,N_8420,N_7876);
xnor U10076 (N_10076,N_6291,N_8919);
and U10077 (N_10077,N_5132,N_7337);
nor U10078 (N_10078,N_5838,N_7553);
xnor U10079 (N_10079,N_8626,N_9168);
or U10080 (N_10080,N_5653,N_9031);
xor U10081 (N_10081,N_6095,N_5151);
or U10082 (N_10082,N_5934,N_6885);
nor U10083 (N_10083,N_8070,N_9384);
xnor U10084 (N_10084,N_8123,N_9175);
nor U10085 (N_10085,N_6140,N_7125);
and U10086 (N_10086,N_9120,N_6709);
and U10087 (N_10087,N_7970,N_9519);
and U10088 (N_10088,N_6535,N_7794);
or U10089 (N_10089,N_9580,N_6720);
or U10090 (N_10090,N_9848,N_9107);
and U10091 (N_10091,N_9412,N_7662);
nand U10092 (N_10092,N_7161,N_5503);
xnor U10093 (N_10093,N_5775,N_9148);
nand U10094 (N_10094,N_5854,N_9515);
and U10095 (N_10095,N_8206,N_7825);
or U10096 (N_10096,N_6481,N_7936);
nor U10097 (N_10097,N_8107,N_5247);
xnor U10098 (N_10098,N_8581,N_9917);
nor U10099 (N_10099,N_5244,N_8477);
xnor U10100 (N_10100,N_9884,N_8543);
and U10101 (N_10101,N_8210,N_9046);
and U10102 (N_10102,N_9663,N_7552);
nand U10103 (N_10103,N_5861,N_9553);
or U10104 (N_10104,N_9740,N_9811);
and U10105 (N_10105,N_8715,N_9859);
and U10106 (N_10106,N_5273,N_8071);
nor U10107 (N_10107,N_6453,N_7291);
and U10108 (N_10108,N_6718,N_6181);
xnor U10109 (N_10109,N_7004,N_5774);
xor U10110 (N_10110,N_6042,N_8122);
xor U10111 (N_10111,N_6405,N_7047);
xor U10112 (N_10112,N_9590,N_9448);
or U10113 (N_10113,N_8601,N_7434);
or U10114 (N_10114,N_5386,N_9332);
or U10115 (N_10115,N_8663,N_8252);
nand U10116 (N_10116,N_9354,N_5624);
and U10117 (N_10117,N_6714,N_7590);
or U10118 (N_10118,N_9621,N_6240);
and U10119 (N_10119,N_8330,N_8610);
xor U10120 (N_10120,N_9616,N_8587);
xnor U10121 (N_10121,N_8850,N_9044);
or U10122 (N_10122,N_8099,N_5435);
nand U10123 (N_10123,N_8625,N_6823);
and U10124 (N_10124,N_9322,N_5166);
nand U10125 (N_10125,N_6342,N_5169);
xor U10126 (N_10126,N_9736,N_9505);
nor U10127 (N_10127,N_9647,N_7623);
xnor U10128 (N_10128,N_8548,N_5530);
nor U10129 (N_10129,N_6911,N_9323);
xor U10130 (N_10130,N_9682,N_9416);
nor U10131 (N_10131,N_9014,N_9636);
nor U10132 (N_10132,N_9678,N_6336);
nand U10133 (N_10133,N_5090,N_8369);
or U10134 (N_10134,N_9508,N_5328);
or U10135 (N_10135,N_8140,N_5253);
or U10136 (N_10136,N_6880,N_8966);
nand U10137 (N_10137,N_7061,N_7028);
nand U10138 (N_10138,N_7181,N_7287);
or U10139 (N_10139,N_6258,N_9121);
nand U10140 (N_10140,N_8905,N_8547);
nand U10141 (N_10141,N_7875,N_8711);
and U10142 (N_10142,N_7527,N_9063);
nor U10143 (N_10143,N_7356,N_9700);
nor U10144 (N_10144,N_7871,N_7220);
or U10145 (N_10145,N_6057,N_5927);
or U10146 (N_10146,N_8474,N_9079);
nor U10147 (N_10147,N_7955,N_6466);
and U10148 (N_10148,N_7615,N_6149);
xnor U10149 (N_10149,N_6440,N_8254);
nand U10150 (N_10150,N_6232,N_5806);
xnor U10151 (N_10151,N_9991,N_7010);
nand U10152 (N_10152,N_8332,N_7868);
xnor U10153 (N_10153,N_5951,N_6077);
and U10154 (N_10154,N_7725,N_5740);
and U10155 (N_10155,N_8333,N_5576);
or U10156 (N_10156,N_9988,N_6087);
nor U10157 (N_10157,N_7756,N_6397);
and U10158 (N_10158,N_9537,N_9411);
nand U10159 (N_10159,N_9229,N_6402);
and U10160 (N_10160,N_6040,N_8238);
nand U10161 (N_10161,N_5623,N_8819);
nand U10162 (N_10162,N_7632,N_9407);
xnor U10163 (N_10163,N_7027,N_9181);
nand U10164 (N_10164,N_8172,N_6340);
and U10165 (N_10165,N_7806,N_5525);
xnor U10166 (N_10166,N_9756,N_8778);
xor U10167 (N_10167,N_7561,N_7585);
xnor U10168 (N_10168,N_5495,N_9455);
nand U10169 (N_10169,N_9057,N_5187);
nand U10170 (N_10170,N_5545,N_5719);
or U10171 (N_10171,N_9345,N_8891);
or U10172 (N_10172,N_9949,N_5498);
or U10173 (N_10173,N_5294,N_9874);
and U10174 (N_10174,N_6015,N_7985);
xor U10175 (N_10175,N_6791,N_7394);
nand U10176 (N_10176,N_7782,N_6706);
nand U10177 (N_10177,N_5613,N_7219);
nand U10178 (N_10178,N_8898,N_9444);
nor U10179 (N_10179,N_8881,N_7389);
or U10180 (N_10180,N_7826,N_9165);
nor U10181 (N_10181,N_6213,N_9822);
nor U10182 (N_10182,N_8239,N_5869);
or U10183 (N_10183,N_5708,N_7895);
nor U10184 (N_10184,N_7041,N_8520);
nor U10185 (N_10185,N_6250,N_7087);
xnor U10186 (N_10186,N_9346,N_8736);
and U10187 (N_10187,N_6686,N_8467);
or U10188 (N_10188,N_7268,N_6632);
xnor U10189 (N_10189,N_5982,N_5104);
or U10190 (N_10190,N_7436,N_7385);
nor U10191 (N_10191,N_7478,N_6226);
xnor U10192 (N_10192,N_7339,N_7019);
nor U10193 (N_10193,N_6903,N_7989);
nor U10194 (N_10194,N_6111,N_6549);
nor U10195 (N_10195,N_5699,N_5426);
and U10196 (N_10196,N_5034,N_6119);
and U10197 (N_10197,N_9719,N_9995);
xnor U10198 (N_10198,N_9920,N_8714);
xnor U10199 (N_10199,N_5636,N_9023);
xnor U10200 (N_10200,N_6949,N_8552);
nor U10201 (N_10201,N_9234,N_7734);
or U10202 (N_10202,N_9645,N_6014);
or U10203 (N_10203,N_9653,N_6004);
nor U10204 (N_10204,N_5730,N_8145);
and U10205 (N_10205,N_8793,N_8777);
nor U10206 (N_10206,N_9711,N_8393);
and U10207 (N_10207,N_8789,N_5536);
and U10208 (N_10208,N_5047,N_6046);
nor U10209 (N_10209,N_5315,N_5960);
and U10210 (N_10210,N_7627,N_9240);
and U10211 (N_10211,N_5942,N_9003);
or U10212 (N_10212,N_5829,N_5288);
and U10213 (N_10213,N_5641,N_6538);
xor U10214 (N_10214,N_7953,N_7792);
nor U10215 (N_10215,N_5881,N_9464);
nor U10216 (N_10216,N_9366,N_8839);
nor U10217 (N_10217,N_6856,N_8506);
or U10218 (N_10218,N_8067,N_7154);
nand U10219 (N_10219,N_5021,N_6383);
nor U10220 (N_10220,N_5984,N_9997);
nand U10221 (N_10221,N_8365,N_7975);
or U10222 (N_10222,N_9237,N_9833);
and U10223 (N_10223,N_6221,N_9527);
or U10224 (N_10224,N_6518,N_7537);
and U10225 (N_10225,N_9461,N_6411);
nand U10226 (N_10226,N_9986,N_7821);
or U10227 (N_10227,N_9823,N_7246);
or U10228 (N_10228,N_6778,N_5896);
xnor U10229 (N_10229,N_9825,N_7702);
and U10230 (N_10230,N_9045,N_6272);
and U10231 (N_10231,N_5424,N_9115);
nor U10232 (N_10232,N_8923,N_7943);
xnor U10233 (N_10233,N_6552,N_8940);
or U10234 (N_10234,N_6787,N_8358);
xnor U10235 (N_10235,N_5857,N_8975);
nor U10236 (N_10236,N_9438,N_5973);
nor U10237 (N_10237,N_7418,N_5916);
nor U10238 (N_10238,N_6229,N_7250);
xor U10239 (N_10239,N_5692,N_9102);
xor U10240 (N_10240,N_8014,N_7766);
and U10241 (N_10241,N_5384,N_6030);
or U10242 (N_10242,N_7050,N_8065);
or U10243 (N_10243,N_6527,N_6700);
nand U10244 (N_10244,N_7018,N_8164);
or U10245 (N_10245,N_7365,N_5417);
nand U10246 (N_10246,N_8093,N_9659);
or U10247 (N_10247,N_5763,N_8622);
nor U10248 (N_10248,N_6051,N_9477);
nor U10249 (N_10249,N_9861,N_8591);
xor U10250 (N_10250,N_9729,N_7071);
or U10251 (N_10251,N_5652,N_5043);
or U10252 (N_10252,N_9992,N_9747);
xnor U10253 (N_10253,N_7267,N_5945);
or U10254 (N_10254,N_6052,N_7395);
and U10255 (N_10255,N_9744,N_9302);
or U10256 (N_10256,N_8804,N_9218);
or U10257 (N_10257,N_7424,N_5620);
xor U10258 (N_10258,N_5142,N_6764);
nor U10259 (N_10259,N_5178,N_8223);
and U10260 (N_10260,N_8539,N_6283);
nor U10261 (N_10261,N_6679,N_6888);
xor U10262 (N_10262,N_6587,N_8951);
or U10263 (N_10263,N_5075,N_9173);
nor U10264 (N_10264,N_5167,N_5372);
or U10265 (N_10265,N_6993,N_9252);
nand U10266 (N_10266,N_9491,N_5972);
and U10267 (N_10267,N_7701,N_6588);
and U10268 (N_10268,N_8931,N_7699);
nor U10269 (N_10269,N_8515,N_9794);
nand U10270 (N_10270,N_8750,N_5914);
xnor U10271 (N_10271,N_7240,N_9692);
or U10272 (N_10272,N_6252,N_9052);
nand U10273 (N_10273,N_6238,N_5000);
or U10274 (N_10274,N_8589,N_7105);
nor U10275 (N_10275,N_9158,N_6912);
nor U10276 (N_10276,N_6581,N_9755);
and U10277 (N_10277,N_7285,N_5326);
and U10278 (N_10278,N_5674,N_5818);
and U10279 (N_10279,N_8730,N_5746);
xor U10280 (N_10280,N_5804,N_6698);
and U10281 (N_10281,N_6950,N_9202);
or U10282 (N_10282,N_7578,N_9867);
nand U10283 (N_10283,N_7428,N_5967);
nor U10284 (N_10284,N_7990,N_9297);
or U10285 (N_10285,N_9803,N_9226);
nand U10286 (N_10286,N_5732,N_8323);
nor U10287 (N_10287,N_9907,N_9906);
nor U10288 (N_10288,N_5546,N_6623);
xor U10289 (N_10289,N_8885,N_6755);
xor U10290 (N_10290,N_6696,N_5461);
xor U10291 (N_10291,N_9029,N_5920);
nand U10292 (N_10292,N_5022,N_5792);
or U10293 (N_10293,N_6933,N_7996);
or U10294 (N_10294,N_7550,N_5462);
nor U10295 (N_10295,N_8036,N_7924);
xor U10296 (N_10296,N_5999,N_6884);
xor U10297 (N_10297,N_6743,N_9314);
or U10298 (N_10298,N_7425,N_9846);
or U10299 (N_10299,N_9881,N_8925);
nor U10300 (N_10300,N_9449,N_6757);
or U10301 (N_10301,N_6355,N_5440);
xor U10302 (N_10302,N_7800,N_7447);
nor U10303 (N_10303,N_6343,N_8655);
or U10304 (N_10304,N_9471,N_5599);
nand U10305 (N_10305,N_9405,N_7074);
xor U10306 (N_10306,N_9073,N_8263);
nor U10307 (N_10307,N_8003,N_5103);
xnor U10308 (N_10308,N_8759,N_6551);
and U10309 (N_10309,N_5617,N_5155);
nand U10310 (N_10310,N_5701,N_8703);
and U10311 (N_10311,N_5301,N_6384);
and U10312 (N_10312,N_5289,N_8376);
nor U10313 (N_10313,N_6670,N_7429);
nor U10314 (N_10314,N_8673,N_9716);
xor U10315 (N_10315,N_6260,N_7148);
nor U10316 (N_10316,N_6779,N_6132);
nand U10317 (N_10317,N_7034,N_5836);
nand U10318 (N_10318,N_6284,N_7313);
and U10319 (N_10319,N_5899,N_7597);
xor U10320 (N_10320,N_5607,N_5670);
nand U10321 (N_10321,N_9386,N_7190);
nor U10322 (N_10322,N_5516,N_6165);
nand U10323 (N_10323,N_9432,N_9064);
or U10324 (N_10324,N_7731,N_6444);
and U10325 (N_10325,N_9009,N_7788);
xnor U10326 (N_10326,N_7145,N_5600);
or U10327 (N_10327,N_6457,N_7006);
and U10328 (N_10328,N_5049,N_9726);
xnor U10329 (N_10329,N_5242,N_7974);
and U10330 (N_10330,N_8943,N_8222);
and U10331 (N_10331,N_6347,N_5824);
and U10332 (N_10332,N_5716,N_7375);
or U10333 (N_10333,N_5229,N_7214);
xor U10334 (N_10334,N_8586,N_6158);
or U10335 (N_10335,N_9257,N_9118);
nand U10336 (N_10336,N_8900,N_7149);
and U10337 (N_10337,N_7841,N_5221);
xor U10338 (N_10338,N_7801,N_8852);
nand U10339 (N_10339,N_5614,N_9761);
xnor U10340 (N_10340,N_8879,N_7070);
nor U10341 (N_10341,N_9315,N_6615);
nor U10342 (N_10342,N_7475,N_7118);
and U10343 (N_10343,N_5092,N_6295);
nor U10344 (N_10344,N_8912,N_5126);
nor U10345 (N_10345,N_6951,N_6338);
xnor U10346 (N_10346,N_8671,N_5482);
or U10347 (N_10347,N_5616,N_5611);
nor U10348 (N_10348,N_8760,N_7231);
or U10349 (N_10349,N_5630,N_9720);
nand U10350 (N_10350,N_6309,N_8380);
nand U10351 (N_10351,N_9520,N_9526);
or U10352 (N_10352,N_6506,N_7864);
and U10353 (N_10353,N_8362,N_7039);
nor U10354 (N_10354,N_8897,N_9143);
or U10355 (N_10355,N_7131,N_5723);
and U10356 (N_10356,N_6633,N_7563);
nand U10357 (N_10357,N_9512,N_9622);
nand U10358 (N_10358,N_8838,N_7830);
nand U10359 (N_10359,N_7515,N_7526);
nand U10360 (N_10360,N_8927,N_7319);
nand U10361 (N_10361,N_5353,N_6974);
or U10362 (N_10362,N_9087,N_7612);
nand U10363 (N_10363,N_8159,N_8536);
nor U10364 (N_10364,N_8614,N_6107);
or U10365 (N_10365,N_8871,N_5695);
or U10366 (N_10366,N_6178,N_8075);
nor U10367 (N_10367,N_9764,N_6450);
xnor U10368 (N_10368,N_8267,N_9836);
and U10369 (N_10369,N_6312,N_9938);
nor U10370 (N_10370,N_6177,N_8157);
nor U10371 (N_10371,N_5484,N_7616);
xor U10372 (N_10372,N_8105,N_7358);
or U10373 (N_10373,N_7491,N_5122);
or U10374 (N_10374,N_6223,N_9042);
nand U10375 (N_10375,N_8865,N_6195);
xor U10376 (N_10376,N_9518,N_5191);
or U10377 (N_10377,N_6275,N_6776);
nand U10378 (N_10378,N_8331,N_8205);
or U10379 (N_10379,N_9664,N_6096);
nor U10380 (N_10380,N_6900,N_7799);
and U10381 (N_10381,N_5281,N_8913);
xnor U10382 (N_10382,N_5394,N_7013);
nor U10383 (N_10383,N_6800,N_6729);
nand U10384 (N_10384,N_7300,N_9066);
xnor U10385 (N_10385,N_9094,N_5296);
xor U10386 (N_10386,N_5448,N_5598);
xor U10387 (N_10387,N_9177,N_7559);
or U10388 (N_10388,N_9383,N_5714);
nor U10389 (N_10389,N_6187,N_8144);
or U10390 (N_10390,N_5754,N_8841);
and U10391 (N_10391,N_7870,N_8475);
xor U10392 (N_10392,N_6973,N_9552);
nor U10393 (N_10393,N_8271,N_5031);
nand U10394 (N_10394,N_8005,N_6483);
nor U10395 (N_10395,N_7003,N_6608);
and U10396 (N_10396,N_5787,N_8337);
nand U10397 (N_10397,N_6786,N_6498);
xnor U10398 (N_10398,N_6832,N_7310);
and U10399 (N_10399,N_7958,N_6862);
or U10400 (N_10400,N_7062,N_5953);
and U10401 (N_10401,N_7560,N_5347);
and U10402 (N_10402,N_5206,N_6618);
and U10403 (N_10403,N_7682,N_9675);
xor U10404 (N_10404,N_9434,N_8173);
nor U10405 (N_10405,N_9262,N_6957);
nor U10406 (N_10406,N_8182,N_6490);
nand U10407 (N_10407,N_6013,N_7290);
xor U10408 (N_10408,N_6710,N_7896);
nor U10409 (N_10409,N_9280,N_5596);
xnor U10410 (N_10410,N_8104,N_8659);
or U10411 (N_10411,N_9810,N_5310);
xor U10412 (N_10412,N_8847,N_9399);
nor U10413 (N_10413,N_6211,N_7237);
and U10414 (N_10414,N_8377,N_9137);
nand U10415 (N_10415,N_7965,N_8867);
or U10416 (N_10416,N_6028,N_7775);
nor U10417 (N_10417,N_5766,N_6246);
and U10418 (N_10418,N_8260,N_9370);
nand U10419 (N_10419,N_8845,N_5805);
or U10420 (N_10420,N_9612,N_7298);
xor U10421 (N_10421,N_7655,N_8848);
and U10422 (N_10422,N_6839,N_5750);
nand U10423 (N_10423,N_6413,N_6108);
and U10424 (N_10424,N_9417,N_7818);
nor U10425 (N_10425,N_5592,N_7493);
nand U10426 (N_10426,N_7419,N_8575);
nor U10427 (N_10427,N_8690,N_9458);
nor U10428 (N_10428,N_8440,N_9556);
nand U10429 (N_10429,N_6674,N_8407);
nand U10430 (N_10430,N_7406,N_7150);
or U10431 (N_10431,N_5139,N_6027);
nor U10432 (N_10432,N_8322,N_6100);
nand U10433 (N_10433,N_5190,N_6917);
nor U10434 (N_10434,N_9032,N_9851);
nand U10435 (N_10435,N_8576,N_5124);
nand U10436 (N_10436,N_5068,N_5593);
nand U10437 (N_10437,N_7111,N_5208);
or U10438 (N_10438,N_8723,N_9531);
xnor U10439 (N_10439,N_5552,N_6846);
nand U10440 (N_10440,N_7348,N_8664);
nand U10441 (N_10441,N_7872,N_7866);
xor U10442 (N_10442,N_7922,N_6179);
and U10443 (N_10443,N_6356,N_7151);
or U10444 (N_10444,N_6896,N_6299);
and U10445 (N_10445,N_5001,N_9789);
or U10446 (N_10446,N_9286,N_5988);
or U10447 (N_10447,N_7384,N_8443);
nand U10448 (N_10448,N_5629,N_8480);
xnor U10449 (N_10449,N_7309,N_8541);
or U10450 (N_10450,N_9685,N_8957);
or U10451 (N_10451,N_7412,N_6889);
or U10452 (N_10452,N_6294,N_8113);
and U10453 (N_10453,N_5477,N_9422);
nor U10454 (N_10454,N_6146,N_9117);
nor U10455 (N_10455,N_8129,N_6688);
xor U10456 (N_10456,N_7017,N_6693);
or U10457 (N_10457,N_8518,N_9065);
nor U10458 (N_10458,N_7022,N_9186);
nor U10459 (N_10459,N_5578,N_9265);
nand U10460 (N_10460,N_9648,N_6886);
and U10461 (N_10461,N_8658,N_6978);
or U10462 (N_10462,N_8438,N_6242);
or U10463 (N_10463,N_7186,N_8218);
nand U10464 (N_10464,N_8230,N_7239);
xor U10465 (N_10465,N_6086,N_5094);
xor U10466 (N_10466,N_6388,N_6593);
or U10467 (N_10467,N_7855,N_5510);
and U10468 (N_10468,N_7551,N_5362);
xnor U10469 (N_10469,N_6834,N_5407);
xor U10470 (N_10470,N_9006,N_6321);
nand U10471 (N_10471,N_9796,N_7226);
nor U10472 (N_10472,N_5404,N_8992);
and U10473 (N_10473,N_8464,N_5496);
nand U10474 (N_10474,N_9958,N_9722);
or U10475 (N_10475,N_6577,N_7667);
xor U10476 (N_10476,N_6500,N_8886);
nand U10477 (N_10477,N_7199,N_6032);
or U10478 (N_10478,N_5538,N_9891);
xnor U10479 (N_10479,N_8651,N_6597);
xnor U10480 (N_10480,N_9221,N_6288);
xnor U10481 (N_10481,N_9116,N_5757);
or U10482 (N_10482,N_9456,N_9011);
nand U10483 (N_10483,N_6006,N_7314);
and U10484 (N_10484,N_6984,N_5375);
nor U10485 (N_10485,N_5688,N_9624);
and U10486 (N_10486,N_5232,N_7328);
xnor U10487 (N_10487,N_5314,N_9957);
nand U10488 (N_10488,N_5891,N_8818);
or U10489 (N_10489,N_7633,N_7410);
xnor U10490 (N_10490,N_8356,N_8195);
nand U10491 (N_10491,N_9813,N_7097);
and U10492 (N_10492,N_7557,N_9785);
and U10493 (N_10493,N_5131,N_8572);
nand U10494 (N_10494,N_6741,N_8784);
xnor U10495 (N_10495,N_9169,N_5282);
nor U10496 (N_10496,N_7863,N_5677);
nor U10497 (N_10497,N_6012,N_8007);
or U10498 (N_10498,N_7432,N_9206);
nand U10499 (N_10499,N_9254,N_6788);
or U10500 (N_10500,N_8521,N_8324);
nor U10501 (N_10501,N_5361,N_8040);
nor U10502 (N_10502,N_5543,N_6110);
xor U10503 (N_10503,N_6809,N_9380);
or U10504 (N_10504,N_7332,N_8458);
xnor U10505 (N_10505,N_5962,N_7113);
and U10506 (N_10506,N_8021,N_6842);
and U10507 (N_10507,N_9487,N_6153);
or U10508 (N_10508,N_9503,N_7416);
or U10509 (N_10509,N_8160,N_8532);
xnor U10510 (N_10510,N_7164,N_8308);
or U10511 (N_10511,N_9348,N_6122);
and U10512 (N_10512,N_6114,N_9754);
xor U10513 (N_10513,N_7343,N_5859);
or U10514 (N_10514,N_9442,N_9249);
and U10515 (N_10515,N_9068,N_8424);
or U10516 (N_10516,N_5589,N_8866);
and U10517 (N_10517,N_5117,N_5006);
xor U10518 (N_10518,N_5064,N_7187);
xnor U10519 (N_10519,N_5364,N_8797);
or U10520 (N_10520,N_9557,N_6997);
nor U10521 (N_10521,N_7907,N_6572);
or U10522 (N_10522,N_9509,N_8455);
and U10523 (N_10523,N_8130,N_9715);
or U10524 (N_10524,N_5200,N_6364);
nand U10525 (N_10525,N_8100,N_9824);
or U10526 (N_10526,N_7078,N_9020);
xnor U10527 (N_10527,N_6760,N_8482);
nor U10528 (N_10528,N_7740,N_8687);
and U10529 (N_10529,N_8816,N_6566);
nor U10530 (N_10530,N_7361,N_8753);
and U10531 (N_10531,N_9521,N_8624);
nor U10532 (N_10532,N_9279,N_9308);
and U10533 (N_10533,N_7433,N_7599);
nand U10534 (N_10534,N_7751,N_6203);
and U10535 (N_10535,N_6962,N_8211);
nor U10536 (N_10536,N_6328,N_8258);
or U10537 (N_10537,N_5291,N_5377);
nand U10538 (N_10538,N_6617,N_7512);
xnor U10539 (N_10539,N_9088,N_9393);
nor U10540 (N_10540,N_7156,N_5924);
nand U10541 (N_10541,N_8108,N_9473);
nor U10542 (N_10542,N_6034,N_5832);
and U10543 (N_10543,N_8570,N_9613);
nand U10544 (N_10544,N_7607,N_5930);
and U10545 (N_10545,N_8135,N_5846);
or U10546 (N_10546,N_8060,N_5844);
nor U10547 (N_10547,N_6395,N_7180);
and U10548 (N_10548,N_8527,N_9800);
nor U10549 (N_10549,N_7538,N_9511);
xor U10550 (N_10550,N_5985,N_6867);
and U10551 (N_10551,N_6590,N_7063);
nand U10552 (N_10552,N_5575,N_6872);
or U10553 (N_10553,N_7874,N_8964);
and U10554 (N_10554,N_8740,N_6408);
and U10555 (N_10555,N_5344,N_7355);
nor U10556 (N_10556,N_5475,N_9862);
and U10557 (N_10557,N_6061,N_9086);
nor U10558 (N_10558,N_9128,N_7140);
and U10559 (N_10559,N_9890,N_5412);
xor U10560 (N_10560,N_7461,N_6514);
nand U10561 (N_10561,N_5045,N_9423);
xnor U10562 (N_10562,N_9452,N_6361);
or U10563 (N_10563,N_7120,N_9530);
nor U10564 (N_10564,N_7718,N_7999);
nor U10565 (N_10565,N_7441,N_9804);
nor U10566 (N_10566,N_6323,N_9050);
and U10567 (N_10567,N_7884,N_6418);
and U10568 (N_10568,N_5571,N_7046);
or U10569 (N_10569,N_6462,N_5192);
or U10570 (N_10570,N_5676,N_9096);
and U10571 (N_10571,N_7203,N_9759);
nand U10572 (N_10572,N_8011,N_8471);
xnor U10573 (N_10573,N_7212,N_7624);
or U10574 (N_10574,N_6540,N_5295);
and U10575 (N_10575,N_8078,N_7102);
nor U10576 (N_10576,N_7969,N_6313);
nor U10577 (N_10577,N_6317,N_7945);
nand U10578 (N_10578,N_9430,N_6319);
nor U10579 (N_10579,N_7869,N_5628);
or U10580 (N_10580,N_8783,N_9609);
xnor U10581 (N_10581,N_6036,N_8580);
nor U10582 (N_10582,N_7128,N_8717);
or U10583 (N_10583,N_7098,N_6184);
nand U10584 (N_10584,N_6793,N_7094);
nor U10585 (N_10585,N_8946,N_7911);
and U10586 (N_10586,N_7347,N_6999);
and U10587 (N_10587,N_6611,N_5520);
and U10588 (N_10588,N_8639,N_5182);
or U10589 (N_10589,N_6599,N_6306);
nor U10590 (N_10590,N_6320,N_9665);
nor U10591 (N_10591,N_6639,N_9931);
or U10592 (N_10592,N_8215,N_5793);
or U10593 (N_10593,N_6847,N_7714);
nand U10594 (N_10594,N_7101,N_9415);
or U10595 (N_10595,N_9787,N_9306);
and U10596 (N_10596,N_7882,N_7205);
or U10597 (N_10597,N_9100,N_8232);
and U10598 (N_10598,N_6484,N_9681);
nor U10599 (N_10599,N_7498,N_7688);
or U10600 (N_10600,N_7230,N_8831);
or U10601 (N_10601,N_9942,N_8261);
or U10602 (N_10602,N_9419,N_9801);
and U10603 (N_10603,N_9000,N_8388);
xnor U10604 (N_10604,N_5831,N_7302);
nor U10605 (N_10605,N_9684,N_8116);
nand U10606 (N_10606,N_8545,N_5185);
nand U10607 (N_10607,N_8106,N_6558);
nor U10608 (N_10608,N_9999,N_9363);
xnor U10609 (N_10609,N_6379,N_6401);
nand U10610 (N_10610,N_6994,N_9197);
nand U10611 (N_10611,N_5040,N_5490);
xor U10612 (N_10612,N_8445,N_8859);
nor U10613 (N_10613,N_6348,N_5308);
and U10614 (N_10614,N_5529,N_9579);
or U10615 (N_10615,N_5579,N_5129);
or U10616 (N_10616,N_7971,N_9205);
and U10617 (N_10617,N_7262,N_7065);
xnor U10618 (N_10618,N_9320,N_6968);
nor U10619 (N_10619,N_5917,N_5882);
xor U10620 (N_10620,N_6681,N_7056);
or U10621 (N_10621,N_7275,N_5059);
or U10622 (N_10622,N_8731,N_6971);
or U10623 (N_10623,N_7431,N_5331);
nor U10624 (N_10624,N_5612,N_8389);
xnor U10625 (N_10625,N_9081,N_8579);
or U10626 (N_10626,N_8513,N_7036);
nand U10627 (N_10627,N_8781,N_8294);
nor U10628 (N_10628,N_8791,N_8079);
xnor U10629 (N_10629,N_6044,N_9849);
and U10630 (N_10630,N_7621,N_5425);
xnor U10631 (N_10631,N_9644,N_9871);
and U10632 (N_10632,N_7088,N_6018);
or U10633 (N_10633,N_7886,N_9394);
and U10634 (N_10634,N_7844,N_5739);
nor U10635 (N_10635,N_8039,N_5243);
xor U10636 (N_10636,N_7916,N_7929);
and U10637 (N_10637,N_9484,N_5447);
nor U10638 (N_10638,N_6605,N_5403);
nand U10639 (N_10639,N_5932,N_6409);
nor U10640 (N_10640,N_7352,N_6647);
and U10641 (N_10641,N_8334,N_9288);
nand U10642 (N_10642,N_7928,N_9799);
or U10643 (N_10643,N_7592,N_6687);
and U10644 (N_10644,N_7918,N_8134);
and U10645 (N_10645,N_7723,N_5002);
nor U10646 (N_10646,N_7719,N_8706);
xnor U10647 (N_10647,N_9277,N_9905);
or U10648 (N_10648,N_9535,N_7086);
xor U10649 (N_10649,N_8439,N_9428);
xnor U10650 (N_10650,N_9689,N_8025);
and U10651 (N_10651,N_6641,N_8873);
nand U10652 (N_10652,N_5085,N_7223);
or U10653 (N_10653,N_5561,N_9601);
nand U10654 (N_10654,N_6059,N_8813);
and U10655 (N_10655,N_8194,N_5238);
or U10656 (N_10656,N_7124,N_5939);
and U10657 (N_10657,N_9204,N_5974);
xor U10658 (N_10658,N_5851,N_8291);
and U10659 (N_10659,N_5736,N_8352);
xor U10660 (N_10660,N_8208,N_6435);
xnor U10661 (N_10661,N_6948,N_6248);
nand U10662 (N_10662,N_9670,N_9704);
and U10663 (N_10663,N_7333,N_6385);
or U10664 (N_10664,N_5171,N_9192);
or U10665 (N_10665,N_5260,N_5401);
nor U10666 (N_10666,N_5210,N_8686);
and U10667 (N_10667,N_6324,N_8976);
nor U10668 (N_10668,N_8229,N_9617);
or U10669 (N_10669,N_7110,N_8030);
and U10670 (N_10670,N_8301,N_9790);
or U10671 (N_10671,N_9333,N_9109);
nor U10672 (N_10672,N_9498,N_9855);
nand U10673 (N_10673,N_6926,N_5885);
nand U10674 (N_10674,N_6797,N_5322);
nor U10675 (N_10675,N_8916,N_6906);
nor U10676 (N_10676,N_6830,N_7605);
or U10677 (N_10677,N_6642,N_8371);
or U10678 (N_10678,N_6875,N_6762);
nand U10679 (N_10679,N_7905,N_6783);
and U10680 (N_10680,N_7889,N_9307);
xor U10681 (N_10681,N_7251,N_7934);
nand U10682 (N_10682,N_5504,N_8953);
and U10683 (N_10683,N_9061,N_9560);
nor U10684 (N_10684,N_6637,N_6624);
xnor U10685 (N_10685,N_7903,N_8459);
nor U10686 (N_10686,N_7255,N_6230);
nand U10687 (N_10687,N_6117,N_7555);
xor U10688 (N_10688,N_7803,N_7194);
and U10689 (N_10689,N_7224,N_7284);
and U10690 (N_10690,N_7233,N_9242);
or U10691 (N_10691,N_5465,N_8348);
xor U10692 (N_10692,N_5821,N_5711);
and U10693 (N_10693,N_9723,N_9607);
and U10694 (N_10694,N_5483,N_8414);
or U10695 (N_10695,N_9651,N_8669);
xor U10696 (N_10696,N_8952,N_8910);
xor U10697 (N_10697,N_8716,N_8735);
xor U10698 (N_10698,N_8220,N_8049);
xnor U10699 (N_10699,N_8341,N_8259);
and U10700 (N_10700,N_7962,N_7571);
and U10701 (N_10701,N_8163,N_7007);
xnor U10702 (N_10702,N_6370,N_6992);
or U10703 (N_10703,N_5745,N_7245);
xnor U10704 (N_10704,N_7009,N_8745);
or U10705 (N_10705,N_8434,N_5170);
nand U10706 (N_10706,N_7211,N_8311);
or U10707 (N_10707,N_5013,N_5833);
nor U10708 (N_10708,N_5202,N_7893);
nand U10709 (N_10709,N_9368,N_9961);
nor U10710 (N_10710,N_9191,N_8903);
nor U10711 (N_10711,N_9077,N_8861);
nor U10712 (N_10712,N_8401,N_8574);
or U10713 (N_10713,N_6390,N_6368);
nand U10714 (N_10714,N_9195,N_9220);
nor U10715 (N_10715,N_7234,N_8098);
nor U10716 (N_10716,N_5511,N_6471);
xor U10717 (N_10717,N_7733,N_9349);
or U10718 (N_10718,N_7308,N_9826);
or U10719 (N_10719,N_9812,N_7448);
nand U10720 (N_10720,N_8009,N_8732);
xnor U10721 (N_10721,N_5095,N_7925);
nor U10722 (N_10722,N_5995,N_8519);
nor U10723 (N_10723,N_6167,N_9593);
nand U10724 (N_10724,N_8954,N_5621);
xor U10725 (N_10725,N_9149,N_7403);
xor U10726 (N_10726,N_7040,N_9290);
nand U10727 (N_10727,N_8084,N_7739);
nand U10728 (N_10728,N_9710,N_9048);
nor U10729 (N_10729,N_9076,N_6222);
xnor U10730 (N_10730,N_7279,N_5505);
xnor U10731 (N_10731,N_8456,N_5637);
and U10732 (N_10732,N_9856,N_8528);
and U10733 (N_10733,N_6346,N_6237);
and U10734 (N_10734,N_5923,N_8353);
or U10735 (N_10735,N_9695,N_5458);
xor U10736 (N_10736,N_5481,N_7509);
or U10737 (N_10737,N_5374,N_8835);
xnor U10738 (N_10738,N_9292,N_8629);
nor U10739 (N_10739,N_8381,N_8326);
or U10740 (N_10740,N_7026,N_6522);
xnor U10741 (N_10741,N_5218,N_8583);
and U10742 (N_10742,N_7619,N_6151);
or U10743 (N_10743,N_9270,N_9247);
or U10744 (N_10744,N_6365,N_6958);
or U10745 (N_10745,N_7165,N_9178);
nor U10746 (N_10746,N_5223,N_6147);
xnor U10747 (N_10747,N_8988,N_6186);
or U10748 (N_10748,N_9465,N_5258);
or U10749 (N_10749,N_6128,N_9582);
nand U10750 (N_10750,N_6467,N_9328);
or U10751 (N_10751,N_6533,N_5906);
xor U10752 (N_10752,N_5383,N_7973);
or U10753 (N_10753,N_7708,N_6802);
nand U10754 (N_10754,N_5473,N_8704);
and U10755 (N_10755,N_5852,N_9721);
xor U10756 (N_10756,N_5519,N_8269);
nor U10757 (N_10757,N_6247,N_6035);
xnor U10758 (N_10758,N_9788,N_6956);
and U10759 (N_10759,N_9971,N_8584);
nor U10760 (N_10760,N_8319,N_9329);
and U10761 (N_10761,N_7331,N_5074);
nand U10762 (N_10762,N_9534,N_6157);
nand U10763 (N_10763,N_9577,N_8729);
xnor U10764 (N_10764,N_5127,N_9475);
or U10765 (N_10765,N_9918,N_6066);
nand U10766 (N_10766,N_6753,N_5121);
nand U10767 (N_10767,N_7104,N_5961);
xor U10768 (N_10768,N_8649,N_8452);
or U10769 (N_10769,N_9300,N_6644);
nand U10770 (N_10770,N_5733,N_7456);
nor U10771 (N_10771,N_6235,N_6078);
nor U10772 (N_10772,N_9596,N_6692);
or U10773 (N_10773,N_8560,N_9967);
xnor U10774 (N_10774,N_6532,N_7179);
and U10775 (N_10775,N_8357,N_5270);
and U10776 (N_10776,N_8908,N_6476);
nand U10777 (N_10777,N_6570,N_5823);
nor U10778 (N_10778,N_8202,N_6560);
xor U10779 (N_10779,N_5922,N_6881);
or U10780 (N_10780,N_5081,N_6695);
or U10781 (N_10781,N_7446,N_8641);
nor U10782 (N_10782,N_5141,N_6118);
nand U10783 (N_10783,N_5493,N_5788);
and U10784 (N_10784,N_6043,N_6416);
or U10785 (N_10785,N_6814,N_9569);
nand U10786 (N_10786,N_8290,N_5204);
and U10787 (N_10787,N_9261,N_8762);
xor U10788 (N_10788,N_8634,N_9814);
xnor U10789 (N_10789,N_5553,N_9236);
xnor U10790 (N_10790,N_7360,N_5125);
nor U10791 (N_10791,N_7318,N_9041);
xnor U10792 (N_10792,N_7344,N_8970);
or U10793 (N_10793,N_5948,N_9540);
and U10794 (N_10794,N_7487,N_8020);
nand U10795 (N_10795,N_8935,N_6202);
and U10796 (N_10796,N_6913,N_7581);
nor U10797 (N_10797,N_7117,N_9281);
and U10798 (N_10798,N_7134,N_9574);
or U10799 (N_10799,N_5143,N_5989);
nand U10800 (N_10800,N_7445,N_6001);
nor U10801 (N_10801,N_9713,N_9657);
xnor U10802 (N_10802,N_9401,N_8068);
nor U10803 (N_10803,N_9774,N_9379);
or U10804 (N_10804,N_7341,N_8743);
xnor U10805 (N_10805,N_9693,N_6511);
xnor U10806 (N_10806,N_5678,N_6735);
nor U10807 (N_10807,N_5399,N_9163);
and U10808 (N_10808,N_7771,N_8012);
xor U10809 (N_10809,N_6738,N_6131);
or U10810 (N_10810,N_8392,N_6120);
nor U10811 (N_10811,N_7082,N_6665);
and U10812 (N_10812,N_8826,N_7264);
and U10813 (N_10813,N_9928,N_9459);
nor U10814 (N_10814,N_7073,N_7422);
xnor U10815 (N_10815,N_5827,N_8811);
or U10816 (N_10816,N_9026,N_8335);
nand U10817 (N_10817,N_6496,N_5605);
xnor U10818 (N_10818,N_6920,N_5120);
and U10819 (N_10819,N_5486,N_9291);
xnor U10820 (N_10820,N_9898,N_5457);
nor U10821 (N_10821,N_5114,N_7947);
or U10822 (N_10822,N_7084,N_7824);
nand U10823 (N_10823,N_7995,N_9233);
nand U10824 (N_10824,N_8316,N_5898);
nand U10825 (N_10825,N_8246,N_9479);
or U10826 (N_10826,N_9176,N_8213);
nor U10827 (N_10827,N_8004,N_6739);
and U10828 (N_10828,N_7735,N_9585);
and U10829 (N_10829,N_8851,N_8944);
and U10830 (N_10830,N_5213,N_9039);
or U10831 (N_10831,N_6509,N_5303);
or U10832 (N_10832,N_6882,N_9282);
and U10833 (N_10833,N_7139,N_9321);
and U10834 (N_10834,N_5152,N_5371);
nor U10835 (N_10835,N_8095,N_8359);
xor U10836 (N_10836,N_5108,N_8197);
nor U10837 (N_10837,N_9742,N_8080);
and U10838 (N_10838,N_5560,N_6640);
and U10839 (N_10839,N_5707,N_5115);
nand U10840 (N_10840,N_8008,N_6367);
nand U10841 (N_10841,N_9310,N_6960);
nand U10842 (N_10842,N_9130,N_8472);
nor U10843 (N_10843,N_7378,N_7042);
nor U10844 (N_10844,N_6567,N_8345);
and U10845 (N_10845,N_8171,N_9259);
or U10846 (N_10846,N_6123,N_8241);
xnor U10847 (N_10847,N_7923,N_7338);
and U10848 (N_10848,N_9198,N_8555);
nor U10849 (N_10849,N_6398,N_7469);
and U10850 (N_10850,N_8611,N_7025);
and U10851 (N_10851,N_6996,N_6600);
and U10852 (N_10852,N_5669,N_6239);
or U10853 (N_10853,N_9301,N_7968);
xor U10854 (N_10854,N_9863,N_8161);
nand U10855 (N_10855,N_8370,N_6979);
xnor U10856 (N_10856,N_5298,N_5548);
nand U10857 (N_10857,N_6631,N_7209);
and U10858 (N_10858,N_8132,N_6908);
nor U10859 (N_10859,N_8343,N_7012);
nor U10860 (N_10860,N_8670,N_8115);
nand U10861 (N_10861,N_6869,N_7236);
nor U10862 (N_10862,N_8674,N_6529);
and U10863 (N_10863,N_8092,N_6883);
or U10864 (N_10864,N_7639,N_6183);
nor U10865 (N_10865,N_9184,N_9690);
or U10866 (N_10866,N_7892,N_7216);
xnor U10867 (N_10867,N_9673,N_5584);
nand U10868 (N_10868,N_6848,N_5373);
or U10869 (N_10869,N_6705,N_6543);
or U10870 (N_10870,N_9615,N_5944);
xor U10871 (N_10871,N_5423,N_5203);
or U10872 (N_10872,N_8128,N_5302);
and U10873 (N_10873,N_7159,N_9746);
or U10874 (N_10874,N_6055,N_8561);
xor U10875 (N_10875,N_6428,N_5153);
and U10876 (N_10876,N_5419,N_6812);
xnor U10877 (N_10877,N_6286,N_7100);
nand U10878 (N_10878,N_7657,N_5531);
nor U10879 (N_10879,N_6925,N_7414);
and U10880 (N_10880,N_9831,N_9620);
and U10881 (N_10881,N_6296,N_9330);
or U10882 (N_10882,N_7109,N_7374);
and U10883 (N_10883,N_7477,N_8045);
xor U10884 (N_10884,N_8103,N_5542);
or U10885 (N_10885,N_5306,N_8338);
xor U10886 (N_10886,N_5500,N_9606);
nand U10887 (N_10887,N_5106,N_8980);
and U10888 (N_10888,N_5791,N_9144);
xnor U10889 (N_10889,N_8372,N_6438);
or U10890 (N_10890,N_5234,N_8056);
or U10891 (N_10891,N_6255,N_5949);
nor U10892 (N_10892,N_8221,N_7933);
nor U10893 (N_10893,N_5897,N_8761);
or U10894 (N_10894,N_7417,N_7847);
xor U10895 (N_10895,N_6497,N_5309);
xnor U10896 (N_10896,N_9040,N_9189);
and U10897 (N_10897,N_6585,N_7201);
or U10898 (N_10898,N_9661,N_5339);
xnor U10899 (N_10899,N_9807,N_8138);
nor U10900 (N_10900,N_8427,N_8284);
or U10901 (N_10901,N_6020,N_8479);
xor U10902 (N_10902,N_5409,N_5915);
xnor U10903 (N_10903,N_5492,N_6188);
nand U10904 (N_10904,N_7514,N_9686);
or U10905 (N_10905,N_5877,N_7126);
nand U10906 (N_10906,N_8096,N_8002);
xnor U10907 (N_10907,N_5537,N_7746);
xnor U10908 (N_10908,N_9099,N_6584);
or U10909 (N_10909,N_7467,N_9598);
nand U10910 (N_10910,N_7752,N_9397);
nand U10911 (N_10911,N_9494,N_9012);
or U10912 (N_10912,N_8118,N_9945);
nand U10913 (N_10913,N_9140,N_7696);
xor U10914 (N_10914,N_7247,N_7951);
or U10915 (N_10915,N_9731,N_5610);
nand U10916 (N_10916,N_6628,N_7501);
nand U10917 (N_10917,N_7146,N_8064);
or U10918 (N_10918,N_9502,N_5802);
nor U10919 (N_10919,N_7541,N_7926);
xnor U10920 (N_10920,N_8240,N_6520);
nor U10921 (N_10921,N_9005,N_5694);
xor U10922 (N_10922,N_7096,N_5058);
xnor U10923 (N_10923,N_6326,N_5452);
and U10924 (N_10924,N_9043,N_6090);
nand U10925 (N_10925,N_8199,N_9642);
nand U10926 (N_10926,N_5267,N_7836);
xor U10927 (N_10927,N_9600,N_5876);
and U10928 (N_10928,N_7948,N_6448);
nor U10929 (N_10929,N_8391,N_8742);
nand U10930 (N_10930,N_6562,N_7177);
nand U10931 (N_10931,N_7289,N_7997);
or U10932 (N_10932,N_7785,N_5188);
xor U10933 (N_10933,N_7804,N_7426);
nor U10934 (N_10934,N_8436,N_6008);
nor U10935 (N_10935,N_9639,N_9683);
xor U10936 (N_10936,N_5342,N_7023);
xor U10937 (N_10937,N_8344,N_5993);
and U10938 (N_10938,N_6763,N_8961);
nor U10939 (N_10939,N_6045,N_6528);
or U10940 (N_10940,N_7850,N_9956);
nand U10941 (N_10941,N_5292,N_7835);
nor U10942 (N_10942,N_8710,N_9632);
nor U10943 (N_10943,N_7543,N_7877);
nor U10944 (N_10944,N_6553,N_6019);
xor U10945 (N_10945,N_6580,N_7470);
nor U10946 (N_10946,N_8073,N_6717);
xnor U10947 (N_10947,N_6477,N_6742);
and U10948 (N_10948,N_7595,N_9467);
xnor U10949 (N_10949,N_6372,N_7227);
and U10950 (N_10950,N_8562,N_9304);
or U10951 (N_10951,N_7742,N_9750);
nand U10952 (N_10952,N_9010,N_7517);
xnor U10953 (N_10953,N_6754,N_9966);
nor U10954 (N_10954,N_9018,N_9866);
nand U10955 (N_10955,N_8399,N_8431);
nor U10956 (N_10956,N_5507,N_8569);
nand U10957 (N_10957,N_5046,N_9797);
or U10958 (N_10958,N_8768,N_9446);
or U10959 (N_10959,N_7465,N_9602);
nand U10960 (N_10960,N_8292,N_6586);
or U10961 (N_10961,N_6810,N_6156);
xnor U10962 (N_10962,N_9203,N_6595);
nand U10963 (N_10963,N_6429,N_6282);
xor U10964 (N_10964,N_7584,N_9293);
or U10965 (N_10965,N_9294,N_6085);
xor U10966 (N_10966,N_6080,N_5562);
xnor U10967 (N_10967,N_7317,N_6423);
nand U10968 (N_10968,N_6541,N_7158);
xnor U10969 (N_10969,N_6643,N_8421);
nor U10970 (N_10970,N_9460,N_9269);
xnor U10971 (N_10971,N_8447,N_8502);
or U10972 (N_10972,N_8306,N_5867);
or U10973 (N_10973,N_8494,N_9743);
and U10974 (N_10974,N_9324,N_9152);
or U10975 (N_10975,N_8400,N_6437);
and U10976 (N_10976,N_7411,N_7271);
nor U10977 (N_10977,N_7408,N_8470);
and U10978 (N_10978,N_9765,N_8198);
or U10979 (N_10979,N_5672,N_9112);
nand U10980 (N_10980,N_5096,N_7980);
or U10981 (N_10981,N_6224,N_9142);
or U10982 (N_10982,N_9980,N_5762);
xor U10983 (N_10983,N_7851,N_9303);
or U10984 (N_10984,N_7859,N_6314);
xnor U10985 (N_10985,N_5443,N_5382);
xor U10986 (N_10986,N_8050,N_7160);
and U10987 (N_10987,N_8530,N_5136);
nand U10988 (N_10988,N_6067,N_9974);
nand U10989 (N_10989,N_7717,N_7631);
and U10990 (N_10990,N_6519,N_9463);
and U10991 (N_10991,N_5783,N_5293);
xor U10992 (N_10992,N_7950,N_7119);
and U10993 (N_10993,N_8450,N_5527);
or U10994 (N_10994,N_5211,N_6963);
or U10995 (N_10995,N_7323,N_5997);
xnor U10996 (N_10996,N_9190,N_9180);
xor U10997 (N_10997,N_5855,N_7858);
xnor U10998 (N_10998,N_5014,N_9762);
or U10999 (N_10999,N_9994,N_6426);
nor U11000 (N_11000,N_8844,N_5179);
nor U11001 (N_11001,N_9542,N_8985);
xor U11002 (N_11002,N_8457,N_9899);
or U11003 (N_11003,N_6144,N_5249);
xnor U11004 (N_11004,N_7654,N_9360);
or U11005 (N_11005,N_7479,N_6400);
and U11006 (N_11006,N_7573,N_5987);
nand U11007 (N_11007,N_7363,N_7813);
nor U11008 (N_11008,N_8914,N_9098);
xor U11009 (N_11009,N_7075,N_7763);
xnor U11010 (N_11010,N_8186,N_9215);
nand U11011 (N_11011,N_8395,N_7758);
nor U11012 (N_11012,N_8630,N_8880);
nor U11013 (N_11013,N_6671,N_6351);
nor U11014 (N_11014,N_9450,N_6773);
or U11015 (N_11015,N_8247,N_8148);
nand U11016 (N_11016,N_6164,N_5903);
or U11017 (N_11017,N_8974,N_9376);
nand U11018 (N_11018,N_8928,N_8636);
nand U11019 (N_11019,N_7144,N_5338);
nand U11020 (N_11020,N_9817,N_9832);
xor U11021 (N_11021,N_5810,N_7396);
or U11022 (N_11022,N_8924,N_7274);
or U11023 (N_11023,N_9439,N_6907);
and U11024 (N_11024,N_5044,N_7940);
or U11025 (N_11025,N_6201,N_6821);
xor U11026 (N_11026,N_8046,N_6751);
and U11027 (N_11027,N_8158,N_8995);
or U11028 (N_11028,N_6205,N_9567);
or U11029 (N_11029,N_9228,N_9272);
xnor U11030 (N_11030,N_8728,N_8027);
nor U11031 (N_11031,N_5389,N_7658);
or U11032 (N_11032,N_6916,N_7353);
or U11033 (N_11033,N_9925,N_9139);
nor U11034 (N_11034,N_8207,N_9440);
nand U11035 (N_11035,N_9340,N_9699);
nand U11036 (N_11036,N_8412,N_9573);
nor U11037 (N_11037,N_7588,N_8397);
xor U11038 (N_11038,N_8538,N_5946);
nand U11039 (N_11039,N_9541,N_7665);
or U11040 (N_11040,N_6573,N_9443);
or U11041 (N_11041,N_5428,N_7894);
nor U11042 (N_11042,N_8225,N_7931);
nor U11043 (N_11043,N_5147,N_6071);
and U11044 (N_11044,N_5618,N_7295);
nor U11045 (N_11045,N_5539,N_8643);
or U11046 (N_11046,N_9603,N_9900);
nor U11047 (N_11047,N_5246,N_8785);
and U11048 (N_11048,N_9305,N_6662);
xnor U11049 (N_11049,N_8984,N_9834);
or U11050 (N_11050,N_8373,N_9365);
or U11051 (N_11051,N_6546,N_9850);
nor U11052 (N_11052,N_5816,N_7340);
nor U11053 (N_11053,N_9445,N_8929);
xor U11054 (N_11054,N_9335,N_8945);
nor U11055 (N_11055,N_5518,N_5168);
nor U11056 (N_11056,N_6563,N_6386);
or U11057 (N_11057,N_9410,N_6601);
or U11058 (N_11058,N_7817,N_8807);
nor U11059 (N_11059,N_7932,N_8114);
xnor U11060 (N_11060,N_6276,N_9802);
or U11061 (N_11061,N_5813,N_6236);
xor U11062 (N_11062,N_6734,N_9245);
and U11063 (N_11063,N_8618,N_9400);
nand U11064 (N_11064,N_8787,N_8683);
and U11065 (N_11065,N_6138,N_9072);
nor U11066 (N_11066,N_7920,N_8755);
nor U11067 (N_11067,N_8177,N_6339);
nand U11068 (N_11068,N_6806,N_9207);
and U11069 (N_11069,N_9660,N_7921);
nand U11070 (N_11070,N_7511,N_5860);
nor U11071 (N_11071,N_9873,N_6952);
nor U11072 (N_11072,N_8978,N_8514);
xor U11073 (N_11073,N_5427,N_6489);
or U11074 (N_11074,N_7848,N_9614);
and U11075 (N_11075,N_6976,N_5866);
and U11076 (N_11076,N_9185,N_7685);
nand U11077 (N_11077,N_7630,N_8764);
nand U11078 (N_11078,N_6664,N_6161);
xor U11079 (N_11079,N_9155,N_5667);
xor U11080 (N_11080,N_5840,N_7176);
xor U11081 (N_11081,N_6070,N_6194);
and U11082 (N_11082,N_9409,N_6799);
nand U11083 (N_11083,N_9160,N_8932);
nand U11084 (N_11084,N_7736,N_7797);
nand U11085 (N_11085,N_9193,N_5352);
or U11086 (N_11086,N_9105,N_6421);
or U11087 (N_11087,N_9371,N_6485);
and U11088 (N_11088,N_6452,N_9637);
nand U11089 (N_11089,N_6154,N_7376);
and U11090 (N_11090,N_5433,N_9141);
and U11091 (N_11091,N_8226,N_8991);
nand U11092 (N_11092,N_5977,N_6029);
nand U11093 (N_11093,N_8498,N_9268);
nor U11094 (N_11094,N_8895,N_9714);
nand U11095 (N_11095,N_8693,N_8286);
xnor U11096 (N_11096,N_8176,N_7079);
nor U11097 (N_11097,N_7377,N_9646);
and U11098 (N_11098,N_5254,N_6375);
or U11099 (N_11099,N_8699,N_6394);
nand U11100 (N_11100,N_7944,N_6961);
nand U11101 (N_11101,N_6417,N_7542);
nand U11102 (N_11102,N_5227,N_8418);
and U11103 (N_11103,N_6134,N_7155);
and U11104 (N_11104,N_6369,N_7127);
nor U11105 (N_11105,N_6873,N_8942);
and U11106 (N_11106,N_9587,N_9341);
nand U11107 (N_11107,N_7217,N_9273);
xnor U11108 (N_11108,N_9256,N_7819);
or U11109 (N_11109,N_6937,N_6327);
or U11110 (N_11110,N_6766,N_6702);
nor U11111 (N_11111,N_5952,N_5722);
or U11112 (N_11112,N_9547,N_5981);
nand U11113 (N_11113,N_5380,N_8681);
nor U11114 (N_11114,N_5795,N_6102);
nand U11115 (N_11115,N_6815,N_9243);
nand U11116 (N_11116,N_8602,N_5397);
and U11117 (N_11117,N_8596,N_9028);
and U11118 (N_11118,N_7562,N_5609);
nand U11119 (N_11119,N_6798,N_8054);
nand U11120 (N_11120,N_9555,N_7596);
nand U11121 (N_11121,N_8692,N_6092);
nand U11122 (N_11122,N_7853,N_5884);
and U11123 (N_11123,N_6921,N_7576);
nand U11124 (N_11124,N_9705,N_7020);
or U11125 (N_11125,N_6332,N_7566);
nand U11126 (N_11126,N_9238,N_8524);
or U11127 (N_11127,N_9730,N_5980);
nor U11128 (N_11128,N_6822,N_8057);
nand U11129 (N_11129,N_6627,N_7191);
and U11130 (N_11130,N_8876,N_5445);
xnor U11131 (N_11131,N_5079,N_6010);
xnor U11132 (N_11132,N_6000,N_7402);
nor U11133 (N_11133,N_7397,N_5908);
nand U11134 (N_11134,N_7099,N_5841);
or U11135 (N_11135,N_8733,N_5012);
or U11136 (N_11136,N_6170,N_5751);
or U11137 (N_11137,N_8656,N_5834);
or U11138 (N_11138,N_6058,N_7371);
or U11139 (N_11139,N_8029,N_9426);
nand U11140 (N_11140,N_7423,N_6136);
or U11141 (N_11141,N_6382,N_9776);
nand U11142 (N_11142,N_7695,N_8268);
and U11143 (N_11143,N_6023,N_6270);
nor U11144 (N_11144,N_7200,N_9629);
nor U11145 (N_11145,N_5564,N_9524);
nor U11146 (N_11146,N_9882,N_9337);
nand U11147 (N_11147,N_8694,N_6733);
nor U11148 (N_11148,N_8295,N_7277);
xnor U11149 (N_11149,N_5767,N_5487);
xor U11150 (N_11150,N_7656,N_7229);
nand U11151 (N_11151,N_8422,N_5690);
nor U11152 (N_11152,N_7459,N_7462);
and U11153 (N_11153,N_7256,N_6208);
nand U11154 (N_11154,N_5324,N_6829);
nand U11155 (N_11155,N_9396,N_9538);
or U11156 (N_11156,N_7325,N_9447);
and U11157 (N_11157,N_8700,N_7915);
or U11158 (N_11158,N_8181,N_6414);
nand U11159 (N_11159,N_7254,N_6305);
and U11160 (N_11160,N_8437,N_7939);
and U11161 (N_11161,N_6612,N_9067);
nand U11162 (N_11162,N_6155,N_7860);
nand U11163 (N_11163,N_9922,N_6130);
nor U11164 (N_11164,N_8554,N_9977);
nand U11165 (N_11165,N_7261,N_9482);
xor U11166 (N_11166,N_7908,N_6932);
and U11167 (N_11167,N_8727,N_8346);
nor U11168 (N_11168,N_7641,N_8137);
and U11169 (N_11169,N_8709,N_5868);
nor U11170 (N_11170,N_6629,N_7802);
nor U11171 (N_11171,N_6172,N_5541);
and U11172 (N_11172,N_8111,N_6934);
and U11173 (N_11173,N_8769,N_6266);
and U11174 (N_11174,N_6331,N_8224);
or U11175 (N_11175,N_5784,N_8019);
and U11176 (N_11176,N_8441,N_6124);
xnor U11177 (N_11177,N_8882,N_7196);
or U11178 (N_11178,N_9114,N_8136);
and U11179 (N_11179,N_9250,N_5055);
nor U11180 (N_11180,N_8280,N_7244);
and U11181 (N_11181,N_5720,N_9049);
or U11182 (N_11182,N_5268,N_5145);
or U11183 (N_11183,N_6303,N_6894);
or U11184 (N_11184,N_8775,N_7949);
xor U11185 (N_11185,N_8806,N_6825);
nand U11186 (N_11186,N_8986,N_5864);
or U11187 (N_11187,N_7037,N_9654);
and U11188 (N_11188,N_8948,N_6076);
xor U11189 (N_11189,N_5350,N_9649);
or U11190 (N_11190,N_5847,N_5285);
nand U11191 (N_11191,N_8585,N_7961);
nor U11192 (N_11192,N_9353,N_8911);
xor U11193 (N_11193,N_9539,N_7720);
and U11194 (N_11194,N_8340,N_7471);
nand U11195 (N_11195,N_8875,N_7495);
or U11196 (N_11196,N_8930,N_5809);
xor U11197 (N_11197,N_9892,N_5675);
and U11198 (N_11198,N_9476,N_5580);
nand U11199 (N_11199,N_5312,N_6406);
or U11200 (N_11200,N_8915,N_7784);
or U11201 (N_11201,N_8250,N_8278);
xor U11202 (N_11202,N_6870,N_8544);
xor U11203 (N_11203,N_9246,N_6377);
or U11204 (N_11204,N_6404,N_9827);
nor U11205 (N_11205,N_9773,N_9883);
xor U11206 (N_11206,N_7650,N_5130);
or U11207 (N_11207,N_6673,N_8722);
xor U11208 (N_11208,N_7480,N_9289);
nor U11209 (N_11209,N_9972,N_7132);
and U11210 (N_11210,N_6910,N_9688);
nor U11211 (N_11211,N_8557,N_6539);
xnor U11212 (N_11212,N_6427,N_6292);
xor U11213 (N_11213,N_6899,N_6677);
xnor U11214 (N_11214,N_6843,N_7259);
nor U11215 (N_11215,N_5661,N_7522);
nand U11216 (N_11216,N_6941,N_6879);
or U11217 (N_11217,N_7452,N_8588);
or U11218 (N_11218,N_7618,N_5174);
nor U11219 (N_11219,N_6876,N_8840);
nor U11220 (N_11220,N_5476,N_7531);
and U11221 (N_11221,N_5497,N_8682);
nand U11222 (N_11222,N_9973,N_8501);
or U11223 (N_11223,N_9691,N_9805);
xor U11224 (N_11224,N_8151,N_8890);
or U11225 (N_11225,N_8902,N_5983);
nand U11226 (N_11226,N_8938,N_7091);
or U11227 (N_11227,N_8874,N_7712);
and U11228 (N_11228,N_6256,N_5594);
and U11229 (N_11229,N_5727,N_8537);
nor U11230 (N_11230,N_6981,N_6504);
and U11231 (N_11231,N_8404,N_9655);
nor U11232 (N_11232,N_7697,N_6160);
nand U11233 (N_11233,N_5655,N_7591);
xnor U11234 (N_11234,N_5772,N_9164);
nor U11235 (N_11235,N_6517,N_8454);
nor U11236 (N_11236,N_7651,N_5526);
nand U11237 (N_11237,N_6267,N_7320);
xor U11238 (N_11238,N_9888,N_7464);
nor U11239 (N_11239,N_6150,N_8265);
or U11240 (N_11240,N_9122,N_5830);
nand U11241 (N_11241,N_5280,N_8662);
xor U11242 (N_11242,N_8244,N_7175);
and U11243 (N_11243,N_8433,N_8565);
nor U11244 (N_11244,N_9965,N_5349);
and U11245 (N_11245,N_8718,N_8059);
or U11246 (N_11246,N_9038,N_7902);
nor U11247 (N_11247,N_7407,N_8321);
nand U11248 (N_11248,N_9134,N_8962);
nor U11249 (N_11249,N_5259,N_8032);
nor U11250 (N_11250,N_8939,N_6897);
and U11251 (N_11251,N_9896,N_7822);
nand U11252 (N_11252,N_7068,N_8442);
and U11253 (N_11253,N_7485,N_7258);
and U11254 (N_11254,N_6048,N_7716);
and U11255 (N_11255,N_8535,N_7185);
nor U11256 (N_11256,N_5378,N_9652);
and U11257 (N_11257,N_5073,N_8497);
and U11258 (N_11258,N_5334,N_9727);
xor U11259 (N_11259,N_7700,N_5027);
nand U11260 (N_11260,N_6568,N_6725);
nor U11261 (N_11261,N_9468,N_9124);
xnor U11262 (N_11262,N_8523,N_5209);
and U11263 (N_11263,N_8815,N_7064);
xor U11264 (N_11264,N_5808,N_9697);
nand U11265 (N_11265,N_5535,N_9919);
nand U11266 (N_11266,N_5685,N_6432);
or U11267 (N_11267,N_7593,N_9499);
xor U11268 (N_11268,N_6817,N_9897);
xor U11269 (N_11269,N_5422,N_5332);
or U11270 (N_11270,N_8737,N_7887);
nor U11271 (N_11271,N_7978,N_5470);
and U11272 (N_11272,N_5311,N_9989);
or U11273 (N_11273,N_8361,N_6125);
or U11274 (N_11274,N_8233,N_5642);
xnor U11275 (N_11275,N_8488,N_5656);
nand U11276 (N_11276,N_8756,N_6127);
nor U11277 (N_11277,N_5588,N_8889);
nand U11278 (N_11278,N_9786,N_7024);
or U11279 (N_11279,N_7174,N_8788);
nor U11280 (N_11280,N_8253,N_8262);
nor U11281 (N_11281,N_9962,N_9424);
xnor U11282 (N_11282,N_5172,N_5540);
and U11283 (N_11283,N_9784,N_8999);
xor U11284 (N_11284,N_7301,N_7638);
nor U11285 (N_11285,N_9878,N_6422);
or U11286 (N_11286,N_6953,N_9934);
or U11287 (N_11287,N_8462,N_6737);
xor U11288 (N_11288,N_9125,N_6168);
and U11289 (N_11289,N_6801,N_5434);
nand U11290 (N_11290,N_9485,N_5333);
nor U11291 (N_11291,N_9554,N_9244);
and U11292 (N_11292,N_6534,N_8606);
nand U11293 (N_11293,N_5721,N_5693);
nand U11294 (N_11294,N_7748,N_6302);
nand U11295 (N_11295,N_5089,N_5189);
xnor U11296 (N_11296,N_9767,N_5107);
or U11297 (N_11297,N_7750,N_5668);
or U11298 (N_11298,N_6970,N_9915);
xor U11299 (N_11299,N_8274,N_8486);
and U11300 (N_11300,N_7823,N_5406);
and U11301 (N_11301,N_8746,N_5648);
nor U11302 (N_11302,N_5446,N_5770);
nand U11303 (N_11303,N_6193,N_7603);
or U11304 (N_11304,N_5735,N_8296);
nand U11305 (N_11305,N_6758,N_6281);
nor U11306 (N_11306,N_5321,N_5442);
or U11307 (N_11307,N_5586,N_7927);
xor U11308 (N_11308,N_7828,N_9078);
nor U11309 (N_11309,N_7218,N_5010);
and U11310 (N_11310,N_7900,N_7586);
nand U11311 (N_11311,N_7820,N_6661);
xor U11312 (N_11312,N_8305,N_7373);
nor U11313 (N_11313,N_7178,N_7912);
and U11314 (N_11314,N_5601,N_7646);
xnor U11315 (N_11315,N_7474,N_6565);
nand U11316 (N_11316,N_6736,N_7401);
nor U11317 (N_11317,N_7207,N_5794);
nor U11318 (N_11318,N_5325,N_5177);
and U11319 (N_11319,N_6098,N_7473);
nand U11320 (N_11320,N_5363,N_6318);
xnor U11321 (N_11321,N_8417,N_7952);
nand U11322 (N_11322,N_9035,N_5902);
xnor U11323 (N_11323,N_8887,N_8668);
xnor U11324 (N_11324,N_8971,N_5615);
nand U11325 (N_11325,N_8053,N_8526);
nand U11326 (N_11326,N_8661,N_6959);
nor U11327 (N_11327,N_5318,N_7917);
nor U11328 (N_11328,N_8097,N_7520);
and U11329 (N_11329,N_8072,N_8085);
nor U11330 (N_11330,N_6694,N_6730);
nor U11331 (N_11331,N_6472,N_8109);
and U11332 (N_11332,N_7984,N_8517);
nor U11333 (N_11333,N_9594,N_7283);
or U11334 (N_11334,N_8191,N_6915);
nor U11335 (N_11335,N_6433,N_5116);
xnor U11336 (N_11336,N_6683,N_5358);
nand U11337 (N_11337,N_9406,N_6507);
and U11338 (N_11338,N_9437,N_5198);
xnor U11339 (N_11339,N_5965,N_6711);
nand U11340 (N_11340,N_9913,N_6989);
nand U11341 (N_11341,N_8383,N_5355);
and U11342 (N_11342,N_5214,N_5937);
xor U11343 (N_11343,N_5801,N_9454);
nor U11344 (N_11344,N_8926,N_6513);
nor U11345 (N_11345,N_6458,N_5513);
nor U11346 (N_11346,N_5271,N_9604);
xor U11347 (N_11347,N_5931,N_7001);
and U11348 (N_11348,N_7404,N_9853);
nor U11349 (N_11349,N_5996,N_9703);
nand U11350 (N_11350,N_6792,N_7568);
nand U11351 (N_11351,N_5489,N_6436);
or U11352 (N_11352,N_9543,N_9929);
xnor U11353 (N_11353,N_7085,N_8426);
nor U11354 (N_11354,N_8892,N_9522);
and U11355 (N_11355,N_5036,N_5574);
nand U11356 (N_11356,N_5509,N_6419);
nand U11357 (N_11357,N_7204,N_9576);
nor U11358 (N_11358,N_5633,N_6234);
xnor U11359 (N_11359,N_8878,N_5215);
and U11360 (N_11360,N_8315,N_5348);
and U11361 (N_11361,N_6503,N_5041);
and U11362 (N_11362,N_5825,N_6715);
and U11363 (N_11363,N_6526,N_6604);
and U11364 (N_11364,N_9053,N_9381);
or U11365 (N_11365,N_5351,N_9578);
nand U11366 (N_11366,N_7677,N_7030);
nor U11367 (N_11367,N_9998,N_5874);
nor U11368 (N_11368,N_7614,N_8758);
and U11369 (N_11369,N_5196,N_7457);
or U11370 (N_11370,N_9640,N_5581);
xnor U11371 (N_11371,N_6176,N_6726);
nand U11372 (N_11372,N_9506,N_6285);
nor U11373 (N_11373,N_8509,N_5393);
xnor U11374 (N_11374,N_5070,N_6845);
nor U11375 (N_11375,N_9717,N_9255);
and U11376 (N_11376,N_6316,N_9210);
and U11377 (N_11377,N_8907,N_5054);
xnor U11378 (N_11378,N_6837,N_8568);
and U11379 (N_11379,N_6828,N_5028);
nand U11380 (N_11380,N_8934,N_9563);
xnor U11381 (N_11381,N_8642,N_6206);
nor U11382 (N_11382,N_6775,N_7798);
or U11383 (N_11383,N_7033,N_8888);
nand U11384 (N_11384,N_9127,N_7232);
nor U11385 (N_11385,N_6583,N_7793);
xor U11386 (N_11386,N_9083,N_8415);
xor U11387 (N_11387,N_8593,N_7387);
xor U11388 (N_11388,N_8153,N_9495);
nand U11389 (N_11389,N_8318,N_5379);
nand U11390 (N_11390,N_8101,N_5666);
xor U11391 (N_11391,N_7738,N_6723);
xor U11392 (N_11392,N_7327,N_6656);
xor U11393 (N_11393,N_5432,N_5431);
nand U11394 (N_11394,N_8354,N_7642);
xnor U11395 (N_11395,N_7533,N_9266);
nor U11396 (N_11396,N_8203,N_8484);
or U11397 (N_11397,N_8043,N_8667);
nor U11398 (N_11398,N_5148,N_7188);
nor U11399 (N_11399,N_5954,N_8684);
and U11400 (N_11400,N_8183,N_5684);
nand U11401 (N_11401,N_5150,N_5051);
nor U11402 (N_11402,N_5368,N_9015);
nand U11403 (N_11403,N_5769,N_5420);
nor U11404 (N_11404,N_9923,N_5307);
or U11405 (N_11405,N_8299,N_9258);
and U11406 (N_11406,N_6964,N_9060);
or U11407 (N_11407,N_6998,N_9643);
nor U11408 (N_11408,N_8023,N_7081);
or U11409 (N_11409,N_6914,N_6112);
nor U11410 (N_11410,N_6074,N_8893);
nand U11411 (N_11411,N_9830,N_8652);
or U11412 (N_11412,N_5665,N_5299);
nand U11413 (N_11413,N_5499,N_6329);
and U11414 (N_11414,N_9951,N_8983);
nor U11415 (N_11415,N_6101,N_6454);
and U11416 (N_11416,N_7238,N_5626);
or U11417 (N_11417,N_8033,N_5263);
nand U11418 (N_11418,N_7051,N_7680);
nor U11419 (N_11419,N_6308,N_6060);
nor U11420 (N_11420,N_9783,N_9561);
nand U11421 (N_11421,N_5112,N_8460);
and U11422 (N_11422,N_9019,N_8977);
and U11423 (N_11423,N_5216,N_5646);
nand U11424 (N_11424,N_6703,N_5912);
nor U11425 (N_11425,N_8854,N_6689);
or U11426 (N_11426,N_5686,N_8563);
or U11427 (N_11427,N_5067,N_6300);
xor U11428 (N_11428,N_7544,N_5639);
nand U11429 (N_11429,N_8773,N_6173);
nand U11430 (N_11430,N_7536,N_7749);
nor U11431 (N_11431,N_5779,N_9489);
nor U11432 (N_11432,N_7496,N_7705);
nand U11433 (N_11433,N_5765,N_5631);
nor U11434 (N_11434,N_7831,N_9860);
xor U11435 (N_11435,N_6449,N_7878);
nand U11436 (N_11436,N_8734,N_9296);
nand U11437 (N_11437,N_9338,N_8402);
or U11438 (N_11438,N_7589,N_5029);
and U11439 (N_11439,N_8285,N_8102);
xor U11440 (N_11440,N_7966,N_8387);
and U11441 (N_11441,N_9975,N_5781);
and U11442 (N_11442,N_6865,N_7005);
nor U11443 (N_11443,N_9775,N_9584);
nor U11444 (N_11444,N_6220,N_5764);
or U11445 (N_11445,N_5042,N_8310);
nor U11446 (N_11446,N_6005,N_6470);
and U11447 (N_11447,N_5710,N_5241);
nor U11448 (N_11448,N_7382,N_6261);
xor U11449 (N_11449,N_8309,N_8169);
nor U11450 (N_11450,N_5634,N_8955);
and U11451 (N_11451,N_9868,N_6407);
xnor U11452 (N_11452,N_8843,N_9154);
nand U11453 (N_11453,N_6396,N_6031);
nor U11454 (N_11454,N_5602,N_7391);
xnor U11455 (N_11455,N_7625,N_9838);
xor U11456 (N_11456,N_5346,N_8384);
nand U11457 (N_11457,N_9738,N_8303);
xnor U11458 (N_11458,N_9343,N_5366);
or U11459 (N_11459,N_7060,N_8495);
or U11460 (N_11460,N_9466,N_5807);
nand U11461 (N_11461,N_9311,N_9382);
or U11462 (N_11462,N_9361,N_7977);
and U11463 (N_11463,N_7637,N_5870);
xnor U11464 (N_11464,N_9791,N_5265);
nand U11465 (N_11465,N_5134,N_6930);
and U11466 (N_11466,N_5460,N_6137);
or U11467 (N_11467,N_9027,N_5193);
xnor U11468 (N_11468,N_7273,N_6376);
nor U11469 (N_11469,N_8941,N_7093);
xnor U11470 (N_11470,N_6555,N_8632);
nand U11471 (N_11471,N_7311,N_5826);
or U11472 (N_11472,N_7791,N_8830);
nor U11473 (N_11473,N_5077,N_6561);
or U11474 (N_11474,N_6578,N_6512);
xor U11475 (N_11475,N_7002,N_7430);
xor U11476 (N_11476,N_8500,N_9470);
xor U11477 (N_11477,N_8038,N_7206);
nand U11478 (N_11478,N_8473,N_9129);
or U11479 (N_11479,N_7346,N_5100);
xor U11480 (N_11480,N_5554,N_9457);
xor U11481 (N_11481,N_6946,N_6322);
and U11482 (N_11482,N_6068,N_8956);
nand U11483 (N_11483,N_6542,N_5164);
or U11484 (N_11484,N_8227,N_8594);
nor U11485 (N_11485,N_9097,N_6818);
xor U11486 (N_11486,N_6646,N_9357);
nand U11487 (N_11487,N_8378,N_8476);
nand U11488 (N_11488,N_9733,N_7303);
nor U11489 (N_11489,N_8754,N_7842);
xor U11490 (N_11490,N_8772,N_9390);
xor U11491 (N_11491,N_5683,N_6972);
nor U11492 (N_11492,N_8795,N_8979);
xnor U11493 (N_11493,N_9954,N_6868);
xnor U11494 (N_11494,N_6790,N_6231);
nor U11495 (N_11495,N_7460,N_7636);
and U11496 (N_11496,N_9635,N_7715);
and U11497 (N_11497,N_7368,N_7349);
xor U11498 (N_11498,N_5354,N_6841);
or U11499 (N_11499,N_8990,N_8688);
xnor U11500 (N_11500,N_7577,N_5272);
xnor U11501 (N_11501,N_6740,N_9362);
or U11502 (N_11502,N_9001,N_8503);
nor U11503 (N_11503,N_9709,N_6657);
xor U11504 (N_11504,N_7476,N_6441);
nand U11505 (N_11505,N_5464,N_5697);
xnor U11506 (N_11506,N_7867,N_7979);
nand U11507 (N_11507,N_9002,N_7982);
xnor U11508 (N_11508,N_7243,N_9145);
or U11509 (N_11509,N_7528,N_5956);
nor U11510 (N_11510,N_6813,N_9627);
xnor U11511 (N_11511,N_6430,N_8726);
or U11512 (N_11512,N_8621,N_9666);
nand U11513 (N_11513,N_5658,N_6218);
nor U11514 (N_11514,N_9667,N_7620);
nand U11515 (N_11515,N_6722,N_5110);
or U11516 (N_11516,N_5632,N_9575);
or U11517 (N_11517,N_9090,N_5176);
nor U11518 (N_11518,N_8336,N_5165);
and U11519 (N_11519,N_7765,N_7732);
and U11520 (N_11520,N_7326,N_8920);
nand U11521 (N_11521,N_7780,N_5494);
nand U11522 (N_11522,N_7095,N_9327);
xnor U11523 (N_11523,N_6654,N_6451);
nor U11524 (N_11524,N_6190,N_6650);
nor U11525 (N_11525,N_9510,N_6545);
nand U11526 (N_11526,N_5084,N_9858);
xor U11527 (N_11527,N_5023,N_5463);
and U11528 (N_11528,N_8849,N_9036);
and U11529 (N_11529,N_7954,N_6245);
nand U11530 (N_11530,N_6002,N_7038);
nor U11531 (N_11531,N_5135,N_7610);
xor U11532 (N_11532,N_6081,N_5625);
or U11533 (N_11533,N_8037,N_7998);
nand U11534 (N_11534,N_9981,N_6796);
nand U11535 (N_11535,N_8573,N_9318);
xnor U11536 (N_11536,N_8398,N_8505);
nand U11537 (N_11537,N_7507,N_8449);
or U11538 (N_11538,N_5297,N_9902);
and U11539 (N_11539,N_6975,N_9350);
and U11540 (N_11540,N_5858,N_7694);
and U11541 (N_11541,N_6863,N_8973);
nor U11542 (N_11542,N_9356,N_5725);
nor U11543 (N_11543,N_6381,N_8631);
and U11544 (N_11544,N_6378,N_5729);
nor U11545 (N_11545,N_6826,N_7392);
or U11546 (N_11546,N_6854,N_6442);
or U11547 (N_11547,N_7466,N_6461);
nor U11548 (N_11548,N_6774,N_7546);
xor U11549 (N_11549,N_6084,N_6487);
xnor U11550 (N_11550,N_5485,N_5453);
or U11551 (N_11551,N_8739,N_7698);
nand U11552 (N_11552,N_6675,N_6902);
and U11553 (N_11553,N_5698,N_6857);
xor U11554 (N_11554,N_9344,N_8605);
or U11555 (N_11555,N_9264,N_7745);
nor U11556 (N_11556,N_5138,N_8550);
or U11557 (N_11557,N_5975,N_8047);
and U11558 (N_11558,N_5638,N_9398);
and U11559 (N_11559,N_5673,N_7729);
nand U11560 (N_11560,N_5450,N_9334);
nand U11561 (N_11561,N_7722,N_9828);
xnor U11562 (N_11562,N_5305,N_5839);
and U11563 (N_11563,N_9325,N_8154);
nor U11564 (N_11564,N_9781,N_9549);
xnor U11565 (N_11565,N_5528,N_6389);
or U11566 (N_11566,N_7129,N_5557);
nor U11567 (N_11567,N_7767,N_8062);
and U11568 (N_11568,N_9108,N_6325);
xnor U11569 (N_11569,N_9103,N_9223);
nor U11570 (N_11570,N_7083,N_9403);
or U11571 (N_11571,N_7683,N_6425);
nand U11572 (N_11572,N_7601,N_5743);
xor U11573 (N_11573,N_7182,N_8744);
or U11574 (N_11574,N_7668,N_9701);
nor U11575 (N_11575,N_6835,N_9298);
nand U11576 (N_11576,N_8188,N_5357);
and U11577 (N_11577,N_5278,N_5327);
and U11578 (N_11578,N_6651,N_8619);
or U11579 (N_11579,N_7879,N_6073);
nand U11580 (N_11580,N_6649,N_5512);
xor U11581 (N_11581,N_9947,N_6699);
nor U11582 (N_11582,N_6263,N_5889);
xor U11583 (N_11583,N_6548,N_8061);
nor U11584 (N_11584,N_9167,N_9908);
nor U11585 (N_11585,N_9389,N_9536);
nand U11586 (N_11586,N_8141,N_7602);
or U11587 (N_11587,N_8058,N_8275);
and U11588 (N_11588,N_9876,N_8972);
or U11589 (N_11589,N_7481,N_6142);
and U11590 (N_11590,N_6393,N_6858);
and U11591 (N_11591,N_8386,N_9583);
nor U11592 (N_11592,N_9523,N_9054);
nor U11593 (N_11593,N_5761,N_7163);
nand U11594 (N_11594,N_6307,N_8917);
and U11595 (N_11595,N_9420,N_8857);
nor U11596 (N_11596,N_7488,N_9564);
nand U11597 (N_11597,N_8792,N_5570);
xor U11598 (N_11598,N_5651,N_8270);
and U11599 (N_11599,N_5038,N_7192);
nor U11600 (N_11600,N_7257,N_6668);
and U11601 (N_11601,N_8094,N_5225);
nor U11602 (N_11602,N_9758,N_6939);
nor U11603 (N_11603,N_9544,N_7413);
nor U11604 (N_11604,N_9151,N_5269);
or U11605 (N_11605,N_8390,N_6616);
nand U11606 (N_11606,N_6180,N_7865);
nand U11607 (N_11607,N_7570,N_6836);
or U11608 (N_11608,N_7490,N_9782);
xnor U11609 (N_11609,N_9216,N_6278);
or U11610 (N_11610,N_5392,N_5786);
nand U11611 (N_11611,N_7930,N_8607);
and U11612 (N_11612,N_9779,N_5025);
or U11613 (N_11613,N_7189,N_5236);
xnor U11614 (N_11614,N_5799,N_8862);
xor U11615 (N_11615,N_6371,N_6569);
nand U11616 (N_11616,N_8802,N_9976);
nand U11617 (N_11617,N_5892,N_5558);
nand U11618 (N_11618,N_5320,N_9150);
nand U11619 (N_11619,N_9926,N_9771);
and U11620 (N_11620,N_9136,N_6944);
xnor U11621 (N_11621,N_5063,N_5469);
nand U11622 (N_11622,N_5878,N_8451);
and U11623 (N_11623,N_7846,N_5005);
xnor U11624 (N_11624,N_7787,N_7208);
or U11625 (N_11625,N_9037,N_7072);
nand U11626 (N_11626,N_7435,N_5252);
xnor U11627 (N_11627,N_8465,N_5796);
nand U11628 (N_11628,N_9507,N_9820);
or U11629 (N_11629,N_7661,N_7486);
or U11630 (N_11630,N_6904,N_7704);
and U11631 (N_11631,N_5197,N_8564);
xnor U11632 (N_11632,N_7594,N_8055);
or U11633 (N_11633,N_8533,N_9106);
nor U11634 (N_11634,N_8877,N_8685);
or U11635 (N_11635,N_9571,N_7713);
and U11636 (N_11636,N_6133,N_6439);
nor U11637 (N_11637,N_8825,N_5966);
nor U11638 (N_11638,N_7519,N_5820);
or U11639 (N_11639,N_6219,N_8026);
xnor U11640 (N_11640,N_8965,N_9725);
xor U11641 (N_11641,N_5219,N_7484);
or U11642 (N_11642,N_8082,N_9987);
or U11643 (N_11643,N_8266,N_5969);
nand U11644 (N_11644,N_9631,N_9533);
and U11645 (N_11645,N_9414,N_5803);
xor U11646 (N_11646,N_5474,N_6909);
nor U11647 (N_11647,N_6621,N_8648);
nor U11648 (N_11648,N_5888,N_7497);
nor U11649 (N_11649,N_6844,N_9932);
and U11650 (N_11650,N_8705,N_8385);
and U11651 (N_11651,N_5053,N_5587);
nor U11652 (N_11652,N_5376,N_6391);
and U11653 (N_11653,N_5284,N_9559);
nor U11654 (N_11654,N_8675,N_6505);
and U11655 (N_11655,N_7910,N_9123);
and U11656 (N_11656,N_5162,N_5217);
nor U11657 (N_11657,N_7500,N_8872);
nor U11658 (N_11658,N_8178,N_7054);
nand U11659 (N_11659,N_7114,N_9847);
and U11660 (N_11660,N_8834,N_7587);
or U11661 (N_11661,N_6728,N_5069);
xor U11662 (N_11662,N_6592,N_7556);
xnor U11663 (N_11663,N_7260,N_6268);
xor U11664 (N_11664,N_9605,N_5715);
or U11665 (N_11665,N_8672,N_5082);
nor U11666 (N_11666,N_5894,N_9753);
nand U11667 (N_11667,N_6891,N_6198);
nor U11668 (N_11668,N_5459,N_5078);
and U11669 (N_11669,N_6877,N_6759);
xnor U11670 (N_11670,N_9772,N_8771);
xor U11671 (N_11671,N_5871,N_9903);
and U11672 (N_11672,N_7076,N_6850);
nor U11673 (N_11673,N_5007,N_8937);
nand U11674 (N_11674,N_6619,N_6121);
or U11675 (N_11675,N_8558,N_6280);
nand U11676 (N_11676,N_9352,N_5955);
and U11677 (N_11677,N_9248,N_8650);
or U11678 (N_11678,N_9656,N_8083);
or U11679 (N_11679,N_8959,N_7090);
nand U11680 (N_11680,N_9113,N_7946);
nand U11681 (N_11681,N_8702,N_5845);
nand U11682 (N_11682,N_8899,N_9170);
nor U11683 (N_11683,N_6626,N_6007);
nand U11684 (N_11684,N_6262,N_9818);
nand U11685 (N_11685,N_6838,N_6105);
xnor U11686 (N_11686,N_9893,N_8212);
nor U11687 (N_11687,N_9351,N_7789);
xnor U11688 (N_11688,N_8091,N_8856);
xor U11689 (N_11689,N_8491,N_6808);
or U11690 (N_11690,N_8360,N_8217);
and U11691 (N_11691,N_5680,N_5709);
or U11692 (N_11692,N_5822,N_7957);
xor U11693 (N_11693,N_5926,N_5317);
nand U11694 (N_11694,N_7263,N_8189);
and U11695 (N_11695,N_8567,N_7221);
and U11696 (N_11696,N_9283,N_5921);
nand U11697 (N_11697,N_5928,N_7786);
nor U11698 (N_11698,N_9626,N_7711);
xnor U11699 (N_11699,N_5522,N_8419);
and U11700 (N_11700,N_5907,N_7781);
and U11701 (N_11701,N_6936,N_7880);
or U11702 (N_11702,N_8780,N_9532);
or U11703 (N_11703,N_5789,N_7080);
or U11704 (N_11704,N_5568,N_6576);
or U11705 (N_11705,N_8921,N_9724);
xnor U11706 (N_11706,N_8712,N_7783);
or U11707 (N_11707,N_8869,N_5207);
nor U11708 (N_11708,N_5091,N_5744);
or U11709 (N_11709,N_6410,N_6982);
and U11710 (N_11710,N_6855,N_6166);
and U11711 (N_11711,N_9267,N_5585);
or U11712 (N_11712,N_6093,N_7393);
xor U11713 (N_11713,N_5086,N_6598);
or U11714 (N_11714,N_7972,N_8571);
and U11715 (N_11715,N_5224,N_6212);
nor U11716 (N_11716,N_9441,N_8013);
nor U11717 (N_11717,N_8124,N_9886);
nor U11718 (N_11718,N_8763,N_6840);
nand U11719 (N_11719,N_8949,N_9935);
xor U11720 (N_11720,N_5341,N_5083);
xor U11721 (N_11721,N_6935,N_6354);
nor U11722 (N_11722,N_8542,N_8024);
or U11723 (N_11723,N_5647,N_7747);
or U11724 (N_11724,N_9241,N_9916);
and U11725 (N_11725,N_8031,N_8676);
or U11726 (N_11726,N_7463,N_9777);
and U11727 (N_11727,N_5682,N_6330);
nor U11728 (N_11728,N_8770,N_5577);
or U11729 (N_11729,N_9894,N_6929);
and U11730 (N_11730,N_6033,N_9806);
or U11731 (N_11731,N_7753,N_7265);
xor U11732 (N_11732,N_7942,N_9299);
or U11733 (N_11733,N_9194,N_8490);
and U11734 (N_11734,N_9792,N_7468);
nor U11735 (N_11735,N_9808,N_6228);
nand U11736 (N_11736,N_8364,N_8066);
nand U11737 (N_11737,N_5287,N_8707);
nor U11738 (N_11738,N_7458,N_8906);
nor U11739 (N_11739,N_5811,N_7242);
nor U11740 (N_11740,N_7307,N_7364);
and U11741 (N_11741,N_6162,N_9462);
and U11742 (N_11742,N_8549,N_9959);
nand U11743 (N_11743,N_6859,N_9059);
nor U11744 (N_11744,N_8551,N_7066);
or U11745 (N_11745,N_6653,N_7483);
nand U11746 (N_11746,N_5929,N_8329);
nor U11747 (N_11747,N_7015,N_5237);
or U11748 (N_11748,N_5408,N_8297);
and U11749 (N_11749,N_9910,N_5517);
xor U11750 (N_11750,N_7647,N_6016);
xor U11751 (N_11751,N_7442,N_9780);
nand U11752 (N_11752,N_5901,N_6659);
nor U11753 (N_11753,N_9769,N_6488);
and U11754 (N_11754,N_6990,N_5978);
xor U11755 (N_11755,N_5065,N_7778);
nor U11756 (N_11756,N_9650,N_6115);
nor U11757 (N_11757,N_6335,N_9815);
or U11758 (N_11758,N_5367,N_9500);
and U11759 (N_11759,N_9844,N_6465);
nor U11760 (N_11760,N_6415,N_8904);
or U11761 (N_11761,N_8613,N_8612);
nand U11762 (N_11762,N_9757,N_8042);
or U11763 (N_11763,N_7993,N_6712);
xnor U11764 (N_11764,N_5071,N_9336);
nor U11765 (N_11765,N_5181,N_8416);
nand U11766 (N_11766,N_6460,N_8540);
nor U11767 (N_11767,N_6274,N_5388);
or U11768 (N_11768,N_7137,N_8633);
and U11769 (N_11769,N_5551,N_9952);
nand U11770 (N_11770,N_9200,N_9982);
nand U11771 (N_11771,N_8896,N_8884);
xnor U11772 (N_11772,N_7523,N_6636);
or U11773 (N_11773,N_6804,N_7499);
and U11774 (N_11774,N_9748,N_7652);
xor U11775 (N_11775,N_7304,N_5248);
or U11776 (N_11776,N_9570,N_9694);
or U11777 (N_11777,N_6805,N_8016);
nand U11778 (N_11778,N_6341,N_5033);
and U11779 (N_11779,N_7438,N_7153);
and U11780 (N_11780,N_6358,N_5466);
nand U11781 (N_11781,N_9339,N_6645);
nor U11782 (N_11782,N_8264,N_6525);
or U11783 (N_11783,N_6362,N_7634);
nand U11784 (N_11784,N_9739,N_9222);
nor U11785 (N_11785,N_5800,N_9588);
nor U11786 (N_11786,N_6721,N_9133);
nor U11787 (N_11787,N_7342,N_8933);
nor U11788 (N_11788,N_5533,N_6464);
xor U11789 (N_11789,N_6672,N_7399);
nor U11790 (N_11790,N_8820,N_9427);
nand U11791 (N_11791,N_7011,N_8996);
xnor U11792 (N_11792,N_8492,N_7755);
or U11793 (N_11793,N_8997,N_5313);
and U11794 (N_11794,N_8469,N_8156);
xor U11795 (N_11795,N_5429,N_5703);
xnor U11796 (N_11796,N_8209,N_6392);
nor U11797 (N_11797,N_7935,N_7121);
or U11798 (N_11798,N_6898,N_9157);
nor U11799 (N_11799,N_6574,N_5502);
or U11800 (N_11800,N_5395,N_7759);
nor U11801 (N_11801,N_9295,N_9912);
and U11802 (N_11802,N_7108,N_9798);
nand U11803 (N_11803,N_5608,N_8413);
nor U11804 (N_11804,N_6022,N_5183);
nor U11805 (N_11805,N_8201,N_6945);
or U11806 (N_11806,N_5837,N_5662);
nor U11807 (N_11807,N_5671,N_7405);
or U11808 (N_11808,N_7649,N_5220);
and U11809 (N_11809,N_5595,N_5873);
or U11810 (N_11810,N_7600,N_7983);
nor U11811 (N_11811,N_8637,N_6667);
nor U11812 (N_11812,N_5925,N_9217);
xor U11813 (N_11813,N_6771,N_5159);
or U11814 (N_11814,N_8168,N_9135);
nor U11815 (N_11815,N_8001,N_7987);
nor U11816 (N_11816,N_9887,N_5752);
nor U11817 (N_11817,N_8125,N_8616);
nor U11818 (N_11818,N_9839,N_7171);
nor U11819 (N_11819,N_9319,N_9199);
xor U11820 (N_11820,N_5230,N_8680);
or U11821 (N_11821,N_9501,N_8150);
nor U11822 (N_11822,N_6011,N_7645);
nor U11823 (N_11823,N_9948,N_5076);
nor U11824 (N_11824,N_7381,N_5583);
or U11825 (N_11825,N_9702,N_8864);
nor U11826 (N_11826,N_5415,N_7811);
or U11827 (N_11827,N_5262,N_7453);
nand U11828 (N_11828,N_6752,N_6337);
xor U11829 (N_11829,N_5566,N_7626);
xor U11830 (N_11830,N_7372,N_7345);
and U11831 (N_11831,N_9857,N_7967);
xnor U11832 (N_11832,N_7992,N_6290);
nor U11833 (N_11833,N_9016,N_9092);
and U11834 (N_11834,N_9674,N_7138);
xnor U11835 (N_11835,N_8276,N_7141);
nand U11836 (N_11836,N_9845,N_7532);
nor U11837 (N_11837,N_7770,N_8598);
or U11838 (N_11838,N_6919,N_6196);
xnor U11839 (N_11839,N_8609,N_5437);
or U11840 (N_11840,N_8814,N_6508);
or U11841 (N_11841,N_6047,N_6860);
xor U11842 (N_11842,N_6524,N_9516);
or U11843 (N_11843,N_9877,N_6556);
nand U11844 (N_11844,N_8922,N_8015);
xor U11845 (N_11845,N_7152,N_6785);
and U11846 (N_11846,N_9829,N_5992);
nand U11847 (N_11847,N_6777,N_9732);
xor U11848 (N_11848,N_8608,N_9599);
nand U11849 (N_11849,N_9968,N_8149);
or U11850 (N_11850,N_7617,N_7388);
and U11851 (N_11851,N_5622,N_9126);
and U11852 (N_11852,N_8342,N_6966);
xor U11853 (N_11853,N_6767,N_6469);
or U11854 (N_11854,N_8406,N_6175);
or U11855 (N_11855,N_5994,N_8251);
or U11856 (N_11856,N_5895,N_7409);
or U11857 (N_11857,N_7330,N_6582);
xor U11858 (N_11858,N_6209,N_5098);
xnor U11859 (N_11859,N_9159,N_8216);
and U11860 (N_11860,N_7810,N_5468);
nor U11861 (N_11861,N_6493,N_5008);
or U11862 (N_11862,N_5416,N_7904);
xor U11863 (N_11863,N_7112,N_5035);
nor U11864 (N_11864,N_5971,N_8640);
and U11865 (N_11865,N_5814,N_7504);
and U11866 (N_11866,N_6691,N_6748);
nor U11867 (N_11867,N_6980,N_7660);
or U11868 (N_11868,N_5345,N_7843);
and U11869 (N_11869,N_5862,N_6159);
nor U11870 (N_11870,N_6669,N_7472);
and U11871 (N_11871,N_5360,N_8483);
nor U11872 (N_11872,N_9051,N_7675);
xnor U11873 (N_11873,N_6893,N_6253);
and U11874 (N_11874,N_5776,N_7891);
or U11875 (N_11875,N_8779,N_7888);
xor U11876 (N_11876,N_7762,N_5195);
nor U11877 (N_11877,N_5097,N_5228);
nor U11878 (N_11878,N_5726,N_8234);
nand U11879 (N_11879,N_8958,N_9735);
xnor U11880 (N_11880,N_6333,N_5251);
nand U11881 (N_11881,N_7197,N_9355);
or U11882 (N_11882,N_9854,N_6009);
xor U11883 (N_11883,N_8741,N_9671);
and U11884 (N_11884,N_6064,N_5140);
or U11885 (N_11885,N_8749,N_8121);
or U11886 (N_11886,N_8696,N_9070);
nand U11887 (N_11887,N_6259,N_8968);
or U11888 (N_11888,N_6824,N_6039);
and U11889 (N_11889,N_8076,N_8166);
or U11890 (N_11890,N_8837,N_5180);
and U11891 (N_11891,N_5534,N_5947);
and U11892 (N_11892,N_6510,N_6564);
or U11893 (N_11893,N_7609,N_6099);
or U11894 (N_11894,N_8279,N_5290);
nor U11895 (N_11895,N_9990,N_6682);
or U11896 (N_11896,N_7444,N_7306);
or U11897 (N_11897,N_8782,N_6853);
xor U11898 (N_11898,N_6871,N_8461);
xnor U11899 (N_11899,N_8801,N_7832);
xnor U11900 (N_11900,N_8603,N_8293);
and U11901 (N_11901,N_6293,N_7103);
xnor U11902 (N_11902,N_8828,N_7366);
or U11903 (N_11903,N_5451,N_5569);
xor U11904 (N_11904,N_8256,N_7252);
or U11905 (N_11905,N_5749,N_5319);
nor U11906 (N_11906,N_5644,N_5056);
nand U11907 (N_11907,N_7266,N_9342);
or U11908 (N_11908,N_7572,N_7726);
xor U11909 (N_11909,N_8281,N_5756);
or U11910 (N_11910,N_6491,N_7913);
and U11911 (N_11911,N_9936,N_8339);
or U11912 (N_11912,N_8236,N_8842);
and U11913 (N_11913,N_6049,N_5390);
and U11914 (N_11914,N_8052,N_9993);
and U11915 (N_11915,N_7184,N_8531);
xnor U11916 (N_11916,N_8219,N_8314);
and U11917 (N_11917,N_5704,N_6761);
or U11918 (N_11918,N_7454,N_6357);
nand U11919 (N_11919,N_6254,N_7829);
xor U11920 (N_11920,N_9172,N_8196);
or U11921 (N_11921,N_9481,N_9712);
or U11922 (N_11922,N_6143,N_6474);
xor U11923 (N_11923,N_5759,N_7664);
nor U11924 (N_11924,N_5910,N_7670);
nor U11925 (N_11925,N_8635,N_8192);
nor U11926 (N_11926,N_8901,N_6315);
or U11927 (N_11927,N_6287,N_8489);
and U11928 (N_11928,N_7170,N_7994);
xor U11929 (N_11929,N_8162,N_6277);
and U11930 (N_11930,N_7455,N_8827);
or U11931 (N_11931,N_6359,N_9469);
or U11932 (N_11932,N_7686,N_7885);
or U11933 (N_11933,N_7420,N_6082);
or U11934 (N_11934,N_6807,N_9737);
nor U11935 (N_11935,N_7909,N_6298);
or U11936 (N_11936,N_7814,N_6169);
or U11937 (N_11937,N_5990,N_9545);
and U11938 (N_11938,N_9213,N_9034);
xor U11939 (N_11939,N_7130,N_7693);
xnor U11940 (N_11940,N_7370,N_6017);
nand U11941 (N_11941,N_7354,N_6750);
nand U11942 (N_11942,N_7202,N_8967);
nor U11943 (N_11943,N_9843,N_5186);
or U11944 (N_11944,N_5449,N_7545);
and U11945 (N_11945,N_5760,N_8185);
xnor U11946 (N_11946,N_5691,N_5556);
xor U11947 (N_11947,N_5635,N_5856);
or U11948 (N_11948,N_7362,N_9595);
nor U11949 (N_11949,N_7684,N_6374);
and U11950 (N_11950,N_5968,N_6827);
and U11951 (N_11951,N_5444,N_7427);
xnor U11952 (N_11952,N_8868,N_8776);
and U11953 (N_11953,N_6141,N_9586);
and U11954 (N_11954,N_6745,N_8653);
xnor U11955 (N_11955,N_6083,N_7606);
nand U11956 (N_11956,N_5728,N_7963);
nand U11957 (N_11957,N_8200,N_8808);
and U11958 (N_11958,N_5275,N_8006);
xor U11959 (N_11959,N_6106,N_6113);
xor U11960 (N_11960,N_9741,N_6024);
and U11961 (N_11961,N_9760,N_8312);
and U11962 (N_11962,N_9869,N_8127);
xor U11963 (N_11963,N_8863,N_7669);
nor U11964 (N_11964,N_6931,N_5659);
xor U11965 (N_11965,N_8184,N_5514);
nand U11966 (N_11966,N_7043,N_6174);
nand U11967 (N_11967,N_8657,N_9369);
nor U11968 (N_11968,N_8766,N_9766);
nand U11969 (N_11969,N_6874,N_6784);
or U11970 (N_11970,N_6225,N_8425);
xnor U11971 (N_11971,N_8034,N_7582);
or U11972 (N_11972,N_8048,N_7580);
or U11973 (N_11973,N_6708,N_9943);
or U11974 (N_11974,N_8448,N_7248);
xnor U11975 (N_11975,N_9451,N_8832);
or U11976 (N_11976,N_8698,N_9879);
and U11977 (N_11977,N_9672,N_9239);
xor U11978 (N_11978,N_6943,N_7440);
or U11979 (N_11979,N_8556,N_5590);
or U11980 (N_11980,N_8074,N_8257);
and U11981 (N_11981,N_6502,N_6210);
or U11982 (N_11982,N_7292,N_6816);
nand U11983 (N_11983,N_5563,N_8546);
nand U11984 (N_11984,N_7648,N_5986);
and U11985 (N_11985,N_9062,N_6557);
or U11986 (N_11986,N_6041,N_8998);
and U11987 (N_11987,N_8288,N_6182);
and U11988 (N_11988,N_8017,N_9069);
or U11989 (N_11989,N_8272,N_7691);
and U11990 (N_11990,N_7583,N_7249);
or U11991 (N_11991,N_8320,N_5842);
nor U11992 (N_11992,N_8112,N_5919);
nand U11993 (N_11993,N_9166,N_8822);
nand U11994 (N_11994,N_9821,N_7513);
or U11995 (N_11995,N_7142,N_5979);
nand U11996 (N_11996,N_9979,N_8522);
xnor U11997 (N_11997,N_5713,N_5790);
or U11998 (N_11998,N_9453,N_9326);
xnor U11999 (N_11999,N_9387,N_6905);
or U12000 (N_12000,N_6353,N_5105);
xor U12001 (N_12001,N_7776,N_8666);
or U12002 (N_12002,N_8466,N_8408);
nand U12003 (N_12003,N_9021,N_5066);
or U12004 (N_12004,N_8375,N_6744);
or U12005 (N_12005,N_8165,N_8510);
and U12006 (N_12006,N_7862,N_7743);
or U12007 (N_12007,N_5011,N_9378);
or U12008 (N_12008,N_9413,N_8660);
and U12009 (N_12009,N_9641,N_9669);
and U12010 (N_12010,N_8824,N_7334);
nand U12011 (N_12011,N_8918,N_8481);
nand U12012 (N_12012,N_9978,N_5119);
and U12013 (N_12013,N_9071,N_6895);
nor U12014 (N_12014,N_7569,N_6575);
or U12015 (N_12015,N_8646,N_8403);
and U12016 (N_12016,N_8511,N_7336);
or U12017 (N_12017,N_8478,N_7890);
xnor U12018 (N_12018,N_9864,N_6901);
xor U12019 (N_12019,N_6241,N_8350);
xor U12020 (N_12020,N_7629,N_6684);
and U12021 (N_12021,N_9131,N_8747);
nand U12022 (N_12022,N_7873,N_9174);
or U12023 (N_12023,N_7089,N_9418);
nand U12024 (N_12024,N_6412,N_7690);
xnor U12025 (N_12025,N_8187,N_9852);
nand U12026 (N_12026,N_9162,N_7761);
nand U12027 (N_12027,N_9504,N_8512);
xor U12028 (N_12028,N_6233,N_6591);
xnor U12029 (N_12029,N_9633,N_8277);
or U12030 (N_12030,N_7383,N_9707);
and U12031 (N_12031,N_9161,N_6191);
or U12032 (N_12032,N_8599,N_5747);
nand U12033 (N_12033,N_5323,N_9377);
or U12034 (N_12034,N_7329,N_9024);
nand U12035 (N_12035,N_8800,N_7049);
nor U12036 (N_12036,N_6571,N_6495);
nand U12037 (N_12037,N_8721,N_6185);
or U12038 (N_12038,N_7492,N_7706);
xor U12039 (N_12039,N_8529,N_9793);
nor U12040 (N_12040,N_8382,N_6387);
nor U12041 (N_12041,N_6589,N_6069);
xor U12042 (N_12042,N_8805,N_5030);
or U12043 (N_12043,N_5128,N_8283);
xnor U12044 (N_12044,N_8485,N_7773);
xor U12045 (N_12045,N_7315,N_5657);
or U12046 (N_12046,N_7827,N_8713);
or U12047 (N_12047,N_5681,N_7790);
xnor U12048 (N_12048,N_6116,N_6701);
xor U12049 (N_12049,N_9483,N_5880);
and U12050 (N_12050,N_7938,N_8701);
or U12051 (N_12051,N_6794,N_9497);
nor U12052 (N_12052,N_6749,N_6475);
and U12053 (N_12053,N_7883,N_6456);
nor U12054 (N_12054,N_5835,N_8379);
or U12055 (N_12055,N_7143,N_8623);
nand U12056 (N_12056,N_8041,N_9985);
and U12057 (N_12057,N_8803,N_5604);
nor U12058 (N_12058,N_5256,N_5797);
xor U12059 (N_12059,N_9514,N_7574);
and U12060 (N_12060,N_7724,N_9388);
nand U12061 (N_12061,N_6304,N_5335);
xor U12062 (N_12062,N_6602,N_6480);
and U12063 (N_12063,N_9231,N_8720);
or U12064 (N_12064,N_5161,N_5555);
or U12065 (N_12065,N_8647,N_9749);
xor U12066 (N_12066,N_6864,N_9271);
nor U12067 (N_12067,N_7269,N_8131);
xnor U12068 (N_12068,N_5643,N_7640);
or U12069 (N_12069,N_9939,N_6782);
or U12070 (N_12070,N_7092,N_6594);
or U12071 (N_12071,N_6663,N_5304);
xor U12072 (N_12072,N_5828,N_7816);
nand U12073 (N_12073,N_5935,N_7421);
or U12074 (N_12074,N_9033,N_6227);
nor U12075 (N_12075,N_9950,N_9662);
xor U12076 (N_12076,N_9591,N_5737);
or U12077 (N_12077,N_6892,N_7976);
xnor U12078 (N_12078,N_6097,N_5009);
nand U12079 (N_12079,N_5381,N_6207);
xnor U12080 (N_12080,N_8833,N_5102);
nand U12081 (N_12081,N_6088,N_5266);
and U12082 (N_12082,N_7503,N_9581);
xnor U12083 (N_12083,N_9768,N_8325);
nor U12084 (N_12084,N_9528,N_7135);
or U12085 (N_12085,N_5113,N_8790);
nand U12086 (N_12086,N_9698,N_6072);
nor U12087 (N_12087,N_8313,N_9225);
nor U12088 (N_12088,N_5016,N_9611);
nor U12089 (N_12089,N_7854,N_9429);
or U12090 (N_12090,N_5742,N_7852);
xor U12091 (N_12091,N_5330,N_7305);
and U12092 (N_12092,N_8748,N_7757);
or U12093 (N_12093,N_7707,N_5544);
or U12094 (N_12094,N_7899,N_8347);
and U12095 (N_12095,N_7044,N_7286);
xnor U12096 (N_12096,N_7807,N_5154);
xor U12097 (N_12097,N_9496,N_6249);
xnor U12098 (N_12098,N_8909,N_6938);
nand U12099 (N_12099,N_9770,N_8179);
or U12100 (N_12100,N_5158,N_5718);
xnor U12101 (N_12101,N_8796,N_8525);
nand U12102 (N_12102,N_9983,N_8644);
or U12103 (N_12103,N_6499,N_6054);
or U12104 (N_12104,N_7116,N_6521);
or U12105 (N_12105,N_6625,N_5819);
xor U12106 (N_12106,N_7518,N_8615);
nor U12107 (N_12107,N_6473,N_7270);
xor U12108 (N_12108,N_9964,N_8963);
nand U12109 (N_12109,N_7643,N_7225);
and U12110 (N_12110,N_7779,N_5817);
xor U12111 (N_12111,N_6927,N_6638);
xnor U12112 (N_12112,N_6655,N_5405);
nor U12113 (N_12113,N_6969,N_9872);
nand U12114 (N_12114,N_9211,N_7450);
or U12115 (N_12115,N_9183,N_7516);
nand U12116 (N_12116,N_9568,N_6660);
and U12117 (N_12117,N_6965,N_8604);
or U12118 (N_12118,N_8516,N_7235);
nor U12119 (N_12119,N_7672,N_8823);
xor U12120 (N_12120,N_7193,N_6942);
nor U12121 (N_12121,N_9927,N_7635);
or U12122 (N_12122,N_5020,N_5369);
xor U12123 (N_12123,N_8870,N_5019);
and U12124 (N_12124,N_9960,N_6025);
or U12125 (N_12125,N_6366,N_6214);
nor U12126 (N_12126,N_5717,N_7956);
and U12127 (N_12127,N_5479,N_7613);
or U12128 (N_12128,N_9680,N_8155);
nand U12129 (N_12129,N_9284,N_7679);
xor U12130 (N_12130,N_6399,N_8077);
and U12131 (N_12131,N_8993,N_9196);
xnor U12132 (N_12132,N_7052,N_6463);
xor U12133 (N_12133,N_5201,N_8590);
or U12134 (N_12134,N_5815,N_7937);
xnor U12135 (N_12135,N_7598,N_5734);
or U12136 (N_12136,N_8028,N_5550);
and U12137 (N_12137,N_5156,N_7067);
or U12138 (N_12138,N_9718,N_6171);
nor U12139 (N_12139,N_5738,N_9013);
or U12140 (N_12140,N_7681,N_9842);
and U12141 (N_12141,N_6537,N_7058);
and U12142 (N_12142,N_8086,N_7045);
and U12143 (N_12143,N_7674,N_8752);
and U12144 (N_12144,N_5785,N_7253);
xor U12145 (N_12145,N_9921,N_8617);
and U12146 (N_12146,N_8366,N_5052);
or U12147 (N_12147,N_9513,N_5918);
or U12148 (N_12148,N_5900,N_7991);
xor U12149 (N_12149,N_8853,N_9840);
xnor U12150 (N_12150,N_8243,N_5712);
xor U12151 (N_12151,N_9316,N_8170);
xnor U12152 (N_12152,N_7297,N_9551);
and U12153 (N_12153,N_9895,N_5940);
nand U12154 (N_12154,N_9364,N_5488);
nand U12155 (N_12155,N_7169,N_5080);
and U12156 (N_12156,N_6363,N_9816);
nor U12157 (N_12157,N_9608,N_7451);
and U12158 (N_12158,N_8665,N_5017);
and U12159 (N_12159,N_5893,N_9914);
xor U12160 (N_12160,N_6849,N_6380);
or U12161 (N_12161,N_7173,N_8368);
and U12162 (N_12162,N_6680,N_6685);
and U12163 (N_12163,N_5523,N_8936);
xnor U12164 (N_12164,N_5753,N_5687);
and U12165 (N_12165,N_6820,N_6089);
or U12166 (N_12166,N_5337,N_8119);
xor U12167 (N_12167,N_8214,N_8582);
or U12168 (N_12168,N_5061,N_6360);
and U12169 (N_12169,N_5890,N_5706);
xnor U12170 (N_12170,N_6924,N_7390);
nand U12171 (N_12171,N_6447,N_8063);
or U12172 (N_12172,N_6271,N_6707);
or U12173 (N_12173,N_9708,N_8534);
xor U12174 (N_12174,N_9795,N_6037);
and U12175 (N_12175,N_5663,N_9008);
nor U12176 (N_12176,N_6197,N_7057);
nor U12177 (N_12177,N_7567,N_7644);
nand U12178 (N_12178,N_6297,N_9395);
and U12179 (N_12179,N_6424,N_7172);
nand U12180 (N_12180,N_5004,N_9550);
nor U12181 (N_12181,N_6603,N_7744);
nand U12182 (N_12182,N_7115,N_5396);
nand U12183 (N_12183,N_7728,N_6104);
and U12184 (N_12184,N_7897,N_6928);
xnor U12185 (N_12185,N_7322,N_9706);
nor U12186 (N_12186,N_5087,N_9385);
nand U12187 (N_12187,N_5702,N_9080);
xor U12188 (N_12188,N_7502,N_5768);
nor U12189 (N_12189,N_7906,N_7133);
nand U12190 (N_12190,N_9084,N_7069);
or U12191 (N_12191,N_5257,N_5413);
or U12192 (N_12192,N_9260,N_5240);
and U12193 (N_12193,N_9597,N_5072);
or U12194 (N_12194,N_8300,N_8142);
or U12195 (N_12195,N_8689,N_7369);
and U12196 (N_12196,N_5619,N_9209);
or U12197 (N_12197,N_5755,N_7689);
xnor U12198 (N_12198,N_7815,N_8245);
nand U12199 (N_12199,N_9421,N_9347);
nand U12200 (N_12200,N_8175,N_5239);
nand U12201 (N_12201,N_5645,N_6334);
and U12202 (N_12202,N_9138,N_9572);
or U12203 (N_12203,N_5491,N_8287);
nor U12204 (N_12204,N_6988,N_5032);
or U12205 (N_12205,N_7494,N_6446);
or U12206 (N_12206,N_5391,N_6204);
and U12207 (N_12207,N_9940,N_5933);
nand U12208 (N_12208,N_8298,N_8081);
nor U12209 (N_12209,N_6666,N_8620);
and U12210 (N_12210,N_9634,N_6091);
xnor U12211 (N_12211,N_9911,N_7579);
or U12212 (N_12212,N_7380,N_6622);
xnor U12213 (N_12213,N_9875,N_8645);
nor U12214 (N_12214,N_9529,N_7769);
nand U12215 (N_12215,N_7241,N_7016);
nand U12216 (N_12216,N_5603,N_5283);
nand U12217 (N_12217,N_6265,N_9865);
and U12218 (N_12218,N_8798,N_9391);
nand U12219 (N_12219,N_9093,N_8204);
nor U12220 (N_12220,N_6918,N_7316);
or U12221 (N_12221,N_6678,N_9372);
nor U12222 (N_12222,N_7534,N_6954);
xnor U12223 (N_12223,N_7768,N_7213);
xor U12224 (N_12224,N_5782,N_7032);
or U12225 (N_12225,N_7379,N_8133);
xor U12226 (N_12226,N_9101,N_5591);
xnor U12227 (N_12227,N_6026,N_9230);
nand U12228 (N_12228,N_6445,N_8559);
xor U12229 (N_12229,N_5905,N_9119);
nor U12230 (N_12230,N_6550,N_7294);
and U12231 (N_12231,N_9374,N_9214);
nand U12232 (N_12232,N_7280,N_9359);
xnor U12233 (N_12233,N_7048,N_7535);
and U12234 (N_12234,N_9517,N_7777);
nand U12235 (N_12235,N_8018,N_7941);
or U12236 (N_12236,N_5279,N_9937);
and U12237 (N_12237,N_7901,N_5850);
or U12238 (N_12238,N_7839,N_9313);
nor U12239 (N_12239,N_6189,N_7505);
nor U12240 (N_12240,N_5964,N_6344);
nand U12241 (N_12241,N_7276,N_9147);
or U12242 (N_12242,N_7228,N_7281);
and U12243 (N_12243,N_7106,N_5508);
and U12244 (N_12244,N_6251,N_8858);
nor U12245 (N_12245,N_7222,N_5111);
and U12246 (N_12246,N_9562,N_7760);
nand U12247 (N_12247,N_9251,N_5173);
nor U12248 (N_12248,N_8468,N_8248);
and U12249 (N_12249,N_9408,N_6967);
or U12250 (N_12250,N_5109,N_6163);
nor U12251 (N_12251,N_9433,N_6038);
and U12252 (N_12252,N_5421,N_7547);
xor U12253 (N_12253,N_8969,N_6579);
nor U12254 (N_12254,N_5909,N_9232);
nor U12255 (N_12255,N_9153,N_7861);
xnor U12256 (N_12256,N_7296,N_8981);
and U12257 (N_12257,N_9030,N_9618);
and U12258 (N_12258,N_8799,N_5863);
nor U12259 (N_12259,N_5003,N_8428);
xnor U12260 (N_12260,N_9402,N_9201);
or U12261 (N_12261,N_7524,N_6103);
nand U12262 (N_12262,N_9525,N_6273);
nor U12263 (N_12263,N_5936,N_7123);
and U12264 (N_12264,N_5343,N_9212);
or U12265 (N_12265,N_7666,N_5524);
nand U12266 (N_12266,N_5430,N_8982);
xnor U12267 (N_12267,N_8677,N_9007);
nand U12268 (N_12268,N_8504,N_9751);
and U12269 (N_12269,N_9955,N_5559);
nor U12270 (N_12270,N_6109,N_5438);
and U12271 (N_12271,N_6494,N_6770);
xor U12272 (N_12272,N_6050,N_6795);
nor U12273 (N_12273,N_9309,N_9331);
and U12274 (N_12274,N_8374,N_8405);
nand U12275 (N_12275,N_7215,N_9436);
or U12276 (N_12276,N_5938,N_8273);
and U12277 (N_12277,N_6310,N_9889);
and U12278 (N_12278,N_7764,N_9132);
and U12279 (N_12279,N_7981,N_7029);
nor U12280 (N_12280,N_7678,N_8846);
xnor U12281 (N_12281,N_6995,N_8487);
nor U12282 (N_12282,N_9565,N_8317);
and U12283 (N_12283,N_8237,N_9546);
and U12284 (N_12284,N_9841,N_7914);
xnor U12285 (N_12285,N_9179,N_9091);
and U12286 (N_12286,N_8809,N_9933);
or U12287 (N_12287,N_5149,N_7183);
or U12288 (N_12288,N_7709,N_6269);
xor U12289 (N_12289,N_8044,N_6887);
or U12290 (N_12290,N_6531,N_8355);
xnor U12291 (N_12291,N_6455,N_5398);
xor U12292 (N_12292,N_8367,N_6724);
nor U12293 (N_12293,N_8989,N_9696);
or U12294 (N_12294,N_5521,N_7210);
nor U12295 (N_12295,N_7659,N_9628);
nor U12296 (N_12296,N_6596,N_9182);
nor U12297 (N_12297,N_7608,N_8836);
nor U12298 (N_12298,N_7558,N_8069);
nor U12299 (N_12299,N_9317,N_8794);
or U12300 (N_12300,N_5235,N_7035);
and U12301 (N_12301,N_7960,N_5700);
nor U12302 (N_12302,N_7059,N_7530);
nor U12303 (N_12303,N_6544,N_8289);
xnor U12304 (N_12304,N_7754,N_6955);
nand U12305 (N_12305,N_6610,N_7510);
nand U12306 (N_12306,N_9885,N_9687);
and U12307 (N_12307,N_8089,N_8553);
xnor U12308 (N_12308,N_5998,N_6732);
nor U12309 (N_12309,N_6851,N_9969);
xnor U12310 (N_12310,N_5175,N_5724);
xor U12311 (N_12311,N_7549,N_6652);
nor U12312 (N_12312,N_8678,N_8578);
nor U12313 (N_12313,N_8786,N_6243);
xor U12314 (N_12314,N_6727,N_6878);
or U12315 (N_12315,N_5356,N_5480);
nand U12316 (N_12316,N_9224,N_9431);
or U12317 (N_12317,N_5222,N_5329);
nand U12318 (N_12318,N_8152,N_6129);
xor U12319 (N_12319,N_7351,N_6200);
nand U12320 (N_12320,N_5970,N_6486);
or U12321 (N_12321,N_9996,N_8351);
xor U12322 (N_12322,N_6264,N_5950);
nor U12323 (N_12323,N_9677,N_8597);
xor U12324 (N_12324,N_6756,N_9287);
nor U12325 (N_12325,N_9017,N_8600);
or U12326 (N_12326,N_9275,N_5887);
or U12327 (N_12327,N_5848,N_7021);
xnor U12328 (N_12328,N_8410,N_9946);
nand U12329 (N_12329,N_8817,N_6635);
and U12330 (N_12330,N_9480,N_5163);
or U12331 (N_12331,N_9909,N_6704);
nand U12332 (N_12332,N_5101,N_5456);
nand U12333 (N_12333,N_7881,N_9025);
nor U12334 (N_12334,N_6554,N_7857);
or U12335 (N_12335,N_9676,N_9901);
nand U12336 (N_12336,N_5478,N_6731);
nand U12337 (N_12337,N_9074,N_7136);
xnor U12338 (N_12338,N_9752,N_8167);
and U12339 (N_12339,N_6126,N_8812);
nor U12340 (N_12340,N_7350,N_9778);
xnor U12341 (N_12341,N_6279,N_8010);
and U12342 (N_12342,N_5118,N_9924);
or U12343 (N_12343,N_9930,N_8638);
nand U12344 (N_12344,N_5705,N_8304);
xnor U12345 (N_12345,N_5286,N_6301);
nand U12346 (N_12346,N_9263,N_8767);
nand U12347 (N_12347,N_8231,N_7167);
nand U12348 (N_12348,N_8411,N_8577);
xnor U12349 (N_12349,N_5099,N_6345);
and U12350 (N_12350,N_7282,N_6769);
nor U12351 (N_12351,N_5037,N_8249);
and U12352 (N_12352,N_7359,N_8190);
or U12353 (N_12353,N_6515,N_8883);
nand U12354 (N_12354,N_7008,N_5088);
or U12355 (N_12355,N_5771,N_8691);
nand U12356 (N_12356,N_8654,N_8022);
nor U12357 (N_12357,N_5454,N_7299);
nor U12358 (N_12358,N_6003,N_6053);
nand U12359 (N_12359,N_8894,N_8146);
nand U12360 (N_12360,N_6479,N_7986);
nand U12361 (N_12361,N_5679,N_8679);
or U12362 (N_12362,N_6478,N_6468);
nand U12363 (N_12363,N_9085,N_9208);
nand U12364 (N_12364,N_5402,N_5026);
nor U12365 (N_12365,N_7014,N_9623);
xnor U12366 (N_12366,N_8088,N_8960);
and U12367 (N_12367,N_9745,N_6459);
or U12368 (N_12368,N_5015,N_6713);
and U12369 (N_12369,N_5231,N_9619);
and U12370 (N_12370,N_6530,N_8139);
xor U12371 (N_12371,N_5137,N_8757);
xnor U12372 (N_12372,N_9835,N_8110);
or U12373 (N_12373,N_6199,N_8087);
nor U12374 (N_12374,N_5439,N_5567);
or U12375 (N_12375,N_7805,N_7845);
nand U12376 (N_12376,N_5316,N_7856);
xnor U12377 (N_12377,N_5250,N_9285);
nand U12378 (N_12378,N_8987,N_7489);
or U12379 (N_12379,N_9058,N_7521);
or U12380 (N_12380,N_5572,N_5050);
xnor U12381 (N_12381,N_6350,N_7168);
nor U12382 (N_12382,N_7671,N_8821);
nor U12383 (N_12383,N_7335,N_5843);
and U12384 (N_12384,N_6609,N_7195);
and U12385 (N_12385,N_6257,N_7367);
nand U12386 (N_12386,N_8994,N_5853);
or U12387 (N_12387,N_7898,N_8396);
xnor U12388 (N_12388,N_7919,N_7628);
nand U12389 (N_12389,N_9004,N_6559);
or U12390 (N_12390,N_9056,N_8147);
or U12391 (N_12391,N_9592,N_9435);
xnor U12392 (N_12392,N_6985,N_5160);
xnor U12393 (N_12393,N_5467,N_8829);
or U12394 (N_12394,N_9075,N_8000);
nand U12395 (N_12395,N_7162,N_9235);
nand U12396 (N_12396,N_9055,N_8738);
or U12397 (N_12397,N_9941,N_9358);
xnor U12398 (N_12398,N_6516,N_8051);
nor U12399 (N_12399,N_9278,N_6620);
xnor U12400 (N_12400,N_9870,N_9944);
nand U12401 (N_12401,N_8507,N_5133);
nor U12402 (N_12402,N_9970,N_5660);
nor U12403 (N_12403,N_6983,N_8180);
nand U12404 (N_12404,N_7611,N_5194);
nand U12405 (N_12405,N_7959,N_6139);
nand U12406 (N_12406,N_8860,N_7198);
and U12407 (N_12407,N_9478,N_8508);
nand U12408 (N_12408,N_5385,N_7272);
nor U12409 (N_12409,N_6607,N_7564);
nor U12410 (N_12410,N_5414,N_9082);
nand U12411 (N_12411,N_7031,N_5731);
nor U12412 (N_12412,N_8627,N_5506);
nand U12413 (N_12413,N_9188,N_5565);
or U12414 (N_12414,N_9589,N_5650);
and U12415 (N_12415,N_7795,N_8328);
or U12416 (N_12416,N_9404,N_5943);
and U12417 (N_12417,N_7710,N_5741);
nand U12418 (N_12418,N_9472,N_8446);
nor U12419 (N_12419,N_5991,N_7774);
xor U12420 (N_12420,N_7604,N_9880);
xor U12421 (N_12421,N_6349,N_5146);
and U12422 (N_12422,N_5062,N_8432);
nor U12423 (N_12423,N_5233,N_9312);
xnor U12424 (N_12424,N_7482,N_9679);
nor U12425 (N_12425,N_9734,N_6833);
nand U12426 (N_12426,N_9146,N_5255);
or U12427 (N_12427,N_7737,N_5941);
and U12428 (N_12428,N_6492,N_8193);
and U12429 (N_12429,N_7293,N_8592);
xnor U12430 (N_12430,N_7622,N_5696);
nand U12431 (N_12431,N_5093,N_5300);
or U12432 (N_12432,N_5689,N_7812);
xor U12433 (N_12433,N_9904,N_9493);
xor U12434 (N_12434,N_9728,N_5582);
or U12435 (N_12435,N_9809,N_6811);
xor U12436 (N_12436,N_6062,N_8174);
or U12437 (N_12437,N_6244,N_8090);
nor U12438 (N_12438,N_5436,N_6501);
and U12439 (N_12439,N_7692,N_6922);
nand U12440 (N_12440,N_6063,N_5547);
or U12441 (N_12441,N_7840,N_7437);
and U12442 (N_12442,N_6215,N_5597);
xor U12443 (N_12443,N_7055,N_7312);
xnor U12444 (N_12444,N_6056,N_5849);
nand U12445 (N_12445,N_5340,N_8363);
and U12446 (N_12446,N_9668,N_9963);
and U12447 (N_12447,N_8423,N_9111);
xnor U12448 (N_12448,N_5798,N_7540);
nand U12449 (N_12449,N_8429,N_5441);
xnor U12450 (N_12450,N_5411,N_7837);
or U12451 (N_12451,N_8228,N_6289);
nor U12452 (N_12452,N_5048,N_9110);
nor U12453 (N_12453,N_6986,N_6523);
xnor U12454 (N_12454,N_9953,N_5274);
or U12455 (N_12455,N_5359,N_9392);
and U12456 (N_12456,N_5365,N_7673);
or U12457 (N_12457,N_9375,N_5277);
and U12458 (N_12458,N_5144,N_5758);
and U12459 (N_12459,N_7575,N_6676);
or U12460 (N_12460,N_6781,N_8719);
nor U12461 (N_12461,N_6803,N_8453);
and U12462 (N_12462,N_8235,N_6630);
nand U12463 (N_12463,N_7772,N_8751);
nor U12464 (N_12464,N_9548,N_8628);
and U12465 (N_12465,N_7730,N_7548);
nor U12466 (N_12466,N_5018,N_5958);
or U12467 (N_12467,N_9022,N_6747);
and U12468 (N_12468,N_6634,N_7398);
xnor U12469 (N_12469,N_6866,N_8126);
nor U12470 (N_12470,N_8499,N_5212);
or U12471 (N_12471,N_5976,N_6403);
and U12472 (N_12472,N_5606,N_5777);
nand U12473 (N_12473,N_5911,N_5261);
nand U12474 (N_12474,N_5773,N_6991);
xnor U12475 (N_12475,N_5654,N_5640);
and U12476 (N_12476,N_6075,N_5865);
or U12477 (N_12477,N_7554,N_6135);
nor U12478 (N_12478,N_9425,N_7053);
nand U12479 (N_12479,N_6606,N_5336);
and U12480 (N_12480,N_6697,N_6021);
or U12481 (N_12481,N_6482,N_9837);
nor U12482 (N_12482,N_6373,N_9367);
xnor U12483 (N_12483,N_9104,N_7386);
or U12484 (N_12484,N_6420,N_5748);
nor U12485 (N_12485,N_5627,N_7157);
xnor U12486 (N_12486,N_7443,N_7288);
or U12487 (N_12487,N_8394,N_5913);
and U12488 (N_12488,N_7166,N_5060);
nor U12489 (N_12489,N_7703,N_8774);
nand U12490 (N_12490,N_9274,N_8855);
xor U12491 (N_12491,N_6987,N_7439);
and U12492 (N_12492,N_9566,N_6746);
or U12493 (N_12493,N_5515,N_8697);
xor U12494 (N_12494,N_6192,N_6613);
nand U12495 (N_12495,N_9630,N_9227);
and U12496 (N_12496,N_9625,N_5387);
and U12497 (N_12497,N_6216,N_8242);
or U12498 (N_12498,N_7529,N_9638);
or U12499 (N_12499,N_8035,N_7663);
xnor U12500 (N_12500,N_7359,N_7517);
xnor U12501 (N_12501,N_7327,N_7524);
xnor U12502 (N_12502,N_7824,N_5122);
nand U12503 (N_12503,N_9980,N_5168);
nor U12504 (N_12504,N_7716,N_9051);
xnor U12505 (N_12505,N_6881,N_5955);
xnor U12506 (N_12506,N_9519,N_5847);
nand U12507 (N_12507,N_7462,N_8862);
nor U12508 (N_12508,N_6102,N_8080);
nand U12509 (N_12509,N_9526,N_9879);
and U12510 (N_12510,N_5894,N_8785);
xor U12511 (N_12511,N_8656,N_9944);
nand U12512 (N_12512,N_7431,N_8590);
nor U12513 (N_12513,N_7015,N_5543);
xor U12514 (N_12514,N_8217,N_7876);
and U12515 (N_12515,N_5389,N_7101);
nand U12516 (N_12516,N_5589,N_9430);
and U12517 (N_12517,N_7966,N_5784);
or U12518 (N_12518,N_8668,N_8106);
or U12519 (N_12519,N_6896,N_7273);
nor U12520 (N_12520,N_9683,N_6973);
or U12521 (N_12521,N_5390,N_5286);
nor U12522 (N_12522,N_9278,N_8601);
xnor U12523 (N_12523,N_7680,N_8039);
or U12524 (N_12524,N_9942,N_8911);
and U12525 (N_12525,N_8368,N_6103);
nor U12526 (N_12526,N_6235,N_5443);
or U12527 (N_12527,N_7776,N_5415);
nor U12528 (N_12528,N_6741,N_5502);
nand U12529 (N_12529,N_5820,N_8377);
or U12530 (N_12530,N_7286,N_8769);
or U12531 (N_12531,N_6927,N_6011);
xnor U12532 (N_12532,N_5401,N_5654);
or U12533 (N_12533,N_5299,N_5119);
and U12534 (N_12534,N_9384,N_9612);
or U12535 (N_12535,N_6971,N_6170);
xor U12536 (N_12536,N_5612,N_7348);
or U12537 (N_12537,N_7218,N_6486);
nor U12538 (N_12538,N_5102,N_5007);
nor U12539 (N_12539,N_7752,N_5412);
xor U12540 (N_12540,N_5886,N_9961);
and U12541 (N_12541,N_9849,N_9194);
or U12542 (N_12542,N_7108,N_7523);
nor U12543 (N_12543,N_8360,N_8895);
or U12544 (N_12544,N_8005,N_9636);
nand U12545 (N_12545,N_8829,N_9807);
or U12546 (N_12546,N_7273,N_8132);
or U12547 (N_12547,N_8386,N_8878);
nor U12548 (N_12548,N_8296,N_7858);
and U12549 (N_12549,N_9688,N_6817);
nor U12550 (N_12550,N_9957,N_6419);
nor U12551 (N_12551,N_8229,N_6884);
nor U12552 (N_12552,N_8411,N_5164);
or U12553 (N_12553,N_7879,N_9532);
xnor U12554 (N_12554,N_6878,N_7993);
nand U12555 (N_12555,N_8755,N_6450);
or U12556 (N_12556,N_6276,N_5877);
nand U12557 (N_12557,N_9454,N_9535);
nand U12558 (N_12558,N_8538,N_6490);
nor U12559 (N_12559,N_9558,N_8630);
xor U12560 (N_12560,N_7317,N_9299);
xnor U12561 (N_12561,N_7588,N_7285);
xor U12562 (N_12562,N_8175,N_6320);
nor U12563 (N_12563,N_6305,N_6699);
nor U12564 (N_12564,N_8928,N_9018);
xor U12565 (N_12565,N_9644,N_5600);
nor U12566 (N_12566,N_6454,N_9241);
nand U12567 (N_12567,N_6993,N_7799);
and U12568 (N_12568,N_6079,N_6601);
nand U12569 (N_12569,N_8480,N_9814);
nor U12570 (N_12570,N_6529,N_5590);
or U12571 (N_12571,N_8507,N_7918);
or U12572 (N_12572,N_8629,N_6987);
or U12573 (N_12573,N_6493,N_9494);
and U12574 (N_12574,N_8332,N_8208);
nand U12575 (N_12575,N_6722,N_7774);
xor U12576 (N_12576,N_6235,N_5230);
or U12577 (N_12577,N_6596,N_8708);
nor U12578 (N_12578,N_9779,N_8106);
nand U12579 (N_12579,N_6513,N_7457);
nand U12580 (N_12580,N_5462,N_8688);
xor U12581 (N_12581,N_6910,N_5597);
and U12582 (N_12582,N_7008,N_9804);
nand U12583 (N_12583,N_7088,N_9506);
or U12584 (N_12584,N_5182,N_6284);
xnor U12585 (N_12585,N_8991,N_9940);
nand U12586 (N_12586,N_8146,N_6666);
or U12587 (N_12587,N_5241,N_5402);
nand U12588 (N_12588,N_8212,N_6432);
nor U12589 (N_12589,N_6025,N_7764);
xor U12590 (N_12590,N_5349,N_8568);
xor U12591 (N_12591,N_7914,N_6447);
or U12592 (N_12592,N_5370,N_9402);
xnor U12593 (N_12593,N_6998,N_5221);
nor U12594 (N_12594,N_9459,N_8040);
xnor U12595 (N_12595,N_6487,N_5873);
and U12596 (N_12596,N_8753,N_5248);
xnor U12597 (N_12597,N_7171,N_9856);
xor U12598 (N_12598,N_9822,N_5157);
or U12599 (N_12599,N_6123,N_9325);
nand U12600 (N_12600,N_9657,N_6149);
or U12601 (N_12601,N_9280,N_8973);
nand U12602 (N_12602,N_7597,N_8840);
xnor U12603 (N_12603,N_9576,N_5344);
and U12604 (N_12604,N_7693,N_5417);
and U12605 (N_12605,N_5918,N_8086);
xnor U12606 (N_12606,N_9514,N_8421);
nand U12607 (N_12607,N_6097,N_8355);
xnor U12608 (N_12608,N_9140,N_8002);
nor U12609 (N_12609,N_5618,N_7281);
nand U12610 (N_12610,N_7515,N_7735);
xor U12611 (N_12611,N_7309,N_8603);
or U12612 (N_12612,N_6985,N_8466);
or U12613 (N_12613,N_5939,N_7822);
nand U12614 (N_12614,N_5810,N_6081);
or U12615 (N_12615,N_7319,N_5554);
nand U12616 (N_12616,N_9210,N_9173);
nor U12617 (N_12617,N_7559,N_8303);
or U12618 (N_12618,N_9476,N_8448);
nand U12619 (N_12619,N_6383,N_8167);
nand U12620 (N_12620,N_8524,N_7868);
nand U12621 (N_12621,N_6482,N_6081);
xor U12622 (N_12622,N_5307,N_5006);
and U12623 (N_12623,N_5164,N_6093);
or U12624 (N_12624,N_6262,N_7507);
nand U12625 (N_12625,N_6746,N_5310);
and U12626 (N_12626,N_8057,N_5058);
nand U12627 (N_12627,N_7918,N_6386);
nand U12628 (N_12628,N_9750,N_7361);
xor U12629 (N_12629,N_8587,N_5654);
and U12630 (N_12630,N_7362,N_7390);
and U12631 (N_12631,N_9652,N_8781);
and U12632 (N_12632,N_6792,N_5299);
or U12633 (N_12633,N_9284,N_9403);
xor U12634 (N_12634,N_8769,N_5462);
nor U12635 (N_12635,N_8802,N_5682);
or U12636 (N_12636,N_5998,N_5241);
or U12637 (N_12637,N_5884,N_5900);
xor U12638 (N_12638,N_9559,N_7343);
and U12639 (N_12639,N_5344,N_6154);
xnor U12640 (N_12640,N_6507,N_8270);
xor U12641 (N_12641,N_9286,N_8274);
and U12642 (N_12642,N_8037,N_6803);
nor U12643 (N_12643,N_7165,N_9089);
or U12644 (N_12644,N_5823,N_5168);
nand U12645 (N_12645,N_9948,N_7416);
and U12646 (N_12646,N_7242,N_7955);
nand U12647 (N_12647,N_5614,N_7554);
or U12648 (N_12648,N_9472,N_7490);
and U12649 (N_12649,N_9246,N_9468);
nor U12650 (N_12650,N_9812,N_9401);
xor U12651 (N_12651,N_8272,N_7288);
xnor U12652 (N_12652,N_6067,N_9565);
xnor U12653 (N_12653,N_9604,N_5179);
or U12654 (N_12654,N_5779,N_9238);
xnor U12655 (N_12655,N_8514,N_8449);
xnor U12656 (N_12656,N_8508,N_5516);
and U12657 (N_12657,N_6153,N_6450);
nand U12658 (N_12658,N_5707,N_7108);
and U12659 (N_12659,N_8913,N_7975);
nand U12660 (N_12660,N_8544,N_8608);
nand U12661 (N_12661,N_9547,N_7751);
or U12662 (N_12662,N_5801,N_9494);
nand U12663 (N_12663,N_7006,N_8217);
xnor U12664 (N_12664,N_8916,N_6144);
or U12665 (N_12665,N_7883,N_5456);
and U12666 (N_12666,N_8693,N_9643);
nor U12667 (N_12667,N_7474,N_5832);
nand U12668 (N_12668,N_7089,N_8178);
nor U12669 (N_12669,N_9925,N_6464);
xnor U12670 (N_12670,N_5141,N_9821);
nand U12671 (N_12671,N_9757,N_6928);
or U12672 (N_12672,N_5755,N_7749);
nand U12673 (N_12673,N_5029,N_5313);
nor U12674 (N_12674,N_6751,N_5145);
nand U12675 (N_12675,N_7052,N_6165);
and U12676 (N_12676,N_8396,N_5543);
nor U12677 (N_12677,N_8329,N_9650);
or U12678 (N_12678,N_6961,N_6381);
nand U12679 (N_12679,N_7826,N_6806);
xor U12680 (N_12680,N_6972,N_5328);
xor U12681 (N_12681,N_7854,N_8479);
nand U12682 (N_12682,N_7057,N_5853);
xor U12683 (N_12683,N_7414,N_8567);
or U12684 (N_12684,N_7713,N_6692);
and U12685 (N_12685,N_7363,N_5457);
and U12686 (N_12686,N_5090,N_6916);
nor U12687 (N_12687,N_8559,N_9437);
or U12688 (N_12688,N_8705,N_7894);
xor U12689 (N_12689,N_7037,N_5840);
and U12690 (N_12690,N_6015,N_8414);
xor U12691 (N_12691,N_5622,N_8711);
or U12692 (N_12692,N_9619,N_7966);
nor U12693 (N_12693,N_5317,N_8097);
xor U12694 (N_12694,N_8463,N_5465);
nand U12695 (N_12695,N_9090,N_5728);
xnor U12696 (N_12696,N_5074,N_6981);
xor U12697 (N_12697,N_9684,N_5634);
xor U12698 (N_12698,N_6642,N_9666);
or U12699 (N_12699,N_8779,N_5304);
and U12700 (N_12700,N_6066,N_5716);
and U12701 (N_12701,N_8938,N_6579);
xor U12702 (N_12702,N_5812,N_6639);
nor U12703 (N_12703,N_5986,N_5621);
nand U12704 (N_12704,N_7581,N_9627);
and U12705 (N_12705,N_7035,N_9811);
or U12706 (N_12706,N_5548,N_7484);
nand U12707 (N_12707,N_9512,N_9779);
or U12708 (N_12708,N_5498,N_6826);
xnor U12709 (N_12709,N_9243,N_6924);
nor U12710 (N_12710,N_6609,N_7567);
nor U12711 (N_12711,N_9016,N_7278);
xor U12712 (N_12712,N_6735,N_5399);
and U12713 (N_12713,N_5548,N_9721);
or U12714 (N_12714,N_9821,N_6468);
nand U12715 (N_12715,N_5611,N_5144);
xor U12716 (N_12716,N_9769,N_9269);
xor U12717 (N_12717,N_8360,N_6466);
xnor U12718 (N_12718,N_9974,N_6000);
nand U12719 (N_12719,N_8542,N_7772);
and U12720 (N_12720,N_6604,N_8643);
or U12721 (N_12721,N_6938,N_5483);
or U12722 (N_12722,N_5512,N_7990);
nor U12723 (N_12723,N_6713,N_5672);
or U12724 (N_12724,N_7631,N_9248);
nand U12725 (N_12725,N_9589,N_5908);
and U12726 (N_12726,N_8682,N_7737);
and U12727 (N_12727,N_9774,N_5972);
nand U12728 (N_12728,N_8802,N_8811);
and U12729 (N_12729,N_7275,N_9542);
nor U12730 (N_12730,N_5240,N_5781);
or U12731 (N_12731,N_9005,N_8036);
and U12732 (N_12732,N_6942,N_6610);
nand U12733 (N_12733,N_8583,N_6130);
and U12734 (N_12734,N_5987,N_9750);
or U12735 (N_12735,N_9526,N_5399);
or U12736 (N_12736,N_8680,N_8195);
nor U12737 (N_12737,N_5163,N_9458);
or U12738 (N_12738,N_9289,N_8106);
and U12739 (N_12739,N_6660,N_6649);
xor U12740 (N_12740,N_9368,N_6136);
and U12741 (N_12741,N_6319,N_9931);
or U12742 (N_12742,N_9742,N_5760);
xnor U12743 (N_12743,N_7027,N_9197);
nor U12744 (N_12744,N_7673,N_8215);
and U12745 (N_12745,N_5741,N_5089);
nand U12746 (N_12746,N_7462,N_8628);
nand U12747 (N_12747,N_7339,N_6783);
nor U12748 (N_12748,N_9337,N_6158);
or U12749 (N_12749,N_7417,N_9867);
nand U12750 (N_12750,N_8829,N_8126);
xnor U12751 (N_12751,N_5819,N_8277);
nand U12752 (N_12752,N_7477,N_6076);
xor U12753 (N_12753,N_5547,N_5167);
nand U12754 (N_12754,N_7404,N_7298);
and U12755 (N_12755,N_7493,N_9470);
and U12756 (N_12756,N_6542,N_8501);
and U12757 (N_12757,N_6501,N_9266);
nand U12758 (N_12758,N_7935,N_9508);
or U12759 (N_12759,N_6617,N_8113);
and U12760 (N_12760,N_7349,N_8498);
nor U12761 (N_12761,N_7347,N_8061);
nor U12762 (N_12762,N_7020,N_6965);
nor U12763 (N_12763,N_9923,N_9214);
xor U12764 (N_12764,N_6701,N_6442);
xnor U12765 (N_12765,N_9740,N_5191);
xor U12766 (N_12766,N_5681,N_9529);
and U12767 (N_12767,N_5486,N_6304);
and U12768 (N_12768,N_7789,N_5098);
xor U12769 (N_12769,N_8266,N_8767);
or U12770 (N_12770,N_5029,N_6034);
nand U12771 (N_12771,N_9770,N_5586);
nand U12772 (N_12772,N_8305,N_8844);
nand U12773 (N_12773,N_9268,N_5570);
nor U12774 (N_12774,N_5287,N_7186);
nand U12775 (N_12775,N_9910,N_8054);
or U12776 (N_12776,N_5933,N_7552);
nor U12777 (N_12777,N_7992,N_9607);
and U12778 (N_12778,N_9317,N_7323);
or U12779 (N_12779,N_6436,N_6681);
nand U12780 (N_12780,N_8999,N_7669);
nand U12781 (N_12781,N_8200,N_5563);
or U12782 (N_12782,N_9153,N_6375);
xnor U12783 (N_12783,N_8170,N_7593);
and U12784 (N_12784,N_6045,N_5150);
and U12785 (N_12785,N_9014,N_6241);
or U12786 (N_12786,N_9187,N_9696);
nand U12787 (N_12787,N_9797,N_6799);
or U12788 (N_12788,N_6878,N_5617);
or U12789 (N_12789,N_6534,N_5237);
xnor U12790 (N_12790,N_9932,N_6300);
or U12791 (N_12791,N_5232,N_7497);
or U12792 (N_12792,N_8829,N_8460);
and U12793 (N_12793,N_7698,N_6277);
and U12794 (N_12794,N_8992,N_7186);
xor U12795 (N_12795,N_6216,N_5935);
xor U12796 (N_12796,N_6657,N_8831);
xor U12797 (N_12797,N_6277,N_6039);
nand U12798 (N_12798,N_5939,N_9076);
nand U12799 (N_12799,N_8748,N_8731);
and U12800 (N_12800,N_5478,N_6615);
and U12801 (N_12801,N_7251,N_5810);
xnor U12802 (N_12802,N_7508,N_6072);
nor U12803 (N_12803,N_5750,N_7701);
or U12804 (N_12804,N_5169,N_5332);
nand U12805 (N_12805,N_5990,N_5439);
or U12806 (N_12806,N_8442,N_9855);
or U12807 (N_12807,N_8030,N_5257);
xor U12808 (N_12808,N_6392,N_7412);
or U12809 (N_12809,N_8149,N_9906);
xnor U12810 (N_12810,N_6942,N_7636);
nor U12811 (N_12811,N_6437,N_6429);
or U12812 (N_12812,N_5300,N_5126);
nand U12813 (N_12813,N_6862,N_8059);
nor U12814 (N_12814,N_6864,N_9307);
and U12815 (N_12815,N_8190,N_6835);
nor U12816 (N_12816,N_8724,N_7426);
nor U12817 (N_12817,N_5846,N_5062);
xnor U12818 (N_12818,N_7494,N_9159);
or U12819 (N_12819,N_5392,N_6123);
or U12820 (N_12820,N_9567,N_8448);
or U12821 (N_12821,N_5672,N_6978);
and U12822 (N_12822,N_6125,N_7792);
nor U12823 (N_12823,N_6923,N_8468);
and U12824 (N_12824,N_7563,N_8090);
and U12825 (N_12825,N_5539,N_5889);
xor U12826 (N_12826,N_5414,N_8759);
nor U12827 (N_12827,N_7016,N_8518);
nand U12828 (N_12828,N_5428,N_7924);
and U12829 (N_12829,N_5778,N_9732);
xnor U12830 (N_12830,N_7241,N_8608);
nor U12831 (N_12831,N_6744,N_7646);
or U12832 (N_12832,N_6552,N_7428);
nor U12833 (N_12833,N_5137,N_6496);
and U12834 (N_12834,N_5810,N_5076);
and U12835 (N_12835,N_7144,N_6428);
nor U12836 (N_12836,N_8481,N_6105);
and U12837 (N_12837,N_9616,N_6507);
nand U12838 (N_12838,N_9060,N_6412);
nand U12839 (N_12839,N_7023,N_6328);
xnor U12840 (N_12840,N_8898,N_8447);
nor U12841 (N_12841,N_5571,N_8026);
xnor U12842 (N_12842,N_7902,N_8591);
and U12843 (N_12843,N_5776,N_6149);
nor U12844 (N_12844,N_7809,N_7643);
nor U12845 (N_12845,N_6902,N_9730);
nand U12846 (N_12846,N_8564,N_6394);
or U12847 (N_12847,N_9761,N_8969);
nor U12848 (N_12848,N_9710,N_7528);
nand U12849 (N_12849,N_5153,N_8600);
nand U12850 (N_12850,N_5574,N_6377);
and U12851 (N_12851,N_8257,N_7150);
xor U12852 (N_12852,N_6565,N_8593);
xor U12853 (N_12853,N_5748,N_5290);
nor U12854 (N_12854,N_5883,N_9287);
nor U12855 (N_12855,N_7906,N_7268);
and U12856 (N_12856,N_8850,N_5271);
xnor U12857 (N_12857,N_8093,N_8516);
xor U12858 (N_12858,N_5462,N_7973);
nand U12859 (N_12859,N_5314,N_8731);
nor U12860 (N_12860,N_5190,N_5112);
nor U12861 (N_12861,N_5991,N_6094);
and U12862 (N_12862,N_6418,N_5219);
xnor U12863 (N_12863,N_7717,N_7170);
nand U12864 (N_12864,N_6189,N_6069);
xor U12865 (N_12865,N_5229,N_7946);
or U12866 (N_12866,N_6338,N_9316);
nor U12867 (N_12867,N_8391,N_8078);
nand U12868 (N_12868,N_9856,N_5175);
or U12869 (N_12869,N_6123,N_5426);
and U12870 (N_12870,N_5686,N_9561);
or U12871 (N_12871,N_6825,N_7744);
or U12872 (N_12872,N_6216,N_9761);
xnor U12873 (N_12873,N_9510,N_9543);
nor U12874 (N_12874,N_6435,N_6088);
nand U12875 (N_12875,N_5936,N_6032);
xnor U12876 (N_12876,N_5785,N_5707);
nor U12877 (N_12877,N_5790,N_7238);
and U12878 (N_12878,N_5280,N_7740);
nor U12879 (N_12879,N_8591,N_9924);
nand U12880 (N_12880,N_9402,N_8908);
and U12881 (N_12881,N_7089,N_5558);
nor U12882 (N_12882,N_5605,N_6079);
and U12883 (N_12883,N_7347,N_5987);
or U12884 (N_12884,N_7072,N_8672);
and U12885 (N_12885,N_7622,N_8045);
xnor U12886 (N_12886,N_6798,N_9064);
or U12887 (N_12887,N_5987,N_5358);
or U12888 (N_12888,N_9616,N_7939);
nand U12889 (N_12889,N_9573,N_5737);
and U12890 (N_12890,N_6282,N_5304);
nand U12891 (N_12891,N_8557,N_9653);
and U12892 (N_12892,N_5554,N_5655);
or U12893 (N_12893,N_6528,N_9834);
xnor U12894 (N_12894,N_8100,N_7346);
xnor U12895 (N_12895,N_9243,N_5509);
nor U12896 (N_12896,N_7987,N_7598);
xor U12897 (N_12897,N_7112,N_6288);
xnor U12898 (N_12898,N_7448,N_7166);
or U12899 (N_12899,N_6152,N_7335);
xor U12900 (N_12900,N_5668,N_8981);
nor U12901 (N_12901,N_9580,N_7411);
nand U12902 (N_12902,N_5446,N_8297);
xnor U12903 (N_12903,N_9177,N_5060);
nand U12904 (N_12904,N_6166,N_7389);
and U12905 (N_12905,N_9465,N_8830);
and U12906 (N_12906,N_8070,N_9846);
nand U12907 (N_12907,N_5113,N_5977);
or U12908 (N_12908,N_6198,N_7605);
or U12909 (N_12909,N_9070,N_7900);
nor U12910 (N_12910,N_7327,N_8441);
nor U12911 (N_12911,N_6251,N_6392);
xnor U12912 (N_12912,N_6282,N_7681);
and U12913 (N_12913,N_8819,N_8492);
nand U12914 (N_12914,N_5274,N_8263);
nor U12915 (N_12915,N_8770,N_6555);
or U12916 (N_12916,N_8041,N_6501);
nor U12917 (N_12917,N_7555,N_9806);
nand U12918 (N_12918,N_8575,N_9611);
xor U12919 (N_12919,N_7056,N_8640);
xnor U12920 (N_12920,N_8477,N_7495);
xnor U12921 (N_12921,N_6874,N_5612);
nor U12922 (N_12922,N_7018,N_9843);
or U12923 (N_12923,N_9997,N_9538);
xnor U12924 (N_12924,N_6065,N_9011);
xnor U12925 (N_12925,N_8189,N_5477);
nor U12926 (N_12926,N_5158,N_8306);
xor U12927 (N_12927,N_7508,N_5519);
nand U12928 (N_12928,N_7780,N_6684);
nor U12929 (N_12929,N_8736,N_9649);
and U12930 (N_12930,N_8337,N_8538);
and U12931 (N_12931,N_8697,N_7810);
nand U12932 (N_12932,N_5816,N_6349);
and U12933 (N_12933,N_8530,N_7160);
nor U12934 (N_12934,N_5791,N_8656);
nand U12935 (N_12935,N_6965,N_7403);
or U12936 (N_12936,N_5403,N_5882);
and U12937 (N_12937,N_9769,N_9187);
and U12938 (N_12938,N_6109,N_9773);
or U12939 (N_12939,N_6155,N_6793);
nor U12940 (N_12940,N_7691,N_7644);
or U12941 (N_12941,N_8633,N_6778);
and U12942 (N_12942,N_8707,N_5255);
nand U12943 (N_12943,N_5414,N_9684);
nor U12944 (N_12944,N_5093,N_6944);
nor U12945 (N_12945,N_5182,N_9720);
nand U12946 (N_12946,N_5819,N_6057);
nand U12947 (N_12947,N_7446,N_7161);
nor U12948 (N_12948,N_8991,N_9031);
and U12949 (N_12949,N_6801,N_5116);
and U12950 (N_12950,N_5586,N_8367);
xnor U12951 (N_12951,N_7164,N_6169);
and U12952 (N_12952,N_9607,N_8855);
or U12953 (N_12953,N_9789,N_9573);
or U12954 (N_12954,N_9754,N_9822);
and U12955 (N_12955,N_6048,N_8588);
nand U12956 (N_12956,N_8820,N_8270);
nand U12957 (N_12957,N_5542,N_9484);
or U12958 (N_12958,N_9086,N_5497);
nand U12959 (N_12959,N_6622,N_9181);
xnor U12960 (N_12960,N_6826,N_6272);
and U12961 (N_12961,N_8238,N_8839);
or U12962 (N_12962,N_8882,N_8569);
nor U12963 (N_12963,N_6605,N_7362);
xor U12964 (N_12964,N_5894,N_6682);
xor U12965 (N_12965,N_5040,N_6748);
xnor U12966 (N_12966,N_7279,N_5609);
nand U12967 (N_12967,N_5813,N_8819);
nand U12968 (N_12968,N_8633,N_9396);
and U12969 (N_12969,N_7310,N_9270);
xor U12970 (N_12970,N_5240,N_5057);
or U12971 (N_12971,N_5059,N_5004);
and U12972 (N_12972,N_8643,N_6076);
nor U12973 (N_12973,N_6039,N_5214);
nand U12974 (N_12974,N_5318,N_6216);
nand U12975 (N_12975,N_7470,N_9530);
and U12976 (N_12976,N_5445,N_9467);
and U12977 (N_12977,N_6090,N_6840);
xor U12978 (N_12978,N_8684,N_8686);
xor U12979 (N_12979,N_9589,N_9282);
or U12980 (N_12980,N_9505,N_5350);
xnor U12981 (N_12981,N_6402,N_7577);
or U12982 (N_12982,N_9597,N_5010);
nand U12983 (N_12983,N_7912,N_7325);
nand U12984 (N_12984,N_7922,N_8644);
nand U12985 (N_12985,N_6335,N_8721);
xor U12986 (N_12986,N_5486,N_6506);
nor U12987 (N_12987,N_8352,N_8141);
nor U12988 (N_12988,N_5555,N_9951);
nand U12989 (N_12989,N_9822,N_7860);
xor U12990 (N_12990,N_8226,N_7089);
nand U12991 (N_12991,N_5279,N_7342);
and U12992 (N_12992,N_7937,N_9797);
or U12993 (N_12993,N_8934,N_7747);
nand U12994 (N_12994,N_7991,N_9286);
xnor U12995 (N_12995,N_6979,N_9596);
xnor U12996 (N_12996,N_6621,N_6121);
nand U12997 (N_12997,N_5235,N_8649);
nor U12998 (N_12998,N_7224,N_9963);
nor U12999 (N_12999,N_8651,N_7158);
nor U13000 (N_13000,N_6927,N_8100);
or U13001 (N_13001,N_7568,N_9941);
and U13002 (N_13002,N_6725,N_8701);
nor U13003 (N_13003,N_7425,N_7063);
nor U13004 (N_13004,N_9913,N_9569);
or U13005 (N_13005,N_7041,N_9310);
nor U13006 (N_13006,N_5686,N_9081);
and U13007 (N_13007,N_5306,N_6842);
xor U13008 (N_13008,N_8806,N_5076);
or U13009 (N_13009,N_8645,N_6402);
nor U13010 (N_13010,N_7363,N_9990);
and U13011 (N_13011,N_6169,N_9100);
nor U13012 (N_13012,N_8913,N_5445);
xnor U13013 (N_13013,N_9384,N_6786);
nor U13014 (N_13014,N_7918,N_6205);
xor U13015 (N_13015,N_6619,N_9780);
xor U13016 (N_13016,N_5220,N_6318);
nand U13017 (N_13017,N_6434,N_6176);
nor U13018 (N_13018,N_6996,N_8985);
and U13019 (N_13019,N_5987,N_5957);
nand U13020 (N_13020,N_5118,N_7447);
nor U13021 (N_13021,N_6152,N_5722);
and U13022 (N_13022,N_9441,N_5795);
xnor U13023 (N_13023,N_6071,N_6483);
nand U13024 (N_13024,N_8798,N_7158);
nand U13025 (N_13025,N_5670,N_7630);
xnor U13026 (N_13026,N_7474,N_5421);
or U13027 (N_13027,N_7935,N_6727);
nand U13028 (N_13028,N_7712,N_7346);
nor U13029 (N_13029,N_7878,N_8052);
xnor U13030 (N_13030,N_8634,N_5917);
and U13031 (N_13031,N_7986,N_6237);
and U13032 (N_13032,N_9396,N_7800);
nand U13033 (N_13033,N_7151,N_6670);
xor U13034 (N_13034,N_8549,N_5774);
or U13035 (N_13035,N_6600,N_5830);
nand U13036 (N_13036,N_7771,N_7229);
nand U13037 (N_13037,N_6501,N_7383);
nor U13038 (N_13038,N_9066,N_6729);
nand U13039 (N_13039,N_6182,N_7341);
and U13040 (N_13040,N_8583,N_9468);
nor U13041 (N_13041,N_8921,N_6961);
xnor U13042 (N_13042,N_9179,N_6996);
xor U13043 (N_13043,N_9000,N_6335);
nor U13044 (N_13044,N_6745,N_5710);
xor U13045 (N_13045,N_9175,N_6764);
and U13046 (N_13046,N_5367,N_9711);
xnor U13047 (N_13047,N_7089,N_5140);
nor U13048 (N_13048,N_5440,N_8907);
and U13049 (N_13049,N_9749,N_7812);
or U13050 (N_13050,N_5997,N_5138);
nor U13051 (N_13051,N_5841,N_9519);
xor U13052 (N_13052,N_6974,N_5266);
or U13053 (N_13053,N_6739,N_6771);
nor U13054 (N_13054,N_6831,N_5726);
nand U13055 (N_13055,N_6903,N_7142);
nor U13056 (N_13056,N_9976,N_9712);
or U13057 (N_13057,N_9077,N_6232);
xnor U13058 (N_13058,N_9247,N_8982);
nor U13059 (N_13059,N_8560,N_6350);
and U13060 (N_13060,N_9547,N_5900);
and U13061 (N_13061,N_7062,N_9697);
or U13062 (N_13062,N_9870,N_6657);
or U13063 (N_13063,N_7220,N_7431);
xnor U13064 (N_13064,N_7920,N_6670);
and U13065 (N_13065,N_8384,N_8221);
or U13066 (N_13066,N_7887,N_5442);
xor U13067 (N_13067,N_5546,N_7425);
and U13068 (N_13068,N_9696,N_6816);
nor U13069 (N_13069,N_9823,N_6020);
or U13070 (N_13070,N_5003,N_6159);
and U13071 (N_13071,N_8340,N_9052);
nand U13072 (N_13072,N_5775,N_7809);
nor U13073 (N_13073,N_7284,N_9380);
nor U13074 (N_13074,N_5606,N_6139);
and U13075 (N_13075,N_9226,N_7883);
and U13076 (N_13076,N_7512,N_7685);
or U13077 (N_13077,N_7202,N_6694);
or U13078 (N_13078,N_7871,N_5151);
nand U13079 (N_13079,N_6409,N_7297);
nor U13080 (N_13080,N_6527,N_9245);
and U13081 (N_13081,N_7033,N_7946);
nand U13082 (N_13082,N_8843,N_5818);
nand U13083 (N_13083,N_8146,N_7369);
nor U13084 (N_13084,N_5318,N_6549);
xor U13085 (N_13085,N_8271,N_5346);
xnor U13086 (N_13086,N_8129,N_6459);
and U13087 (N_13087,N_7667,N_9064);
or U13088 (N_13088,N_6092,N_7278);
or U13089 (N_13089,N_7510,N_7463);
or U13090 (N_13090,N_9965,N_7769);
nor U13091 (N_13091,N_6231,N_7613);
or U13092 (N_13092,N_9400,N_6986);
nand U13093 (N_13093,N_5080,N_8390);
nor U13094 (N_13094,N_5126,N_7161);
and U13095 (N_13095,N_5370,N_5105);
or U13096 (N_13096,N_8259,N_6737);
nor U13097 (N_13097,N_5924,N_8379);
xor U13098 (N_13098,N_5961,N_8223);
nand U13099 (N_13099,N_5065,N_7733);
nand U13100 (N_13100,N_6441,N_8685);
xnor U13101 (N_13101,N_9711,N_9740);
or U13102 (N_13102,N_9251,N_7462);
and U13103 (N_13103,N_6208,N_8820);
xnor U13104 (N_13104,N_6211,N_8384);
or U13105 (N_13105,N_9360,N_5869);
xnor U13106 (N_13106,N_7393,N_7747);
nor U13107 (N_13107,N_9974,N_9033);
nand U13108 (N_13108,N_6067,N_7144);
nor U13109 (N_13109,N_5050,N_8657);
xor U13110 (N_13110,N_9430,N_6796);
xnor U13111 (N_13111,N_7589,N_9819);
nand U13112 (N_13112,N_7048,N_5835);
xnor U13113 (N_13113,N_8316,N_7518);
xor U13114 (N_13114,N_8538,N_5129);
xnor U13115 (N_13115,N_6777,N_7174);
xor U13116 (N_13116,N_8336,N_5966);
nor U13117 (N_13117,N_6506,N_6551);
or U13118 (N_13118,N_7107,N_8261);
nor U13119 (N_13119,N_7663,N_7310);
nor U13120 (N_13120,N_9163,N_8162);
and U13121 (N_13121,N_8645,N_5693);
xnor U13122 (N_13122,N_8217,N_9626);
xnor U13123 (N_13123,N_6983,N_5865);
nor U13124 (N_13124,N_7368,N_8581);
or U13125 (N_13125,N_8711,N_8427);
and U13126 (N_13126,N_5823,N_8674);
xor U13127 (N_13127,N_8264,N_5501);
xnor U13128 (N_13128,N_9760,N_5084);
nand U13129 (N_13129,N_5927,N_6408);
nand U13130 (N_13130,N_5287,N_5496);
or U13131 (N_13131,N_8546,N_8569);
nor U13132 (N_13132,N_8387,N_7057);
nor U13133 (N_13133,N_6701,N_7169);
nand U13134 (N_13134,N_8362,N_9746);
and U13135 (N_13135,N_8430,N_7534);
xor U13136 (N_13136,N_8133,N_6726);
nand U13137 (N_13137,N_6691,N_8503);
xnor U13138 (N_13138,N_5956,N_7009);
nand U13139 (N_13139,N_7617,N_8719);
or U13140 (N_13140,N_9940,N_5414);
nand U13141 (N_13141,N_7640,N_9416);
xnor U13142 (N_13142,N_8496,N_6005);
and U13143 (N_13143,N_5685,N_7812);
or U13144 (N_13144,N_6836,N_7023);
nor U13145 (N_13145,N_6044,N_5444);
and U13146 (N_13146,N_7840,N_6282);
nand U13147 (N_13147,N_7547,N_9693);
nor U13148 (N_13148,N_7865,N_8164);
nand U13149 (N_13149,N_6165,N_8559);
or U13150 (N_13150,N_9972,N_7632);
nor U13151 (N_13151,N_9021,N_5268);
xor U13152 (N_13152,N_5004,N_9115);
or U13153 (N_13153,N_7169,N_6751);
xnor U13154 (N_13154,N_6512,N_9090);
or U13155 (N_13155,N_7824,N_7957);
and U13156 (N_13156,N_7340,N_7427);
and U13157 (N_13157,N_7241,N_7824);
xor U13158 (N_13158,N_8706,N_5654);
or U13159 (N_13159,N_6545,N_6354);
and U13160 (N_13160,N_7783,N_5330);
xnor U13161 (N_13161,N_6622,N_7661);
xnor U13162 (N_13162,N_6984,N_5409);
or U13163 (N_13163,N_5091,N_8396);
and U13164 (N_13164,N_6678,N_8691);
nor U13165 (N_13165,N_8762,N_6887);
nand U13166 (N_13166,N_6964,N_7698);
nand U13167 (N_13167,N_6845,N_5842);
nand U13168 (N_13168,N_7615,N_5133);
nand U13169 (N_13169,N_5399,N_6512);
or U13170 (N_13170,N_6643,N_9667);
nand U13171 (N_13171,N_6915,N_7804);
xor U13172 (N_13172,N_5478,N_8815);
xnor U13173 (N_13173,N_6085,N_7146);
nor U13174 (N_13174,N_9034,N_8686);
or U13175 (N_13175,N_6002,N_7892);
nand U13176 (N_13176,N_6202,N_7561);
nand U13177 (N_13177,N_7517,N_6566);
and U13178 (N_13178,N_5855,N_8351);
xnor U13179 (N_13179,N_9082,N_9695);
nand U13180 (N_13180,N_6380,N_9851);
xor U13181 (N_13181,N_7253,N_8922);
nor U13182 (N_13182,N_5523,N_7675);
nand U13183 (N_13183,N_6612,N_5819);
or U13184 (N_13184,N_5548,N_7071);
xor U13185 (N_13185,N_7107,N_9861);
and U13186 (N_13186,N_8044,N_5986);
nand U13187 (N_13187,N_7783,N_6390);
and U13188 (N_13188,N_7735,N_8027);
and U13189 (N_13189,N_8515,N_7130);
nand U13190 (N_13190,N_6148,N_6119);
or U13191 (N_13191,N_8933,N_9408);
and U13192 (N_13192,N_7701,N_6070);
nand U13193 (N_13193,N_6937,N_8540);
xnor U13194 (N_13194,N_7607,N_6519);
and U13195 (N_13195,N_9792,N_8825);
xor U13196 (N_13196,N_9933,N_9481);
or U13197 (N_13197,N_7863,N_9609);
or U13198 (N_13198,N_9577,N_7536);
nand U13199 (N_13199,N_9876,N_8904);
and U13200 (N_13200,N_8440,N_8173);
nand U13201 (N_13201,N_6936,N_7114);
nand U13202 (N_13202,N_9591,N_7119);
and U13203 (N_13203,N_8322,N_6260);
nor U13204 (N_13204,N_8680,N_8048);
nor U13205 (N_13205,N_7462,N_8885);
nor U13206 (N_13206,N_6202,N_6145);
xnor U13207 (N_13207,N_9429,N_5390);
nor U13208 (N_13208,N_8898,N_7883);
nand U13209 (N_13209,N_5900,N_7855);
xor U13210 (N_13210,N_8778,N_6400);
xor U13211 (N_13211,N_7622,N_8143);
nor U13212 (N_13212,N_6663,N_6992);
nor U13213 (N_13213,N_9539,N_8854);
and U13214 (N_13214,N_5369,N_9331);
or U13215 (N_13215,N_6961,N_6452);
or U13216 (N_13216,N_6475,N_8430);
and U13217 (N_13217,N_9636,N_6398);
xnor U13218 (N_13218,N_6803,N_9305);
nor U13219 (N_13219,N_7267,N_9751);
xnor U13220 (N_13220,N_9418,N_8257);
nor U13221 (N_13221,N_8296,N_8491);
or U13222 (N_13222,N_8619,N_5458);
nand U13223 (N_13223,N_7018,N_7318);
nor U13224 (N_13224,N_8826,N_9270);
and U13225 (N_13225,N_8185,N_8298);
nor U13226 (N_13226,N_9509,N_9345);
nand U13227 (N_13227,N_9893,N_5511);
and U13228 (N_13228,N_8687,N_8205);
and U13229 (N_13229,N_8714,N_7438);
or U13230 (N_13230,N_6967,N_6949);
xnor U13231 (N_13231,N_8841,N_5216);
and U13232 (N_13232,N_7499,N_9637);
or U13233 (N_13233,N_9375,N_6154);
or U13234 (N_13234,N_7301,N_5221);
and U13235 (N_13235,N_7084,N_9556);
or U13236 (N_13236,N_7104,N_9411);
nand U13237 (N_13237,N_8477,N_7946);
and U13238 (N_13238,N_8287,N_6387);
or U13239 (N_13239,N_8917,N_6063);
xor U13240 (N_13240,N_5007,N_5882);
nand U13241 (N_13241,N_9812,N_7045);
or U13242 (N_13242,N_8624,N_5305);
nor U13243 (N_13243,N_8940,N_9541);
nor U13244 (N_13244,N_7712,N_6020);
xnor U13245 (N_13245,N_5547,N_7281);
nor U13246 (N_13246,N_6058,N_7748);
and U13247 (N_13247,N_5488,N_6091);
nor U13248 (N_13248,N_5508,N_5382);
nor U13249 (N_13249,N_8777,N_7826);
and U13250 (N_13250,N_6497,N_6352);
nand U13251 (N_13251,N_5148,N_6414);
or U13252 (N_13252,N_6063,N_5559);
and U13253 (N_13253,N_8372,N_7615);
nor U13254 (N_13254,N_7199,N_9595);
nor U13255 (N_13255,N_6513,N_8144);
nor U13256 (N_13256,N_5919,N_9327);
and U13257 (N_13257,N_5060,N_5762);
nand U13258 (N_13258,N_7457,N_9690);
or U13259 (N_13259,N_7860,N_5850);
and U13260 (N_13260,N_6569,N_8688);
nor U13261 (N_13261,N_8862,N_8448);
nand U13262 (N_13262,N_6514,N_6404);
nor U13263 (N_13263,N_9463,N_6409);
nand U13264 (N_13264,N_9320,N_9542);
nor U13265 (N_13265,N_5931,N_7562);
nor U13266 (N_13266,N_7899,N_9295);
nor U13267 (N_13267,N_8954,N_6379);
nand U13268 (N_13268,N_9966,N_8648);
nand U13269 (N_13269,N_8898,N_6447);
nand U13270 (N_13270,N_9329,N_8718);
nor U13271 (N_13271,N_7904,N_6423);
xnor U13272 (N_13272,N_9854,N_6726);
and U13273 (N_13273,N_7638,N_9373);
and U13274 (N_13274,N_8801,N_7255);
nor U13275 (N_13275,N_5948,N_5497);
xor U13276 (N_13276,N_5341,N_5615);
or U13277 (N_13277,N_7821,N_5436);
nand U13278 (N_13278,N_9455,N_5103);
nor U13279 (N_13279,N_5450,N_9153);
nor U13280 (N_13280,N_6808,N_6583);
and U13281 (N_13281,N_9728,N_6114);
and U13282 (N_13282,N_9243,N_7061);
and U13283 (N_13283,N_6253,N_7550);
xnor U13284 (N_13284,N_6090,N_7604);
nand U13285 (N_13285,N_6134,N_6969);
xnor U13286 (N_13286,N_6661,N_5528);
nand U13287 (N_13287,N_7312,N_6282);
nor U13288 (N_13288,N_8401,N_9417);
xnor U13289 (N_13289,N_5377,N_5030);
nand U13290 (N_13290,N_8222,N_5166);
nand U13291 (N_13291,N_5842,N_5468);
xnor U13292 (N_13292,N_5270,N_6434);
and U13293 (N_13293,N_7157,N_7114);
nand U13294 (N_13294,N_8435,N_6912);
nor U13295 (N_13295,N_9333,N_6721);
and U13296 (N_13296,N_8272,N_6715);
nor U13297 (N_13297,N_7742,N_5984);
and U13298 (N_13298,N_6447,N_6118);
xnor U13299 (N_13299,N_8331,N_5251);
and U13300 (N_13300,N_9969,N_6294);
xor U13301 (N_13301,N_7007,N_6454);
and U13302 (N_13302,N_9219,N_5109);
nand U13303 (N_13303,N_7965,N_5645);
xor U13304 (N_13304,N_7355,N_9244);
nand U13305 (N_13305,N_5801,N_8610);
nand U13306 (N_13306,N_7443,N_6089);
and U13307 (N_13307,N_8409,N_8660);
nand U13308 (N_13308,N_7436,N_9985);
and U13309 (N_13309,N_5665,N_6866);
and U13310 (N_13310,N_7079,N_5696);
xnor U13311 (N_13311,N_5078,N_5601);
xor U13312 (N_13312,N_6733,N_5547);
xor U13313 (N_13313,N_6572,N_5905);
or U13314 (N_13314,N_7696,N_9120);
xor U13315 (N_13315,N_5683,N_9860);
xor U13316 (N_13316,N_5782,N_7867);
or U13317 (N_13317,N_5265,N_5567);
xor U13318 (N_13318,N_6902,N_7230);
nor U13319 (N_13319,N_5904,N_8217);
and U13320 (N_13320,N_8763,N_6138);
nand U13321 (N_13321,N_7833,N_8693);
xnor U13322 (N_13322,N_5598,N_8158);
xnor U13323 (N_13323,N_8743,N_8939);
or U13324 (N_13324,N_7646,N_8963);
nand U13325 (N_13325,N_9432,N_7314);
nand U13326 (N_13326,N_8492,N_7250);
xnor U13327 (N_13327,N_7315,N_5178);
xnor U13328 (N_13328,N_6251,N_9309);
nor U13329 (N_13329,N_9546,N_5071);
nor U13330 (N_13330,N_7095,N_9058);
and U13331 (N_13331,N_7883,N_5892);
nand U13332 (N_13332,N_8925,N_8058);
and U13333 (N_13333,N_5627,N_6306);
and U13334 (N_13334,N_6858,N_7015);
and U13335 (N_13335,N_9733,N_8985);
and U13336 (N_13336,N_7232,N_5163);
xor U13337 (N_13337,N_5886,N_6235);
and U13338 (N_13338,N_5169,N_7100);
xnor U13339 (N_13339,N_9344,N_6401);
or U13340 (N_13340,N_6819,N_5084);
and U13341 (N_13341,N_6267,N_5327);
nand U13342 (N_13342,N_9776,N_6451);
nor U13343 (N_13343,N_9440,N_7392);
or U13344 (N_13344,N_8752,N_7684);
nand U13345 (N_13345,N_5873,N_8389);
nand U13346 (N_13346,N_8334,N_8053);
nand U13347 (N_13347,N_9574,N_7013);
xnor U13348 (N_13348,N_8468,N_6709);
nand U13349 (N_13349,N_8174,N_8726);
and U13350 (N_13350,N_5020,N_6468);
nand U13351 (N_13351,N_6677,N_8995);
or U13352 (N_13352,N_8145,N_9365);
or U13353 (N_13353,N_8271,N_6551);
and U13354 (N_13354,N_6495,N_7610);
and U13355 (N_13355,N_7049,N_6692);
nor U13356 (N_13356,N_7415,N_6171);
nand U13357 (N_13357,N_9986,N_6159);
nand U13358 (N_13358,N_7550,N_9569);
or U13359 (N_13359,N_8296,N_5782);
or U13360 (N_13360,N_7423,N_8623);
and U13361 (N_13361,N_6293,N_9802);
nor U13362 (N_13362,N_6076,N_5667);
and U13363 (N_13363,N_5374,N_6132);
nand U13364 (N_13364,N_9795,N_7361);
xor U13365 (N_13365,N_8529,N_5822);
xnor U13366 (N_13366,N_7837,N_8143);
and U13367 (N_13367,N_5620,N_6697);
nor U13368 (N_13368,N_7285,N_6576);
and U13369 (N_13369,N_5311,N_5957);
nand U13370 (N_13370,N_6703,N_6381);
or U13371 (N_13371,N_9340,N_7783);
and U13372 (N_13372,N_6504,N_6725);
nor U13373 (N_13373,N_6641,N_6898);
or U13374 (N_13374,N_9719,N_7469);
xor U13375 (N_13375,N_5160,N_7041);
xnor U13376 (N_13376,N_5940,N_5728);
or U13377 (N_13377,N_7128,N_5966);
and U13378 (N_13378,N_8457,N_7722);
or U13379 (N_13379,N_9003,N_7776);
nand U13380 (N_13380,N_6862,N_8699);
xnor U13381 (N_13381,N_6670,N_8180);
or U13382 (N_13382,N_6932,N_9979);
nand U13383 (N_13383,N_5178,N_5622);
and U13384 (N_13384,N_5848,N_6914);
xor U13385 (N_13385,N_7091,N_9014);
or U13386 (N_13386,N_9594,N_7958);
or U13387 (N_13387,N_9442,N_6891);
or U13388 (N_13388,N_6162,N_7933);
and U13389 (N_13389,N_9557,N_7558);
nand U13390 (N_13390,N_5211,N_8768);
and U13391 (N_13391,N_9867,N_9440);
nand U13392 (N_13392,N_7164,N_7427);
nor U13393 (N_13393,N_6306,N_8644);
and U13394 (N_13394,N_8071,N_8405);
nand U13395 (N_13395,N_5616,N_5845);
and U13396 (N_13396,N_7624,N_5926);
and U13397 (N_13397,N_6383,N_7037);
nand U13398 (N_13398,N_6108,N_7325);
and U13399 (N_13399,N_9508,N_8131);
nor U13400 (N_13400,N_9848,N_9044);
nor U13401 (N_13401,N_6056,N_8075);
or U13402 (N_13402,N_5132,N_9727);
or U13403 (N_13403,N_7769,N_8946);
xor U13404 (N_13404,N_7603,N_6507);
and U13405 (N_13405,N_8523,N_7396);
nor U13406 (N_13406,N_5552,N_5897);
nand U13407 (N_13407,N_7099,N_7345);
nor U13408 (N_13408,N_6515,N_9650);
xor U13409 (N_13409,N_8654,N_5743);
or U13410 (N_13410,N_5800,N_5271);
or U13411 (N_13411,N_6045,N_7130);
or U13412 (N_13412,N_8057,N_5935);
and U13413 (N_13413,N_6732,N_9585);
or U13414 (N_13414,N_9891,N_5075);
nand U13415 (N_13415,N_8858,N_6237);
xnor U13416 (N_13416,N_9874,N_9954);
xnor U13417 (N_13417,N_7564,N_7061);
and U13418 (N_13418,N_8926,N_8698);
xor U13419 (N_13419,N_6215,N_5417);
xor U13420 (N_13420,N_6165,N_6361);
nor U13421 (N_13421,N_6447,N_6512);
nand U13422 (N_13422,N_7974,N_9404);
nand U13423 (N_13423,N_6387,N_8074);
and U13424 (N_13424,N_6855,N_8524);
xor U13425 (N_13425,N_9902,N_7034);
xor U13426 (N_13426,N_7034,N_7508);
and U13427 (N_13427,N_5568,N_7536);
and U13428 (N_13428,N_7775,N_7686);
xor U13429 (N_13429,N_7764,N_8906);
and U13430 (N_13430,N_5795,N_7237);
xnor U13431 (N_13431,N_7406,N_6682);
xor U13432 (N_13432,N_5870,N_9487);
or U13433 (N_13433,N_7289,N_9943);
nand U13434 (N_13434,N_5022,N_5398);
or U13435 (N_13435,N_8973,N_9082);
and U13436 (N_13436,N_9860,N_6415);
nor U13437 (N_13437,N_8342,N_6062);
and U13438 (N_13438,N_5937,N_6308);
and U13439 (N_13439,N_6937,N_8705);
or U13440 (N_13440,N_6135,N_6211);
xor U13441 (N_13441,N_9017,N_9548);
and U13442 (N_13442,N_5915,N_5081);
nor U13443 (N_13443,N_9898,N_5711);
xnor U13444 (N_13444,N_7227,N_8695);
xnor U13445 (N_13445,N_9256,N_9775);
nor U13446 (N_13446,N_8906,N_7925);
nor U13447 (N_13447,N_7549,N_8747);
or U13448 (N_13448,N_7489,N_5382);
or U13449 (N_13449,N_6322,N_6137);
nand U13450 (N_13450,N_8864,N_6521);
or U13451 (N_13451,N_5403,N_9657);
nand U13452 (N_13452,N_9612,N_5205);
nor U13453 (N_13453,N_5685,N_7247);
xor U13454 (N_13454,N_5297,N_6552);
or U13455 (N_13455,N_5728,N_5236);
or U13456 (N_13456,N_5216,N_7867);
or U13457 (N_13457,N_8368,N_6895);
nor U13458 (N_13458,N_7935,N_9533);
and U13459 (N_13459,N_6661,N_8292);
nor U13460 (N_13460,N_8197,N_8979);
nor U13461 (N_13461,N_8343,N_9891);
and U13462 (N_13462,N_9005,N_5187);
nand U13463 (N_13463,N_9177,N_7729);
nand U13464 (N_13464,N_9786,N_5501);
or U13465 (N_13465,N_8900,N_9645);
and U13466 (N_13466,N_8574,N_8336);
or U13467 (N_13467,N_6131,N_5496);
xor U13468 (N_13468,N_9400,N_7366);
xnor U13469 (N_13469,N_8731,N_6001);
and U13470 (N_13470,N_7633,N_8404);
nor U13471 (N_13471,N_5686,N_8549);
xnor U13472 (N_13472,N_9537,N_9770);
and U13473 (N_13473,N_7533,N_5350);
or U13474 (N_13474,N_7081,N_9701);
nor U13475 (N_13475,N_6617,N_8738);
or U13476 (N_13476,N_6277,N_6040);
nor U13477 (N_13477,N_8390,N_6029);
nand U13478 (N_13478,N_5145,N_6088);
nor U13479 (N_13479,N_8254,N_7927);
nand U13480 (N_13480,N_8469,N_8864);
nor U13481 (N_13481,N_5676,N_5610);
nand U13482 (N_13482,N_5759,N_6852);
and U13483 (N_13483,N_5507,N_9263);
and U13484 (N_13484,N_5135,N_6814);
and U13485 (N_13485,N_9507,N_6775);
nand U13486 (N_13486,N_9897,N_6748);
nand U13487 (N_13487,N_9723,N_7432);
or U13488 (N_13488,N_9781,N_7037);
nand U13489 (N_13489,N_8401,N_6247);
or U13490 (N_13490,N_6001,N_7421);
or U13491 (N_13491,N_9064,N_5568);
nand U13492 (N_13492,N_6152,N_5549);
nor U13493 (N_13493,N_6499,N_9670);
and U13494 (N_13494,N_5235,N_5497);
xor U13495 (N_13495,N_5605,N_8531);
nand U13496 (N_13496,N_5615,N_8631);
and U13497 (N_13497,N_7027,N_9567);
and U13498 (N_13498,N_6541,N_5925);
and U13499 (N_13499,N_9636,N_6091);
xnor U13500 (N_13500,N_7194,N_8964);
nor U13501 (N_13501,N_7544,N_6424);
or U13502 (N_13502,N_5632,N_5907);
nor U13503 (N_13503,N_9533,N_5571);
and U13504 (N_13504,N_5450,N_6848);
and U13505 (N_13505,N_9480,N_5736);
xnor U13506 (N_13506,N_5508,N_5378);
and U13507 (N_13507,N_6077,N_8088);
nand U13508 (N_13508,N_9474,N_8921);
nor U13509 (N_13509,N_7918,N_6046);
nand U13510 (N_13510,N_8240,N_8673);
xnor U13511 (N_13511,N_7469,N_6110);
and U13512 (N_13512,N_6991,N_5071);
and U13513 (N_13513,N_7627,N_8494);
or U13514 (N_13514,N_7850,N_9662);
and U13515 (N_13515,N_6532,N_9983);
nor U13516 (N_13516,N_6107,N_5434);
and U13517 (N_13517,N_5485,N_5545);
and U13518 (N_13518,N_5605,N_5321);
xor U13519 (N_13519,N_9667,N_7048);
nor U13520 (N_13520,N_8287,N_9816);
xor U13521 (N_13521,N_8051,N_9303);
xnor U13522 (N_13522,N_8001,N_9028);
xnor U13523 (N_13523,N_5472,N_8054);
or U13524 (N_13524,N_8996,N_6224);
and U13525 (N_13525,N_7150,N_8042);
and U13526 (N_13526,N_9826,N_9541);
or U13527 (N_13527,N_5738,N_9023);
nor U13528 (N_13528,N_6363,N_7870);
nor U13529 (N_13529,N_7249,N_8700);
xnor U13530 (N_13530,N_5234,N_5511);
and U13531 (N_13531,N_9704,N_6803);
and U13532 (N_13532,N_7829,N_7948);
nand U13533 (N_13533,N_9111,N_6713);
nor U13534 (N_13534,N_8402,N_6311);
and U13535 (N_13535,N_5081,N_6554);
xnor U13536 (N_13536,N_7881,N_7373);
xor U13537 (N_13537,N_6767,N_7227);
nand U13538 (N_13538,N_8636,N_7634);
and U13539 (N_13539,N_7008,N_5206);
nand U13540 (N_13540,N_9987,N_7115);
xnor U13541 (N_13541,N_7017,N_8222);
nor U13542 (N_13542,N_8243,N_9658);
or U13543 (N_13543,N_5515,N_6393);
and U13544 (N_13544,N_9923,N_8473);
xor U13545 (N_13545,N_8278,N_5645);
or U13546 (N_13546,N_5659,N_8061);
xor U13547 (N_13547,N_5916,N_9241);
or U13548 (N_13548,N_8593,N_5868);
nor U13549 (N_13549,N_6144,N_7280);
nand U13550 (N_13550,N_9515,N_5848);
xnor U13551 (N_13551,N_5872,N_8504);
nand U13552 (N_13552,N_7012,N_9683);
nor U13553 (N_13553,N_7432,N_7527);
xnor U13554 (N_13554,N_5266,N_6854);
and U13555 (N_13555,N_9827,N_9522);
xor U13556 (N_13556,N_7791,N_5191);
nor U13557 (N_13557,N_6499,N_5277);
nand U13558 (N_13558,N_9492,N_6479);
xor U13559 (N_13559,N_6296,N_7199);
and U13560 (N_13560,N_5362,N_9136);
nor U13561 (N_13561,N_9300,N_6355);
xor U13562 (N_13562,N_9275,N_5008);
xor U13563 (N_13563,N_6923,N_7336);
nor U13564 (N_13564,N_6281,N_9934);
or U13565 (N_13565,N_9554,N_6159);
or U13566 (N_13566,N_9722,N_9314);
or U13567 (N_13567,N_8926,N_5215);
xor U13568 (N_13568,N_8881,N_6124);
and U13569 (N_13569,N_6448,N_7471);
nand U13570 (N_13570,N_8609,N_5299);
nor U13571 (N_13571,N_7070,N_5796);
or U13572 (N_13572,N_6596,N_8257);
nand U13573 (N_13573,N_6683,N_8576);
xnor U13574 (N_13574,N_6273,N_6973);
xnor U13575 (N_13575,N_5047,N_6485);
nor U13576 (N_13576,N_9671,N_6716);
nand U13577 (N_13577,N_7383,N_6048);
nor U13578 (N_13578,N_9709,N_5673);
nor U13579 (N_13579,N_6338,N_7972);
and U13580 (N_13580,N_7129,N_6382);
and U13581 (N_13581,N_6868,N_6528);
or U13582 (N_13582,N_6260,N_5100);
xnor U13583 (N_13583,N_5789,N_6205);
nand U13584 (N_13584,N_6278,N_8998);
xor U13585 (N_13585,N_7410,N_8988);
and U13586 (N_13586,N_7937,N_7600);
nor U13587 (N_13587,N_8524,N_7547);
and U13588 (N_13588,N_9498,N_9388);
and U13589 (N_13589,N_6945,N_9870);
nor U13590 (N_13590,N_5074,N_8622);
and U13591 (N_13591,N_5849,N_9199);
nor U13592 (N_13592,N_9390,N_6486);
and U13593 (N_13593,N_9393,N_8528);
xnor U13594 (N_13594,N_8469,N_6617);
and U13595 (N_13595,N_7629,N_7784);
xor U13596 (N_13596,N_6277,N_9595);
and U13597 (N_13597,N_9497,N_7487);
nor U13598 (N_13598,N_9607,N_6860);
nor U13599 (N_13599,N_5484,N_8799);
or U13600 (N_13600,N_7918,N_5205);
xnor U13601 (N_13601,N_8321,N_6665);
xor U13602 (N_13602,N_5170,N_7748);
nand U13603 (N_13603,N_8713,N_5027);
and U13604 (N_13604,N_7534,N_7188);
nand U13605 (N_13605,N_5463,N_7730);
nand U13606 (N_13606,N_7392,N_8679);
and U13607 (N_13607,N_8980,N_6931);
nand U13608 (N_13608,N_7389,N_7132);
nor U13609 (N_13609,N_8820,N_9799);
or U13610 (N_13610,N_9318,N_6735);
and U13611 (N_13611,N_9390,N_7900);
nor U13612 (N_13612,N_5538,N_9661);
or U13613 (N_13613,N_6483,N_5229);
or U13614 (N_13614,N_7278,N_5182);
nor U13615 (N_13615,N_5496,N_9745);
and U13616 (N_13616,N_9394,N_8072);
xor U13617 (N_13617,N_5180,N_8238);
xnor U13618 (N_13618,N_8053,N_6094);
and U13619 (N_13619,N_5390,N_5142);
xor U13620 (N_13620,N_9296,N_7635);
nand U13621 (N_13621,N_6891,N_5051);
nor U13622 (N_13622,N_8951,N_5179);
or U13623 (N_13623,N_6198,N_6525);
and U13624 (N_13624,N_9263,N_6035);
nand U13625 (N_13625,N_8251,N_5279);
nor U13626 (N_13626,N_5470,N_7524);
xor U13627 (N_13627,N_8237,N_6198);
nor U13628 (N_13628,N_8807,N_7768);
nor U13629 (N_13629,N_7700,N_8183);
nor U13630 (N_13630,N_6049,N_9492);
xor U13631 (N_13631,N_5125,N_6635);
and U13632 (N_13632,N_9522,N_8082);
xor U13633 (N_13633,N_9554,N_8002);
xnor U13634 (N_13634,N_6051,N_5766);
and U13635 (N_13635,N_8886,N_5299);
nand U13636 (N_13636,N_7739,N_9696);
and U13637 (N_13637,N_6157,N_8095);
nor U13638 (N_13638,N_5335,N_7793);
nand U13639 (N_13639,N_5969,N_5314);
nor U13640 (N_13640,N_7478,N_9669);
nor U13641 (N_13641,N_7570,N_9208);
xor U13642 (N_13642,N_9501,N_7341);
and U13643 (N_13643,N_5707,N_8585);
or U13644 (N_13644,N_8605,N_6738);
and U13645 (N_13645,N_6675,N_9563);
nor U13646 (N_13646,N_6988,N_5896);
or U13647 (N_13647,N_9316,N_7663);
xnor U13648 (N_13648,N_5186,N_5333);
or U13649 (N_13649,N_7575,N_8157);
or U13650 (N_13650,N_7050,N_5516);
and U13651 (N_13651,N_5545,N_5130);
nand U13652 (N_13652,N_5536,N_6322);
nand U13653 (N_13653,N_7996,N_6654);
and U13654 (N_13654,N_5160,N_9004);
or U13655 (N_13655,N_6706,N_9383);
and U13656 (N_13656,N_7471,N_9455);
xor U13657 (N_13657,N_9953,N_6851);
nor U13658 (N_13658,N_8010,N_5044);
and U13659 (N_13659,N_5319,N_5960);
or U13660 (N_13660,N_6619,N_5558);
xor U13661 (N_13661,N_9800,N_9324);
nor U13662 (N_13662,N_5937,N_7368);
xnor U13663 (N_13663,N_8776,N_6586);
or U13664 (N_13664,N_6520,N_5858);
or U13665 (N_13665,N_7911,N_6495);
or U13666 (N_13666,N_9210,N_7278);
or U13667 (N_13667,N_7601,N_7329);
xor U13668 (N_13668,N_9107,N_7269);
nand U13669 (N_13669,N_8303,N_9544);
or U13670 (N_13670,N_9562,N_6872);
nor U13671 (N_13671,N_9964,N_6642);
and U13672 (N_13672,N_8572,N_8683);
nor U13673 (N_13673,N_7234,N_7291);
or U13674 (N_13674,N_9178,N_8464);
or U13675 (N_13675,N_7946,N_6429);
nand U13676 (N_13676,N_5849,N_9050);
or U13677 (N_13677,N_8706,N_5918);
xor U13678 (N_13678,N_9317,N_7891);
nand U13679 (N_13679,N_8899,N_8204);
xnor U13680 (N_13680,N_6121,N_5140);
nor U13681 (N_13681,N_5320,N_6254);
and U13682 (N_13682,N_6552,N_6160);
and U13683 (N_13683,N_5019,N_7393);
or U13684 (N_13684,N_5470,N_7934);
nor U13685 (N_13685,N_8137,N_8946);
nand U13686 (N_13686,N_9060,N_9728);
nor U13687 (N_13687,N_7293,N_6157);
xor U13688 (N_13688,N_7601,N_5948);
and U13689 (N_13689,N_6543,N_5728);
nor U13690 (N_13690,N_7748,N_7119);
nand U13691 (N_13691,N_6260,N_8795);
xor U13692 (N_13692,N_7029,N_5699);
and U13693 (N_13693,N_6887,N_9504);
or U13694 (N_13694,N_6538,N_6150);
nand U13695 (N_13695,N_7675,N_7737);
or U13696 (N_13696,N_8096,N_7323);
and U13697 (N_13697,N_9323,N_6422);
nand U13698 (N_13698,N_9754,N_9303);
nand U13699 (N_13699,N_6317,N_8001);
or U13700 (N_13700,N_5863,N_5728);
xnor U13701 (N_13701,N_7148,N_5956);
xor U13702 (N_13702,N_5222,N_9797);
nand U13703 (N_13703,N_8459,N_5668);
or U13704 (N_13704,N_6974,N_5141);
nand U13705 (N_13705,N_9862,N_8337);
xor U13706 (N_13706,N_5501,N_5254);
xor U13707 (N_13707,N_5414,N_6287);
xor U13708 (N_13708,N_5419,N_8981);
xnor U13709 (N_13709,N_8351,N_8977);
or U13710 (N_13710,N_7423,N_8244);
nor U13711 (N_13711,N_6354,N_6077);
nor U13712 (N_13712,N_5797,N_9874);
xnor U13713 (N_13713,N_9350,N_8208);
and U13714 (N_13714,N_6257,N_5062);
or U13715 (N_13715,N_9909,N_9399);
nand U13716 (N_13716,N_6057,N_6932);
nor U13717 (N_13717,N_6366,N_9579);
and U13718 (N_13718,N_8645,N_6250);
or U13719 (N_13719,N_5692,N_9463);
and U13720 (N_13720,N_7903,N_9672);
xor U13721 (N_13721,N_9381,N_5161);
nor U13722 (N_13722,N_9165,N_9625);
or U13723 (N_13723,N_5743,N_8931);
nor U13724 (N_13724,N_5859,N_6225);
and U13725 (N_13725,N_5550,N_8527);
nand U13726 (N_13726,N_9010,N_5687);
xor U13727 (N_13727,N_5253,N_7603);
xor U13728 (N_13728,N_6797,N_6743);
nand U13729 (N_13729,N_9785,N_5919);
and U13730 (N_13730,N_6764,N_7158);
nor U13731 (N_13731,N_9530,N_9459);
nand U13732 (N_13732,N_5009,N_6941);
nand U13733 (N_13733,N_7035,N_5915);
or U13734 (N_13734,N_9061,N_7700);
or U13735 (N_13735,N_6828,N_7665);
xnor U13736 (N_13736,N_5857,N_8931);
and U13737 (N_13737,N_5173,N_5719);
nor U13738 (N_13738,N_9771,N_9307);
or U13739 (N_13739,N_8721,N_7440);
or U13740 (N_13740,N_6482,N_7400);
xor U13741 (N_13741,N_5980,N_9481);
xor U13742 (N_13742,N_9900,N_6258);
or U13743 (N_13743,N_9314,N_5762);
and U13744 (N_13744,N_6386,N_7001);
nor U13745 (N_13745,N_8159,N_8191);
and U13746 (N_13746,N_8755,N_6314);
xor U13747 (N_13747,N_5434,N_9544);
and U13748 (N_13748,N_7405,N_9498);
nand U13749 (N_13749,N_7211,N_7737);
nand U13750 (N_13750,N_8835,N_5965);
and U13751 (N_13751,N_9488,N_7692);
and U13752 (N_13752,N_5539,N_7258);
or U13753 (N_13753,N_8772,N_7825);
nand U13754 (N_13754,N_8755,N_5786);
nor U13755 (N_13755,N_5374,N_9080);
and U13756 (N_13756,N_8306,N_8273);
xnor U13757 (N_13757,N_6151,N_5192);
nor U13758 (N_13758,N_9920,N_5946);
nor U13759 (N_13759,N_7497,N_5758);
xnor U13760 (N_13760,N_7383,N_9375);
nand U13761 (N_13761,N_7698,N_5491);
and U13762 (N_13762,N_7594,N_5445);
xnor U13763 (N_13763,N_6140,N_8352);
and U13764 (N_13764,N_9766,N_5397);
nor U13765 (N_13765,N_9250,N_5832);
xor U13766 (N_13766,N_7822,N_5159);
or U13767 (N_13767,N_5825,N_9555);
and U13768 (N_13768,N_5036,N_8444);
or U13769 (N_13769,N_8264,N_5626);
nand U13770 (N_13770,N_8968,N_7353);
nor U13771 (N_13771,N_6347,N_5253);
xor U13772 (N_13772,N_9621,N_6714);
nor U13773 (N_13773,N_5070,N_8582);
or U13774 (N_13774,N_8392,N_7558);
and U13775 (N_13775,N_8861,N_6957);
nor U13776 (N_13776,N_5785,N_7631);
xor U13777 (N_13777,N_8843,N_8231);
or U13778 (N_13778,N_8931,N_7801);
nand U13779 (N_13779,N_5886,N_5705);
or U13780 (N_13780,N_8144,N_5151);
xor U13781 (N_13781,N_7720,N_8674);
and U13782 (N_13782,N_5812,N_8723);
xnor U13783 (N_13783,N_9264,N_6829);
nor U13784 (N_13784,N_6340,N_7513);
xnor U13785 (N_13785,N_9195,N_6431);
xor U13786 (N_13786,N_5230,N_7583);
and U13787 (N_13787,N_5861,N_5534);
nand U13788 (N_13788,N_7132,N_6697);
nand U13789 (N_13789,N_7175,N_6619);
and U13790 (N_13790,N_9946,N_8116);
or U13791 (N_13791,N_5605,N_8928);
and U13792 (N_13792,N_8135,N_5446);
nand U13793 (N_13793,N_5203,N_5837);
nor U13794 (N_13794,N_6972,N_8535);
nand U13795 (N_13795,N_5678,N_6963);
nor U13796 (N_13796,N_5493,N_9189);
nor U13797 (N_13797,N_6368,N_8104);
xnor U13798 (N_13798,N_7843,N_6073);
and U13799 (N_13799,N_9836,N_5374);
nor U13800 (N_13800,N_5274,N_9583);
xor U13801 (N_13801,N_9816,N_5712);
xor U13802 (N_13802,N_9205,N_6715);
nor U13803 (N_13803,N_9448,N_9499);
or U13804 (N_13804,N_9120,N_5795);
nor U13805 (N_13805,N_9334,N_5550);
xor U13806 (N_13806,N_8440,N_8983);
nor U13807 (N_13807,N_9333,N_5206);
nand U13808 (N_13808,N_8240,N_5588);
or U13809 (N_13809,N_9662,N_7599);
nand U13810 (N_13810,N_8882,N_8554);
nor U13811 (N_13811,N_5195,N_5673);
or U13812 (N_13812,N_9087,N_7046);
xor U13813 (N_13813,N_8731,N_7695);
xor U13814 (N_13814,N_6547,N_5618);
and U13815 (N_13815,N_8076,N_7974);
nand U13816 (N_13816,N_5263,N_8586);
nor U13817 (N_13817,N_5812,N_7196);
or U13818 (N_13818,N_5559,N_5689);
and U13819 (N_13819,N_7189,N_5208);
nand U13820 (N_13820,N_7340,N_8224);
or U13821 (N_13821,N_6231,N_5614);
xor U13822 (N_13822,N_9203,N_7371);
nand U13823 (N_13823,N_8543,N_9632);
nor U13824 (N_13824,N_7996,N_6295);
xnor U13825 (N_13825,N_8515,N_5382);
nor U13826 (N_13826,N_9629,N_6464);
nor U13827 (N_13827,N_8406,N_5220);
nand U13828 (N_13828,N_7053,N_8312);
nor U13829 (N_13829,N_8714,N_6292);
nor U13830 (N_13830,N_7884,N_8295);
or U13831 (N_13831,N_8049,N_7133);
xor U13832 (N_13832,N_9922,N_9631);
xor U13833 (N_13833,N_6326,N_8106);
nand U13834 (N_13834,N_7447,N_7183);
xnor U13835 (N_13835,N_5472,N_9800);
or U13836 (N_13836,N_5155,N_8512);
and U13837 (N_13837,N_6489,N_9416);
and U13838 (N_13838,N_7220,N_9911);
xor U13839 (N_13839,N_7331,N_5337);
nand U13840 (N_13840,N_6677,N_6201);
xnor U13841 (N_13841,N_8598,N_5946);
or U13842 (N_13842,N_9410,N_8852);
xnor U13843 (N_13843,N_8482,N_6341);
xnor U13844 (N_13844,N_9233,N_7569);
nor U13845 (N_13845,N_8898,N_9974);
or U13846 (N_13846,N_6267,N_5941);
and U13847 (N_13847,N_9359,N_7820);
xnor U13848 (N_13848,N_5182,N_5351);
or U13849 (N_13849,N_6659,N_5272);
and U13850 (N_13850,N_6524,N_7077);
and U13851 (N_13851,N_7043,N_9017);
nor U13852 (N_13852,N_9020,N_6031);
xnor U13853 (N_13853,N_7267,N_9102);
nor U13854 (N_13854,N_8449,N_7290);
nand U13855 (N_13855,N_9501,N_9040);
nand U13856 (N_13856,N_6828,N_8109);
nor U13857 (N_13857,N_8095,N_8888);
nand U13858 (N_13858,N_5308,N_7133);
xnor U13859 (N_13859,N_6737,N_5775);
xor U13860 (N_13860,N_6170,N_8187);
or U13861 (N_13861,N_5249,N_5745);
or U13862 (N_13862,N_9872,N_7859);
or U13863 (N_13863,N_6040,N_5861);
nor U13864 (N_13864,N_6451,N_7189);
or U13865 (N_13865,N_9794,N_9713);
nand U13866 (N_13866,N_7523,N_8719);
nand U13867 (N_13867,N_6676,N_8809);
nor U13868 (N_13868,N_9672,N_8269);
and U13869 (N_13869,N_6239,N_9364);
xnor U13870 (N_13870,N_5038,N_6342);
xnor U13871 (N_13871,N_8370,N_6147);
or U13872 (N_13872,N_5391,N_9690);
xnor U13873 (N_13873,N_8616,N_6009);
nor U13874 (N_13874,N_5053,N_5815);
or U13875 (N_13875,N_6187,N_9116);
and U13876 (N_13876,N_8292,N_8472);
nor U13877 (N_13877,N_7849,N_9415);
or U13878 (N_13878,N_6080,N_9826);
xnor U13879 (N_13879,N_8725,N_6447);
or U13880 (N_13880,N_6793,N_7378);
nor U13881 (N_13881,N_5395,N_7883);
nor U13882 (N_13882,N_8526,N_8754);
and U13883 (N_13883,N_7938,N_7344);
nand U13884 (N_13884,N_8603,N_9864);
nand U13885 (N_13885,N_7459,N_8398);
and U13886 (N_13886,N_9557,N_9838);
or U13887 (N_13887,N_7726,N_9596);
nand U13888 (N_13888,N_5912,N_6593);
nand U13889 (N_13889,N_7818,N_9572);
nor U13890 (N_13890,N_6804,N_9109);
or U13891 (N_13891,N_5169,N_7367);
nor U13892 (N_13892,N_7564,N_9178);
or U13893 (N_13893,N_6931,N_9821);
nor U13894 (N_13894,N_6941,N_8169);
nor U13895 (N_13895,N_9861,N_5446);
nor U13896 (N_13896,N_8958,N_6888);
nand U13897 (N_13897,N_5351,N_6368);
xor U13898 (N_13898,N_7648,N_9644);
nor U13899 (N_13899,N_5230,N_6465);
and U13900 (N_13900,N_5839,N_9673);
or U13901 (N_13901,N_5680,N_5180);
nor U13902 (N_13902,N_9637,N_6822);
nand U13903 (N_13903,N_9350,N_9257);
or U13904 (N_13904,N_7532,N_5314);
and U13905 (N_13905,N_6593,N_7464);
xnor U13906 (N_13906,N_5912,N_8369);
xor U13907 (N_13907,N_9939,N_8858);
nor U13908 (N_13908,N_9891,N_9416);
nor U13909 (N_13909,N_6699,N_5627);
xnor U13910 (N_13910,N_7924,N_6517);
nor U13911 (N_13911,N_6753,N_8668);
and U13912 (N_13912,N_7108,N_6321);
nand U13913 (N_13913,N_5581,N_7441);
and U13914 (N_13914,N_7693,N_7794);
xor U13915 (N_13915,N_9999,N_8717);
and U13916 (N_13916,N_8413,N_9235);
and U13917 (N_13917,N_5525,N_6364);
and U13918 (N_13918,N_9568,N_6064);
nor U13919 (N_13919,N_5705,N_8939);
nor U13920 (N_13920,N_5286,N_9920);
nand U13921 (N_13921,N_7510,N_9294);
xnor U13922 (N_13922,N_9573,N_9615);
xor U13923 (N_13923,N_6510,N_5784);
nand U13924 (N_13924,N_8652,N_6589);
nand U13925 (N_13925,N_5615,N_6366);
nor U13926 (N_13926,N_6488,N_8944);
nand U13927 (N_13927,N_7267,N_5682);
or U13928 (N_13928,N_6788,N_8316);
or U13929 (N_13929,N_6422,N_9116);
and U13930 (N_13930,N_8643,N_8886);
xor U13931 (N_13931,N_5448,N_6023);
nand U13932 (N_13932,N_5344,N_9704);
nor U13933 (N_13933,N_6289,N_5674);
nand U13934 (N_13934,N_9121,N_9740);
or U13935 (N_13935,N_5832,N_7132);
nor U13936 (N_13936,N_9750,N_6776);
nor U13937 (N_13937,N_8234,N_7932);
or U13938 (N_13938,N_5279,N_9373);
nor U13939 (N_13939,N_8639,N_8960);
and U13940 (N_13940,N_8486,N_6397);
and U13941 (N_13941,N_6957,N_8753);
and U13942 (N_13942,N_6869,N_5050);
nand U13943 (N_13943,N_9974,N_7497);
and U13944 (N_13944,N_5470,N_7699);
nor U13945 (N_13945,N_8784,N_6960);
and U13946 (N_13946,N_8290,N_6818);
nor U13947 (N_13947,N_7606,N_9676);
and U13948 (N_13948,N_5998,N_8871);
nor U13949 (N_13949,N_6419,N_6329);
nand U13950 (N_13950,N_6505,N_8028);
xor U13951 (N_13951,N_6957,N_9811);
nand U13952 (N_13952,N_8222,N_9210);
nand U13953 (N_13953,N_7135,N_9922);
nor U13954 (N_13954,N_7895,N_9562);
and U13955 (N_13955,N_9484,N_7171);
or U13956 (N_13956,N_9796,N_8109);
nand U13957 (N_13957,N_9054,N_7078);
or U13958 (N_13958,N_6791,N_8063);
or U13959 (N_13959,N_8577,N_6565);
or U13960 (N_13960,N_5212,N_8315);
nand U13961 (N_13961,N_7433,N_5484);
or U13962 (N_13962,N_8265,N_6765);
nand U13963 (N_13963,N_7319,N_5579);
and U13964 (N_13964,N_5506,N_5903);
and U13965 (N_13965,N_8496,N_7795);
nor U13966 (N_13966,N_6104,N_8246);
and U13967 (N_13967,N_7941,N_9692);
nand U13968 (N_13968,N_7406,N_6068);
and U13969 (N_13969,N_7187,N_8890);
xnor U13970 (N_13970,N_8467,N_9086);
or U13971 (N_13971,N_8163,N_6788);
nor U13972 (N_13972,N_5948,N_8538);
nor U13973 (N_13973,N_7644,N_8861);
or U13974 (N_13974,N_8012,N_6692);
xor U13975 (N_13975,N_8586,N_9473);
nor U13976 (N_13976,N_8133,N_6605);
and U13977 (N_13977,N_6451,N_9069);
or U13978 (N_13978,N_9178,N_7397);
nand U13979 (N_13979,N_8951,N_6016);
nor U13980 (N_13980,N_6478,N_5148);
or U13981 (N_13981,N_9926,N_6999);
and U13982 (N_13982,N_5257,N_5013);
nand U13983 (N_13983,N_7461,N_7840);
nor U13984 (N_13984,N_5489,N_7729);
xnor U13985 (N_13985,N_6905,N_6615);
and U13986 (N_13986,N_8672,N_6004);
or U13987 (N_13987,N_7940,N_8604);
xnor U13988 (N_13988,N_9289,N_7857);
and U13989 (N_13989,N_9443,N_5671);
xnor U13990 (N_13990,N_8993,N_9577);
nand U13991 (N_13991,N_9645,N_7278);
or U13992 (N_13992,N_6561,N_8540);
and U13993 (N_13993,N_7792,N_7094);
nor U13994 (N_13994,N_5346,N_6797);
xor U13995 (N_13995,N_9733,N_7514);
or U13996 (N_13996,N_6247,N_6271);
xnor U13997 (N_13997,N_7261,N_6949);
xnor U13998 (N_13998,N_9742,N_7717);
nor U13999 (N_13999,N_6673,N_6900);
and U14000 (N_14000,N_5654,N_5643);
xor U14001 (N_14001,N_5778,N_5270);
nor U14002 (N_14002,N_5159,N_6022);
xor U14003 (N_14003,N_5744,N_7386);
nand U14004 (N_14004,N_7538,N_9400);
and U14005 (N_14005,N_5224,N_7832);
and U14006 (N_14006,N_9425,N_8345);
xor U14007 (N_14007,N_6051,N_8017);
and U14008 (N_14008,N_9812,N_9744);
xnor U14009 (N_14009,N_8328,N_9771);
nand U14010 (N_14010,N_5976,N_7646);
and U14011 (N_14011,N_9493,N_5444);
nor U14012 (N_14012,N_8306,N_6370);
xor U14013 (N_14013,N_8215,N_5317);
and U14014 (N_14014,N_6399,N_9705);
or U14015 (N_14015,N_5774,N_7292);
nor U14016 (N_14016,N_6935,N_6434);
and U14017 (N_14017,N_9126,N_5430);
xor U14018 (N_14018,N_8091,N_6012);
xor U14019 (N_14019,N_6664,N_6371);
nand U14020 (N_14020,N_9654,N_8775);
nand U14021 (N_14021,N_7309,N_8389);
or U14022 (N_14022,N_9898,N_6481);
or U14023 (N_14023,N_5999,N_6706);
and U14024 (N_14024,N_9597,N_9925);
nand U14025 (N_14025,N_9857,N_5847);
or U14026 (N_14026,N_6834,N_9149);
xnor U14027 (N_14027,N_6069,N_9769);
nor U14028 (N_14028,N_5670,N_6497);
nor U14029 (N_14029,N_6990,N_5201);
nand U14030 (N_14030,N_9890,N_8139);
nor U14031 (N_14031,N_8170,N_9117);
nor U14032 (N_14032,N_9580,N_8369);
xnor U14033 (N_14033,N_9047,N_6575);
nand U14034 (N_14034,N_9146,N_7538);
and U14035 (N_14035,N_6385,N_5649);
or U14036 (N_14036,N_9261,N_8801);
xnor U14037 (N_14037,N_6491,N_5921);
or U14038 (N_14038,N_5935,N_5922);
nand U14039 (N_14039,N_7454,N_8718);
nor U14040 (N_14040,N_7407,N_8001);
nor U14041 (N_14041,N_6747,N_7405);
or U14042 (N_14042,N_9740,N_9512);
or U14043 (N_14043,N_7284,N_6119);
nor U14044 (N_14044,N_9899,N_8100);
nor U14045 (N_14045,N_5088,N_7413);
xnor U14046 (N_14046,N_6201,N_9133);
and U14047 (N_14047,N_9025,N_8162);
and U14048 (N_14048,N_9904,N_7398);
or U14049 (N_14049,N_8352,N_9201);
or U14050 (N_14050,N_8890,N_5527);
nand U14051 (N_14051,N_6600,N_8869);
and U14052 (N_14052,N_9547,N_7759);
and U14053 (N_14053,N_9731,N_9090);
and U14054 (N_14054,N_7828,N_8907);
nor U14055 (N_14055,N_7054,N_5700);
and U14056 (N_14056,N_7019,N_6779);
nand U14057 (N_14057,N_9598,N_8615);
nand U14058 (N_14058,N_9215,N_5930);
xnor U14059 (N_14059,N_7636,N_8931);
and U14060 (N_14060,N_8371,N_6002);
xnor U14061 (N_14061,N_5882,N_5141);
xnor U14062 (N_14062,N_5761,N_6168);
nor U14063 (N_14063,N_6310,N_8520);
and U14064 (N_14064,N_6246,N_7529);
and U14065 (N_14065,N_7895,N_9724);
nand U14066 (N_14066,N_7528,N_5719);
or U14067 (N_14067,N_5296,N_6017);
nand U14068 (N_14068,N_6435,N_7174);
xnor U14069 (N_14069,N_8123,N_6636);
nor U14070 (N_14070,N_9273,N_7506);
nand U14071 (N_14071,N_5197,N_5386);
nand U14072 (N_14072,N_5982,N_8487);
or U14073 (N_14073,N_5457,N_8959);
and U14074 (N_14074,N_8612,N_8566);
nor U14075 (N_14075,N_5155,N_7219);
nor U14076 (N_14076,N_6827,N_5025);
and U14077 (N_14077,N_9995,N_6716);
nand U14078 (N_14078,N_9081,N_8525);
and U14079 (N_14079,N_9129,N_8794);
nand U14080 (N_14080,N_7701,N_9465);
xnor U14081 (N_14081,N_5852,N_7692);
nand U14082 (N_14082,N_5016,N_5632);
nand U14083 (N_14083,N_8623,N_5767);
xnor U14084 (N_14084,N_8988,N_6103);
or U14085 (N_14085,N_5033,N_7473);
nand U14086 (N_14086,N_5629,N_6509);
or U14087 (N_14087,N_5755,N_9170);
nor U14088 (N_14088,N_5483,N_7501);
xnor U14089 (N_14089,N_8618,N_6734);
nor U14090 (N_14090,N_7839,N_5249);
or U14091 (N_14091,N_7722,N_5852);
nand U14092 (N_14092,N_7479,N_6078);
nor U14093 (N_14093,N_6290,N_6560);
nor U14094 (N_14094,N_7206,N_9124);
and U14095 (N_14095,N_5620,N_5401);
xor U14096 (N_14096,N_6716,N_7376);
xor U14097 (N_14097,N_9783,N_6237);
nand U14098 (N_14098,N_5529,N_8673);
xnor U14099 (N_14099,N_9669,N_9517);
nor U14100 (N_14100,N_9604,N_5783);
xnor U14101 (N_14101,N_5429,N_9642);
and U14102 (N_14102,N_5078,N_8768);
xnor U14103 (N_14103,N_8440,N_6195);
or U14104 (N_14104,N_7648,N_5753);
xnor U14105 (N_14105,N_9871,N_9999);
nand U14106 (N_14106,N_5249,N_8567);
nor U14107 (N_14107,N_8761,N_7933);
nand U14108 (N_14108,N_6438,N_5054);
nand U14109 (N_14109,N_6992,N_8510);
nand U14110 (N_14110,N_9666,N_6508);
nand U14111 (N_14111,N_6716,N_5408);
xor U14112 (N_14112,N_9535,N_8927);
nor U14113 (N_14113,N_8166,N_6822);
nor U14114 (N_14114,N_5193,N_7087);
and U14115 (N_14115,N_5193,N_7639);
nand U14116 (N_14116,N_8531,N_6050);
nand U14117 (N_14117,N_6490,N_6521);
and U14118 (N_14118,N_8408,N_9960);
nand U14119 (N_14119,N_7452,N_5407);
nor U14120 (N_14120,N_8408,N_9597);
and U14121 (N_14121,N_5409,N_9426);
and U14122 (N_14122,N_8940,N_9479);
nor U14123 (N_14123,N_8267,N_6530);
or U14124 (N_14124,N_5669,N_9292);
nor U14125 (N_14125,N_6958,N_9715);
nor U14126 (N_14126,N_5116,N_6735);
nor U14127 (N_14127,N_7927,N_9530);
xnor U14128 (N_14128,N_9633,N_5413);
xnor U14129 (N_14129,N_9298,N_9526);
nor U14130 (N_14130,N_9051,N_6858);
xnor U14131 (N_14131,N_7085,N_5309);
or U14132 (N_14132,N_5237,N_6603);
and U14133 (N_14133,N_6164,N_7822);
and U14134 (N_14134,N_5118,N_8623);
or U14135 (N_14135,N_7289,N_7755);
and U14136 (N_14136,N_8958,N_8653);
and U14137 (N_14137,N_6151,N_6767);
or U14138 (N_14138,N_9736,N_6054);
nor U14139 (N_14139,N_6303,N_9669);
or U14140 (N_14140,N_5841,N_5303);
xnor U14141 (N_14141,N_5974,N_8306);
and U14142 (N_14142,N_9967,N_6091);
nor U14143 (N_14143,N_6101,N_8628);
nand U14144 (N_14144,N_8134,N_8447);
nand U14145 (N_14145,N_8761,N_8633);
nor U14146 (N_14146,N_5989,N_6340);
and U14147 (N_14147,N_6355,N_7000);
or U14148 (N_14148,N_9274,N_6837);
and U14149 (N_14149,N_6950,N_8690);
nor U14150 (N_14150,N_9790,N_5158);
and U14151 (N_14151,N_8858,N_7470);
nor U14152 (N_14152,N_8368,N_8027);
nor U14153 (N_14153,N_8708,N_8242);
nor U14154 (N_14154,N_7301,N_8414);
or U14155 (N_14155,N_5179,N_9780);
and U14156 (N_14156,N_7633,N_5574);
nand U14157 (N_14157,N_7199,N_8403);
xor U14158 (N_14158,N_8797,N_5383);
xnor U14159 (N_14159,N_6285,N_7041);
xnor U14160 (N_14160,N_5456,N_6282);
xor U14161 (N_14161,N_5023,N_6972);
nor U14162 (N_14162,N_9689,N_9676);
xnor U14163 (N_14163,N_8611,N_9767);
nor U14164 (N_14164,N_7027,N_8947);
nand U14165 (N_14165,N_6067,N_7223);
or U14166 (N_14166,N_6564,N_8549);
nor U14167 (N_14167,N_7454,N_7010);
xor U14168 (N_14168,N_7277,N_8394);
or U14169 (N_14169,N_6539,N_9414);
nor U14170 (N_14170,N_8493,N_9314);
xor U14171 (N_14171,N_6068,N_8435);
or U14172 (N_14172,N_5270,N_9222);
nor U14173 (N_14173,N_5082,N_9808);
nor U14174 (N_14174,N_8861,N_7986);
nor U14175 (N_14175,N_5325,N_9865);
and U14176 (N_14176,N_7822,N_6286);
or U14177 (N_14177,N_6734,N_5516);
nand U14178 (N_14178,N_8456,N_5906);
nand U14179 (N_14179,N_8663,N_6151);
or U14180 (N_14180,N_9682,N_9123);
and U14181 (N_14181,N_9656,N_6212);
xnor U14182 (N_14182,N_5252,N_6620);
nor U14183 (N_14183,N_8180,N_8383);
xor U14184 (N_14184,N_6663,N_8206);
nand U14185 (N_14185,N_6411,N_5035);
xor U14186 (N_14186,N_9237,N_7914);
or U14187 (N_14187,N_5338,N_9936);
xnor U14188 (N_14188,N_7541,N_7970);
or U14189 (N_14189,N_8597,N_7160);
and U14190 (N_14190,N_7836,N_6910);
xor U14191 (N_14191,N_7766,N_7820);
and U14192 (N_14192,N_6120,N_5197);
nand U14193 (N_14193,N_6092,N_8672);
nand U14194 (N_14194,N_5471,N_8236);
and U14195 (N_14195,N_7650,N_6229);
nor U14196 (N_14196,N_8041,N_8620);
nor U14197 (N_14197,N_7674,N_8330);
and U14198 (N_14198,N_7870,N_6984);
or U14199 (N_14199,N_8820,N_5691);
and U14200 (N_14200,N_7892,N_6950);
xor U14201 (N_14201,N_8512,N_6698);
nor U14202 (N_14202,N_6560,N_8584);
nand U14203 (N_14203,N_9535,N_7792);
or U14204 (N_14204,N_8128,N_5164);
and U14205 (N_14205,N_5783,N_9201);
or U14206 (N_14206,N_5967,N_9422);
nand U14207 (N_14207,N_5252,N_5778);
nand U14208 (N_14208,N_5550,N_5685);
xnor U14209 (N_14209,N_5994,N_6927);
xor U14210 (N_14210,N_8530,N_5934);
nor U14211 (N_14211,N_6753,N_6950);
and U14212 (N_14212,N_7517,N_7780);
xnor U14213 (N_14213,N_6250,N_6640);
or U14214 (N_14214,N_6726,N_5392);
and U14215 (N_14215,N_7096,N_9527);
and U14216 (N_14216,N_9000,N_6272);
or U14217 (N_14217,N_7466,N_5959);
or U14218 (N_14218,N_5625,N_9485);
xnor U14219 (N_14219,N_9362,N_8472);
nand U14220 (N_14220,N_9188,N_7625);
nand U14221 (N_14221,N_9458,N_6491);
or U14222 (N_14222,N_5771,N_7103);
nor U14223 (N_14223,N_7395,N_9313);
xor U14224 (N_14224,N_6730,N_5424);
or U14225 (N_14225,N_8621,N_8194);
xor U14226 (N_14226,N_6607,N_9750);
xor U14227 (N_14227,N_7354,N_5526);
nor U14228 (N_14228,N_8805,N_7073);
nand U14229 (N_14229,N_7250,N_7369);
nor U14230 (N_14230,N_7175,N_5924);
xor U14231 (N_14231,N_6815,N_9410);
nor U14232 (N_14232,N_7861,N_6312);
nor U14233 (N_14233,N_9207,N_9357);
nand U14234 (N_14234,N_6016,N_5876);
nand U14235 (N_14235,N_6669,N_5051);
or U14236 (N_14236,N_6120,N_8794);
nand U14237 (N_14237,N_6730,N_6847);
xnor U14238 (N_14238,N_8933,N_5089);
xor U14239 (N_14239,N_9008,N_6908);
xnor U14240 (N_14240,N_8830,N_6173);
or U14241 (N_14241,N_9302,N_9041);
nand U14242 (N_14242,N_5405,N_7257);
nor U14243 (N_14243,N_8817,N_7130);
nor U14244 (N_14244,N_6764,N_9159);
or U14245 (N_14245,N_8743,N_5392);
nor U14246 (N_14246,N_8028,N_6312);
xor U14247 (N_14247,N_9418,N_6227);
or U14248 (N_14248,N_6252,N_6806);
xor U14249 (N_14249,N_7402,N_5026);
nand U14250 (N_14250,N_6226,N_8816);
xnor U14251 (N_14251,N_5205,N_9946);
nand U14252 (N_14252,N_6868,N_9248);
or U14253 (N_14253,N_7017,N_9003);
nand U14254 (N_14254,N_7059,N_8042);
nor U14255 (N_14255,N_6336,N_7812);
nand U14256 (N_14256,N_7230,N_7117);
nor U14257 (N_14257,N_5220,N_5856);
or U14258 (N_14258,N_6420,N_8743);
and U14259 (N_14259,N_9655,N_6881);
and U14260 (N_14260,N_9992,N_7758);
xor U14261 (N_14261,N_8247,N_5030);
or U14262 (N_14262,N_6811,N_9560);
xnor U14263 (N_14263,N_8734,N_5562);
xnor U14264 (N_14264,N_6988,N_7316);
xnor U14265 (N_14265,N_5414,N_5541);
nor U14266 (N_14266,N_7752,N_8225);
and U14267 (N_14267,N_6566,N_9002);
nor U14268 (N_14268,N_8799,N_9248);
nor U14269 (N_14269,N_7747,N_8441);
nand U14270 (N_14270,N_8951,N_6764);
or U14271 (N_14271,N_5455,N_5264);
and U14272 (N_14272,N_8275,N_5201);
xor U14273 (N_14273,N_9510,N_6659);
and U14274 (N_14274,N_7445,N_9141);
xnor U14275 (N_14275,N_5121,N_6022);
or U14276 (N_14276,N_5821,N_6961);
nor U14277 (N_14277,N_5453,N_7491);
xor U14278 (N_14278,N_6344,N_9676);
xnor U14279 (N_14279,N_6862,N_6697);
nor U14280 (N_14280,N_8513,N_7705);
and U14281 (N_14281,N_7228,N_7297);
or U14282 (N_14282,N_5273,N_5051);
or U14283 (N_14283,N_5194,N_7699);
nor U14284 (N_14284,N_8745,N_7495);
xor U14285 (N_14285,N_5043,N_6938);
or U14286 (N_14286,N_5723,N_5752);
nor U14287 (N_14287,N_9904,N_8521);
nor U14288 (N_14288,N_6868,N_6747);
or U14289 (N_14289,N_6692,N_8157);
nor U14290 (N_14290,N_8036,N_8851);
nor U14291 (N_14291,N_6240,N_5168);
xor U14292 (N_14292,N_8986,N_8157);
nand U14293 (N_14293,N_8963,N_7735);
xor U14294 (N_14294,N_6200,N_7517);
or U14295 (N_14295,N_5896,N_9491);
xor U14296 (N_14296,N_9745,N_8002);
and U14297 (N_14297,N_6779,N_7926);
and U14298 (N_14298,N_8473,N_8293);
nor U14299 (N_14299,N_7198,N_8244);
and U14300 (N_14300,N_8719,N_5765);
and U14301 (N_14301,N_6093,N_6953);
or U14302 (N_14302,N_6066,N_5940);
nor U14303 (N_14303,N_5657,N_5924);
nor U14304 (N_14304,N_5727,N_6664);
or U14305 (N_14305,N_6531,N_7756);
xnor U14306 (N_14306,N_9771,N_6276);
nor U14307 (N_14307,N_8415,N_9170);
nor U14308 (N_14308,N_6617,N_8481);
nor U14309 (N_14309,N_9605,N_5852);
nor U14310 (N_14310,N_7182,N_5407);
and U14311 (N_14311,N_7472,N_7571);
nand U14312 (N_14312,N_8882,N_8165);
xor U14313 (N_14313,N_7389,N_8924);
and U14314 (N_14314,N_9631,N_7398);
and U14315 (N_14315,N_5118,N_8948);
and U14316 (N_14316,N_8150,N_9232);
xnor U14317 (N_14317,N_6852,N_7074);
or U14318 (N_14318,N_7320,N_7862);
or U14319 (N_14319,N_5158,N_8322);
or U14320 (N_14320,N_6245,N_5767);
nor U14321 (N_14321,N_7878,N_8589);
xnor U14322 (N_14322,N_8693,N_9823);
or U14323 (N_14323,N_6389,N_7683);
or U14324 (N_14324,N_7910,N_7541);
or U14325 (N_14325,N_5343,N_5338);
and U14326 (N_14326,N_8227,N_5682);
and U14327 (N_14327,N_6740,N_7973);
or U14328 (N_14328,N_5729,N_5291);
nor U14329 (N_14329,N_6132,N_8192);
xnor U14330 (N_14330,N_9508,N_9039);
nand U14331 (N_14331,N_9322,N_5826);
xor U14332 (N_14332,N_9295,N_8726);
or U14333 (N_14333,N_5259,N_6183);
xor U14334 (N_14334,N_9856,N_9120);
and U14335 (N_14335,N_5941,N_5625);
nand U14336 (N_14336,N_7963,N_9033);
or U14337 (N_14337,N_9842,N_7627);
nor U14338 (N_14338,N_5267,N_7792);
and U14339 (N_14339,N_9348,N_6750);
xnor U14340 (N_14340,N_8515,N_6068);
nor U14341 (N_14341,N_5420,N_9876);
nand U14342 (N_14342,N_9289,N_8440);
or U14343 (N_14343,N_6097,N_8572);
and U14344 (N_14344,N_5207,N_9448);
xor U14345 (N_14345,N_8655,N_8881);
nor U14346 (N_14346,N_7529,N_9777);
xnor U14347 (N_14347,N_5809,N_9090);
and U14348 (N_14348,N_8640,N_6760);
nand U14349 (N_14349,N_8670,N_8247);
nand U14350 (N_14350,N_6938,N_5256);
nor U14351 (N_14351,N_8783,N_8076);
nor U14352 (N_14352,N_8251,N_7004);
nand U14353 (N_14353,N_7135,N_6843);
xor U14354 (N_14354,N_7449,N_7234);
xor U14355 (N_14355,N_9831,N_8747);
nor U14356 (N_14356,N_8753,N_6679);
nand U14357 (N_14357,N_6103,N_6529);
nor U14358 (N_14358,N_9100,N_7182);
nand U14359 (N_14359,N_7839,N_6293);
or U14360 (N_14360,N_7925,N_9281);
xor U14361 (N_14361,N_9252,N_9791);
xor U14362 (N_14362,N_8514,N_5912);
nor U14363 (N_14363,N_7468,N_9911);
or U14364 (N_14364,N_7496,N_6938);
xor U14365 (N_14365,N_8941,N_6821);
nand U14366 (N_14366,N_6586,N_8403);
nand U14367 (N_14367,N_8449,N_6119);
nand U14368 (N_14368,N_8333,N_6037);
or U14369 (N_14369,N_5816,N_7088);
or U14370 (N_14370,N_7923,N_9343);
xnor U14371 (N_14371,N_7091,N_7349);
or U14372 (N_14372,N_6953,N_8626);
xor U14373 (N_14373,N_8674,N_6263);
or U14374 (N_14374,N_7131,N_8513);
nand U14375 (N_14375,N_8043,N_8297);
nand U14376 (N_14376,N_6266,N_7237);
nand U14377 (N_14377,N_7375,N_9877);
and U14378 (N_14378,N_9207,N_5734);
nor U14379 (N_14379,N_9274,N_6059);
xnor U14380 (N_14380,N_5722,N_5138);
nand U14381 (N_14381,N_9592,N_8261);
or U14382 (N_14382,N_8265,N_9067);
nand U14383 (N_14383,N_8757,N_7111);
xor U14384 (N_14384,N_9445,N_8715);
xnor U14385 (N_14385,N_9565,N_6335);
nand U14386 (N_14386,N_5632,N_7065);
nor U14387 (N_14387,N_6168,N_5809);
and U14388 (N_14388,N_6992,N_8178);
or U14389 (N_14389,N_8839,N_9620);
and U14390 (N_14390,N_7767,N_6373);
and U14391 (N_14391,N_7292,N_7030);
and U14392 (N_14392,N_8991,N_8726);
nand U14393 (N_14393,N_8176,N_5349);
or U14394 (N_14394,N_5657,N_9439);
or U14395 (N_14395,N_8963,N_6817);
xnor U14396 (N_14396,N_6706,N_9591);
or U14397 (N_14397,N_5434,N_8822);
or U14398 (N_14398,N_5281,N_7062);
nand U14399 (N_14399,N_5267,N_8915);
xnor U14400 (N_14400,N_8656,N_7838);
or U14401 (N_14401,N_8087,N_7877);
or U14402 (N_14402,N_8107,N_5200);
and U14403 (N_14403,N_5869,N_8335);
nand U14404 (N_14404,N_5854,N_8111);
and U14405 (N_14405,N_5611,N_5730);
nand U14406 (N_14406,N_6663,N_9377);
xnor U14407 (N_14407,N_8382,N_6587);
or U14408 (N_14408,N_7551,N_9679);
xnor U14409 (N_14409,N_9621,N_8866);
nor U14410 (N_14410,N_6972,N_5933);
nand U14411 (N_14411,N_8048,N_5248);
and U14412 (N_14412,N_8940,N_9773);
and U14413 (N_14413,N_5949,N_7727);
nand U14414 (N_14414,N_8036,N_6225);
nand U14415 (N_14415,N_5610,N_6138);
and U14416 (N_14416,N_6027,N_8024);
nor U14417 (N_14417,N_7678,N_8661);
and U14418 (N_14418,N_6946,N_5939);
or U14419 (N_14419,N_8022,N_9599);
or U14420 (N_14420,N_5788,N_7470);
nor U14421 (N_14421,N_8056,N_9785);
xnor U14422 (N_14422,N_5078,N_7648);
nand U14423 (N_14423,N_6351,N_9627);
xnor U14424 (N_14424,N_5331,N_7831);
nor U14425 (N_14425,N_6919,N_5146);
nor U14426 (N_14426,N_6139,N_9446);
nand U14427 (N_14427,N_9745,N_5620);
xor U14428 (N_14428,N_8994,N_5428);
nand U14429 (N_14429,N_7095,N_6168);
nor U14430 (N_14430,N_5086,N_8074);
nand U14431 (N_14431,N_8710,N_6015);
nand U14432 (N_14432,N_9758,N_5229);
nor U14433 (N_14433,N_9724,N_8652);
or U14434 (N_14434,N_5631,N_6905);
xor U14435 (N_14435,N_7795,N_5647);
and U14436 (N_14436,N_9162,N_5690);
and U14437 (N_14437,N_7834,N_7142);
xnor U14438 (N_14438,N_9632,N_6654);
and U14439 (N_14439,N_8193,N_9266);
xnor U14440 (N_14440,N_6603,N_5993);
or U14441 (N_14441,N_8665,N_6452);
or U14442 (N_14442,N_5536,N_5443);
xnor U14443 (N_14443,N_5018,N_9723);
or U14444 (N_14444,N_6051,N_7616);
nand U14445 (N_14445,N_9956,N_9042);
nand U14446 (N_14446,N_9300,N_9416);
nand U14447 (N_14447,N_8152,N_5884);
nor U14448 (N_14448,N_6786,N_8838);
and U14449 (N_14449,N_7592,N_7455);
xnor U14450 (N_14450,N_8094,N_6061);
or U14451 (N_14451,N_9358,N_7552);
nor U14452 (N_14452,N_7467,N_6420);
nor U14453 (N_14453,N_6026,N_8029);
or U14454 (N_14454,N_7012,N_9693);
nand U14455 (N_14455,N_8551,N_8039);
and U14456 (N_14456,N_5665,N_9090);
or U14457 (N_14457,N_5530,N_8103);
nand U14458 (N_14458,N_9045,N_7648);
and U14459 (N_14459,N_5141,N_5797);
nor U14460 (N_14460,N_7782,N_8119);
nand U14461 (N_14461,N_6138,N_6934);
xor U14462 (N_14462,N_9292,N_8606);
nor U14463 (N_14463,N_7516,N_8843);
or U14464 (N_14464,N_5505,N_6461);
or U14465 (N_14465,N_8387,N_6535);
nand U14466 (N_14466,N_5682,N_8688);
xor U14467 (N_14467,N_5114,N_8067);
nor U14468 (N_14468,N_5381,N_9582);
and U14469 (N_14469,N_9470,N_7818);
nand U14470 (N_14470,N_7328,N_9856);
nor U14471 (N_14471,N_8105,N_9661);
and U14472 (N_14472,N_5080,N_6660);
xor U14473 (N_14473,N_6701,N_5227);
xor U14474 (N_14474,N_8170,N_8470);
or U14475 (N_14475,N_6413,N_7473);
nor U14476 (N_14476,N_7792,N_5429);
nor U14477 (N_14477,N_5395,N_6110);
nor U14478 (N_14478,N_9910,N_6971);
nand U14479 (N_14479,N_9042,N_6532);
and U14480 (N_14480,N_6964,N_7492);
or U14481 (N_14481,N_5390,N_5572);
and U14482 (N_14482,N_9539,N_8262);
and U14483 (N_14483,N_6607,N_5437);
xor U14484 (N_14484,N_5595,N_8665);
nand U14485 (N_14485,N_6889,N_5122);
and U14486 (N_14486,N_9476,N_6701);
nand U14487 (N_14487,N_5907,N_6456);
and U14488 (N_14488,N_5418,N_7378);
or U14489 (N_14489,N_6146,N_9527);
nor U14490 (N_14490,N_8867,N_8714);
nor U14491 (N_14491,N_8228,N_7095);
nor U14492 (N_14492,N_5886,N_6995);
or U14493 (N_14493,N_5345,N_9477);
or U14494 (N_14494,N_6436,N_5191);
nand U14495 (N_14495,N_8030,N_9391);
or U14496 (N_14496,N_6391,N_8178);
nand U14497 (N_14497,N_6949,N_8379);
nand U14498 (N_14498,N_8395,N_5578);
nand U14499 (N_14499,N_5798,N_6658);
xor U14500 (N_14500,N_9780,N_8844);
xnor U14501 (N_14501,N_5889,N_9911);
and U14502 (N_14502,N_9633,N_8679);
nand U14503 (N_14503,N_9581,N_7133);
and U14504 (N_14504,N_8733,N_7917);
xor U14505 (N_14505,N_6420,N_8072);
and U14506 (N_14506,N_8700,N_8097);
or U14507 (N_14507,N_7725,N_9930);
or U14508 (N_14508,N_7587,N_9515);
xor U14509 (N_14509,N_7452,N_9674);
or U14510 (N_14510,N_6383,N_7722);
nand U14511 (N_14511,N_8497,N_8248);
or U14512 (N_14512,N_6507,N_6398);
or U14513 (N_14513,N_5421,N_6350);
and U14514 (N_14514,N_5214,N_7036);
and U14515 (N_14515,N_7407,N_7092);
and U14516 (N_14516,N_5917,N_5974);
nor U14517 (N_14517,N_7512,N_6208);
and U14518 (N_14518,N_6418,N_5527);
or U14519 (N_14519,N_9205,N_7635);
or U14520 (N_14520,N_8993,N_7713);
or U14521 (N_14521,N_6770,N_6007);
or U14522 (N_14522,N_8323,N_6725);
and U14523 (N_14523,N_5127,N_5335);
nand U14524 (N_14524,N_7242,N_7334);
nor U14525 (N_14525,N_6190,N_5040);
or U14526 (N_14526,N_9533,N_8751);
nand U14527 (N_14527,N_9810,N_6789);
nand U14528 (N_14528,N_9267,N_6982);
xnor U14529 (N_14529,N_7436,N_8915);
xnor U14530 (N_14530,N_7531,N_9372);
nor U14531 (N_14531,N_7077,N_7977);
and U14532 (N_14532,N_7144,N_8603);
nand U14533 (N_14533,N_5042,N_5177);
xor U14534 (N_14534,N_9956,N_9659);
and U14535 (N_14535,N_7846,N_6699);
nand U14536 (N_14536,N_9071,N_6277);
nor U14537 (N_14537,N_9194,N_8420);
nor U14538 (N_14538,N_5499,N_9582);
nor U14539 (N_14539,N_9623,N_9080);
and U14540 (N_14540,N_9005,N_9020);
and U14541 (N_14541,N_8386,N_5253);
and U14542 (N_14542,N_6718,N_9672);
or U14543 (N_14543,N_8977,N_6168);
xnor U14544 (N_14544,N_7366,N_7510);
nor U14545 (N_14545,N_9864,N_9954);
and U14546 (N_14546,N_6828,N_8584);
xnor U14547 (N_14547,N_7761,N_9232);
nand U14548 (N_14548,N_6956,N_5870);
and U14549 (N_14549,N_5819,N_8180);
or U14550 (N_14550,N_6710,N_6041);
xnor U14551 (N_14551,N_6472,N_8137);
nand U14552 (N_14552,N_7137,N_8924);
and U14553 (N_14553,N_9857,N_8195);
nor U14554 (N_14554,N_6559,N_5198);
xnor U14555 (N_14555,N_6692,N_8673);
and U14556 (N_14556,N_5440,N_6037);
xnor U14557 (N_14557,N_6266,N_5336);
nand U14558 (N_14558,N_7887,N_7799);
nor U14559 (N_14559,N_7189,N_6404);
or U14560 (N_14560,N_7539,N_9142);
nor U14561 (N_14561,N_5715,N_7014);
or U14562 (N_14562,N_9378,N_7595);
or U14563 (N_14563,N_9721,N_6215);
xor U14564 (N_14564,N_8856,N_9350);
xnor U14565 (N_14565,N_6429,N_7082);
xor U14566 (N_14566,N_6641,N_5495);
and U14567 (N_14567,N_9805,N_7071);
xnor U14568 (N_14568,N_7830,N_5329);
and U14569 (N_14569,N_8521,N_8970);
or U14570 (N_14570,N_9323,N_8686);
xor U14571 (N_14571,N_5420,N_9436);
nor U14572 (N_14572,N_6676,N_9447);
and U14573 (N_14573,N_5565,N_7726);
xnor U14574 (N_14574,N_9058,N_6355);
or U14575 (N_14575,N_7937,N_6023);
nor U14576 (N_14576,N_8026,N_8030);
nand U14577 (N_14577,N_7000,N_8425);
and U14578 (N_14578,N_9029,N_8409);
nand U14579 (N_14579,N_7876,N_5435);
or U14580 (N_14580,N_6661,N_9708);
and U14581 (N_14581,N_5475,N_9451);
xnor U14582 (N_14582,N_7007,N_9820);
nor U14583 (N_14583,N_8445,N_5135);
and U14584 (N_14584,N_9735,N_7749);
xor U14585 (N_14585,N_8216,N_5274);
and U14586 (N_14586,N_8221,N_5454);
xnor U14587 (N_14587,N_9459,N_7231);
nor U14588 (N_14588,N_6151,N_9877);
nand U14589 (N_14589,N_5261,N_5772);
nand U14590 (N_14590,N_8696,N_7737);
or U14591 (N_14591,N_5165,N_8894);
and U14592 (N_14592,N_9649,N_7858);
or U14593 (N_14593,N_8546,N_5085);
and U14594 (N_14594,N_7572,N_9784);
and U14595 (N_14595,N_6396,N_5821);
nor U14596 (N_14596,N_5240,N_7726);
xnor U14597 (N_14597,N_5518,N_7078);
or U14598 (N_14598,N_6576,N_8180);
xnor U14599 (N_14599,N_5797,N_9051);
and U14600 (N_14600,N_5832,N_9906);
xnor U14601 (N_14601,N_9493,N_6945);
xnor U14602 (N_14602,N_8563,N_7971);
nor U14603 (N_14603,N_9432,N_7763);
nand U14604 (N_14604,N_9596,N_7036);
xnor U14605 (N_14605,N_7824,N_6247);
or U14606 (N_14606,N_7575,N_6494);
xor U14607 (N_14607,N_8659,N_8610);
nor U14608 (N_14608,N_6071,N_6729);
nor U14609 (N_14609,N_5980,N_7067);
xor U14610 (N_14610,N_8398,N_6489);
xnor U14611 (N_14611,N_7127,N_8263);
or U14612 (N_14612,N_8537,N_7883);
nand U14613 (N_14613,N_8810,N_6045);
or U14614 (N_14614,N_5290,N_5628);
or U14615 (N_14615,N_5820,N_6190);
nor U14616 (N_14616,N_8743,N_5910);
and U14617 (N_14617,N_9320,N_5905);
xnor U14618 (N_14618,N_6470,N_8936);
and U14619 (N_14619,N_5761,N_5716);
nor U14620 (N_14620,N_9239,N_7791);
xnor U14621 (N_14621,N_9653,N_9645);
nand U14622 (N_14622,N_6073,N_7068);
xnor U14623 (N_14623,N_5770,N_8268);
nor U14624 (N_14624,N_5531,N_6436);
nor U14625 (N_14625,N_7274,N_9839);
nor U14626 (N_14626,N_7618,N_8431);
nand U14627 (N_14627,N_7593,N_8570);
or U14628 (N_14628,N_7803,N_8487);
nor U14629 (N_14629,N_5306,N_5234);
and U14630 (N_14630,N_7048,N_7464);
or U14631 (N_14631,N_5051,N_5215);
xnor U14632 (N_14632,N_7296,N_7131);
nor U14633 (N_14633,N_6969,N_9526);
xor U14634 (N_14634,N_7833,N_9980);
nand U14635 (N_14635,N_7177,N_5040);
nor U14636 (N_14636,N_8659,N_9114);
nand U14637 (N_14637,N_7108,N_7651);
xnor U14638 (N_14638,N_7803,N_6087);
nor U14639 (N_14639,N_5774,N_5407);
nand U14640 (N_14640,N_9586,N_7855);
nor U14641 (N_14641,N_5191,N_5001);
or U14642 (N_14642,N_6441,N_6442);
nor U14643 (N_14643,N_9636,N_6355);
nand U14644 (N_14644,N_5299,N_6389);
xor U14645 (N_14645,N_6569,N_6193);
xnor U14646 (N_14646,N_5705,N_5360);
nand U14647 (N_14647,N_8003,N_9445);
and U14648 (N_14648,N_9184,N_8665);
xnor U14649 (N_14649,N_7522,N_7325);
nand U14650 (N_14650,N_9529,N_7935);
and U14651 (N_14651,N_7005,N_6652);
xnor U14652 (N_14652,N_8735,N_6558);
or U14653 (N_14653,N_5195,N_6064);
nor U14654 (N_14654,N_8520,N_6734);
or U14655 (N_14655,N_6184,N_8926);
nand U14656 (N_14656,N_9133,N_5556);
or U14657 (N_14657,N_8088,N_9957);
nand U14658 (N_14658,N_9290,N_5530);
and U14659 (N_14659,N_7507,N_8583);
xnor U14660 (N_14660,N_9795,N_5982);
nor U14661 (N_14661,N_7481,N_8647);
or U14662 (N_14662,N_7012,N_8636);
and U14663 (N_14663,N_6984,N_9487);
nand U14664 (N_14664,N_6182,N_6363);
xor U14665 (N_14665,N_8780,N_5933);
nand U14666 (N_14666,N_9691,N_7183);
xnor U14667 (N_14667,N_6390,N_7479);
and U14668 (N_14668,N_7230,N_9486);
nand U14669 (N_14669,N_6813,N_6871);
or U14670 (N_14670,N_9074,N_9452);
nor U14671 (N_14671,N_5191,N_7146);
and U14672 (N_14672,N_9497,N_7754);
nand U14673 (N_14673,N_8840,N_9191);
nor U14674 (N_14674,N_6567,N_5216);
xor U14675 (N_14675,N_5578,N_5658);
nand U14676 (N_14676,N_5171,N_6087);
nand U14677 (N_14677,N_9898,N_5109);
nor U14678 (N_14678,N_9801,N_7391);
and U14679 (N_14679,N_5369,N_6678);
or U14680 (N_14680,N_9093,N_9774);
nand U14681 (N_14681,N_6927,N_9755);
xnor U14682 (N_14682,N_6564,N_5801);
nand U14683 (N_14683,N_8724,N_7188);
nand U14684 (N_14684,N_6457,N_9715);
and U14685 (N_14685,N_5661,N_6529);
nor U14686 (N_14686,N_7004,N_5142);
nor U14687 (N_14687,N_6553,N_9149);
or U14688 (N_14688,N_5532,N_9329);
xor U14689 (N_14689,N_8885,N_8119);
nand U14690 (N_14690,N_8208,N_9839);
nor U14691 (N_14691,N_6268,N_8002);
nor U14692 (N_14692,N_9248,N_5463);
and U14693 (N_14693,N_9153,N_8103);
xor U14694 (N_14694,N_6721,N_6970);
xor U14695 (N_14695,N_8967,N_8332);
or U14696 (N_14696,N_6388,N_5397);
xor U14697 (N_14697,N_9102,N_7839);
nor U14698 (N_14698,N_7905,N_8904);
or U14699 (N_14699,N_9784,N_8038);
nand U14700 (N_14700,N_9496,N_8581);
or U14701 (N_14701,N_7834,N_5248);
and U14702 (N_14702,N_9847,N_9386);
nor U14703 (N_14703,N_6770,N_6506);
xnor U14704 (N_14704,N_7619,N_9147);
xnor U14705 (N_14705,N_7404,N_6924);
xnor U14706 (N_14706,N_5822,N_7801);
nand U14707 (N_14707,N_8847,N_9656);
xor U14708 (N_14708,N_6587,N_5018);
nand U14709 (N_14709,N_8922,N_5780);
xor U14710 (N_14710,N_9713,N_8073);
and U14711 (N_14711,N_9457,N_8116);
xor U14712 (N_14712,N_9384,N_9595);
xnor U14713 (N_14713,N_8963,N_5712);
nand U14714 (N_14714,N_5403,N_9465);
xnor U14715 (N_14715,N_5239,N_7217);
xnor U14716 (N_14716,N_8679,N_8515);
and U14717 (N_14717,N_5435,N_7179);
nand U14718 (N_14718,N_7497,N_8196);
and U14719 (N_14719,N_8969,N_9911);
and U14720 (N_14720,N_8554,N_7208);
and U14721 (N_14721,N_8894,N_8627);
and U14722 (N_14722,N_6641,N_5926);
xnor U14723 (N_14723,N_9117,N_9761);
nand U14724 (N_14724,N_5127,N_7550);
nand U14725 (N_14725,N_7053,N_8063);
and U14726 (N_14726,N_5170,N_6056);
xnor U14727 (N_14727,N_5215,N_8273);
nand U14728 (N_14728,N_7806,N_6450);
xor U14729 (N_14729,N_5006,N_9483);
nand U14730 (N_14730,N_6358,N_5812);
or U14731 (N_14731,N_7387,N_8077);
nor U14732 (N_14732,N_8099,N_6861);
or U14733 (N_14733,N_8536,N_9701);
or U14734 (N_14734,N_5949,N_5809);
and U14735 (N_14735,N_6758,N_9909);
xor U14736 (N_14736,N_9624,N_9782);
and U14737 (N_14737,N_7934,N_8751);
nand U14738 (N_14738,N_5822,N_8789);
nor U14739 (N_14739,N_8937,N_9777);
nor U14740 (N_14740,N_9920,N_7948);
or U14741 (N_14741,N_6171,N_7895);
xnor U14742 (N_14742,N_6739,N_6815);
xnor U14743 (N_14743,N_6862,N_8318);
or U14744 (N_14744,N_8076,N_9549);
nor U14745 (N_14745,N_9131,N_5159);
nand U14746 (N_14746,N_7458,N_8891);
and U14747 (N_14747,N_5635,N_5793);
nand U14748 (N_14748,N_7976,N_7435);
nand U14749 (N_14749,N_7598,N_7267);
and U14750 (N_14750,N_5315,N_8973);
and U14751 (N_14751,N_8687,N_6886);
xor U14752 (N_14752,N_7137,N_7557);
nor U14753 (N_14753,N_9610,N_7219);
nand U14754 (N_14754,N_6032,N_5596);
nand U14755 (N_14755,N_5401,N_7965);
or U14756 (N_14756,N_6091,N_8744);
nand U14757 (N_14757,N_6813,N_7026);
and U14758 (N_14758,N_8292,N_6156);
and U14759 (N_14759,N_6083,N_9755);
or U14760 (N_14760,N_7509,N_5229);
or U14761 (N_14761,N_9080,N_8216);
or U14762 (N_14762,N_7325,N_9908);
xnor U14763 (N_14763,N_5440,N_8306);
nand U14764 (N_14764,N_5769,N_7179);
nand U14765 (N_14765,N_5314,N_8064);
nand U14766 (N_14766,N_9801,N_5856);
nor U14767 (N_14767,N_8134,N_9460);
or U14768 (N_14768,N_7279,N_9353);
xor U14769 (N_14769,N_6450,N_7458);
nor U14770 (N_14770,N_6176,N_5821);
and U14771 (N_14771,N_8031,N_7368);
and U14772 (N_14772,N_7284,N_8530);
xor U14773 (N_14773,N_7930,N_6575);
nor U14774 (N_14774,N_9530,N_9608);
or U14775 (N_14775,N_9938,N_9802);
and U14776 (N_14776,N_9377,N_6229);
xnor U14777 (N_14777,N_9030,N_9450);
or U14778 (N_14778,N_9127,N_7299);
xnor U14779 (N_14779,N_7720,N_8239);
or U14780 (N_14780,N_6665,N_8697);
and U14781 (N_14781,N_9972,N_9785);
or U14782 (N_14782,N_6030,N_8093);
nand U14783 (N_14783,N_6747,N_7783);
and U14784 (N_14784,N_6135,N_8758);
xor U14785 (N_14785,N_8690,N_9779);
and U14786 (N_14786,N_6995,N_9686);
nand U14787 (N_14787,N_7716,N_6712);
xnor U14788 (N_14788,N_6387,N_6033);
and U14789 (N_14789,N_7512,N_6188);
or U14790 (N_14790,N_6783,N_8543);
and U14791 (N_14791,N_8984,N_6013);
nand U14792 (N_14792,N_7016,N_7704);
and U14793 (N_14793,N_9066,N_8134);
and U14794 (N_14794,N_7687,N_5346);
or U14795 (N_14795,N_8254,N_8473);
nand U14796 (N_14796,N_5865,N_7663);
and U14797 (N_14797,N_6432,N_7797);
nand U14798 (N_14798,N_9673,N_8291);
or U14799 (N_14799,N_8225,N_6855);
nand U14800 (N_14800,N_8512,N_5635);
and U14801 (N_14801,N_9129,N_9801);
or U14802 (N_14802,N_5218,N_6549);
xnor U14803 (N_14803,N_5472,N_8386);
or U14804 (N_14804,N_9602,N_7593);
or U14805 (N_14805,N_6015,N_8120);
or U14806 (N_14806,N_9482,N_7320);
or U14807 (N_14807,N_7299,N_8168);
and U14808 (N_14808,N_9851,N_6730);
nor U14809 (N_14809,N_5214,N_6437);
xor U14810 (N_14810,N_9284,N_8423);
xnor U14811 (N_14811,N_7934,N_7506);
or U14812 (N_14812,N_5315,N_7682);
nor U14813 (N_14813,N_6794,N_7329);
and U14814 (N_14814,N_7638,N_7756);
and U14815 (N_14815,N_5319,N_8321);
xor U14816 (N_14816,N_6334,N_9309);
xnor U14817 (N_14817,N_5848,N_9510);
nand U14818 (N_14818,N_9523,N_9414);
nor U14819 (N_14819,N_6931,N_6709);
xor U14820 (N_14820,N_8772,N_9880);
or U14821 (N_14821,N_6805,N_6137);
and U14822 (N_14822,N_9364,N_9191);
or U14823 (N_14823,N_5986,N_7569);
nor U14824 (N_14824,N_6756,N_6757);
and U14825 (N_14825,N_8421,N_9892);
nor U14826 (N_14826,N_6296,N_8613);
xnor U14827 (N_14827,N_8302,N_8275);
or U14828 (N_14828,N_8252,N_7729);
xor U14829 (N_14829,N_9747,N_6215);
and U14830 (N_14830,N_9390,N_9797);
xor U14831 (N_14831,N_5950,N_5905);
nor U14832 (N_14832,N_6265,N_5018);
nand U14833 (N_14833,N_6057,N_9772);
and U14834 (N_14834,N_9853,N_7054);
or U14835 (N_14835,N_7140,N_6654);
xnor U14836 (N_14836,N_9388,N_7616);
and U14837 (N_14837,N_9109,N_8294);
nand U14838 (N_14838,N_7902,N_6048);
nand U14839 (N_14839,N_5645,N_9277);
or U14840 (N_14840,N_6512,N_6857);
or U14841 (N_14841,N_7447,N_9465);
or U14842 (N_14842,N_6450,N_6955);
or U14843 (N_14843,N_8724,N_7401);
nand U14844 (N_14844,N_9863,N_5764);
or U14845 (N_14845,N_6203,N_8992);
nor U14846 (N_14846,N_6980,N_6337);
xor U14847 (N_14847,N_6185,N_6889);
nand U14848 (N_14848,N_8411,N_9685);
and U14849 (N_14849,N_8168,N_9343);
and U14850 (N_14850,N_8688,N_5071);
xor U14851 (N_14851,N_6014,N_5776);
nand U14852 (N_14852,N_6638,N_6276);
and U14853 (N_14853,N_9018,N_8354);
and U14854 (N_14854,N_7497,N_9953);
xnor U14855 (N_14855,N_5174,N_7016);
nor U14856 (N_14856,N_6846,N_6816);
nor U14857 (N_14857,N_6394,N_9292);
nand U14858 (N_14858,N_6806,N_7293);
xor U14859 (N_14859,N_9081,N_7068);
nor U14860 (N_14860,N_9023,N_6068);
xnor U14861 (N_14861,N_8707,N_7665);
nand U14862 (N_14862,N_5471,N_8896);
and U14863 (N_14863,N_6318,N_6855);
xor U14864 (N_14864,N_9913,N_8000);
nand U14865 (N_14865,N_5534,N_9196);
or U14866 (N_14866,N_9060,N_9072);
xor U14867 (N_14867,N_9691,N_5993);
xor U14868 (N_14868,N_7000,N_8085);
nor U14869 (N_14869,N_6613,N_6360);
nor U14870 (N_14870,N_7327,N_5896);
nor U14871 (N_14871,N_9112,N_5199);
or U14872 (N_14872,N_9155,N_8565);
or U14873 (N_14873,N_7151,N_5014);
or U14874 (N_14874,N_6853,N_7863);
xnor U14875 (N_14875,N_5784,N_7093);
nor U14876 (N_14876,N_7770,N_5146);
and U14877 (N_14877,N_8969,N_5472);
nor U14878 (N_14878,N_6338,N_9250);
or U14879 (N_14879,N_9671,N_9339);
xor U14880 (N_14880,N_5459,N_8692);
and U14881 (N_14881,N_9237,N_5701);
and U14882 (N_14882,N_8767,N_9511);
nor U14883 (N_14883,N_6841,N_5841);
nand U14884 (N_14884,N_7230,N_7767);
nand U14885 (N_14885,N_5601,N_7405);
nor U14886 (N_14886,N_9029,N_9559);
nor U14887 (N_14887,N_8660,N_7638);
and U14888 (N_14888,N_7906,N_7039);
or U14889 (N_14889,N_5040,N_5299);
nor U14890 (N_14890,N_9479,N_6021);
nand U14891 (N_14891,N_5996,N_7867);
xnor U14892 (N_14892,N_7132,N_8376);
nor U14893 (N_14893,N_6964,N_9246);
nand U14894 (N_14894,N_7753,N_8451);
xnor U14895 (N_14895,N_8245,N_6991);
or U14896 (N_14896,N_5798,N_9796);
and U14897 (N_14897,N_5826,N_8230);
nor U14898 (N_14898,N_5786,N_8098);
xnor U14899 (N_14899,N_9819,N_8020);
nor U14900 (N_14900,N_9507,N_9700);
nor U14901 (N_14901,N_9033,N_5126);
xnor U14902 (N_14902,N_7660,N_7562);
or U14903 (N_14903,N_9681,N_8495);
nand U14904 (N_14904,N_6940,N_6319);
xnor U14905 (N_14905,N_9817,N_9710);
xor U14906 (N_14906,N_8423,N_8916);
nor U14907 (N_14907,N_7114,N_8787);
xnor U14908 (N_14908,N_6028,N_7117);
xnor U14909 (N_14909,N_9899,N_8363);
nand U14910 (N_14910,N_5177,N_9376);
nor U14911 (N_14911,N_7975,N_7423);
xnor U14912 (N_14912,N_5997,N_5668);
nor U14913 (N_14913,N_5174,N_8772);
or U14914 (N_14914,N_6811,N_9038);
or U14915 (N_14915,N_6386,N_5479);
and U14916 (N_14916,N_6770,N_7642);
nand U14917 (N_14917,N_7457,N_6905);
nor U14918 (N_14918,N_6567,N_9040);
xor U14919 (N_14919,N_5752,N_5652);
xnor U14920 (N_14920,N_5589,N_7870);
xnor U14921 (N_14921,N_6873,N_9318);
and U14922 (N_14922,N_9182,N_5261);
or U14923 (N_14923,N_5345,N_5580);
nand U14924 (N_14924,N_9592,N_6540);
nor U14925 (N_14925,N_5991,N_5420);
nor U14926 (N_14926,N_5532,N_6195);
xor U14927 (N_14927,N_6898,N_5180);
or U14928 (N_14928,N_9184,N_6715);
and U14929 (N_14929,N_8171,N_8025);
or U14930 (N_14930,N_5682,N_9562);
xnor U14931 (N_14931,N_8531,N_8849);
nor U14932 (N_14932,N_7790,N_7406);
nor U14933 (N_14933,N_7090,N_7645);
xnor U14934 (N_14934,N_5805,N_9843);
nand U14935 (N_14935,N_8079,N_8959);
or U14936 (N_14936,N_6741,N_5190);
nand U14937 (N_14937,N_9359,N_5031);
or U14938 (N_14938,N_6270,N_5206);
nand U14939 (N_14939,N_5076,N_6971);
nand U14940 (N_14940,N_6369,N_8130);
nand U14941 (N_14941,N_5896,N_5582);
xor U14942 (N_14942,N_9494,N_8507);
nand U14943 (N_14943,N_6048,N_9915);
nor U14944 (N_14944,N_7804,N_9440);
or U14945 (N_14945,N_5729,N_6340);
nor U14946 (N_14946,N_7203,N_8585);
xnor U14947 (N_14947,N_5646,N_9205);
xnor U14948 (N_14948,N_9473,N_8212);
xor U14949 (N_14949,N_8781,N_8344);
and U14950 (N_14950,N_9808,N_9343);
xnor U14951 (N_14951,N_8100,N_5925);
xnor U14952 (N_14952,N_9775,N_6062);
nor U14953 (N_14953,N_5956,N_7558);
nor U14954 (N_14954,N_9303,N_7413);
and U14955 (N_14955,N_5125,N_6499);
or U14956 (N_14956,N_8656,N_7010);
or U14957 (N_14957,N_9336,N_6316);
nand U14958 (N_14958,N_8554,N_9406);
nor U14959 (N_14959,N_6883,N_6132);
and U14960 (N_14960,N_9182,N_8793);
nor U14961 (N_14961,N_6027,N_6202);
nor U14962 (N_14962,N_5892,N_8371);
nand U14963 (N_14963,N_7698,N_5773);
nand U14964 (N_14964,N_6761,N_9649);
nand U14965 (N_14965,N_8293,N_9869);
xnor U14966 (N_14966,N_7727,N_7528);
or U14967 (N_14967,N_9786,N_6010);
nor U14968 (N_14968,N_5320,N_9306);
nor U14969 (N_14969,N_8780,N_8293);
nand U14970 (N_14970,N_9499,N_5875);
or U14971 (N_14971,N_9845,N_6406);
and U14972 (N_14972,N_7862,N_6946);
and U14973 (N_14973,N_6053,N_8914);
nor U14974 (N_14974,N_6675,N_5862);
and U14975 (N_14975,N_8817,N_9383);
xor U14976 (N_14976,N_9153,N_6687);
nand U14977 (N_14977,N_8770,N_7354);
and U14978 (N_14978,N_7437,N_7241);
nand U14979 (N_14979,N_8799,N_5910);
nand U14980 (N_14980,N_6983,N_7488);
or U14981 (N_14981,N_7365,N_8904);
xor U14982 (N_14982,N_8423,N_5147);
or U14983 (N_14983,N_7200,N_8786);
or U14984 (N_14984,N_8594,N_5388);
xor U14985 (N_14985,N_6483,N_6966);
or U14986 (N_14986,N_7520,N_5399);
or U14987 (N_14987,N_6996,N_6896);
nand U14988 (N_14988,N_7207,N_8235);
nand U14989 (N_14989,N_5969,N_9770);
or U14990 (N_14990,N_6944,N_5898);
xor U14991 (N_14991,N_7992,N_7923);
and U14992 (N_14992,N_8728,N_5211);
or U14993 (N_14993,N_6746,N_8280);
and U14994 (N_14994,N_8580,N_5205);
and U14995 (N_14995,N_5434,N_6217);
xnor U14996 (N_14996,N_8869,N_8233);
xor U14997 (N_14997,N_9766,N_9895);
or U14998 (N_14998,N_5108,N_5213);
nand U14999 (N_14999,N_9677,N_7714);
xor U15000 (N_15000,N_12964,N_13511);
or U15001 (N_15001,N_12383,N_13795);
and U15002 (N_15002,N_12929,N_14949);
nand U15003 (N_15003,N_14703,N_10955);
nand U15004 (N_15004,N_11685,N_10590);
nor U15005 (N_15005,N_14893,N_13285);
nand U15006 (N_15006,N_11225,N_12327);
xnor U15007 (N_15007,N_11532,N_11339);
xor U15008 (N_15008,N_13225,N_11233);
nand U15009 (N_15009,N_11141,N_10142);
xnor U15010 (N_15010,N_14952,N_10589);
or U15011 (N_15011,N_10722,N_11013);
or U15012 (N_15012,N_14255,N_12716);
nand U15013 (N_15013,N_12572,N_11594);
nand U15014 (N_15014,N_14785,N_10726);
or U15015 (N_15015,N_14782,N_12022);
and U15016 (N_15016,N_12786,N_14103);
nand U15017 (N_15017,N_11147,N_11336);
and U15018 (N_15018,N_10634,N_12349);
nor U15019 (N_15019,N_12185,N_14627);
and U15020 (N_15020,N_11278,N_13145);
nand U15021 (N_15021,N_13377,N_12799);
nor U15022 (N_15022,N_13973,N_14095);
xor U15023 (N_15023,N_13555,N_12027);
or U15024 (N_15024,N_10040,N_14573);
nand U15025 (N_15025,N_12497,N_12151);
nor U15026 (N_15026,N_10700,N_14894);
nor U15027 (N_15027,N_14825,N_13359);
xor U15028 (N_15028,N_14840,N_10222);
nor U15029 (N_15029,N_11898,N_13294);
nand U15030 (N_15030,N_10158,N_13545);
nand U15031 (N_15031,N_13263,N_11374);
or U15032 (N_15032,N_12251,N_11519);
xnor U15033 (N_15033,N_11097,N_13358);
xnor U15034 (N_15034,N_14432,N_11796);
and U15035 (N_15035,N_14836,N_14137);
xor U15036 (N_15036,N_14768,N_13443);
xnor U15037 (N_15037,N_10267,N_14352);
xnor U15038 (N_15038,N_11211,N_12605);
nand U15039 (N_15039,N_12390,N_10563);
xnor U15040 (N_15040,N_10831,N_14364);
nand U15041 (N_15041,N_11879,N_12548);
and U15042 (N_15042,N_12517,N_10095);
and U15043 (N_15043,N_14972,N_10471);
nor U15044 (N_15044,N_10845,N_10062);
nand U15045 (N_15045,N_11188,N_14168);
nand U15046 (N_15046,N_14610,N_10058);
nor U15047 (N_15047,N_10778,N_12459);
nor U15048 (N_15048,N_10692,N_11775);
nor U15049 (N_15049,N_13402,N_14899);
xor U15050 (N_15050,N_10024,N_13475);
or U15051 (N_15051,N_13078,N_10398);
or U15052 (N_15052,N_11073,N_11379);
nand U15053 (N_15053,N_10376,N_14908);
and U15054 (N_15054,N_14913,N_10909);
and U15055 (N_15055,N_11417,N_11235);
and U15056 (N_15056,N_10309,N_14463);
xnor U15057 (N_15057,N_13192,N_14822);
or U15058 (N_15058,N_10496,N_12375);
and U15059 (N_15059,N_14687,N_12587);
or U15060 (N_15060,N_10349,N_10195);
and U15061 (N_15061,N_10363,N_11162);
nor U15062 (N_15062,N_12313,N_11032);
and U15063 (N_15063,N_11588,N_13603);
nor U15064 (N_15064,N_13637,N_11101);
or U15065 (N_15065,N_13512,N_13076);
or U15066 (N_15066,N_10628,N_14329);
nand U15067 (N_15067,N_11944,N_10560);
xnor U15068 (N_15068,N_13298,N_13862);
xnor U15069 (N_15069,N_11824,N_11790);
nand U15070 (N_15070,N_12692,N_14163);
and U15071 (N_15071,N_10210,N_10649);
nor U15072 (N_15072,N_14957,N_12109);
nor U15073 (N_15073,N_14494,N_14931);
or U15074 (N_15074,N_11029,N_14268);
nand U15075 (N_15075,N_13820,N_14224);
nand U15076 (N_15076,N_12616,N_11507);
nor U15077 (N_15077,N_10096,N_14421);
or U15078 (N_15078,N_11381,N_14151);
nand U15079 (N_15079,N_11177,N_11576);
or U15080 (N_15080,N_14533,N_12366);
nor U15081 (N_15081,N_12886,N_14123);
xnor U15082 (N_15082,N_11783,N_13749);
nor U15083 (N_15083,N_14764,N_10678);
and U15084 (N_15084,N_13827,N_14150);
and U15085 (N_15085,N_11117,N_13431);
xor U15086 (N_15086,N_14727,N_14511);
and U15087 (N_15087,N_14404,N_10979);
xor U15088 (N_15088,N_14057,N_12300);
xor U15089 (N_15089,N_12393,N_10602);
and U15090 (N_15090,N_14692,N_10872);
xor U15091 (N_15091,N_13237,N_10161);
nand U15092 (N_15092,N_11825,N_14688);
xor U15093 (N_15093,N_10346,N_12636);
or U15094 (N_15094,N_12555,N_14049);
nand U15095 (N_15095,N_14482,N_10295);
or U15096 (N_15096,N_10554,N_11150);
or U15097 (N_15097,N_10420,N_11546);
nor U15098 (N_15098,N_11355,N_10412);
or U15099 (N_15099,N_13928,N_12681);
or U15100 (N_15100,N_13244,N_10596);
nand U15101 (N_15101,N_13420,N_14125);
nor U15102 (N_15102,N_14261,N_12642);
nand U15103 (N_15103,N_14447,N_13978);
nor U15104 (N_15104,N_13178,N_10547);
or U15105 (N_15105,N_14603,N_10520);
and U15106 (N_15106,N_14721,N_12610);
nand U15107 (N_15107,N_11208,N_11660);
or U15108 (N_15108,N_13049,N_13905);
nand U15109 (N_15109,N_10663,N_12210);
nand U15110 (N_15110,N_12701,N_13945);
and U15111 (N_15111,N_12117,N_13976);
and U15112 (N_15112,N_11031,N_14347);
or U15113 (N_15113,N_13961,N_13654);
and U15114 (N_15114,N_13213,N_13997);
nand U15115 (N_15115,N_13360,N_12891);
nand U15116 (N_15116,N_10952,N_10307);
xnor U15117 (N_15117,N_11108,N_14531);
nand U15118 (N_15118,N_11292,N_13700);
xor U15119 (N_15119,N_11595,N_11988);
xor U15120 (N_15120,N_14718,N_12316);
nand U15121 (N_15121,N_14536,N_14177);
xor U15122 (N_15122,N_11301,N_10773);
and U15123 (N_15123,N_12672,N_14522);
or U15124 (N_15124,N_13843,N_14632);
or U15125 (N_15125,N_11544,N_14301);
or U15126 (N_15126,N_14269,N_13129);
or U15127 (N_15127,N_14328,N_14334);
xnor U15128 (N_15128,N_14325,N_10552);
nor U15129 (N_15129,N_11493,N_14789);
nor U15130 (N_15130,N_12032,N_10861);
and U15131 (N_15131,N_14932,N_10584);
and U15132 (N_15132,N_10390,N_12887);
and U15133 (N_15133,N_10459,N_14921);
nor U15134 (N_15134,N_13874,N_12706);
or U15135 (N_15135,N_13342,N_10898);
xor U15136 (N_15136,N_12595,N_12078);
xnor U15137 (N_15137,N_12246,N_14165);
xnor U15138 (N_15138,N_10667,N_14503);
or U15139 (N_15139,N_14986,N_12689);
and U15140 (N_15140,N_11137,N_11267);
and U15141 (N_15141,N_13745,N_14655);
xor U15142 (N_15142,N_13607,N_11993);
xnor U15143 (N_15143,N_12319,N_13430);
nor U15144 (N_15144,N_12332,N_13794);
nand U15145 (N_15145,N_10237,N_11492);
xnor U15146 (N_15146,N_11288,N_12391);
or U15147 (N_15147,N_12979,N_11724);
nor U15148 (N_15148,N_12485,N_10915);
and U15149 (N_15149,N_12728,N_12167);
xor U15150 (N_15150,N_11348,N_14405);
nand U15151 (N_15151,N_10467,N_11470);
nor U15152 (N_15152,N_13268,N_14420);
nor U15153 (N_15153,N_13733,N_12395);
and U15154 (N_15154,N_12470,N_10859);
nor U15155 (N_15155,N_12667,N_14951);
or U15156 (N_15156,N_10483,N_14378);
nand U15157 (N_15157,N_11817,N_12164);
or U15158 (N_15158,N_12045,N_14176);
and U15159 (N_15159,N_13209,N_11322);
and U15160 (N_15160,N_11464,N_13707);
nand U15161 (N_15161,N_11501,N_10929);
xnor U15162 (N_15162,N_14792,N_14833);
or U15163 (N_15163,N_11787,N_12488);
xnor U15164 (N_15164,N_10739,N_13343);
and U15165 (N_15165,N_13458,N_12248);
or U15166 (N_15166,N_14476,N_14348);
nand U15167 (N_15167,N_14698,N_10291);
and U15168 (N_15168,N_10418,N_13015);
xor U15169 (N_15169,N_14526,N_10652);
nand U15170 (N_15170,N_13481,N_14067);
xnor U15171 (N_15171,N_12193,N_11036);
or U15172 (N_15172,N_13524,N_10636);
nand U15173 (N_15173,N_12344,N_12204);
nand U15174 (N_15174,N_14973,N_11627);
nor U15175 (N_15175,N_12064,N_14766);
nand U15176 (N_15176,N_14315,N_12108);
and U15177 (N_15177,N_11516,N_10710);
or U15178 (N_15178,N_14413,N_14635);
and U15179 (N_15179,N_10101,N_11420);
xor U15180 (N_15180,N_11894,N_11066);
or U15181 (N_15181,N_12206,N_13572);
or U15182 (N_15182,N_12918,N_12369);
xnor U15183 (N_15183,N_13964,N_13946);
nor U15184 (N_15184,N_10292,N_14280);
nand U15185 (N_15185,N_13867,N_14449);
xor U15186 (N_15186,N_12169,N_11466);
xnor U15187 (N_15187,N_11549,N_12745);
or U15188 (N_15188,N_11372,N_11949);
nor U15189 (N_15189,N_11525,N_10847);
or U15190 (N_15190,N_11762,N_13471);
nor U15191 (N_15191,N_10993,N_12453);
nand U15192 (N_15192,N_12850,N_13855);
xnor U15193 (N_15193,N_10816,N_14445);
and U15194 (N_15194,N_11473,N_12593);
nand U15195 (N_15195,N_13943,N_12474);
nor U15196 (N_15196,N_11881,N_11020);
xnor U15197 (N_15197,N_14898,N_14461);
xnor U15198 (N_15198,N_11643,N_11294);
xor U15199 (N_15199,N_10597,N_14978);
or U15200 (N_15200,N_10016,N_11967);
nand U15201 (N_15201,N_13418,N_14853);
and U15202 (N_15202,N_12469,N_10744);
or U15203 (N_15203,N_13930,N_11377);
nor U15204 (N_15204,N_13882,N_11165);
nand U15205 (N_15205,N_13799,N_13510);
or U15206 (N_15206,N_12287,N_10469);
xnor U15207 (N_15207,N_11465,N_11127);
or U15208 (N_15208,N_12569,N_14650);
xor U15209 (N_15209,N_14529,N_12427);
and U15210 (N_15210,N_13688,N_12877);
and U15211 (N_15211,N_10765,N_11264);
nor U15212 (N_15212,N_12450,N_11043);
and U15213 (N_15213,N_12530,N_10511);
or U15214 (N_15214,N_11435,N_10767);
and U15215 (N_15215,N_11099,N_10379);
nor U15216 (N_15216,N_13550,N_14528);
xor U15217 (N_15217,N_14771,N_14388);
or U15218 (N_15218,N_13156,N_12471);
or U15219 (N_15219,N_14143,N_12789);
nor U15220 (N_15220,N_12201,N_10896);
nand U15221 (N_15221,N_13438,N_13502);
xnor U15222 (N_15222,N_11149,N_10509);
nand U15223 (N_15223,N_14945,N_13123);
nand U15224 (N_15224,N_14832,N_14873);
xnor U15225 (N_15225,N_11412,N_12126);
and U15226 (N_15226,N_12992,N_11620);
and U15227 (N_15227,N_11648,N_12950);
xnor U15228 (N_15228,N_13281,N_12059);
or U15229 (N_15229,N_13066,N_13303);
xor U15230 (N_15230,N_13551,N_11940);
xnor U15231 (N_15231,N_10913,N_14954);
and U15232 (N_15232,N_12568,N_10997);
nor U15233 (N_15233,N_10685,N_12999);
nand U15234 (N_15234,N_14953,N_13547);
nand U15235 (N_15235,N_14346,N_10711);
nor U15236 (N_15236,N_11171,N_12919);
nand U15237 (N_15237,N_13762,N_13063);
nand U15238 (N_15238,N_14600,N_10974);
and U15239 (N_15239,N_13863,N_11917);
nor U15240 (N_15240,N_10729,N_10169);
xor U15241 (N_15241,N_12675,N_14097);
xor U15242 (N_15242,N_10912,N_12409);
xor U15243 (N_15243,N_14201,N_11258);
and U15244 (N_15244,N_10903,N_13927);
nor U15245 (N_15245,N_14468,N_14229);
and U15246 (N_15246,N_14085,N_13200);
nand U15247 (N_15247,N_12826,N_11652);
xor U15248 (N_15248,N_14985,N_10426);
nand U15249 (N_15249,N_13683,N_14896);
or U15250 (N_15250,N_11059,N_12447);
nand U15251 (N_15251,N_10757,N_11703);
nor U15252 (N_15252,N_12356,N_10894);
nor U15253 (N_15253,N_11132,N_12034);
nor U15254 (N_15254,N_14772,N_13922);
and U15255 (N_15255,N_11715,N_12107);
and U15256 (N_15256,N_14530,N_10423);
xor U15257 (N_15257,N_13877,N_14379);
nor U15258 (N_15258,N_13424,N_13333);
and U15259 (N_15259,N_10437,N_12718);
nor U15260 (N_15260,N_14171,N_13125);
and U15261 (N_15261,N_14015,N_11863);
nand U15262 (N_15262,N_13439,N_11340);
nor U15263 (N_15263,N_11399,N_12779);
or U15264 (N_15264,N_14885,N_13426);
and U15265 (N_15265,N_13891,N_10198);
nor U15266 (N_15266,N_11402,N_10247);
or U15267 (N_15267,N_12732,N_12969);
nand U15268 (N_15268,N_10111,N_10824);
or U15269 (N_15269,N_10555,N_10294);
xnor U15270 (N_15270,N_10190,N_13613);
xnor U15271 (N_15271,N_11971,N_11959);
nor U15272 (N_15272,N_13926,N_10372);
nand U15273 (N_15273,N_11913,N_14206);
or U15274 (N_15274,N_11027,N_12884);
xnor U15275 (N_15275,N_12773,N_11864);
xor U15276 (N_15276,N_12602,N_11404);
xor U15277 (N_15277,N_11996,N_11587);
and U15278 (N_15278,N_11873,N_13786);
xnor U15279 (N_15279,N_11789,N_13159);
nand U15280 (N_15280,N_10300,N_13714);
nand U15281 (N_15281,N_10830,N_10867);
nand U15282 (N_15282,N_14733,N_13632);
or U15283 (N_15283,N_10605,N_14197);
or U15284 (N_15284,N_13215,N_14009);
nor U15285 (N_15285,N_12446,N_11236);
nand U15286 (N_15286,N_13509,N_11401);
xor U15287 (N_15287,N_11976,N_10234);
xnor U15288 (N_15288,N_10638,N_12230);
and U15289 (N_15289,N_11803,N_12532);
nor U15290 (N_15290,N_12721,N_11287);
or U15291 (N_15291,N_12696,N_13187);
xor U15292 (N_15292,N_13672,N_12995);
xor U15293 (N_15293,N_11369,N_10644);
nand U15294 (N_15294,N_14656,N_10537);
nor U15295 (N_15295,N_14955,N_10617);
nand U15296 (N_15296,N_10647,N_11343);
or U15297 (N_15297,N_11909,N_10592);
nor U15298 (N_15298,N_11063,N_10808);
nor U15299 (N_15299,N_13923,N_11540);
and U15300 (N_15300,N_12484,N_10821);
xor U15301 (N_15301,N_13616,N_14377);
nand U15302 (N_15302,N_13288,N_12996);
nor U15303 (N_15303,N_11529,N_12054);
nand U15304 (N_15304,N_14363,N_14619);
nand U15305 (N_15305,N_13484,N_10461);
xor U15306 (N_15306,N_10166,N_12277);
nor U15307 (N_15307,N_10524,N_12067);
nand U15308 (N_15308,N_11094,N_13530);
xor U15309 (N_15309,N_14738,N_11897);
nor U15310 (N_15310,N_14475,N_11812);
or U15311 (N_15311,N_11541,N_11609);
nand U15312 (N_15312,N_13691,N_12902);
or U15313 (N_15313,N_13436,N_10255);
nor U15314 (N_15314,N_14866,N_12284);
nor U15315 (N_15315,N_13025,N_14800);
xnor U15316 (N_15316,N_12521,N_12702);
and U15317 (N_15317,N_13167,N_12425);
or U15318 (N_15318,N_13692,N_12410);
nand U15319 (N_15319,N_11397,N_13705);
or U15320 (N_15320,N_11745,N_13950);
and U15321 (N_15321,N_11347,N_14689);
or U15322 (N_15322,N_10801,N_13531);
nor U15323 (N_15323,N_12498,N_11052);
or U15324 (N_15324,N_11628,N_11337);
xnor U15325 (N_15325,N_14070,N_14002);
xnor U15326 (N_15326,N_11157,N_11123);
nor U15327 (N_15327,N_11770,N_13105);
nor U15328 (N_15328,N_12601,N_13222);
and U15329 (N_15329,N_14695,N_13223);
nand U15330 (N_15330,N_10521,N_14033);
nor U15331 (N_15331,N_11054,N_12763);
nor U15332 (N_15332,N_13212,N_12741);
and U15333 (N_15333,N_12867,N_12239);
and U15334 (N_15334,N_10193,N_12691);
nand U15335 (N_15335,N_14310,N_13642);
nand U15336 (N_15336,N_12567,N_10180);
nor U15337 (N_15337,N_12796,N_14725);
or U15338 (N_15338,N_13035,N_14005);
and U15339 (N_15339,N_11567,N_14044);
nor U15340 (N_15340,N_11077,N_12559);
nor U15341 (N_15341,N_14118,N_12035);
nor U15342 (N_15342,N_11018,N_13061);
and U15343 (N_15343,N_12767,N_14936);
nand U15344 (N_15344,N_11647,N_10782);
nand U15345 (N_15345,N_10699,N_13506);
or U15346 (N_15346,N_11736,N_14107);
nor U15347 (N_15347,N_13102,N_14906);
nor U15348 (N_15348,N_13047,N_13816);
and U15349 (N_15349,N_11217,N_11952);
nor U15350 (N_15350,N_10144,N_12677);
nand U15351 (N_15351,N_12268,N_11344);
xnor U15352 (N_15352,N_10562,N_12250);
nand U15353 (N_15353,N_10174,N_10028);
xnor U15354 (N_15354,N_10740,N_11624);
and U15355 (N_15355,N_12822,N_14161);
or U15356 (N_15356,N_12942,N_13437);
xor U15357 (N_15357,N_13190,N_11923);
nor U15358 (N_15358,N_13069,N_10764);
nor U15359 (N_15359,N_11445,N_13925);
nand U15360 (N_15360,N_11633,N_11279);
or U15361 (N_15361,N_13042,N_14036);
or U15362 (N_15362,N_13638,N_11857);
nand U15363 (N_15363,N_14467,N_12270);
and U15364 (N_15364,N_14916,N_13114);
nor U15365 (N_15365,N_12180,N_10301);
or U15366 (N_15366,N_12703,N_12159);
and U15367 (N_15367,N_13340,N_11120);
xor U15368 (N_15368,N_14676,N_12573);
or U15369 (N_15369,N_12331,N_13407);
or U15370 (N_15370,N_11689,N_10984);
or U15371 (N_15371,N_10341,N_11542);
and U15372 (N_15372,N_14540,N_10728);
nand U15373 (N_15373,N_14061,N_13173);
nand U15374 (N_15374,N_11290,N_10573);
nand U15375 (N_15375,N_13847,N_11433);
nand U15376 (N_15376,N_10356,N_12845);
nand U15377 (N_15377,N_11273,N_12576);
xnor U15378 (N_15378,N_10789,N_10565);
nor U15379 (N_15379,N_11823,N_11552);
or U15380 (N_15380,N_11742,N_11152);
xnor U15381 (N_15381,N_11721,N_12232);
nand U15382 (N_15382,N_10591,N_10574);
nand U15383 (N_15383,N_12906,N_13236);
xnor U15384 (N_15384,N_11191,N_12993);
and U15385 (N_15385,N_12515,N_11760);
or U15386 (N_15386,N_14779,N_10855);
xor U15387 (N_15387,N_12611,N_11874);
or U15388 (N_15388,N_12039,N_13028);
and U15389 (N_15389,N_11170,N_11781);
or U15390 (N_15390,N_12192,N_13957);
xnor U15391 (N_15391,N_10790,N_11616);
or U15392 (N_15392,N_10799,N_12042);
xor U15393 (N_15393,N_12790,N_10038);
and U15394 (N_15394,N_13844,N_11030);
xor U15395 (N_15395,N_10250,N_13544);
nor U15396 (N_15396,N_13203,N_14863);
and U15397 (N_15397,N_10570,N_12468);
xnor U15398 (N_15398,N_14281,N_10064);
and U15399 (N_15399,N_11670,N_10559);
and U15400 (N_15400,N_11534,N_13627);
or U15401 (N_15401,N_14356,N_11843);
and U15402 (N_15402,N_11256,N_11835);
xnor U15403 (N_15403,N_11777,N_10545);
or U15404 (N_15404,N_10397,N_11320);
or U15405 (N_15405,N_12781,N_14966);
or U15406 (N_15406,N_10084,N_12968);
and U15407 (N_15407,N_11304,N_12758);
and U15408 (N_15408,N_13180,N_12129);
or U15409 (N_15409,N_13866,N_10077);
xnor U15410 (N_15410,N_14994,N_10967);
or U15411 (N_15411,N_12755,N_12553);
nand U15412 (N_15412,N_14905,N_14767);
nand U15413 (N_15413,N_10529,N_10454);
nand U15414 (N_15414,N_10625,N_13994);
and U15415 (N_15415,N_11237,N_12833);
or U15416 (N_15416,N_12063,N_13489);
xor U15417 (N_15417,N_10449,N_12868);
xor U15418 (N_15418,N_12203,N_10175);
and U15419 (N_15419,N_12374,N_12695);
nor U15420 (N_15420,N_14382,N_14109);
nand U15421 (N_15421,N_14265,N_12462);
nor U15422 (N_15422,N_10494,N_13919);
xnor U15423 (N_15423,N_14093,N_13831);
and U15424 (N_15424,N_11793,N_10853);
or U15425 (N_15425,N_14060,N_14045);
nand U15426 (N_15426,N_11346,N_13146);
or U15427 (N_15427,N_14317,N_12678);
nor U15428 (N_15428,N_10873,N_10057);
or U15429 (N_15429,N_14104,N_14842);
and U15430 (N_15430,N_10433,N_13787);
and U15431 (N_15431,N_14625,N_14336);
and U15432 (N_15432,N_11382,N_11637);
xnor U15433 (N_15433,N_13837,N_12843);
xor U15434 (N_15434,N_12306,N_14648);
nand U15435 (N_15435,N_11116,N_14318);
and U15436 (N_15436,N_11164,N_14572);
xnor U15437 (N_15437,N_10092,N_13767);
nor U15438 (N_15438,N_10150,N_10138);
nand U15439 (N_15439,N_12719,N_12861);
xnor U15440 (N_15440,N_10274,N_13110);
and U15441 (N_15441,N_12258,N_14474);
nor U15442 (N_15442,N_12988,N_14158);
and U15443 (N_15443,N_14874,N_14839);
nand U15444 (N_15444,N_13269,N_14642);
or U15445 (N_15445,N_10709,N_11155);
xnor U15446 (N_15446,N_12442,N_13202);
nor U15447 (N_15447,N_11615,N_13953);
xor U15448 (N_15448,N_14728,N_11593);
nand U15449 (N_15449,N_11297,N_14845);
xnor U15450 (N_15450,N_12388,N_13088);
nand U15451 (N_15451,N_12176,N_14222);
and U15452 (N_15452,N_14277,N_13456);
nand U15453 (N_15453,N_13365,N_10128);
and U15454 (N_15454,N_11598,N_11386);
xor U15455 (N_15455,N_10503,N_12265);
nand U15456 (N_15456,N_10844,N_14236);
nor U15457 (N_15457,N_13163,N_10962);
nor U15458 (N_15458,N_11428,N_14576);
xnor U15459 (N_15459,N_11318,N_14391);
xnor U15460 (N_15460,N_10104,N_14081);
xor U15461 (N_15461,N_11836,N_14758);
nor U15462 (N_15462,N_13322,N_13954);
nor U15463 (N_15463,N_14697,N_14759);
or U15464 (N_15464,N_12604,N_13419);
xor U15465 (N_15465,N_14791,N_12307);
xnor U15466 (N_15466,N_13783,N_10681);
xnor U15467 (N_15467,N_13195,N_11130);
or U15468 (N_15468,N_13518,N_14244);
xor U15469 (N_15469,N_11193,N_12663);
xor U15470 (N_15470,N_12544,N_10080);
xnor U15471 (N_15471,N_12749,N_12564);
or U15472 (N_15472,N_11599,N_14918);
xor U15473 (N_15473,N_14867,N_13247);
xnor U15474 (N_15474,N_11449,N_10048);
xor U15475 (N_15475,N_14562,N_12435);
nand U15476 (N_15476,N_11497,N_13046);
nand U15477 (N_15477,N_12247,N_10856);
xnor U15478 (N_15478,N_12197,N_10436);
and U15479 (N_15479,N_10173,N_11509);
and U15480 (N_15480,N_11642,N_12314);
and U15481 (N_15481,N_11143,N_13653);
and U15482 (N_15482,N_10023,N_11167);
and U15483 (N_15483,N_10034,N_10703);
and U15484 (N_15484,N_11220,N_10120);
xor U15485 (N_15485,N_11938,N_14958);
nand U15486 (N_15486,N_12679,N_10164);
xor U15487 (N_15487,N_11559,N_10876);
and U15488 (N_15488,N_14581,N_13310);
nand U15489 (N_15489,N_13680,N_11392);
xor U15490 (N_15490,N_13472,N_13258);
or U15491 (N_15491,N_14122,N_12873);
nor U15492 (N_15492,N_11808,N_14233);
nand U15493 (N_15493,N_14570,N_14911);
xnor U15494 (N_15494,N_14948,N_14929);
and U15495 (N_15495,N_10310,N_13806);
xnor U15496 (N_15496,N_11677,N_14284);
xor U15497 (N_15497,N_14322,N_10067);
xnor U15498 (N_15498,N_12637,N_12328);
nand U15499 (N_15499,N_11126,N_12693);
or U15500 (N_15500,N_12088,N_11302);
or U15501 (N_15501,N_10124,N_12399);
or U15502 (N_15502,N_10707,N_10424);
nor U15503 (N_15503,N_12002,N_12281);
or U15504 (N_15504,N_10388,N_13324);
nor U15505 (N_15505,N_14205,N_13622);
or U15506 (N_15506,N_14232,N_10994);
nor U15507 (N_15507,N_10833,N_13341);
and U15508 (N_15508,N_10313,N_11042);
nor U15509 (N_15509,N_11496,N_10694);
xor U15510 (N_15510,N_13559,N_12785);
and U15511 (N_15511,N_10725,N_12953);
nor U15512 (N_15512,N_12512,N_14199);
and U15513 (N_15513,N_14547,N_11315);
and U15514 (N_15514,N_14128,N_13211);
and U15515 (N_15515,N_10796,N_14018);
and U15516 (N_15516,N_11345,N_11792);
nor U15517 (N_15517,N_12997,N_14838);
and U15518 (N_15518,N_11075,N_14466);
nor U15519 (N_15519,N_14561,N_13573);
nor U15520 (N_15520,N_11558,N_12155);
and U15521 (N_15521,N_10624,N_14302);
xor U15522 (N_15522,N_13248,N_11946);
nand U15523 (N_15523,N_13620,N_13461);
or U15524 (N_15524,N_12924,N_14471);
or U15525 (N_15525,N_12536,N_14719);
or U15526 (N_15526,N_13574,N_11600);
or U15527 (N_15527,N_14793,N_12960);
and U15528 (N_15528,N_13589,N_11842);
or U15529 (N_15529,N_14820,N_14069);
nand U15530 (N_15530,N_14492,N_10956);
nor U15531 (N_15531,N_11753,N_10156);
xor U15532 (N_15532,N_13083,N_10007);
nand U15533 (N_15533,N_13729,N_10304);
nand U15534 (N_15534,N_12365,N_10192);
nand U15535 (N_15535,N_13353,N_11138);
nor U15536 (N_15536,N_13395,N_12980);
xnor U15537 (N_15537,N_10795,N_14127);
and U15538 (N_15538,N_13916,N_13280);
xnor U15539 (N_15539,N_12050,N_14702);
and U15540 (N_15540,N_12492,N_10339);
or U15541 (N_15541,N_11640,N_13869);
and U15542 (N_15542,N_12226,N_10297);
xnor U15543 (N_15543,N_10293,N_14657);
nand U15544 (N_15544,N_13164,N_14464);
nor U15545 (N_15545,N_10528,N_14801);
or U15546 (N_15546,N_13630,N_11102);
or U15547 (N_15547,N_14699,N_11907);
xnor U15548 (N_15548,N_14849,N_11231);
or U15549 (N_15549,N_11666,N_11727);
nand U15550 (N_15550,N_11696,N_14493);
nand U15551 (N_15551,N_12628,N_10618);
or U15552 (N_15552,N_14734,N_12614);
and U15553 (N_15553,N_11764,N_14664);
xnor U15554 (N_15554,N_12320,N_13271);
and U15555 (N_15555,N_11717,N_11527);
xor U15556 (N_15556,N_12674,N_10910);
or U15557 (N_15557,N_12046,N_13940);
xor U15558 (N_15558,N_14852,N_10041);
nor U15559 (N_15559,N_11081,N_13266);
or U15560 (N_15560,N_13805,N_12486);
or U15561 (N_15561,N_14508,N_14480);
xnor U15562 (N_15562,N_11611,N_14074);
or U15563 (N_15563,N_12212,N_13516);
xor U15564 (N_15564,N_10010,N_12998);
nor U15565 (N_15565,N_11895,N_13161);
nor U15566 (N_15566,N_10961,N_14257);
nand U15567 (N_15567,N_14937,N_14204);
xor U15568 (N_15568,N_14011,N_11688);
nor U15569 (N_15569,N_13910,N_13526);
or U15570 (N_15570,N_11456,N_13681);
nor U15571 (N_15571,N_13447,N_13775);
and U15572 (N_15572,N_11748,N_13763);
nor U15573 (N_15573,N_12487,N_13554);
nand U15574 (N_15574,N_11517,N_11644);
xor U15575 (N_15575,N_11104,N_12771);
xor U15576 (N_15576,N_13659,N_10836);
nor U15577 (N_15577,N_14035,N_11706);
nand U15578 (N_15578,N_11145,N_14102);
xor U15579 (N_15579,N_12848,N_14380);
and U15580 (N_15580,N_12858,N_14705);
or U15581 (N_15581,N_14510,N_12917);
xor U15582 (N_15582,N_13480,N_11479);
or U15583 (N_15583,N_14130,N_11869);
nand U15584 (N_15584,N_11209,N_14170);
or U15585 (N_15585,N_11769,N_10788);
xnor U15586 (N_15586,N_13245,N_13966);
and U15587 (N_15587,N_13425,N_12113);
xnor U15588 (N_15588,N_11367,N_11205);
xor U15589 (N_15589,N_10286,N_13153);
nor U15590 (N_15590,N_10608,N_13104);
nor U15591 (N_15591,N_13391,N_11385);
and U15592 (N_15592,N_11608,N_10977);
nand U15593 (N_15593,N_13583,N_12895);
nor U15594 (N_15594,N_11072,N_12188);
nor U15595 (N_15595,N_10514,N_10784);
or U15596 (N_15596,N_10172,N_14512);
and U15597 (N_15597,N_10407,N_12400);
and U15598 (N_15598,N_10908,N_10680);
nor U15599 (N_15599,N_14136,N_11914);
nor U15600 (N_15600,N_10553,N_14979);
nor U15601 (N_15601,N_10693,N_12903);
nand U15602 (N_15602,N_12121,N_10140);
xnor U15603 (N_15603,N_14495,N_12297);
xor U15604 (N_15604,N_14537,N_11071);
nand U15605 (N_15605,N_14569,N_13534);
and U15606 (N_15606,N_11396,N_12658);
nand U15607 (N_15607,N_13062,N_14630);
nand U15608 (N_15608,N_10899,N_13140);
nor U15609 (N_15609,N_10452,N_14487);
and U15610 (N_15610,N_12939,N_10862);
nand U15611 (N_15611,N_14544,N_12940);
nor U15612 (N_15612,N_10588,N_14477);
nand U15613 (N_15613,N_13290,N_14462);
nor U15614 (N_15614,N_14134,N_12419);
xnor U15615 (N_15615,N_13639,N_14580);
and U15616 (N_15616,N_11661,N_11484);
and U15617 (N_15617,N_11841,N_12191);
or U15618 (N_15618,N_10254,N_13537);
or U15619 (N_15619,N_11530,N_12264);
and U15620 (N_15620,N_11729,N_14663);
nand U15621 (N_15621,N_12336,N_12526);
and U15622 (N_15622,N_11092,N_11065);
nand U15623 (N_15623,N_14964,N_11405);
and U15624 (N_15624,N_14938,N_11524);
xnor U15625 (N_15625,N_14194,N_14740);
nand U15626 (N_15626,N_12049,N_13821);
xnor U15627 (N_15627,N_14659,N_14409);
nor U15628 (N_15628,N_13181,N_13406);
nand U15629 (N_15629,N_13802,N_11806);
and U15630 (N_15630,N_11011,N_11747);
and U15631 (N_15631,N_14735,N_12591);
xor U15632 (N_15632,N_10047,N_11555);
xnor U15633 (N_15633,N_13948,N_14567);
and U15634 (N_15634,N_12099,N_10924);
and U15635 (N_15635,N_14187,N_11270);
and U15636 (N_15636,N_10999,N_13890);
nor U15637 (N_15637,N_11105,N_11118);
nand U15638 (N_15638,N_14080,N_11639);
nor U15639 (N_15639,N_12102,N_13538);
nand U15640 (N_15640,N_10276,N_14998);
nor U15641 (N_15641,N_14427,N_12136);
or U15642 (N_15642,N_12676,N_10475);
nand U15643 (N_15643,N_10935,N_11296);
and U15644 (N_15644,N_12735,N_10296);
nand U15645 (N_15645,N_13713,N_14647);
or U15646 (N_15646,N_12178,N_13598);
and U15647 (N_15647,N_12303,N_10655);
nor U15648 (N_15648,N_10148,N_11480);
nand U15649 (N_15649,N_12086,N_10432);
nand U15650 (N_15650,N_10727,N_12851);
or U15651 (N_15651,N_11780,N_12819);
xnor U15652 (N_15652,N_12343,N_14691);
or U15653 (N_15653,N_10708,N_11954);
and U15654 (N_15654,N_11195,N_14757);
xnor U15655 (N_15655,N_10619,N_11674);
nor U15656 (N_15656,N_13201,N_12842);
nor U15657 (N_15657,N_12132,N_10330);
xnor U15658 (N_15658,N_11908,N_10259);
xnor U15659 (N_15659,N_12590,N_12948);
or U15660 (N_15660,N_14995,N_10311);
and U15661 (N_15661,N_11033,N_11389);
nand U15662 (N_15662,N_12900,N_14773);
or U15663 (N_15663,N_13336,N_14411);
nand U15664 (N_15664,N_13120,N_12956);
or U15665 (N_15665,N_14860,N_14987);
nand U15666 (N_15666,N_11210,N_12172);
and U15667 (N_15667,N_12480,N_11431);
or U15668 (N_15668,N_14827,N_12615);
xor U15669 (N_15669,N_12632,N_13982);
xnor U15670 (N_15670,N_10575,N_10137);
or U15671 (N_15671,N_10980,N_10567);
nand U15672 (N_15672,N_10448,N_13094);
nor U15673 (N_15673,N_14794,N_12872);
nand U15674 (N_15674,N_11927,N_12158);
and U15675 (N_15675,N_10539,N_11046);
nand U15676 (N_15676,N_12346,N_14403);
nor U15677 (N_15677,N_12537,N_13975);
xnor U15678 (N_15678,N_14871,N_12715);
xor U15679 (N_15679,N_11390,N_14670);
xor U15680 (N_15680,N_12808,N_11463);
and U15681 (N_15681,N_13362,N_12489);
and U15682 (N_15682,N_11740,N_11360);
or U15683 (N_15683,N_11249,N_13698);
and U15684 (N_15684,N_12584,N_12147);
and U15685 (N_15685,N_12818,N_13467);
xor U15686 (N_15686,N_11667,N_13117);
and U15687 (N_15687,N_12778,N_10127);
and U15688 (N_15688,N_11617,N_14841);
or U15689 (N_15689,N_11618,N_14888);
nand U15690 (N_15690,N_11266,N_12751);
xnor U15691 (N_15691,N_14338,N_10202);
xnor U15692 (N_15692,N_14271,N_10087);
xnor U15693 (N_15693,N_14928,N_14481);
and U15694 (N_15694,N_13283,N_11603);
and U15695 (N_15695,N_14030,N_13776);
xnor U15696 (N_15696,N_13924,N_12205);
nand U15697 (N_15697,N_13468,N_14374);
nand U15698 (N_15698,N_14981,N_14398);
nor U15699 (N_15699,N_10525,N_10004);
xor U15700 (N_15700,N_10018,N_12661);
and U15701 (N_15701,N_14654,N_11111);
nor U15702 (N_15702,N_12134,N_12464);
and U15703 (N_15703,N_12361,N_13540);
or U15704 (N_15704,N_14278,N_12062);
xnor U15705 (N_15705,N_13541,N_13373);
and U15706 (N_15706,N_12019,N_10181);
nand U15707 (N_15707,N_14690,N_10081);
nand U15708 (N_15708,N_11862,N_12820);
nand U15709 (N_15709,N_13103,N_10800);
nand U15710 (N_15710,N_10561,N_12358);
nor U15711 (N_15711,N_11978,N_12018);
and U15712 (N_15712,N_10809,N_12334);
and U15713 (N_15713,N_14882,N_12617);
and U15714 (N_15714,N_12016,N_13896);
nor U15715 (N_15715,N_10919,N_11083);
xnor U15716 (N_15716,N_11912,N_14554);
xnor U15717 (N_15717,N_13500,N_13548);
nor U15718 (N_15718,N_10743,N_10717);
nand U15719 (N_15719,N_11774,N_14636);
or U15720 (N_15720,N_13249,N_14519);
nand U15721 (N_15721,N_12142,N_10535);
or U15722 (N_15722,N_13356,N_12913);
and U15723 (N_15723,N_10675,N_12523);
and U15724 (N_15724,N_10052,N_14961);
xnor U15725 (N_15725,N_13457,N_13641);
nand U15726 (N_15726,N_12404,N_13759);
nand U15727 (N_15727,N_12766,N_14276);
nor U15728 (N_15728,N_10938,N_14549);
and U15729 (N_15729,N_10218,N_10612);
nand U15730 (N_15730,N_10118,N_11638);
and U15731 (N_15731,N_12345,N_13053);
nand U15732 (N_15732,N_11441,N_12413);
and U15733 (N_15733,N_11941,N_11429);
or U15734 (N_15734,N_10585,N_10671);
xor U15735 (N_15735,N_14881,N_11983);
nor U15736 (N_15736,N_14947,N_13326);
nor U15737 (N_15737,N_12550,N_11543);
nor U15738 (N_15738,N_14666,N_10277);
xnor U15739 (N_15739,N_14333,N_13319);
xnor U15740 (N_15740,N_12357,N_11438);
nand U15741 (N_15741,N_13284,N_13040);
nor U15742 (N_15742,N_11458,N_12240);
and U15743 (N_15743,N_13807,N_14020);
or U15744 (N_15744,N_13760,N_13179);
and U15745 (N_15745,N_13351,N_10507);
or U15746 (N_15746,N_11001,N_13274);
and U15747 (N_15747,N_10664,N_10695);
and U15748 (N_15748,N_10840,N_11649);
xor U15749 (N_15749,N_12516,N_11457);
and U15750 (N_15750,N_13119,N_14884);
nor U15751 (N_15751,N_13375,N_11248);
nor U15752 (N_15752,N_10954,N_13564);
and U15753 (N_15753,N_12869,N_10630);
or U15754 (N_15754,N_11686,N_13999);
xor U15755 (N_15755,N_14350,N_12295);
and U15756 (N_15756,N_14564,N_13278);
and U15757 (N_15757,N_11733,N_12140);
nor U15758 (N_15758,N_12020,N_12920);
and U15759 (N_15759,N_14708,N_14907);
nand U15760 (N_15760,N_14672,N_11169);
nor U15761 (N_15761,N_14668,N_12299);
nand U15762 (N_15762,N_14681,N_11476);
and U15763 (N_15763,N_14146,N_13984);
and U15764 (N_15764,N_10223,N_13977);
nand U15765 (N_15765,N_10691,N_11921);
or U15766 (N_15766,N_11380,N_12682);
nor U15767 (N_15767,N_13969,N_14217);
or U15768 (N_15768,N_12966,N_11012);
nor U15769 (N_15769,N_14798,N_10813);
nand U15770 (N_15770,N_13856,N_13724);
nor U15771 (N_15771,N_10907,N_11291);
nand U15772 (N_15772,N_10990,N_10761);
xnor U15773 (N_15773,N_14596,N_13731);
xor U15774 (N_15774,N_11477,N_14747);
xor U15775 (N_15775,N_14730,N_13399);
or U15776 (N_15776,N_13016,N_11260);
and U15777 (N_15777,N_10316,N_12430);
or U15778 (N_15778,N_14601,N_13711);
nand U15779 (N_15779,N_14514,N_14919);
nor U15780 (N_15780,N_11110,N_12283);
and U15781 (N_15781,N_14307,N_14816);
xor U15782 (N_15782,N_11212,N_11659);
nand U15783 (N_15783,N_14414,N_11395);
nor U15784 (N_15784,N_12925,N_12222);
or U15785 (N_15785,N_11482,N_10093);
or U15786 (N_15786,N_13568,N_13096);
and U15787 (N_15787,N_14072,N_10697);
nand U15788 (N_15788,N_10843,N_12742);
xnor U15789 (N_15789,N_13264,N_10822);
and U15790 (N_15790,N_11213,N_14289);
nand U15791 (N_15791,N_10457,N_10474);
nand U15792 (N_15792,N_12829,N_14682);
or U15793 (N_15793,N_10261,N_10425);
and U15794 (N_15794,N_11680,N_13220);
nand U15795 (N_15795,N_13815,N_12467);
xnor U15796 (N_15796,N_13836,N_13935);
or U15797 (N_15797,N_12244,N_14942);
or U15798 (N_15798,N_13095,N_12744);
xor U15799 (N_15799,N_10530,N_13979);
nand U15800 (N_15800,N_13851,N_10826);
or U15801 (N_15801,N_10290,N_13282);
or U15802 (N_15802,N_10783,N_12079);
or U15803 (N_15803,N_14628,N_10829);
nor U15804 (N_15804,N_11654,N_11454);
and U15805 (N_15805,N_11426,N_13171);
and U15806 (N_15806,N_11312,N_13682);
xor U15807 (N_15807,N_10232,N_11720);
xor U15808 (N_15808,N_13868,N_10620);
and U15809 (N_15809,N_10668,N_13817);
nand U15810 (N_15810,N_11310,N_11916);
or U15811 (N_15811,N_10838,N_11329);
xnor U15812 (N_15812,N_12641,N_10989);
and U15813 (N_15813,N_10531,N_14077);
nor U15814 (N_15814,N_13558,N_11303);
nor U15815 (N_15815,N_11265,N_10768);
and U15816 (N_15816,N_12618,N_11810);
nand U15817 (N_15817,N_10009,N_12262);
nor U15818 (N_15818,N_10019,N_14343);
xor U15819 (N_15819,N_13137,N_11766);
nor U15820 (N_15820,N_12511,N_10421);
nand U15821 (N_15821,N_14368,N_11815);
or U15822 (N_15822,N_12426,N_11704);
or U15823 (N_15823,N_14804,N_13350);
or U15824 (N_15824,N_13592,N_14260);
or U15825 (N_15825,N_10332,N_11121);
xor U15826 (N_15826,N_14927,N_12800);
or U15827 (N_15827,N_14351,N_11252);
or U15828 (N_15828,N_11788,N_13034);
nor U15829 (N_15829,N_14988,N_12394);
nor U15830 (N_15830,N_13014,N_13355);
and U15831 (N_15831,N_10405,N_10661);
or U15832 (N_15832,N_12128,N_14160);
or U15833 (N_15833,N_14683,N_13533);
or U15834 (N_15834,N_13686,N_13291);
nor U15835 (N_15835,N_13937,N_13838);
and U15836 (N_15836,N_10686,N_13903);
nor U15837 (N_15837,N_12124,N_13904);
and U15838 (N_15838,N_14591,N_12671);
and U15839 (N_15839,N_10216,N_13671);
and U15840 (N_15840,N_14751,N_10951);
and U15841 (N_15841,N_14525,N_10947);
and U15842 (N_15842,N_14453,N_14967);
and U15843 (N_15843,N_13386,N_12803);
nand U15844 (N_15844,N_10996,N_11816);
and U15845 (N_15845,N_12865,N_10888);
and U15846 (N_15846,N_10071,N_10749);
and U15847 (N_15847,N_12945,N_14605);
and U15848 (N_15848,N_11794,N_13658);
nand U15849 (N_15849,N_12153,N_11631);
or U15850 (N_15850,N_11306,N_10600);
xnor U15851 (N_15851,N_13077,N_14577);
and U15852 (N_15852,N_14408,N_11430);
and U15853 (N_15853,N_14117,N_14064);
nor U15854 (N_15854,N_11230,N_10226);
or U15855 (N_15855,N_10289,N_11321);
nand U15856 (N_15856,N_11577,N_14539);
nor U15857 (N_15857,N_12104,N_12673);
and U15858 (N_15858,N_10738,N_13774);
or U15859 (N_15859,N_13238,N_13728);
or U15860 (N_15860,N_12814,N_14148);
nand U15861 (N_15861,N_12087,N_12444);
nor U15862 (N_15862,N_13304,N_11166);
and U15863 (N_15863,N_10526,N_13496);
nor U15864 (N_15864,N_11883,N_13051);
and U15865 (N_15865,N_10315,N_11784);
nor U15866 (N_15866,N_13834,N_13677);
or U15867 (N_15867,N_10239,N_13007);
and U15868 (N_15868,N_10604,N_13858);
nand U15869 (N_15869,N_13477,N_11942);
nor U15870 (N_15870,N_14478,N_10603);
nor U15871 (N_15871,N_12729,N_13566);
nor U15872 (N_15872,N_12768,N_13273);
nor U15873 (N_15873,N_11695,N_12607);
nor U15874 (N_15874,N_14052,N_11103);
or U15875 (N_15875,N_10770,N_11447);
nor U15876 (N_15876,N_12839,N_13645);
xnor U15877 (N_15877,N_13824,N_12603);
nor U15878 (N_15878,N_11804,N_10005);
xor U15879 (N_15879,N_14710,N_14593);
and U15880 (N_15880,N_12805,N_12440);
xor U15881 (N_15881,N_14761,N_10564);
nand U15882 (N_15882,N_13260,N_11754);
or U15883 (N_15883,N_14909,N_10230);
nor U15884 (N_15884,N_10544,N_11716);
or U15885 (N_15885,N_14303,N_13678);
nand U15886 (N_15886,N_13751,N_14488);
or U15887 (N_15887,N_11767,N_12528);
or U15888 (N_15888,N_11289,N_12387);
xnor U15889 (N_15889,N_11752,N_11100);
nor U15890 (N_15890,N_13138,N_10443);
nor U15891 (N_15891,N_10143,N_13958);
xor U15892 (N_15892,N_14043,N_10026);
nor U15893 (N_15893,N_14939,N_14607);
and U15894 (N_15894,N_12077,N_11698);
or U15895 (N_15895,N_11682,N_10191);
xnor U15896 (N_15896,N_12223,N_12890);
nand U15897 (N_15897,N_13228,N_10519);
and U15898 (N_15898,N_12910,N_10260);
nand U15899 (N_15899,N_14644,N_11311);
nor U15900 (N_15900,N_13004,N_14360);
and U15901 (N_15901,N_11768,N_11274);
and U15902 (N_15902,N_11737,N_14202);
nor U15903 (N_15903,N_13981,N_12080);
nor U15904 (N_15904,N_13112,N_13990);
nand U15905 (N_15905,N_14039,N_11936);
or U15906 (N_15906,N_10627,N_13970);
nand U15907 (N_15907,N_10501,N_12631);
nand U15908 (N_15908,N_10429,N_14989);
and U15909 (N_15909,N_13813,N_12200);
xor U15910 (N_15910,N_11006,N_10932);
nand U15911 (N_15911,N_14256,N_14763);
or U15912 (N_15912,N_12912,N_14220);
nand U15913 (N_15913,N_14181,N_12011);
and U15914 (N_15914,N_10981,N_13543);
nor U15915 (N_15915,N_14588,N_10086);
and U15916 (N_15916,N_10430,N_12967);
nor U15917 (N_15917,N_14565,N_11450);
and U15918 (N_15918,N_10670,N_13828);
and U15919 (N_15919,N_10576,N_12139);
xor U15920 (N_15920,N_11929,N_11192);
xor U15921 (N_15921,N_13587,N_14667);
nand U15922 (N_15922,N_10037,N_10450);
and U15923 (N_15923,N_13750,N_12699);
nand U15924 (N_15924,N_14071,N_12263);
and U15925 (N_15925,N_13508,N_10074);
and U15926 (N_15926,N_11341,N_10455);
nand U15927 (N_15927,N_11148,N_10460);
nand U15928 (N_15928,N_11945,N_11090);
or U15929 (N_15929,N_12074,N_13239);
xnor U15930 (N_15930,N_11738,N_11522);
nor U15931 (N_15931,N_12285,N_12793);
nand U15932 (N_15932,N_10413,N_13801);
xnor U15933 (N_15933,N_12213,N_12520);
xor U15934 (N_15934,N_14386,N_13569);
nand U15935 (N_15935,N_14837,N_14606);
nor U15936 (N_15936,N_12652,N_14633);
or U15937 (N_15937,N_14436,N_14568);
nand U15938 (N_15938,N_14502,N_10123);
nor U15939 (N_15939,N_13348,N_13670);
and U15940 (N_15940,N_11699,N_10416);
xor U15941 (N_15941,N_14819,N_12580);
or U15942 (N_15942,N_14895,N_12043);
nor U15943 (N_15943,N_12448,N_13071);
xor U15944 (N_15944,N_12272,N_14566);
nand U15945 (N_15945,N_12775,N_13716);
nand U15946 (N_15946,N_10914,N_14019);
nand U15947 (N_15947,N_11511,N_14314);
nor U15948 (N_15948,N_10078,N_12686);
or U15949 (N_15949,N_11741,N_12522);
xnor U15950 (N_15950,N_14812,N_12482);
or U15951 (N_15951,N_11335,N_13084);
nand U15952 (N_15952,N_13757,N_14308);
xnor U15953 (N_15953,N_11047,N_13091);
and U15954 (N_15954,N_10365,N_13299);
nand U15955 (N_15955,N_11502,N_14634);
xor U15956 (N_15956,N_10747,N_10171);
nor U15957 (N_15957,N_13734,N_10248);
nor U15958 (N_15958,N_10470,N_12882);
or U15959 (N_15959,N_10392,N_10109);
and U15960 (N_15960,N_11676,N_11584);
xor U15961 (N_15961,N_13871,N_13722);
and U15962 (N_15962,N_13060,N_13210);
xor U15963 (N_15963,N_14267,N_12036);
or U15964 (N_15964,N_14341,N_10194);
or U15965 (N_15965,N_10066,N_10852);
xnor U15966 (N_15966,N_13738,N_10441);
or U15967 (N_15967,N_11154,N_11349);
xnor U15968 (N_15968,N_11761,N_12457);
or U15969 (N_15969,N_14431,N_12606);
nand U15970 (N_15970,N_10263,N_11151);
xor U15971 (N_15971,N_12111,N_13251);
and U15972 (N_15972,N_10964,N_11641);
and U15973 (N_15973,N_10760,N_14711);
xor U15974 (N_15974,N_12832,N_11363);
or U15975 (N_15975,N_14774,N_13732);
and U15976 (N_15976,N_10050,N_13106);
xnor U15977 (N_15977,N_10482,N_10165);
xor U15978 (N_15978,N_14159,N_14183);
xor U15979 (N_15979,N_13772,N_11325);
nor U15980 (N_15980,N_14465,N_13079);
nand U15981 (N_15981,N_11601,N_14920);
or U15982 (N_15982,N_13427,N_10170);
nand U15983 (N_15983,N_11370,N_12171);
xnor U15984 (N_15984,N_11613,N_13328);
nand U15985 (N_15985,N_11467,N_10854);
nor U15986 (N_15986,N_10285,N_14754);
nand U15987 (N_15987,N_11697,N_11338);
nor U15988 (N_15988,N_10622,N_10442);
nor U15989 (N_15989,N_11612,N_14991);
nand U15990 (N_15990,N_14615,N_14182);
nand U15991 (N_15991,N_14700,N_11896);
or U15992 (N_15992,N_13697,N_10763);
nor U15993 (N_15993,N_13704,N_10209);
or U15994 (N_15994,N_12417,N_12893);
xor U15995 (N_15995,N_14149,N_14614);
nor U15996 (N_15996,N_13452,N_10730);
nor U15997 (N_15997,N_10488,N_13032);
and U15998 (N_15998,N_14900,N_14479);
nand U15999 (N_15999,N_13073,N_13886);
nand U16000 (N_16000,N_10130,N_14621);
and U16001 (N_16001,N_12322,N_11560);
and U16002 (N_16002,N_14399,N_14821);
nor U16003 (N_16003,N_13148,N_13219);
xnor U16004 (N_16004,N_14319,N_12137);
nor U16005 (N_16005,N_10944,N_11427);
nor U16006 (N_16006,N_10724,N_12897);
nand U16007 (N_16007,N_12994,N_13379);
xnor U16008 (N_16008,N_13908,N_11868);
and U16009 (N_16009,N_12531,N_14456);
and U16010 (N_16010,N_14861,N_10581);
nand U16011 (N_16011,N_11453,N_13143);
and U16012 (N_16012,N_12382,N_11809);
nand U16013 (N_16013,N_14762,N_13715);
nor U16014 (N_16014,N_13445,N_12752);
xor U16015 (N_16015,N_14755,N_10721);
and U16016 (N_16016,N_10324,N_14891);
nor U16017 (N_16017,N_10329,N_13183);
and U16018 (N_16018,N_12234,N_11730);
nand U16019 (N_16019,N_12711,N_11356);
nand U16020 (N_16020,N_11219,N_14631);
nor U16021 (N_16021,N_13401,N_11713);
nand U16022 (N_16022,N_13441,N_13405);
and U16023 (N_16023,N_11472,N_12982);
and U16024 (N_16024,N_14598,N_11726);
or U16025 (N_16025,N_12748,N_13606);
xor U16026 (N_16026,N_10643,N_13773);
and U16027 (N_16027,N_14520,N_13694);
nand U16028 (N_16028,N_13501,N_14392);
nand U16029 (N_16029,N_10049,N_10920);
and U16030 (N_16030,N_12952,N_14062);
or U16031 (N_16031,N_12380,N_14883);
or U16032 (N_16032,N_12243,N_10476);
xnor U16033 (N_16033,N_12533,N_14661);
and U16034 (N_16034,N_12071,N_14320);
nor U16035 (N_16035,N_13830,N_10549);
or U16036 (N_16036,N_11773,N_12235);
nor U16037 (N_16037,N_11022,N_13412);
nor U16038 (N_16038,N_14976,N_12508);
and U16039 (N_16039,N_10792,N_11106);
nor U16040 (N_16040,N_10648,N_12985);
and U16041 (N_16041,N_10771,N_13364);
or U16042 (N_16042,N_13621,N_11979);
nand U16043 (N_16043,N_13859,N_14746);
and U16044 (N_16044,N_13989,N_14144);
and U16045 (N_16045,N_13124,N_10508);
nand U16046 (N_16046,N_13579,N_14752);
xnor U16047 (N_16047,N_11388,N_10672);
nor U16048 (N_16048,N_12150,N_10769);
and U16049 (N_16049,N_12278,N_10933);
xnor U16050 (N_16050,N_12451,N_13064);
nand U16051 (N_16051,N_11972,N_13906);
xnor U16052 (N_16052,N_13043,N_14749);
or U16053 (N_16053,N_10646,N_12739);
nand U16054 (N_16054,N_14450,N_11142);
and U16055 (N_16055,N_13019,N_11829);
xor U16056 (N_16056,N_14831,N_14297);
xnor U16057 (N_16057,N_14396,N_10184);
and U16058 (N_16058,N_11876,N_10152);
nand U16059 (N_16059,N_11610,N_10345);
or U16060 (N_16060,N_11692,N_13038);
and U16061 (N_16061,N_14426,N_14584);
or U16062 (N_16062,N_12625,N_10839);
and U16063 (N_16063,N_11425,N_14188);
and U16064 (N_16064,N_14083,N_12415);
xnor U16065 (N_16065,N_11771,N_14068);
xor U16066 (N_16066,N_14869,N_14221);
or U16067 (N_16067,N_12855,N_11621);
xnor U16068 (N_16068,N_13563,N_14162);
or U16069 (N_16069,N_10359,N_14864);
nor U16070 (N_16070,N_10734,N_10960);
or U16071 (N_16071,N_11280,N_13486);
or U16072 (N_16072,N_12725,N_14370);
xnor U16073 (N_16073,N_12040,N_13422);
xor U16074 (N_16074,N_10870,N_10404);
xor U16075 (N_16075,N_12666,N_10008);
and U16076 (N_16076,N_10523,N_14722);
or U16077 (N_16077,N_14678,N_10238);
or U16078 (N_16078,N_10848,N_13796);
xor U16079 (N_16079,N_11095,N_14418);
xor U16080 (N_16080,N_13968,N_13567);
xor U16081 (N_16081,N_11244,N_13879);
nor U16082 (N_16082,N_14589,N_12225);
nand U16083 (N_16083,N_10776,N_11570);
xor U16084 (N_16084,N_10614,N_14507);
nand U16085 (N_16085,N_11316,N_14324);
xor U16086 (N_16086,N_12065,N_13081);
or U16087 (N_16087,N_14407,N_10271);
or U16088 (N_16088,N_12983,N_10543);
and U16089 (N_16089,N_10399,N_10201);
or U16090 (N_16090,N_11391,N_14486);
xor U16091 (N_16091,N_11653,N_10106);
nor U16092 (N_16092,N_14583,N_13693);
and U16093 (N_16093,N_10033,N_11739);
xor U16094 (N_16094,N_13149,N_10682);
nand U16095 (N_16095,N_10107,N_14677);
or U16096 (N_16096,N_13352,N_12000);
or U16097 (N_16097,N_13381,N_14796);
xor U16098 (N_16098,N_13535,N_13597);
nand U16099 (N_16099,N_14879,N_11565);
nand U16100 (N_16100,N_10586,N_10212);
nor U16101 (N_16101,N_12707,N_11950);
xor U16102 (N_16102,N_12423,N_11051);
or U16103 (N_16103,N_11384,N_14359);
and U16104 (N_16104,N_11039,N_11866);
nor U16105 (N_16105,N_14034,N_12827);
xor U16106 (N_16106,N_14558,N_11185);
nand U16107 (N_16107,N_14933,N_14875);
nor U16108 (N_16108,N_12312,N_10003);
or U16109 (N_16109,N_10723,N_11705);
or U16110 (N_16110,N_13860,N_10378);
nand U16111 (N_16111,N_14311,N_13302);
and U16112 (N_16112,N_11911,N_11872);
and U16113 (N_16113,N_12935,N_12740);
xnor U16114 (N_16114,N_10930,N_13701);
nor U16115 (N_16115,N_10163,N_12236);
xor U16116 (N_16116,N_14028,N_14497);
nor U16117 (N_16117,N_13320,N_10484);
nand U16118 (N_16118,N_11495,N_11197);
xnor U16119 (N_16119,N_14604,N_12629);
nand U16120 (N_16120,N_10215,N_12310);
nor U16121 (N_16121,N_14496,N_14330);
or U16122 (N_16122,N_12600,N_13382);
xnor U16123 (N_16123,N_11554,N_11134);
and U16124 (N_16124,N_10518,N_14287);
nand U16125 (N_16125,N_12598,N_12863);
nor U16126 (N_16126,N_10417,N_10121);
and U16127 (N_16127,N_11364,N_11376);
nand U16128 (N_16128,N_13718,N_14675);
nor U16129 (N_16129,N_12411,N_12914);
nor U16130 (N_16130,N_14595,N_12282);
nor U16131 (N_16131,N_13657,N_13504);
nand U16132 (N_16132,N_11224,N_10902);
xor U16133 (N_16133,N_13565,N_11407);
nor U16134 (N_16134,N_11175,N_13933);
and U16135 (N_16135,N_14053,N_10931);
and U16136 (N_16136,N_11475,N_14169);
and U16137 (N_16137,N_11460,N_12228);
xnor U16138 (N_16138,N_13666,N_11393);
or U16139 (N_16139,N_12026,N_14805);
nor U16140 (N_16140,N_11067,N_14099);
and U16141 (N_16141,N_10492,N_13898);
xnor U16142 (N_16142,N_14131,N_13218);
nand U16143 (N_16143,N_10090,N_10035);
and U16144 (N_16144,N_11867,N_10477);
or U16145 (N_16145,N_10408,N_13497);
and U16146 (N_16146,N_14559,N_12438);
and U16147 (N_16147,N_10965,N_13041);
nand U16148 (N_16148,N_11571,N_10340);
nor U16149 (N_16149,N_14208,N_12029);
nor U16150 (N_16150,N_13020,N_13136);
and U16151 (N_16151,N_12094,N_11853);
or U16152 (N_16152,N_14982,N_10645);
or U16153 (N_16153,N_12259,N_14808);
nand U16154 (N_16154,N_12298,N_12597);
nor U16155 (N_16155,N_13434,N_11798);
xnor U16156 (N_16156,N_12504,N_10265);
nor U16157 (N_16157,N_13725,N_13577);
and U16158 (N_16158,N_14813,N_14098);
nor U16159 (N_16159,N_14546,N_13610);
or U16160 (N_16160,N_12770,N_14440);
nand U16161 (N_16161,N_10918,N_11424);
and U16162 (N_16162,N_12461,N_12329);
nor U16163 (N_16163,N_14215,N_12455);
nor U16164 (N_16164,N_11061,N_13099);
xor U16165 (N_16165,N_12127,N_12296);
and U16166 (N_16166,N_10139,N_11206);
and U16167 (N_16167,N_10595,N_13792);
nand U16168 (N_16168,N_10712,N_13523);
or U16169 (N_16169,N_10522,N_12743);
and U16170 (N_16170,N_13988,N_10462);
nand U16171 (N_16171,N_11658,N_10249);
nor U16172 (N_16172,N_14375,N_14997);
or U16173 (N_16173,N_10435,N_10396);
nand U16174 (N_16174,N_13082,N_10558);
nor U16175 (N_16175,N_10214,N_14084);
xnor U16176 (N_16176,N_12353,N_13667);
xor U16177 (N_16177,N_13934,N_11523);
xnor U16178 (N_16178,N_14291,N_12443);
nor U16179 (N_16179,N_11899,N_11683);
xnor U16180 (N_16180,N_10533,N_13221);
nand U16181 (N_16181,N_11634,N_11243);
and U16182 (N_16182,N_11547,N_12592);
nor U16183 (N_16183,N_11956,N_10168);
or U16184 (N_16184,N_11085,N_11515);
and U16185 (N_16185,N_13026,N_12305);
nor U16186 (N_16186,N_14299,N_11722);
or U16187 (N_16187,N_12688,N_11007);
nor U16188 (N_16188,N_11758,N_13170);
nor U16189 (N_16189,N_14780,N_13995);
or U16190 (N_16190,N_10091,N_13253);
and U16191 (N_16191,N_12582,N_10353);
xor U16192 (N_16192,N_12211,N_13494);
nand U16193 (N_16193,N_12651,N_12143);
or U16194 (N_16194,N_11814,N_10705);
xor U16195 (N_16195,N_12558,N_12105);
nor U16196 (N_16196,N_14517,N_11285);
and U16197 (N_16197,N_13470,N_11136);
nand U16198 (N_16198,N_13893,N_13086);
or U16199 (N_16199,N_12783,N_12866);
or U16200 (N_16200,N_12753,N_10837);
or U16201 (N_16201,N_14145,N_10061);
nor U16202 (N_16202,N_14505,N_13314);
or U16203 (N_16203,N_13250,N_10897);
nand U16204 (N_16204,N_11107,N_13897);
xnor U16205 (N_16205,N_10126,N_10688);
nand U16206 (N_16206,N_10299,N_10986);
nand U16207 (N_16207,N_14200,N_11202);
nor U16208 (N_16208,N_13735,N_10995);
xnor U16209 (N_16209,N_12166,N_13582);
and U16210 (N_16210,N_10401,N_13003);
nand U16211 (N_16211,N_10716,N_10270);
and U16212 (N_16212,N_11974,N_12539);
nand U16213 (N_16213,N_14575,N_13482);
or U16214 (N_16214,N_14295,N_10613);
and U16215 (N_16215,N_14094,N_13131);
and U16216 (N_16216,N_11062,N_14904);
nand U16217 (N_16217,N_11830,N_10568);
nor U16218 (N_16218,N_10042,N_12021);
or U16219 (N_16219,N_11284,N_13367);
nor U16220 (N_16220,N_14397,N_12012);
and U16221 (N_16221,N_12685,N_13649);
and U16222 (N_16222,N_13634,N_10021);
xor U16223 (N_16223,N_14003,N_10866);
xnor U16224 (N_16224,N_14935,N_10427);
nor U16225 (N_16225,N_10361,N_13012);
or U16226 (N_16226,N_12747,N_12546);
or U16227 (N_16227,N_14425,N_14385);
or U16228 (N_16228,N_10103,N_11901);
nor U16229 (N_16229,N_12946,N_10719);
or U16230 (N_16230,N_11440,N_13542);
nor U16231 (N_16231,N_13135,N_10516);
and U16232 (N_16232,N_11975,N_11003);
xor U16233 (N_16233,N_14189,N_12791);
or U16234 (N_16234,N_11746,N_12981);
or U16235 (N_16235,N_12005,N_13741);
xor U16236 (N_16236,N_13396,N_13329);
xor U16237 (N_16237,N_13960,N_11551);
or U16238 (N_16238,N_12535,N_10674);
and U16239 (N_16239,N_13665,N_12368);
and U16240 (N_16240,N_14856,N_11045);
nor U16241 (N_16241,N_14608,N_11779);
and U16242 (N_16242,N_14643,N_10434);
xnor U16243 (N_16243,N_10633,N_11553);
or U16244 (N_16244,N_13029,N_13243);
or U16245 (N_16245,N_11446,N_12289);
or U16246 (N_16246,N_14846,N_10781);
and U16247 (N_16247,N_14886,N_10053);
or U16248 (N_16248,N_11187,N_12609);
nand U16249 (N_16249,N_13044,N_10465);
xnor U16250 (N_16250,N_13991,N_10207);
xor U16251 (N_16251,N_12309,N_13633);
and U16252 (N_16252,N_10958,N_14959);
xnor U16253 (N_16253,N_12061,N_10885);
nand U16254 (N_16254,N_14415,N_11928);
nand U16255 (N_16255,N_14887,N_12549);
nor U16256 (N_16256,N_14716,N_13765);
xor U16257 (N_16257,N_13947,N_10953);
xor U16258 (N_16258,N_10060,N_13663);
nor U16259 (N_16259,N_14639,N_14858);
or U16260 (N_16260,N_13575,N_11023);
or U16261 (N_16261,N_13685,N_10926);
nor U16262 (N_16262,N_11579,N_13624);
nor U16263 (N_16263,N_10601,N_14611);
and U16264 (N_16264,N_13972,N_12904);
and U16265 (N_16265,N_10065,N_10335);
and U16266 (N_16266,N_13661,N_14219);
or U16267 (N_16267,N_11034,N_10972);
nand U16268 (N_16268,N_14665,N_11707);
and U16269 (N_16269,N_12254,N_13098);
nand U16270 (N_16270,N_10387,N_11700);
and U16271 (N_16271,N_10863,N_12003);
or U16272 (N_16272,N_11194,N_12503);
and U16273 (N_16273,N_13812,N_12901);
nand U16274 (N_16274,N_13588,N_14444);
nand U16275 (N_16275,N_10456,N_13307);
and U16276 (N_16276,N_14592,N_13782);
xor U16277 (N_16277,N_10527,N_14400);
or U16278 (N_16278,N_12575,N_10676);
xor U16279 (N_16279,N_13414,N_14880);
nand U16280 (N_16280,N_10438,N_14741);
xnor U16281 (N_16281,N_14047,N_14455);
nor U16282 (N_16282,N_11822,N_11383);
nor U16283 (N_16283,N_13527,N_12571);
and U16284 (N_16284,N_14059,N_10446);
or U16285 (N_16285,N_10354,N_10242);
and U16286 (N_16286,N_13027,N_10205);
xor U16287 (N_16287,N_12001,N_11275);
or U16288 (N_16288,N_10370,N_10110);
and U16289 (N_16289,N_10323,N_13743);
and U16290 (N_16290,N_12574,N_11556);
or U16291 (N_16291,N_11886,N_13507);
nor U16292 (N_16292,N_11904,N_13217);
nor U16293 (N_16293,N_11221,N_11906);
or U16294 (N_16294,N_13899,N_11669);
or U16295 (N_16295,N_12170,N_14114);
and U16296 (N_16296,N_14999,N_10141);
nand U16297 (N_16297,N_11261,N_13938);
or U16298 (N_16298,N_11295,N_12053);
nor U16299 (N_16299,N_14765,N_10011);
or U16300 (N_16300,N_10834,N_10656);
xor U16301 (N_16301,N_12970,N_14327);
or U16302 (N_16302,N_13067,N_10325);
and U16303 (N_16303,N_12965,N_13719);
or U16304 (N_16304,N_11690,N_10850);
xnor U16305 (N_16305,N_13885,N_12157);
nor U16306 (N_16306,N_13374,N_11905);
nand U16307 (N_16307,N_11889,N_14054);
xnor U16308 (N_16308,N_11079,N_13522);
xnor U16309 (N_16309,N_10225,N_11299);
nand U16310 (N_16310,N_12162,N_11259);
xor U16311 (N_16311,N_10264,N_12759);
xor U16312 (N_16312,N_14903,N_10338);
nand U16313 (N_16313,N_13031,N_13673);
xor U16314 (N_16314,N_11702,N_14451);
nand U16315 (N_16315,N_10020,N_11581);
xnor U16316 (N_16316,N_11334,N_10105);
or U16317 (N_16317,N_12372,N_11885);
or U16318 (N_16318,N_14775,N_13469);
nor U16319 (N_16319,N_13476,N_14658);
xor U16320 (N_16320,N_11998,N_13462);
or U16321 (N_16321,N_10445,N_13739);
xnor U16322 (N_16322,N_13308,N_10428);
and U16323 (N_16323,N_13804,N_10068);
and U16324 (N_16324,N_13295,N_14731);
xor U16325 (N_16325,N_10278,N_12708);
and U16326 (N_16326,N_14063,N_13036);
nor U16327 (N_16327,N_12030,N_14983);
or U16328 (N_16328,N_10383,N_13617);
xor U16329 (N_16329,N_10217,N_13644);
xor U16330 (N_16330,N_12115,N_13818);
nor U16331 (N_16331,N_11489,N_10946);
and U16332 (N_16332,N_13113,N_13109);
and U16333 (N_16333,N_11245,N_10182);
xnor U16334 (N_16334,N_11846,N_12765);
nand U16335 (N_16335,N_12055,N_11328);
xor U16336 (N_16336,N_10640,N_11743);
nand U16337 (N_16337,N_10253,N_11597);
nor U16338 (N_16338,N_12874,N_12186);
or U16339 (N_16339,N_10794,N_10732);
nand U16340 (N_16340,N_11807,N_12141);
nor U16341 (N_16341,N_12017,N_12547);
nor U16342 (N_16342,N_11088,N_12870);
nand U16343 (N_16343,N_11526,N_13139);
or U16344 (N_16344,N_12351,N_10364);
xor U16345 (N_16345,N_11091,N_11182);
xnor U16346 (N_16346,N_12290,N_12817);
nand U16347 (N_16347,N_14458,N_13107);
nand U16348 (N_16348,N_12377,N_13525);
xor U16349 (N_16349,N_14963,N_10639);
xnor U16350 (N_16350,N_14283,N_11068);
xnor U16351 (N_16351,N_14807,N_11277);
or U16352 (N_16352,N_11005,N_14737);
or U16353 (N_16353,N_13781,N_13093);
and U16354 (N_16354,N_10819,N_10153);
or U16355 (N_16355,N_11050,N_10487);
nand U16356 (N_16356,N_10151,N_10257);
or U16357 (N_16357,N_11093,N_11227);
or U16358 (N_16358,N_11019,N_11204);
nor U16359 (N_16359,N_11684,N_13174);
or U16360 (N_16360,N_11888,N_10495);
xnor U16361 (N_16361,N_11422,N_12933);
nor U16362 (N_16362,N_13549,N_13428);
or U16363 (N_16363,N_12165,N_13746);
and U16364 (N_16364,N_10326,N_10022);
nand U16365 (N_16365,N_11196,N_11387);
or U16366 (N_16366,N_11870,N_10654);
xor U16367 (N_16367,N_10312,N_14198);
nor U16368 (N_16368,N_12648,N_12875);
and U16369 (N_16369,N_10992,N_12626);
nand U16370 (N_16370,N_11406,N_12784);
nor U16371 (N_16371,N_10606,N_13361);
xnor U16372 (N_16372,N_12577,N_12083);
nand U16373 (N_16373,N_12209,N_14140);
or U16374 (N_16374,N_14868,N_12534);
nor U16375 (N_16375,N_10302,N_12101);
and U16376 (N_16376,N_10051,N_11930);
xnor U16377 (N_16377,N_13411,N_12273);
nor U16378 (N_16378,N_10698,N_13793);
xor U16379 (N_16379,N_10116,N_10317);
nand U16380 (N_16380,N_13921,N_11626);
xor U16381 (N_16381,N_13357,N_13252);
and U16382 (N_16382,N_11986,N_13154);
or U16383 (N_16383,N_10880,N_13246);
or U16384 (N_16384,N_14305,N_10832);
or U16385 (N_16385,N_10689,N_14941);
nand U16386 (N_16386,N_13454,N_13660);
or U16387 (N_16387,N_14340,N_11418);
and U16388 (N_16388,N_14662,N_14344);
nand U16389 (N_16389,N_13383,N_12801);
and U16390 (N_16390,N_12974,N_14714);
and U16391 (N_16391,N_12048,N_11300);
nand U16392 (N_16392,N_13791,N_11184);
or U16393 (N_16393,N_10791,N_14212);
or U16394 (N_16394,N_13232,N_13520);
nor U16395 (N_16395,N_11973,N_11353);
or U16396 (N_16396,N_10478,N_10031);
xor U16397 (N_16397,N_10045,N_12378);
nor U16398 (N_16398,N_12179,N_13030);
or U16399 (N_16399,N_10088,N_10733);
and U16400 (N_16400,N_14292,N_12846);
nand U16401 (N_16401,N_11309,N_14025);
or U16402 (N_16402,N_14078,N_12233);
nand U16403 (N_16403,N_13257,N_10089);
or U16404 (N_16404,N_13385,N_13409);
xor U16405 (N_16405,N_11892,N_14142);
nor U16406 (N_16406,N_14092,N_13087);
nor U16407 (N_16407,N_11190,N_11662);
and U16408 (N_16408,N_13444,N_12144);
and U16409 (N_16409,N_10384,N_13894);
nor U16410 (N_16410,N_12338,N_14141);
or U16411 (N_16411,N_12189,N_11605);
nor U16412 (N_16412,N_11313,N_11989);
or U16413 (N_16413,N_14501,N_11575);
nand U16414 (N_16414,N_14264,N_10548);
nor U16415 (N_16415,N_12655,N_14361);
xor U16416 (N_16416,N_11871,N_14743);
nand U16417 (N_16417,N_11763,N_11257);
nand U16418 (N_16418,N_11744,N_13561);
nor U16419 (N_16419,N_14156,N_14532);
nand U16420 (N_16420,N_12821,N_11847);
and U16421 (N_16421,N_12586,N_11651);
nand U16422 (N_16422,N_11827,N_10882);
xor U16423 (N_16423,N_10197,N_13277);
nor U16424 (N_16424,N_11630,N_14362);
and U16425 (N_16425,N_14339,N_12376);
nand U16426 (N_16426,N_13840,N_12363);
nand U16427 (N_16427,N_14429,N_11216);
or U16428 (N_16428,N_12973,N_12095);
or U16429 (N_16429,N_14193,N_11915);
xor U16430 (N_16430,N_13121,N_12422);
xnor U16431 (N_16431,N_10135,N_11776);
and U16432 (N_16432,N_13515,N_14878);
nand U16433 (N_16433,N_11234,N_13455);
xnor U16434 (N_16434,N_10657,N_11021);
and U16435 (N_16435,N_10374,N_10012);
and U16436 (N_16436,N_14235,N_12633);
or U16437 (N_16437,N_14649,N_13240);
or U16438 (N_16438,N_13712,N_13915);
nand U16439 (N_16439,N_12406,N_14285);
or U16440 (N_16440,N_14617,N_11373);
nand U16441 (N_16441,N_12183,N_14835);
nand U16442 (N_16442,N_10377,N_10976);
or U16443 (N_16443,N_12859,N_13625);
nor U16444 (N_16444,N_14389,N_13883);
nand U16445 (N_16445,N_14126,N_11991);
or U16446 (N_16446,N_12072,N_13323);
and U16447 (N_16447,N_10884,N_13744);
nand U16448 (N_16448,N_14504,N_12698);
nor U16449 (N_16449,N_12138,N_13394);
nor U16450 (N_16450,N_10358,N_10044);
and U16451 (N_16451,N_10117,N_12931);
nor U16452 (N_16452,N_11557,N_12727);
or U16453 (N_16453,N_12596,N_10122);
xor U16454 (N_16454,N_10610,N_11572);
and U16455 (N_16455,N_14237,N_11413);
or U16456 (N_16456,N_13911,N_13557);
or U16457 (N_16457,N_12133,N_11161);
and U16458 (N_16458,N_11518,N_13306);
nand U16459 (N_16459,N_10660,N_10288);
nand U16460 (N_16460,N_10268,N_12905);
nand U16461 (N_16461,N_10258,N_13165);
or U16462 (N_16462,N_10817,N_10188);
nand U16463 (N_16463,N_13058,N_13798);
xor U16464 (N_16464,N_10942,N_10756);
xnor U16465 (N_16465,N_14124,N_10684);
xnor U16466 (N_16466,N_10616,N_11332);
nor U16467 (N_16467,N_13270,N_10043);
xor U16468 (N_16468,N_11561,N_12110);
xor U16469 (N_16469,N_11084,N_10303);
nor U16470 (N_16470,N_14349,N_12881);
nand U16471 (N_16471,N_10419,N_12321);
xnor U16472 (N_16472,N_11947,N_13529);
nand U16473 (N_16473,N_13055,N_14410);
xor U16474 (N_16474,N_10642,N_11564);
and U16475 (N_16475,N_13460,N_11750);
or U16476 (N_16476,N_13080,N_14924);
nor U16477 (N_16477,N_13057,N_13726);
nand U16478 (N_16478,N_11718,N_11060);
nor U16479 (N_16479,N_11663,N_11795);
or U16480 (N_16480,N_14066,N_11671);
and U16481 (N_16481,N_13839,N_11176);
and U16482 (N_16482,N_11539,N_13949);
or U16483 (N_16483,N_13870,N_11650);
nand U16484 (N_16484,N_14454,N_14321);
xnor U16485 (N_16485,N_12664,N_14384);
nand U16486 (N_16486,N_12015,N_13227);
and U16487 (N_16487,N_11491,N_12119);
xor U16488 (N_16488,N_13296,N_14902);
and U16489 (N_16489,N_10385,N_14524);
xor U16490 (N_16490,N_12481,N_13519);
and U16491 (N_16491,N_13626,N_10869);
xnor U16492 (N_16492,N_13152,N_14437);
or U16493 (N_16493,N_14781,N_14965);
and U16494 (N_16494,N_13596,N_14129);
nor U16495 (N_16495,N_13331,N_10481);
nor U16496 (N_16496,N_11681,N_12085);
nor U16497 (N_16497,N_11968,N_12857);
and U16498 (N_16498,N_13155,N_14353);
or U16499 (N_16499,N_10079,N_13376);
xnor U16500 (N_16500,N_11082,N_12844);
nor U16501 (N_16501,N_10298,N_13160);
nand U16502 (N_16502,N_10256,N_12475);
or U16503 (N_16503,N_10231,N_12730);
or U16504 (N_16504,N_10355,N_14523);
and U16505 (N_16505,N_14164,N_10860);
and U16506 (N_16506,N_10281,N_12669);
nand U16507 (N_16507,N_11498,N_12854);
or U16508 (N_16508,N_12009,N_14186);
xor U16509 (N_16509,N_10892,N_10851);
xnor U16510 (N_16510,N_10895,N_12123);
xor U16511 (N_16511,N_10718,N_12871);
and U16512 (N_16512,N_11179,N_11982);
and U16513 (N_16513,N_12986,N_12657);
xor U16514 (N_16514,N_11801,N_13259);
and U16515 (N_16515,N_14179,N_14473);
and U16516 (N_16516,N_11668,N_13074);
xnor U16517 (N_16517,N_11238,N_14620);
xor U16518 (N_16518,N_14694,N_10607);
xnor U16519 (N_16519,N_10114,N_10753);
nand U16520 (N_16520,N_14275,N_12660);
or U16521 (N_16521,N_13176,N_10865);
or U16522 (N_16522,N_13992,N_13878);
xor U16523 (N_16523,N_12524,N_13846);
xnor U16524 (N_16524,N_11444,N_14889);
xnor U16525 (N_16525,N_12227,N_11694);
nor U16526 (N_16526,N_12830,N_10319);
nor U16527 (N_16527,N_10085,N_13208);
nor U16528 (N_16528,N_12405,N_13442);
nand U16529 (N_16529,N_12883,N_11791);
nor U16530 (N_16530,N_10988,N_12552);
xnor U16531 (N_16531,N_13615,N_14489);
nand U16532 (N_16532,N_12506,N_14401);
xnor U16533 (N_16533,N_14660,N_11421);
nand U16534 (N_16534,N_13652,N_12069);
xor U16535 (N_16535,N_12028,N_13231);
nand U16536 (N_16536,N_13914,N_13909);
nand U16537 (N_16537,N_12943,N_14227);
or U16538 (N_16538,N_10669,N_14646);
nor U16539 (N_16539,N_14290,N_11174);
nand U16540 (N_16540,N_13888,N_10746);
xor U16541 (N_16541,N_12722,N_12292);
and U16542 (N_16542,N_12229,N_11308);
or U16543 (N_16543,N_13400,N_11451);
xnor U16544 (N_16544,N_13313,N_10076);
nand U16545 (N_16545,N_10745,N_12333);
xnor U16546 (N_16546,N_10485,N_12878);
xor U16547 (N_16547,N_10132,N_10963);
or U16548 (N_16548,N_12723,N_10775);
and U16549 (N_16549,N_14014,N_14586);
nor U16550 (N_16550,N_14406,N_12990);
nand U16551 (N_16551,N_14195,N_11882);
and U16552 (N_16552,N_13369,N_11293);
or U16553 (N_16553,N_12989,N_14744);
nor U16554 (N_16554,N_13842,N_11089);
xor U16555 (N_16555,N_14922,N_10982);
or U16556 (N_16556,N_11228,N_11317);
nor U16557 (N_16557,N_12930,N_11183);
nand U16558 (N_16558,N_13643,N_14304);
xnor U16559 (N_16559,N_10001,N_13614);
xnor U16560 (N_16560,N_13951,N_12670);
and U16561 (N_16561,N_10075,N_12726);
or U16562 (N_16562,N_12341,N_12160);
or U16563 (N_16563,N_11725,N_14100);
xnor U16564 (N_16564,N_11483,N_12977);
xor U16565 (N_16565,N_14173,N_12928);
xnor U16566 (N_16566,N_11966,N_13463);
nand U16567 (N_16567,N_11538,N_14892);
or U16568 (N_16568,N_11934,N_13706);
nand U16569 (N_16569,N_11331,N_13664);
and U16570 (N_16570,N_12588,N_12196);
xor U16571 (N_16571,N_13709,N_10532);
nor U16572 (N_16572,N_14175,N_10368);
xnor U16573 (N_16573,N_11592,N_13876);
xnor U16574 (N_16574,N_11240,N_12428);
nand U16575 (N_16575,N_12713,N_11582);
and U16576 (N_16576,N_13488,N_14001);
or U16577 (N_16577,N_12014,N_14613);
nor U16578 (N_16578,N_11933,N_10731);
and U16579 (N_16579,N_10134,N_10679);
nor U16580 (N_16580,N_11163,N_12975);
xnor U16581 (N_16581,N_14712,N_11931);
or U16582 (N_16582,N_10968,N_10422);
or U16583 (N_16583,N_11632,N_13286);
and U16584 (N_16584,N_13389,N_11826);
xor U16585 (N_16585,N_14483,N_14865);
or U16586 (N_16586,N_11323,N_13967);
nand U16587 (N_16587,N_13771,N_13498);
and U16588 (N_16588,N_14653,N_13393);
or U16589 (N_16589,N_14073,N_13122);
nor U16590 (N_16590,N_10046,N_13090);
nand U16591 (N_16591,N_12367,N_13595);
nor U16592 (N_16592,N_10957,N_12653);
nor U16593 (N_16593,N_13214,N_14446);
xor U16594 (N_16594,N_10803,N_12949);
nand U16595 (N_16595,N_11877,N_11995);
nand U16596 (N_16596,N_10969,N_10410);
xor U16597 (N_16597,N_10887,N_13578);
xor U16598 (N_16598,N_12414,N_10949);
or U16599 (N_16599,N_10499,N_13371);
xor U16600 (N_16600,N_10097,N_11135);
xor U16601 (N_16601,N_13604,N_10948);
nand U16602 (N_16602,N_14412,N_11887);
xnor U16603 (N_16603,N_10715,N_13986);
nor U16604 (N_16604,N_13800,N_14574);
or U16605 (N_16605,N_13446,N_12731);
nor U16606 (N_16606,N_11125,N_14000);
or U16607 (N_16607,N_11562,N_12984);
xor U16608 (N_16608,N_11282,N_11215);
or U16609 (N_16609,N_13499,N_12938);
or U16610 (N_16610,N_10513,N_11223);
xor U16611 (N_16611,N_10550,N_13449);
and U16612 (N_16612,N_10245,N_12280);
nand U16613 (N_16613,N_14844,N_10069);
nand U16614 (N_16614,N_11645,N_11962);
and U16615 (N_16615,N_14192,N_12025);
xor U16616 (N_16616,N_13590,N_14106);
xor U16617 (N_16617,N_12218,N_14809);
xor U16618 (N_16618,N_13378,N_13605);
nor U16619 (N_16619,N_13528,N_13297);
or U16620 (N_16620,N_10211,N_13305);
xnor U16621 (N_16621,N_14940,N_12291);
nor U16622 (N_16622,N_14830,N_12118);
and U16623 (N_16623,N_10157,N_14416);
or U16624 (N_16624,N_13204,N_11159);
nand U16625 (N_16625,N_14213,N_12649);
or U16626 (N_16626,N_10886,N_11797);
nor U16627 (N_16627,N_13116,N_13895);
and U16628 (N_16628,N_10029,N_11452);
and U16629 (N_16629,N_14371,N_10380);
nor U16630 (N_16630,N_11900,N_13727);
nor U16631 (N_16631,N_14848,N_14110);
xnor U16632 (N_16632,N_10362,N_10240);
nand U16633 (N_16633,N_11408,N_13474);
or U16634 (N_16634,N_13849,N_10742);
nand U16635 (N_16635,N_11903,N_13147);
nor U16636 (N_16636,N_11880,N_14394);
nor U16637 (N_16637,N_10635,N_10825);
nand U16638 (N_16638,N_11358,N_12831);
and U16639 (N_16639,N_12070,N_14538);
nand U16640 (N_16640,N_12024,N_12662);
nor U16641 (N_16641,N_13300,N_13881);
nand U16642 (N_16642,N_11144,N_11925);
nor U16643 (N_16643,N_14029,N_10814);
xnor U16644 (N_16644,N_11985,N_12066);
xnor U16645 (N_16645,N_10973,N_14203);
and U16646 (N_16646,N_10883,N_11352);
or U16647 (N_16647,N_12738,N_10403);
xnor U16648 (N_16648,N_13944,N_13423);
xor U16649 (N_16649,N_14355,N_11180);
and U16650 (N_16650,N_12421,N_12561);
xnor U16651 (N_16651,N_11573,N_10147);
and U16652 (N_16652,N_11160,N_14890);
or U16653 (N_16653,N_12221,N_10357);
nand U16654 (N_16654,N_10754,N_12551);
nand U16655 (N_16655,N_12932,N_10431);
nor U16656 (N_16656,N_11673,N_10395);
and U16657 (N_16657,N_14372,N_10159);
or U16658 (N_16658,N_14017,N_14249);
nor U16659 (N_16659,N_13338,N_10406);
nand U16660 (N_16660,N_12772,N_14332);
nand U16661 (N_16661,N_14769,N_14038);
or U16662 (N_16662,N_10131,N_14240);
or U16663 (N_16663,N_11201,N_12276);
nand U16664 (N_16664,N_13546,N_12472);
nand U16665 (N_16665,N_11712,N_13702);
nand U16666 (N_16666,N_14946,N_13464);
and U16667 (N_16667,N_13065,N_11286);
and U16668 (N_16668,N_11935,N_14231);
xnor U16669 (N_16669,N_11607,N_14742);
xor U16670 (N_16670,N_13965,N_14112);
xor U16671 (N_16671,N_14223,N_14582);
nand U16672 (N_16672,N_11058,N_13822);
nand U16673 (N_16673,N_12962,N_11574);
nor U16674 (N_16674,N_11069,N_10082);
nor U16675 (N_16675,N_12589,N_13018);
and U16676 (N_16676,N_10273,N_14962);
nor U16677 (N_16677,N_11200,N_12452);
nand U16678 (N_16678,N_12454,N_10350);
xnor U16679 (N_16679,N_14178,N_10827);
and U16680 (N_16680,N_10244,N_14266);
xnor U16681 (N_16681,N_14506,N_10987);
and U16682 (N_16682,N_13602,N_13435);
nor U16683 (N_16683,N_11269,N_10805);
nor U16684 (N_16684,N_11015,N_11009);
or U16685 (N_16685,N_14553,N_14241);
nor U16686 (N_16686,N_11772,N_10985);
nor U16687 (N_16687,N_11048,N_12624);
or U16688 (N_16688,N_11056,N_11875);
xor U16689 (N_16689,N_11487,N_13832);
xor U16690 (N_16690,N_12199,N_14091);
nand U16691 (N_16691,N_11378,N_12659);
nor U16692 (N_16692,N_10704,N_11578);
or U16693 (N_16693,N_10334,N_13756);
nand U16694 (N_16694,N_10224,N_12402);
nand U16695 (N_16695,N_11481,N_14753);
nor U16696 (N_16696,N_14087,N_14850);
nand U16697 (N_16697,N_13415,N_14238);
xor U16698 (N_16698,N_13942,N_13169);
nand U16699 (N_16699,N_12112,N_12293);
and U16700 (N_16700,N_11604,N_14252);
nor U16701 (N_16701,N_13823,N_14923);
nor U16702 (N_16702,N_10342,N_12373);
nor U16703 (N_16703,N_13392,N_11723);
or U16704 (N_16704,N_11535,N_14910);
nand U16705 (N_16705,N_14857,N_12853);
or U16706 (N_16706,N_11276,N_12168);
nand U16707 (N_16707,N_10490,N_13325);
and U16708 (N_16708,N_11112,N_11965);
xnor U16709 (N_16709,N_13479,N_13675);
nand U16710 (N_16710,N_12527,N_10206);
nor U16711 (N_16711,N_11550,N_10806);
nand U16712 (N_16712,N_13730,N_10580);
nand U16713 (N_16713,N_11856,N_10497);
nor U16714 (N_16714,N_12640,N_14810);
nor U16715 (N_16715,N_11679,N_14709);
nand U16716 (N_16716,N_13753,N_10720);
or U16717 (N_16717,N_14645,N_10842);
xor U16718 (N_16718,N_12944,N_12456);
xnor U16719 (N_16719,N_10735,N_14776);
nand U16720 (N_16720,N_10468,N_12896);
or U16721 (N_16721,N_11838,N_13687);
nor U16722 (N_16722,N_13611,N_14726);
nor U16723 (N_16723,N_10246,N_10510);
and U16724 (N_16724,N_12214,N_10344);
and U16725 (N_16725,N_14790,N_14797);
xnor U16726 (N_16726,N_13230,N_11813);
nand U16727 (N_16727,N_10306,N_13182);
nand U16728 (N_16728,N_11890,N_12694);
xnor U16729 (N_16729,N_14357,N_11865);
and U16730 (N_16730,N_12704,N_13408);
or U16731 (N_16731,N_10480,N_11939);
nor U16732 (N_16732,N_10599,N_11924);
xnor U16733 (N_16733,N_14042,N_10167);
xor U16734 (N_16734,N_11129,N_14732);
or U16735 (N_16735,N_11239,N_12304);
xnor U16736 (N_16736,N_14253,N_11281);
and U16737 (N_16737,N_10736,N_10083);
and U16738 (N_16738,N_10582,N_14803);
nor U16739 (N_16739,N_14135,N_12379);
xor U16740 (N_16740,N_12776,N_12315);
nor U16741 (N_16741,N_12294,N_12433);
or U16742 (N_16742,N_14132,N_12841);
xor U16743 (N_16743,N_13002,N_14701);
or U16744 (N_16744,N_10025,N_11619);
and U16745 (N_16745,N_10369,N_14500);
and U16746 (N_16746,N_13309,N_10464);
xnor U16747 (N_16747,N_11851,N_11755);
xnor U16748 (N_16748,N_14251,N_11044);
nor U16749 (N_16749,N_11342,N_12350);
xnor U16750 (N_16750,N_12407,N_14551);
and U16751 (N_16751,N_11434,N_12798);
nor U16752 (N_16752,N_12004,N_12389);
and U16753 (N_16753,N_14736,N_14704);
nor U16754 (N_16754,N_13421,N_11932);
nand U16755 (N_16755,N_11327,N_10473);
nand U16756 (N_16756,N_12560,N_12646);
nand U16757 (N_16757,N_13478,N_10983);
nand U16758 (N_16758,N_11756,N_11186);
xnor U16759 (N_16759,N_12505,N_10186);
nor U16760 (N_16760,N_10593,N_10611);
and U16761 (N_16761,N_14209,N_10331);
nand U16762 (N_16762,N_12013,N_14534);
nor U16763 (N_16763,N_14434,N_13189);
xor U16764 (N_16764,N_12502,N_11964);
or U16765 (N_16765,N_11734,N_12894);
xor U16766 (N_16766,N_13172,N_14050);
nor U16767 (N_16767,N_12923,N_13608);
nor U16768 (N_16768,N_11860,N_14119);
or U16769 (N_16769,N_14521,N_12934);
xor U16770 (N_16770,N_13466,N_13696);
nor U16771 (N_16771,N_14686,N_13809);
or U16772 (N_16772,N_12635,N_12545);
nor U16773 (N_16773,N_10812,N_12645);
nand U16774 (N_16774,N_13045,N_12352);
and U16775 (N_16775,N_10056,N_10998);
nor U16776 (N_16776,N_14516,N_12921);
nor U16777 (N_16777,N_11999,N_10683);
xor U16778 (N_16778,N_14390,N_14548);
or U16779 (N_16779,N_10927,N_14815);
or U16780 (N_16780,N_13440,N_10200);
or U16781 (N_16781,N_14108,N_13289);
nand U16782 (N_16782,N_12705,N_12418);
nor U16783 (N_16783,N_11471,N_14787);
or U16784 (N_16784,N_13006,N_12700);
or U16785 (N_16785,N_11955,N_14230);
nand U16786 (N_16786,N_11513,N_10696);
xnor U16787 (N_16787,N_12566,N_14041);
nor U16788 (N_16788,N_12279,N_10321);
xor U16789 (N_16789,N_12255,N_13723);
nand U16790 (N_16790,N_10389,N_10039);
nand U16791 (N_16791,N_12613,N_11416);
nor U16792 (N_16792,N_11858,N_12823);
and U16793 (N_16793,N_13917,N_13085);
nor U16794 (N_16794,N_13983,N_13150);
nor U16795 (N_16795,N_13514,N_12215);
nor U16796 (N_16796,N_11229,N_12181);
and U16797 (N_16797,N_11436,N_11850);
and U16798 (N_16798,N_13560,N_13432);
or U16799 (N_16799,N_14843,N_11181);
xnor U16800 (N_16800,N_13001,N_14680);
and U16801 (N_16801,N_11563,N_14259);
or U16802 (N_16802,N_13118,N_11351);
nor U16803 (N_16803,N_11854,N_11656);
xnor U16804 (N_16804,N_10129,N_10505);
xor U16805 (N_16805,N_13936,N_13955);
and U16806 (N_16806,N_13168,N_14174);
nor U16807 (N_16807,N_10786,N_10073);
or U16808 (N_16808,N_14460,N_14513);
nand U16809 (N_16809,N_13689,N_11844);
and U16810 (N_16810,N_13517,N_12889);
nor U16811 (N_16811,N_12325,N_12146);
nand U16812 (N_16812,N_10917,N_12267);
nand U16813 (N_16813,N_14599,N_10386);
nand U16814 (N_16814,N_11222,N_11891);
nor U16815 (N_16815,N_14373,N_11153);
nor U16816 (N_16816,N_14419,N_14541);
nor U16817 (N_16817,N_11778,N_12037);
nand U16818 (N_16818,N_12557,N_10714);
or U16819 (N_16819,N_10393,N_10815);
nand U16820 (N_16820,N_10351,N_14428);
xor U16821 (N_16821,N_12639,N_12060);
and U16822 (N_16822,N_10266,N_12182);
nand U16823 (N_16823,N_12836,N_11596);
nand U16824 (N_16824,N_12499,N_12058);
or U16825 (N_16825,N_14138,N_11459);
xor U16826 (N_16826,N_11504,N_10015);
nor U16827 (N_16827,N_10287,N_11691);
nor U16828 (N_16828,N_14184,N_12495);
nand U16829 (N_16829,N_10400,N_13941);
and U16830 (N_16830,N_14139,N_14579);
and U16831 (N_16831,N_11298,N_11818);
and U16832 (N_16832,N_13755,N_13024);
or U16833 (N_16833,N_12006,N_14376);
nor U16834 (N_16834,N_12525,N_10213);
nor U16835 (N_16835,N_12441,N_13332);
and U16836 (N_16836,N_14234,N_11545);
nor U16837 (N_16837,N_11948,N_12207);
nand U16838 (N_16838,N_11859,N_10557);
nor U16839 (N_16839,N_12275,N_14216);
and U16840 (N_16840,N_11214,N_14022);
and U16841 (N_16841,N_11623,N_13902);
or U16842 (N_16842,N_12408,N_10541);
nor U16843 (N_16843,N_12041,N_12824);
or U16844 (N_16844,N_13841,N_14395);
nand U16845 (N_16845,N_10970,N_10327);
xor U16846 (N_16846,N_14629,N_10002);
and U16847 (N_16847,N_13315,N_13108);
xor U16848 (N_16848,N_13416,N_14226);
or U16849 (N_16849,N_13612,N_12978);
or U16850 (N_16850,N_12838,N_12135);
xnor U16851 (N_16851,N_10780,N_12466);
nand U16852 (N_16852,N_12579,N_13403);
and U16853 (N_16853,N_12797,N_11035);
and U16854 (N_16854,N_11970,N_14443);
nand U16855 (N_16855,N_14638,N_12326);
or U16856 (N_16856,N_14246,N_10687);
xnor U16857 (N_16857,N_12804,N_14296);
nor U16858 (N_16858,N_12149,N_14956);
or U16859 (N_16859,N_11514,N_14626);
xor U16860 (N_16860,N_11017,N_12384);
or U16861 (N_16861,N_14974,N_14358);
or U16862 (N_16862,N_14651,N_12684);
nor U16863 (N_16863,N_10512,N_12023);
or U16864 (N_16864,N_10846,N_14046);
xor U16865 (N_16865,N_12081,N_14306);
and U16866 (N_16866,N_12465,N_14051);
or U16867 (N_16867,N_12416,N_11969);
nor U16868 (N_16868,N_11080,N_14652);
nand U16869 (N_16869,N_11362,N_10227);
xnor U16870 (N_16870,N_12802,N_10027);
nor U16871 (N_16871,N_10975,N_14817);
xor U16872 (N_16872,N_12252,N_11719);
or U16873 (N_16873,N_13754,N_13631);
or U16874 (N_16874,N_12810,N_12807);
xor U16875 (N_16875,N_13788,N_13758);
and U16876 (N_16876,N_10347,N_12038);
and U16877 (N_16877,N_10314,N_13233);
nand U16878 (N_16878,N_14723,N_14335);
nand U16879 (N_16879,N_13562,N_14293);
or U16880 (N_16880,N_10229,N_13581);
nand U16881 (N_16881,N_14618,N_14720);
xnor U16882 (N_16882,N_11398,N_11115);
and U16883 (N_16883,N_12432,N_13033);
nand U16884 (N_16884,N_11984,N_11606);
or U16885 (N_16885,N_12241,N_13487);
nand U16886 (N_16886,N_13873,N_10713);
and U16887 (N_16887,N_12420,N_10160);
nor U16888 (N_16888,N_13872,N_14274);
nor U16889 (N_16889,N_12370,N_13335);
nand U16890 (N_16890,N_13267,N_14970);
nor U16891 (N_16891,N_10868,N_14760);
xnor U16892 (N_16892,N_14172,N_11485);
or U16893 (N_16893,N_11811,N_14089);
xor U16894 (N_16894,N_13370,N_10874);
nor U16895 (N_16895,N_13177,N_13052);
and U16896 (N_16896,N_14847,N_13912);
and U16897 (N_16897,N_10893,N_11711);
or U16898 (N_16898,N_13591,N_13742);
and U16899 (N_16899,N_10032,N_12190);
and U16900 (N_16900,N_13703,N_12491);
or U16901 (N_16901,N_10235,N_13334);
and U16902 (N_16902,N_10538,N_10900);
nor U16903 (N_16903,N_12362,N_11024);
xor U16904 (N_16904,N_12828,N_13144);
xnor U16905 (N_16905,N_11000,N_14671);
xor U16906 (N_16906,N_10373,N_12073);
and U16907 (N_16907,N_14105,N_13429);
nor U16908 (N_16908,N_10879,N_14342);
or U16909 (N_16909,N_11503,N_12911);
xnor U16910 (N_16910,N_14286,N_11586);
and U16911 (N_16911,N_10690,N_13318);
nor U16912 (N_16912,N_14006,N_14472);
xor U16913 (N_16913,N_13829,N_12397);
and U16914 (N_16914,N_11646,N_14442);
nor U16915 (N_16915,N_13008,N_12885);
nor U16916 (N_16916,N_11002,N_14824);
xor U16917 (N_16917,N_12837,N_12392);
xor U16918 (N_16918,N_11852,N_11251);
nand U16919 (N_16919,N_14778,N_14872);
or U16920 (N_16920,N_10779,N_10243);
nand U16921 (N_16921,N_13229,N_10737);
and U16922 (N_16922,N_13651,N_11994);
nand U16923 (N_16923,N_10305,N_14556);
or U16924 (N_16924,N_12476,N_11665);
nor U16925 (N_16925,N_14055,N_10219);
nand U16926 (N_16926,N_13410,N_11845);
nor U16927 (N_16927,N_10145,N_12339);
and U16928 (N_16928,N_14417,N_13684);
nand U16929 (N_16929,N_10322,N_12068);
xnor U16930 (N_16930,N_13808,N_13593);
and U16931 (N_16931,N_10233,N_11922);
and U16932 (N_16932,N_11963,N_10063);
or U16933 (N_16933,N_14004,N_11765);
nand U16934 (N_16934,N_13777,N_14323);
and U16935 (N_16935,N_14282,N_11086);
xor U16936 (N_16936,N_13317,N_11394);
or U16937 (N_16937,N_12490,N_14518);
nand U16938 (N_16938,N_14439,N_11977);
nand U16939 (N_16939,N_13880,N_12585);
or U16940 (N_16940,N_13623,N_13861);
xnor U16941 (N_16941,N_11520,N_12360);
or U16942 (N_16942,N_11992,N_12668);
nand U16943 (N_16943,N_10133,N_10411);
or U16944 (N_16944,N_12052,N_12496);
nand U16945 (N_16945,N_14552,N_14788);
nand U16946 (N_16946,N_13483,N_12008);
and U16947 (N_16947,N_11614,N_13655);
xnor U16948 (N_16948,N_13126,N_14612);
nand U16949 (N_16949,N_11403,N_14834);
or U16950 (N_16950,N_13629,N_10189);
nand U16951 (N_16951,N_12680,N_12543);
nand U16952 (N_16952,N_13985,N_13339);
or U16953 (N_16953,N_12231,N_13072);
nor U16954 (N_16954,N_12583,N_12880);
and U16955 (N_16955,N_14484,N_14926);
or U16956 (N_16956,N_12302,N_10943);
and U16957 (N_16957,N_11437,N_11131);
xnor U16958 (N_16958,N_13186,N_10835);
and U16959 (N_16959,N_13380,N_10906);
nand U16960 (N_16960,N_13128,N_12509);
nand U16961 (N_16961,N_14901,N_10221);
or U16962 (N_16962,N_10178,N_11819);
xnor U16963 (N_16963,N_12761,N_13321);
nand U16964 (N_16964,N_14433,N_14075);
nor U16965 (N_16965,N_14245,N_11709);
nand U16966 (N_16966,N_11254,N_11333);
nor U16967 (N_16967,N_11537,N_11124);
or U16968 (N_16968,N_12927,N_11469);
nor U16969 (N_16969,N_12847,N_12096);
xnor U16970 (N_16970,N_11751,N_11585);
xor U16971 (N_16971,N_10070,N_11548);
and U16972 (N_16972,N_12541,N_12825);
nand U16973 (N_16973,N_11536,N_12876);
and U16974 (N_16974,N_12852,N_12091);
xor U16975 (N_16975,N_10766,N_11629);
nand U16976 (N_16976,N_11049,N_12187);
and U16977 (N_16977,N_14509,N_10594);
nor U16978 (N_16978,N_11365,N_14784);
nand U16979 (N_16979,N_10099,N_10658);
xor U16980 (N_16980,N_10774,N_14930);
and U16981 (N_16981,N_10569,N_11232);
and U16982 (N_16982,N_14402,N_12712);
nand U16983 (N_16983,N_10556,N_14116);
nor U16984 (N_16984,N_14491,N_14031);
nand U16985 (N_16985,N_12654,N_10391);
xnor U16986 (N_16986,N_11884,N_11028);
or U16987 (N_16987,N_12811,N_10320);
nand U16988 (N_16988,N_13009,N_14056);
nand U16989 (N_16989,N_11728,N_10615);
nor U16990 (N_16990,N_14802,N_10479);
or U16991 (N_16991,N_10811,N_10451);
nand U16992 (N_16992,N_10706,N_10916);
nand U16993 (N_16993,N_13316,N_11037);
nor U16994 (N_16994,N_10036,N_11832);
nor U16995 (N_16995,N_14422,N_10154);
xor U16996 (N_16996,N_13130,N_14196);
nor U16997 (N_16997,N_14944,N_10220);
nand U16998 (N_16998,N_10155,N_11902);
and U16999 (N_16999,N_11262,N_13959);
nor U17000 (N_17000,N_13852,N_11008);
or U17001 (N_17001,N_14026,N_11283);
xnor U17002 (N_17002,N_10677,N_10804);
xnor U17003 (N_17003,N_13766,N_11010);
and U17004 (N_17004,N_10136,N_12815);
nand U17005 (N_17005,N_10176,N_14624);
and U17006 (N_17006,N_13996,N_12737);
nand U17007 (N_17007,N_13803,N_12010);
or U17008 (N_17008,N_14369,N_12812);
xnor U17009 (N_17009,N_14147,N_14977);
xnor U17010 (N_17010,N_13618,N_13070);
and U17011 (N_17011,N_11242,N_12318);
nand U17012 (N_17012,N_14133,N_12436);
or U17013 (N_17013,N_12621,N_13261);
and U17014 (N_17014,N_13157,N_14669);
xnor U17015 (N_17015,N_11400,N_12746);
nor U17016 (N_17016,N_12274,N_12510);
xnor U17017 (N_17017,N_10950,N_13736);
nor U17018 (N_17018,N_14499,N_11981);
nand U17019 (N_17019,N_13013,N_12092);
nor U17020 (N_17020,N_14013,N_14366);
nand U17021 (N_17021,N_10785,N_12774);
and U17022 (N_17022,N_13601,N_11785);
and U17023 (N_17023,N_10598,N_13301);
nor U17024 (N_17024,N_13492,N_11468);
nand U17025 (N_17025,N_12216,N_13505);
or U17026 (N_17026,N_13198,N_11848);
or U17027 (N_17027,N_10318,N_14316);
or U17028 (N_17028,N_13553,N_12340);
nor U17029 (N_17029,N_11655,N_11198);
nor U17030 (N_17030,N_13287,N_13276);
or U17031 (N_17031,N_13194,N_12760);
nand U17032 (N_17032,N_11893,N_10493);
or U17033 (N_17033,N_13330,N_13115);
and U17034 (N_17034,N_13790,N_14950);
nand U17035 (N_17035,N_10536,N_14828);
nand U17036 (N_17036,N_14424,N_13272);
xnor U17037 (N_17037,N_11087,N_12792);
and U17038 (N_17038,N_10371,N_13312);
nand U17039 (N_17039,N_13789,N_13552);
nand U17040 (N_17040,N_11247,N_14685);
nand U17041 (N_17041,N_10810,N_10402);
nand U17042 (N_17042,N_13586,N_14337);
nand U17043 (N_17043,N_11158,N_11074);
nor U17044 (N_17044,N_10650,N_13737);
nand U17045 (N_17045,N_12098,N_14917);
and U17046 (N_17046,N_14448,N_11218);
xor U17047 (N_17047,N_11041,N_10631);
nor U17048 (N_17048,N_12097,N_14365);
nor U17049 (N_17049,N_13344,N_14609);
or U17050 (N_17050,N_12044,N_14180);
nor U17051 (N_17051,N_12764,N_12337);
nor U17052 (N_17052,N_10701,N_12717);
and U17053 (N_17053,N_11531,N_10641);
nand U17054 (N_17054,N_10659,N_10626);
nand U17055 (N_17055,N_11026,N_12795);
xnor U17056 (N_17056,N_10623,N_13717);
and U17057 (N_17057,N_14190,N_11474);
or U17058 (N_17058,N_14076,N_11521);
nor U17059 (N_17059,N_12794,N_12385);
or U17060 (N_17060,N_10991,N_10199);
or U17061 (N_17061,N_12458,N_13784);
and U17062 (N_17062,N_13490,N_12806);
xnor U17063 (N_17063,N_12620,N_13459);
or U17064 (N_17064,N_11114,N_11350);
nor U17065 (N_17065,N_14345,N_14441);
and U17066 (N_17066,N_14674,N_12093);
nand U17067 (N_17067,N_14023,N_13811);
or U17068 (N_17068,N_12439,N_10203);
and U17069 (N_17069,N_14367,N_10054);
or U17070 (N_17070,N_10653,N_14490);
nor U17071 (N_17071,N_12963,N_12219);
and U17072 (N_17072,N_11834,N_13810);
and U17073 (N_17073,N_14783,N_12082);
nand U17074 (N_17074,N_11528,N_10517);
nand U17075 (N_17075,N_12253,N_10491);
and U17076 (N_17076,N_12518,N_10113);
xor U17077 (N_17077,N_12581,N_13039);
nand U17078 (N_17078,N_13337,N_14037);
and U17079 (N_17079,N_14354,N_13050);
or U17080 (N_17080,N_10108,N_11128);
xor U17081 (N_17081,N_11510,N_10875);
nor U17082 (N_17082,N_10849,N_10343);
xor U17083 (N_17083,N_13216,N_13769);
nor U17084 (N_17084,N_12813,N_10000);
nor U17085 (N_17085,N_13853,N_12540);
xor U17086 (N_17086,N_10251,N_13699);
xnor U17087 (N_17087,N_12371,N_13235);
and U17088 (N_17088,N_12359,N_11849);
and U17089 (N_17089,N_10284,N_13918);
xnor U17090 (N_17090,N_10382,N_12710);
and U17091 (N_17091,N_11271,N_11199);
nor U17092 (N_17092,N_10125,N_13539);
and U17093 (N_17093,N_13068,N_12342);
xnor U17094 (N_17094,N_13679,N_12242);
nor U17095 (N_17095,N_10308,N_14984);
nor U17096 (N_17096,N_12271,N_12131);
or U17097 (N_17097,N_14684,N_11119);
nand U17098 (N_17098,N_12961,N_14925);
nor U17099 (N_17099,N_14210,N_13932);
or U17100 (N_17100,N_10440,N_14326);
xor U17101 (N_17101,N_14912,N_10094);
nand U17102 (N_17102,N_13397,N_12623);
xnor U17103 (N_17103,N_14262,N_13075);
or U17104 (N_17104,N_12154,N_12311);
xor U17105 (N_17105,N_12324,N_13599);
or U17106 (N_17106,N_10283,N_13279);
and U17107 (N_17107,N_13768,N_10904);
or U17108 (N_17108,N_13398,N_10439);
xnor U17109 (N_17109,N_13162,N_13993);
nand U17110 (N_17110,N_14980,N_13451);
xnor U17111 (N_17111,N_13100,N_10758);
nand U17112 (N_17112,N_14152,N_13133);
or U17113 (N_17113,N_10629,N_12538);
and U17114 (N_17114,N_11494,N_10798);
nand U17115 (N_17115,N_10666,N_14806);
or U17116 (N_17116,N_14777,N_13347);
nor U17117 (N_17117,N_13205,N_11098);
and U17118 (N_17118,N_14960,N_13193);
or U17119 (N_17119,N_10500,N_14027);
xor U17120 (N_17120,N_13721,N_13848);
nor U17121 (N_17121,N_10871,N_13005);
nor U17122 (N_17122,N_11625,N_10272);
nand U17123 (N_17123,N_12208,N_13797);
nand U17124 (N_17124,N_12056,N_12260);
or U17125 (N_17125,N_11488,N_12224);
and U17126 (N_17126,N_12941,N_12634);
or U17127 (N_17127,N_11505,N_11701);
nand U17128 (N_17128,N_13662,N_12500);
xnor U17129 (N_17129,N_13963,N_13491);
and U17130 (N_17130,N_13234,N_12578);
or U17131 (N_17131,N_11263,N_12317);
or U17132 (N_17132,N_11990,N_14254);
nand U17133 (N_17133,N_13349,N_12269);
xor U17134 (N_17134,N_11831,N_12720);
and U17135 (N_17135,N_13054,N_12733);
or U17136 (N_17136,N_11189,N_10546);
nor U17137 (N_17137,N_14423,N_12937);
xnor U17138 (N_17138,N_10858,N_13778);
and U17139 (N_17139,N_11411,N_12335);
nand U17140 (N_17140,N_11980,N_14207);
and U17141 (N_17141,N_14545,N_13097);
nor U17142 (N_17142,N_10498,N_13011);
nor U17143 (N_17143,N_12860,N_13962);
and U17144 (N_17144,N_11241,N_12643);
nor U17145 (N_17145,N_14012,N_14191);
nand U17146 (N_17146,N_14571,N_13262);
nand U17147 (N_17147,N_13532,N_13850);
nor U17148 (N_17148,N_10269,N_10262);
nor U17149 (N_17149,N_14673,N_12145);
or U17150 (N_17150,N_14724,N_14312);
nand U17151 (N_17151,N_14225,N_13956);
xor U17152 (N_17152,N_10252,N_10755);
or U17153 (N_17153,N_14313,N_12816);
xor U17154 (N_17154,N_11319,N_11139);
xor U17155 (N_17155,N_11687,N_10030);
or U17156 (N_17156,N_14706,N_11314);
and U17157 (N_17157,N_10275,N_13929);
and U17158 (N_17158,N_11636,N_11419);
or U17159 (N_17159,N_12434,N_13720);
or U17160 (N_17160,N_11508,N_10577);
xor U17161 (N_17161,N_11076,N_12161);
and U17162 (N_17162,N_13779,N_10183);
and U17163 (N_17163,N_11038,N_14010);
nor U17164 (N_17164,N_10502,N_10941);
nor U17165 (N_17165,N_11786,N_12862);
nand U17166 (N_17166,N_11987,N_14829);
nor U17167 (N_17167,N_13907,N_12431);
xnor U17168 (N_17168,N_13254,N_10750);
xnor U17169 (N_17169,N_14679,N_11109);
nand U17170 (N_17170,N_10059,N_12114);
and U17171 (N_17171,N_13892,N_14770);
nand U17172 (N_17172,N_13708,N_12529);
xor U17173 (N_17173,N_12424,N_12622);
nand U17174 (N_17174,N_10415,N_10006);
xor U17175 (N_17175,N_11307,N_12090);
nor U17176 (N_17176,N_11455,N_11462);
xor U17177 (N_17177,N_10204,N_11448);
or U17178 (N_17178,N_10146,N_10651);
or U17179 (N_17179,N_13576,N_12076);
nand U17180 (N_17180,N_14823,N_14040);
xor U17181 (N_17181,N_13184,N_12976);
or U17182 (N_17182,N_14111,N_11053);
nand U17183 (N_17183,N_14270,N_10013);
xnor U17184 (N_17184,N_12429,N_14485);
nand U17185 (N_17185,N_14739,N_14637);
nor U17186 (N_17186,N_10877,N_13656);
and U17187 (N_17187,N_11461,N_13513);
or U17188 (N_17188,N_13417,N_13022);
nand U17189 (N_17189,N_12840,N_10891);
xnor U17190 (N_17190,N_11113,N_12266);
nand U17191 (N_17191,N_13752,N_14243);
nor U17192 (N_17192,N_11172,N_13748);
nor U17193 (N_17193,N_10797,N_13650);
nor U17194 (N_17194,N_10328,N_13473);
nand U17195 (N_17195,N_10901,N_13920);
nor U17196 (N_17196,N_11589,N_14120);
nor U17197 (N_17197,N_10162,N_14811);
nand U17198 (N_17198,N_12007,N_11958);
and U17199 (N_17199,N_13092,N_10702);
and U17200 (N_17200,N_12650,N_13448);
nor U17201 (N_17201,N_10282,N_10978);
or U17202 (N_17202,N_14470,N_13556);
xnor U17203 (N_17203,N_12563,N_12697);
and U17204 (N_17204,N_12130,N_10911);
nand U17205 (N_17205,N_10890,N_10571);
nand U17206 (N_17206,N_14993,N_13764);
nor U17207 (N_17207,N_12477,N_10864);
nand U17208 (N_17208,N_12864,N_10905);
or U17209 (N_17209,N_13127,N_14717);
and U17210 (N_17210,N_12173,N_11735);
xnor U17211 (N_17211,N_11040,N_14016);
or U17212 (N_17212,N_13206,N_11635);
nor U17213 (N_17213,N_14915,N_10394);
or U17214 (N_17214,N_10928,N_12556);
nand U17215 (N_17215,N_13134,N_13256);
nand U17216 (N_17216,N_12057,N_10336);
nand U17217 (N_17217,N_11226,N_10115);
xnor U17218 (N_17218,N_13635,N_14058);
nand U17219 (N_17219,N_12493,N_13690);
nor U17220 (N_17220,N_11442,N_12031);
xor U17221 (N_17221,N_10179,N_13887);
or U17222 (N_17222,N_11566,N_10583);
and U17223 (N_17223,N_10673,N_12238);
and U17224 (N_17224,N_10280,N_13366);
nand U17225 (N_17225,N_10820,N_10333);
nand U17226 (N_17226,N_12501,N_13585);
nand U17227 (N_17227,N_14242,N_10665);
nor U17228 (N_17228,N_13864,N_12565);
nand U17229 (N_17229,N_13584,N_12638);
xor U17230 (N_17230,N_11250,N_14862);
nor U17231 (N_17231,N_12724,N_12301);
or U17232 (N_17232,N_13255,N_11025);
and U17233 (N_17233,N_13345,N_13939);
or U17234 (N_17234,N_10572,N_12323);
xnor U17235 (N_17235,N_10279,N_13900);
and U17236 (N_17236,N_13676,N_13037);
and U17237 (N_17237,N_13197,N_14452);
nor U17238 (N_17238,N_12788,N_14877);
or U17239 (N_17239,N_13648,N_12656);
nand U17240 (N_17240,N_11805,N_13242);
or U17241 (N_17241,N_12959,N_14934);
and U17242 (N_17242,N_10662,N_11960);
xnor U17243 (N_17243,N_10751,N_12972);
nand U17244 (N_17244,N_10463,N_13600);
and U17245 (N_17245,N_13710,N_14587);
and U17246 (N_17246,N_11368,N_12951);
nor U17247 (N_17247,N_11833,N_14641);
and U17248 (N_17248,N_14300,N_12926);
nor U17249 (N_17249,N_10823,N_13640);
xnor U17250 (N_17250,N_14228,N_10185);
xnor U17251 (N_17251,N_10579,N_14814);
xnor U17252 (N_17252,N_12644,N_11837);
nand U17253 (N_17253,N_14498,N_11732);
nand U17254 (N_17254,N_10119,N_11953);
nor U17255 (N_17255,N_12152,N_12936);
nand U17256 (N_17256,N_13390,N_11926);
nor U17257 (N_17257,N_12075,N_12958);
xnor U17258 (N_17258,N_12120,N_14298);
and U17259 (N_17259,N_14090,N_10925);
nor U17260 (N_17260,N_14272,N_11207);
and U17261 (N_17261,N_12780,N_14550);
nor U17262 (N_17262,N_14707,N_13674);
and U17263 (N_17263,N_12116,N_12084);
xnor U17264 (N_17264,N_11366,N_11714);
nand U17265 (N_17265,N_10793,N_10149);
nor U17266 (N_17266,N_12401,N_12777);
nor U17267 (N_17267,N_10945,N_10841);
and U17268 (N_17268,N_14247,N_13132);
or U17269 (N_17269,N_12683,N_10637);
xnor U17270 (N_17270,N_13363,N_14387);
xor U17271 (N_17271,N_14113,N_13521);
xnor U17272 (N_17272,N_14870,N_11918);
or U17273 (N_17273,N_12991,N_14854);
xnor U17274 (N_17274,N_13224,N_14167);
xnor U17275 (N_17275,N_13740,N_14032);
nand U17276 (N_17276,N_10472,N_13952);
and U17277 (N_17277,N_13594,N_13021);
xor U17278 (N_17278,N_13668,N_13493);
nor U17279 (N_17279,N_10352,N_14381);
or U17280 (N_17280,N_10208,N_14279);
or U17281 (N_17281,N_14101,N_14021);
or U17282 (N_17282,N_13971,N_11004);
nand U17283 (N_17283,N_11064,N_11672);
and U17284 (N_17284,N_11710,N_10937);
and U17285 (N_17285,N_13000,N_14288);
and U17286 (N_17286,N_13835,N_11910);
nand U17287 (N_17287,N_12175,N_10453);
nand U17288 (N_17288,N_13010,N_14239);
and U17289 (N_17289,N_14153,N_12769);
xnor U17290 (N_17290,N_12460,N_10409);
nor U17291 (N_17291,N_13931,N_13571);
nand U17292 (N_17292,N_11506,N_14560);
nor U17293 (N_17293,N_14693,N_14007);
nand U17294 (N_17294,N_12907,N_11055);
nand U17295 (N_17295,N_13311,N_14457);
nor U17296 (N_17296,N_14185,N_14602);
and U17297 (N_17297,N_14578,N_11802);
and U17298 (N_17298,N_13628,N_13747);
nor U17299 (N_17299,N_13293,N_13151);
nor U17300 (N_17300,N_14048,N_12570);
xor U17301 (N_17301,N_14211,N_13695);
and U17302 (N_17302,N_12955,N_13865);
or U17303 (N_17303,N_11657,N_13226);
nor U17304 (N_17304,N_11409,N_13636);
nand U17305 (N_17305,N_11622,N_11253);
nand U17306 (N_17306,N_10367,N_13647);
xor U17307 (N_17307,N_13619,N_14082);
or U17308 (N_17308,N_12261,N_10100);
and U17309 (N_17309,N_13770,N_13974);
and U17310 (N_17310,N_13646,N_14990);
nand U17311 (N_17311,N_12879,N_12330);
nor U17312 (N_17312,N_13265,N_14897);
nor U17313 (N_17313,N_10381,N_14713);
and U17314 (N_17314,N_13327,N_12734);
xor U17315 (N_17315,N_10177,N_11057);
nand U17316 (N_17316,N_11423,N_13854);
nor U17317 (N_17317,N_13889,N_10762);
or U17318 (N_17318,N_14542,N_11330);
nand U17319 (N_17319,N_13761,N_12198);
and U17320 (N_17320,N_14622,N_13609);
nor U17321 (N_17321,N_12483,N_13059);
nor U17322 (N_17322,N_13354,N_12174);
nor U17323 (N_17323,N_12513,N_12437);
and U17324 (N_17324,N_12217,N_11943);
nor U17325 (N_17325,N_13901,N_14623);
nand U17326 (N_17326,N_10966,N_13111);
and U17327 (N_17327,N_10014,N_12612);
or U17328 (N_17328,N_14876,N_12849);
and U17329 (N_17329,N_11375,N_13056);
and U17330 (N_17330,N_14263,N_12355);
and U17331 (N_17331,N_14597,N_13450);
or U17332 (N_17332,N_12286,N_13017);
nor U17333 (N_17333,N_12809,N_13913);
or U17334 (N_17334,N_12051,N_11268);
or U17335 (N_17335,N_11432,N_11414);
nand U17336 (N_17336,N_12687,N_10940);
xnor U17337 (N_17337,N_13207,N_14294);
nor U17338 (N_17338,N_12106,N_12245);
or U17339 (N_17339,N_13536,N_11731);
xor U17340 (N_17340,N_14729,N_13465);
nand U17341 (N_17341,N_12519,N_10878);
nand U17342 (N_17342,N_14331,N_12787);
xor U17343 (N_17343,N_11133,N_13833);
or U17344 (N_17344,N_11957,N_14557);
or U17345 (N_17345,N_11591,N_11490);
and U17346 (N_17346,N_12892,N_11203);
nor U17347 (N_17347,N_12449,N_13453);
xor U17348 (N_17348,N_10922,N_12750);
and U17349 (N_17349,N_12987,N_14826);
or U17350 (N_17350,N_10936,N_12089);
nand U17351 (N_17351,N_10787,N_11255);
nor U17352 (N_17352,N_10072,N_11146);
or U17353 (N_17353,N_10881,N_12736);
nor U17354 (N_17354,N_14515,N_10447);
nand U17355 (N_17355,N_13826,N_12899);
nor U17356 (N_17356,N_14563,N_14543);
nand U17357 (N_17357,N_14166,N_13495);
and U17358 (N_17358,N_14065,N_14121);
and U17359 (N_17359,N_14943,N_12033);
xnor U17360 (N_17360,N_12177,N_11602);
nand U17361 (N_17361,N_12888,N_11486);
nand U17362 (N_17362,N_10566,N_13166);
or U17363 (N_17363,N_12690,N_11168);
and U17364 (N_17364,N_11861,N_11590);
or U17365 (N_17365,N_10504,N_14795);
or U17366 (N_17366,N_11821,N_10939);
nand U17367 (N_17367,N_11305,N_12619);
or U17368 (N_17368,N_13669,N_13388);
nor U17369 (N_17369,N_13142,N_13485);
nor U17370 (N_17370,N_13101,N_12627);
nor U17371 (N_17371,N_11840,N_12599);
nand U17372 (N_17372,N_11324,N_12386);
nor U17373 (N_17373,N_12125,N_14258);
and U17374 (N_17374,N_11512,N_13998);
xnor U17375 (N_17375,N_14594,N_11820);
xor U17376 (N_17376,N_14535,N_13780);
nand U17377 (N_17377,N_14155,N_12249);
nand U17378 (N_17378,N_10348,N_12288);
and U17379 (N_17379,N_10241,N_11961);
nor U17380 (N_17380,N_13023,N_14756);
or U17381 (N_17381,N_12754,N_11951);
and U17382 (N_17382,N_12122,N_12148);
xor U17383 (N_17383,N_14640,N_11500);
xor U17384 (N_17384,N_14786,N_12403);
nand U17385 (N_17385,N_13241,N_14250);
nor U17386 (N_17386,N_14024,N_14115);
or U17387 (N_17387,N_11499,N_10621);
or U17388 (N_17388,N_10587,N_10337);
xor U17389 (N_17389,N_12756,N_11178);
and U17390 (N_17390,N_13875,N_12782);
and U17391 (N_17391,N_12478,N_12709);
nor U17392 (N_17392,N_10414,N_10489);
xnor U17393 (N_17393,N_11919,N_12714);
nand U17394 (N_17394,N_12398,N_12473);
xor U17395 (N_17395,N_12381,N_14008);
xnor U17396 (N_17396,N_11140,N_13089);
and U17397 (N_17397,N_11443,N_13185);
nand U17398 (N_17398,N_12348,N_14968);
xor U17399 (N_17399,N_13570,N_12412);
nand U17400 (N_17400,N_12665,N_10889);
nand U17401 (N_17401,N_11678,N_13814);
nor U17402 (N_17402,N_12856,N_13857);
or U17403 (N_17403,N_12184,N_10506);
or U17404 (N_17404,N_12257,N_11759);
xor U17405 (N_17405,N_13884,N_10540);
or U17406 (N_17406,N_12954,N_13845);
or U17407 (N_17407,N_14914,N_14855);
and U17408 (N_17408,N_11664,N_10802);
or U17409 (N_17409,N_13387,N_10818);
and U17410 (N_17410,N_11828,N_10458);
nand U17411 (N_17411,N_13384,N_12630);
or U17412 (N_17412,N_10228,N_12514);
nor U17413 (N_17413,N_11361,N_10578);
xor U17414 (N_17414,N_14715,N_14750);
nor U17415 (N_17415,N_10923,N_11478);
or U17416 (N_17416,N_14079,N_10828);
nand U17417 (N_17417,N_13503,N_14430);
xor U17418 (N_17418,N_12237,N_11078);
and U17419 (N_17419,N_10102,N_10187);
nand U17420 (N_17420,N_12347,N_12100);
and U17421 (N_17421,N_10534,N_11997);
xor U17422 (N_17422,N_14818,N_14696);
xnor U17423 (N_17423,N_12163,N_14157);
or U17424 (N_17424,N_12542,N_10112);
nand U17425 (N_17425,N_12922,N_13175);
xor U17426 (N_17426,N_13048,N_14971);
and U17427 (N_17427,N_12220,N_11272);
nor U17428 (N_17428,N_13188,N_12947);
nand U17429 (N_17429,N_12047,N_14383);
nor U17430 (N_17430,N_11568,N_10515);
nor U17431 (N_17431,N_10741,N_10360);
xnor U17432 (N_17432,N_14555,N_11246);
xor U17433 (N_17433,N_13580,N_10971);
nand U17434 (N_17434,N_14096,N_13825);
xor U17435 (N_17435,N_12971,N_14218);
nor U17436 (N_17436,N_11070,N_12308);
nor U17437 (N_17437,N_11569,N_10807);
and U17438 (N_17438,N_13433,N_12834);
or U17439 (N_17439,N_11920,N_10542);
and U17440 (N_17440,N_11749,N_14748);
and U17441 (N_17441,N_14585,N_12479);
xnor U17442 (N_17442,N_10366,N_13141);
nor U17443 (N_17443,N_12195,N_10444);
or U17444 (N_17444,N_12762,N_14086);
and U17445 (N_17445,N_11410,N_10551);
xnor U17446 (N_17446,N_14214,N_14851);
nor U17447 (N_17447,N_10857,N_10375);
or U17448 (N_17448,N_14992,N_10772);
nor U17449 (N_17449,N_14616,N_12156);
nor U17450 (N_17450,N_11580,N_12835);
and U17451 (N_17451,N_11533,N_10236);
and U17452 (N_17452,N_11855,N_12608);
nand U17453 (N_17453,N_14969,N_14590);
nand U17454 (N_17454,N_11326,N_13346);
or U17455 (N_17455,N_13987,N_11799);
and U17456 (N_17456,N_11757,N_13819);
nand U17457 (N_17457,N_12757,N_12898);
or U17458 (N_17458,N_13292,N_12562);
nor U17459 (N_17459,N_14248,N_10934);
xor U17460 (N_17460,N_10752,N_10017);
and U17461 (N_17461,N_11357,N_11415);
and U17462 (N_17462,N_11173,N_10777);
and U17463 (N_17463,N_11122,N_14859);
and U17464 (N_17464,N_13785,N_14469);
or U17465 (N_17465,N_13372,N_10959);
nor U17466 (N_17466,N_11937,N_13368);
and U17467 (N_17467,N_14393,N_13275);
and U17468 (N_17468,N_10632,N_12494);
nor U17469 (N_17469,N_11359,N_12463);
nand U17470 (N_17470,N_14527,N_10759);
and U17471 (N_17471,N_12957,N_14154);
xnor U17472 (N_17472,N_10486,N_12916);
nor U17473 (N_17473,N_13158,N_13199);
and U17474 (N_17474,N_11878,N_10196);
xnor U17475 (N_17475,N_12256,N_12194);
or U17476 (N_17476,N_13196,N_10098);
or U17477 (N_17477,N_12507,N_12647);
xnor U17478 (N_17478,N_10748,N_11583);
xnor U17479 (N_17479,N_11839,N_11782);
nor U17480 (N_17480,N_11708,N_14273);
or U17481 (N_17481,N_11439,N_10466);
and U17482 (N_17482,N_11800,N_12554);
nand U17483 (N_17483,N_13413,N_14435);
nor U17484 (N_17484,N_12103,N_13980);
nand U17485 (N_17485,N_12364,N_12396);
nor U17486 (N_17486,N_12354,N_11675);
nor U17487 (N_17487,N_13191,N_12915);
or U17488 (N_17488,N_12909,N_10055);
or U17489 (N_17489,N_14088,N_11693);
xnor U17490 (N_17490,N_11354,N_11096);
nand U17491 (N_17491,N_12908,N_12594);
and U17492 (N_17492,N_14975,N_14745);
xnor U17493 (N_17493,N_12202,N_11156);
or U17494 (N_17494,N_14309,N_14799);
nand U17495 (N_17495,N_14438,N_12445);
xnor U17496 (N_17496,N_14996,N_10921);
xor U17497 (N_17497,N_11016,N_14459);
nand U17498 (N_17498,N_11014,N_11371);
or U17499 (N_17499,N_13404,N_10609);
and U17500 (N_17500,N_13380,N_11477);
nor U17501 (N_17501,N_10148,N_13660);
nand U17502 (N_17502,N_13025,N_10139);
and U17503 (N_17503,N_11160,N_13704);
or U17504 (N_17504,N_12975,N_14061);
and U17505 (N_17505,N_11175,N_11858);
nand U17506 (N_17506,N_13448,N_11767);
nand U17507 (N_17507,N_14270,N_13386);
nor U17508 (N_17508,N_11077,N_10673);
and U17509 (N_17509,N_12903,N_10481);
and U17510 (N_17510,N_11789,N_12557);
nor U17511 (N_17511,N_13973,N_14939);
xnor U17512 (N_17512,N_13760,N_12345);
nand U17513 (N_17513,N_11420,N_14451);
xor U17514 (N_17514,N_11501,N_11178);
and U17515 (N_17515,N_12352,N_14723);
and U17516 (N_17516,N_13299,N_13315);
nor U17517 (N_17517,N_13871,N_11956);
nand U17518 (N_17518,N_13092,N_11625);
nor U17519 (N_17519,N_14222,N_13802);
nand U17520 (N_17520,N_11006,N_11009);
or U17521 (N_17521,N_14127,N_10298);
xor U17522 (N_17522,N_12765,N_10726);
nor U17523 (N_17523,N_12289,N_10230);
and U17524 (N_17524,N_13141,N_12301);
xor U17525 (N_17525,N_12801,N_14023);
and U17526 (N_17526,N_14411,N_13571);
nor U17527 (N_17527,N_10915,N_12624);
or U17528 (N_17528,N_11759,N_13295);
or U17529 (N_17529,N_13999,N_11050);
xor U17530 (N_17530,N_10994,N_13668);
and U17531 (N_17531,N_12690,N_10718);
or U17532 (N_17532,N_10247,N_14902);
nor U17533 (N_17533,N_12514,N_14912);
or U17534 (N_17534,N_11002,N_12785);
nand U17535 (N_17535,N_14778,N_12010);
nor U17536 (N_17536,N_14358,N_14804);
nand U17537 (N_17537,N_10703,N_10088);
xnor U17538 (N_17538,N_14794,N_10938);
and U17539 (N_17539,N_10063,N_11818);
xnor U17540 (N_17540,N_11236,N_14259);
xnor U17541 (N_17541,N_13907,N_13897);
nand U17542 (N_17542,N_14392,N_10550);
or U17543 (N_17543,N_14084,N_11956);
and U17544 (N_17544,N_13824,N_12374);
xor U17545 (N_17545,N_10818,N_11100);
or U17546 (N_17546,N_12161,N_11081);
nor U17547 (N_17547,N_14241,N_12436);
or U17548 (N_17548,N_13446,N_12021);
nor U17549 (N_17549,N_12421,N_10622);
or U17550 (N_17550,N_11366,N_13532);
nor U17551 (N_17551,N_12308,N_12204);
or U17552 (N_17552,N_11965,N_12841);
xnor U17553 (N_17553,N_14739,N_12285);
or U17554 (N_17554,N_11771,N_14024);
or U17555 (N_17555,N_12994,N_11117);
xor U17556 (N_17556,N_11683,N_11819);
and U17557 (N_17557,N_11143,N_14773);
nor U17558 (N_17558,N_12260,N_14906);
xor U17559 (N_17559,N_12801,N_10223);
nand U17560 (N_17560,N_14231,N_14475);
nand U17561 (N_17561,N_10992,N_13108);
nor U17562 (N_17562,N_10800,N_11402);
nor U17563 (N_17563,N_14716,N_14045);
xnor U17564 (N_17564,N_12896,N_11807);
and U17565 (N_17565,N_10098,N_13404);
nand U17566 (N_17566,N_14355,N_10940);
nor U17567 (N_17567,N_14354,N_11783);
nand U17568 (N_17568,N_13555,N_14597);
nor U17569 (N_17569,N_11102,N_11033);
nor U17570 (N_17570,N_11316,N_10517);
and U17571 (N_17571,N_10034,N_12885);
nor U17572 (N_17572,N_13617,N_14423);
nor U17573 (N_17573,N_12914,N_10418);
and U17574 (N_17574,N_13370,N_14992);
and U17575 (N_17575,N_14822,N_14430);
xnor U17576 (N_17576,N_11891,N_14004);
xnor U17577 (N_17577,N_11900,N_12916);
nand U17578 (N_17578,N_10400,N_11692);
and U17579 (N_17579,N_10396,N_14624);
and U17580 (N_17580,N_13784,N_12270);
nor U17581 (N_17581,N_14939,N_11203);
nand U17582 (N_17582,N_11531,N_10836);
nand U17583 (N_17583,N_13957,N_11403);
and U17584 (N_17584,N_12806,N_11003);
xor U17585 (N_17585,N_13013,N_10357);
nand U17586 (N_17586,N_12811,N_10080);
or U17587 (N_17587,N_13498,N_12856);
and U17588 (N_17588,N_13072,N_13046);
nand U17589 (N_17589,N_11549,N_12928);
xor U17590 (N_17590,N_12820,N_13907);
xnor U17591 (N_17591,N_11700,N_10804);
nand U17592 (N_17592,N_12756,N_10274);
nand U17593 (N_17593,N_12461,N_12897);
xnor U17594 (N_17594,N_10644,N_10180);
nand U17595 (N_17595,N_13442,N_10186);
xnor U17596 (N_17596,N_11252,N_11590);
or U17597 (N_17597,N_13998,N_10646);
and U17598 (N_17598,N_12217,N_13303);
and U17599 (N_17599,N_12806,N_13476);
nand U17600 (N_17600,N_13319,N_13823);
or U17601 (N_17601,N_12410,N_10697);
nand U17602 (N_17602,N_13563,N_14264);
nor U17603 (N_17603,N_14204,N_13679);
and U17604 (N_17604,N_13639,N_10505);
or U17605 (N_17605,N_10758,N_13504);
xnor U17606 (N_17606,N_14658,N_14141);
and U17607 (N_17607,N_12796,N_13099);
or U17608 (N_17608,N_12578,N_13165);
xnor U17609 (N_17609,N_10016,N_13042);
nor U17610 (N_17610,N_10946,N_11114);
xnor U17611 (N_17611,N_13750,N_12353);
nand U17612 (N_17612,N_10180,N_13884);
xnor U17613 (N_17613,N_10895,N_11593);
and U17614 (N_17614,N_10033,N_14804);
nand U17615 (N_17615,N_14795,N_12000);
xnor U17616 (N_17616,N_14588,N_11454);
nor U17617 (N_17617,N_10629,N_14974);
nor U17618 (N_17618,N_10384,N_14158);
nor U17619 (N_17619,N_13924,N_11232);
nand U17620 (N_17620,N_13769,N_14970);
nor U17621 (N_17621,N_14232,N_10193);
xnor U17622 (N_17622,N_10566,N_13383);
nor U17623 (N_17623,N_12869,N_14658);
xor U17624 (N_17624,N_10392,N_14099);
nor U17625 (N_17625,N_11747,N_10684);
or U17626 (N_17626,N_11243,N_14111);
nor U17627 (N_17627,N_11639,N_14814);
nand U17628 (N_17628,N_11681,N_11262);
or U17629 (N_17629,N_14944,N_14233);
and U17630 (N_17630,N_11810,N_13835);
xor U17631 (N_17631,N_13158,N_13284);
nor U17632 (N_17632,N_11391,N_14948);
nor U17633 (N_17633,N_10088,N_12397);
nand U17634 (N_17634,N_10201,N_13939);
nand U17635 (N_17635,N_12966,N_14866);
xor U17636 (N_17636,N_11536,N_14367);
nand U17637 (N_17637,N_12210,N_14856);
xor U17638 (N_17638,N_12863,N_10521);
or U17639 (N_17639,N_11523,N_14683);
nor U17640 (N_17640,N_13581,N_12042);
or U17641 (N_17641,N_14883,N_14230);
xor U17642 (N_17642,N_12270,N_11414);
nand U17643 (N_17643,N_10890,N_13880);
xor U17644 (N_17644,N_10223,N_13100);
nand U17645 (N_17645,N_12368,N_10236);
or U17646 (N_17646,N_13129,N_14362);
nor U17647 (N_17647,N_13476,N_13417);
nor U17648 (N_17648,N_10353,N_10882);
or U17649 (N_17649,N_13134,N_13616);
xor U17650 (N_17650,N_14409,N_13483);
xnor U17651 (N_17651,N_14679,N_13763);
nand U17652 (N_17652,N_13338,N_14917);
and U17653 (N_17653,N_10040,N_11605);
and U17654 (N_17654,N_14608,N_14681);
xor U17655 (N_17655,N_11419,N_11798);
nor U17656 (N_17656,N_10321,N_12661);
and U17657 (N_17657,N_11739,N_10871);
or U17658 (N_17658,N_11611,N_10470);
nand U17659 (N_17659,N_12666,N_14731);
nor U17660 (N_17660,N_14101,N_10979);
or U17661 (N_17661,N_14495,N_13200);
nor U17662 (N_17662,N_13483,N_12851);
xnor U17663 (N_17663,N_12566,N_12662);
xor U17664 (N_17664,N_13907,N_10016);
nor U17665 (N_17665,N_10040,N_14000);
or U17666 (N_17666,N_10910,N_12675);
xnor U17667 (N_17667,N_10146,N_10219);
or U17668 (N_17668,N_12392,N_10294);
xnor U17669 (N_17669,N_14132,N_12006);
xnor U17670 (N_17670,N_13424,N_12338);
or U17671 (N_17671,N_11206,N_13590);
xnor U17672 (N_17672,N_11835,N_14556);
nand U17673 (N_17673,N_13222,N_10113);
or U17674 (N_17674,N_11482,N_10417);
nor U17675 (N_17675,N_12643,N_14282);
or U17676 (N_17676,N_14481,N_13449);
nor U17677 (N_17677,N_10150,N_13069);
or U17678 (N_17678,N_13102,N_10206);
xnor U17679 (N_17679,N_11384,N_14538);
nor U17680 (N_17680,N_13581,N_14519);
or U17681 (N_17681,N_12749,N_11692);
or U17682 (N_17682,N_10140,N_12798);
nor U17683 (N_17683,N_13075,N_10111);
nand U17684 (N_17684,N_13188,N_11357);
and U17685 (N_17685,N_12165,N_10928);
nor U17686 (N_17686,N_12574,N_12834);
xnor U17687 (N_17687,N_13665,N_14897);
nor U17688 (N_17688,N_14428,N_13147);
or U17689 (N_17689,N_10828,N_13616);
or U17690 (N_17690,N_10462,N_14437);
nand U17691 (N_17691,N_11244,N_10322);
or U17692 (N_17692,N_13721,N_12046);
nand U17693 (N_17693,N_14956,N_12378);
nand U17694 (N_17694,N_12192,N_13139);
xnor U17695 (N_17695,N_11721,N_14007);
xnor U17696 (N_17696,N_11874,N_14898);
xnor U17697 (N_17697,N_14965,N_11838);
and U17698 (N_17698,N_11464,N_11189);
xnor U17699 (N_17699,N_13652,N_14731);
xor U17700 (N_17700,N_13706,N_10904);
or U17701 (N_17701,N_10487,N_11314);
and U17702 (N_17702,N_12149,N_12871);
and U17703 (N_17703,N_14502,N_13183);
nand U17704 (N_17704,N_13050,N_14702);
nor U17705 (N_17705,N_11463,N_14719);
xnor U17706 (N_17706,N_10887,N_12612);
or U17707 (N_17707,N_11223,N_12764);
nand U17708 (N_17708,N_13534,N_10217);
or U17709 (N_17709,N_13114,N_14577);
nand U17710 (N_17710,N_12807,N_13676);
or U17711 (N_17711,N_12309,N_10343);
or U17712 (N_17712,N_14943,N_11774);
nand U17713 (N_17713,N_12482,N_14177);
or U17714 (N_17714,N_11950,N_11824);
nand U17715 (N_17715,N_14454,N_10906);
nand U17716 (N_17716,N_11976,N_10950);
xnor U17717 (N_17717,N_14114,N_13605);
nand U17718 (N_17718,N_13111,N_13652);
xor U17719 (N_17719,N_11492,N_10844);
or U17720 (N_17720,N_14491,N_10875);
nor U17721 (N_17721,N_10311,N_14749);
xor U17722 (N_17722,N_11378,N_14957);
or U17723 (N_17723,N_11565,N_13667);
nor U17724 (N_17724,N_13550,N_11378);
nor U17725 (N_17725,N_10751,N_12374);
xnor U17726 (N_17726,N_13796,N_13934);
xor U17727 (N_17727,N_14314,N_10686);
xnor U17728 (N_17728,N_12043,N_11012);
xnor U17729 (N_17729,N_14249,N_12498);
nand U17730 (N_17730,N_14505,N_12591);
or U17731 (N_17731,N_13903,N_13731);
or U17732 (N_17732,N_12626,N_11726);
and U17733 (N_17733,N_12151,N_14975);
xnor U17734 (N_17734,N_11546,N_11943);
xor U17735 (N_17735,N_10673,N_10572);
nand U17736 (N_17736,N_14111,N_13308);
and U17737 (N_17737,N_10324,N_13059);
or U17738 (N_17738,N_12516,N_10634);
nand U17739 (N_17739,N_14153,N_11385);
or U17740 (N_17740,N_11782,N_12596);
nor U17741 (N_17741,N_14909,N_14544);
nor U17742 (N_17742,N_14755,N_13472);
or U17743 (N_17743,N_11533,N_11339);
nor U17744 (N_17744,N_14695,N_12947);
xnor U17745 (N_17745,N_11680,N_13980);
or U17746 (N_17746,N_10900,N_10520);
xor U17747 (N_17747,N_12219,N_12552);
or U17748 (N_17748,N_10185,N_12105);
nand U17749 (N_17749,N_10990,N_12739);
nor U17750 (N_17750,N_12088,N_11635);
nand U17751 (N_17751,N_14676,N_11052);
xor U17752 (N_17752,N_10365,N_12231);
xnor U17753 (N_17753,N_10636,N_14825);
xor U17754 (N_17754,N_13989,N_12392);
or U17755 (N_17755,N_13709,N_11256);
nor U17756 (N_17756,N_13642,N_14215);
and U17757 (N_17757,N_13559,N_14083);
or U17758 (N_17758,N_12151,N_13515);
xor U17759 (N_17759,N_13368,N_12462);
or U17760 (N_17760,N_11705,N_12357);
xor U17761 (N_17761,N_11750,N_12760);
nor U17762 (N_17762,N_12059,N_13425);
nand U17763 (N_17763,N_12551,N_11806);
or U17764 (N_17764,N_12468,N_10959);
and U17765 (N_17765,N_11535,N_10948);
xnor U17766 (N_17766,N_12902,N_12408);
nor U17767 (N_17767,N_14718,N_10660);
or U17768 (N_17768,N_14907,N_12439);
and U17769 (N_17769,N_10007,N_10573);
nand U17770 (N_17770,N_13845,N_12200);
nor U17771 (N_17771,N_11485,N_14148);
nand U17772 (N_17772,N_10306,N_12031);
nor U17773 (N_17773,N_14389,N_11982);
and U17774 (N_17774,N_13445,N_12959);
and U17775 (N_17775,N_12525,N_11282);
xor U17776 (N_17776,N_14369,N_10291);
xnor U17777 (N_17777,N_10449,N_14318);
or U17778 (N_17778,N_11963,N_14910);
nor U17779 (N_17779,N_11203,N_12176);
or U17780 (N_17780,N_13601,N_12425);
nand U17781 (N_17781,N_10852,N_14278);
nand U17782 (N_17782,N_13132,N_14558);
and U17783 (N_17783,N_10427,N_12846);
and U17784 (N_17784,N_11579,N_10857);
xnor U17785 (N_17785,N_14118,N_13915);
and U17786 (N_17786,N_10297,N_10805);
or U17787 (N_17787,N_13044,N_11095);
or U17788 (N_17788,N_14179,N_11768);
nand U17789 (N_17789,N_10867,N_11679);
xor U17790 (N_17790,N_10386,N_14980);
nand U17791 (N_17791,N_11971,N_14096);
nand U17792 (N_17792,N_13357,N_14374);
xor U17793 (N_17793,N_10428,N_13013);
or U17794 (N_17794,N_12316,N_11064);
or U17795 (N_17795,N_12312,N_13870);
nor U17796 (N_17796,N_11680,N_14267);
nor U17797 (N_17797,N_10602,N_10834);
xnor U17798 (N_17798,N_12998,N_10428);
xnor U17799 (N_17799,N_13341,N_11861);
xor U17800 (N_17800,N_12974,N_12435);
and U17801 (N_17801,N_12827,N_12524);
xnor U17802 (N_17802,N_10845,N_14114);
and U17803 (N_17803,N_12694,N_13120);
or U17804 (N_17804,N_11662,N_14504);
and U17805 (N_17805,N_12443,N_13482);
nand U17806 (N_17806,N_13931,N_10104);
and U17807 (N_17807,N_14404,N_11501);
or U17808 (N_17808,N_13498,N_11856);
and U17809 (N_17809,N_11011,N_14940);
nor U17810 (N_17810,N_12178,N_10485);
xnor U17811 (N_17811,N_11583,N_10660);
nor U17812 (N_17812,N_11639,N_13473);
nor U17813 (N_17813,N_12426,N_13393);
xnor U17814 (N_17814,N_14957,N_12850);
nor U17815 (N_17815,N_11261,N_14107);
xnor U17816 (N_17816,N_13474,N_13581);
nor U17817 (N_17817,N_10396,N_10966);
nand U17818 (N_17818,N_11828,N_12661);
nand U17819 (N_17819,N_10620,N_14607);
xor U17820 (N_17820,N_13357,N_14613);
xnor U17821 (N_17821,N_11207,N_13765);
xnor U17822 (N_17822,N_13575,N_12202);
and U17823 (N_17823,N_13590,N_11592);
nor U17824 (N_17824,N_14332,N_10099);
nand U17825 (N_17825,N_10255,N_11338);
and U17826 (N_17826,N_14893,N_14210);
or U17827 (N_17827,N_10227,N_11682);
and U17828 (N_17828,N_14146,N_11673);
xnor U17829 (N_17829,N_13813,N_14340);
and U17830 (N_17830,N_11527,N_14485);
and U17831 (N_17831,N_12027,N_13877);
and U17832 (N_17832,N_11841,N_12708);
nand U17833 (N_17833,N_14898,N_12873);
and U17834 (N_17834,N_12225,N_13155);
and U17835 (N_17835,N_13651,N_10506);
or U17836 (N_17836,N_12718,N_14613);
or U17837 (N_17837,N_10618,N_11821);
nand U17838 (N_17838,N_12430,N_14345);
and U17839 (N_17839,N_13911,N_13456);
xnor U17840 (N_17840,N_14545,N_10040);
or U17841 (N_17841,N_10610,N_10689);
nand U17842 (N_17842,N_11299,N_11720);
nor U17843 (N_17843,N_10423,N_12067);
and U17844 (N_17844,N_14920,N_14634);
or U17845 (N_17845,N_12546,N_11811);
and U17846 (N_17846,N_10193,N_12145);
xnor U17847 (N_17847,N_12050,N_10439);
nand U17848 (N_17848,N_14679,N_11269);
or U17849 (N_17849,N_12549,N_11199);
nor U17850 (N_17850,N_11962,N_12420);
xnor U17851 (N_17851,N_12771,N_12035);
nor U17852 (N_17852,N_13868,N_14766);
nor U17853 (N_17853,N_14048,N_14901);
nor U17854 (N_17854,N_10115,N_13317);
xor U17855 (N_17855,N_12704,N_13013);
xnor U17856 (N_17856,N_11849,N_10138);
nand U17857 (N_17857,N_13790,N_12031);
and U17858 (N_17858,N_14748,N_12641);
or U17859 (N_17859,N_13724,N_13508);
and U17860 (N_17860,N_12101,N_11946);
or U17861 (N_17861,N_10918,N_13734);
and U17862 (N_17862,N_11147,N_10146);
or U17863 (N_17863,N_13212,N_10483);
and U17864 (N_17864,N_13345,N_10199);
xnor U17865 (N_17865,N_13851,N_14057);
nor U17866 (N_17866,N_12286,N_13743);
nand U17867 (N_17867,N_12427,N_14443);
xor U17868 (N_17868,N_10585,N_12017);
nor U17869 (N_17869,N_14740,N_11453);
and U17870 (N_17870,N_12076,N_12214);
nor U17871 (N_17871,N_11385,N_14201);
nor U17872 (N_17872,N_13134,N_12260);
and U17873 (N_17873,N_13991,N_11395);
xor U17874 (N_17874,N_11449,N_13416);
nand U17875 (N_17875,N_13668,N_13661);
and U17876 (N_17876,N_10088,N_12738);
nand U17877 (N_17877,N_12854,N_14581);
xnor U17878 (N_17878,N_10358,N_10975);
or U17879 (N_17879,N_14936,N_11746);
and U17880 (N_17880,N_13542,N_10711);
xnor U17881 (N_17881,N_12326,N_14250);
or U17882 (N_17882,N_13576,N_13990);
and U17883 (N_17883,N_10877,N_14588);
nor U17884 (N_17884,N_10862,N_14420);
xor U17885 (N_17885,N_11442,N_14571);
nor U17886 (N_17886,N_13932,N_12432);
xor U17887 (N_17887,N_13316,N_11731);
nor U17888 (N_17888,N_12300,N_12445);
nand U17889 (N_17889,N_12747,N_12725);
nor U17890 (N_17890,N_13041,N_11185);
xor U17891 (N_17891,N_10192,N_14327);
nand U17892 (N_17892,N_13092,N_14240);
or U17893 (N_17893,N_10670,N_13670);
nand U17894 (N_17894,N_12309,N_11945);
xor U17895 (N_17895,N_11763,N_10672);
or U17896 (N_17896,N_14347,N_14129);
and U17897 (N_17897,N_12909,N_14703);
xor U17898 (N_17898,N_12724,N_10183);
xor U17899 (N_17899,N_12230,N_10035);
nor U17900 (N_17900,N_14977,N_12596);
or U17901 (N_17901,N_10069,N_14728);
xnor U17902 (N_17902,N_10596,N_13190);
nor U17903 (N_17903,N_13323,N_10570);
and U17904 (N_17904,N_11848,N_14594);
xor U17905 (N_17905,N_13362,N_10272);
nor U17906 (N_17906,N_14119,N_13498);
nor U17907 (N_17907,N_13630,N_10145);
nor U17908 (N_17908,N_14148,N_13731);
nand U17909 (N_17909,N_11070,N_14363);
xor U17910 (N_17910,N_12588,N_12772);
nor U17911 (N_17911,N_10128,N_14972);
and U17912 (N_17912,N_12410,N_13825);
nand U17913 (N_17913,N_13700,N_10470);
or U17914 (N_17914,N_13611,N_14279);
and U17915 (N_17915,N_13072,N_11262);
nor U17916 (N_17916,N_13868,N_14426);
or U17917 (N_17917,N_11562,N_14276);
xnor U17918 (N_17918,N_10558,N_11910);
nor U17919 (N_17919,N_14057,N_13323);
xor U17920 (N_17920,N_12632,N_13857);
and U17921 (N_17921,N_13878,N_12273);
nand U17922 (N_17922,N_14820,N_13387);
nand U17923 (N_17923,N_10828,N_12902);
and U17924 (N_17924,N_14393,N_10082);
or U17925 (N_17925,N_12528,N_13923);
xor U17926 (N_17926,N_10851,N_12812);
nor U17927 (N_17927,N_12573,N_12148);
and U17928 (N_17928,N_11541,N_11648);
nor U17929 (N_17929,N_12027,N_10313);
and U17930 (N_17930,N_10133,N_14185);
nor U17931 (N_17931,N_13070,N_11213);
nand U17932 (N_17932,N_10142,N_11051);
or U17933 (N_17933,N_10857,N_13638);
nor U17934 (N_17934,N_12609,N_10598);
xnor U17935 (N_17935,N_12694,N_14768);
and U17936 (N_17936,N_11055,N_13741);
nand U17937 (N_17937,N_14927,N_10800);
xnor U17938 (N_17938,N_14007,N_10513);
and U17939 (N_17939,N_10646,N_12754);
nand U17940 (N_17940,N_11524,N_10405);
and U17941 (N_17941,N_11125,N_13739);
nor U17942 (N_17942,N_11513,N_12427);
nor U17943 (N_17943,N_13158,N_11153);
or U17944 (N_17944,N_11710,N_14489);
nand U17945 (N_17945,N_14459,N_10081);
xnor U17946 (N_17946,N_11092,N_14890);
nand U17947 (N_17947,N_12629,N_14304);
nand U17948 (N_17948,N_13743,N_14571);
and U17949 (N_17949,N_10994,N_14746);
or U17950 (N_17950,N_12699,N_11221);
nor U17951 (N_17951,N_10546,N_11593);
xor U17952 (N_17952,N_12289,N_11608);
nand U17953 (N_17953,N_14479,N_12516);
or U17954 (N_17954,N_14002,N_11498);
or U17955 (N_17955,N_14696,N_14647);
nor U17956 (N_17956,N_13083,N_14324);
nor U17957 (N_17957,N_11692,N_14167);
nand U17958 (N_17958,N_12887,N_13261);
nor U17959 (N_17959,N_12986,N_14449);
or U17960 (N_17960,N_10259,N_12733);
or U17961 (N_17961,N_10931,N_13151);
and U17962 (N_17962,N_14585,N_10164);
xor U17963 (N_17963,N_11768,N_13152);
or U17964 (N_17964,N_12430,N_11036);
and U17965 (N_17965,N_14926,N_14909);
xor U17966 (N_17966,N_14929,N_11318);
or U17967 (N_17967,N_12558,N_13824);
or U17968 (N_17968,N_10827,N_11146);
nand U17969 (N_17969,N_12248,N_10476);
and U17970 (N_17970,N_11661,N_11943);
nand U17971 (N_17971,N_11968,N_10129);
nor U17972 (N_17972,N_10588,N_11831);
nand U17973 (N_17973,N_13875,N_14117);
or U17974 (N_17974,N_12114,N_14074);
nand U17975 (N_17975,N_13142,N_13541);
xnor U17976 (N_17976,N_13585,N_10808);
or U17977 (N_17977,N_11816,N_14458);
xor U17978 (N_17978,N_11069,N_10089);
or U17979 (N_17979,N_10433,N_14232);
nor U17980 (N_17980,N_14939,N_14875);
nor U17981 (N_17981,N_14422,N_10946);
nand U17982 (N_17982,N_11078,N_10149);
nor U17983 (N_17983,N_14426,N_10941);
nor U17984 (N_17984,N_12455,N_14149);
xor U17985 (N_17985,N_13335,N_12231);
or U17986 (N_17986,N_14560,N_11685);
and U17987 (N_17987,N_10562,N_11165);
or U17988 (N_17988,N_11297,N_12080);
nor U17989 (N_17989,N_14887,N_12481);
nor U17990 (N_17990,N_12841,N_11399);
nor U17991 (N_17991,N_12233,N_13489);
nor U17992 (N_17992,N_12841,N_11975);
or U17993 (N_17993,N_11138,N_14354);
or U17994 (N_17994,N_11304,N_10673);
or U17995 (N_17995,N_13846,N_10534);
or U17996 (N_17996,N_14547,N_12109);
or U17997 (N_17997,N_13914,N_14447);
xor U17998 (N_17998,N_11714,N_11334);
nor U17999 (N_17999,N_12254,N_11583);
xnor U18000 (N_18000,N_12005,N_14037);
xnor U18001 (N_18001,N_10366,N_13904);
and U18002 (N_18002,N_10775,N_12281);
or U18003 (N_18003,N_11995,N_11387);
nand U18004 (N_18004,N_10975,N_10256);
xor U18005 (N_18005,N_11307,N_11577);
nor U18006 (N_18006,N_11678,N_14837);
and U18007 (N_18007,N_10529,N_10526);
nand U18008 (N_18008,N_11045,N_11963);
or U18009 (N_18009,N_12317,N_10562);
nand U18010 (N_18010,N_12794,N_12796);
and U18011 (N_18011,N_14247,N_10474);
xnor U18012 (N_18012,N_12728,N_13852);
or U18013 (N_18013,N_13900,N_14154);
nor U18014 (N_18014,N_14026,N_12398);
or U18015 (N_18015,N_13746,N_12061);
nand U18016 (N_18016,N_10010,N_11718);
or U18017 (N_18017,N_10658,N_11437);
and U18018 (N_18018,N_14095,N_11684);
and U18019 (N_18019,N_13409,N_13018);
nand U18020 (N_18020,N_10203,N_14396);
nand U18021 (N_18021,N_13472,N_14529);
and U18022 (N_18022,N_11133,N_11015);
and U18023 (N_18023,N_12904,N_13028);
and U18024 (N_18024,N_11767,N_10280);
nor U18025 (N_18025,N_10558,N_11567);
or U18026 (N_18026,N_10336,N_14757);
nand U18027 (N_18027,N_11268,N_10017);
nand U18028 (N_18028,N_13228,N_11968);
xor U18029 (N_18029,N_13781,N_10977);
xor U18030 (N_18030,N_12453,N_13587);
or U18031 (N_18031,N_10739,N_12686);
nand U18032 (N_18032,N_11315,N_12991);
or U18033 (N_18033,N_11837,N_11458);
or U18034 (N_18034,N_13672,N_13546);
and U18035 (N_18035,N_10227,N_10458);
nor U18036 (N_18036,N_11079,N_13057);
nor U18037 (N_18037,N_13076,N_13571);
xor U18038 (N_18038,N_12449,N_11799);
nor U18039 (N_18039,N_12381,N_11949);
nand U18040 (N_18040,N_12926,N_10816);
xor U18041 (N_18041,N_11742,N_14979);
or U18042 (N_18042,N_13557,N_12724);
nor U18043 (N_18043,N_10092,N_12731);
nor U18044 (N_18044,N_11151,N_13658);
nand U18045 (N_18045,N_13245,N_14640);
xor U18046 (N_18046,N_12256,N_13533);
or U18047 (N_18047,N_12658,N_10338);
xor U18048 (N_18048,N_10512,N_12020);
xnor U18049 (N_18049,N_13296,N_13225);
nor U18050 (N_18050,N_10523,N_10426);
nor U18051 (N_18051,N_13283,N_12678);
and U18052 (N_18052,N_11694,N_11222);
or U18053 (N_18053,N_12999,N_13722);
or U18054 (N_18054,N_12703,N_13077);
and U18055 (N_18055,N_12939,N_11779);
xnor U18056 (N_18056,N_10053,N_14912);
nand U18057 (N_18057,N_14237,N_13764);
nand U18058 (N_18058,N_11725,N_14499);
nor U18059 (N_18059,N_13788,N_11743);
and U18060 (N_18060,N_11163,N_10456);
and U18061 (N_18061,N_10933,N_14996);
nand U18062 (N_18062,N_14883,N_14271);
or U18063 (N_18063,N_10653,N_11070);
or U18064 (N_18064,N_14515,N_12405);
nor U18065 (N_18065,N_10046,N_10327);
nor U18066 (N_18066,N_11440,N_13115);
and U18067 (N_18067,N_12547,N_11994);
or U18068 (N_18068,N_10425,N_10010);
and U18069 (N_18069,N_11089,N_14232);
or U18070 (N_18070,N_10417,N_12752);
xnor U18071 (N_18071,N_11032,N_14231);
nor U18072 (N_18072,N_14070,N_14661);
and U18073 (N_18073,N_13173,N_10149);
nor U18074 (N_18074,N_12198,N_13451);
and U18075 (N_18075,N_12335,N_12730);
or U18076 (N_18076,N_12057,N_14166);
and U18077 (N_18077,N_10261,N_14749);
xor U18078 (N_18078,N_13502,N_11054);
xnor U18079 (N_18079,N_10804,N_12596);
xnor U18080 (N_18080,N_13792,N_11072);
and U18081 (N_18081,N_11665,N_10844);
xor U18082 (N_18082,N_10685,N_10832);
and U18083 (N_18083,N_13852,N_11989);
xnor U18084 (N_18084,N_11841,N_14253);
nand U18085 (N_18085,N_12603,N_14332);
or U18086 (N_18086,N_11657,N_14269);
or U18087 (N_18087,N_14358,N_11648);
and U18088 (N_18088,N_10418,N_14453);
or U18089 (N_18089,N_13492,N_11125);
or U18090 (N_18090,N_12405,N_13539);
or U18091 (N_18091,N_13916,N_12080);
or U18092 (N_18092,N_13277,N_13191);
or U18093 (N_18093,N_13206,N_11757);
and U18094 (N_18094,N_13875,N_13787);
nor U18095 (N_18095,N_14811,N_14609);
or U18096 (N_18096,N_10458,N_11227);
nand U18097 (N_18097,N_12228,N_14074);
xor U18098 (N_18098,N_13977,N_11984);
nor U18099 (N_18099,N_13037,N_11783);
nand U18100 (N_18100,N_11468,N_10895);
and U18101 (N_18101,N_11011,N_12443);
and U18102 (N_18102,N_12848,N_11566);
xor U18103 (N_18103,N_13787,N_13423);
or U18104 (N_18104,N_12182,N_14215);
nand U18105 (N_18105,N_13603,N_10172);
nor U18106 (N_18106,N_11124,N_10385);
and U18107 (N_18107,N_13081,N_13808);
or U18108 (N_18108,N_14333,N_12796);
nor U18109 (N_18109,N_10716,N_10659);
xnor U18110 (N_18110,N_10361,N_14436);
or U18111 (N_18111,N_14826,N_11962);
nor U18112 (N_18112,N_11786,N_12031);
nor U18113 (N_18113,N_14251,N_11661);
nor U18114 (N_18114,N_13080,N_13855);
nor U18115 (N_18115,N_11892,N_14859);
nand U18116 (N_18116,N_10774,N_14373);
and U18117 (N_18117,N_10381,N_11306);
nor U18118 (N_18118,N_12395,N_14244);
xnor U18119 (N_18119,N_13808,N_13912);
or U18120 (N_18120,N_13011,N_14877);
xor U18121 (N_18121,N_11864,N_14610);
nor U18122 (N_18122,N_13698,N_10842);
xnor U18123 (N_18123,N_13928,N_12630);
xnor U18124 (N_18124,N_12550,N_12115);
xor U18125 (N_18125,N_12558,N_10444);
nand U18126 (N_18126,N_12234,N_14507);
and U18127 (N_18127,N_11246,N_10838);
and U18128 (N_18128,N_11941,N_12179);
nor U18129 (N_18129,N_14778,N_11202);
or U18130 (N_18130,N_11204,N_11999);
nor U18131 (N_18131,N_11683,N_12739);
nor U18132 (N_18132,N_11136,N_13200);
and U18133 (N_18133,N_11456,N_13021);
nor U18134 (N_18134,N_12576,N_12785);
xor U18135 (N_18135,N_12203,N_11999);
nand U18136 (N_18136,N_12709,N_14063);
nand U18137 (N_18137,N_12621,N_13604);
and U18138 (N_18138,N_13444,N_12922);
nand U18139 (N_18139,N_11461,N_10483);
xnor U18140 (N_18140,N_13702,N_11383);
and U18141 (N_18141,N_13947,N_12788);
xnor U18142 (N_18142,N_11059,N_10895);
nor U18143 (N_18143,N_14870,N_13130);
or U18144 (N_18144,N_13808,N_13094);
or U18145 (N_18145,N_11411,N_14111);
xnor U18146 (N_18146,N_11372,N_10198);
nand U18147 (N_18147,N_13700,N_10643);
nand U18148 (N_18148,N_12527,N_14022);
and U18149 (N_18149,N_10748,N_10053);
nand U18150 (N_18150,N_13051,N_11902);
nor U18151 (N_18151,N_14178,N_10534);
nand U18152 (N_18152,N_10242,N_11562);
or U18153 (N_18153,N_12251,N_12356);
nor U18154 (N_18154,N_12166,N_11670);
nor U18155 (N_18155,N_11150,N_13383);
nor U18156 (N_18156,N_13213,N_13286);
nand U18157 (N_18157,N_14083,N_12617);
or U18158 (N_18158,N_13789,N_11881);
nor U18159 (N_18159,N_11859,N_10109);
xnor U18160 (N_18160,N_14326,N_12621);
nand U18161 (N_18161,N_14173,N_14844);
xor U18162 (N_18162,N_14927,N_11721);
xor U18163 (N_18163,N_11351,N_12883);
and U18164 (N_18164,N_12132,N_10107);
or U18165 (N_18165,N_11311,N_13072);
nand U18166 (N_18166,N_12225,N_10614);
or U18167 (N_18167,N_13115,N_11386);
or U18168 (N_18168,N_11562,N_11304);
xor U18169 (N_18169,N_11028,N_14560);
nand U18170 (N_18170,N_10392,N_11814);
nand U18171 (N_18171,N_10756,N_10518);
and U18172 (N_18172,N_12568,N_13572);
xor U18173 (N_18173,N_13666,N_12573);
nor U18174 (N_18174,N_12274,N_12796);
nor U18175 (N_18175,N_12697,N_14667);
nand U18176 (N_18176,N_11184,N_11007);
and U18177 (N_18177,N_12042,N_12419);
nor U18178 (N_18178,N_13390,N_10688);
nand U18179 (N_18179,N_12522,N_14980);
and U18180 (N_18180,N_11366,N_14328);
nand U18181 (N_18181,N_12709,N_11297);
xor U18182 (N_18182,N_11950,N_13452);
nor U18183 (N_18183,N_12385,N_14472);
nand U18184 (N_18184,N_12990,N_11838);
nor U18185 (N_18185,N_14696,N_10063);
or U18186 (N_18186,N_14107,N_10337);
or U18187 (N_18187,N_13783,N_12758);
and U18188 (N_18188,N_13161,N_14861);
nor U18189 (N_18189,N_10114,N_13405);
xnor U18190 (N_18190,N_13115,N_12980);
or U18191 (N_18191,N_13019,N_12216);
nand U18192 (N_18192,N_13434,N_10905);
nand U18193 (N_18193,N_12442,N_12056);
nor U18194 (N_18194,N_11361,N_12878);
xnor U18195 (N_18195,N_13839,N_14637);
or U18196 (N_18196,N_12666,N_13406);
xor U18197 (N_18197,N_10860,N_10339);
xnor U18198 (N_18198,N_13132,N_14113);
or U18199 (N_18199,N_13869,N_12359);
or U18200 (N_18200,N_13619,N_14699);
xor U18201 (N_18201,N_10760,N_14865);
and U18202 (N_18202,N_11696,N_13086);
nor U18203 (N_18203,N_10884,N_10147);
xor U18204 (N_18204,N_10126,N_13299);
xnor U18205 (N_18205,N_10803,N_11010);
xor U18206 (N_18206,N_14255,N_13106);
nor U18207 (N_18207,N_13040,N_13527);
and U18208 (N_18208,N_14569,N_10828);
or U18209 (N_18209,N_11079,N_14764);
xor U18210 (N_18210,N_11818,N_12232);
or U18211 (N_18211,N_10037,N_10066);
or U18212 (N_18212,N_10988,N_14928);
xor U18213 (N_18213,N_10506,N_11442);
nor U18214 (N_18214,N_10574,N_13206);
nand U18215 (N_18215,N_14950,N_11440);
nand U18216 (N_18216,N_12605,N_10847);
nand U18217 (N_18217,N_13918,N_11464);
nand U18218 (N_18218,N_12946,N_11027);
or U18219 (N_18219,N_11144,N_11558);
and U18220 (N_18220,N_12478,N_12854);
nand U18221 (N_18221,N_14648,N_10123);
nand U18222 (N_18222,N_13229,N_10711);
xnor U18223 (N_18223,N_11642,N_14236);
and U18224 (N_18224,N_14352,N_14554);
and U18225 (N_18225,N_10849,N_11952);
or U18226 (N_18226,N_11854,N_10564);
and U18227 (N_18227,N_11499,N_11159);
or U18228 (N_18228,N_10606,N_10008);
or U18229 (N_18229,N_13258,N_14124);
or U18230 (N_18230,N_14815,N_14928);
xnor U18231 (N_18231,N_11531,N_14815);
nor U18232 (N_18232,N_10194,N_14760);
nand U18233 (N_18233,N_13670,N_14119);
and U18234 (N_18234,N_11689,N_13569);
nand U18235 (N_18235,N_14811,N_12215);
and U18236 (N_18236,N_13811,N_12516);
and U18237 (N_18237,N_12393,N_13693);
or U18238 (N_18238,N_14772,N_11066);
or U18239 (N_18239,N_14003,N_11773);
nor U18240 (N_18240,N_13457,N_13608);
nand U18241 (N_18241,N_14953,N_14049);
nand U18242 (N_18242,N_10938,N_10257);
xnor U18243 (N_18243,N_10847,N_12139);
nand U18244 (N_18244,N_12700,N_11871);
xor U18245 (N_18245,N_11352,N_10038);
or U18246 (N_18246,N_12933,N_11431);
nor U18247 (N_18247,N_11952,N_11772);
and U18248 (N_18248,N_10568,N_11782);
and U18249 (N_18249,N_10546,N_14751);
xor U18250 (N_18250,N_14678,N_14153);
nand U18251 (N_18251,N_14856,N_12699);
nand U18252 (N_18252,N_10165,N_13752);
or U18253 (N_18253,N_10425,N_13608);
nor U18254 (N_18254,N_14242,N_13973);
nor U18255 (N_18255,N_13976,N_12863);
nor U18256 (N_18256,N_13121,N_10680);
nor U18257 (N_18257,N_11877,N_14174);
nand U18258 (N_18258,N_10219,N_14585);
and U18259 (N_18259,N_11711,N_13778);
nand U18260 (N_18260,N_13437,N_12526);
nor U18261 (N_18261,N_11422,N_12125);
or U18262 (N_18262,N_11149,N_11033);
or U18263 (N_18263,N_13992,N_11628);
xnor U18264 (N_18264,N_13918,N_14282);
nor U18265 (N_18265,N_12509,N_10974);
nor U18266 (N_18266,N_12809,N_12299);
and U18267 (N_18267,N_14276,N_14069);
and U18268 (N_18268,N_10340,N_14063);
and U18269 (N_18269,N_12960,N_10540);
xnor U18270 (N_18270,N_10987,N_12868);
or U18271 (N_18271,N_11695,N_12950);
or U18272 (N_18272,N_11993,N_13674);
nor U18273 (N_18273,N_10531,N_10768);
nand U18274 (N_18274,N_10777,N_10231);
nand U18275 (N_18275,N_11524,N_11138);
nand U18276 (N_18276,N_11193,N_13198);
or U18277 (N_18277,N_14962,N_14553);
or U18278 (N_18278,N_12687,N_14872);
xor U18279 (N_18279,N_11362,N_14344);
nand U18280 (N_18280,N_12151,N_13296);
or U18281 (N_18281,N_13974,N_11227);
and U18282 (N_18282,N_10935,N_10928);
xor U18283 (N_18283,N_11830,N_11406);
nand U18284 (N_18284,N_14120,N_11088);
nor U18285 (N_18285,N_13667,N_13457);
or U18286 (N_18286,N_10856,N_10881);
and U18287 (N_18287,N_10147,N_14438);
and U18288 (N_18288,N_10875,N_13676);
nor U18289 (N_18289,N_13377,N_11301);
xor U18290 (N_18290,N_14367,N_12802);
nor U18291 (N_18291,N_14646,N_10678);
xnor U18292 (N_18292,N_13252,N_14139);
and U18293 (N_18293,N_14721,N_14367);
xor U18294 (N_18294,N_12908,N_11142);
nand U18295 (N_18295,N_13584,N_10732);
or U18296 (N_18296,N_10250,N_11272);
xnor U18297 (N_18297,N_11529,N_11926);
nor U18298 (N_18298,N_11846,N_13343);
or U18299 (N_18299,N_14113,N_11894);
nand U18300 (N_18300,N_14001,N_14683);
and U18301 (N_18301,N_12018,N_14871);
nor U18302 (N_18302,N_13265,N_13765);
or U18303 (N_18303,N_13074,N_11761);
and U18304 (N_18304,N_10520,N_14479);
nand U18305 (N_18305,N_12289,N_11700);
xor U18306 (N_18306,N_10539,N_14608);
or U18307 (N_18307,N_12838,N_10692);
xnor U18308 (N_18308,N_14855,N_14937);
nand U18309 (N_18309,N_11905,N_13224);
nand U18310 (N_18310,N_11514,N_11527);
or U18311 (N_18311,N_12388,N_12551);
xor U18312 (N_18312,N_13064,N_14507);
nand U18313 (N_18313,N_13753,N_13309);
nand U18314 (N_18314,N_11982,N_11417);
or U18315 (N_18315,N_14772,N_12975);
nand U18316 (N_18316,N_12691,N_13426);
xor U18317 (N_18317,N_10308,N_11019);
and U18318 (N_18318,N_13371,N_10289);
xnor U18319 (N_18319,N_12502,N_10272);
xnor U18320 (N_18320,N_12801,N_12989);
nor U18321 (N_18321,N_11228,N_11408);
or U18322 (N_18322,N_10685,N_13422);
or U18323 (N_18323,N_13551,N_14145);
nand U18324 (N_18324,N_12684,N_10466);
or U18325 (N_18325,N_13349,N_10599);
or U18326 (N_18326,N_14627,N_14926);
nor U18327 (N_18327,N_13207,N_12592);
nor U18328 (N_18328,N_12005,N_12974);
nor U18329 (N_18329,N_14376,N_14315);
xnor U18330 (N_18330,N_13773,N_10783);
and U18331 (N_18331,N_10502,N_14412);
xnor U18332 (N_18332,N_11491,N_12960);
nor U18333 (N_18333,N_10752,N_14458);
xor U18334 (N_18334,N_13718,N_14529);
or U18335 (N_18335,N_12919,N_10166);
and U18336 (N_18336,N_10734,N_13105);
or U18337 (N_18337,N_10067,N_12792);
xnor U18338 (N_18338,N_14808,N_12977);
nor U18339 (N_18339,N_12784,N_14714);
nand U18340 (N_18340,N_12762,N_13144);
and U18341 (N_18341,N_12466,N_12091);
xor U18342 (N_18342,N_11652,N_13045);
nor U18343 (N_18343,N_14759,N_10317);
and U18344 (N_18344,N_13447,N_14186);
or U18345 (N_18345,N_14491,N_13214);
nor U18346 (N_18346,N_11912,N_13201);
and U18347 (N_18347,N_13274,N_10528);
xor U18348 (N_18348,N_14280,N_12189);
xnor U18349 (N_18349,N_14439,N_12173);
or U18350 (N_18350,N_12523,N_14257);
xor U18351 (N_18351,N_13313,N_11765);
or U18352 (N_18352,N_10280,N_13233);
and U18353 (N_18353,N_11584,N_12978);
xnor U18354 (N_18354,N_10595,N_13443);
and U18355 (N_18355,N_13763,N_12020);
or U18356 (N_18356,N_12691,N_14756);
nand U18357 (N_18357,N_14687,N_14228);
nand U18358 (N_18358,N_12351,N_12757);
nand U18359 (N_18359,N_13011,N_14100);
nand U18360 (N_18360,N_13182,N_12148);
nor U18361 (N_18361,N_12780,N_12668);
nor U18362 (N_18362,N_14216,N_12444);
and U18363 (N_18363,N_13518,N_11317);
nor U18364 (N_18364,N_12951,N_13758);
nor U18365 (N_18365,N_13863,N_13315);
xnor U18366 (N_18366,N_13696,N_10017);
or U18367 (N_18367,N_11974,N_11348);
and U18368 (N_18368,N_12045,N_11370);
and U18369 (N_18369,N_11159,N_10489);
nor U18370 (N_18370,N_13193,N_12019);
nand U18371 (N_18371,N_10949,N_10718);
and U18372 (N_18372,N_14183,N_14168);
or U18373 (N_18373,N_12485,N_14656);
xnor U18374 (N_18374,N_10385,N_13333);
xor U18375 (N_18375,N_12958,N_10758);
or U18376 (N_18376,N_11422,N_12976);
or U18377 (N_18377,N_11405,N_10623);
nand U18378 (N_18378,N_11952,N_12057);
or U18379 (N_18379,N_13002,N_11071);
or U18380 (N_18380,N_12969,N_10469);
xor U18381 (N_18381,N_14836,N_13187);
xor U18382 (N_18382,N_14171,N_12528);
or U18383 (N_18383,N_13043,N_14935);
nor U18384 (N_18384,N_10899,N_13239);
or U18385 (N_18385,N_13422,N_11609);
and U18386 (N_18386,N_10548,N_10623);
and U18387 (N_18387,N_11792,N_11336);
xnor U18388 (N_18388,N_11570,N_13037);
nand U18389 (N_18389,N_11429,N_10503);
and U18390 (N_18390,N_10613,N_11191);
and U18391 (N_18391,N_14200,N_11208);
nor U18392 (N_18392,N_10084,N_10337);
nand U18393 (N_18393,N_11792,N_14606);
xor U18394 (N_18394,N_10182,N_14205);
and U18395 (N_18395,N_14708,N_11787);
xor U18396 (N_18396,N_13360,N_10866);
and U18397 (N_18397,N_12784,N_11490);
nand U18398 (N_18398,N_11846,N_14282);
nand U18399 (N_18399,N_11143,N_13809);
and U18400 (N_18400,N_13703,N_10673);
or U18401 (N_18401,N_12331,N_11384);
and U18402 (N_18402,N_12547,N_13517);
nand U18403 (N_18403,N_10540,N_12984);
or U18404 (N_18404,N_10469,N_12207);
nand U18405 (N_18405,N_11873,N_14428);
xor U18406 (N_18406,N_10705,N_10085);
or U18407 (N_18407,N_13525,N_12032);
or U18408 (N_18408,N_14908,N_10345);
nor U18409 (N_18409,N_11050,N_11943);
xnor U18410 (N_18410,N_13911,N_13720);
and U18411 (N_18411,N_11566,N_10409);
nand U18412 (N_18412,N_13145,N_14187);
xor U18413 (N_18413,N_10300,N_12366);
and U18414 (N_18414,N_13654,N_13763);
nand U18415 (N_18415,N_12689,N_10531);
and U18416 (N_18416,N_13274,N_14739);
nand U18417 (N_18417,N_12753,N_10337);
and U18418 (N_18418,N_11729,N_14088);
nor U18419 (N_18419,N_14454,N_11133);
and U18420 (N_18420,N_13715,N_12092);
or U18421 (N_18421,N_10517,N_12372);
nor U18422 (N_18422,N_14938,N_10262);
nor U18423 (N_18423,N_10110,N_10589);
nor U18424 (N_18424,N_11144,N_10680);
nand U18425 (N_18425,N_14651,N_13438);
and U18426 (N_18426,N_13101,N_12323);
nand U18427 (N_18427,N_10414,N_13442);
and U18428 (N_18428,N_12655,N_14421);
nand U18429 (N_18429,N_13887,N_11425);
or U18430 (N_18430,N_13911,N_10247);
nand U18431 (N_18431,N_13018,N_14777);
nand U18432 (N_18432,N_13277,N_12188);
nor U18433 (N_18433,N_12851,N_11362);
xnor U18434 (N_18434,N_12558,N_12216);
or U18435 (N_18435,N_12179,N_14248);
nor U18436 (N_18436,N_13803,N_11257);
or U18437 (N_18437,N_14928,N_10029);
nor U18438 (N_18438,N_12662,N_10102);
or U18439 (N_18439,N_11125,N_14254);
and U18440 (N_18440,N_11928,N_13695);
xnor U18441 (N_18441,N_13266,N_14433);
and U18442 (N_18442,N_11847,N_14224);
nor U18443 (N_18443,N_14807,N_10272);
nand U18444 (N_18444,N_11192,N_11624);
xor U18445 (N_18445,N_13356,N_12197);
nor U18446 (N_18446,N_10397,N_11366);
nand U18447 (N_18447,N_10501,N_13396);
or U18448 (N_18448,N_14950,N_11376);
xor U18449 (N_18449,N_11156,N_11428);
nor U18450 (N_18450,N_12735,N_10964);
xor U18451 (N_18451,N_11154,N_14570);
and U18452 (N_18452,N_12171,N_13812);
xor U18453 (N_18453,N_11877,N_14071);
nand U18454 (N_18454,N_13882,N_14719);
nand U18455 (N_18455,N_11416,N_11713);
and U18456 (N_18456,N_12394,N_10640);
or U18457 (N_18457,N_14023,N_12491);
and U18458 (N_18458,N_13099,N_11447);
nand U18459 (N_18459,N_12437,N_12325);
nor U18460 (N_18460,N_12633,N_11865);
nor U18461 (N_18461,N_13285,N_12456);
nand U18462 (N_18462,N_11525,N_10162);
or U18463 (N_18463,N_11863,N_12584);
and U18464 (N_18464,N_13976,N_10994);
nand U18465 (N_18465,N_10228,N_11363);
xor U18466 (N_18466,N_12748,N_11242);
nor U18467 (N_18467,N_11402,N_12701);
nor U18468 (N_18468,N_11918,N_11181);
nor U18469 (N_18469,N_13253,N_10601);
xor U18470 (N_18470,N_10510,N_14414);
or U18471 (N_18471,N_13842,N_13643);
nor U18472 (N_18472,N_11707,N_13481);
and U18473 (N_18473,N_12032,N_13476);
nand U18474 (N_18474,N_13099,N_10890);
or U18475 (N_18475,N_14570,N_11887);
or U18476 (N_18476,N_13394,N_13203);
xor U18477 (N_18477,N_11119,N_12768);
xnor U18478 (N_18478,N_12349,N_14992);
xnor U18479 (N_18479,N_14604,N_13013);
and U18480 (N_18480,N_14242,N_12886);
nand U18481 (N_18481,N_13758,N_10652);
and U18482 (N_18482,N_10204,N_12027);
nand U18483 (N_18483,N_10918,N_11939);
or U18484 (N_18484,N_10840,N_13548);
nand U18485 (N_18485,N_12127,N_14480);
and U18486 (N_18486,N_11383,N_12357);
and U18487 (N_18487,N_12288,N_11434);
nand U18488 (N_18488,N_13920,N_10149);
or U18489 (N_18489,N_14945,N_10164);
nor U18490 (N_18490,N_14642,N_11989);
or U18491 (N_18491,N_13330,N_10036);
nor U18492 (N_18492,N_11391,N_13058);
or U18493 (N_18493,N_13292,N_10189);
and U18494 (N_18494,N_11711,N_13066);
or U18495 (N_18495,N_12041,N_14961);
or U18496 (N_18496,N_13685,N_10247);
or U18497 (N_18497,N_13635,N_11004);
and U18498 (N_18498,N_14600,N_14734);
nor U18499 (N_18499,N_14372,N_12048);
and U18500 (N_18500,N_13802,N_12722);
nand U18501 (N_18501,N_14726,N_14308);
nand U18502 (N_18502,N_13159,N_13653);
nand U18503 (N_18503,N_11256,N_12711);
nand U18504 (N_18504,N_11885,N_11833);
nand U18505 (N_18505,N_10966,N_13426);
and U18506 (N_18506,N_12860,N_11767);
and U18507 (N_18507,N_10191,N_11137);
or U18508 (N_18508,N_12554,N_12392);
nor U18509 (N_18509,N_10891,N_13184);
or U18510 (N_18510,N_14426,N_10997);
or U18511 (N_18511,N_10578,N_14272);
xnor U18512 (N_18512,N_14529,N_13289);
xnor U18513 (N_18513,N_13788,N_13511);
or U18514 (N_18514,N_12257,N_14778);
or U18515 (N_18515,N_12167,N_14745);
and U18516 (N_18516,N_14277,N_11294);
nor U18517 (N_18517,N_10225,N_12219);
xor U18518 (N_18518,N_10463,N_14012);
nor U18519 (N_18519,N_12853,N_12522);
nor U18520 (N_18520,N_10830,N_10108);
and U18521 (N_18521,N_12067,N_11496);
and U18522 (N_18522,N_10153,N_12231);
or U18523 (N_18523,N_11714,N_10304);
nand U18524 (N_18524,N_14228,N_14978);
and U18525 (N_18525,N_10387,N_11117);
and U18526 (N_18526,N_11413,N_12195);
and U18527 (N_18527,N_10212,N_13724);
xnor U18528 (N_18528,N_14603,N_13669);
nor U18529 (N_18529,N_14261,N_11720);
nor U18530 (N_18530,N_10269,N_11581);
nand U18531 (N_18531,N_11665,N_13494);
xor U18532 (N_18532,N_12579,N_11407);
and U18533 (N_18533,N_14528,N_10651);
xnor U18534 (N_18534,N_10439,N_14677);
xnor U18535 (N_18535,N_12845,N_14409);
nor U18536 (N_18536,N_11108,N_11908);
nand U18537 (N_18537,N_13910,N_13339);
nor U18538 (N_18538,N_10901,N_14363);
nand U18539 (N_18539,N_11704,N_14698);
or U18540 (N_18540,N_12788,N_11328);
or U18541 (N_18541,N_14820,N_10129);
xor U18542 (N_18542,N_10342,N_10415);
nand U18543 (N_18543,N_11775,N_14546);
xor U18544 (N_18544,N_13298,N_14276);
nor U18545 (N_18545,N_13103,N_10768);
nand U18546 (N_18546,N_14963,N_10757);
nand U18547 (N_18547,N_14983,N_13665);
nand U18548 (N_18548,N_13551,N_13996);
and U18549 (N_18549,N_12675,N_13537);
xnor U18550 (N_18550,N_10609,N_14608);
or U18551 (N_18551,N_13674,N_10137);
nand U18552 (N_18552,N_13525,N_11243);
xnor U18553 (N_18553,N_13111,N_11017);
and U18554 (N_18554,N_14817,N_12493);
nand U18555 (N_18555,N_14877,N_13835);
xnor U18556 (N_18556,N_11795,N_10655);
nor U18557 (N_18557,N_14101,N_14398);
or U18558 (N_18558,N_13553,N_11318);
xor U18559 (N_18559,N_11567,N_12449);
nor U18560 (N_18560,N_10616,N_12914);
xor U18561 (N_18561,N_14962,N_11386);
nor U18562 (N_18562,N_14829,N_13232);
nor U18563 (N_18563,N_14744,N_13428);
nor U18564 (N_18564,N_10796,N_14209);
and U18565 (N_18565,N_10077,N_11917);
nand U18566 (N_18566,N_10161,N_12200);
nand U18567 (N_18567,N_11600,N_10034);
nand U18568 (N_18568,N_14028,N_13802);
nor U18569 (N_18569,N_11821,N_13089);
nand U18570 (N_18570,N_10675,N_13983);
and U18571 (N_18571,N_13687,N_12995);
nor U18572 (N_18572,N_13752,N_13016);
nand U18573 (N_18573,N_13881,N_13204);
nor U18574 (N_18574,N_10497,N_14935);
or U18575 (N_18575,N_14254,N_12857);
nand U18576 (N_18576,N_10170,N_10411);
xnor U18577 (N_18577,N_12556,N_13228);
nand U18578 (N_18578,N_10246,N_10400);
nor U18579 (N_18579,N_10249,N_12433);
or U18580 (N_18580,N_10199,N_13755);
nand U18581 (N_18581,N_13984,N_10108);
or U18582 (N_18582,N_10971,N_12523);
nand U18583 (N_18583,N_11291,N_14380);
and U18584 (N_18584,N_11381,N_11405);
nand U18585 (N_18585,N_10243,N_14018);
xnor U18586 (N_18586,N_10099,N_13353);
nand U18587 (N_18587,N_11550,N_12996);
nand U18588 (N_18588,N_12298,N_10808);
nor U18589 (N_18589,N_12238,N_11998);
nand U18590 (N_18590,N_12279,N_12284);
xnor U18591 (N_18591,N_14994,N_11489);
or U18592 (N_18592,N_13821,N_10369);
xor U18593 (N_18593,N_11207,N_11789);
or U18594 (N_18594,N_11882,N_13711);
nor U18595 (N_18595,N_13033,N_12822);
or U18596 (N_18596,N_13614,N_10322);
nor U18597 (N_18597,N_13393,N_13302);
and U18598 (N_18598,N_14713,N_13159);
nand U18599 (N_18599,N_11383,N_13828);
xor U18600 (N_18600,N_12436,N_11748);
or U18601 (N_18601,N_13485,N_11596);
nor U18602 (N_18602,N_10172,N_10947);
and U18603 (N_18603,N_10575,N_10973);
or U18604 (N_18604,N_10719,N_14426);
nand U18605 (N_18605,N_12338,N_13174);
xor U18606 (N_18606,N_14934,N_14268);
or U18607 (N_18607,N_14474,N_10251);
nor U18608 (N_18608,N_11276,N_14920);
nand U18609 (N_18609,N_10952,N_10282);
or U18610 (N_18610,N_14492,N_12567);
or U18611 (N_18611,N_12078,N_12815);
xnor U18612 (N_18612,N_13108,N_10803);
nor U18613 (N_18613,N_12804,N_14464);
xor U18614 (N_18614,N_14708,N_11078);
or U18615 (N_18615,N_12065,N_12338);
nand U18616 (N_18616,N_11117,N_13525);
and U18617 (N_18617,N_12094,N_12428);
xor U18618 (N_18618,N_13426,N_13182);
and U18619 (N_18619,N_13160,N_13847);
and U18620 (N_18620,N_13299,N_12118);
xnor U18621 (N_18621,N_13842,N_14506);
and U18622 (N_18622,N_12934,N_11267);
xnor U18623 (N_18623,N_12706,N_12726);
and U18624 (N_18624,N_14472,N_11645);
or U18625 (N_18625,N_14234,N_13023);
nor U18626 (N_18626,N_13531,N_13540);
nor U18627 (N_18627,N_11544,N_12461);
nor U18628 (N_18628,N_12524,N_14845);
nor U18629 (N_18629,N_14989,N_10975);
nor U18630 (N_18630,N_12290,N_14336);
and U18631 (N_18631,N_12598,N_13942);
nand U18632 (N_18632,N_13333,N_10637);
and U18633 (N_18633,N_14853,N_12128);
nor U18634 (N_18634,N_12264,N_13513);
and U18635 (N_18635,N_10878,N_12987);
xor U18636 (N_18636,N_14906,N_14255);
or U18637 (N_18637,N_11430,N_10429);
and U18638 (N_18638,N_14652,N_11026);
and U18639 (N_18639,N_12224,N_12275);
and U18640 (N_18640,N_14700,N_14102);
nor U18641 (N_18641,N_14441,N_13097);
or U18642 (N_18642,N_11579,N_13862);
xor U18643 (N_18643,N_14944,N_12936);
xnor U18644 (N_18644,N_12412,N_11681);
xor U18645 (N_18645,N_10296,N_10955);
or U18646 (N_18646,N_12200,N_10911);
or U18647 (N_18647,N_11536,N_13271);
or U18648 (N_18648,N_13499,N_10322);
and U18649 (N_18649,N_13639,N_12712);
and U18650 (N_18650,N_14381,N_12580);
or U18651 (N_18651,N_14676,N_12248);
nor U18652 (N_18652,N_13917,N_10123);
or U18653 (N_18653,N_12580,N_13742);
or U18654 (N_18654,N_12602,N_10467);
and U18655 (N_18655,N_14918,N_14176);
and U18656 (N_18656,N_10964,N_14349);
xor U18657 (N_18657,N_12421,N_12791);
or U18658 (N_18658,N_10050,N_11200);
or U18659 (N_18659,N_11177,N_10096);
and U18660 (N_18660,N_14503,N_10470);
and U18661 (N_18661,N_13847,N_13425);
nor U18662 (N_18662,N_12936,N_14476);
and U18663 (N_18663,N_14574,N_11926);
and U18664 (N_18664,N_14471,N_11598);
and U18665 (N_18665,N_14092,N_10861);
nand U18666 (N_18666,N_11865,N_10100);
or U18667 (N_18667,N_14395,N_13782);
nand U18668 (N_18668,N_14547,N_12650);
nand U18669 (N_18669,N_14206,N_13298);
nand U18670 (N_18670,N_11407,N_12071);
or U18671 (N_18671,N_11034,N_13234);
nand U18672 (N_18672,N_11645,N_10137);
or U18673 (N_18673,N_12068,N_13425);
nand U18674 (N_18674,N_10844,N_10963);
xor U18675 (N_18675,N_12887,N_13610);
or U18676 (N_18676,N_13458,N_11072);
or U18677 (N_18677,N_13726,N_10819);
and U18678 (N_18678,N_13215,N_11701);
and U18679 (N_18679,N_12291,N_10924);
xor U18680 (N_18680,N_10039,N_11122);
or U18681 (N_18681,N_14664,N_12074);
or U18682 (N_18682,N_14764,N_13574);
and U18683 (N_18683,N_11951,N_11435);
xnor U18684 (N_18684,N_13661,N_10951);
or U18685 (N_18685,N_14998,N_12832);
or U18686 (N_18686,N_10050,N_11586);
nand U18687 (N_18687,N_11090,N_14768);
nor U18688 (N_18688,N_11290,N_11354);
or U18689 (N_18689,N_13024,N_12901);
and U18690 (N_18690,N_10036,N_10376);
nor U18691 (N_18691,N_13864,N_11721);
and U18692 (N_18692,N_10885,N_11877);
xor U18693 (N_18693,N_12557,N_11871);
xnor U18694 (N_18694,N_13412,N_14450);
xnor U18695 (N_18695,N_13834,N_10092);
or U18696 (N_18696,N_12113,N_13164);
nand U18697 (N_18697,N_11720,N_11155);
and U18698 (N_18698,N_11278,N_12327);
nand U18699 (N_18699,N_11884,N_13645);
and U18700 (N_18700,N_13055,N_13882);
nand U18701 (N_18701,N_10357,N_12944);
nor U18702 (N_18702,N_12212,N_10594);
or U18703 (N_18703,N_13644,N_13914);
nor U18704 (N_18704,N_13316,N_12465);
nor U18705 (N_18705,N_13667,N_13077);
nor U18706 (N_18706,N_10807,N_12870);
nand U18707 (N_18707,N_10126,N_13211);
xor U18708 (N_18708,N_11476,N_11962);
or U18709 (N_18709,N_14114,N_14090);
xnor U18710 (N_18710,N_10854,N_10710);
nor U18711 (N_18711,N_13850,N_13555);
nor U18712 (N_18712,N_12004,N_12965);
nor U18713 (N_18713,N_11232,N_14624);
nand U18714 (N_18714,N_13821,N_12854);
or U18715 (N_18715,N_13467,N_11481);
and U18716 (N_18716,N_14313,N_14586);
nor U18717 (N_18717,N_13686,N_11103);
nor U18718 (N_18718,N_13819,N_12354);
nand U18719 (N_18719,N_11931,N_13019);
and U18720 (N_18720,N_14713,N_14586);
and U18721 (N_18721,N_14248,N_11034);
or U18722 (N_18722,N_12448,N_10795);
xor U18723 (N_18723,N_14007,N_12546);
nor U18724 (N_18724,N_11830,N_10092);
nand U18725 (N_18725,N_10215,N_13215);
and U18726 (N_18726,N_13636,N_14743);
and U18727 (N_18727,N_14905,N_11281);
xnor U18728 (N_18728,N_10595,N_13427);
xor U18729 (N_18729,N_14310,N_14821);
or U18730 (N_18730,N_14612,N_12378);
xnor U18731 (N_18731,N_11034,N_14672);
nor U18732 (N_18732,N_14598,N_13584);
or U18733 (N_18733,N_11903,N_14594);
xor U18734 (N_18734,N_10759,N_12641);
nand U18735 (N_18735,N_13467,N_14725);
and U18736 (N_18736,N_11543,N_11816);
or U18737 (N_18737,N_14368,N_14642);
xnor U18738 (N_18738,N_13805,N_10181);
or U18739 (N_18739,N_11641,N_14317);
and U18740 (N_18740,N_11671,N_13619);
xnor U18741 (N_18741,N_10062,N_13510);
or U18742 (N_18742,N_14781,N_14074);
and U18743 (N_18743,N_12385,N_12176);
and U18744 (N_18744,N_10623,N_12524);
nor U18745 (N_18745,N_10396,N_10079);
or U18746 (N_18746,N_14358,N_12601);
nor U18747 (N_18747,N_13919,N_14358);
or U18748 (N_18748,N_12322,N_10572);
or U18749 (N_18749,N_14402,N_11941);
or U18750 (N_18750,N_13459,N_11576);
or U18751 (N_18751,N_11503,N_12860);
or U18752 (N_18752,N_13549,N_14074);
xor U18753 (N_18753,N_14621,N_12938);
nor U18754 (N_18754,N_13121,N_13167);
xor U18755 (N_18755,N_12285,N_12445);
nand U18756 (N_18756,N_12200,N_12397);
nor U18757 (N_18757,N_13930,N_10469);
nor U18758 (N_18758,N_10242,N_12640);
and U18759 (N_18759,N_11748,N_10951);
xnor U18760 (N_18760,N_10175,N_14835);
and U18761 (N_18761,N_12709,N_12608);
xor U18762 (N_18762,N_10225,N_14046);
and U18763 (N_18763,N_14619,N_14579);
and U18764 (N_18764,N_10204,N_10250);
nor U18765 (N_18765,N_12768,N_13988);
xor U18766 (N_18766,N_14261,N_11890);
nand U18767 (N_18767,N_12776,N_11276);
and U18768 (N_18768,N_13500,N_11092);
and U18769 (N_18769,N_12317,N_13125);
nor U18770 (N_18770,N_12167,N_10804);
nor U18771 (N_18771,N_12534,N_13241);
nor U18772 (N_18772,N_11874,N_11200);
nor U18773 (N_18773,N_13397,N_10011);
nor U18774 (N_18774,N_11611,N_14667);
nor U18775 (N_18775,N_14536,N_11281);
or U18776 (N_18776,N_12190,N_10957);
xor U18777 (N_18777,N_10073,N_14396);
nand U18778 (N_18778,N_13021,N_14068);
nor U18779 (N_18779,N_10955,N_11149);
nand U18780 (N_18780,N_11419,N_13396);
nor U18781 (N_18781,N_12809,N_12143);
nand U18782 (N_18782,N_14267,N_13644);
or U18783 (N_18783,N_10402,N_13014);
nor U18784 (N_18784,N_10264,N_14477);
nand U18785 (N_18785,N_12305,N_12101);
nor U18786 (N_18786,N_11278,N_11776);
or U18787 (N_18787,N_14499,N_14467);
nor U18788 (N_18788,N_12792,N_13796);
nor U18789 (N_18789,N_11566,N_10938);
and U18790 (N_18790,N_14159,N_10540);
nor U18791 (N_18791,N_13637,N_14254);
nand U18792 (N_18792,N_11545,N_11638);
and U18793 (N_18793,N_14026,N_10504);
and U18794 (N_18794,N_13568,N_10247);
and U18795 (N_18795,N_12008,N_10335);
xnor U18796 (N_18796,N_10535,N_11188);
and U18797 (N_18797,N_12341,N_13501);
nor U18798 (N_18798,N_11047,N_13048);
nor U18799 (N_18799,N_11420,N_12171);
or U18800 (N_18800,N_14619,N_11895);
nand U18801 (N_18801,N_11458,N_12175);
nand U18802 (N_18802,N_12922,N_14599);
nand U18803 (N_18803,N_11899,N_10890);
nand U18804 (N_18804,N_13209,N_12345);
xor U18805 (N_18805,N_10731,N_14453);
or U18806 (N_18806,N_13112,N_13297);
nand U18807 (N_18807,N_12021,N_14854);
xnor U18808 (N_18808,N_13970,N_14294);
or U18809 (N_18809,N_13703,N_12621);
or U18810 (N_18810,N_11910,N_11011);
xor U18811 (N_18811,N_10543,N_12793);
and U18812 (N_18812,N_12237,N_14780);
xor U18813 (N_18813,N_13576,N_14518);
xnor U18814 (N_18814,N_12139,N_10867);
nand U18815 (N_18815,N_10021,N_13209);
nand U18816 (N_18816,N_11930,N_11901);
nand U18817 (N_18817,N_10539,N_12868);
nor U18818 (N_18818,N_12182,N_11373);
nor U18819 (N_18819,N_12988,N_12477);
or U18820 (N_18820,N_12952,N_11554);
nand U18821 (N_18821,N_13301,N_10311);
nor U18822 (N_18822,N_12208,N_12360);
nand U18823 (N_18823,N_14912,N_12662);
nand U18824 (N_18824,N_11951,N_10711);
xor U18825 (N_18825,N_12335,N_10883);
and U18826 (N_18826,N_13943,N_11162);
or U18827 (N_18827,N_14015,N_10340);
nand U18828 (N_18828,N_11554,N_13440);
or U18829 (N_18829,N_11881,N_11362);
nor U18830 (N_18830,N_14293,N_14271);
and U18831 (N_18831,N_10132,N_13800);
nand U18832 (N_18832,N_13841,N_11511);
nand U18833 (N_18833,N_14614,N_13078);
nand U18834 (N_18834,N_13396,N_11545);
xor U18835 (N_18835,N_14331,N_14875);
nor U18836 (N_18836,N_11591,N_14039);
or U18837 (N_18837,N_10192,N_10617);
nor U18838 (N_18838,N_11496,N_10997);
xnor U18839 (N_18839,N_10676,N_12155);
xnor U18840 (N_18840,N_10830,N_13485);
or U18841 (N_18841,N_12690,N_14291);
or U18842 (N_18842,N_10117,N_11944);
or U18843 (N_18843,N_12725,N_13173);
nand U18844 (N_18844,N_13386,N_10785);
nor U18845 (N_18845,N_11235,N_13421);
and U18846 (N_18846,N_13015,N_10056);
or U18847 (N_18847,N_10349,N_14584);
or U18848 (N_18848,N_11152,N_13111);
nand U18849 (N_18849,N_10733,N_13973);
and U18850 (N_18850,N_11448,N_13340);
nand U18851 (N_18851,N_12695,N_13067);
and U18852 (N_18852,N_11136,N_12907);
nor U18853 (N_18853,N_14653,N_11002);
or U18854 (N_18854,N_14714,N_12638);
nor U18855 (N_18855,N_11422,N_13643);
xnor U18856 (N_18856,N_10403,N_11776);
nand U18857 (N_18857,N_14824,N_10661);
and U18858 (N_18858,N_13186,N_10636);
and U18859 (N_18859,N_13884,N_13520);
nand U18860 (N_18860,N_12243,N_13100);
nand U18861 (N_18861,N_11311,N_13092);
or U18862 (N_18862,N_10221,N_11096);
nor U18863 (N_18863,N_12654,N_12467);
or U18864 (N_18864,N_14549,N_11357);
or U18865 (N_18865,N_12505,N_11500);
or U18866 (N_18866,N_14390,N_14461);
xor U18867 (N_18867,N_13097,N_10991);
nor U18868 (N_18868,N_14714,N_11178);
xor U18869 (N_18869,N_11702,N_13491);
nand U18870 (N_18870,N_10914,N_12844);
nor U18871 (N_18871,N_10137,N_13115);
nand U18872 (N_18872,N_12674,N_13105);
and U18873 (N_18873,N_13570,N_10194);
or U18874 (N_18874,N_10095,N_13679);
and U18875 (N_18875,N_11694,N_10979);
xor U18876 (N_18876,N_11957,N_13458);
xnor U18877 (N_18877,N_11969,N_14449);
xor U18878 (N_18878,N_13170,N_12321);
nand U18879 (N_18879,N_13080,N_13309);
nor U18880 (N_18880,N_11335,N_10968);
nand U18881 (N_18881,N_11710,N_14356);
nand U18882 (N_18882,N_11178,N_10649);
or U18883 (N_18883,N_10926,N_13145);
nand U18884 (N_18884,N_10698,N_13026);
or U18885 (N_18885,N_11404,N_13644);
or U18886 (N_18886,N_14398,N_14484);
or U18887 (N_18887,N_13120,N_12576);
or U18888 (N_18888,N_10110,N_14808);
nand U18889 (N_18889,N_12823,N_11547);
or U18890 (N_18890,N_11272,N_12017);
nor U18891 (N_18891,N_13734,N_13097);
or U18892 (N_18892,N_10710,N_13201);
nor U18893 (N_18893,N_14452,N_14032);
nor U18894 (N_18894,N_11696,N_11689);
nand U18895 (N_18895,N_10491,N_11229);
nor U18896 (N_18896,N_13245,N_14747);
xor U18897 (N_18897,N_13072,N_14901);
nor U18898 (N_18898,N_14683,N_14326);
and U18899 (N_18899,N_14436,N_14822);
and U18900 (N_18900,N_14508,N_12038);
or U18901 (N_18901,N_12806,N_11818);
or U18902 (N_18902,N_13575,N_12627);
or U18903 (N_18903,N_13310,N_12996);
or U18904 (N_18904,N_12880,N_11349);
nor U18905 (N_18905,N_10395,N_11356);
or U18906 (N_18906,N_11912,N_10281);
nor U18907 (N_18907,N_13736,N_14547);
nand U18908 (N_18908,N_13091,N_12032);
nor U18909 (N_18909,N_13222,N_12566);
xnor U18910 (N_18910,N_14366,N_13262);
xor U18911 (N_18911,N_13139,N_13453);
xnor U18912 (N_18912,N_13707,N_14838);
nand U18913 (N_18913,N_10791,N_10978);
xor U18914 (N_18914,N_11390,N_14692);
nand U18915 (N_18915,N_13105,N_14288);
nand U18916 (N_18916,N_11992,N_14374);
or U18917 (N_18917,N_10791,N_13546);
xnor U18918 (N_18918,N_12552,N_11439);
xnor U18919 (N_18919,N_11285,N_11258);
and U18920 (N_18920,N_14772,N_10270);
and U18921 (N_18921,N_13042,N_10546);
nor U18922 (N_18922,N_14446,N_12701);
xnor U18923 (N_18923,N_14857,N_14476);
nor U18924 (N_18924,N_11596,N_12077);
or U18925 (N_18925,N_14647,N_12318);
xor U18926 (N_18926,N_13630,N_14906);
and U18927 (N_18927,N_11503,N_11515);
and U18928 (N_18928,N_13162,N_14168);
nor U18929 (N_18929,N_12873,N_10992);
or U18930 (N_18930,N_12317,N_10338);
nand U18931 (N_18931,N_10923,N_13488);
xor U18932 (N_18932,N_13111,N_14609);
or U18933 (N_18933,N_10409,N_10144);
xor U18934 (N_18934,N_12500,N_13652);
xor U18935 (N_18935,N_11393,N_13102);
or U18936 (N_18936,N_13322,N_14544);
nor U18937 (N_18937,N_11110,N_10782);
nand U18938 (N_18938,N_11094,N_13614);
nor U18939 (N_18939,N_11140,N_12981);
xnor U18940 (N_18940,N_11134,N_12759);
nor U18941 (N_18941,N_11566,N_11344);
nand U18942 (N_18942,N_14863,N_12752);
or U18943 (N_18943,N_11449,N_10788);
xor U18944 (N_18944,N_12313,N_13088);
nand U18945 (N_18945,N_12239,N_14779);
or U18946 (N_18946,N_11920,N_14595);
or U18947 (N_18947,N_12330,N_14640);
nor U18948 (N_18948,N_14498,N_10401);
nor U18949 (N_18949,N_14095,N_11139);
and U18950 (N_18950,N_12069,N_14294);
and U18951 (N_18951,N_13049,N_10927);
nor U18952 (N_18952,N_12073,N_13688);
nor U18953 (N_18953,N_10634,N_11408);
and U18954 (N_18954,N_11555,N_13180);
nand U18955 (N_18955,N_11333,N_10293);
and U18956 (N_18956,N_11362,N_12628);
or U18957 (N_18957,N_14312,N_13562);
xnor U18958 (N_18958,N_11823,N_12715);
and U18959 (N_18959,N_11768,N_12794);
and U18960 (N_18960,N_10427,N_11153);
nor U18961 (N_18961,N_10082,N_12783);
nor U18962 (N_18962,N_12662,N_10316);
nand U18963 (N_18963,N_14201,N_12343);
xnor U18964 (N_18964,N_13926,N_11578);
nor U18965 (N_18965,N_11408,N_11331);
nand U18966 (N_18966,N_11177,N_11798);
nand U18967 (N_18967,N_12572,N_11893);
nor U18968 (N_18968,N_14420,N_13278);
or U18969 (N_18969,N_11627,N_11867);
nor U18970 (N_18970,N_12309,N_11342);
nor U18971 (N_18971,N_10472,N_10126);
nand U18972 (N_18972,N_11143,N_14492);
and U18973 (N_18973,N_13803,N_14346);
nand U18974 (N_18974,N_10344,N_11693);
nor U18975 (N_18975,N_10373,N_11225);
xnor U18976 (N_18976,N_11093,N_12797);
nand U18977 (N_18977,N_12390,N_14994);
nor U18978 (N_18978,N_13159,N_11102);
or U18979 (N_18979,N_11476,N_11140);
nor U18980 (N_18980,N_10991,N_13088);
nor U18981 (N_18981,N_10169,N_11013);
xor U18982 (N_18982,N_12262,N_11232);
nand U18983 (N_18983,N_11193,N_13651);
or U18984 (N_18984,N_13038,N_14373);
and U18985 (N_18985,N_11585,N_13656);
nand U18986 (N_18986,N_14167,N_13110);
xnor U18987 (N_18987,N_13815,N_12586);
nor U18988 (N_18988,N_12553,N_10868);
nand U18989 (N_18989,N_10424,N_13907);
or U18990 (N_18990,N_11283,N_10570);
nor U18991 (N_18991,N_11152,N_12432);
nor U18992 (N_18992,N_12181,N_13138);
or U18993 (N_18993,N_14189,N_11181);
nor U18994 (N_18994,N_11795,N_10553);
nand U18995 (N_18995,N_13646,N_14842);
and U18996 (N_18996,N_13004,N_11625);
or U18997 (N_18997,N_14669,N_11416);
and U18998 (N_18998,N_11550,N_11620);
xor U18999 (N_18999,N_12666,N_11428);
nand U19000 (N_19000,N_10104,N_10198);
nor U19001 (N_19001,N_13194,N_10432);
and U19002 (N_19002,N_13810,N_11755);
xor U19003 (N_19003,N_11844,N_14947);
nor U19004 (N_19004,N_13381,N_14724);
or U19005 (N_19005,N_14662,N_13647);
nand U19006 (N_19006,N_14713,N_14554);
nor U19007 (N_19007,N_14768,N_12925);
nand U19008 (N_19008,N_12136,N_12011);
nor U19009 (N_19009,N_10189,N_13028);
xnor U19010 (N_19010,N_10630,N_14943);
xor U19011 (N_19011,N_10088,N_14604);
nor U19012 (N_19012,N_14864,N_13116);
nand U19013 (N_19013,N_12411,N_12115);
or U19014 (N_19014,N_11541,N_11726);
nor U19015 (N_19015,N_11805,N_13932);
nor U19016 (N_19016,N_11726,N_13108);
nor U19017 (N_19017,N_11450,N_11587);
and U19018 (N_19018,N_12601,N_11584);
nor U19019 (N_19019,N_11480,N_11142);
nor U19020 (N_19020,N_14269,N_12883);
xor U19021 (N_19021,N_10088,N_14522);
xnor U19022 (N_19022,N_11019,N_14823);
nor U19023 (N_19023,N_14336,N_10977);
and U19024 (N_19024,N_11153,N_13921);
or U19025 (N_19025,N_14928,N_14688);
nor U19026 (N_19026,N_11674,N_11988);
nor U19027 (N_19027,N_13706,N_10394);
and U19028 (N_19028,N_13588,N_11817);
or U19029 (N_19029,N_10737,N_14291);
nand U19030 (N_19030,N_12865,N_13186);
xnor U19031 (N_19031,N_10651,N_12432);
and U19032 (N_19032,N_13677,N_11626);
and U19033 (N_19033,N_13956,N_13709);
xnor U19034 (N_19034,N_12584,N_10291);
nand U19035 (N_19035,N_11694,N_11663);
xor U19036 (N_19036,N_13901,N_13965);
xor U19037 (N_19037,N_10882,N_14130);
nor U19038 (N_19038,N_12943,N_11037);
nor U19039 (N_19039,N_10028,N_13118);
or U19040 (N_19040,N_13914,N_11496);
and U19041 (N_19041,N_13052,N_13189);
nand U19042 (N_19042,N_14202,N_10911);
nor U19043 (N_19043,N_10283,N_14457);
nand U19044 (N_19044,N_14635,N_14184);
or U19045 (N_19045,N_10330,N_13943);
nor U19046 (N_19046,N_14122,N_14409);
and U19047 (N_19047,N_11497,N_11866);
and U19048 (N_19048,N_14258,N_14101);
nand U19049 (N_19049,N_11971,N_13462);
nor U19050 (N_19050,N_13776,N_14147);
xnor U19051 (N_19051,N_11164,N_11335);
and U19052 (N_19052,N_10066,N_10145);
or U19053 (N_19053,N_12137,N_14656);
and U19054 (N_19054,N_14203,N_14891);
and U19055 (N_19055,N_13735,N_13260);
xor U19056 (N_19056,N_11627,N_14100);
and U19057 (N_19057,N_13502,N_13948);
and U19058 (N_19058,N_13258,N_14637);
or U19059 (N_19059,N_13800,N_10844);
and U19060 (N_19060,N_11528,N_10541);
nand U19061 (N_19061,N_13502,N_13052);
xor U19062 (N_19062,N_10746,N_13213);
xor U19063 (N_19063,N_14095,N_11141);
nor U19064 (N_19064,N_12277,N_14868);
xnor U19065 (N_19065,N_10569,N_14086);
xor U19066 (N_19066,N_11029,N_12068);
and U19067 (N_19067,N_12341,N_12752);
or U19068 (N_19068,N_12901,N_10602);
xnor U19069 (N_19069,N_12070,N_12552);
and U19070 (N_19070,N_11000,N_10073);
nor U19071 (N_19071,N_13360,N_13362);
or U19072 (N_19072,N_13213,N_11263);
nand U19073 (N_19073,N_14426,N_12775);
nor U19074 (N_19074,N_14541,N_13569);
xnor U19075 (N_19075,N_12627,N_13715);
and U19076 (N_19076,N_13144,N_11009);
xor U19077 (N_19077,N_14403,N_13378);
xor U19078 (N_19078,N_11820,N_11471);
xnor U19079 (N_19079,N_10663,N_14766);
nor U19080 (N_19080,N_12124,N_14124);
and U19081 (N_19081,N_13026,N_12748);
or U19082 (N_19082,N_10130,N_10411);
nor U19083 (N_19083,N_12318,N_10440);
or U19084 (N_19084,N_12532,N_10807);
nor U19085 (N_19085,N_13891,N_12828);
or U19086 (N_19086,N_11150,N_14104);
nand U19087 (N_19087,N_13265,N_13914);
nand U19088 (N_19088,N_13789,N_10513);
and U19089 (N_19089,N_14557,N_11884);
or U19090 (N_19090,N_10182,N_14535);
nand U19091 (N_19091,N_12124,N_10214);
nand U19092 (N_19092,N_14116,N_13552);
or U19093 (N_19093,N_10657,N_11997);
nor U19094 (N_19094,N_13621,N_14159);
nor U19095 (N_19095,N_12509,N_10549);
or U19096 (N_19096,N_14617,N_12601);
xor U19097 (N_19097,N_10267,N_13472);
nand U19098 (N_19098,N_13028,N_10006);
xor U19099 (N_19099,N_13923,N_11993);
nor U19100 (N_19100,N_13197,N_12803);
nand U19101 (N_19101,N_11863,N_13579);
xor U19102 (N_19102,N_14798,N_10086);
or U19103 (N_19103,N_13701,N_11560);
nand U19104 (N_19104,N_13521,N_11962);
nand U19105 (N_19105,N_14203,N_11201);
nor U19106 (N_19106,N_10768,N_11237);
nor U19107 (N_19107,N_14761,N_14139);
or U19108 (N_19108,N_14621,N_11322);
xnor U19109 (N_19109,N_11909,N_12008);
nand U19110 (N_19110,N_12338,N_14228);
and U19111 (N_19111,N_12989,N_14838);
nand U19112 (N_19112,N_13487,N_14466);
nor U19113 (N_19113,N_14223,N_14706);
and U19114 (N_19114,N_12174,N_14486);
xor U19115 (N_19115,N_10530,N_14647);
nand U19116 (N_19116,N_10952,N_12146);
xnor U19117 (N_19117,N_14777,N_11184);
xnor U19118 (N_19118,N_11475,N_13849);
nor U19119 (N_19119,N_12595,N_10468);
nor U19120 (N_19120,N_12805,N_14113);
nor U19121 (N_19121,N_10534,N_13455);
and U19122 (N_19122,N_13350,N_11231);
xor U19123 (N_19123,N_10807,N_13291);
and U19124 (N_19124,N_13373,N_10596);
and U19125 (N_19125,N_10007,N_12363);
nand U19126 (N_19126,N_11344,N_14980);
and U19127 (N_19127,N_10237,N_11838);
nand U19128 (N_19128,N_14540,N_11080);
and U19129 (N_19129,N_12099,N_13090);
or U19130 (N_19130,N_13459,N_13027);
xor U19131 (N_19131,N_12659,N_10641);
nand U19132 (N_19132,N_12226,N_13975);
and U19133 (N_19133,N_12901,N_13141);
nand U19134 (N_19134,N_11114,N_10040);
nor U19135 (N_19135,N_12578,N_13034);
or U19136 (N_19136,N_12633,N_14821);
or U19137 (N_19137,N_11133,N_10943);
or U19138 (N_19138,N_11599,N_13476);
or U19139 (N_19139,N_12500,N_14823);
xor U19140 (N_19140,N_10620,N_14512);
xnor U19141 (N_19141,N_13883,N_13360);
xnor U19142 (N_19142,N_10561,N_14865);
nand U19143 (N_19143,N_10036,N_14487);
nand U19144 (N_19144,N_10475,N_11178);
nand U19145 (N_19145,N_14659,N_11103);
and U19146 (N_19146,N_13088,N_12001);
nand U19147 (N_19147,N_13187,N_10293);
xnor U19148 (N_19148,N_14164,N_14690);
and U19149 (N_19149,N_12293,N_10709);
nand U19150 (N_19150,N_12242,N_13746);
and U19151 (N_19151,N_12281,N_13104);
and U19152 (N_19152,N_14183,N_11784);
nor U19153 (N_19153,N_10458,N_13337);
nand U19154 (N_19154,N_11659,N_11051);
nor U19155 (N_19155,N_10519,N_12372);
xor U19156 (N_19156,N_14163,N_10952);
and U19157 (N_19157,N_12566,N_14947);
nor U19158 (N_19158,N_14824,N_11926);
nand U19159 (N_19159,N_14852,N_12414);
and U19160 (N_19160,N_13496,N_11980);
xnor U19161 (N_19161,N_14065,N_11972);
nand U19162 (N_19162,N_10253,N_12147);
and U19163 (N_19163,N_10471,N_13432);
xnor U19164 (N_19164,N_10030,N_10252);
nand U19165 (N_19165,N_14112,N_12904);
xor U19166 (N_19166,N_13301,N_10090);
nand U19167 (N_19167,N_11909,N_12233);
and U19168 (N_19168,N_10277,N_10786);
or U19169 (N_19169,N_12338,N_14763);
or U19170 (N_19170,N_13790,N_13851);
nor U19171 (N_19171,N_14771,N_11897);
or U19172 (N_19172,N_14400,N_11070);
nand U19173 (N_19173,N_11077,N_10193);
xor U19174 (N_19174,N_13446,N_10463);
and U19175 (N_19175,N_10011,N_12718);
nor U19176 (N_19176,N_11926,N_11144);
nor U19177 (N_19177,N_13152,N_11747);
nand U19178 (N_19178,N_10781,N_13093);
nor U19179 (N_19179,N_14599,N_14744);
or U19180 (N_19180,N_13872,N_10425);
xor U19181 (N_19181,N_14157,N_10446);
and U19182 (N_19182,N_12270,N_12638);
nand U19183 (N_19183,N_12578,N_13991);
nand U19184 (N_19184,N_14025,N_10667);
or U19185 (N_19185,N_10903,N_13588);
nand U19186 (N_19186,N_11457,N_13968);
or U19187 (N_19187,N_13876,N_13986);
nor U19188 (N_19188,N_10796,N_10729);
and U19189 (N_19189,N_10433,N_11702);
nand U19190 (N_19190,N_11587,N_12125);
nor U19191 (N_19191,N_13012,N_13242);
nand U19192 (N_19192,N_11388,N_11378);
nor U19193 (N_19193,N_14364,N_11028);
or U19194 (N_19194,N_12051,N_13900);
nor U19195 (N_19195,N_13681,N_11271);
xnor U19196 (N_19196,N_13195,N_11600);
or U19197 (N_19197,N_13223,N_12860);
or U19198 (N_19198,N_14351,N_13420);
xnor U19199 (N_19199,N_12474,N_13776);
nand U19200 (N_19200,N_11468,N_13604);
nor U19201 (N_19201,N_10258,N_11331);
or U19202 (N_19202,N_10674,N_14849);
nor U19203 (N_19203,N_13103,N_14685);
nand U19204 (N_19204,N_10777,N_14783);
xor U19205 (N_19205,N_10311,N_10822);
and U19206 (N_19206,N_11340,N_13440);
xnor U19207 (N_19207,N_10601,N_12142);
and U19208 (N_19208,N_12957,N_12297);
or U19209 (N_19209,N_11230,N_10432);
nand U19210 (N_19210,N_14295,N_11407);
xor U19211 (N_19211,N_12540,N_10543);
or U19212 (N_19212,N_12187,N_12829);
nor U19213 (N_19213,N_11133,N_10284);
nand U19214 (N_19214,N_14413,N_13434);
xor U19215 (N_19215,N_13206,N_10976);
and U19216 (N_19216,N_11050,N_11132);
nand U19217 (N_19217,N_14484,N_13524);
nor U19218 (N_19218,N_14181,N_11227);
and U19219 (N_19219,N_14153,N_10615);
and U19220 (N_19220,N_13404,N_12911);
nor U19221 (N_19221,N_13523,N_14641);
nand U19222 (N_19222,N_10064,N_12206);
and U19223 (N_19223,N_14875,N_12660);
xnor U19224 (N_19224,N_14750,N_14764);
and U19225 (N_19225,N_14889,N_12154);
nor U19226 (N_19226,N_12674,N_12768);
nand U19227 (N_19227,N_11409,N_10915);
xnor U19228 (N_19228,N_11935,N_14070);
nor U19229 (N_19229,N_11120,N_12133);
xor U19230 (N_19230,N_13691,N_11486);
xor U19231 (N_19231,N_14491,N_12910);
and U19232 (N_19232,N_11475,N_13981);
or U19233 (N_19233,N_13465,N_10827);
or U19234 (N_19234,N_11677,N_10422);
nand U19235 (N_19235,N_12589,N_10654);
xor U19236 (N_19236,N_13272,N_14689);
or U19237 (N_19237,N_10378,N_12904);
xor U19238 (N_19238,N_12878,N_11173);
nand U19239 (N_19239,N_10881,N_12591);
and U19240 (N_19240,N_12830,N_13320);
xnor U19241 (N_19241,N_12356,N_14932);
and U19242 (N_19242,N_11390,N_13241);
nor U19243 (N_19243,N_11175,N_10760);
or U19244 (N_19244,N_11985,N_14833);
nand U19245 (N_19245,N_10505,N_10553);
xor U19246 (N_19246,N_12291,N_12085);
nor U19247 (N_19247,N_11772,N_11030);
nor U19248 (N_19248,N_12353,N_12781);
and U19249 (N_19249,N_10904,N_14536);
nand U19250 (N_19250,N_14668,N_11980);
nor U19251 (N_19251,N_11176,N_11954);
or U19252 (N_19252,N_14815,N_13515);
or U19253 (N_19253,N_11039,N_10224);
nand U19254 (N_19254,N_10947,N_13343);
nand U19255 (N_19255,N_11410,N_12652);
nand U19256 (N_19256,N_12081,N_12833);
nand U19257 (N_19257,N_14294,N_14871);
nand U19258 (N_19258,N_13305,N_10915);
or U19259 (N_19259,N_11528,N_11787);
and U19260 (N_19260,N_12957,N_11119);
or U19261 (N_19261,N_14170,N_10371);
nand U19262 (N_19262,N_13006,N_12327);
xor U19263 (N_19263,N_13167,N_14379);
nor U19264 (N_19264,N_12438,N_13828);
nand U19265 (N_19265,N_11855,N_13735);
xnor U19266 (N_19266,N_14880,N_10178);
nor U19267 (N_19267,N_12686,N_14470);
and U19268 (N_19268,N_11909,N_14979);
nand U19269 (N_19269,N_14596,N_10940);
nor U19270 (N_19270,N_12302,N_10512);
and U19271 (N_19271,N_11703,N_10435);
nor U19272 (N_19272,N_10482,N_10580);
or U19273 (N_19273,N_10349,N_10743);
xor U19274 (N_19274,N_13946,N_10836);
xor U19275 (N_19275,N_13371,N_14072);
nor U19276 (N_19276,N_10587,N_13090);
nor U19277 (N_19277,N_10298,N_10967);
nor U19278 (N_19278,N_10798,N_10147);
or U19279 (N_19279,N_11002,N_13708);
and U19280 (N_19280,N_12965,N_13950);
or U19281 (N_19281,N_10721,N_10201);
nand U19282 (N_19282,N_13976,N_11258);
and U19283 (N_19283,N_14371,N_10677);
xnor U19284 (N_19284,N_14886,N_11990);
nand U19285 (N_19285,N_13697,N_12379);
nor U19286 (N_19286,N_12377,N_14298);
nand U19287 (N_19287,N_10923,N_14538);
nor U19288 (N_19288,N_12453,N_13111);
nor U19289 (N_19289,N_12521,N_10531);
nor U19290 (N_19290,N_13731,N_10093);
xnor U19291 (N_19291,N_14980,N_11643);
nand U19292 (N_19292,N_11792,N_11994);
xor U19293 (N_19293,N_14583,N_12942);
xor U19294 (N_19294,N_12799,N_12987);
or U19295 (N_19295,N_11034,N_13307);
or U19296 (N_19296,N_10854,N_14837);
nor U19297 (N_19297,N_12559,N_10155);
or U19298 (N_19298,N_13833,N_13097);
nor U19299 (N_19299,N_11504,N_11862);
xnor U19300 (N_19300,N_10098,N_11106);
or U19301 (N_19301,N_12247,N_14300);
nand U19302 (N_19302,N_14646,N_14127);
or U19303 (N_19303,N_12777,N_12436);
or U19304 (N_19304,N_10362,N_14888);
nand U19305 (N_19305,N_12461,N_14622);
nor U19306 (N_19306,N_11882,N_11613);
and U19307 (N_19307,N_12848,N_12126);
nand U19308 (N_19308,N_13204,N_11940);
and U19309 (N_19309,N_14096,N_11446);
or U19310 (N_19310,N_10623,N_13699);
xor U19311 (N_19311,N_12781,N_12027);
nand U19312 (N_19312,N_12659,N_14804);
nor U19313 (N_19313,N_12816,N_13257);
nor U19314 (N_19314,N_14846,N_14804);
nand U19315 (N_19315,N_12741,N_13697);
nand U19316 (N_19316,N_14390,N_14388);
xnor U19317 (N_19317,N_13684,N_14649);
nor U19318 (N_19318,N_12738,N_14329);
and U19319 (N_19319,N_14682,N_12444);
nand U19320 (N_19320,N_11474,N_10960);
and U19321 (N_19321,N_11797,N_14979);
and U19322 (N_19322,N_10133,N_13371);
nand U19323 (N_19323,N_14364,N_12646);
xor U19324 (N_19324,N_11669,N_11220);
xor U19325 (N_19325,N_11480,N_12540);
and U19326 (N_19326,N_11887,N_13672);
nand U19327 (N_19327,N_13329,N_12460);
nand U19328 (N_19328,N_14527,N_14560);
nand U19329 (N_19329,N_13763,N_12671);
nor U19330 (N_19330,N_14328,N_14241);
nand U19331 (N_19331,N_12159,N_12024);
and U19332 (N_19332,N_10412,N_13935);
nor U19333 (N_19333,N_11273,N_13009);
nand U19334 (N_19334,N_12758,N_13590);
and U19335 (N_19335,N_13831,N_13556);
xnor U19336 (N_19336,N_13182,N_14297);
or U19337 (N_19337,N_13698,N_10477);
or U19338 (N_19338,N_12677,N_10923);
xnor U19339 (N_19339,N_13959,N_14325);
xor U19340 (N_19340,N_11733,N_11635);
or U19341 (N_19341,N_13508,N_12070);
nor U19342 (N_19342,N_12147,N_12918);
or U19343 (N_19343,N_11970,N_10176);
nor U19344 (N_19344,N_11004,N_13239);
nand U19345 (N_19345,N_12578,N_13153);
xnor U19346 (N_19346,N_11988,N_13546);
nand U19347 (N_19347,N_13706,N_14415);
nand U19348 (N_19348,N_13821,N_13798);
xor U19349 (N_19349,N_14664,N_14707);
and U19350 (N_19350,N_13459,N_11510);
xor U19351 (N_19351,N_12896,N_11664);
nor U19352 (N_19352,N_14600,N_13494);
and U19353 (N_19353,N_14220,N_13536);
nor U19354 (N_19354,N_11784,N_12096);
nand U19355 (N_19355,N_12402,N_10074);
or U19356 (N_19356,N_13522,N_13385);
and U19357 (N_19357,N_11838,N_12989);
and U19358 (N_19358,N_11764,N_13102);
xnor U19359 (N_19359,N_11111,N_14653);
and U19360 (N_19360,N_10522,N_11294);
and U19361 (N_19361,N_14520,N_14349);
nor U19362 (N_19362,N_13370,N_13202);
or U19363 (N_19363,N_13734,N_13580);
nor U19364 (N_19364,N_11431,N_12573);
xnor U19365 (N_19365,N_14671,N_10624);
and U19366 (N_19366,N_14814,N_12667);
and U19367 (N_19367,N_11032,N_14876);
nand U19368 (N_19368,N_11807,N_10153);
xor U19369 (N_19369,N_14382,N_13331);
nand U19370 (N_19370,N_13680,N_13323);
nand U19371 (N_19371,N_14620,N_11520);
nor U19372 (N_19372,N_10109,N_11087);
and U19373 (N_19373,N_10157,N_13240);
or U19374 (N_19374,N_10366,N_10947);
nand U19375 (N_19375,N_13261,N_14889);
nand U19376 (N_19376,N_10639,N_12724);
nor U19377 (N_19377,N_12083,N_14301);
nand U19378 (N_19378,N_12690,N_14836);
and U19379 (N_19379,N_14142,N_13359);
nand U19380 (N_19380,N_10372,N_13255);
and U19381 (N_19381,N_11982,N_10871);
and U19382 (N_19382,N_14144,N_10495);
xnor U19383 (N_19383,N_11631,N_12900);
and U19384 (N_19384,N_10947,N_12315);
or U19385 (N_19385,N_12351,N_11621);
xnor U19386 (N_19386,N_10565,N_12698);
xor U19387 (N_19387,N_10426,N_12798);
nor U19388 (N_19388,N_11758,N_12776);
or U19389 (N_19389,N_14987,N_13051);
and U19390 (N_19390,N_13088,N_10630);
xnor U19391 (N_19391,N_13695,N_13608);
xnor U19392 (N_19392,N_13380,N_14207);
and U19393 (N_19393,N_14369,N_10202);
nand U19394 (N_19394,N_10520,N_13977);
nor U19395 (N_19395,N_14480,N_10398);
nor U19396 (N_19396,N_10826,N_14060);
xnor U19397 (N_19397,N_11278,N_11843);
and U19398 (N_19398,N_11308,N_14348);
nand U19399 (N_19399,N_11294,N_14452);
nor U19400 (N_19400,N_13834,N_12900);
nor U19401 (N_19401,N_12848,N_10708);
nand U19402 (N_19402,N_14966,N_11032);
xor U19403 (N_19403,N_13045,N_11709);
xnor U19404 (N_19404,N_12194,N_14136);
nand U19405 (N_19405,N_14507,N_14610);
and U19406 (N_19406,N_10067,N_12263);
xnor U19407 (N_19407,N_13631,N_11902);
nor U19408 (N_19408,N_14311,N_14064);
nor U19409 (N_19409,N_10345,N_11069);
xnor U19410 (N_19410,N_10672,N_10683);
xnor U19411 (N_19411,N_12683,N_10920);
and U19412 (N_19412,N_11029,N_13511);
xor U19413 (N_19413,N_12343,N_12852);
or U19414 (N_19414,N_10535,N_14999);
xnor U19415 (N_19415,N_11002,N_13039);
and U19416 (N_19416,N_12121,N_12165);
or U19417 (N_19417,N_10656,N_14979);
and U19418 (N_19418,N_14381,N_14090);
xor U19419 (N_19419,N_10879,N_13329);
or U19420 (N_19420,N_13814,N_14321);
nand U19421 (N_19421,N_11524,N_13219);
nor U19422 (N_19422,N_14061,N_13137);
nand U19423 (N_19423,N_11608,N_10654);
nor U19424 (N_19424,N_10356,N_12540);
nor U19425 (N_19425,N_14819,N_14900);
nor U19426 (N_19426,N_12980,N_13869);
xor U19427 (N_19427,N_11012,N_10969);
and U19428 (N_19428,N_13183,N_12830);
nor U19429 (N_19429,N_14271,N_13337);
or U19430 (N_19430,N_11471,N_12781);
nor U19431 (N_19431,N_10702,N_11229);
nor U19432 (N_19432,N_13105,N_13683);
or U19433 (N_19433,N_12716,N_11482);
nand U19434 (N_19434,N_14397,N_14380);
and U19435 (N_19435,N_10907,N_10305);
nor U19436 (N_19436,N_12371,N_14941);
and U19437 (N_19437,N_13456,N_12410);
nand U19438 (N_19438,N_14276,N_12708);
nand U19439 (N_19439,N_12442,N_12623);
nand U19440 (N_19440,N_12076,N_12031);
or U19441 (N_19441,N_14170,N_14056);
and U19442 (N_19442,N_12560,N_11612);
or U19443 (N_19443,N_10215,N_12145);
nand U19444 (N_19444,N_13221,N_11871);
nand U19445 (N_19445,N_13017,N_12305);
xor U19446 (N_19446,N_10311,N_10863);
and U19447 (N_19447,N_12001,N_10869);
nand U19448 (N_19448,N_14533,N_11245);
nor U19449 (N_19449,N_11456,N_11841);
xor U19450 (N_19450,N_12370,N_11547);
nor U19451 (N_19451,N_13868,N_13465);
nand U19452 (N_19452,N_10302,N_10691);
xnor U19453 (N_19453,N_13728,N_10394);
xor U19454 (N_19454,N_14569,N_14818);
and U19455 (N_19455,N_13881,N_12865);
and U19456 (N_19456,N_14683,N_10137);
or U19457 (N_19457,N_10863,N_14352);
xnor U19458 (N_19458,N_11584,N_11225);
and U19459 (N_19459,N_11141,N_11836);
nor U19460 (N_19460,N_10797,N_11904);
nand U19461 (N_19461,N_11502,N_10498);
nand U19462 (N_19462,N_10354,N_10851);
xnor U19463 (N_19463,N_13232,N_13025);
or U19464 (N_19464,N_10746,N_14665);
xor U19465 (N_19465,N_12595,N_11472);
xor U19466 (N_19466,N_14779,N_11196);
or U19467 (N_19467,N_14644,N_12871);
nand U19468 (N_19468,N_14368,N_12182);
or U19469 (N_19469,N_12222,N_13746);
or U19470 (N_19470,N_12905,N_12015);
xnor U19471 (N_19471,N_14194,N_11219);
or U19472 (N_19472,N_13672,N_13623);
nor U19473 (N_19473,N_12422,N_11731);
and U19474 (N_19474,N_11194,N_12939);
nand U19475 (N_19475,N_10497,N_13746);
xor U19476 (N_19476,N_14439,N_14823);
nand U19477 (N_19477,N_13435,N_10239);
nor U19478 (N_19478,N_13864,N_13209);
nand U19479 (N_19479,N_10683,N_11931);
and U19480 (N_19480,N_12054,N_13103);
and U19481 (N_19481,N_11054,N_11229);
nor U19482 (N_19482,N_13252,N_11637);
nand U19483 (N_19483,N_14774,N_10949);
or U19484 (N_19484,N_11886,N_12134);
nor U19485 (N_19485,N_10120,N_11647);
nand U19486 (N_19486,N_12345,N_11385);
nor U19487 (N_19487,N_14711,N_14812);
or U19488 (N_19488,N_14036,N_14662);
xor U19489 (N_19489,N_14657,N_12263);
or U19490 (N_19490,N_13276,N_12356);
and U19491 (N_19491,N_14728,N_13395);
or U19492 (N_19492,N_13801,N_12135);
and U19493 (N_19493,N_12579,N_13534);
xor U19494 (N_19494,N_10829,N_11728);
nand U19495 (N_19495,N_10310,N_11229);
or U19496 (N_19496,N_14030,N_14288);
or U19497 (N_19497,N_10171,N_13845);
nand U19498 (N_19498,N_14220,N_14620);
and U19499 (N_19499,N_12717,N_13588);
xor U19500 (N_19500,N_10572,N_14379);
xor U19501 (N_19501,N_14562,N_10026);
nand U19502 (N_19502,N_12077,N_11114);
or U19503 (N_19503,N_10030,N_10864);
nor U19504 (N_19504,N_10483,N_10566);
and U19505 (N_19505,N_13944,N_12364);
nor U19506 (N_19506,N_10458,N_14747);
and U19507 (N_19507,N_10124,N_10297);
and U19508 (N_19508,N_11391,N_11684);
nor U19509 (N_19509,N_12434,N_10837);
xnor U19510 (N_19510,N_10368,N_13196);
nor U19511 (N_19511,N_10553,N_13336);
and U19512 (N_19512,N_13345,N_10739);
or U19513 (N_19513,N_12347,N_10074);
xor U19514 (N_19514,N_13169,N_12081);
nand U19515 (N_19515,N_13027,N_12439);
or U19516 (N_19516,N_12926,N_10351);
nor U19517 (N_19517,N_11595,N_10331);
and U19518 (N_19518,N_14607,N_14054);
nand U19519 (N_19519,N_13370,N_11037);
xor U19520 (N_19520,N_10566,N_10541);
nand U19521 (N_19521,N_10101,N_11236);
xor U19522 (N_19522,N_11341,N_10818);
nand U19523 (N_19523,N_14118,N_11752);
xor U19524 (N_19524,N_13446,N_10902);
nor U19525 (N_19525,N_13352,N_14680);
or U19526 (N_19526,N_10830,N_12505);
or U19527 (N_19527,N_11026,N_14334);
or U19528 (N_19528,N_13731,N_12516);
nor U19529 (N_19529,N_13813,N_14586);
nand U19530 (N_19530,N_11969,N_10819);
and U19531 (N_19531,N_13336,N_14232);
and U19532 (N_19532,N_13076,N_10537);
and U19533 (N_19533,N_10712,N_11772);
nor U19534 (N_19534,N_10637,N_13018);
or U19535 (N_19535,N_11462,N_14849);
nand U19536 (N_19536,N_12490,N_13938);
and U19537 (N_19537,N_11809,N_10285);
nand U19538 (N_19538,N_13657,N_11934);
xnor U19539 (N_19539,N_14190,N_10736);
xnor U19540 (N_19540,N_14699,N_12392);
nor U19541 (N_19541,N_14368,N_14942);
xor U19542 (N_19542,N_14020,N_13526);
and U19543 (N_19543,N_10437,N_13754);
and U19544 (N_19544,N_11102,N_14937);
or U19545 (N_19545,N_12624,N_14180);
xnor U19546 (N_19546,N_10901,N_11300);
and U19547 (N_19547,N_12381,N_13538);
and U19548 (N_19548,N_10890,N_13954);
nand U19549 (N_19549,N_11124,N_10725);
nand U19550 (N_19550,N_11188,N_12673);
or U19551 (N_19551,N_13414,N_12306);
nor U19552 (N_19552,N_14910,N_13515);
or U19553 (N_19553,N_10699,N_13088);
xnor U19554 (N_19554,N_10418,N_14265);
or U19555 (N_19555,N_11206,N_12645);
or U19556 (N_19556,N_13822,N_11458);
nor U19557 (N_19557,N_12693,N_14035);
or U19558 (N_19558,N_13879,N_13554);
and U19559 (N_19559,N_14024,N_13386);
xnor U19560 (N_19560,N_10731,N_12959);
and U19561 (N_19561,N_12280,N_11629);
nand U19562 (N_19562,N_13786,N_10837);
xnor U19563 (N_19563,N_13715,N_14275);
nor U19564 (N_19564,N_10207,N_12023);
nor U19565 (N_19565,N_10588,N_13007);
nor U19566 (N_19566,N_13969,N_14569);
or U19567 (N_19567,N_12183,N_11633);
nor U19568 (N_19568,N_14729,N_14124);
nand U19569 (N_19569,N_12093,N_13465);
and U19570 (N_19570,N_13703,N_12881);
and U19571 (N_19571,N_14248,N_11741);
xnor U19572 (N_19572,N_14313,N_11464);
and U19573 (N_19573,N_11936,N_10296);
or U19574 (N_19574,N_11323,N_14765);
or U19575 (N_19575,N_14370,N_10088);
nand U19576 (N_19576,N_11212,N_10506);
and U19577 (N_19577,N_14822,N_13686);
and U19578 (N_19578,N_11240,N_13554);
or U19579 (N_19579,N_10521,N_11801);
and U19580 (N_19580,N_10446,N_11923);
and U19581 (N_19581,N_12605,N_10257);
nor U19582 (N_19582,N_12689,N_10610);
nand U19583 (N_19583,N_11310,N_14028);
or U19584 (N_19584,N_14689,N_12752);
nor U19585 (N_19585,N_13383,N_11812);
xor U19586 (N_19586,N_14646,N_11728);
xor U19587 (N_19587,N_14423,N_10800);
and U19588 (N_19588,N_13726,N_11302);
and U19589 (N_19589,N_14128,N_10812);
or U19590 (N_19590,N_12925,N_11206);
nand U19591 (N_19591,N_11361,N_11360);
xnor U19592 (N_19592,N_14802,N_10939);
xor U19593 (N_19593,N_13325,N_12223);
or U19594 (N_19594,N_14025,N_13957);
nand U19595 (N_19595,N_10984,N_13080);
nand U19596 (N_19596,N_14163,N_10964);
nor U19597 (N_19597,N_11073,N_13643);
xnor U19598 (N_19598,N_14311,N_13023);
or U19599 (N_19599,N_14368,N_13163);
nand U19600 (N_19600,N_13735,N_12099);
nand U19601 (N_19601,N_10790,N_14245);
nor U19602 (N_19602,N_10322,N_14268);
xnor U19603 (N_19603,N_10937,N_12706);
nand U19604 (N_19604,N_14465,N_10999);
xor U19605 (N_19605,N_12219,N_13175);
and U19606 (N_19606,N_12263,N_13921);
nor U19607 (N_19607,N_12892,N_10433);
or U19608 (N_19608,N_12812,N_10219);
or U19609 (N_19609,N_14692,N_10827);
nand U19610 (N_19610,N_10799,N_13489);
or U19611 (N_19611,N_10943,N_11077);
and U19612 (N_19612,N_10385,N_13293);
nor U19613 (N_19613,N_14243,N_14664);
nand U19614 (N_19614,N_14310,N_14829);
nand U19615 (N_19615,N_11815,N_11549);
and U19616 (N_19616,N_12886,N_11629);
nand U19617 (N_19617,N_11815,N_13895);
nor U19618 (N_19618,N_14542,N_10315);
nand U19619 (N_19619,N_13156,N_10405);
nand U19620 (N_19620,N_13904,N_11683);
or U19621 (N_19621,N_11447,N_14435);
nor U19622 (N_19622,N_11125,N_10759);
and U19623 (N_19623,N_12989,N_12236);
nor U19624 (N_19624,N_10119,N_13582);
and U19625 (N_19625,N_12997,N_14923);
or U19626 (N_19626,N_11026,N_11456);
and U19627 (N_19627,N_13657,N_11900);
and U19628 (N_19628,N_10504,N_14505);
or U19629 (N_19629,N_13901,N_11042);
and U19630 (N_19630,N_10652,N_10092);
and U19631 (N_19631,N_10395,N_13720);
or U19632 (N_19632,N_13025,N_13514);
nand U19633 (N_19633,N_14080,N_12837);
and U19634 (N_19634,N_10540,N_12476);
xor U19635 (N_19635,N_13201,N_14783);
nor U19636 (N_19636,N_13729,N_11943);
or U19637 (N_19637,N_11000,N_12059);
and U19638 (N_19638,N_14983,N_14160);
and U19639 (N_19639,N_13360,N_12884);
or U19640 (N_19640,N_11829,N_13013);
xnor U19641 (N_19641,N_11456,N_14127);
nand U19642 (N_19642,N_13101,N_12810);
or U19643 (N_19643,N_14321,N_13252);
nand U19644 (N_19644,N_13639,N_14176);
xor U19645 (N_19645,N_11450,N_12567);
nand U19646 (N_19646,N_13481,N_12310);
nor U19647 (N_19647,N_11800,N_11344);
xor U19648 (N_19648,N_13207,N_10603);
nor U19649 (N_19649,N_13865,N_14809);
xnor U19650 (N_19650,N_13142,N_11276);
nand U19651 (N_19651,N_13436,N_14451);
and U19652 (N_19652,N_14230,N_14933);
or U19653 (N_19653,N_10861,N_12260);
and U19654 (N_19654,N_11792,N_10582);
xor U19655 (N_19655,N_10842,N_13595);
or U19656 (N_19656,N_13758,N_11504);
and U19657 (N_19657,N_11897,N_11044);
or U19658 (N_19658,N_13905,N_11130);
xnor U19659 (N_19659,N_11533,N_14035);
nor U19660 (N_19660,N_12211,N_14663);
xor U19661 (N_19661,N_12660,N_12081);
nor U19662 (N_19662,N_14564,N_11935);
or U19663 (N_19663,N_14052,N_14075);
xor U19664 (N_19664,N_13957,N_12606);
and U19665 (N_19665,N_11623,N_12336);
nand U19666 (N_19666,N_13870,N_10003);
xnor U19667 (N_19667,N_10079,N_10690);
or U19668 (N_19668,N_11976,N_14963);
xor U19669 (N_19669,N_14429,N_10347);
or U19670 (N_19670,N_11099,N_14325);
nand U19671 (N_19671,N_13074,N_13423);
or U19672 (N_19672,N_11848,N_14729);
nor U19673 (N_19673,N_12518,N_14400);
and U19674 (N_19674,N_12239,N_14327);
or U19675 (N_19675,N_14218,N_12899);
and U19676 (N_19676,N_12383,N_11564);
or U19677 (N_19677,N_13601,N_12413);
nand U19678 (N_19678,N_12248,N_13240);
and U19679 (N_19679,N_14790,N_11272);
nor U19680 (N_19680,N_11799,N_11977);
nand U19681 (N_19681,N_11627,N_12233);
xor U19682 (N_19682,N_11383,N_12658);
nand U19683 (N_19683,N_14408,N_13468);
or U19684 (N_19684,N_13264,N_10231);
and U19685 (N_19685,N_14444,N_14656);
xor U19686 (N_19686,N_11308,N_14582);
nand U19687 (N_19687,N_11934,N_11714);
nor U19688 (N_19688,N_12126,N_13000);
or U19689 (N_19689,N_12848,N_10982);
nor U19690 (N_19690,N_14866,N_14039);
xnor U19691 (N_19691,N_13819,N_12161);
or U19692 (N_19692,N_12025,N_12891);
and U19693 (N_19693,N_10484,N_13146);
xor U19694 (N_19694,N_12190,N_13212);
nor U19695 (N_19695,N_11795,N_11048);
nor U19696 (N_19696,N_13780,N_14162);
xnor U19697 (N_19697,N_12932,N_11977);
nand U19698 (N_19698,N_11174,N_14819);
xnor U19699 (N_19699,N_12399,N_13254);
or U19700 (N_19700,N_11243,N_14202);
or U19701 (N_19701,N_13795,N_14641);
nor U19702 (N_19702,N_11356,N_11672);
nor U19703 (N_19703,N_10318,N_12111);
nor U19704 (N_19704,N_13045,N_12206);
nand U19705 (N_19705,N_14345,N_12560);
or U19706 (N_19706,N_11514,N_12910);
nor U19707 (N_19707,N_10288,N_10797);
nor U19708 (N_19708,N_13817,N_10677);
or U19709 (N_19709,N_10035,N_13167);
nor U19710 (N_19710,N_12183,N_10973);
nand U19711 (N_19711,N_11429,N_14631);
xnor U19712 (N_19712,N_13347,N_13184);
and U19713 (N_19713,N_12345,N_13038);
xnor U19714 (N_19714,N_10351,N_14878);
nand U19715 (N_19715,N_14004,N_11489);
nand U19716 (N_19716,N_10416,N_12157);
nor U19717 (N_19717,N_13236,N_10872);
nand U19718 (N_19718,N_10060,N_14237);
xnor U19719 (N_19719,N_12870,N_13584);
or U19720 (N_19720,N_12979,N_11779);
nand U19721 (N_19721,N_10819,N_11769);
or U19722 (N_19722,N_13439,N_13888);
or U19723 (N_19723,N_12455,N_14498);
xnor U19724 (N_19724,N_13720,N_14660);
nor U19725 (N_19725,N_10254,N_11222);
xnor U19726 (N_19726,N_10684,N_10221);
nor U19727 (N_19727,N_14479,N_13408);
nand U19728 (N_19728,N_11363,N_11990);
xor U19729 (N_19729,N_11909,N_10813);
nor U19730 (N_19730,N_13515,N_14701);
nand U19731 (N_19731,N_11217,N_10621);
and U19732 (N_19732,N_14897,N_14603);
xor U19733 (N_19733,N_13576,N_11287);
or U19734 (N_19734,N_14039,N_14755);
xnor U19735 (N_19735,N_11213,N_13183);
and U19736 (N_19736,N_10369,N_14587);
and U19737 (N_19737,N_13806,N_13723);
or U19738 (N_19738,N_11298,N_13143);
and U19739 (N_19739,N_13024,N_12059);
xnor U19740 (N_19740,N_11057,N_10961);
and U19741 (N_19741,N_12724,N_12674);
nand U19742 (N_19742,N_12488,N_14824);
and U19743 (N_19743,N_12890,N_14016);
xor U19744 (N_19744,N_13576,N_14327);
nor U19745 (N_19745,N_14740,N_14977);
nor U19746 (N_19746,N_12264,N_14282);
nand U19747 (N_19747,N_13880,N_10472);
or U19748 (N_19748,N_14005,N_14327);
or U19749 (N_19749,N_13559,N_11860);
nor U19750 (N_19750,N_11739,N_10302);
nand U19751 (N_19751,N_13178,N_11051);
xor U19752 (N_19752,N_12433,N_10539);
nand U19753 (N_19753,N_13755,N_13904);
or U19754 (N_19754,N_12304,N_11350);
or U19755 (N_19755,N_11782,N_11386);
or U19756 (N_19756,N_12923,N_12409);
nand U19757 (N_19757,N_10953,N_12826);
and U19758 (N_19758,N_12716,N_11593);
nand U19759 (N_19759,N_14500,N_12221);
and U19760 (N_19760,N_11121,N_11666);
nand U19761 (N_19761,N_10424,N_14513);
nor U19762 (N_19762,N_12738,N_14272);
nand U19763 (N_19763,N_10737,N_10486);
xor U19764 (N_19764,N_10838,N_10751);
nand U19765 (N_19765,N_11455,N_11641);
nor U19766 (N_19766,N_14621,N_13066);
and U19767 (N_19767,N_13334,N_10575);
nand U19768 (N_19768,N_12473,N_14095);
or U19769 (N_19769,N_12430,N_11719);
and U19770 (N_19770,N_13756,N_10534);
and U19771 (N_19771,N_12261,N_11442);
nor U19772 (N_19772,N_11954,N_11273);
xor U19773 (N_19773,N_14898,N_14128);
nand U19774 (N_19774,N_14619,N_10806);
nor U19775 (N_19775,N_14379,N_14727);
and U19776 (N_19776,N_13115,N_13781);
or U19777 (N_19777,N_14595,N_12934);
and U19778 (N_19778,N_12422,N_10584);
nor U19779 (N_19779,N_13387,N_12210);
xnor U19780 (N_19780,N_14853,N_14542);
xnor U19781 (N_19781,N_10478,N_12282);
nor U19782 (N_19782,N_12060,N_10211);
nor U19783 (N_19783,N_10119,N_10206);
xor U19784 (N_19784,N_10024,N_11917);
or U19785 (N_19785,N_14553,N_14914);
nand U19786 (N_19786,N_14993,N_11725);
xnor U19787 (N_19787,N_14972,N_11436);
or U19788 (N_19788,N_10728,N_11216);
nor U19789 (N_19789,N_12908,N_10482);
and U19790 (N_19790,N_12876,N_10824);
xnor U19791 (N_19791,N_10179,N_12763);
or U19792 (N_19792,N_11009,N_11368);
or U19793 (N_19793,N_12527,N_11451);
and U19794 (N_19794,N_14293,N_14621);
xnor U19795 (N_19795,N_13751,N_13793);
nor U19796 (N_19796,N_13257,N_13007);
and U19797 (N_19797,N_12235,N_14110);
nand U19798 (N_19798,N_14447,N_11137);
or U19799 (N_19799,N_11570,N_12821);
nand U19800 (N_19800,N_12000,N_10329);
and U19801 (N_19801,N_11123,N_14789);
nand U19802 (N_19802,N_11278,N_12410);
or U19803 (N_19803,N_12490,N_10782);
nor U19804 (N_19804,N_10700,N_13395);
or U19805 (N_19805,N_14762,N_14881);
xor U19806 (N_19806,N_11390,N_10288);
nor U19807 (N_19807,N_13694,N_10881);
nor U19808 (N_19808,N_11286,N_14711);
xor U19809 (N_19809,N_13088,N_10064);
nor U19810 (N_19810,N_14109,N_10379);
nand U19811 (N_19811,N_14301,N_13247);
nor U19812 (N_19812,N_12601,N_14823);
xnor U19813 (N_19813,N_13161,N_10121);
or U19814 (N_19814,N_11413,N_10285);
and U19815 (N_19815,N_14166,N_14189);
or U19816 (N_19816,N_10173,N_11599);
xor U19817 (N_19817,N_13947,N_11935);
and U19818 (N_19818,N_13797,N_10165);
nand U19819 (N_19819,N_11844,N_11914);
xnor U19820 (N_19820,N_14257,N_11373);
nand U19821 (N_19821,N_12961,N_12051);
xor U19822 (N_19822,N_14255,N_12678);
and U19823 (N_19823,N_11467,N_11004);
and U19824 (N_19824,N_10931,N_10446);
and U19825 (N_19825,N_11488,N_12977);
nor U19826 (N_19826,N_10356,N_11286);
nand U19827 (N_19827,N_10098,N_12140);
and U19828 (N_19828,N_13842,N_10535);
or U19829 (N_19829,N_10591,N_14412);
nor U19830 (N_19830,N_11020,N_14462);
nand U19831 (N_19831,N_10879,N_10070);
nor U19832 (N_19832,N_14302,N_10702);
nor U19833 (N_19833,N_12888,N_10170);
or U19834 (N_19834,N_10049,N_10188);
or U19835 (N_19835,N_11736,N_11540);
xor U19836 (N_19836,N_12329,N_10023);
and U19837 (N_19837,N_12851,N_12241);
xnor U19838 (N_19838,N_14954,N_14569);
xnor U19839 (N_19839,N_11050,N_10686);
xor U19840 (N_19840,N_13284,N_11385);
or U19841 (N_19841,N_11683,N_10747);
and U19842 (N_19842,N_14870,N_13230);
or U19843 (N_19843,N_11087,N_13549);
or U19844 (N_19844,N_12596,N_14469);
xor U19845 (N_19845,N_11565,N_10891);
or U19846 (N_19846,N_12441,N_11147);
xor U19847 (N_19847,N_10199,N_11764);
nor U19848 (N_19848,N_14689,N_11755);
or U19849 (N_19849,N_14199,N_12181);
nand U19850 (N_19850,N_13770,N_11807);
or U19851 (N_19851,N_14006,N_14978);
nand U19852 (N_19852,N_10487,N_11522);
or U19853 (N_19853,N_10928,N_12515);
nor U19854 (N_19854,N_12048,N_13076);
and U19855 (N_19855,N_14684,N_13477);
nand U19856 (N_19856,N_12036,N_11488);
nor U19857 (N_19857,N_14943,N_12135);
and U19858 (N_19858,N_14285,N_13351);
xor U19859 (N_19859,N_14975,N_11414);
nor U19860 (N_19860,N_11528,N_12988);
or U19861 (N_19861,N_10294,N_13253);
nor U19862 (N_19862,N_11751,N_10608);
or U19863 (N_19863,N_14077,N_10451);
nand U19864 (N_19864,N_10744,N_13401);
and U19865 (N_19865,N_13672,N_12306);
and U19866 (N_19866,N_12953,N_10635);
and U19867 (N_19867,N_13964,N_14010);
and U19868 (N_19868,N_13750,N_11770);
and U19869 (N_19869,N_14269,N_10580);
or U19870 (N_19870,N_10358,N_13908);
xnor U19871 (N_19871,N_13330,N_14228);
xnor U19872 (N_19872,N_10336,N_10959);
nor U19873 (N_19873,N_14055,N_11287);
nand U19874 (N_19874,N_10757,N_10136);
nand U19875 (N_19875,N_11004,N_11692);
xnor U19876 (N_19876,N_10754,N_11384);
and U19877 (N_19877,N_12296,N_13099);
or U19878 (N_19878,N_14818,N_10880);
xor U19879 (N_19879,N_10790,N_10133);
and U19880 (N_19880,N_13850,N_12157);
and U19881 (N_19881,N_14246,N_10793);
nor U19882 (N_19882,N_14358,N_14830);
nand U19883 (N_19883,N_10741,N_11660);
nand U19884 (N_19884,N_11524,N_12121);
nand U19885 (N_19885,N_12663,N_10611);
xnor U19886 (N_19886,N_14452,N_13541);
nor U19887 (N_19887,N_11429,N_10516);
nor U19888 (N_19888,N_12022,N_12071);
nor U19889 (N_19889,N_12213,N_11248);
and U19890 (N_19890,N_14006,N_13935);
nor U19891 (N_19891,N_14418,N_14971);
and U19892 (N_19892,N_12057,N_10497);
nor U19893 (N_19893,N_11914,N_12603);
and U19894 (N_19894,N_10672,N_14780);
or U19895 (N_19895,N_10978,N_11433);
and U19896 (N_19896,N_13143,N_13996);
nand U19897 (N_19897,N_11600,N_12998);
nand U19898 (N_19898,N_14378,N_14522);
xor U19899 (N_19899,N_12682,N_10838);
nor U19900 (N_19900,N_10223,N_10450);
nor U19901 (N_19901,N_11742,N_12820);
and U19902 (N_19902,N_12120,N_11678);
nand U19903 (N_19903,N_11335,N_12228);
nor U19904 (N_19904,N_13776,N_14752);
xnor U19905 (N_19905,N_11809,N_11242);
nor U19906 (N_19906,N_11773,N_13040);
and U19907 (N_19907,N_14819,N_10292);
and U19908 (N_19908,N_11686,N_12991);
xor U19909 (N_19909,N_14220,N_13431);
and U19910 (N_19910,N_12591,N_13599);
and U19911 (N_19911,N_10092,N_12258);
nand U19912 (N_19912,N_14487,N_10727);
and U19913 (N_19913,N_14876,N_13408);
or U19914 (N_19914,N_10995,N_12954);
xor U19915 (N_19915,N_10159,N_12033);
xnor U19916 (N_19916,N_14537,N_11995);
or U19917 (N_19917,N_11003,N_10625);
or U19918 (N_19918,N_13400,N_13322);
nor U19919 (N_19919,N_12548,N_10170);
nor U19920 (N_19920,N_12681,N_12455);
xor U19921 (N_19921,N_14853,N_11280);
xor U19922 (N_19922,N_10144,N_14231);
or U19923 (N_19923,N_14197,N_12238);
or U19924 (N_19924,N_14169,N_11493);
nand U19925 (N_19925,N_11334,N_11333);
nor U19926 (N_19926,N_13740,N_14421);
nand U19927 (N_19927,N_10295,N_11960);
xnor U19928 (N_19928,N_13023,N_12287);
or U19929 (N_19929,N_13790,N_14428);
nand U19930 (N_19930,N_11132,N_13056);
and U19931 (N_19931,N_11934,N_11061);
xor U19932 (N_19932,N_13897,N_13665);
nor U19933 (N_19933,N_11204,N_12331);
nand U19934 (N_19934,N_10705,N_14986);
and U19935 (N_19935,N_13510,N_10978);
nor U19936 (N_19936,N_13429,N_12116);
and U19937 (N_19937,N_11009,N_10519);
nand U19938 (N_19938,N_11387,N_11024);
or U19939 (N_19939,N_14854,N_10343);
nand U19940 (N_19940,N_12137,N_10100);
or U19941 (N_19941,N_11337,N_11934);
and U19942 (N_19942,N_12482,N_13413);
xor U19943 (N_19943,N_10748,N_14043);
or U19944 (N_19944,N_11872,N_12319);
or U19945 (N_19945,N_14547,N_10279);
xnor U19946 (N_19946,N_14749,N_10312);
or U19947 (N_19947,N_13596,N_11943);
or U19948 (N_19948,N_13908,N_14623);
xnor U19949 (N_19949,N_12932,N_12688);
xor U19950 (N_19950,N_10283,N_11806);
nand U19951 (N_19951,N_10778,N_11831);
nor U19952 (N_19952,N_14666,N_14392);
nand U19953 (N_19953,N_10187,N_11020);
nor U19954 (N_19954,N_11525,N_14068);
xor U19955 (N_19955,N_12725,N_10195);
and U19956 (N_19956,N_12450,N_10070);
or U19957 (N_19957,N_13581,N_12138);
nor U19958 (N_19958,N_13346,N_13506);
or U19959 (N_19959,N_12089,N_12157);
nor U19960 (N_19960,N_11926,N_13417);
and U19961 (N_19961,N_13231,N_12837);
nand U19962 (N_19962,N_11074,N_10593);
xnor U19963 (N_19963,N_12400,N_10817);
nand U19964 (N_19964,N_14792,N_13925);
and U19965 (N_19965,N_12940,N_10206);
or U19966 (N_19966,N_14007,N_11958);
or U19967 (N_19967,N_10357,N_13064);
xor U19968 (N_19968,N_10736,N_12171);
nor U19969 (N_19969,N_12866,N_11770);
or U19970 (N_19970,N_14871,N_14101);
nand U19971 (N_19971,N_12421,N_10623);
or U19972 (N_19972,N_13418,N_10131);
xor U19973 (N_19973,N_10296,N_12964);
nand U19974 (N_19974,N_10616,N_12716);
xor U19975 (N_19975,N_14249,N_14014);
or U19976 (N_19976,N_10280,N_13772);
and U19977 (N_19977,N_10945,N_14601);
nor U19978 (N_19978,N_14922,N_14639);
or U19979 (N_19979,N_13839,N_11483);
nor U19980 (N_19980,N_14678,N_11690);
xor U19981 (N_19981,N_13228,N_10683);
and U19982 (N_19982,N_11708,N_13708);
or U19983 (N_19983,N_10321,N_11606);
nor U19984 (N_19984,N_13534,N_13977);
or U19985 (N_19985,N_12691,N_10637);
or U19986 (N_19986,N_14827,N_10677);
and U19987 (N_19987,N_14204,N_12054);
or U19988 (N_19988,N_14452,N_12100);
nand U19989 (N_19989,N_11683,N_12361);
nand U19990 (N_19990,N_13748,N_14195);
xnor U19991 (N_19991,N_14715,N_14236);
or U19992 (N_19992,N_11586,N_13203);
nor U19993 (N_19993,N_12438,N_14712);
and U19994 (N_19994,N_10504,N_11468);
or U19995 (N_19995,N_10934,N_14189);
nor U19996 (N_19996,N_11044,N_11950);
xor U19997 (N_19997,N_13427,N_10813);
or U19998 (N_19998,N_12729,N_11799);
nor U19999 (N_19999,N_13251,N_14020);
or UO_0 (O_0,N_17860,N_18433);
nor UO_1 (O_1,N_16230,N_16595);
nor UO_2 (O_2,N_17622,N_18979);
xor UO_3 (O_3,N_18645,N_18815);
xor UO_4 (O_4,N_19914,N_19557);
and UO_5 (O_5,N_17301,N_15670);
and UO_6 (O_6,N_18475,N_15457);
or UO_7 (O_7,N_17970,N_19950);
xnor UO_8 (O_8,N_15872,N_15924);
and UO_9 (O_9,N_18393,N_17379);
and UO_10 (O_10,N_16178,N_17107);
nand UO_11 (O_11,N_16929,N_18081);
and UO_12 (O_12,N_15747,N_18176);
nor UO_13 (O_13,N_17114,N_15028);
nor UO_14 (O_14,N_17817,N_19697);
nor UO_15 (O_15,N_18830,N_17778);
and UO_16 (O_16,N_16234,N_19569);
or UO_17 (O_17,N_19738,N_15752);
xor UO_18 (O_18,N_18558,N_16353);
nor UO_19 (O_19,N_16747,N_19735);
nor UO_20 (O_20,N_15013,N_15915);
and UO_21 (O_21,N_18262,N_17461);
xor UO_22 (O_22,N_17734,N_18297);
nor UO_23 (O_23,N_17939,N_16279);
and UO_24 (O_24,N_19367,N_19902);
xnor UO_25 (O_25,N_16823,N_19217);
xnor UO_26 (O_26,N_18694,N_17774);
or UO_27 (O_27,N_16422,N_15651);
xnor UO_28 (O_28,N_18652,N_16618);
xor UO_29 (O_29,N_18070,N_17748);
and UO_30 (O_30,N_15765,N_19023);
nand UO_31 (O_31,N_16839,N_17450);
and UO_32 (O_32,N_19817,N_16419);
or UO_33 (O_33,N_19422,N_19712);
nand UO_34 (O_34,N_19140,N_19517);
xnor UO_35 (O_35,N_16143,N_15685);
nor UO_36 (O_36,N_18446,N_18035);
or UO_37 (O_37,N_15462,N_18267);
and UO_38 (O_38,N_17535,N_19453);
or UO_39 (O_39,N_19595,N_16381);
nor UO_40 (O_40,N_17957,N_19154);
nand UO_41 (O_41,N_19737,N_19324);
xor UO_42 (O_42,N_17271,N_18419);
and UO_43 (O_43,N_19520,N_15214);
and UO_44 (O_44,N_19560,N_18423);
nor UO_45 (O_45,N_16566,N_18106);
xor UO_46 (O_46,N_15690,N_15154);
and UO_47 (O_47,N_16849,N_18921);
xor UO_48 (O_48,N_17581,N_19810);
and UO_49 (O_49,N_17109,N_18405);
or UO_50 (O_50,N_15314,N_18024);
and UO_51 (O_51,N_15504,N_18834);
or UO_52 (O_52,N_16673,N_18950);
nor UO_53 (O_53,N_15005,N_16284);
nor UO_54 (O_54,N_17449,N_15088);
xnor UO_55 (O_55,N_15282,N_17967);
nor UO_56 (O_56,N_16003,N_19605);
nand UO_57 (O_57,N_18115,N_16660);
nand UO_58 (O_58,N_18014,N_16063);
nand UO_59 (O_59,N_18511,N_19183);
nand UO_60 (O_60,N_19402,N_16456);
nor UO_61 (O_61,N_16104,N_19187);
nand UO_62 (O_62,N_19503,N_19506);
nand UO_63 (O_63,N_15461,N_16399);
or UO_64 (O_64,N_19878,N_17527);
nor UO_65 (O_65,N_19652,N_15642);
and UO_66 (O_66,N_17524,N_18096);
nand UO_67 (O_67,N_19119,N_19285);
or UO_68 (O_68,N_17665,N_16168);
xor UO_69 (O_69,N_19479,N_17278);
and UO_70 (O_70,N_15992,N_16352);
nor UO_71 (O_71,N_19143,N_16240);
nand UO_72 (O_72,N_18227,N_17146);
xor UO_73 (O_73,N_18266,N_19661);
nand UO_74 (O_74,N_16067,N_15466);
or UO_75 (O_75,N_17982,N_18930);
xnor UO_76 (O_76,N_19028,N_17306);
or UO_77 (O_77,N_17833,N_17862);
nand UO_78 (O_78,N_18480,N_17378);
xnor UO_79 (O_79,N_19429,N_18365);
nand UO_80 (O_80,N_16702,N_17344);
nor UO_81 (O_81,N_15696,N_15615);
or UO_82 (O_82,N_19856,N_17809);
nand UO_83 (O_83,N_19237,N_15876);
and UO_84 (O_84,N_18723,N_18717);
and UO_85 (O_85,N_18064,N_15603);
xnor UO_86 (O_86,N_15261,N_18289);
nand UO_87 (O_87,N_15675,N_16206);
or UO_88 (O_88,N_15553,N_19978);
xor UO_89 (O_89,N_15026,N_17600);
nor UO_90 (O_90,N_15896,N_17380);
nand UO_91 (O_91,N_15280,N_18172);
xor UO_92 (O_92,N_18698,N_18478);
nor UO_93 (O_93,N_18051,N_17245);
and UO_94 (O_94,N_19206,N_17536);
xnor UO_95 (O_95,N_17233,N_17139);
or UO_96 (O_96,N_17744,N_16524);
xnor UO_97 (O_97,N_17779,N_16584);
or UO_98 (O_98,N_19260,N_16360);
nor UO_99 (O_99,N_19800,N_17101);
xnor UO_100 (O_100,N_19133,N_17965);
and UO_101 (O_101,N_17217,N_18610);
xnor UO_102 (O_102,N_18258,N_17545);
nand UO_103 (O_103,N_15938,N_15350);
nand UO_104 (O_104,N_19536,N_17376);
and UO_105 (O_105,N_15489,N_17607);
nand UO_106 (O_106,N_19087,N_19590);
or UO_107 (O_107,N_15239,N_19547);
xor UO_108 (O_108,N_16531,N_19778);
or UO_109 (O_109,N_19854,N_17171);
nor UO_110 (O_110,N_15993,N_17408);
nor UO_111 (O_111,N_15304,N_16836);
or UO_112 (O_112,N_19869,N_17123);
nand UO_113 (O_113,N_18640,N_18908);
xnor UO_114 (O_114,N_18592,N_18263);
xor UO_115 (O_115,N_19678,N_18667);
nor UO_116 (O_116,N_15066,N_17364);
xnor UO_117 (O_117,N_15930,N_16626);
nand UO_118 (O_118,N_18758,N_15391);
xor UO_119 (O_119,N_19879,N_15961);
or UO_120 (O_120,N_16526,N_16184);
nor UO_121 (O_121,N_17058,N_16869);
nand UO_122 (O_122,N_19955,N_17574);
nand UO_123 (O_123,N_15016,N_18788);
xor UO_124 (O_124,N_19431,N_17293);
xnor UO_125 (O_125,N_15439,N_16989);
nor UO_126 (O_126,N_17385,N_18056);
nor UO_127 (O_127,N_18838,N_17304);
and UO_128 (O_128,N_19939,N_17717);
or UO_129 (O_129,N_16964,N_17668);
nor UO_130 (O_130,N_17025,N_17081);
xnor UO_131 (O_131,N_18370,N_18944);
and UO_132 (O_132,N_15926,N_15021);
and UO_133 (O_133,N_15476,N_16275);
xnor UO_134 (O_134,N_19215,N_16932);
and UO_135 (O_135,N_19870,N_18119);
nand UO_136 (O_136,N_19516,N_17090);
and UO_137 (O_137,N_18006,N_19256);
or UO_138 (O_138,N_18941,N_17371);
nand UO_139 (O_139,N_15023,N_16333);
xor UO_140 (O_140,N_19226,N_19178);
or UO_141 (O_141,N_17009,N_19663);
or UO_142 (O_142,N_15233,N_18767);
nand UO_143 (O_143,N_16805,N_18681);
or UO_144 (O_144,N_16078,N_17940);
and UO_145 (O_145,N_17707,N_17129);
nor UO_146 (O_146,N_15890,N_19495);
nand UO_147 (O_147,N_17182,N_15098);
nor UO_148 (O_148,N_17203,N_17749);
or UO_149 (O_149,N_17764,N_15894);
nand UO_150 (O_150,N_18940,N_16040);
nor UO_151 (O_151,N_18749,N_15602);
nor UO_152 (O_152,N_18848,N_19081);
nor UO_153 (O_153,N_19907,N_19499);
nand UO_154 (O_154,N_15585,N_17667);
nand UO_155 (O_155,N_15137,N_18460);
nor UO_156 (O_156,N_19204,N_17054);
xor UO_157 (O_157,N_15315,N_17465);
or UO_158 (O_158,N_16358,N_17452);
nor UO_159 (O_159,N_19910,N_19155);
nor UO_160 (O_160,N_17026,N_17598);
xor UO_161 (O_161,N_17260,N_17288);
nand UO_162 (O_162,N_16301,N_19413);
or UO_163 (O_163,N_15119,N_16935);
or UO_164 (O_164,N_15164,N_15040);
nand UO_165 (O_165,N_18129,N_15617);
nand UO_166 (O_166,N_15086,N_17196);
xor UO_167 (O_167,N_17137,N_17281);
or UO_168 (O_168,N_19476,N_15837);
nand UO_169 (O_169,N_17213,N_19197);
xnor UO_170 (O_170,N_16493,N_16972);
or UO_171 (O_171,N_17396,N_16314);
nand UO_172 (O_172,N_16560,N_18503);
nor UO_173 (O_173,N_17354,N_16926);
nand UO_174 (O_174,N_15133,N_19241);
xnor UO_175 (O_175,N_18962,N_17525);
or UO_176 (O_176,N_15730,N_17892);
nor UO_177 (O_177,N_18973,N_15296);
or UO_178 (O_178,N_17893,N_16995);
and UO_179 (O_179,N_15318,N_16950);
or UO_180 (O_180,N_18657,N_19244);
xor UO_181 (O_181,N_16198,N_18541);
or UO_182 (O_182,N_16476,N_19015);
and UO_183 (O_183,N_18823,N_18642);
or UO_184 (O_184,N_15432,N_16377);
and UO_185 (O_185,N_19968,N_18217);
nand UO_186 (O_186,N_16973,N_16440);
nand UO_187 (O_187,N_17074,N_15900);
or UO_188 (O_188,N_16763,N_15147);
and UO_189 (O_189,N_17195,N_17653);
xnor UO_190 (O_190,N_16996,N_15948);
nor UO_191 (O_191,N_17199,N_19103);
nand UO_192 (O_192,N_16686,N_15606);
or UO_193 (O_193,N_17898,N_18508);
nor UO_194 (O_194,N_17246,N_15204);
nor UO_195 (O_195,N_19224,N_16281);
nor UO_196 (O_196,N_18875,N_17888);
or UO_197 (O_197,N_18027,N_18138);
xor UO_198 (O_198,N_19608,N_18658);
nor UO_199 (O_199,N_17554,N_19981);
nor UO_200 (O_200,N_15799,N_15820);
xor UO_201 (O_201,N_19451,N_18917);
nand UO_202 (O_202,N_15437,N_16154);
or UO_203 (O_203,N_17285,N_18529);
and UO_204 (O_204,N_15500,N_15917);
nand UO_205 (O_205,N_15259,N_16817);
or UO_206 (O_206,N_15763,N_19489);
or UO_207 (O_207,N_19296,N_18968);
nor UO_208 (O_208,N_17874,N_15366);
xnor UO_209 (O_209,N_16006,N_18726);
xor UO_210 (O_210,N_17126,N_16776);
xnor UO_211 (O_211,N_15008,N_17896);
nand UO_212 (O_212,N_18918,N_16244);
or UO_213 (O_213,N_17855,N_17181);
and UO_214 (O_214,N_17803,N_15779);
and UO_215 (O_215,N_17954,N_15145);
or UO_216 (O_216,N_18421,N_19942);
nor UO_217 (O_217,N_18967,N_17176);
nand UO_218 (O_218,N_16803,N_17695);
nor UO_219 (O_219,N_15785,N_16986);
or UO_220 (O_220,N_19567,N_17721);
nor UO_221 (O_221,N_17520,N_17144);
and UO_222 (O_222,N_18149,N_19196);
xor UO_223 (O_223,N_19483,N_18826);
nor UO_224 (O_224,N_16915,N_18379);
or UO_225 (O_225,N_17027,N_15046);
nor UO_226 (O_226,N_15446,N_17840);
and UO_227 (O_227,N_15482,N_19934);
or UO_228 (O_228,N_19032,N_19524);
nand UO_229 (O_229,N_19995,N_19316);
nor UO_230 (O_230,N_16411,N_19356);
xor UO_231 (O_231,N_16273,N_19535);
nand UO_232 (O_232,N_15390,N_15174);
nand UO_233 (O_233,N_15134,N_17522);
and UO_234 (O_234,N_18567,N_18257);
or UO_235 (O_235,N_18672,N_19598);
xor UO_236 (O_236,N_15297,N_15006);
nor UO_237 (O_237,N_15004,N_16228);
and UO_238 (O_238,N_19374,N_16743);
xnor UO_239 (O_239,N_17773,N_19670);
or UO_240 (O_240,N_18811,N_19044);
or UO_241 (O_241,N_15289,N_19504);
nor UO_242 (O_242,N_19419,N_17122);
nand UO_243 (O_243,N_18026,N_15762);
nor UO_244 (O_244,N_18005,N_19207);
and UO_245 (O_245,N_17656,N_16080);
and UO_246 (O_246,N_18911,N_19986);
and UO_247 (O_247,N_19975,N_17343);
xor UO_248 (O_248,N_18191,N_15228);
or UO_249 (O_249,N_18268,N_18605);
nand UO_250 (O_250,N_15731,N_17041);
nor UO_251 (O_251,N_17990,N_19623);
nor UO_252 (O_252,N_17185,N_16896);
nor UO_253 (O_253,N_16372,N_17983);
nor UO_254 (O_254,N_15727,N_17366);
and UO_255 (O_255,N_19548,N_18884);
nand UO_256 (O_256,N_18265,N_17457);
and UO_257 (O_257,N_17407,N_16406);
xnor UO_258 (O_258,N_19077,N_15749);
or UO_259 (O_259,N_19365,N_19390);
or UO_260 (O_260,N_16748,N_17722);
nor UO_261 (O_261,N_18317,N_17799);
nor UO_262 (O_262,N_16313,N_15887);
or UO_263 (O_263,N_18234,N_19864);
or UO_264 (O_264,N_15030,N_16039);
and UO_265 (O_265,N_18739,N_19128);
nand UO_266 (O_266,N_16548,N_19011);
or UO_267 (O_267,N_17445,N_17120);
and UO_268 (O_268,N_15469,N_15808);
nand UO_269 (O_269,N_19046,N_18641);
or UO_270 (O_270,N_19667,N_17859);
nor UO_271 (O_271,N_15575,N_18988);
nor UO_272 (O_272,N_16151,N_17095);
xnor UO_273 (O_273,N_18107,N_18057);
xnor UO_274 (O_274,N_16933,N_19675);
xnor UO_275 (O_275,N_19501,N_15502);
nor UO_276 (O_276,N_16768,N_19076);
nand UO_277 (O_277,N_18915,N_19362);
nand UO_278 (O_278,N_18184,N_15031);
nand UO_279 (O_279,N_15569,N_17214);
nor UO_280 (O_280,N_15377,N_18678);
nand UO_281 (O_281,N_18703,N_16255);
nor UO_282 (O_282,N_17089,N_19475);
and UO_283 (O_283,N_19126,N_18286);
or UO_284 (O_284,N_18556,N_19732);
nor UO_285 (O_285,N_18814,N_18891);
or UO_286 (O_286,N_17111,N_18000);
and UO_287 (O_287,N_18562,N_16064);
nand UO_288 (O_288,N_18103,N_17516);
nand UO_289 (O_289,N_16231,N_17775);
nand UO_290 (O_290,N_17549,N_17350);
or UO_291 (O_291,N_18909,N_17875);
or UO_292 (O_292,N_18235,N_15657);
and UO_293 (O_293,N_16388,N_18974);
and UO_294 (O_294,N_16642,N_15153);
nand UO_295 (O_295,N_17415,N_15689);
xnor UO_296 (O_296,N_19245,N_15686);
nand UO_297 (O_297,N_18148,N_18361);
and UO_298 (O_298,N_18679,N_17531);
and UO_299 (O_299,N_16141,N_15015);
and UO_300 (O_300,N_16646,N_16183);
nor UO_301 (O_301,N_16450,N_18137);
or UO_302 (O_302,N_18894,N_15798);
and UO_303 (O_303,N_18292,N_18253);
nor UO_304 (O_304,N_19194,N_19181);
or UO_305 (O_305,N_15532,N_18886);
nor UO_306 (O_306,N_18426,N_19287);
xor UO_307 (O_307,N_16523,N_18187);
or UO_308 (O_308,N_17927,N_19725);
xnor UO_309 (O_309,N_15002,N_19442);
xnor UO_310 (O_310,N_19223,N_16857);
nand UO_311 (O_311,N_16386,N_15591);
xor UO_312 (O_312,N_16821,N_17492);
or UO_313 (O_313,N_18994,N_16838);
xor UO_314 (O_314,N_19049,N_18887);
nand UO_315 (O_315,N_16786,N_16305);
or UO_316 (O_316,N_16378,N_17234);
and UO_317 (O_317,N_18568,N_19600);
xor UO_318 (O_318,N_19612,N_17412);
nand UO_319 (O_319,N_18799,N_19284);
and UO_320 (O_320,N_15202,N_15175);
xor UO_321 (O_321,N_19289,N_16813);
xor UO_322 (O_322,N_15370,N_16976);
xnor UO_323 (O_323,N_15494,N_15627);
and UO_324 (O_324,N_18618,N_18113);
xnor UO_325 (O_325,N_15076,N_16431);
xor UO_326 (O_326,N_19384,N_16402);
and UO_327 (O_327,N_17780,N_16518);
and UO_328 (O_328,N_19082,N_16041);
nand UO_329 (O_329,N_16343,N_19294);
nand UO_330 (O_330,N_15378,N_19893);
and UO_331 (O_331,N_17963,N_15358);
nand UO_332 (O_332,N_18464,N_18506);
and UO_333 (O_333,N_17034,N_15913);
and UO_334 (O_334,N_15570,N_16514);
xor UO_335 (O_335,N_19871,N_16021);
nand UO_336 (O_336,N_16497,N_15144);
or UO_337 (O_337,N_19331,N_16201);
nand UO_338 (O_338,N_19065,N_17071);
and UO_339 (O_339,N_18879,N_19167);
or UO_340 (O_340,N_15839,N_17998);
or UO_341 (O_341,N_16014,N_19010);
nor UO_342 (O_342,N_16057,N_18841);
xnor UO_343 (O_343,N_17459,N_15135);
nor UO_344 (O_344,N_18590,N_15760);
or UO_345 (O_345,N_16429,N_18920);
nor UO_346 (O_346,N_19382,N_16445);
or UO_347 (O_347,N_15552,N_19736);
nor UO_348 (O_348,N_19649,N_15042);
xnor UO_349 (O_349,N_17348,N_19397);
and UO_350 (O_350,N_18321,N_16068);
nand UO_351 (O_351,N_18049,N_19683);
xnor UO_352 (O_352,N_15975,N_15250);
nor UO_353 (O_353,N_16772,N_15235);
nor UO_354 (O_354,N_19676,N_19043);
nor UO_355 (O_355,N_15867,N_15351);
or UO_356 (O_356,N_16349,N_18538);
nor UO_357 (O_357,N_19347,N_15847);
nand UO_358 (O_358,N_19936,N_17154);
and UO_359 (O_359,N_16017,N_15320);
and UO_360 (O_360,N_17877,N_16004);
and UO_361 (O_361,N_19890,N_15758);
nand UO_362 (O_362,N_19466,N_15372);
nand UO_363 (O_363,N_16008,N_15712);
xor UO_364 (O_364,N_17367,N_15538);
nand UO_365 (O_365,N_15737,N_18314);
nand UO_366 (O_366,N_16187,N_18414);
or UO_367 (O_367,N_19733,N_15085);
and UO_368 (O_368,N_18260,N_15513);
or UO_369 (O_369,N_16199,N_16729);
nand UO_370 (O_370,N_19789,N_15554);
xor UO_371 (O_371,N_17497,N_18507);
and UO_372 (O_372,N_15354,N_16226);
nand UO_373 (O_373,N_19363,N_15518);
nand UO_374 (O_374,N_19407,N_15984);
xnor UO_375 (O_375,N_17273,N_19430);
nand UO_376 (O_376,N_16542,N_15947);
and UO_377 (O_377,N_19545,N_18801);
nand UO_378 (O_378,N_15664,N_16106);
nor UO_379 (O_379,N_15982,N_15179);
xnor UO_380 (O_380,N_19468,N_18435);
xor UO_381 (O_381,N_17130,N_15925);
or UO_382 (O_382,N_16046,N_18980);
and UO_383 (O_383,N_19759,N_17724);
or UO_384 (O_384,N_18987,N_18223);
nor UO_385 (O_385,N_18502,N_18704);
xnor UO_386 (O_386,N_15804,N_18048);
xor UO_387 (O_387,N_15769,N_18589);
and UO_388 (O_388,N_17991,N_18494);
nor UO_389 (O_389,N_18984,N_19826);
nand UO_390 (O_390,N_17552,N_18416);
nand UO_391 (O_391,N_16794,N_15526);
or UO_392 (O_392,N_15613,N_16454);
and UO_393 (O_393,N_16549,N_16264);
xor UO_394 (O_394,N_19309,N_17719);
nor UO_395 (O_395,N_19443,N_19912);
xor UO_396 (O_396,N_17346,N_18545);
nand UO_397 (O_397,N_17868,N_18722);
and UO_398 (O_398,N_19299,N_18334);
and UO_399 (O_399,N_16999,N_16738);
xnor UO_400 (O_400,N_15454,N_19270);
nor UO_401 (O_401,N_19057,N_17012);
or UO_402 (O_402,N_17710,N_18169);
nor UO_403 (O_403,N_16227,N_17190);
nand UO_404 (O_404,N_17197,N_19319);
xnor UO_405 (O_405,N_15208,N_19069);
nand UO_406 (O_406,N_16623,N_16121);
or UO_407 (O_407,N_18104,N_18923);
nor UO_408 (O_408,N_15285,N_19346);
or UO_409 (O_409,N_16847,N_19297);
or UO_410 (O_410,N_15220,N_18151);
nor UO_411 (O_411,N_19777,N_17479);
xor UO_412 (O_412,N_16452,N_18874);
or UO_413 (O_413,N_19563,N_16829);
xor UO_414 (O_414,N_15155,N_16118);
xor UO_415 (O_415,N_19177,N_19905);
nor UO_416 (O_416,N_18491,N_15247);
nor UO_417 (O_417,N_18636,N_15962);
nand UO_418 (O_418,N_15053,N_18033);
xor UO_419 (O_419,N_16961,N_17061);
or UO_420 (O_420,N_19399,N_18910);
and UO_421 (O_421,N_15449,N_19099);
and UO_422 (O_422,N_18624,N_16174);
nand UO_423 (O_423,N_18152,N_15932);
or UO_424 (O_424,N_17956,N_16749);
or UO_425 (O_425,N_19385,N_18183);
or UO_426 (O_426,N_17615,N_17272);
or UO_427 (O_427,N_15877,N_15367);
nor UO_428 (O_428,N_16047,N_16661);
and UO_429 (O_429,N_15997,N_15114);
or UO_430 (O_430,N_15519,N_17252);
nor UO_431 (O_431,N_18328,N_19259);
nand UO_432 (O_432,N_16718,N_17905);
xnor UO_433 (O_433,N_16942,N_18588);
or UO_434 (O_434,N_19710,N_15802);
and UO_435 (O_435,N_17669,N_17951);
and UO_436 (O_436,N_17894,N_19549);
nor UO_437 (O_437,N_19423,N_15191);
or UO_438 (O_438,N_18531,N_19677);
xor UO_439 (O_439,N_19131,N_15495);
nand UO_440 (O_440,N_18036,N_19231);
and UO_441 (O_441,N_16886,N_18481);
nand UO_442 (O_442,N_16656,N_16001);
xor UO_443 (O_443,N_15786,N_18298);
xnor UO_444 (O_444,N_18876,N_16577);
and UO_445 (O_445,N_15599,N_17436);
xor UO_446 (O_446,N_19266,N_19768);
and UO_447 (O_447,N_15678,N_18214);
and UO_448 (O_448,N_19631,N_18959);
nor UO_449 (O_449,N_18252,N_18937);
or UO_450 (O_450,N_15311,N_16808);
nand UO_451 (O_451,N_15420,N_16195);
nor UO_452 (O_452,N_18742,N_19498);
or UO_453 (O_453,N_18824,N_19774);
nor UO_454 (O_454,N_16681,N_15382);
or UO_455 (O_455,N_15534,N_19491);
nand UO_456 (O_456,N_15922,N_16905);
xnor UO_457 (O_457,N_15362,N_17046);
nor UO_458 (O_458,N_17121,N_16400);
nand UO_459 (O_459,N_15195,N_15022);
or UO_460 (O_460,N_18582,N_19348);
and UO_461 (O_461,N_16024,N_19092);
xnor UO_462 (O_462,N_18631,N_18261);
nor UO_463 (O_463,N_18804,N_19690);
or UO_464 (O_464,N_18397,N_19421);
nor UO_465 (O_465,N_19964,N_18425);
nor UO_466 (O_466,N_15100,N_19416);
nor UO_467 (O_467,N_17663,N_17422);
xnor UO_468 (O_468,N_19997,N_19274);
or UO_469 (O_469,N_19926,N_16674);
or UO_470 (O_470,N_17259,N_19551);
nand UO_471 (O_471,N_19992,N_19750);
nor UO_472 (O_472,N_16393,N_18181);
nor UO_473 (O_473,N_18904,N_16752);
nor UO_474 (O_474,N_18727,N_16750);
nand UO_475 (O_475,N_18845,N_19037);
or UO_476 (O_476,N_16156,N_18073);
and UO_477 (O_477,N_17478,N_16512);
xor UO_478 (O_478,N_19460,N_17289);
xnor UO_479 (O_479,N_15971,N_18175);
and UO_480 (O_480,N_18294,N_19261);
xnor UO_481 (O_481,N_18109,N_16269);
and UO_482 (O_482,N_17317,N_17808);
and UO_483 (O_483,N_17079,N_18851);
or UO_484 (O_484,N_15931,N_18131);
nand UO_485 (O_485,N_15159,N_16731);
nor UO_486 (O_486,N_16798,N_15866);
nand UO_487 (O_487,N_19574,N_15481);
xnor UO_488 (O_488,N_17928,N_18381);
or UO_489 (O_489,N_16510,N_19314);
nor UO_490 (O_490,N_19444,N_15187);
or UO_491 (O_491,N_18714,N_18774);
or UO_492 (O_492,N_16220,N_19005);
and UO_493 (O_493,N_19762,N_17362);
xor UO_494 (O_494,N_15265,N_18522);
nor UO_495 (O_495,N_15484,N_19664);
nand UO_496 (O_496,N_16654,N_15733);
xnor UO_497 (O_497,N_15636,N_15793);
or UO_498 (O_498,N_17091,N_17431);
xor UO_499 (O_499,N_18695,N_17563);
xnor UO_500 (O_500,N_16394,N_18548);
or UO_501 (O_501,N_18170,N_16815);
nand UO_502 (O_502,N_18740,N_16814);
and UO_503 (O_503,N_19016,N_17319);
or UO_504 (O_504,N_19695,N_18593);
xnor UO_505 (O_505,N_18795,N_16755);
or UO_506 (O_506,N_16648,N_18601);
nor UO_507 (O_507,N_16906,N_18552);
nor UO_508 (O_508,N_18971,N_16318);
nand UO_509 (O_509,N_17321,N_16608);
xor UO_510 (O_510,N_16538,N_16913);
or UO_511 (O_511,N_18118,N_16086);
nor UO_512 (O_512,N_16028,N_17692);
nor UO_513 (O_513,N_15121,N_15400);
or UO_514 (O_514,N_18960,N_18518);
nor UO_515 (O_515,N_15907,N_19593);
nor UO_516 (O_516,N_16267,N_19317);
xnor UO_517 (O_517,N_16107,N_16820);
nand UO_518 (O_518,N_19280,N_18357);
nor UO_519 (O_519,N_15665,N_17086);
or UO_520 (O_520,N_15507,N_15262);
and UO_521 (O_521,N_15716,N_18822);
nor UO_522 (O_522,N_16979,N_16076);
or UO_523 (O_523,N_15267,N_18474);
and UO_524 (O_524,N_18747,N_18270);
nor UO_525 (O_525,N_15976,N_17846);
xnor UO_526 (O_526,N_18347,N_15918);
or UO_527 (O_527,N_19078,N_16423);
nor UO_528 (O_528,N_18333,N_16248);
or UO_529 (O_529,N_15317,N_19139);
nand UO_530 (O_530,N_19618,N_16945);
or UO_531 (O_531,N_19149,N_18243);
nor UO_532 (O_532,N_17687,N_16978);
nor UO_533 (O_533,N_19185,N_17383);
and UO_534 (O_534,N_19748,N_16398);
or UO_535 (O_535,N_18530,N_18825);
nor UO_536 (O_536,N_19841,N_19828);
nor UO_537 (O_537,N_17472,N_16022);
or UO_538 (O_538,N_18244,N_16477);
or UO_539 (O_539,N_15058,N_18970);
nand UO_540 (O_540,N_17451,N_15697);
xnor UO_541 (O_541,N_17205,N_19671);
and UO_542 (O_542,N_16435,N_16294);
nand UO_543 (O_543,N_15954,N_15899);
or UO_544 (O_544,N_17603,N_17406);
xor UO_545 (O_545,N_15215,N_18721);
and UO_546 (O_546,N_18769,N_18866);
xor UO_547 (O_547,N_17539,N_17537);
and UO_548 (O_548,N_15775,N_18630);
or UO_549 (O_549,N_16527,N_16534);
xor UO_550 (O_550,N_16736,N_15392);
or UO_551 (O_551,N_19801,N_15969);
nor UO_552 (O_552,N_19214,N_19354);
nor UO_553 (O_553,N_19723,N_15142);
xnor UO_554 (O_554,N_16324,N_19436);
xnor UO_555 (O_555,N_15269,N_16016);
and UO_556 (O_556,N_17232,N_17930);
nor UO_557 (O_557,N_15433,N_18543);
nand UO_558 (O_558,N_15107,N_18933);
or UO_559 (O_559,N_19478,N_17094);
xnor UO_560 (O_560,N_16136,N_19990);
nand UO_561 (O_561,N_18623,N_18756);
or UO_562 (O_562,N_18364,N_15474);
and UO_563 (O_563,N_18061,N_15387);
xnor UO_564 (O_564,N_17946,N_17819);
and UO_565 (O_565,N_16918,N_15498);
and UO_566 (O_566,N_19221,N_15791);
and UO_567 (O_567,N_15855,N_16270);
nand UO_568 (O_568,N_15699,N_19655);
and UO_569 (O_569,N_15090,N_18403);
and UO_570 (O_570,N_18046,N_15240);
xnor UO_571 (O_571,N_19812,N_16874);
nand UO_572 (O_572,N_17861,N_15882);
nand UO_573 (O_573,N_18813,N_16011);
xnor UO_574 (O_574,N_19722,N_15829);
nand UO_575 (O_575,N_17747,N_18476);
nor UO_576 (O_576,N_15169,N_15755);
and UO_577 (O_577,N_19279,N_15693);
nand UO_578 (O_578,N_18755,N_15337);
nor UO_579 (O_579,N_15356,N_17363);
or UO_580 (O_580,N_15124,N_15794);
and UO_581 (O_581,N_16730,N_17767);
xor UO_582 (O_582,N_15863,N_16590);
or UO_583 (O_583,N_16927,N_18493);
xnor UO_584 (O_584,N_19747,N_17766);
and UO_585 (O_585,N_18088,N_18706);
and UO_586 (O_586,N_17736,N_16142);
xnor UO_587 (O_587,N_19298,N_16052);
nand UO_588 (O_588,N_18094,N_17761);
xnor UO_589 (O_589,N_16437,N_16977);
nor UO_590 (O_590,N_19919,N_15522);
and UO_591 (O_591,N_16898,N_19659);
and UO_592 (O_592,N_19823,N_17386);
nand UO_593 (O_593,N_17230,N_16810);
and UO_594 (O_594,N_15966,N_18074);
xnor UO_595 (O_595,N_17326,N_15879);
or UO_596 (O_596,N_19195,N_19071);
nand UO_597 (O_597,N_19959,N_17322);
or UO_598 (O_598,N_16715,N_18132);
or UO_599 (O_599,N_15115,N_19829);
and UO_600 (O_600,N_17482,N_18546);
nor UO_601 (O_601,N_19328,N_19689);
xnor UO_602 (O_602,N_18514,N_16427);
nand UO_603 (O_603,N_16460,N_17238);
nand UO_604 (O_604,N_16347,N_16578);
xnor UO_605 (O_605,N_18455,N_16628);
or UO_606 (O_606,N_17879,N_16638);
or UO_607 (O_607,N_19275,N_19171);
nor UO_608 (O_608,N_19606,N_18587);
xor UO_609 (O_609,N_16340,N_18828);
and UO_610 (O_610,N_19749,N_16179);
xnor UO_611 (O_611,N_16096,N_15949);
nand UO_612 (O_612,N_15610,N_19783);
nand UO_613 (O_613,N_16941,N_18544);
nand UO_614 (O_614,N_15645,N_18185);
nand UO_615 (O_615,N_17941,N_17659);
xor UO_616 (O_616,N_16556,N_15380);
or UO_617 (O_617,N_15736,N_17709);
and UO_618 (O_618,N_15549,N_15229);
xnor UO_619 (O_619,N_15422,N_15643);
and UO_620 (O_620,N_16059,N_16591);
and UO_621 (O_621,N_19465,N_18043);
or UO_622 (O_622,N_16037,N_15757);
and UO_623 (O_623,N_17599,N_16533);
or UO_624 (O_624,N_19692,N_17295);
and UO_625 (O_625,N_19007,N_19201);
xnor UO_626 (O_626,N_19130,N_17100);
nand UO_627 (O_627,N_18312,N_15713);
and UO_628 (O_628,N_17037,N_16951);
nor UO_629 (O_629,N_16509,N_16921);
nor UO_630 (O_630,N_15505,N_16925);
nand UO_631 (O_631,N_17538,N_18765);
or UO_632 (O_632,N_18928,N_15940);
and UO_633 (O_633,N_15376,N_17872);
xnor UO_634 (O_634,N_19116,N_17138);
and UO_635 (O_635,N_15274,N_19349);
nand UO_636 (O_636,N_18520,N_17099);
nand UO_637 (O_637,N_15342,N_19072);
xor UO_638 (O_638,N_17670,N_19360);
or UO_639 (O_639,N_19534,N_19622);
or UO_640 (O_640,N_16116,N_16344);
nor UO_641 (O_641,N_16647,N_15990);
or UO_642 (O_642,N_18408,N_17514);
xnor UO_643 (O_643,N_15272,N_18130);
and UO_644 (O_644,N_16883,N_15117);
or UO_645 (O_645,N_17610,N_16229);
nor UO_646 (O_646,N_16545,N_16844);
xnor UO_647 (O_647,N_18540,N_16291);
nand UO_648 (O_648,N_16616,N_19301);
or UO_649 (O_649,N_17430,N_19079);
nand UO_650 (O_650,N_17688,N_17003);
xor UO_651 (O_651,N_18855,N_18114);
and UO_652 (O_652,N_16089,N_17324);
or UO_653 (O_653,N_17679,N_18369);
nand UO_654 (O_654,N_18178,N_19586);
xor UO_655 (O_655,N_19510,N_19165);
xor UO_656 (O_656,N_16271,N_15740);
xor UO_657 (O_657,N_16696,N_17648);
nor UO_658 (O_658,N_19896,N_16887);
nand UO_659 (O_659,N_17337,N_18071);
and UO_660 (O_660,N_17978,N_15258);
nand UO_661 (O_661,N_17562,N_19490);
nor UO_662 (O_662,N_19881,N_19448);
nand UO_663 (O_663,N_19379,N_18355);
and UO_664 (O_664,N_16543,N_16818);
or UO_665 (O_665,N_18086,N_18764);
or UO_666 (O_666,N_19310,N_18078);
nor UO_667 (O_667,N_17727,N_18961);
xor UO_668 (O_668,N_17592,N_15901);
xor UO_669 (O_669,N_17758,N_15054);
or UO_670 (O_670,N_17216,N_17116);
xnor UO_671 (O_671,N_15097,N_19656);
and UO_672 (O_672,N_15225,N_18275);
or UO_673 (O_673,N_17828,N_15560);
nand UO_674 (O_674,N_19064,N_15338);
xnor UO_675 (O_675,N_19286,N_16165);
nand UO_676 (O_676,N_17308,N_15849);
xor UO_677 (O_677,N_17513,N_18793);
nand UO_678 (O_678,N_17740,N_16936);
nor UO_679 (O_679,N_18391,N_19323);
xor UO_680 (O_680,N_17175,N_17517);
or UO_681 (O_681,N_19632,N_17698);
and UO_682 (O_682,N_17134,N_19956);
nor UO_683 (O_683,N_15952,N_18300);
and UO_684 (O_684,N_19615,N_17274);
xnor UO_685 (O_685,N_17305,N_16265);
or UO_686 (O_686,N_16023,N_18445);
nand UO_687 (O_687,N_15414,N_18389);
nor UO_688 (O_688,N_19066,N_16410);
xor UO_689 (O_689,N_19089,N_15047);
nor UO_690 (O_690,N_17439,N_15355);
nand UO_691 (O_691,N_16380,N_15029);
or UO_692 (O_692,N_18313,N_17624);
nand UO_693 (O_693,N_17136,N_18687);
nand UO_694 (O_694,N_17638,N_15806);
nand UO_695 (O_695,N_18413,N_17481);
and UO_696 (O_696,N_18065,N_16561);
xnor UO_697 (O_697,N_19420,N_16633);
nand UO_698 (O_698,N_18797,N_16446);
nand UO_699 (O_699,N_19537,N_18311);
and UO_700 (O_700,N_16732,N_17635);
and UO_701 (O_701,N_18604,N_16311);
or UO_702 (O_702,N_19393,N_19727);
or UO_703 (O_703,N_17448,N_16965);
and UO_704 (O_704,N_18609,N_17469);
or UO_705 (O_705,N_18232,N_16899);
and UO_706 (O_706,N_17835,N_19439);
xnor UO_707 (O_707,N_16778,N_18100);
and UO_708 (O_708,N_17634,N_16722);
and UO_709 (O_709,N_18105,N_17823);
nor UO_710 (O_710,N_18054,N_19575);
nor UO_711 (O_711,N_18422,N_17542);
xor UO_712 (O_712,N_19858,N_16487);
nand UO_713 (O_713,N_19054,N_17249);
or UO_714 (O_714,N_15111,N_17885);
and UO_715 (O_715,N_18483,N_19114);
and UO_716 (O_716,N_19930,N_18194);
nor UO_717 (O_717,N_19027,N_17639);
xnor UO_718 (O_718,N_15227,N_19486);
nand UO_719 (O_719,N_17193,N_15373);
nor UO_720 (O_720,N_15172,N_16484);
nor UO_721 (O_721,N_16797,N_18513);
xnor UO_722 (O_722,N_17508,N_18812);
nand UO_723 (O_723,N_16541,N_17277);
or UO_724 (O_724,N_15150,N_15050);
xnor UO_725 (O_725,N_16330,N_17063);
nor UO_726 (O_726,N_19400,N_15632);
and UO_727 (O_727,N_17680,N_18537);
xnor UO_728 (O_728,N_17887,N_19220);
xnor UO_729 (O_729,N_15951,N_18869);
nor UO_730 (O_730,N_15881,N_18807);
and UO_731 (O_731,N_15634,N_16773);
nor UO_732 (O_732,N_15974,N_15795);
and UO_733 (O_733,N_17938,N_18741);
and UO_734 (O_734,N_18750,N_18066);
xnor UO_735 (O_735,N_15864,N_19614);
or UO_736 (O_736,N_17160,N_16300);
and UO_737 (O_737,N_16366,N_16053);
or UO_738 (O_738,N_16990,N_17287);
and UO_739 (O_739,N_17526,N_18158);
xor UO_740 (O_740,N_15118,N_17880);
nor UO_741 (O_741,N_16771,N_18343);
or UO_742 (O_742,N_15941,N_18432);
nor UO_743 (O_743,N_17529,N_18492);
nor UO_744 (O_744,N_16412,N_16546);
and UO_745 (O_745,N_16756,N_15994);
xor UO_746 (O_746,N_15910,N_19189);
nand UO_747 (O_747,N_16678,N_17674);
or UO_748 (O_748,N_18569,N_16554);
nor UO_749 (O_749,N_16205,N_16137);
nor UO_750 (O_750,N_18635,N_19666);
nor UO_751 (O_751,N_16088,N_18477);
nand UO_752 (O_752,N_16631,N_18574);
nand UO_753 (O_753,N_18533,N_17088);
or UO_754 (O_754,N_16880,N_16383);
nand UO_755 (O_755,N_19740,N_16373);
nand UO_756 (O_756,N_16155,N_18193);
nor UO_757 (O_757,N_17399,N_17657);
or UO_758 (O_758,N_16392,N_17921);
or UO_759 (O_759,N_17435,N_17886);
nand UO_760 (O_760,N_19282,N_15719);
and UO_761 (O_761,N_19726,N_17863);
and UO_762 (O_762,N_15146,N_19819);
nand UO_763 (O_763,N_18356,N_19035);
xor UO_764 (O_764,N_15612,N_15548);
or UO_765 (O_765,N_18019,N_18331);
and UO_766 (O_766,N_19474,N_15905);
nand UO_767 (O_767,N_19638,N_19884);
nor UO_768 (O_768,N_16405,N_17672);
nand UO_769 (O_769,N_16726,N_19650);
and UO_770 (O_770,N_16213,N_18319);
nand UO_771 (O_771,N_18964,N_18735);
or UO_772 (O_772,N_17625,N_15991);
or UO_773 (O_773,N_16414,N_15909);
or UO_774 (O_774,N_17907,N_17510);
xnor UO_775 (O_775,N_17824,N_19265);
nor UO_776 (O_776,N_15361,N_18143);
nor UO_777 (O_777,N_18565,N_16285);
nand UO_778 (O_778,N_16035,N_17523);
xnor UO_779 (O_779,N_17673,N_15044);
or UO_780 (O_780,N_16337,N_15406);
nor UO_781 (O_781,N_16559,N_19582);
or UO_782 (O_782,N_16790,N_17426);
nand UO_783 (O_783,N_19619,N_18737);
and UO_784 (O_784,N_15254,N_16734);
nor UO_785 (O_785,N_16853,N_16479);
xnor UO_786 (O_786,N_16841,N_17268);
and UO_787 (O_787,N_17323,N_17493);
nor UO_788 (O_788,N_18079,N_18827);
and UO_789 (O_789,N_18829,N_15875);
nand UO_790 (O_790,N_17056,N_18806);
or UO_791 (O_791,N_19440,N_16525);
nand UO_792 (O_792,N_19313,N_19398);
nor UO_793 (O_793,N_18045,N_18616);
and UO_794 (O_794,N_17059,N_18885);
and UO_795 (O_795,N_15701,N_15903);
nor UO_796 (O_796,N_15253,N_15830);
nand UO_797 (O_797,N_16157,N_16071);
or UO_798 (O_798,N_15856,N_19724);
and UO_799 (O_799,N_18847,N_15102);
or UO_800 (O_800,N_18135,N_15805);
or UO_801 (O_801,N_16669,N_16766);
xor UO_802 (O_802,N_15563,N_16774);
and UO_803 (O_803,N_16048,N_19963);
nand UO_804 (O_804,N_18712,N_15633);
xnor UO_805 (O_805,N_16049,N_15171);
or UO_806 (O_806,N_15486,N_16084);
xor UO_807 (O_807,N_16127,N_16789);
xor UO_808 (O_808,N_15623,N_18628);
and UO_809 (O_809,N_18210,N_15558);
or UO_810 (O_810,N_19966,N_16562);
or UO_811 (O_811,N_15478,N_17616);
nor UO_812 (O_812,N_19457,N_17753);
xnor UO_813 (O_813,N_17708,N_17309);
and UO_814 (O_814,N_19558,N_18133);
nor UO_815 (O_815,N_18926,N_15788);
nand UO_816 (O_816,N_17904,N_19030);
and UO_817 (O_817,N_16581,N_19635);
nor UO_818 (O_818,N_17443,N_19719);
nor UO_819 (O_819,N_17291,N_15496);
nor UO_820 (O_820,N_17968,N_19052);
nand UO_821 (O_821,N_15163,N_18693);
nand UO_822 (O_822,N_19651,N_17275);
and UO_823 (O_823,N_18309,N_15161);
or UO_824 (O_824,N_19705,N_17551);
and UO_825 (O_825,N_19790,N_18673);
nor UO_826 (O_826,N_17515,N_18783);
nand UO_827 (O_827,N_19967,N_16901);
and UO_828 (O_828,N_18182,N_15578);
nand UO_829 (O_829,N_16676,N_16570);
or UO_830 (O_830,N_17628,N_15451);
nand UO_831 (O_831,N_19074,N_19529);
or UO_832 (O_832,N_17977,N_17300);
nand UO_833 (O_833,N_19332,N_17836);
nand UO_834 (O_834,N_19228,N_19707);
nor UO_835 (O_835,N_18701,N_17791);
and UO_836 (O_836,N_17693,N_18780);
nand UO_837 (O_837,N_18898,N_16162);
or UO_838 (O_838,N_16251,N_16605);
nor UO_839 (O_839,N_18863,N_19086);
or UO_840 (O_840,N_18504,N_15942);
nand UO_841 (O_841,N_18166,N_16919);
xnor UO_842 (O_842,N_18903,N_16150);
or UO_843 (O_843,N_18720,N_19232);
and UO_844 (O_844,N_17864,N_18302);
nor UO_845 (O_845,N_16110,N_18174);
nor UO_846 (O_846,N_15649,N_17512);
nor UO_847 (O_847,N_16200,N_15782);
or UO_848 (O_848,N_18710,N_16421);
or UO_849 (O_849,N_15681,N_15025);
nor UO_850 (O_850,N_15790,N_16516);
nor UO_851 (O_851,N_17891,N_18412);
or UO_852 (O_852,N_16224,N_19368);
or UO_853 (O_853,N_16627,N_18380);
or UO_854 (O_854,N_16125,N_15270);
nor UO_855 (O_855,N_17735,N_19252);
nand UO_856 (O_856,N_18161,N_19470);
or UO_857 (O_857,N_17765,N_19508);
nand UO_858 (O_858,N_17499,N_17757);
nand UO_859 (O_859,N_19359,N_16448);
xor UO_860 (O_860,N_18192,N_15019);
xor UO_861 (O_861,N_17413,N_17555);
nor UO_862 (O_862,N_18862,N_18978);
and UO_863 (O_863,N_18611,N_17307);
nor UO_864 (O_864,N_17878,N_15405);
nand UO_865 (O_865,N_16519,N_18805);
nand UO_866 (O_866,N_16625,N_16612);
nor UO_867 (O_867,N_16592,N_17935);
xnor UO_868 (O_868,N_19243,N_15524);
nand UO_869 (O_869,N_19395,N_19518);
or UO_870 (O_870,N_15768,N_16261);
nor UO_871 (O_871,N_18870,N_16441);
and UO_872 (O_872,N_19960,N_15464);
nor UO_873 (O_873,N_17206,N_17594);
xor UO_874 (O_874,N_19162,N_17224);
nand UO_875 (O_875,N_15988,N_16708);
xnor UO_876 (O_876,N_16404,N_19624);
or UO_877 (O_877,N_16115,N_17867);
nand UO_878 (O_878,N_19639,N_19308);
nor UO_879 (O_879,N_15838,N_17677);
and UO_880 (O_880,N_18329,N_16530);
nand UO_881 (O_881,N_17395,N_18246);
and UO_882 (O_882,N_15197,N_19459);
xor UO_883 (O_883,N_16573,N_15112);
nor UO_884 (O_884,N_17373,N_19467);
nor UO_885 (O_885,N_19672,N_19958);
xor UO_886 (O_886,N_19170,N_19318);
xor UO_887 (O_887,N_18981,N_19472);
or UO_888 (O_888,N_19060,N_18378);
and UO_889 (O_889,N_18449,N_19779);
and UO_890 (O_890,N_17636,N_17704);
nor UO_891 (O_891,N_18625,N_19578);
nor UO_892 (O_892,N_19255,N_19713);
or UO_893 (O_893,N_17068,N_19977);
or UO_894 (O_894,N_17115,N_19337);
and UO_895 (O_895,N_19357,N_17528);
nor UO_896 (O_896,N_18454,N_19438);
or UO_897 (O_897,N_17495,N_19061);
nor UO_898 (O_898,N_17805,N_18516);
xnor UO_899 (O_899,N_17098,N_17794);
and UO_900 (O_900,N_15468,N_15448);
xor UO_901 (O_901,N_18594,N_15963);
xor UO_902 (O_902,N_16482,N_16356);
nand UO_903 (O_903,N_17434,N_16904);
or UO_904 (O_904,N_16042,N_18345);
nand UO_905 (O_905,N_19404,N_19602);
xnor UO_906 (O_906,N_15138,N_17486);
nand UO_907 (O_907,N_17897,N_17077);
nand UO_908 (O_908,N_15087,N_19708);
nand UO_909 (O_909,N_18542,N_15278);
nor UO_910 (O_910,N_17796,N_16700);
xnor UO_911 (O_911,N_18690,N_19118);
nand UO_912 (O_912,N_19645,N_16504);
xnor UO_913 (O_913,N_18833,N_18008);
nand UO_914 (O_914,N_18383,N_17577);
nand UO_915 (O_915,N_15479,N_19511);
nor UO_916 (O_916,N_16050,N_16532);
nand UO_917 (O_917,N_16288,N_17652);
and UO_918 (O_918,N_16784,N_18547);
nand UO_919 (O_919,N_18215,N_19129);
nand UO_920 (O_920,N_19432,N_17349);
or UO_921 (O_921,N_17831,N_15635);
xnor UO_922 (O_922,N_19212,N_16303);
or UO_923 (O_923,N_18993,N_18360);
xnor UO_924 (O_924,N_17429,N_19839);
nor UO_925 (O_925,N_18938,N_16258);
or UO_926 (O_926,N_17858,N_15978);
xor UO_927 (O_927,N_19018,N_18377);
or UO_928 (O_928,N_19888,N_18853);
and UO_929 (O_929,N_17979,N_15323);
nand UO_930 (O_930,N_18566,N_18042);
xor UO_931 (O_931,N_15041,N_19625);
and UO_932 (O_932,N_16266,N_16489);
nor UO_933 (O_933,N_16449,N_19424);
nor UO_934 (O_934,N_16363,N_15581);
nor UO_935 (O_935,N_18167,N_18949);
nor UO_936 (O_936,N_19378,N_16948);
xnor UO_937 (O_937,N_17686,N_17320);
and UO_938 (O_938,N_19091,N_19388);
xor UO_939 (O_939,N_19152,N_17496);
xor UO_940 (O_940,N_15148,N_16465);
nand UO_941 (O_941,N_18707,N_17647);
or UO_942 (O_942,N_15024,N_17959);
or UO_943 (O_943,N_16552,N_18977);
or UO_944 (O_944,N_19865,N_18264);
and UO_945 (O_945,N_16801,N_18336);
xor UO_946 (O_946,N_16218,N_18147);
and UO_947 (O_947,N_19961,N_19264);
or UO_948 (O_948,N_17454,N_19874);
or UO_949 (O_949,N_16242,N_19492);
and UO_950 (O_950,N_16474,N_18247);
xor UO_951 (O_951,N_15252,N_16346);
xnor UO_952 (O_952,N_19862,N_15168);
or UO_953 (O_953,N_15718,N_15739);
nand UO_954 (O_954,N_16547,N_19372);
or UO_955 (O_955,N_15902,N_17950);
or UO_956 (O_956,N_15661,N_19555);
nand UO_957 (O_957,N_19445,N_15596);
xnor UO_958 (O_958,N_16597,N_17557);
and UO_959 (O_959,N_16415,N_17611);
or UO_960 (O_960,N_17746,N_15770);
xor UO_961 (O_961,N_19853,N_16881);
xnor UO_962 (O_962,N_15572,N_15286);
nand UO_963 (O_963,N_16909,N_16407);
nand UO_964 (O_964,N_15165,N_16401);
nand UO_965 (O_965,N_15722,N_18688);
xor UO_966 (O_966,N_15604,N_19144);
xor UO_967 (O_967,N_16739,N_18952);
nor UO_968 (O_968,N_19611,N_18963);
nand UO_969 (O_969,N_17483,N_16535);
nor UO_970 (O_970,N_15608,N_17505);
nand UO_971 (O_971,N_19025,N_16210);
nor UO_972 (O_972,N_19895,N_18586);
nor UO_973 (O_973,N_18168,N_17632);
nor UO_974 (O_974,N_16196,N_18090);
and UO_975 (O_975,N_17028,N_19031);
nor UO_976 (O_976,N_18802,N_17064);
and UO_977 (O_977,N_18632,N_18337);
and UO_978 (O_978,N_18819,N_16505);
and UO_979 (O_979,N_16807,N_18434);
nand UO_980 (O_980,N_19882,N_18942);
and UO_981 (O_981,N_16317,N_17255);
and UO_982 (O_982,N_19141,N_16871);
or UO_983 (O_983,N_15659,N_15567);
nand UO_984 (O_984,N_16108,N_16754);
nor UO_985 (O_985,N_16362,N_19816);
nand UO_986 (O_986,N_15063,N_17235);
nor UO_987 (O_987,N_19633,N_19951);
and UO_988 (O_988,N_15210,N_17795);
xor UO_989 (O_989,N_15415,N_18075);
xnor UO_990 (O_990,N_15527,N_17062);
and UO_991 (O_991,N_15514,N_16690);
or UO_992 (O_992,N_19580,N_16169);
nand UO_993 (O_993,N_16243,N_18398);
xor UO_994 (O_994,N_16276,N_17313);
xnor UO_995 (O_995,N_19320,N_18584);
xor UO_996 (O_996,N_17384,N_16846);
or UO_997 (O_997,N_17992,N_19983);
nand UO_998 (O_998,N_17438,N_17650);
nor UO_999 (O_999,N_16705,N_19418);
nand UO_1000 (O_1000,N_19276,N_16293);
or UO_1001 (O_1001,N_16128,N_18010);
xor UO_1002 (O_1002,N_16019,N_16987);
or UO_1003 (O_1003,N_19304,N_18608);
and UO_1004 (O_1004,N_16055,N_17030);
xor UO_1005 (O_1005,N_18985,N_19570);
and UO_1006 (O_1006,N_15605,N_18245);
or UO_1007 (O_1007,N_15557,N_17558);
nor UO_1008 (O_1008,N_16852,N_16148);
xnor UO_1009 (O_1009,N_18634,N_15655);
nand UO_1010 (O_1010,N_15503,N_18719);
nand UO_1011 (O_1011,N_15721,N_17713);
and UO_1012 (O_1012,N_15402,N_16634);
xor UO_1013 (O_1013,N_17702,N_18452);
or UO_1014 (O_1014,N_17140,N_15352);
and UO_1015 (O_1015,N_18761,N_16120);
nand UO_1016 (O_1016,N_16101,N_18117);
and UO_1017 (O_1017,N_18484,N_16464);
or UO_1018 (O_1018,N_15868,N_19741);
xnor UO_1019 (O_1019,N_15621,N_16032);
nor UO_1020 (O_1020,N_16079,N_16177);
nand UO_1021 (O_1021,N_16176,N_16498);
or UO_1022 (O_1022,N_17165,N_15720);
nor UO_1023 (O_1023,N_19435,N_15309);
nor UO_1024 (O_1024,N_19694,N_17020);
nor UO_1025 (O_1025,N_19932,N_18883);
nor UO_1026 (O_1026,N_18836,N_17358);
nor UO_1027 (O_1027,N_16600,N_17390);
nor UO_1028 (O_1028,N_15920,N_15205);
nor UO_1029 (O_1029,N_16697,N_19894);
nand UO_1030 (O_1030,N_17394,N_17446);
nand UO_1031 (O_1031,N_17919,N_18482);
nor UO_1032 (O_1032,N_17593,N_16762);
and UO_1033 (O_1033,N_16007,N_15281);
nor UO_1034 (O_1034,N_19267,N_18407);
or UO_1035 (O_1035,N_19040,N_17911);
nor UO_1036 (O_1036,N_17404,N_18083);
and UO_1037 (O_1037,N_16860,N_18563);
or UO_1038 (O_1038,N_17145,N_18173);
or UO_1039 (O_1039,N_18663,N_16928);
xnor UO_1040 (O_1040,N_15708,N_19767);
nand UO_1041 (O_1041,N_17789,N_19833);
and UO_1042 (O_1042,N_16868,N_19851);
xor UO_1043 (O_1043,N_18803,N_16912);
nor UO_1044 (O_1044,N_15395,N_16606);
or UO_1045 (O_1045,N_17585,N_18301);
or UO_1046 (O_1046,N_15442,N_15520);
xor UO_1047 (O_1047,N_17788,N_18470);
nand UO_1048 (O_1048,N_16015,N_15300);
xor UO_1049 (O_1049,N_17751,N_19485);
xnor UO_1050 (O_1050,N_16765,N_18015);
xnor UO_1051 (O_1051,N_15221,N_17106);
xnor UO_1052 (O_1052,N_15236,N_18099);
nand UO_1053 (O_1053,N_18122,N_18955);
nor UO_1054 (O_1054,N_18521,N_16699);
nand UO_1055 (O_1055,N_19208,N_17944);
or UO_1056 (O_1056,N_16643,N_17814);
nand UO_1057 (O_1057,N_15038,N_15276);
xnor UO_1058 (O_1058,N_16212,N_16861);
and UO_1059 (O_1059,N_16903,N_18831);
xnor UO_1060 (O_1060,N_15698,N_15964);
and UO_1061 (O_1061,N_15618,N_16332);
nor UO_1062 (O_1062,N_15874,N_19366);
nor UO_1063 (O_1063,N_17910,N_16207);
or UO_1064 (O_1064,N_18203,N_15419);
nor UO_1065 (O_1065,N_19561,N_15684);
or UO_1066 (O_1066,N_16072,N_17784);
nor UO_1067 (O_1067,N_18617,N_18859);
xnor UO_1068 (O_1068,N_16884,N_16069);
xor UO_1069 (O_1069,N_18156,N_15573);
nand UO_1070 (O_1070,N_18620,N_19654);
nor UO_1071 (O_1071,N_15933,N_19755);
nand UO_1072 (O_1072,N_19804,N_17595);
and UO_1073 (O_1073,N_17299,N_16054);
and UO_1074 (O_1074,N_16970,N_16036);
nand UO_1075 (O_1075,N_18459,N_17587);
nand UO_1076 (O_1076,N_16286,N_16391);
or UO_1077 (O_1077,N_15508,N_16225);
xnor UO_1078 (O_1078,N_15628,N_19137);
xor UO_1079 (O_1079,N_19373,N_17502);
xor UO_1080 (O_1080,N_17664,N_17400);
nand UO_1081 (O_1081,N_16713,N_18020);
and UO_1082 (O_1082,N_15037,N_15738);
xor UO_1083 (O_1083,N_16704,N_15417);
and UO_1084 (O_1084,N_16364,N_17578);
and UO_1085 (O_1085,N_17829,N_15450);
or UO_1086 (O_1086,N_16579,N_19835);
or UO_1087 (O_1087,N_17820,N_15330);
xnor UO_1088 (O_1088,N_16571,N_18076);
or UO_1089 (O_1089,N_17675,N_18839);
xor UO_1090 (O_1090,N_19020,N_18120);
or UO_1091 (O_1091,N_18087,N_16237);
nand UO_1092 (O_1092,N_16158,N_15374);
xor UO_1093 (O_1093,N_17000,N_15561);
nand UO_1094 (O_1094,N_17398,N_19355);
or UO_1095 (O_1095,N_18585,N_15663);
nor UO_1096 (O_1096,N_16253,N_15588);
nor UO_1097 (O_1097,N_18366,N_17017);
and UO_1098 (O_1098,N_15842,N_19039);
or UO_1099 (O_1099,N_19085,N_16639);
or UO_1100 (O_1100,N_19151,N_16867);
nor UO_1101 (O_1101,N_17783,N_15091);
and UO_1102 (O_1102,N_15184,N_19480);
or UO_1103 (O_1103,N_16075,N_17402);
nor UO_1104 (O_1104,N_19757,N_15436);
and UO_1105 (O_1105,N_15700,N_15695);
xnor UO_1106 (O_1106,N_18892,N_15216);
nand UO_1107 (O_1107,N_15523,N_17804);
xor UO_1108 (O_1108,N_15365,N_19982);
nand UO_1109 (O_1109,N_17699,N_17643);
xnor UO_1110 (O_1110,N_17209,N_16670);
and UO_1111 (O_1111,N_19192,N_18818);
and UO_1112 (O_1112,N_15521,N_19166);
nand UO_1113 (O_1113,N_16342,N_15332);
nand UO_1114 (O_1114,N_18889,N_19802);
nand UO_1115 (O_1115,N_16295,N_18912);
and UO_1116 (O_1116,N_19901,N_17655);
and UO_1117 (O_1117,N_15110,N_18591);
nor UO_1118 (O_1118,N_16727,N_16802);
nor UO_1119 (O_1119,N_17540,N_15562);
nor UO_1120 (O_1120,N_15598,N_17641);
nor UO_1121 (O_1121,N_15290,N_18753);
or UO_1122 (O_1122,N_19962,N_17902);
xor UO_1123 (O_1123,N_17569,N_18251);
and UO_1124 (O_1124,N_15735,N_17818);
nand UO_1125 (O_1125,N_18577,N_17382);
xnor UO_1126 (O_1126,N_15157,N_16780);
nand UO_1127 (O_1127,N_18715,N_17676);
xnor UO_1128 (O_1128,N_18488,N_17980);
or UO_1129 (O_1129,N_15823,N_16665);
or UO_1130 (O_1130,N_18134,N_19627);
nand UO_1131 (O_1131,N_16900,N_16947);
nor UO_1132 (O_1132,N_15064,N_19004);
and UO_1133 (O_1133,N_16934,N_18259);
and UO_1134 (O_1134,N_15835,N_18274);
or UO_1135 (O_1135,N_15409,N_18786);
xnor UO_1136 (O_1136,N_15357,N_19892);
nand UO_1137 (O_1137,N_16828,N_18241);
and UO_1138 (O_1138,N_15347,N_16650);
and UO_1139 (O_1139,N_15796,N_17153);
or UO_1140 (O_1140,N_15828,N_15586);
xor UO_1141 (O_1141,N_17884,N_15927);
or UO_1142 (O_1142,N_19553,N_18468);
xnor UO_1143 (O_1143,N_16485,N_16599);
and UO_1144 (O_1144,N_17842,N_16409);
and UO_1145 (O_1145,N_15629,N_17045);
nand UO_1146 (O_1146,N_19744,N_19277);
nor UO_1147 (O_1147,N_15139,N_16723);
nand UO_1148 (O_1148,N_15692,N_15893);
and UO_1149 (O_1149,N_15717,N_19952);
and UO_1150 (O_1150,N_19859,N_16420);
or UO_1151 (O_1151,N_16254,N_19288);
xnor UO_1152 (O_1152,N_19599,N_16152);
nor UO_1153 (O_1153,N_17768,N_16922);
and UO_1154 (O_1154,N_18789,N_17080);
nor UO_1155 (O_1155,N_17264,N_16682);
nand UO_1156 (O_1156,N_15783,N_17521);
or UO_1157 (O_1157,N_19326,N_16209);
and UO_1158 (O_1158,N_16012,N_18060);
or UO_1159 (O_1159,N_15243,N_17755);
or UO_1160 (O_1160,N_19247,N_18752);
nand UO_1161 (O_1161,N_19127,N_16816);
or UO_1162 (O_1162,N_18598,N_16160);
and UO_1163 (O_1163,N_19703,N_18856);
or UO_1164 (O_1164,N_15288,N_17974);
nand UO_1165 (O_1165,N_19696,N_15244);
nor UO_1166 (O_1166,N_19920,N_16074);
nand UO_1167 (O_1167,N_16764,N_16496);
nand UO_1168 (O_1168,N_16038,N_16308);
nand UO_1169 (O_1169,N_15488,N_17559);
nor UO_1170 (O_1170,N_17798,N_18084);
and UO_1171 (O_1171,N_16508,N_18666);
and UO_1172 (O_1172,N_17646,N_16675);
and UO_1173 (O_1173,N_16467,N_16355);
xor UO_1174 (O_1174,N_19704,N_19164);
and UO_1175 (O_1175,N_17726,N_19452);
nor UO_1176 (O_1176,N_17561,N_16361);
nand UO_1177 (O_1177,N_18919,N_16826);
or UO_1178 (O_1178,N_17546,N_16782);
xnor UO_1179 (O_1179,N_19837,N_16733);
or UO_1180 (O_1180,N_18017,N_15497);
nand UO_1181 (O_1181,N_15430,N_19108);
nor UO_1182 (O_1182,N_17503,N_16544);
or UO_1183 (O_1183,N_17167,N_18226);
xnor UO_1184 (O_1184,N_17912,N_16236);
xor UO_1185 (O_1185,N_16492,N_19715);
xor UO_1186 (O_1186,N_19150,N_16568);
or UO_1187 (O_1187,N_15609,N_18925);
xor UO_1188 (O_1188,N_16963,N_17423);
xnor UO_1189 (O_1189,N_17550,N_15389);
xor UO_1190 (O_1190,N_16795,N_19145);
nand UO_1191 (O_1191,N_15327,N_19840);
and UO_1192 (O_1192,N_15537,N_19184);
or UO_1193 (O_1193,N_15819,N_19875);
nand UO_1194 (O_1194,N_18600,N_15424);
nor UO_1195 (O_1195,N_15095,N_16463);
or UO_1196 (O_1196,N_17785,N_15945);
and UO_1197 (O_1197,N_15099,N_16914);
xnor UO_1198 (O_1198,N_19820,N_15580);
nor UO_1199 (O_1199,N_16287,N_18479);
xnor UO_1200 (O_1200,N_18239,N_19509);
xnor UO_1201 (O_1201,N_19773,N_15108);
nor UO_1202 (O_1202,N_19917,N_19993);
and UO_1203 (O_1203,N_15965,N_19369);
and UO_1204 (O_1204,N_17462,N_18648);
nor UO_1205 (O_1205,N_18485,N_16123);
xor UO_1206 (O_1206,N_19809,N_15646);
or UO_1207 (O_1207,N_19249,N_18966);
and UO_1208 (O_1208,N_16189,N_15167);
xnor UO_1209 (O_1209,N_19088,N_17381);
or UO_1210 (O_1210,N_15032,N_19098);
xnor UO_1211 (O_1211,N_19953,N_17631);
nor UO_1212 (O_1212,N_15766,N_16632);
xor UO_1213 (O_1213,N_16744,N_17955);
xnor UO_1214 (O_1214,N_16893,N_17975);
or UO_1215 (O_1215,N_19572,N_17368);
or UO_1216 (O_1216,N_15619,N_15622);
xnor UO_1217 (O_1217,N_15703,N_16359);
nand UO_1218 (O_1218,N_15065,N_19515);
xnor UO_1219 (O_1219,N_15452,N_19514);
xor UO_1220 (O_1220,N_16974,N_16767);
nor UO_1221 (O_1221,N_17762,N_17660);
or UO_1222 (O_1222,N_18284,N_19101);
nand UO_1223 (O_1223,N_18165,N_19268);
nand UO_1224 (O_1224,N_17839,N_17697);
and UO_1225 (O_1225,N_18810,N_19538);
nand UO_1226 (O_1226,N_19182,N_17018);
nor UO_1227 (O_1227,N_18653,N_15105);
nor UO_1228 (O_1228,N_16043,N_18579);
or UO_1229 (O_1229,N_18009,N_15445);
nor UO_1230 (O_1230,N_15851,N_18058);
or UO_1231 (O_1231,N_15306,N_19487);
and UO_1232 (O_1232,N_18865,N_18487);
or UO_1233 (O_1233,N_17701,N_16013);
and UO_1234 (O_1234,N_18559,N_16192);
nor UO_1235 (O_1235,N_18127,N_17332);
and UO_1236 (O_1236,N_17943,N_19924);
xor UO_1237 (O_1237,N_18583,N_16471);
or UO_1238 (O_1238,N_17760,N_17575);
and UO_1239 (O_1239,N_16567,N_18733);
xnor UO_1240 (O_1240,N_15132,N_15544);
or UO_1241 (O_1241,N_17534,N_16000);
or UO_1242 (O_1242,N_16331,N_17036);
xnor UO_1243 (O_1243,N_19084,N_17776);
nand UO_1244 (O_1244,N_17739,N_16760);
or UO_1245 (O_1245,N_16351,N_15084);
or UO_1246 (O_1246,N_15660,N_17032);
and UO_1247 (O_1247,N_18729,N_18011);
nand UO_1248 (O_1248,N_15914,N_16862);
and UO_1249 (O_1249,N_18212,N_15850);
nor UO_1250 (O_1250,N_17334,N_15753);
or UO_1251 (O_1251,N_18128,N_17690);
xnor UO_1252 (O_1252,N_15418,N_17338);
xor UO_1253 (O_1253,N_15809,N_17039);
and UO_1254 (O_1254,N_18237,N_17793);
xnor UO_1255 (O_1255,N_15620,N_15546);
or UO_1256 (O_1256,N_17029,N_16939);
or UO_1257 (O_1257,N_19094,N_16629);
xnor UO_1258 (O_1258,N_16741,N_15944);
and UO_1259 (O_1259,N_15582,N_19913);
or UO_1260 (O_1260,N_17414,N_18762);
xnor UO_1261 (O_1261,N_18231,N_16652);
nor UO_1262 (O_1262,N_19764,N_19945);
xor UO_1263 (O_1263,N_15045,N_15957);
nor UO_1264 (O_1264,N_16172,N_16746);
nor UO_1265 (O_1265,N_17103,N_17458);
nor UO_1266 (O_1266,N_17057,N_19805);
xor UO_1267 (O_1267,N_19120,N_19029);
or UO_1268 (O_1268,N_15547,N_15081);
nand UO_1269 (O_1269,N_17876,N_15043);
and UO_1270 (O_1270,N_16958,N_15857);
or UO_1271 (O_1271,N_15816,N_17608);
xnor UO_1272 (O_1272,N_17261,N_17035);
and UO_1273 (O_1273,N_17769,N_19674);
and UO_1274 (O_1274,N_17984,N_18575);
nand UO_1275 (O_1275,N_18606,N_16433);
and UO_1276 (O_1276,N_15375,N_17662);
nand UO_1277 (O_1277,N_16259,N_19842);
nand UO_1278 (O_1278,N_17156,N_16031);
or UO_1279 (O_1279,N_19617,N_18835);
and UO_1280 (O_1280,N_15542,N_16163);
nor UO_1281 (O_1281,N_16777,N_19646);
xor UO_1282 (O_1282,N_17015,N_19883);
xor UO_1283 (O_1283,N_16910,N_17085);
xnor UO_1284 (O_1284,N_17102,N_15069);
and UO_1285 (O_1285,N_17811,N_16991);
and UO_1286 (O_1286,N_19329,N_18821);
or UO_1287 (O_1287,N_16438,N_19716);
xnor UO_1288 (O_1288,N_16737,N_19577);
and UO_1289 (O_1289,N_18013,N_19743);
or UO_1290 (O_1290,N_17725,N_18111);
nand UO_1291 (O_1291,N_19434,N_15861);
or UO_1292 (O_1292,N_15334,N_16601);
nor UO_1293 (O_1293,N_15109,N_18050);
nor UO_1294 (O_1294,N_18418,N_19322);
nor UO_1295 (O_1295,N_17759,N_18708);
or UO_1296 (O_1296,N_18599,N_15792);
nand UO_1297 (O_1297,N_18288,N_18091);
nor UO_1298 (O_1298,N_15891,N_17005);
nand UO_1299 (O_1299,N_16223,N_16611);
nand UO_1300 (O_1300,N_17571,N_17335);
nand UO_1301 (O_1301,N_15691,N_15339);
and UO_1302 (O_1302,N_15295,N_19106);
or UO_1303 (O_1303,N_16025,N_18293);
nor UO_1304 (O_1304,N_19643,N_17294);
and UO_1305 (O_1305,N_17179,N_16133);
xor UO_1306 (O_1306,N_19701,N_18154);
xnor UO_1307 (O_1307,N_18510,N_16073);
or UO_1308 (O_1308,N_17553,N_16114);
or UO_1309 (O_1309,N_19775,N_19821);
xnor UO_1310 (O_1310,N_19693,N_17916);
nor UO_1311 (O_1311,N_16598,N_16701);
nand UO_1312 (O_1312,N_15012,N_19583);
nand UO_1313 (O_1313,N_16507,N_19425);
and UO_1314 (O_1314,N_15937,N_17019);
xor UO_1315 (O_1315,N_15399,N_16960);
xor UO_1316 (O_1316,N_19370,N_16720);
nor UO_1317 (O_1317,N_15487,N_17158);
and UO_1318 (O_1318,N_19568,N_18238);
or UO_1319 (O_1319,N_15056,N_18306);
nor UO_1320 (O_1320,N_18136,N_19925);
or UO_1321 (O_1321,N_15231,N_16382);
and UO_1322 (O_1322,N_19647,N_16434);
or UO_1323 (O_1323,N_18362,N_17256);
xor UO_1324 (O_1324,N_19785,N_19552);
nand UO_1325 (O_1325,N_15443,N_15251);
and UO_1326 (O_1326,N_17180,N_19073);
and UO_1327 (O_1327,N_16480,N_16424);
xnor UO_1328 (O_1328,N_17743,N_15319);
and UO_1329 (O_1329,N_15656,N_19482);
or UO_1330 (O_1330,N_17229,N_17821);
nand UO_1331 (O_1331,N_19269,N_17613);
and UO_1332 (O_1332,N_17750,N_16946);
nand UO_1333 (O_1333,N_17174,N_16326);
or UO_1334 (O_1334,N_16943,N_16955);
nand UO_1335 (O_1335,N_15360,N_15143);
or UO_1336 (O_1336,N_17391,N_17573);
nor UO_1337 (O_1337,N_17298,N_19947);
nor UO_1338 (O_1338,N_19603,N_16594);
nand UO_1339 (O_1339,N_18872,N_19272);
and UO_1340 (O_1340,N_16569,N_15149);
or UO_1341 (O_1341,N_16182,N_19739);
nand UO_1342 (O_1342,N_18409,N_18420);
and UO_1343 (O_1343,N_18840,N_15490);
or UO_1344 (O_1344,N_18052,N_15465);
nand UO_1345 (O_1345,N_15345,N_19161);
xnor UO_1346 (O_1346,N_16811,N_18472);
nor UO_1347 (O_1347,N_17375,N_15207);
xor UO_1348 (O_1348,N_18401,N_18465);
nor UO_1349 (O_1349,N_15483,N_17339);
or UO_1350 (O_1350,N_16694,N_19493);
and UO_1351 (O_1351,N_17960,N_18999);
nand UO_1352 (O_1352,N_16280,N_18034);
and UO_1353 (O_1353,N_17802,N_17883);
xnor UO_1354 (O_1354,N_17627,N_16283);
and UO_1355 (O_1355,N_17487,N_17311);
and UO_1356 (O_1356,N_17427,N_15641);
or UO_1357 (O_1357,N_16185,N_16336);
nor UO_1358 (O_1358,N_19657,N_17689);
nand UO_1359 (O_1359,N_15846,N_18249);
nand UO_1360 (O_1360,N_18002,N_17333);
nand UO_1361 (O_1361,N_16998,N_15781);
xor UO_1362 (O_1362,N_19873,N_15888);
and UO_1363 (O_1363,N_18768,N_15728);
or UO_1364 (O_1364,N_18890,N_19844);
xnor UO_1365 (O_1365,N_18759,N_16387);
nor UO_1366 (O_1366,N_19488,N_15501);
nor UO_1367 (O_1367,N_19014,N_19283);
nor UO_1368 (O_1368,N_18085,N_17617);
nand UO_1369 (O_1369,N_15061,N_19426);
nor UO_1370 (O_1370,N_16403,N_19984);
nor UO_1371 (O_1371,N_16565,N_18602);
and UO_1372 (O_1372,N_17411,N_18934);
nand UO_1373 (O_1373,N_17254,N_18387);
or UO_1374 (O_1374,N_16967,N_16298);
nor UO_1375 (O_1375,N_18201,N_18431);
nand UO_1376 (O_1376,N_19036,N_15904);
xnor UO_1377 (O_1377,N_17504,N_15889);
and UO_1378 (O_1378,N_18554,N_17096);
xnor UO_1379 (O_1379,N_18451,N_19688);
and UO_1380 (O_1380,N_19100,N_15177);
nor UO_1381 (O_1381,N_17630,N_19765);
and UO_1382 (O_1382,N_15840,N_16250);
or UO_1383 (O_1383,N_19251,N_15780);
nand UO_1384 (O_1384,N_18018,N_17489);
nand UO_1385 (O_1385,N_18947,N_18341);
or UO_1386 (O_1386,N_18637,N_18155);
xor UO_1387 (O_1387,N_18417,N_19899);
or UO_1388 (O_1388,N_16164,N_19845);
nand UO_1389 (O_1389,N_15884,N_16703);
and UO_1390 (O_1390,N_19559,N_16307);
xor UO_1391 (O_1391,N_17937,N_16792);
nor UO_1392 (O_1392,N_18954,N_18140);
or UO_1393 (O_1393,N_19234,N_18082);
or UO_1394 (O_1394,N_15741,N_17251);
and UO_1395 (O_1395,N_17812,N_18906);
or UO_1396 (O_1396,N_16640,N_16027);
nand UO_1397 (O_1397,N_15571,N_18732);
or UO_1398 (O_1398,N_15219,N_15648);
xnor UO_1399 (O_1399,N_18561,N_17929);
xor UO_1400 (O_1400,N_19957,N_18385);
nand UO_1401 (O_1401,N_16834,N_16139);
and UO_1402 (O_1402,N_17606,N_16451);
and UO_1403 (O_1403,N_17810,N_16481);
xor UO_1404 (O_1404,N_15584,N_17447);
and UO_1405 (O_1405,N_15127,N_17284);
and UO_1406 (O_1406,N_15870,N_18386);
or UO_1407 (O_1407,N_19242,N_19218);
or UO_1408 (O_1408,N_19616,N_15470);
nand UO_1409 (O_1409,N_15074,N_18660);
nand UO_1410 (O_1410,N_17848,N_15667);
nand UO_1411 (O_1411,N_15082,N_17917);
nor UO_1412 (O_1412,N_17369,N_16962);
and UO_1413 (O_1413,N_16214,N_17623);
and UO_1414 (O_1414,N_16056,N_18025);
and UO_1415 (O_1415,N_17401,N_17947);
or UO_1416 (O_1416,N_19055,N_16129);
xnor UO_1417 (O_1417,N_15200,N_15595);
and UO_1418 (O_1418,N_18395,N_17792);
or UO_1419 (O_1419,N_16033,N_16895);
xnor UO_1420 (O_1420,N_18438,N_17327);
xor UO_1421 (O_1421,N_19941,N_15335);
xor UO_1422 (O_1422,N_16083,N_15248);
nand UO_1423 (O_1423,N_18924,N_19889);
nor UO_1424 (O_1424,N_15625,N_18526);
or UO_1425 (O_1425,N_15412,N_16791);
or UO_1426 (O_1426,N_17942,N_17290);
nand UO_1427 (O_1427,N_16457,N_19531);
nand UO_1428 (O_1428,N_17854,N_18458);
nand UO_1429 (O_1429,N_18442,N_19782);
xor UO_1430 (O_1430,N_17049,N_17051);
and UO_1431 (O_1431,N_16418,N_18867);
nor UO_1432 (O_1432,N_16208,N_18473);
nand UO_1433 (O_1433,N_16520,N_16725);
nor UO_1434 (O_1434,N_17226,N_16289);
or UO_1435 (O_1435,N_15089,N_16645);
nor UO_1436 (O_1436,N_17485,N_15062);
nand UO_1437 (O_1437,N_16740,N_19146);
xnor UO_1438 (O_1438,N_15859,N_19589);
xnor UO_1439 (O_1439,N_19303,N_15156);
xnor UO_1440 (O_1440,N_18230,N_19302);
nand UO_1441 (O_1441,N_17869,N_19573);
or UO_1442 (O_1442,N_17186,N_19588);
xor UO_1443 (O_1443,N_16354,N_19996);
or UO_1444 (O_1444,N_19525,N_16937);
and UO_1445 (O_1445,N_16026,N_17237);
xor UO_1446 (O_1446,N_18322,N_16604);
and UO_1447 (O_1447,N_16328,N_19846);
and UO_1448 (O_1448,N_17745,N_19473);
nor UO_1449 (O_1449,N_16113,N_15672);
or UO_1450 (O_1450,N_18463,N_18638);
or UO_1451 (O_1451,N_16348,N_16428);
or UO_1452 (O_1452,N_16173,N_17491);
and UO_1453 (O_1453,N_17112,N_19898);
nor UO_1454 (O_1454,N_16770,N_16540);
and UO_1455 (O_1455,N_19172,N_19877);
or UO_1456 (O_1456,N_18571,N_16020);
and UO_1457 (O_1457,N_16126,N_15616);
and UO_1458 (O_1458,N_15093,N_18038);
nand UO_1459 (O_1459,N_15211,N_18498);
or UO_1460 (O_1460,N_15313,N_18798);
and UO_1461 (O_1461,N_18325,N_16029);
or UO_1462 (O_1462,N_18820,N_18705);
xor UO_1463 (O_1463,N_19918,N_15967);
and UO_1464 (O_1464,N_19792,N_18581);
nand UO_1465 (O_1465,N_18164,N_17310);
xor UO_1466 (O_1466,N_19262,N_16320);
or UO_1467 (O_1467,N_16252,N_19233);
xor UO_1468 (O_1468,N_17711,N_19433);
nand UO_1469 (O_1469,N_17547,N_15396);
or UO_1470 (O_1470,N_19377,N_15256);
or UO_1471 (O_1471,N_15176,N_18527);
nand UO_1472 (O_1472,N_15410,N_15640);
and UO_1473 (O_1473,N_19381,N_16146);
nand UO_1474 (O_1474,N_15349,N_15404);
nor UO_1475 (O_1475,N_17421,N_16876);
nor UO_1476 (O_1476,N_15407,N_17142);
and UO_1477 (O_1477,N_19565,N_16499);
nand UO_1478 (O_1478,N_16045,N_18796);
or UO_1479 (O_1479,N_15614,N_17403);
and UO_1480 (O_1480,N_15973,N_15116);
xor UO_1481 (O_1481,N_15822,N_16688);
or UO_1482 (O_1482,N_16296,N_18776);
nand UO_1483 (O_1483,N_16138,N_18578);
xor UO_1484 (O_1484,N_17164,N_18809);
nor UO_1485 (O_1485,N_15242,N_17282);
or UO_1486 (O_1486,N_18914,N_18059);
nand UO_1487 (O_1487,N_16475,N_17532);
nor UO_1488 (O_1488,N_15336,N_15626);
nor UO_1489 (O_1489,N_19973,N_15671);
and UO_1490 (O_1490,N_15958,N_19780);
or UO_1491 (O_1491,N_19341,N_19411);
or UO_1492 (O_1492,N_16558,N_16443);
or UO_1493 (O_1493,N_19068,N_16436);
nand UO_1494 (O_1494,N_18228,N_18457);
or UO_1495 (O_1495,N_15600,N_17852);
and UO_1496 (O_1496,N_15516,N_17279);
nor UO_1497 (O_1497,N_15152,N_19891);
nand UO_1498 (O_1498,N_19686,N_19604);
or UO_1499 (O_1499,N_15858,N_17331);
and UO_1500 (O_1500,N_15654,N_19648);
or UO_1501 (O_1501,N_17168,N_15384);
xor UO_1502 (O_1502,N_16263,N_15883);
xnor UO_1503 (O_1503,N_19169,N_16257);
xnor UO_1504 (O_1504,N_18685,N_17069);
xnor UO_1505 (O_1505,N_16082,N_17895);
or UO_1506 (O_1506,N_16297,N_18406);
nand UO_1507 (O_1507,N_15531,N_19391);
and UO_1508 (O_1508,N_16683,N_18121);
xnor UO_1509 (O_1509,N_19186,N_19971);
and UO_1510 (O_1510,N_18352,N_18808);
xor UO_1511 (O_1511,N_16833,N_18093);
xor UO_1512 (O_1512,N_16721,N_18619);
xor UO_1513 (O_1513,N_18443,N_15434);
nor UO_1514 (O_1514,N_15180,N_19728);
and UO_1515 (O_1515,N_17807,N_17741);
and UO_1516 (O_1516,N_18388,N_18697);
nand UO_1517 (O_1517,N_15151,N_18124);
nand UO_1518 (O_1518,N_16593,N_19684);
and UO_1519 (O_1519,N_18778,N_18290);
or UO_1520 (O_1520,N_16831,N_18144);
or UO_1521 (O_1521,N_19291,N_19928);
nand UO_1522 (O_1522,N_17903,N_16147);
xor UO_1523 (O_1523,N_17067,N_18982);
xor UO_1524 (O_1524,N_17845,N_15238);
and UO_1525 (O_1525,N_19921,N_16325);
and UO_1526 (O_1526,N_18022,N_18656);
xnor UO_1527 (O_1527,N_18953,N_16742);
and UO_1528 (O_1528,N_17296,N_15677);
xor UO_1529 (O_1529,N_17700,N_17683);
nand UO_1530 (O_1530,N_17906,N_17257);
nand UO_1531 (O_1531,N_19352,N_15385);
xnor UO_1532 (O_1532,N_16663,N_19250);
nor UO_1533 (O_1533,N_18340,N_18196);
or UO_1534 (O_1534,N_17021,N_16329);
xor UO_1535 (O_1535,N_15305,N_15818);
and UO_1536 (O_1536,N_18692,N_18375);
nor UO_1537 (O_1537,N_19637,N_16180);
or UO_1538 (O_1538,N_19263,N_19122);
nor UO_1539 (O_1539,N_18935,N_17913);
xnor UO_1540 (O_1540,N_16397,N_15539);
nand UO_1541 (O_1541,N_18850,N_15778);
xnor UO_1542 (O_1542,N_17651,N_19897);
xor UO_1543 (O_1543,N_15249,N_15293);
or UO_1544 (O_1544,N_16954,N_18394);
nand UO_1545 (O_1545,N_15072,N_17374);
and UO_1546 (O_1546,N_16491,N_16655);
or UO_1547 (O_1547,N_16827,N_19544);
nand UO_1548 (O_1548,N_18785,N_19642);
xor UO_1549 (O_1549,N_16641,N_16885);
and UO_1550 (O_1550,N_15831,N_15383);
nand UO_1551 (O_1551,N_16649,N_18951);
nand UO_1552 (O_1552,N_19900,N_19799);
xnor UO_1553 (O_1553,N_17437,N_19699);
or UO_1554 (O_1554,N_16090,N_17932);
and UO_1555 (O_1555,N_15662,N_18384);
xnor UO_1556 (O_1556,N_18644,N_15746);
nand UO_1557 (O_1557,N_19198,N_18471);
nor UO_1558 (O_1558,N_19188,N_18643);
nand UO_1559 (O_1559,N_15068,N_16620);
or UO_1560 (O_1560,N_19339,N_19387);
xnor UO_1561 (O_1561,N_17844,N_19375);
and UO_1562 (O_1562,N_16095,N_15566);
and UO_1563 (O_1563,N_17463,N_18816);
nor UO_1564 (O_1564,N_16130,N_19160);
nor UO_1565 (O_1565,N_17360,N_18437);
nor UO_1566 (O_1566,N_17161,N_15756);
and UO_1567 (O_1567,N_19481,N_19758);
or UO_1568 (O_1568,N_15773,N_18142);
or UO_1569 (O_1569,N_17582,N_19042);
xnor UO_1570 (O_1570,N_15075,N_17355);
and UO_1571 (O_1571,N_18528,N_15706);
or UO_1572 (O_1572,N_15748,N_19358);
nand UO_1573 (O_1573,N_19974,N_16239);
or UO_1574 (O_1574,N_17715,N_15854);
xnor UO_1575 (O_1575,N_17584,N_16902);
or UO_1576 (O_1576,N_18063,N_17614);
nand UO_1577 (O_1577,N_16241,N_16855);
and UO_1578 (O_1578,N_15000,N_19540);
nor UO_1579 (O_1579,N_17220,N_15083);
and UO_1580 (O_1580,N_15682,N_15428);
nor UO_1581 (O_1581,N_15797,N_18163);
and UO_1582 (O_1582,N_16500,N_18441);
nor UO_1583 (O_1583,N_17006,N_16060);
nor UO_1584 (O_1584,N_16506,N_16783);
xor UO_1585 (O_1585,N_16968,N_15460);
nor UO_1586 (O_1586,N_15368,N_18519);
xor UO_1587 (O_1587,N_18069,N_19211);
nand UO_1588 (O_1588,N_18411,N_15477);
xor UO_1589 (O_1589,N_15303,N_15865);
and UO_1590 (O_1590,N_17330,N_17328);
nand UO_1591 (O_1591,N_18760,N_17500);
xnor UO_1592 (O_1592,N_16395,N_17889);
nor UO_1593 (O_1593,N_15939,N_17372);
nand UO_1594 (O_1594,N_19254,N_16085);
and UO_1595 (O_1595,N_18424,N_16975);
nor UO_1596 (O_1596,N_17666,N_15669);
or UO_1597 (O_1597,N_19335,N_15506);
nor UO_1598 (O_1598,N_17016,N_18969);
and UO_1599 (O_1599,N_19502,N_18157);
and UO_1600 (O_1600,N_19857,N_18956);
and UO_1601 (O_1601,N_17988,N_18888);
nand UO_1602 (O_1602,N_16350,N_19887);
or UO_1603 (O_1603,N_17597,N_16931);
nor UO_1604 (O_1604,N_19067,N_16426);
nor UO_1605 (O_1605,N_15998,N_17357);
or UO_1606 (O_1606,N_16194,N_19807);
and UO_1607 (O_1607,N_15485,N_16822);
or UO_1608 (O_1608,N_17694,N_18126);
nor UO_1609 (O_1609,N_19662,N_18596);
or UO_1610 (O_1610,N_19706,N_19566);
and UO_1611 (O_1611,N_19609,N_16985);
and UO_1612 (O_1612,N_19371,N_16145);
and UO_1613 (O_1613,N_18269,N_18041);
nand UO_1614 (O_1614,N_15079,N_15096);
xnor UO_1615 (O_1615,N_19868,N_17022);
nand UO_1616 (O_1616,N_17737,N_19808);
or UO_1617 (O_1617,N_17637,N_19886);
xnor UO_1618 (O_1618,N_16102,N_16809);
and UO_1619 (O_1619,N_18532,N_17936);
nor UO_1620 (O_1620,N_15310,N_15754);
xor UO_1621 (O_1621,N_17276,N_18188);
xor UO_1622 (O_1622,N_16501,N_18023);
xor UO_1623 (O_1623,N_17303,N_19711);
xor UO_1624 (O_1624,N_18895,N_17604);
xor UO_1625 (O_1625,N_19048,N_19849);
xnor UO_1626 (O_1626,N_16551,N_18555);
and UO_1627 (O_1627,N_15067,N_16971);
or UO_1628 (O_1628,N_16830,N_15980);
nand UO_1629 (O_1629,N_15245,N_19062);
xor UO_1630 (O_1630,N_15986,N_16100);
or UO_1631 (O_1631,N_17055,N_17219);
and UO_1632 (O_1632,N_17052,N_15388);
xor UO_1633 (O_1633,N_18757,N_18731);
and UO_1634 (O_1634,N_17242,N_15381);
or UO_1635 (O_1635,N_17262,N_18858);
xor UO_1636 (O_1636,N_17442,N_16091);
xor UO_1637 (O_1637,N_15128,N_19093);
xor UO_1638 (O_1638,N_19168,N_18102);
nand UO_1639 (O_1639,N_17474,N_17838);
xor UO_1640 (O_1640,N_18689,N_18342);
and UO_1641 (O_1641,N_18775,N_15589);
nand UO_1642 (O_1642,N_17915,N_19594);
or UO_1643 (O_1643,N_17619,N_17958);
nor UO_1644 (O_1644,N_18199,N_19412);
nor UO_1645 (O_1645,N_15196,N_16062);
xor UO_1646 (O_1646,N_16166,N_16260);
nor UO_1647 (O_1647,N_16684,N_19383);
xnor UO_1648 (O_1648,N_17853,N_19142);
or UO_1649 (O_1649,N_17948,N_15010);
xor UO_1650 (O_1650,N_15230,N_17377);
nand UO_1651 (O_1651,N_19469,N_16217);
nand UO_1652 (O_1652,N_16444,N_17873);
nand UO_1653 (O_1653,N_17352,N_18975);
xnor UO_1654 (O_1654,N_18211,N_19685);
xor UO_1655 (O_1655,N_16034,N_19938);
or UO_1656 (O_1656,N_15977,N_17718);
xnor UO_1657 (O_1657,N_19522,N_17177);
and UO_1658 (O_1658,N_16621,N_15852);
and UO_1659 (O_1659,N_15972,N_19989);
and UO_1660 (O_1660,N_16897,N_16490);
or UO_1661 (O_1661,N_16872,N_16536);
nor UO_1662 (O_1662,N_19056,N_18677);
nand UO_1663 (O_1663,N_18539,N_16203);
nor UO_1664 (O_1664,N_15764,N_16268);
nand UO_1665 (O_1665,N_15801,N_17189);
nor UO_1666 (O_1666,N_17908,N_17084);
nand UO_1667 (O_1667,N_16635,N_15203);
and UO_1668 (O_1668,N_15441,N_16586);
nor UO_1669 (O_1669,N_18209,N_17771);
nor UO_1670 (O_1670,N_16134,N_19949);
nand UO_1671 (O_1671,N_19788,N_16233);
or UO_1672 (O_1672,N_18564,N_19389);
nand UO_1673 (O_1673,N_16277,N_15453);
and UO_1674 (O_1674,N_18236,N_16430);
nand UO_1675 (O_1675,N_16061,N_16537);
and UO_1676 (O_1676,N_16944,N_16468);
and UO_1677 (O_1677,N_16602,N_17155);
nor UO_1678 (O_1678,N_18461,N_16093);
nor UO_1679 (O_1679,N_19850,N_18777);
nand UO_1680 (O_1680,N_15140,N_18936);
and UO_1681 (O_1681,N_15162,N_17359);
nor UO_1682 (O_1682,N_16879,N_16367);
nor UO_1683 (O_1683,N_18159,N_17849);
nor UO_1684 (O_1684,N_18622,N_15194);
nand UO_1685 (O_1685,N_18373,N_15455);
nor UO_1686 (O_1686,N_15411,N_16181);
nor UO_1687 (O_1687,N_17754,N_18651);
and UO_1688 (O_1688,N_16186,N_19872);
xnor UO_1689 (O_1689,N_19281,N_17800);
xor UO_1690 (O_1690,N_18916,N_15246);
nor UO_1691 (O_1691,N_17183,N_19943);
and UO_1692 (O_1692,N_17455,N_15639);
or UO_1693 (O_1693,N_18004,N_19513);
and UO_1694 (O_1694,N_15565,N_18743);
nor UO_1695 (O_1695,N_19134,N_15955);
xor UO_1696 (O_1696,N_16959,N_16502);
nor UO_1697 (O_1697,N_16109,N_17093);
nand UO_1698 (O_1698,N_17173,N_17602);
and UO_1699 (O_1699,N_17832,N_17989);
and UO_1700 (O_1700,N_16653,N_18108);
nand UO_1701 (O_1701,N_18535,N_18400);
and UO_1702 (O_1702,N_18913,N_19781);
nor UO_1703 (O_1703,N_17225,N_15346);
nor UO_1704 (O_1704,N_17464,N_17926);
or UO_1705 (O_1705,N_16193,N_17393);
nor UO_1706 (O_1706,N_16716,N_17590);
and UO_1707 (O_1707,N_17031,N_15551);
nor UO_1708 (O_1708,N_15833,N_15970);
nand UO_1709 (O_1709,N_17149,N_15647);
or UO_1710 (O_1710,N_19806,N_19315);
nor UO_1711 (O_1711,N_18781,N_15908);
xnor UO_1712 (O_1712,N_19428,N_17466);
xnor UO_1713 (O_1713,N_17841,N_16171);
and UO_1714 (O_1714,N_18505,N_19401);
nor UO_1715 (O_1715,N_18160,N_18931);
and UO_1716 (O_1716,N_17047,N_19414);
xnor UO_1717 (O_1717,N_19058,N_19403);
xor UO_1718 (O_1718,N_19756,N_15853);
or UO_1719 (O_1719,N_17589,N_16575);
nand UO_1720 (O_1720,N_15587,N_16375);
and UO_1721 (O_1721,N_19083,N_18272);
nand UO_1722 (O_1722,N_18702,N_19124);
and UO_1723 (O_1723,N_19307,N_16891);
xor UO_1724 (O_1724,N_16787,N_19000);
nand UO_1725 (O_1725,N_19754,N_16615);
nor UO_1726 (O_1726,N_15509,N_15673);
nor UO_1727 (O_1727,N_15364,N_19202);
xnor UO_1728 (O_1728,N_17777,N_18674);
or UO_1729 (O_1729,N_18725,N_15039);
or UO_1730 (O_1730,N_19673,N_17135);
and UO_1731 (O_1731,N_18668,N_15825);
or UO_1732 (O_1732,N_15767,N_16888);
nor UO_1733 (O_1733,N_15607,N_18649);
or UO_1734 (O_1734,N_17105,N_17530);
xnor UO_1735 (O_1735,N_15676,N_15744);
nor UO_1736 (O_1736,N_15321,N_15653);
xnor UO_1737 (O_1737,N_18572,N_18428);
nand UO_1738 (O_1738,N_18092,N_18989);
or UO_1739 (O_1739,N_15226,N_18280);
or UO_1740 (O_1740,N_17432,N_16587);
xor UO_1741 (O_1741,N_19763,N_17023);
xnor UO_1742 (O_1742,N_19229,N_15723);
xor UO_1743 (O_1743,N_17871,N_19909);
and UO_1744 (O_1744,N_17329,N_18754);
nor UO_1745 (O_1745,N_15886,N_16585);
nand UO_1746 (O_1746,N_17204,N_18323);
xnor UO_1747 (O_1747,N_18299,N_18929);
nand UO_1748 (O_1748,N_18031,N_19461);
and UO_1749 (O_1749,N_15919,N_19532);
or UO_1750 (O_1750,N_15702,N_16389);
nor UO_1751 (O_1751,N_17494,N_15995);
nor UO_1752 (O_1752,N_17208,N_16917);
xnor UO_1753 (O_1753,N_17280,N_19427);
nor UO_1754 (O_1754,N_18208,N_17468);
nor UO_1755 (O_1755,N_17920,N_15130);
nor UO_1756 (O_1756,N_16002,N_18390);
nor UO_1757 (O_1757,N_16753,N_18077);
nor UO_1758 (O_1758,N_18902,N_17850);
and UO_1759 (O_1759,N_17576,N_19811);
nor UO_1760 (O_1760,N_17043,N_17519);
nor UO_1761 (O_1761,N_16170,N_18358);
or UO_1762 (O_1762,N_16522,N_19148);
nand UO_1763 (O_1763,N_19731,N_15666);
nor UO_1764 (O_1764,N_19752,N_19447);
or UO_1765 (O_1765,N_15960,N_15834);
nand UO_1766 (O_1766,N_15217,N_15182);
and UO_1767 (O_1767,N_15018,N_18700);
xor UO_1768 (O_1768,N_15860,N_18713);
nand UO_1769 (O_1769,N_16459,N_16472);
and UO_1770 (O_1770,N_19392,N_18112);
and UO_1771 (O_1771,N_16728,N_17243);
and UO_1772 (O_1772,N_16097,N_17110);
or UO_1773 (O_1773,N_17467,N_18320);
xor UO_1774 (O_1774,N_18171,N_15510);
and UO_1775 (O_1775,N_15279,N_16322);
nor UO_1776 (O_1776,N_16235,N_17042);
nand UO_1777 (O_1777,N_15679,N_18205);
xor UO_1778 (O_1778,N_19105,N_17013);
or UO_1779 (O_1779,N_16390,N_15789);
nor UO_1780 (O_1780,N_19601,N_18430);
nor UO_1781 (O_1781,N_15275,N_15577);
and UO_1782 (O_1782,N_17070,N_18145);
nor UO_1783 (O_1783,N_15815,N_18991);
xnor UO_1784 (O_1784,N_19787,N_16589);
or UO_1785 (O_1785,N_17649,N_17564);
and UO_1786 (O_1786,N_17985,N_18551);
and UO_1787 (O_1787,N_16966,N_16310);
xnor UO_1788 (O_1788,N_18028,N_19542);
and UO_1789 (O_1789,N_17716,N_15435);
or UO_1790 (O_1790,N_15750,N_19554);
or UO_1791 (O_1791,N_19745,N_18467);
nor UO_1792 (O_1792,N_16315,N_18860);
nor UO_1793 (O_1793,N_15386,N_19679);
or UO_1794 (O_1794,N_16371,N_15943);
nor UO_1795 (O_1795,N_17621,N_19257);
nor UO_1796 (O_1796,N_16081,N_18512);
xnor UO_1797 (O_1797,N_19063,N_18560);
and UO_1798 (O_1798,N_16865,N_17918);
nand UO_1799 (O_1799,N_17924,N_18281);
xor UO_1800 (O_1800,N_19766,N_16785);
nand UO_1801 (O_1801,N_15821,N_15057);
nand UO_1802 (O_1802,N_17728,N_19209);
and UO_1803 (O_1803,N_19832,N_19640);
nor UO_1804 (O_1804,N_16553,N_17417);
or UO_1805 (O_1805,N_17267,N_18791);
or UO_1806 (O_1806,N_18110,N_15438);
or UO_1807 (O_1807,N_15536,N_18368);
nor UO_1808 (O_1808,N_18728,N_17428);
nor UO_1809 (O_1809,N_18067,N_17433);
or UO_1810 (O_1810,N_19904,N_16246);
and UO_1811 (O_1811,N_15218,N_17834);
nand UO_1812 (O_1812,N_19729,N_15104);
nor UO_1813 (O_1813,N_18040,N_16483);
nand UO_1814 (O_1814,N_18255,N_17424);
xor UO_1815 (O_1815,N_18224,N_19969);
nor UO_1816 (O_1816,N_19225,N_16278);
and UO_1817 (O_1817,N_16651,N_15843);
nand UO_1818 (O_1818,N_19380,N_15020);
xor UO_1819 (O_1819,N_16949,N_16916);
nor UO_1820 (O_1820,N_19539,N_17456);
xnor UO_1821 (O_1821,N_16980,N_16111);
xnor UO_1822 (O_1822,N_18399,N_15472);
nor UO_1823 (O_1823,N_15989,N_15475);
or UO_1824 (O_1824,N_17732,N_19095);
nand UO_1825 (O_1825,N_17566,N_18576);
xnor UO_1826 (O_1826,N_16687,N_17738);
nand UO_1827 (O_1827,N_15774,N_15745);
nor UO_1828 (O_1828,N_18499,N_19246);
or UO_1829 (O_1829,N_17202,N_19838);
nand UO_1830 (O_1830,N_15687,N_15459);
or UO_1831 (O_1831,N_19636,N_16622);
nand UO_1832 (O_1832,N_17075,N_17712);
nor UO_1833 (O_1833,N_15447,N_15911);
nor UO_1834 (O_1834,N_17756,N_19113);
nor UO_1835 (O_1835,N_19293,N_15052);
nand UO_1836 (O_1836,N_17104,N_19836);
xor UO_1837 (O_1837,N_17342,N_19824);
xnor UO_1838 (O_1838,N_16667,N_17720);
and UO_1839 (O_1839,N_19550,N_19830);
nor UO_1840 (O_1840,N_18372,N_17511);
nand UO_1841 (O_1841,N_19342,N_15183);
nor UO_1842 (O_1842,N_17822,N_16576);
xor UO_1843 (O_1843,N_16202,N_19592);
nor UO_1844 (O_1844,N_15027,N_17498);
xor UO_1845 (O_1845,N_16851,N_17588);
nor UO_1846 (O_1846,N_17986,N_17826);
nand UO_1847 (O_1847,N_19855,N_16804);
or UO_1848 (O_1848,N_16691,N_19700);
and UO_1849 (O_1849,N_19579,N_19607);
nand UO_1850 (O_1850,N_18439,N_16122);
nor UO_1851 (O_1851,N_18367,N_15326);
or UO_1852 (O_1852,N_15325,N_15841);
and UO_1853 (O_1853,N_18003,N_19123);
nand UO_1854 (O_1854,N_19394,N_18730);
or UO_1855 (O_1855,N_16478,N_19791);
and UO_1856 (O_1856,N_17087,N_17801);
xor UO_1857 (O_1857,N_18496,N_18296);
and UO_1858 (O_1858,N_19937,N_19235);
or UO_1859 (O_1859,N_17827,N_16619);
nand UO_1860 (O_1860,N_16609,N_16292);
xnor UO_1861 (O_1861,N_18772,N_15559);
xnor UO_1862 (O_1862,N_16662,N_15103);
nand UO_1863 (O_1863,N_17228,N_17236);
or UO_1864 (O_1864,N_15912,N_18326);
nand UO_1865 (O_1865,N_19494,N_15543);
nor UO_1866 (O_1866,N_16112,N_16637);
and UO_1867 (O_1867,N_19998,N_17132);
and UO_1868 (O_1868,N_16461,N_16923);
or UO_1869 (O_1869,N_16788,N_15556);
xor UO_1870 (O_1870,N_19361,N_15824);
or UO_1871 (O_1871,N_18349,N_19405);
or UO_1872 (O_1872,N_16832,N_17119);
and UO_1873 (O_1873,N_15188,N_19680);
xnor UO_1874 (O_1874,N_17221,N_16521);
nand UO_1875 (O_1875,N_19053,N_17609);
xor UO_1876 (O_1876,N_18318,N_17073);
or UO_1877 (O_1877,N_17082,N_19746);
nor UO_1878 (O_1878,N_19587,N_19922);
or UO_1879 (O_1879,N_16759,N_17556);
xnor UO_1880 (O_1880,N_16327,N_19641);
and UO_1881 (O_1881,N_18204,N_19861);
or UO_1882 (O_1882,N_18699,N_16969);
xnor UO_1883 (O_1883,N_15193,N_16370);
and UO_1884 (O_1884,N_16707,N_18986);
and UO_1885 (O_1885,N_16124,N_17645);
nand UO_1886 (O_1886,N_19097,N_19163);
nand UO_1887 (O_1887,N_18882,N_17389);
nand UO_1888 (O_1888,N_18162,N_18837);
xnor UO_1889 (O_1889,N_19376,N_16796);
nor UO_1890 (O_1890,N_15141,N_18976);
xnor UO_1891 (O_1891,N_17014,N_16907);
nor UO_1892 (O_1892,N_19772,N_19001);
nand UO_1893 (O_1893,N_18039,N_15456);
or UO_1894 (O_1894,N_16863,N_19717);
nor UO_1895 (O_1895,N_18817,N_17730);
xnor UO_1896 (O_1896,N_15131,N_15515);
or UO_1897 (O_1897,N_19455,N_18517);
or UO_1898 (O_1898,N_18570,N_19556);
or UO_1899 (O_1899,N_17409,N_18972);
nand UO_1900 (O_1900,N_18101,N_19273);
or UO_1901 (O_1901,N_15985,N_19019);
xnor UO_1902 (O_1902,N_17816,N_19769);
nor UO_1903 (O_1903,N_17033,N_16473);
xor UO_1904 (O_1904,N_15550,N_18905);
and UO_1905 (O_1905,N_17397,N_19230);
and UO_1906 (O_1906,N_15101,N_15060);
and UO_1907 (O_1907,N_18116,N_17270);
xnor UO_1908 (O_1908,N_15255,N_16238);
xor UO_1909 (O_1909,N_19629,N_19523);
xnor UO_1910 (O_1910,N_19831,N_17856);
xnor UO_1911 (O_1911,N_19464,N_16385);
and UO_1912 (O_1912,N_19321,N_16866);
xor UO_1913 (O_1913,N_17923,N_16799);
xnor UO_1914 (O_1914,N_18354,N_19644);
nor UO_1915 (O_1915,N_18557,N_16167);
and UO_1916 (O_1916,N_19687,N_16850);
nor UO_1917 (O_1917,N_18327,N_16009);
xor UO_1918 (O_1918,N_18233,N_17612);
xnor UO_1919 (O_1919,N_15694,N_19795);
nand UO_1920 (O_1920,N_15921,N_18684);
and UO_1921 (O_1921,N_18946,N_16664);
xnor UO_1922 (O_1922,N_15897,N_16092);
nor UO_1923 (O_1923,N_15458,N_19022);
xor UO_1924 (O_1924,N_16245,N_17453);
or UO_1925 (O_1925,N_16983,N_19976);
xor UO_1926 (O_1926,N_18218,N_18573);
and UO_1927 (O_1927,N_17187,N_19596);
and UO_1928 (O_1928,N_17786,N_18646);
and UO_1929 (O_1929,N_16190,N_19903);
nor UO_1930 (O_1930,N_18125,N_17053);
or UO_1931 (O_1931,N_15059,N_15186);
xnor UO_1932 (O_1932,N_16930,N_19003);
nor UO_1933 (O_1933,N_16706,N_15807);
or UO_1934 (O_1934,N_17507,N_19115);
and UO_1935 (O_1935,N_17484,N_15898);
nand UO_1936 (O_1936,N_18509,N_19571);
or UO_1937 (O_1937,N_18427,N_15292);
xnor UO_1938 (O_1938,N_15181,N_17163);
or UO_1939 (O_1939,N_17117,N_16215);
nand UO_1940 (O_1940,N_15291,N_15946);
and UO_1941 (O_1941,N_19350,N_15403);
or UO_1942 (O_1942,N_19533,N_15055);
xnor UO_1943 (O_1943,N_16341,N_16894);
xnor UO_1944 (O_1944,N_18899,N_17925);
nor UO_1945 (O_1945,N_19075,N_16379);
nor UO_1946 (O_1946,N_15011,N_18846);
xnor UO_1947 (O_1947,N_15711,N_18436);
nor UO_1948 (O_1948,N_15080,N_19620);
or UO_1949 (O_1949,N_17866,N_15999);
xnor UO_1950 (O_1950,N_17644,N_18363);
xnor UO_1951 (O_1951,N_15206,N_18177);
xnor UO_1952 (O_1952,N_16957,N_18225);
or UO_1953 (O_1953,N_15848,N_17240);
and UO_1954 (O_1954,N_18614,N_19336);
or UO_1955 (O_1955,N_16066,N_19834);
and UO_1956 (O_1956,N_15234,N_15007);
xnor UO_1957 (O_1957,N_18771,N_15423);
or UO_1958 (O_1958,N_17441,N_19325);
and UO_1959 (O_1959,N_18629,N_17825);
and UO_1960 (O_1960,N_18189,N_15517);
nor UO_1961 (O_1961,N_16249,N_18665);
nor UO_1962 (O_1962,N_16221,N_17490);
and UO_1963 (O_1963,N_18948,N_19292);
and UO_1964 (O_1964,N_18682,N_15601);
or UO_1965 (O_1965,N_16175,N_19512);
or UO_1966 (O_1966,N_17040,N_17007);
xor UO_1967 (O_1967,N_17533,N_16993);
and UO_1968 (O_1968,N_19980,N_17770);
nor UO_1969 (O_1969,N_15528,N_15094);
nor UO_1970 (O_1970,N_16396,N_16994);
nor UO_1971 (O_1971,N_16555,N_18068);
or UO_1972 (O_1972,N_18444,N_18012);
nor UO_1973 (O_1973,N_16132,N_17999);
and UO_1974 (O_1974,N_18308,N_18410);
nand UO_1975 (O_1975,N_16769,N_16365);
and UO_1976 (O_1976,N_18901,N_15817);
nor UO_1977 (O_1977,N_19923,N_15343);
and UO_1978 (O_1978,N_16735,N_16940);
and UO_1979 (O_1979,N_18995,N_19908);
nor UO_1980 (O_1980,N_17388,N_19863);
nor UO_1981 (O_1981,N_17731,N_16105);
or UO_1982 (O_1982,N_19070,N_17351);
nand UO_1983 (O_1983,N_17253,N_16384);
and UO_1984 (O_1984,N_19987,N_15631);
nor UO_1985 (O_1985,N_19718,N_19333);
nor UO_1986 (O_1986,N_18179,N_19135);
or UO_1987 (O_1987,N_16582,N_15237);
and UO_1988 (O_1988,N_17605,N_19771);
nor UO_1989 (O_1989,N_17806,N_16659);
xor UO_1990 (O_1990,N_15071,N_19034);
and UO_1991 (O_1991,N_19541,N_19415);
nand UO_1992 (O_1992,N_18868,N_17882);
nor UO_1993 (O_1993,N_15224,N_15198);
or UO_1994 (O_1994,N_17596,N_16952);
or UO_1995 (O_1995,N_16724,N_18792);
xnor UO_1996 (O_1996,N_19311,N_16806);
nor UO_1997 (O_1997,N_16455,N_15440);
nand UO_1998 (O_1998,N_15512,N_16140);
nand UO_1999 (O_1999,N_19770,N_18032);
nor UO_2000 (O_2000,N_16689,N_19038);
and UO_2001 (O_2001,N_15307,N_17148);
and UO_2002 (O_2002,N_15120,N_18659);
nor UO_2003 (O_2003,N_16316,N_18766);
nand UO_2004 (O_2004,N_17851,N_17987);
xnor UO_2005 (O_2005,N_17420,N_15298);
nor UO_2006 (O_2006,N_17933,N_16920);
nand UO_2007 (O_2007,N_16617,N_15363);
nor UO_2008 (O_2008,N_19630,N_16745);
or UO_2009 (O_2009,N_15590,N_17361);
nand UO_2010 (O_2010,N_18794,N_15742);
and UO_2011 (O_2011,N_19876,N_18779);
or UO_2012 (O_2012,N_16131,N_16588);
nand UO_2013 (O_2013,N_15761,N_18007);
and UO_2014 (O_2014,N_18315,N_15593);
nand UO_2015 (O_2015,N_17292,N_18515);
xor UO_2016 (O_2016,N_19860,N_16758);
or UO_2017 (O_2017,N_17151,N_19179);
nor UO_2018 (O_2018,N_16714,N_16159);
or UO_2019 (O_2019,N_16099,N_16873);
and UO_2020 (O_2020,N_17642,N_19526);
nand UO_2021 (O_2021,N_15344,N_18524);
or UO_2022 (O_2022,N_19253,N_15827);
nor UO_2023 (O_2023,N_15416,N_19954);
nor UO_2024 (O_2024,N_17972,N_17865);
and UO_2025 (O_2025,N_16882,N_16864);
and UO_2026 (O_2026,N_15729,N_19312);
nor UO_2027 (O_2027,N_19176,N_17580);
nor UO_2028 (O_2028,N_19999,N_16812);
or UO_2029 (O_2029,N_17440,N_17966);
and UO_2030 (O_2030,N_18206,N_15525);
nor UO_2031 (O_2031,N_18664,N_16877);
or UO_2032 (O_2032,N_16911,N_15530);
and UO_2033 (O_2033,N_19852,N_16338);
xnor UO_2034 (O_2034,N_19110,N_15644);
xnor UO_2035 (O_2035,N_18490,N_19033);
xor UO_2036 (O_2036,N_16374,N_19203);
or UO_2037 (O_2037,N_18897,N_18671);
nand UO_2038 (O_2038,N_16672,N_19798);
xor UO_2039 (O_2039,N_19660,N_18304);
nor UO_2040 (O_2040,N_17953,N_15271);
xor UO_2041 (O_2041,N_18348,N_15185);
nor UO_2042 (O_2042,N_15862,N_17365);
xnor UO_2043 (O_2043,N_19965,N_19507);
nand UO_2044 (O_2044,N_17318,N_15800);
xor UO_2045 (O_2045,N_16997,N_18429);
and UO_2046 (O_2046,N_16824,N_18291);
nor UO_2047 (O_2047,N_15892,N_18900);
xnor UO_2048 (O_2048,N_19576,N_15480);
or UO_2049 (O_2049,N_19521,N_17147);
nand UO_2050 (O_2050,N_17922,N_19417);
and UO_2051 (O_2051,N_17962,N_17729);
and UO_2052 (O_2052,N_17159,N_16956);
xor UO_2053 (O_2053,N_18745,N_18864);
and UO_2054 (O_2054,N_16197,N_16191);
nand UO_2055 (O_2055,N_16272,N_17733);
nor UO_2056 (O_2056,N_18857,N_16698);
nor UO_2057 (O_2057,N_19345,N_18098);
and UO_2058 (O_2058,N_15776,N_17405);
xnor UO_2059 (O_2059,N_17416,N_15704);
or UO_2060 (O_2060,N_19300,N_19236);
and UO_2061 (O_2061,N_15777,N_16299);
and UO_2062 (O_2062,N_17570,N_15241);
nor UO_2063 (O_2063,N_17870,N_15726);
or UO_2064 (O_2064,N_15873,N_16135);
xor UO_2065 (O_2065,N_17157,N_15878);
nor UO_2066 (O_2066,N_16835,N_17004);
or UO_2067 (O_2067,N_18922,N_18072);
nand UO_2068 (O_2068,N_16819,N_18650);
or UO_2069 (O_2069,N_15592,N_15263);
nand UO_2070 (O_2070,N_18998,N_15953);
or UO_2071 (O_2071,N_17969,N_19669);
nor UO_2072 (O_2072,N_18195,N_19584);
nand UO_2073 (O_2073,N_18053,N_16775);
xor UO_2074 (O_2074,N_18278,N_18880);
nand UO_2075 (O_2075,N_16442,N_18550);
and UO_2076 (O_2076,N_18939,N_18871);
nor UO_2077 (O_2077,N_16094,N_18097);
nand UO_2078 (O_2078,N_15929,N_16077);
and UO_2079 (O_2079,N_16528,N_19219);
xor UO_2080 (O_2080,N_19698,N_16878);
nand UO_2081 (O_2081,N_17269,N_17166);
or UO_2082 (O_2082,N_16607,N_17010);
nor UO_2083 (O_2083,N_19916,N_17218);
xor UO_2084 (O_2084,N_18447,N_18220);
and UO_2085 (O_2085,N_16712,N_15869);
or UO_2086 (O_2086,N_18744,N_17210);
nor UO_2087 (O_2087,N_15579,N_19994);
xnor UO_2088 (O_2088,N_19714,N_15287);
nor UO_2089 (O_2089,N_17011,N_19591);
nor UO_2090 (O_2090,N_19059,N_18927);
and UO_2091 (O_2091,N_17567,N_16256);
nor UO_2092 (O_2092,N_16709,N_19450);
nor UO_2093 (O_2093,N_19458,N_19006);
and UO_2094 (O_2094,N_15732,N_17201);
xor UO_2095 (O_2095,N_17341,N_18016);
and UO_2096 (O_2096,N_18392,N_16369);
nand UO_2097 (O_2097,N_16044,N_15533);
nor UO_2098 (O_2098,N_19157,N_17543);
nand UO_2099 (O_2099,N_18957,N_18307);
nor UO_2100 (O_2100,N_19132,N_16717);
nor UO_2101 (O_2101,N_18198,N_18139);
nor UO_2102 (O_2102,N_19985,N_18448);
nor UO_2103 (O_2103,N_19751,N_19112);
and UO_2104 (O_2104,N_17200,N_16425);
xor UO_2105 (O_2105,N_17654,N_18683);
nor UO_2106 (O_2106,N_18146,N_19929);
nand UO_2107 (O_2107,N_15968,N_17128);
and UO_2108 (O_2108,N_18849,N_19761);
and UO_2109 (O_2109,N_18376,N_19935);
xor UO_2110 (O_2110,N_18415,N_15710);
xnor UO_2111 (O_2111,N_18627,N_17601);
nand UO_2112 (O_2112,N_15545,N_16416);
xnor UO_2113 (O_2113,N_18466,N_15178);
or UO_2114 (O_2114,N_17347,N_15725);
and UO_2115 (O_2115,N_15845,N_15158);
and UO_2116 (O_2116,N_16495,N_15223);
or UO_2117 (O_2117,N_19497,N_18335);
and UO_2118 (O_2118,N_17044,N_18655);
xor UO_2119 (O_2119,N_17696,N_18353);
and UO_2120 (O_2120,N_18639,N_16761);
nor UO_2121 (O_2121,N_18186,N_16458);
xnor UO_2122 (O_2122,N_16842,N_17518);
and UO_2123 (O_2123,N_18197,N_16636);
and UO_2124 (O_2124,N_19159,N_16870);
nor UO_2125 (O_2125,N_16188,N_19199);
nand UO_2126 (O_2126,N_19305,N_19437);
nor UO_2127 (O_2127,N_17579,N_18222);
or UO_2128 (O_2128,N_18770,N_18219);
nor UO_2129 (O_2129,N_18997,N_18597);
nor UO_2130 (O_2130,N_16557,N_19008);
and UO_2131 (O_2131,N_16677,N_17961);
nor UO_2132 (O_2132,N_18287,N_17222);
and UO_2133 (O_2133,N_15212,N_16624);
and UO_2134 (O_2134,N_18633,N_15421);
nor UO_2135 (O_2135,N_19847,N_17618);
or UO_2136 (O_2136,N_18404,N_15035);
nand UO_2137 (O_2137,N_19946,N_17286);
nand UO_2138 (O_2138,N_17315,N_18893);
and UO_2139 (O_2139,N_16010,N_19866);
and UO_2140 (O_2140,N_16211,N_15916);
or UO_2141 (O_2141,N_17685,N_17191);
xnor UO_2142 (O_2142,N_18842,N_18180);
nor UO_2143 (O_2143,N_18062,N_15426);
nor UO_2144 (O_2144,N_18844,N_19239);
nor UO_2145 (O_2145,N_18709,N_15493);
or UO_2146 (O_2146,N_17881,N_18216);
xor UO_2147 (O_2147,N_16098,N_16984);
and UO_2148 (O_2148,N_17239,N_16494);
or UO_2149 (O_2149,N_16583,N_19190);
and UO_2150 (O_2150,N_17837,N_18965);
xor UO_2151 (O_2151,N_17976,N_16065);
or UO_2152 (O_2152,N_15113,N_19543);
xnor UO_2153 (O_2153,N_15652,N_18141);
nor UO_2154 (O_2154,N_15491,N_17583);
and UO_2155 (O_2155,N_19880,N_19794);
nor UO_2156 (O_2156,N_19867,N_18316);
xnor UO_2157 (O_2157,N_16614,N_16119);
or UO_2158 (O_2158,N_16658,N_16856);
nor UO_2159 (O_2159,N_18351,N_16030);
xnor UO_2160 (O_2160,N_17392,N_15751);
xnor UO_2161 (O_2161,N_19153,N_18332);
and UO_2162 (O_2162,N_18790,N_16563);
or UO_2163 (O_2163,N_17914,N_19668);
and UO_2164 (O_2164,N_15624,N_18256);
nand UO_2165 (O_2165,N_17172,N_19047);
xnor UO_2166 (O_2166,N_18350,N_16357);
or UO_2167 (O_2167,N_19471,N_16466);
xnor UO_2168 (O_2168,N_19446,N_18716);
nor UO_2169 (O_2169,N_16005,N_17572);
xnor UO_2170 (O_2170,N_16274,N_17097);
and UO_2171 (O_2171,N_16517,N_19012);
nor UO_2172 (O_2172,N_18676,N_15294);
and UO_2173 (O_2173,N_19248,N_16117);
xnor UO_2174 (O_2174,N_16825,N_18273);
or UO_2175 (O_2175,N_16232,N_16290);
and UO_2176 (O_2176,N_17152,N_17162);
and UO_2177 (O_2177,N_19449,N_19216);
xor UO_2178 (O_2178,N_18751,N_16564);
and UO_2179 (O_2179,N_18943,N_19530);
and UO_2180 (O_2180,N_19519,N_19613);
nor UO_2181 (O_2181,N_19191,N_15467);
and UO_2182 (O_2182,N_19505,N_15273);
nand UO_2183 (O_2183,N_15213,N_15714);
and UO_2184 (O_2184,N_15078,N_15871);
or UO_2185 (O_2185,N_16657,N_17971);
nand UO_2186 (O_2186,N_18240,N_17356);
and UO_2187 (O_2187,N_17370,N_15312);
or UO_2188 (O_2188,N_17763,N_15268);
xor UO_2189 (O_2189,N_18462,N_15895);
or UO_2190 (O_2190,N_15709,N_15928);
nand UO_2191 (O_2191,N_16018,N_15836);
and UO_2192 (O_2192,N_18250,N_18787);
nor UO_2193 (O_2193,N_19147,N_19906);
xor UO_2194 (O_2194,N_18453,N_15814);
or UO_2195 (O_2195,N_17008,N_18282);
xnor UO_2196 (O_2196,N_17620,N_16470);
xor UO_2197 (O_2197,N_19408,N_17661);
and UO_2198 (O_2198,N_17782,N_16630);
xnor UO_2199 (O_2199,N_18854,N_19940);
nor UO_2200 (O_2200,N_15232,N_18305);
xor UO_2201 (O_2201,N_18932,N_19818);
and UO_2202 (O_2202,N_15674,N_15427);
or UO_2203 (O_2203,N_19125,N_16580);
nand UO_2204 (O_2204,N_15394,N_17125);
or UO_2205 (O_2205,N_15885,N_15329);
xor UO_2206 (O_2206,N_18276,N_19343);
nor UO_2207 (O_2207,N_17215,N_17150);
xor UO_2208 (O_2208,N_19634,N_17065);
xnor UO_2209 (O_2209,N_18861,N_17314);
xnor UO_2210 (O_2210,N_19104,N_18310);
nor UO_2211 (O_2211,N_17890,N_19205);
or UO_2212 (O_2212,N_17353,N_18654);
and UO_2213 (O_2213,N_15906,N_16319);
nor UO_2214 (O_2214,N_19240,N_18248);
and UO_2215 (O_2215,N_17847,N_19045);
nand UO_2216 (O_2216,N_17002,N_18324);
or UO_2217 (O_2217,N_18440,N_17568);
xnor UO_2218 (O_2218,N_15341,N_18992);
nor UO_2219 (O_2219,N_19109,N_17169);
nor UO_2220 (O_2220,N_17681,N_19121);
nand UO_2221 (O_2221,N_17212,N_19527);
nor UO_2222 (O_2222,N_15413,N_16692);
nor UO_2223 (O_2223,N_19691,N_19174);
and UO_2224 (O_2224,N_18832,N_17488);
and UO_2225 (O_2225,N_15574,N_19136);
nor UO_2226 (O_2226,N_18607,N_16144);
xor UO_2227 (O_2227,N_19793,N_18647);
nand UO_2228 (O_2228,N_19915,N_18095);
xnor UO_2229 (O_2229,N_16153,N_19610);
nand UO_2230 (O_2230,N_19585,N_15077);
xor UO_2231 (O_2231,N_15981,N_19564);
nor UO_2232 (O_2232,N_16321,N_19753);
nand UO_2233 (O_2233,N_19295,N_18271);
and UO_2234 (O_2234,N_17336,N_15331);
nor UO_2235 (O_2235,N_17325,N_15555);
nor UO_2236 (O_2236,N_15070,N_15302);
or UO_2237 (O_2237,N_17297,N_18044);
nand UO_2238 (O_2238,N_18495,N_17460);
nor UO_2239 (O_2239,N_17048,N_19051);
or UO_2240 (O_2240,N_15987,N_15369);
nand UO_2241 (O_2241,N_18456,N_18207);
or UO_2242 (O_2242,N_16447,N_17283);
nand UO_2243 (O_2243,N_16892,N_17723);
nand UO_2244 (O_2244,N_17931,N_18295);
or UO_2245 (O_2245,N_16845,N_16890);
and UO_2246 (O_2246,N_18736,N_16453);
and UO_2247 (O_2247,N_17909,N_18782);
or UO_2248 (O_2248,N_18724,N_17244);
and UO_2249 (O_2249,N_17316,N_15126);
xor UO_2250 (O_2250,N_18359,N_16596);
or UO_2251 (O_2251,N_17113,N_15199);
and UO_2252 (O_2252,N_17108,N_18843);
nor UO_2253 (O_2253,N_16462,N_18346);
nor UO_2254 (O_2254,N_19338,N_16858);
or UO_2255 (O_2255,N_18371,N_19972);
nand UO_2256 (O_2256,N_15787,N_15529);
and UO_2257 (O_2257,N_15444,N_15936);
or UO_2258 (O_2258,N_17133,N_17076);
nand UO_2259 (O_2259,N_17425,N_19927);
nand UO_2260 (O_2260,N_19702,N_19278);
nor UO_2261 (O_2261,N_17964,N_18691);
or UO_2262 (O_2262,N_19597,N_15348);
xor UO_2263 (O_2263,N_19021,N_15398);
and UO_2264 (O_2264,N_16550,N_19682);
xor UO_2265 (O_2265,N_16680,N_19827);
nor UO_2266 (O_2266,N_19158,N_19386);
nand UO_2267 (O_2267,N_16889,N_19410);
or UO_2268 (O_2268,N_17797,N_16981);
nand UO_2269 (O_2269,N_15668,N_19200);
xnor UO_2270 (O_2270,N_15073,N_15463);
and UO_2271 (O_2271,N_16610,N_16282);
nand UO_2272 (O_2272,N_18001,N_17678);
and UO_2273 (O_2273,N_17410,N_16613);
xnor UO_2274 (O_2274,N_18945,N_18800);
or UO_2275 (O_2275,N_19156,N_18553);
and UO_2276 (O_2276,N_16719,N_15771);
or UO_2277 (O_2277,N_17560,N_18254);
xor UO_2278 (O_2278,N_19462,N_19813);
or UO_2279 (O_2279,N_17475,N_18374);
xnor UO_2280 (O_2280,N_16757,N_17781);
xnor UO_2281 (O_2281,N_17247,N_15379);
nand UO_2282 (O_2282,N_15803,N_15036);
and UO_2283 (O_2283,N_15328,N_15597);
or UO_2284 (O_2284,N_17994,N_17995);
and UO_2285 (O_2285,N_16432,N_19628);
nor UO_2286 (O_2286,N_19409,N_19944);
or UO_2287 (O_2287,N_19786,N_19441);
nand UO_2288 (O_2288,N_16837,N_19090);
and UO_2289 (O_2289,N_16572,N_15935);
nand UO_2290 (O_2290,N_15683,N_16103);
nand UO_2291 (O_2291,N_17899,N_19107);
and UO_2292 (O_2292,N_18675,N_17078);
nand UO_2293 (O_2293,N_17473,N_19213);
and UO_2294 (O_2294,N_15260,N_16666);
and UO_2295 (O_2295,N_19848,N_16306);
nor UO_2296 (O_2296,N_15170,N_18878);
or UO_2297 (O_2297,N_16644,N_17194);
nand UO_2298 (O_2298,N_18603,N_16875);
and UO_2299 (O_2299,N_16312,N_15594);
xnor UO_2300 (O_2300,N_15316,N_17706);
or UO_2301 (O_2301,N_16848,N_19306);
or UO_2302 (O_2302,N_18242,N_16334);
and UO_2303 (O_2303,N_17714,N_16216);
nor UO_2304 (O_2304,N_19080,N_18626);
or UO_2305 (O_2305,N_17586,N_19991);
xor UO_2306 (O_2306,N_15844,N_18047);
or UO_2307 (O_2307,N_15583,N_16515);
and UO_2308 (O_2308,N_15340,N_17705);
nand UO_2309 (O_2309,N_16503,N_18277);
xor UO_2310 (O_2310,N_19484,N_18190);
nor UO_2311 (O_2311,N_19009,N_19175);
nor UO_2312 (O_2312,N_15431,N_17949);
or UO_2313 (O_2313,N_15511,N_19948);
nand UO_2314 (O_2314,N_15630,N_15934);
nand UO_2315 (O_2315,N_15811,N_19562);
or UO_2316 (O_2316,N_17223,N_17996);
nand UO_2317 (O_2317,N_19271,N_19734);
xor UO_2318 (O_2318,N_19041,N_17658);
nor UO_2319 (O_2319,N_15979,N_15308);
and UO_2320 (O_2320,N_15277,N_18718);
and UO_2321 (O_2321,N_19796,N_16710);
and UO_2322 (O_2322,N_18123,N_17973);
or UO_2323 (O_2323,N_17480,N_18303);
and UO_2324 (O_2324,N_15322,N_19500);
nand UO_2325 (O_2325,N_19784,N_17266);
nor UO_2326 (O_2326,N_15535,N_19454);
nor UO_2327 (O_2327,N_18525,N_17470);
and UO_2328 (O_2328,N_19024,N_17192);
nor UO_2329 (O_2329,N_16711,N_16486);
xor UO_2330 (O_2330,N_15003,N_15189);
xor UO_2331 (O_2331,N_19002,N_17188);
or UO_2332 (O_2332,N_16908,N_18612);
and UO_2333 (O_2333,N_18696,N_16408);
or UO_2334 (O_2334,N_15429,N_17691);
xor UO_2335 (O_2335,N_18029,N_18873);
or UO_2336 (O_2336,N_16988,N_15688);
or UO_2337 (O_2337,N_17092,N_19111);
nand UO_2338 (O_2338,N_19173,N_17207);
or UO_2339 (O_2339,N_16309,N_17857);
and UO_2340 (O_2340,N_18402,N_17640);
nor UO_2341 (O_2341,N_17050,N_16779);
and UO_2342 (O_2342,N_18469,N_17178);
nor UO_2343 (O_2343,N_15266,N_15743);
or UO_2344 (O_2344,N_17198,N_15812);
or UO_2345 (O_2345,N_17001,N_18382);
xor UO_2346 (O_2346,N_15759,N_16368);
xor UO_2347 (O_2347,N_18339,N_15209);
nand UO_2348 (O_2348,N_15125,N_15192);
nand UO_2349 (O_2349,N_17703,N_15707);
or UO_2350 (O_2350,N_17387,N_17258);
xnor UO_2351 (O_2351,N_15880,N_15190);
nor UO_2352 (O_2352,N_17477,N_15772);
or UO_2353 (O_2353,N_18330,N_19681);
nand UO_2354 (O_2354,N_15813,N_16953);
nand UO_2355 (O_2355,N_17506,N_18662);
or UO_2356 (O_2356,N_15576,N_18996);
and UO_2357 (O_2357,N_17124,N_17418);
nand UO_2358 (O_2358,N_15564,N_19180);
or UO_2359 (O_2359,N_18763,N_18711);
nor UO_2360 (O_2360,N_17591,N_17901);
and UO_2361 (O_2361,N_17813,N_16693);
nand UO_2362 (O_2362,N_16793,N_19803);
or UO_2363 (O_2363,N_16840,N_19406);
and UO_2364 (O_2364,N_15650,N_17565);
or UO_2365 (O_2365,N_18080,N_19709);
nor UO_2366 (O_2366,N_17083,N_16345);
or UO_2367 (O_2367,N_15393,N_19222);
nor UO_2368 (O_2368,N_17419,N_19364);
xor UO_2369 (O_2369,N_19026,N_18773);
nor UO_2370 (O_2370,N_19528,N_16222);
nand UO_2371 (O_2371,N_17934,N_19330);
xnor UO_2372 (O_2372,N_18852,N_18200);
and UO_2373 (O_2373,N_17945,N_18907);
nor UO_2374 (O_2374,N_16087,N_15001);
nand UO_2375 (O_2375,N_16671,N_17684);
or UO_2376 (O_2376,N_19117,N_18283);
nand UO_2377 (O_2377,N_17038,N_17742);
nand UO_2378 (O_2378,N_17211,N_18285);
xnor UO_2379 (O_2379,N_15425,N_16376);
nor UO_2380 (O_2380,N_16417,N_15359);
xor UO_2381 (O_2381,N_17131,N_19885);
xor UO_2382 (O_2382,N_17952,N_18613);
nor UO_2383 (O_2383,N_19210,N_18983);
and UO_2384 (O_2384,N_18680,N_16668);
or UO_2385 (O_2385,N_19290,N_19721);
nand UO_2386 (O_2386,N_17671,N_16247);
nand UO_2387 (O_2387,N_17981,N_19344);
nor UO_2388 (O_2388,N_16469,N_16339);
and UO_2389 (O_2389,N_15956,N_17501);
xor UO_2390 (O_2390,N_17476,N_15106);
and UO_2391 (O_2391,N_19353,N_18344);
xnor UO_2392 (O_2392,N_19843,N_18089);
nand UO_2393 (O_2393,N_16781,N_19396);
xnor UO_2394 (O_2394,N_16439,N_17772);
and UO_2395 (O_2395,N_16219,N_19496);
or UO_2396 (O_2396,N_19334,N_15715);
or UO_2397 (O_2397,N_15284,N_17541);
nor UO_2398 (O_2398,N_18881,N_15401);
nor UO_2399 (O_2399,N_19653,N_16603);
nand UO_2400 (O_2400,N_16511,N_15123);
xor UO_2401 (O_2401,N_17843,N_18279);
nor UO_2402 (O_2402,N_19096,N_15173);
nor UO_2403 (O_2403,N_17231,N_17444);
and UO_2404 (O_2404,N_17790,N_18669);
nand UO_2405 (O_2405,N_18661,N_18958);
and UO_2406 (O_2406,N_15299,N_17340);
nand UO_2407 (O_2407,N_17548,N_17629);
xor UO_2408 (O_2408,N_15353,N_16695);
and UO_2409 (O_2409,N_15324,N_19327);
xnor UO_2410 (O_2410,N_18877,N_18489);
and UO_2411 (O_2411,N_16051,N_15996);
nand UO_2412 (O_2412,N_19825,N_17241);
nor UO_2413 (O_2413,N_17127,N_18580);
and UO_2414 (O_2414,N_18221,N_16304);
nand UO_2415 (O_2415,N_18213,N_19815);
xnor UO_2416 (O_2416,N_19463,N_16982);
or UO_2417 (O_2417,N_19193,N_19979);
and UO_2418 (O_2418,N_18486,N_19911);
or UO_2419 (O_2419,N_19760,N_17544);
xor UO_2420 (O_2420,N_17900,N_17633);
xor UO_2421 (O_2421,N_18501,N_18150);
and UO_2422 (O_2422,N_18595,N_15734);
nand UO_2423 (O_2423,N_19017,N_18784);
nand UO_2424 (O_2424,N_15222,N_15009);
or UO_2425 (O_2425,N_15301,N_17170);
nand UO_2426 (O_2426,N_19665,N_16302);
and UO_2427 (O_2427,N_18670,N_17184);
or UO_2428 (O_2428,N_15637,N_15397);
or UO_2429 (O_2429,N_16751,N_18615);
xor UO_2430 (O_2430,N_18621,N_15983);
nand UO_2431 (O_2431,N_15136,N_18990);
and UO_2432 (O_2432,N_17024,N_16413);
nor UO_2433 (O_2433,N_15129,N_17509);
nor UO_2434 (O_2434,N_19970,N_18229);
and UO_2435 (O_2435,N_16938,N_18534);
nand UO_2436 (O_2436,N_19742,N_15408);
and UO_2437 (O_2437,N_15959,N_16539);
or UO_2438 (O_2438,N_17302,N_17993);
or UO_2439 (O_2439,N_18536,N_19814);
nor UO_2440 (O_2440,N_19546,N_19351);
nor UO_2441 (O_2441,N_19988,N_18021);
nand UO_2442 (O_2442,N_19238,N_15283);
or UO_2443 (O_2443,N_17626,N_16800);
and UO_2444 (O_2444,N_15658,N_15705);
xnor UO_2445 (O_2445,N_15680,N_15264);
xor UO_2446 (O_2446,N_16859,N_15371);
nand UO_2447 (O_2447,N_17066,N_18450);
xnor UO_2448 (O_2448,N_15092,N_19013);
or UO_2449 (O_2449,N_19730,N_17752);
nor UO_2450 (O_2450,N_16529,N_15049);
and UO_2451 (O_2451,N_19102,N_17060);
nand UO_2452 (O_2452,N_17815,N_18055);
xnor UO_2453 (O_2453,N_18500,N_19581);
nand UO_2454 (O_2454,N_19776,N_18686);
nand UO_2455 (O_2455,N_19258,N_17250);
nor UO_2456 (O_2456,N_19822,N_17997);
nand UO_2457 (O_2457,N_16843,N_15122);
nand UO_2458 (O_2458,N_15201,N_16161);
and UO_2459 (O_2459,N_15541,N_15333);
xnor UO_2460 (O_2460,N_18497,N_18153);
xnor UO_2461 (O_2461,N_15950,N_15540);
nand UO_2462 (O_2462,N_16262,N_15051);
and UO_2463 (O_2463,N_18037,N_18523);
xnor UO_2464 (O_2464,N_17312,N_16992);
or UO_2465 (O_2465,N_15471,N_15923);
or UO_2466 (O_2466,N_16058,N_19456);
nand UO_2467 (O_2467,N_19477,N_18734);
nand UO_2468 (O_2468,N_19931,N_16679);
or UO_2469 (O_2469,N_15810,N_15166);
and UO_2470 (O_2470,N_16513,N_17345);
xor UO_2471 (O_2471,N_19658,N_15784);
nor UO_2472 (O_2472,N_19227,N_16149);
xor UO_2473 (O_2473,N_18202,N_15033);
nand UO_2474 (O_2474,N_19626,N_18746);
nor UO_2475 (O_2475,N_15017,N_18338);
or UO_2476 (O_2476,N_15568,N_17141);
nor UO_2477 (O_2477,N_17787,N_15473);
nand UO_2478 (O_2478,N_16924,N_16685);
or UO_2479 (O_2479,N_15724,N_15034);
xnor UO_2480 (O_2480,N_18738,N_17143);
and UO_2481 (O_2481,N_17072,N_18396);
and UO_2482 (O_2482,N_15492,N_17263);
nor UO_2483 (O_2483,N_18030,N_19340);
or UO_2484 (O_2484,N_17227,N_17682);
xnor UO_2485 (O_2485,N_15826,N_16574);
nor UO_2486 (O_2486,N_16335,N_17118);
nor UO_2487 (O_2487,N_16854,N_15638);
or UO_2488 (O_2488,N_19621,N_17471);
nor UO_2489 (O_2489,N_19720,N_16488);
or UO_2490 (O_2490,N_17830,N_19050);
nor UO_2491 (O_2491,N_19138,N_19797);
nor UO_2492 (O_2492,N_18896,N_19933);
and UO_2493 (O_2493,N_16070,N_15014);
or UO_2494 (O_2494,N_16204,N_15611);
and UO_2495 (O_2495,N_18748,N_15499);
nand UO_2496 (O_2496,N_15048,N_16323);
or UO_2497 (O_2497,N_15257,N_17265);
nand UO_2498 (O_2498,N_15832,N_18549);
xnor UO_2499 (O_2499,N_17248,N_15160);
endmodule