module basic_500_3000_500_3_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_365,In_139);
nor U1 (N_1,In_163,In_313);
xnor U2 (N_2,In_473,In_128);
nor U3 (N_3,In_253,In_434);
xnor U4 (N_4,In_226,In_36);
or U5 (N_5,In_414,In_421);
or U6 (N_6,In_146,In_111);
nor U7 (N_7,In_138,In_420);
and U8 (N_8,In_415,In_378);
nor U9 (N_9,In_45,In_57);
or U10 (N_10,In_21,In_323);
nor U11 (N_11,In_471,In_364);
and U12 (N_12,In_393,In_204);
and U13 (N_13,In_379,In_217);
nand U14 (N_14,In_145,In_133);
nor U15 (N_15,In_2,In_126);
or U16 (N_16,In_429,In_108);
nor U17 (N_17,In_93,In_412);
or U18 (N_18,In_293,In_302);
nand U19 (N_19,In_453,In_181);
or U20 (N_20,In_458,In_372);
xor U21 (N_21,In_148,In_477);
and U22 (N_22,In_123,In_152);
xnor U23 (N_23,In_284,In_220);
or U24 (N_24,In_349,In_416);
nor U25 (N_25,In_258,In_292);
nor U26 (N_26,In_10,In_265);
or U27 (N_27,In_358,In_362);
nor U28 (N_28,In_306,In_264);
nor U29 (N_29,In_81,In_476);
xnor U30 (N_30,In_244,In_374);
xor U31 (N_31,In_316,In_247);
and U32 (N_32,In_350,In_41);
and U33 (N_33,In_483,In_248);
and U34 (N_34,In_96,In_74);
and U35 (N_35,In_337,In_418);
xnor U36 (N_36,In_427,In_67);
or U37 (N_37,In_219,In_94);
nand U38 (N_38,In_1,In_147);
nand U39 (N_39,In_407,In_328);
xnor U40 (N_40,In_12,In_485);
xor U41 (N_41,In_66,In_245);
xor U42 (N_42,In_326,In_327);
xnor U43 (N_43,In_363,In_272);
and U44 (N_44,In_209,In_411);
nor U45 (N_45,In_406,In_17);
nand U46 (N_46,In_353,In_54);
or U47 (N_47,In_428,In_391);
xor U48 (N_48,In_63,In_296);
nor U49 (N_49,In_381,In_491);
nand U50 (N_50,In_396,In_212);
or U51 (N_51,In_444,In_165);
or U52 (N_52,In_334,In_84);
nor U53 (N_53,In_62,In_461);
and U54 (N_54,In_102,In_210);
nand U55 (N_55,In_154,In_254);
nor U56 (N_56,In_143,In_311);
and U57 (N_57,In_120,In_338);
xnor U58 (N_58,In_125,In_443);
and U59 (N_59,In_73,In_236);
nor U60 (N_60,In_256,In_282);
nand U61 (N_61,In_371,In_179);
and U62 (N_62,In_270,In_164);
or U63 (N_63,In_26,In_392);
xnor U64 (N_64,In_35,In_127);
xnor U65 (N_65,In_169,In_174);
nand U66 (N_66,In_95,In_50);
nand U67 (N_67,In_42,In_425);
and U68 (N_68,In_173,In_86);
xor U69 (N_69,In_319,In_118);
nand U70 (N_70,In_184,In_195);
nand U71 (N_71,In_69,In_442);
nor U72 (N_72,In_439,In_330);
and U73 (N_73,In_250,In_99);
nand U74 (N_74,In_33,In_225);
and U75 (N_75,In_7,In_390);
nor U76 (N_76,In_433,In_333);
or U77 (N_77,In_101,In_497);
nand U78 (N_78,In_355,In_494);
xor U79 (N_79,In_5,In_263);
xor U80 (N_80,In_80,In_377);
and U81 (N_81,In_214,In_159);
xnor U82 (N_82,In_186,In_470);
xnor U83 (N_83,In_499,In_322);
nor U84 (N_84,In_329,In_395);
nor U85 (N_85,In_142,In_397);
nand U86 (N_86,In_233,In_340);
xnor U87 (N_87,In_230,In_277);
or U88 (N_88,In_175,In_375);
and U89 (N_89,In_274,In_246);
nand U90 (N_90,In_177,In_75);
and U91 (N_91,In_493,In_287);
nor U92 (N_92,In_198,In_281);
nor U93 (N_93,In_369,In_388);
xnor U94 (N_94,In_417,In_294);
nor U95 (N_95,In_200,In_279);
nor U96 (N_96,In_64,In_71);
or U97 (N_97,In_20,In_240);
nor U98 (N_98,In_110,In_347);
or U99 (N_99,In_280,In_76);
xor U100 (N_100,In_467,In_91);
or U101 (N_101,In_342,In_426);
nand U102 (N_102,In_44,In_484);
or U103 (N_103,In_6,In_43);
and U104 (N_104,In_47,In_180);
or U105 (N_105,In_162,In_8);
or U106 (N_106,In_314,In_399);
or U107 (N_107,In_114,In_90);
xor U108 (N_108,In_141,In_83);
or U109 (N_109,In_380,In_295);
nand U110 (N_110,In_432,In_131);
nor U111 (N_111,In_239,In_482);
nand U112 (N_112,In_341,In_437);
and U113 (N_113,In_384,In_359);
or U114 (N_114,In_385,In_413);
nor U115 (N_115,In_304,In_52);
nand U116 (N_116,In_24,In_495);
or U117 (N_117,In_419,In_53);
and U118 (N_118,In_194,In_273);
nand U119 (N_119,In_153,In_121);
nor U120 (N_120,In_234,In_29);
nor U121 (N_121,In_197,In_192);
or U122 (N_122,In_58,In_171);
nor U123 (N_123,In_452,In_130);
nand U124 (N_124,In_367,In_344);
or U125 (N_125,In_100,In_435);
nand U126 (N_126,In_106,In_321);
xor U127 (N_127,In_144,In_136);
and U128 (N_128,In_0,In_278);
or U129 (N_129,In_223,In_262);
or U130 (N_130,In_455,In_157);
nor U131 (N_131,In_325,In_46);
xnor U132 (N_132,In_469,In_454);
and U133 (N_133,In_283,In_423);
nand U134 (N_134,In_215,In_348);
and U135 (N_135,In_436,In_297);
nand U136 (N_136,In_410,In_105);
xnor U137 (N_137,In_486,In_447);
nand U138 (N_138,In_109,In_431);
and U139 (N_139,In_383,In_16);
and U140 (N_140,In_150,In_261);
nand U141 (N_141,In_56,In_464);
nand U142 (N_142,In_113,In_68);
or U143 (N_143,In_373,In_267);
nand U144 (N_144,In_361,In_259);
nand U145 (N_145,In_465,In_370);
nor U146 (N_146,In_79,In_271);
or U147 (N_147,In_160,In_28);
nor U148 (N_148,In_88,In_14);
and U149 (N_149,In_167,In_22);
and U150 (N_150,In_199,In_360);
and U151 (N_151,In_85,In_156);
xnor U152 (N_152,In_135,In_496);
nor U153 (N_153,In_366,In_356);
nand U154 (N_154,In_13,In_104);
or U155 (N_155,In_51,In_237);
nor U156 (N_156,In_203,In_3);
nand U157 (N_157,In_345,In_227);
nor U158 (N_158,In_31,In_103);
nor U159 (N_159,In_404,In_206);
xor U160 (N_160,In_405,In_249);
nand U161 (N_161,In_290,In_300);
nand U162 (N_162,In_291,In_275);
and U163 (N_163,In_172,In_185);
and U164 (N_164,In_251,In_324);
or U165 (N_165,In_368,In_242);
nand U166 (N_166,In_232,In_107);
and U167 (N_167,In_309,In_466);
or U168 (N_168,In_424,In_401);
xnor U169 (N_169,In_55,In_346);
and U170 (N_170,In_307,In_243);
nor U171 (N_171,In_196,In_122);
nand U172 (N_172,In_301,In_389);
nor U173 (N_173,In_438,In_124);
nor U174 (N_174,In_305,In_409);
xor U175 (N_175,In_354,In_134);
nor U176 (N_176,In_229,In_216);
nor U177 (N_177,In_474,In_315);
or U178 (N_178,In_218,In_32);
nor U179 (N_179,In_288,In_317);
and U180 (N_180,In_11,In_176);
nand U181 (N_181,In_289,In_332);
xnor U182 (N_182,In_286,In_61);
nor U183 (N_183,In_459,In_137);
and U184 (N_184,In_231,In_190);
and U185 (N_185,In_201,In_463);
nor U186 (N_186,In_92,In_255);
or U187 (N_187,In_207,In_18);
or U188 (N_188,In_193,In_213);
xor U189 (N_189,In_49,In_205);
and U190 (N_190,In_40,In_394);
nand U191 (N_191,In_490,In_276);
and U192 (N_192,In_151,In_252);
nor U193 (N_193,In_402,In_158);
xnor U194 (N_194,In_189,In_89);
nor U195 (N_195,In_285,In_266);
or U196 (N_196,In_224,In_343);
nor U197 (N_197,In_446,In_422);
xor U198 (N_198,In_82,In_238);
nor U199 (N_199,In_87,In_450);
or U200 (N_200,In_487,In_257);
and U201 (N_201,In_38,In_187);
or U202 (N_202,In_30,In_166);
xnor U203 (N_203,In_312,In_129);
xor U204 (N_204,In_269,In_449);
or U205 (N_205,In_400,In_492);
xnor U206 (N_206,In_440,In_472);
or U207 (N_207,In_115,In_468);
or U208 (N_208,In_456,In_72);
nor U209 (N_209,In_116,In_132);
nor U210 (N_210,In_310,In_318);
xnor U211 (N_211,In_303,In_112);
xnor U212 (N_212,In_228,In_335);
or U213 (N_213,In_19,In_59);
xnor U214 (N_214,In_149,In_117);
xnor U215 (N_215,In_119,In_320);
xor U216 (N_216,In_48,In_60);
nand U217 (N_217,In_140,In_357);
nand U218 (N_218,In_479,In_408);
or U219 (N_219,In_386,In_268);
xor U220 (N_220,In_308,In_235);
or U221 (N_221,In_191,In_298);
and U222 (N_222,In_445,In_382);
or U223 (N_223,In_448,In_25);
nor U224 (N_224,In_481,In_65);
xnor U225 (N_225,In_488,In_498);
nand U226 (N_226,In_168,In_241);
and U227 (N_227,In_183,In_331);
or U228 (N_228,In_352,In_155);
xor U229 (N_229,In_182,In_480);
xnor U230 (N_230,In_387,In_34);
or U231 (N_231,In_15,In_462);
nor U232 (N_232,In_460,In_430);
and U233 (N_233,In_170,In_37);
xnor U234 (N_234,In_475,In_77);
xor U235 (N_235,In_489,In_457);
nor U236 (N_236,In_70,In_202);
xor U237 (N_237,In_451,In_403);
or U238 (N_238,In_441,In_188);
nor U239 (N_239,In_221,In_23);
nand U240 (N_240,In_97,In_78);
or U241 (N_241,In_336,In_478);
nor U242 (N_242,In_178,In_376);
nand U243 (N_243,In_161,In_9);
or U244 (N_244,In_4,In_27);
nor U245 (N_245,In_98,In_39);
or U246 (N_246,In_299,In_222);
nand U247 (N_247,In_398,In_351);
nor U248 (N_248,In_208,In_260);
nor U249 (N_249,In_339,In_211);
xor U250 (N_250,In_105,In_224);
or U251 (N_251,In_406,In_472);
nand U252 (N_252,In_362,In_488);
or U253 (N_253,In_275,In_478);
nand U254 (N_254,In_233,In_133);
and U255 (N_255,In_224,In_333);
xor U256 (N_256,In_119,In_162);
xor U257 (N_257,In_144,In_347);
xnor U258 (N_258,In_395,In_289);
and U259 (N_259,In_460,In_385);
nor U260 (N_260,In_103,In_454);
nor U261 (N_261,In_228,In_264);
or U262 (N_262,In_307,In_479);
and U263 (N_263,In_41,In_92);
nand U264 (N_264,In_423,In_104);
and U265 (N_265,In_32,In_172);
nand U266 (N_266,In_255,In_64);
or U267 (N_267,In_128,In_29);
nor U268 (N_268,In_323,In_372);
or U269 (N_269,In_401,In_486);
nor U270 (N_270,In_396,In_65);
and U271 (N_271,In_39,In_324);
xor U272 (N_272,In_225,In_180);
and U273 (N_273,In_276,In_217);
xor U274 (N_274,In_429,In_265);
and U275 (N_275,In_460,In_310);
xor U276 (N_276,In_477,In_412);
nor U277 (N_277,In_134,In_314);
or U278 (N_278,In_269,In_353);
nor U279 (N_279,In_395,In_401);
xnor U280 (N_280,In_58,In_168);
or U281 (N_281,In_76,In_10);
xnor U282 (N_282,In_138,In_499);
or U283 (N_283,In_344,In_175);
or U284 (N_284,In_265,In_313);
or U285 (N_285,In_108,In_128);
and U286 (N_286,In_144,In_141);
or U287 (N_287,In_282,In_409);
and U288 (N_288,In_19,In_366);
nand U289 (N_289,In_494,In_103);
or U290 (N_290,In_394,In_49);
xnor U291 (N_291,In_386,In_59);
nand U292 (N_292,In_125,In_45);
xor U293 (N_293,In_481,In_314);
xor U294 (N_294,In_433,In_245);
nand U295 (N_295,In_367,In_467);
or U296 (N_296,In_303,In_196);
and U297 (N_297,In_153,In_386);
xor U298 (N_298,In_493,In_200);
and U299 (N_299,In_216,In_17);
and U300 (N_300,In_281,In_64);
xor U301 (N_301,In_152,In_378);
nand U302 (N_302,In_212,In_220);
and U303 (N_303,In_213,In_258);
nor U304 (N_304,In_458,In_352);
or U305 (N_305,In_464,In_280);
nand U306 (N_306,In_340,In_47);
or U307 (N_307,In_299,In_386);
xor U308 (N_308,In_98,In_351);
or U309 (N_309,In_440,In_278);
nor U310 (N_310,In_286,In_20);
xor U311 (N_311,In_119,In_225);
and U312 (N_312,In_378,In_160);
nand U313 (N_313,In_47,In_204);
nand U314 (N_314,In_401,In_83);
nand U315 (N_315,In_42,In_179);
and U316 (N_316,In_266,In_336);
or U317 (N_317,In_434,In_292);
or U318 (N_318,In_307,In_75);
or U319 (N_319,In_266,In_308);
or U320 (N_320,In_370,In_233);
xor U321 (N_321,In_199,In_339);
nor U322 (N_322,In_37,In_430);
and U323 (N_323,In_171,In_362);
or U324 (N_324,In_120,In_113);
or U325 (N_325,In_141,In_204);
xnor U326 (N_326,In_245,In_464);
nor U327 (N_327,In_185,In_355);
xnor U328 (N_328,In_490,In_88);
or U329 (N_329,In_368,In_4);
xnor U330 (N_330,In_426,In_9);
nor U331 (N_331,In_197,In_339);
or U332 (N_332,In_190,In_176);
xor U333 (N_333,In_23,In_357);
xor U334 (N_334,In_254,In_24);
or U335 (N_335,In_397,In_411);
and U336 (N_336,In_42,In_88);
xnor U337 (N_337,In_98,In_151);
nor U338 (N_338,In_340,In_367);
or U339 (N_339,In_326,In_342);
and U340 (N_340,In_459,In_196);
nand U341 (N_341,In_73,In_365);
and U342 (N_342,In_238,In_314);
nor U343 (N_343,In_413,In_22);
xnor U344 (N_344,In_453,In_481);
nor U345 (N_345,In_152,In_294);
nor U346 (N_346,In_261,In_16);
nand U347 (N_347,In_368,In_450);
nor U348 (N_348,In_155,In_84);
xnor U349 (N_349,In_188,In_349);
nor U350 (N_350,In_296,In_17);
nor U351 (N_351,In_338,In_432);
nand U352 (N_352,In_19,In_138);
xor U353 (N_353,In_378,In_265);
and U354 (N_354,In_276,In_404);
nor U355 (N_355,In_268,In_32);
xnor U356 (N_356,In_479,In_60);
and U357 (N_357,In_234,In_309);
and U358 (N_358,In_259,In_485);
xor U359 (N_359,In_201,In_481);
nor U360 (N_360,In_236,In_477);
nor U361 (N_361,In_400,In_427);
or U362 (N_362,In_198,In_434);
xor U363 (N_363,In_55,In_181);
nand U364 (N_364,In_317,In_155);
xnor U365 (N_365,In_288,In_444);
xor U366 (N_366,In_333,In_123);
nor U367 (N_367,In_486,In_254);
or U368 (N_368,In_46,In_65);
or U369 (N_369,In_129,In_453);
and U370 (N_370,In_482,In_387);
xor U371 (N_371,In_84,In_290);
and U372 (N_372,In_342,In_348);
nor U373 (N_373,In_373,In_423);
or U374 (N_374,In_49,In_166);
xnor U375 (N_375,In_213,In_131);
nand U376 (N_376,In_162,In_149);
nand U377 (N_377,In_404,In_218);
xnor U378 (N_378,In_141,In_299);
and U379 (N_379,In_319,In_30);
and U380 (N_380,In_74,In_262);
nor U381 (N_381,In_257,In_129);
and U382 (N_382,In_155,In_135);
or U383 (N_383,In_364,In_128);
nand U384 (N_384,In_453,In_480);
xnor U385 (N_385,In_361,In_376);
or U386 (N_386,In_273,In_298);
nor U387 (N_387,In_102,In_441);
xnor U388 (N_388,In_276,In_284);
nand U389 (N_389,In_131,In_224);
or U390 (N_390,In_19,In_205);
nor U391 (N_391,In_438,In_148);
nor U392 (N_392,In_54,In_19);
and U393 (N_393,In_467,In_149);
or U394 (N_394,In_371,In_19);
xor U395 (N_395,In_362,In_294);
or U396 (N_396,In_48,In_15);
nand U397 (N_397,In_1,In_390);
nand U398 (N_398,In_419,In_86);
or U399 (N_399,In_303,In_323);
xor U400 (N_400,In_401,In_286);
nand U401 (N_401,In_387,In_173);
xnor U402 (N_402,In_245,In_19);
or U403 (N_403,In_293,In_233);
xnor U404 (N_404,In_266,In_286);
and U405 (N_405,In_462,In_391);
nor U406 (N_406,In_417,In_286);
nor U407 (N_407,In_7,In_332);
or U408 (N_408,In_177,In_322);
nand U409 (N_409,In_232,In_386);
and U410 (N_410,In_241,In_98);
or U411 (N_411,In_73,In_252);
nand U412 (N_412,In_82,In_331);
and U413 (N_413,In_41,In_31);
xnor U414 (N_414,In_337,In_148);
nor U415 (N_415,In_66,In_113);
xnor U416 (N_416,In_484,In_220);
nor U417 (N_417,In_57,In_442);
xor U418 (N_418,In_283,In_489);
nand U419 (N_419,In_161,In_251);
nor U420 (N_420,In_167,In_368);
xor U421 (N_421,In_477,In_344);
nand U422 (N_422,In_282,In_170);
nand U423 (N_423,In_106,In_164);
nand U424 (N_424,In_466,In_44);
or U425 (N_425,In_245,In_107);
nand U426 (N_426,In_380,In_210);
or U427 (N_427,In_207,In_275);
and U428 (N_428,In_13,In_179);
nor U429 (N_429,In_479,In_84);
xor U430 (N_430,In_355,In_215);
nand U431 (N_431,In_135,In_484);
xnor U432 (N_432,In_74,In_256);
nor U433 (N_433,In_373,In_453);
xnor U434 (N_434,In_285,In_332);
or U435 (N_435,In_87,In_391);
nor U436 (N_436,In_371,In_75);
nand U437 (N_437,In_267,In_243);
nand U438 (N_438,In_243,In_334);
xor U439 (N_439,In_234,In_300);
xor U440 (N_440,In_425,In_99);
or U441 (N_441,In_318,In_393);
and U442 (N_442,In_284,In_437);
or U443 (N_443,In_16,In_371);
nor U444 (N_444,In_209,In_132);
or U445 (N_445,In_342,In_483);
or U446 (N_446,In_358,In_174);
nand U447 (N_447,In_381,In_101);
nor U448 (N_448,In_481,In_361);
xnor U449 (N_449,In_238,In_84);
nor U450 (N_450,In_368,In_77);
and U451 (N_451,In_37,In_284);
or U452 (N_452,In_38,In_293);
nor U453 (N_453,In_136,In_149);
nor U454 (N_454,In_369,In_201);
nor U455 (N_455,In_388,In_410);
xnor U456 (N_456,In_406,In_59);
nor U457 (N_457,In_347,In_496);
xor U458 (N_458,In_48,In_315);
or U459 (N_459,In_122,In_396);
and U460 (N_460,In_478,In_413);
and U461 (N_461,In_131,In_236);
nand U462 (N_462,In_90,In_359);
nand U463 (N_463,In_170,In_419);
xnor U464 (N_464,In_65,In_169);
xor U465 (N_465,In_474,In_465);
or U466 (N_466,In_333,In_117);
nor U467 (N_467,In_88,In_457);
nor U468 (N_468,In_88,In_54);
and U469 (N_469,In_489,In_2);
nor U470 (N_470,In_205,In_119);
and U471 (N_471,In_336,In_119);
xnor U472 (N_472,In_480,In_457);
nand U473 (N_473,In_416,In_145);
nand U474 (N_474,In_136,In_59);
nand U475 (N_475,In_436,In_485);
and U476 (N_476,In_396,In_36);
and U477 (N_477,In_126,In_336);
nor U478 (N_478,In_118,In_222);
xnor U479 (N_479,In_97,In_277);
or U480 (N_480,In_62,In_400);
nand U481 (N_481,In_55,In_248);
nand U482 (N_482,In_69,In_378);
and U483 (N_483,In_232,In_199);
xnor U484 (N_484,In_7,In_350);
nand U485 (N_485,In_419,In_238);
xor U486 (N_486,In_97,In_127);
nand U487 (N_487,In_171,In_330);
or U488 (N_488,In_249,In_146);
or U489 (N_489,In_217,In_248);
nor U490 (N_490,In_425,In_338);
nor U491 (N_491,In_42,In_193);
nor U492 (N_492,In_12,In_283);
nor U493 (N_493,In_435,In_436);
or U494 (N_494,In_455,In_273);
nand U495 (N_495,In_258,In_124);
and U496 (N_496,In_407,In_406);
nand U497 (N_497,In_116,In_344);
nand U498 (N_498,In_334,In_283);
or U499 (N_499,In_434,In_258);
and U500 (N_500,In_352,In_357);
nor U501 (N_501,In_206,In_215);
or U502 (N_502,In_334,In_32);
xnor U503 (N_503,In_339,In_379);
or U504 (N_504,In_285,In_172);
xor U505 (N_505,In_99,In_217);
nand U506 (N_506,In_318,In_62);
nor U507 (N_507,In_95,In_369);
or U508 (N_508,In_190,In_322);
nand U509 (N_509,In_321,In_260);
nor U510 (N_510,In_384,In_424);
nor U511 (N_511,In_32,In_56);
nor U512 (N_512,In_444,In_470);
nand U513 (N_513,In_300,In_132);
nor U514 (N_514,In_138,In_488);
or U515 (N_515,In_171,In_426);
nor U516 (N_516,In_452,In_125);
nand U517 (N_517,In_235,In_113);
xnor U518 (N_518,In_437,In_325);
nand U519 (N_519,In_13,In_411);
nor U520 (N_520,In_136,In_389);
nor U521 (N_521,In_235,In_100);
nand U522 (N_522,In_166,In_410);
and U523 (N_523,In_167,In_116);
nor U524 (N_524,In_124,In_84);
nand U525 (N_525,In_381,In_170);
nand U526 (N_526,In_171,In_251);
xnor U527 (N_527,In_29,In_493);
and U528 (N_528,In_0,In_382);
nand U529 (N_529,In_359,In_197);
nand U530 (N_530,In_156,In_40);
or U531 (N_531,In_295,In_9);
nor U532 (N_532,In_423,In_327);
or U533 (N_533,In_250,In_293);
and U534 (N_534,In_36,In_366);
nor U535 (N_535,In_230,In_368);
nand U536 (N_536,In_117,In_152);
or U537 (N_537,In_299,In_237);
xor U538 (N_538,In_497,In_465);
or U539 (N_539,In_465,In_58);
and U540 (N_540,In_103,In_221);
nand U541 (N_541,In_395,In_480);
or U542 (N_542,In_16,In_415);
or U543 (N_543,In_462,In_336);
nand U544 (N_544,In_391,In_284);
nand U545 (N_545,In_368,In_84);
or U546 (N_546,In_385,In_30);
xor U547 (N_547,In_443,In_302);
or U548 (N_548,In_146,In_287);
xnor U549 (N_549,In_214,In_390);
nor U550 (N_550,In_390,In_14);
xnor U551 (N_551,In_484,In_166);
and U552 (N_552,In_444,In_56);
nor U553 (N_553,In_470,In_133);
xor U554 (N_554,In_244,In_152);
xnor U555 (N_555,In_85,In_74);
nor U556 (N_556,In_38,In_492);
nor U557 (N_557,In_160,In_3);
nand U558 (N_558,In_466,In_355);
and U559 (N_559,In_182,In_358);
xnor U560 (N_560,In_95,In_92);
nor U561 (N_561,In_152,In_462);
nor U562 (N_562,In_454,In_166);
xor U563 (N_563,In_462,In_107);
or U564 (N_564,In_124,In_144);
and U565 (N_565,In_258,In_225);
nor U566 (N_566,In_114,In_319);
nor U567 (N_567,In_228,In_265);
or U568 (N_568,In_492,In_295);
and U569 (N_569,In_319,In_3);
nor U570 (N_570,In_143,In_381);
xnor U571 (N_571,In_179,In_240);
nor U572 (N_572,In_41,In_166);
nand U573 (N_573,In_195,In_413);
nor U574 (N_574,In_309,In_468);
and U575 (N_575,In_170,In_130);
and U576 (N_576,In_306,In_335);
nor U577 (N_577,In_456,In_104);
and U578 (N_578,In_447,In_182);
nor U579 (N_579,In_9,In_122);
nand U580 (N_580,In_410,In_93);
and U581 (N_581,In_491,In_32);
and U582 (N_582,In_44,In_106);
or U583 (N_583,In_154,In_247);
nand U584 (N_584,In_198,In_262);
nor U585 (N_585,In_17,In_45);
nor U586 (N_586,In_296,In_406);
nand U587 (N_587,In_318,In_210);
nor U588 (N_588,In_412,In_73);
or U589 (N_589,In_421,In_236);
nor U590 (N_590,In_99,In_23);
or U591 (N_591,In_478,In_286);
or U592 (N_592,In_246,In_214);
nor U593 (N_593,In_152,In_97);
or U594 (N_594,In_279,In_485);
xnor U595 (N_595,In_302,In_39);
nand U596 (N_596,In_438,In_210);
xnor U597 (N_597,In_156,In_84);
or U598 (N_598,In_103,In_87);
nor U599 (N_599,In_323,In_498);
nor U600 (N_600,In_353,In_405);
xor U601 (N_601,In_284,In_170);
nor U602 (N_602,In_14,In_381);
and U603 (N_603,In_381,In_249);
nor U604 (N_604,In_341,In_388);
nand U605 (N_605,In_250,In_399);
or U606 (N_606,In_98,In_138);
or U607 (N_607,In_311,In_368);
nor U608 (N_608,In_289,In_339);
xnor U609 (N_609,In_315,In_91);
and U610 (N_610,In_62,In_69);
or U611 (N_611,In_208,In_339);
xnor U612 (N_612,In_66,In_329);
nand U613 (N_613,In_166,In_143);
nand U614 (N_614,In_365,In_87);
nor U615 (N_615,In_61,In_106);
xor U616 (N_616,In_187,In_173);
and U617 (N_617,In_404,In_178);
nor U618 (N_618,In_69,In_244);
nand U619 (N_619,In_160,In_49);
or U620 (N_620,In_94,In_22);
xnor U621 (N_621,In_268,In_295);
nand U622 (N_622,In_170,In_239);
nor U623 (N_623,In_35,In_326);
and U624 (N_624,In_396,In_100);
or U625 (N_625,In_137,In_119);
xnor U626 (N_626,In_252,In_341);
nor U627 (N_627,In_38,In_195);
xor U628 (N_628,In_27,In_79);
or U629 (N_629,In_329,In_227);
and U630 (N_630,In_81,In_271);
nand U631 (N_631,In_354,In_364);
or U632 (N_632,In_241,In_103);
nor U633 (N_633,In_181,In_141);
and U634 (N_634,In_319,In_268);
or U635 (N_635,In_343,In_82);
nand U636 (N_636,In_333,In_29);
xor U637 (N_637,In_267,In_91);
and U638 (N_638,In_140,In_112);
nor U639 (N_639,In_246,In_380);
and U640 (N_640,In_372,In_54);
xor U641 (N_641,In_300,In_359);
and U642 (N_642,In_342,In_36);
nor U643 (N_643,In_10,In_401);
nor U644 (N_644,In_458,In_178);
and U645 (N_645,In_310,In_270);
nand U646 (N_646,In_295,In_329);
or U647 (N_647,In_167,In_177);
nor U648 (N_648,In_472,In_288);
and U649 (N_649,In_394,In_459);
nand U650 (N_650,In_104,In_265);
nand U651 (N_651,In_301,In_156);
or U652 (N_652,In_95,In_154);
nand U653 (N_653,In_32,In_344);
or U654 (N_654,In_10,In_440);
nand U655 (N_655,In_180,In_419);
nor U656 (N_656,In_399,In_258);
or U657 (N_657,In_105,In_336);
nor U658 (N_658,In_51,In_485);
or U659 (N_659,In_213,In_374);
or U660 (N_660,In_468,In_306);
nor U661 (N_661,In_182,In_113);
and U662 (N_662,In_262,In_101);
nand U663 (N_663,In_491,In_127);
and U664 (N_664,In_195,In_69);
and U665 (N_665,In_5,In_86);
and U666 (N_666,In_404,In_70);
or U667 (N_667,In_125,In_326);
and U668 (N_668,In_243,In_251);
xor U669 (N_669,In_127,In_315);
nor U670 (N_670,In_424,In_144);
nor U671 (N_671,In_212,In_313);
and U672 (N_672,In_492,In_32);
nand U673 (N_673,In_109,In_289);
nand U674 (N_674,In_445,In_441);
xor U675 (N_675,In_202,In_13);
or U676 (N_676,In_132,In_382);
nand U677 (N_677,In_481,In_349);
nand U678 (N_678,In_314,In_429);
and U679 (N_679,In_339,In_446);
or U680 (N_680,In_337,In_261);
xnor U681 (N_681,In_126,In_317);
nor U682 (N_682,In_269,In_339);
nand U683 (N_683,In_445,In_136);
or U684 (N_684,In_182,In_49);
and U685 (N_685,In_251,In_94);
xor U686 (N_686,In_397,In_165);
or U687 (N_687,In_39,In_309);
or U688 (N_688,In_140,In_226);
or U689 (N_689,In_222,In_418);
xnor U690 (N_690,In_111,In_388);
xor U691 (N_691,In_344,In_472);
and U692 (N_692,In_33,In_305);
nand U693 (N_693,In_259,In_86);
nand U694 (N_694,In_164,In_63);
xnor U695 (N_695,In_473,In_109);
or U696 (N_696,In_386,In_74);
nor U697 (N_697,In_435,In_249);
and U698 (N_698,In_468,In_3);
and U699 (N_699,In_146,In_399);
nor U700 (N_700,In_66,In_417);
or U701 (N_701,In_20,In_185);
xor U702 (N_702,In_407,In_493);
xnor U703 (N_703,In_126,In_233);
nand U704 (N_704,In_125,In_414);
or U705 (N_705,In_248,In_477);
and U706 (N_706,In_27,In_340);
xor U707 (N_707,In_450,In_362);
and U708 (N_708,In_448,In_423);
xor U709 (N_709,In_436,In_168);
xnor U710 (N_710,In_319,In_28);
xnor U711 (N_711,In_456,In_397);
xnor U712 (N_712,In_16,In_8);
xor U713 (N_713,In_267,In_309);
and U714 (N_714,In_300,In_331);
nor U715 (N_715,In_28,In_213);
nor U716 (N_716,In_480,In_452);
or U717 (N_717,In_119,In_59);
nor U718 (N_718,In_239,In_127);
and U719 (N_719,In_402,In_439);
nand U720 (N_720,In_129,In_29);
nand U721 (N_721,In_212,In_364);
or U722 (N_722,In_412,In_120);
and U723 (N_723,In_174,In_240);
nand U724 (N_724,In_57,In_435);
and U725 (N_725,In_378,In_179);
or U726 (N_726,In_375,In_68);
nand U727 (N_727,In_90,In_272);
or U728 (N_728,In_398,In_309);
or U729 (N_729,In_301,In_12);
or U730 (N_730,In_298,In_400);
or U731 (N_731,In_81,In_153);
nor U732 (N_732,In_362,In_217);
or U733 (N_733,In_339,In_484);
or U734 (N_734,In_72,In_436);
or U735 (N_735,In_36,In_47);
nor U736 (N_736,In_59,In_357);
nor U737 (N_737,In_120,In_465);
and U738 (N_738,In_238,In_152);
or U739 (N_739,In_248,In_438);
or U740 (N_740,In_285,In_248);
xnor U741 (N_741,In_443,In_212);
nor U742 (N_742,In_490,In_23);
nand U743 (N_743,In_70,In_235);
xor U744 (N_744,In_243,In_301);
and U745 (N_745,In_341,In_274);
and U746 (N_746,In_497,In_28);
or U747 (N_747,In_294,In_358);
or U748 (N_748,In_349,In_232);
or U749 (N_749,In_109,In_258);
and U750 (N_750,In_416,In_273);
nand U751 (N_751,In_234,In_367);
or U752 (N_752,In_220,In_253);
and U753 (N_753,In_473,In_201);
nor U754 (N_754,In_415,In_220);
nand U755 (N_755,In_75,In_342);
nor U756 (N_756,In_418,In_7);
xor U757 (N_757,In_170,In_21);
nand U758 (N_758,In_469,In_263);
xor U759 (N_759,In_6,In_201);
or U760 (N_760,In_28,In_375);
nor U761 (N_761,In_441,In_350);
and U762 (N_762,In_103,In_118);
nor U763 (N_763,In_338,In_30);
nor U764 (N_764,In_143,In_38);
and U765 (N_765,In_224,In_326);
xor U766 (N_766,In_385,In_246);
or U767 (N_767,In_452,In_254);
or U768 (N_768,In_423,In_383);
xnor U769 (N_769,In_251,In_375);
xnor U770 (N_770,In_73,In_328);
xnor U771 (N_771,In_282,In_274);
xnor U772 (N_772,In_422,In_159);
nand U773 (N_773,In_93,In_100);
xnor U774 (N_774,In_305,In_306);
nor U775 (N_775,In_294,In_38);
nor U776 (N_776,In_271,In_331);
and U777 (N_777,In_7,In_414);
nor U778 (N_778,In_29,In_456);
nand U779 (N_779,In_79,In_42);
xor U780 (N_780,In_269,In_229);
xor U781 (N_781,In_173,In_418);
and U782 (N_782,In_38,In_151);
and U783 (N_783,In_87,In_116);
nand U784 (N_784,In_466,In_105);
or U785 (N_785,In_77,In_139);
or U786 (N_786,In_339,In_64);
or U787 (N_787,In_337,In_136);
nand U788 (N_788,In_206,In_91);
or U789 (N_789,In_14,In_306);
nor U790 (N_790,In_241,In_14);
or U791 (N_791,In_88,In_359);
and U792 (N_792,In_201,In_177);
or U793 (N_793,In_499,In_188);
and U794 (N_794,In_73,In_1);
nand U795 (N_795,In_447,In_333);
nand U796 (N_796,In_127,In_328);
or U797 (N_797,In_381,In_95);
nor U798 (N_798,In_361,In_194);
and U799 (N_799,In_400,In_179);
xor U800 (N_800,In_458,In_398);
and U801 (N_801,In_172,In_169);
and U802 (N_802,In_185,In_319);
xnor U803 (N_803,In_308,In_275);
nor U804 (N_804,In_126,In_390);
nand U805 (N_805,In_332,In_478);
and U806 (N_806,In_233,In_162);
nand U807 (N_807,In_429,In_262);
nor U808 (N_808,In_404,In_489);
nand U809 (N_809,In_151,In_220);
nor U810 (N_810,In_318,In_375);
nor U811 (N_811,In_14,In_482);
nor U812 (N_812,In_113,In_318);
nor U813 (N_813,In_481,In_342);
nand U814 (N_814,In_139,In_389);
nand U815 (N_815,In_151,In_269);
nor U816 (N_816,In_493,In_385);
nand U817 (N_817,In_92,In_258);
xor U818 (N_818,In_495,In_134);
nand U819 (N_819,In_67,In_200);
nor U820 (N_820,In_276,In_302);
and U821 (N_821,In_116,In_33);
xor U822 (N_822,In_24,In_368);
and U823 (N_823,In_480,In_442);
nor U824 (N_824,In_344,In_449);
nor U825 (N_825,In_4,In_181);
nor U826 (N_826,In_222,In_173);
nor U827 (N_827,In_142,In_165);
xnor U828 (N_828,In_362,In_102);
xnor U829 (N_829,In_473,In_43);
and U830 (N_830,In_139,In_89);
nand U831 (N_831,In_344,In_379);
nand U832 (N_832,In_260,In_147);
xnor U833 (N_833,In_498,In_341);
xnor U834 (N_834,In_189,In_265);
and U835 (N_835,In_276,In_425);
nand U836 (N_836,In_75,In_383);
nand U837 (N_837,In_163,In_268);
xor U838 (N_838,In_441,In_489);
nor U839 (N_839,In_133,In_389);
xnor U840 (N_840,In_442,In_122);
xor U841 (N_841,In_313,In_25);
xnor U842 (N_842,In_74,In_59);
nand U843 (N_843,In_277,In_257);
xor U844 (N_844,In_212,In_330);
or U845 (N_845,In_203,In_5);
or U846 (N_846,In_462,In_296);
nor U847 (N_847,In_131,In_246);
and U848 (N_848,In_122,In_253);
or U849 (N_849,In_58,In_411);
nand U850 (N_850,In_138,In_480);
xnor U851 (N_851,In_484,In_260);
nor U852 (N_852,In_451,In_326);
nor U853 (N_853,In_157,In_318);
and U854 (N_854,In_107,In_382);
xor U855 (N_855,In_90,In_414);
nand U856 (N_856,In_251,In_39);
nand U857 (N_857,In_164,In_428);
xor U858 (N_858,In_405,In_357);
or U859 (N_859,In_195,In_262);
nor U860 (N_860,In_46,In_468);
xnor U861 (N_861,In_80,In_284);
nand U862 (N_862,In_485,In_392);
and U863 (N_863,In_252,In_367);
or U864 (N_864,In_415,In_87);
nand U865 (N_865,In_403,In_188);
or U866 (N_866,In_148,In_478);
or U867 (N_867,In_206,In_368);
nand U868 (N_868,In_325,In_115);
and U869 (N_869,In_391,In_19);
xnor U870 (N_870,In_451,In_168);
or U871 (N_871,In_174,In_24);
or U872 (N_872,In_332,In_394);
and U873 (N_873,In_81,In_366);
nor U874 (N_874,In_91,In_486);
and U875 (N_875,In_286,In_98);
and U876 (N_876,In_128,In_103);
and U877 (N_877,In_20,In_349);
or U878 (N_878,In_236,In_136);
or U879 (N_879,In_261,In_9);
nand U880 (N_880,In_190,In_308);
xnor U881 (N_881,In_21,In_463);
and U882 (N_882,In_112,In_136);
or U883 (N_883,In_175,In_255);
xnor U884 (N_884,In_217,In_56);
and U885 (N_885,In_105,In_211);
nor U886 (N_886,In_207,In_162);
nand U887 (N_887,In_270,In_265);
and U888 (N_888,In_18,In_481);
or U889 (N_889,In_77,In_358);
xnor U890 (N_890,In_342,In_112);
and U891 (N_891,In_485,In_380);
and U892 (N_892,In_346,In_66);
or U893 (N_893,In_65,In_298);
and U894 (N_894,In_239,In_195);
nor U895 (N_895,In_257,In_238);
and U896 (N_896,In_48,In_32);
xnor U897 (N_897,In_457,In_368);
or U898 (N_898,In_244,In_428);
xor U899 (N_899,In_23,In_9);
and U900 (N_900,In_80,In_477);
and U901 (N_901,In_93,In_306);
xnor U902 (N_902,In_17,In_118);
nor U903 (N_903,In_21,In_89);
and U904 (N_904,In_468,In_260);
nor U905 (N_905,In_167,In_56);
or U906 (N_906,In_448,In_116);
or U907 (N_907,In_122,In_397);
or U908 (N_908,In_69,In_474);
xor U909 (N_909,In_407,In_59);
nor U910 (N_910,In_177,In_463);
xor U911 (N_911,In_351,In_126);
nor U912 (N_912,In_16,In_446);
nor U913 (N_913,In_226,In_4);
xor U914 (N_914,In_287,In_267);
or U915 (N_915,In_170,In_234);
and U916 (N_916,In_68,In_141);
nor U917 (N_917,In_244,In_21);
xnor U918 (N_918,In_437,In_199);
or U919 (N_919,In_85,In_148);
nand U920 (N_920,In_310,In_462);
xor U921 (N_921,In_325,In_20);
nand U922 (N_922,In_5,In_15);
or U923 (N_923,In_127,In_449);
nor U924 (N_924,In_167,In_391);
nand U925 (N_925,In_40,In_62);
and U926 (N_926,In_494,In_252);
xnor U927 (N_927,In_193,In_8);
nand U928 (N_928,In_117,In_119);
or U929 (N_929,In_88,In_399);
nand U930 (N_930,In_263,In_107);
and U931 (N_931,In_96,In_330);
xnor U932 (N_932,In_303,In_219);
nand U933 (N_933,In_107,In_97);
and U934 (N_934,In_160,In_444);
and U935 (N_935,In_193,In_125);
nor U936 (N_936,In_449,In_21);
or U937 (N_937,In_411,In_10);
and U938 (N_938,In_331,In_339);
or U939 (N_939,In_343,In_307);
and U940 (N_940,In_66,In_405);
nor U941 (N_941,In_139,In_84);
and U942 (N_942,In_89,In_96);
and U943 (N_943,In_414,In_137);
nand U944 (N_944,In_168,In_177);
nor U945 (N_945,In_455,In_358);
nor U946 (N_946,In_309,In_99);
and U947 (N_947,In_169,In_290);
nor U948 (N_948,In_328,In_162);
nor U949 (N_949,In_7,In_88);
nor U950 (N_950,In_153,In_244);
nor U951 (N_951,In_176,In_204);
nand U952 (N_952,In_18,In_423);
or U953 (N_953,In_223,In_98);
xnor U954 (N_954,In_47,In_168);
nor U955 (N_955,In_277,In_382);
nand U956 (N_956,In_249,In_485);
nor U957 (N_957,In_83,In_29);
nor U958 (N_958,In_299,In_80);
xnor U959 (N_959,In_318,In_20);
nor U960 (N_960,In_396,In_255);
nor U961 (N_961,In_396,In_136);
nor U962 (N_962,In_385,In_251);
nor U963 (N_963,In_357,In_428);
nor U964 (N_964,In_306,In_107);
nand U965 (N_965,In_102,In_159);
nand U966 (N_966,In_282,In_223);
or U967 (N_967,In_212,In_149);
and U968 (N_968,In_77,In_472);
and U969 (N_969,In_481,In_39);
nor U970 (N_970,In_97,In_172);
and U971 (N_971,In_483,In_114);
nor U972 (N_972,In_401,In_416);
xor U973 (N_973,In_10,In_367);
xor U974 (N_974,In_491,In_267);
or U975 (N_975,In_128,In_441);
xnor U976 (N_976,In_287,In_94);
or U977 (N_977,In_352,In_188);
nor U978 (N_978,In_317,In_413);
or U979 (N_979,In_243,In_158);
xnor U980 (N_980,In_181,In_249);
or U981 (N_981,In_68,In_470);
nor U982 (N_982,In_464,In_213);
and U983 (N_983,In_148,In_348);
xnor U984 (N_984,In_394,In_41);
nand U985 (N_985,In_398,In_467);
nor U986 (N_986,In_286,In_29);
and U987 (N_987,In_166,In_78);
and U988 (N_988,In_463,In_34);
nand U989 (N_989,In_51,In_24);
nor U990 (N_990,In_493,In_236);
and U991 (N_991,In_478,In_52);
xnor U992 (N_992,In_319,In_77);
nand U993 (N_993,In_229,In_301);
nand U994 (N_994,In_147,In_67);
nor U995 (N_995,In_183,In_233);
nor U996 (N_996,In_0,In_184);
xnor U997 (N_997,In_474,In_304);
nor U998 (N_998,In_49,In_275);
or U999 (N_999,In_390,In_11);
and U1000 (N_1000,N_866,N_153);
or U1001 (N_1001,N_584,N_771);
or U1002 (N_1002,N_593,N_420);
nand U1003 (N_1003,N_100,N_849);
and U1004 (N_1004,N_394,N_271);
nor U1005 (N_1005,N_66,N_257);
nor U1006 (N_1006,N_510,N_119);
nor U1007 (N_1007,N_506,N_450);
and U1008 (N_1008,N_497,N_10);
nor U1009 (N_1009,N_594,N_905);
nand U1010 (N_1010,N_609,N_799);
and U1011 (N_1011,N_143,N_174);
xor U1012 (N_1012,N_286,N_165);
and U1013 (N_1013,N_992,N_336);
nor U1014 (N_1014,N_5,N_562);
nor U1015 (N_1015,N_47,N_109);
and U1016 (N_1016,N_129,N_695);
nand U1017 (N_1017,N_735,N_163);
and U1018 (N_1018,N_534,N_171);
nand U1019 (N_1019,N_466,N_603);
and U1020 (N_1020,N_685,N_617);
and U1021 (N_1021,N_610,N_911);
nor U1022 (N_1022,N_488,N_242);
nand U1023 (N_1023,N_991,N_699);
or U1024 (N_1024,N_199,N_503);
nand U1025 (N_1025,N_878,N_983);
nand U1026 (N_1026,N_73,N_761);
or U1027 (N_1027,N_934,N_486);
nor U1028 (N_1028,N_445,N_106);
xor U1029 (N_1029,N_754,N_891);
and U1030 (N_1030,N_93,N_639);
xor U1031 (N_1031,N_181,N_985);
and U1032 (N_1032,N_736,N_720);
or U1033 (N_1033,N_104,N_46);
nand U1034 (N_1034,N_330,N_869);
or U1035 (N_1035,N_338,N_904);
and U1036 (N_1036,N_378,N_28);
xnor U1037 (N_1037,N_427,N_572);
and U1038 (N_1038,N_363,N_653);
or U1039 (N_1039,N_69,N_932);
or U1040 (N_1040,N_17,N_437);
nor U1041 (N_1041,N_600,N_725);
nand U1042 (N_1042,N_980,N_969);
and U1043 (N_1043,N_342,N_155);
xnor U1044 (N_1044,N_813,N_555);
and U1045 (N_1045,N_894,N_60);
nand U1046 (N_1046,N_842,N_647);
nand U1047 (N_1047,N_586,N_507);
xnor U1048 (N_1048,N_606,N_879);
nand U1049 (N_1049,N_241,N_172);
or U1050 (N_1050,N_938,N_775);
nor U1051 (N_1051,N_796,N_779);
nand U1052 (N_1052,N_467,N_370);
or U1053 (N_1053,N_947,N_392);
or U1054 (N_1054,N_846,N_851);
and U1055 (N_1055,N_304,N_840);
xnor U1056 (N_1056,N_218,N_780);
or U1057 (N_1057,N_990,N_585);
nand U1058 (N_1058,N_976,N_128);
nand U1059 (N_1059,N_288,N_833);
and U1060 (N_1060,N_113,N_354);
and U1061 (N_1061,N_388,N_255);
nand U1062 (N_1062,N_327,N_299);
xor U1063 (N_1063,N_335,N_893);
xor U1064 (N_1064,N_25,N_334);
nand U1065 (N_1065,N_810,N_249);
nand U1066 (N_1066,N_117,N_292);
xor U1067 (N_1067,N_326,N_0);
nor U1068 (N_1068,N_713,N_195);
or U1069 (N_1069,N_688,N_818);
xor U1070 (N_1070,N_864,N_669);
xor U1071 (N_1071,N_480,N_649);
nand U1072 (N_1072,N_791,N_341);
nor U1073 (N_1073,N_386,N_641);
nand U1074 (N_1074,N_419,N_268);
or U1075 (N_1075,N_34,N_704);
and U1076 (N_1076,N_170,N_22);
nand U1077 (N_1077,N_579,N_783);
nor U1078 (N_1078,N_638,N_156);
nand U1079 (N_1079,N_789,N_727);
or U1080 (N_1080,N_829,N_374);
nand U1081 (N_1081,N_84,N_375);
nand U1082 (N_1082,N_132,N_471);
nand U1083 (N_1083,N_705,N_321);
xnor U1084 (N_1084,N_886,N_513);
xor U1085 (N_1085,N_655,N_708);
and U1086 (N_1086,N_279,N_308);
or U1087 (N_1087,N_677,N_193);
or U1088 (N_1088,N_665,N_558);
and U1089 (N_1089,N_663,N_322);
nand U1090 (N_1090,N_591,N_532);
or U1091 (N_1091,N_964,N_541);
or U1092 (N_1092,N_732,N_739);
xor U1093 (N_1093,N_920,N_184);
nand U1094 (N_1094,N_456,N_97);
nor U1095 (N_1095,N_913,N_148);
or U1096 (N_1096,N_207,N_778);
nand U1097 (N_1097,N_762,N_616);
nor U1098 (N_1098,N_183,N_848);
nor U1099 (N_1099,N_144,N_896);
and U1100 (N_1100,N_626,N_409);
or U1101 (N_1101,N_131,N_765);
nor U1102 (N_1102,N_403,N_23);
nand U1103 (N_1103,N_212,N_125);
nor U1104 (N_1104,N_393,N_99);
nand U1105 (N_1105,N_668,N_475);
nand U1106 (N_1106,N_993,N_40);
xor U1107 (N_1107,N_58,N_366);
nand U1108 (N_1108,N_728,N_582);
xnor U1109 (N_1109,N_747,N_531);
nand U1110 (N_1110,N_596,N_952);
nand U1111 (N_1111,N_566,N_12);
nand U1112 (N_1112,N_970,N_229);
nand U1113 (N_1113,N_114,N_627);
or U1114 (N_1114,N_824,N_492);
nand U1115 (N_1115,N_464,N_973);
or U1116 (N_1116,N_547,N_645);
xnor U1117 (N_1117,N_908,N_194);
nor U1118 (N_1118,N_362,N_927);
xor U1119 (N_1119,N_903,N_790);
nand U1120 (N_1120,N_38,N_753);
nor U1121 (N_1121,N_935,N_383);
nor U1122 (N_1122,N_161,N_887);
nand U1123 (N_1123,N_43,N_368);
or U1124 (N_1124,N_118,N_455);
and U1125 (N_1125,N_280,N_127);
nor U1126 (N_1126,N_272,N_382);
and U1127 (N_1127,N_828,N_15);
and U1128 (N_1128,N_666,N_701);
nor U1129 (N_1129,N_244,N_770);
nand U1130 (N_1130,N_331,N_536);
or U1131 (N_1131,N_8,N_11);
or U1132 (N_1132,N_644,N_785);
and U1133 (N_1133,N_406,N_89);
or U1134 (N_1134,N_700,N_633);
nand U1135 (N_1135,N_216,N_683);
xor U1136 (N_1136,N_423,N_202);
and U1137 (N_1137,N_760,N_13);
xor U1138 (N_1138,N_781,N_847);
nand U1139 (N_1139,N_431,N_517);
xnor U1140 (N_1140,N_340,N_516);
nor U1141 (N_1141,N_235,N_265);
nand U1142 (N_1142,N_347,N_226);
xnor U1143 (N_1143,N_324,N_709);
or U1144 (N_1144,N_915,N_294);
nand U1145 (N_1145,N_634,N_188);
or U1146 (N_1146,N_41,N_629);
or U1147 (N_1147,N_469,N_950);
nor U1148 (N_1148,N_830,N_614);
and U1149 (N_1149,N_214,N_495);
nor U1150 (N_1150,N_693,N_673);
nor U1151 (N_1151,N_411,N_454);
nor U1152 (N_1152,N_929,N_519);
or U1153 (N_1153,N_948,N_731);
nand U1154 (N_1154,N_70,N_457);
or U1155 (N_1155,N_316,N_458);
xnor U1156 (N_1156,N_64,N_751);
nor U1157 (N_1157,N_399,N_160);
xnor U1158 (N_1158,N_92,N_329);
nor U1159 (N_1159,N_530,N_227);
nor U1160 (N_1160,N_504,N_422);
nor U1161 (N_1161,N_997,N_296);
nand U1162 (N_1162,N_391,N_544);
xor U1163 (N_1163,N_734,N_525);
and U1164 (N_1164,N_314,N_477);
nor U1165 (N_1165,N_877,N_3);
nand U1166 (N_1166,N_961,N_944);
nor U1167 (N_1167,N_744,N_396);
nand U1168 (N_1168,N_50,N_141);
or U1169 (N_1169,N_769,N_599);
and U1170 (N_1170,N_468,N_230);
xor U1171 (N_1171,N_130,N_278);
nand U1172 (N_1172,N_801,N_180);
and U1173 (N_1173,N_196,N_910);
nand U1174 (N_1174,N_169,N_563);
or U1175 (N_1175,N_35,N_812);
xnor U1176 (N_1176,N_206,N_256);
nand U1177 (N_1177,N_277,N_494);
and U1178 (N_1178,N_712,N_658);
and U1179 (N_1179,N_446,N_576);
or U1180 (N_1180,N_524,N_385);
xor U1181 (N_1181,N_679,N_592);
and U1182 (N_1182,N_860,N_900);
xor U1183 (N_1183,N_743,N_573);
nor U1184 (N_1184,N_146,N_250);
nor U1185 (N_1185,N_618,N_266);
xor U1186 (N_1186,N_756,N_398);
and U1187 (N_1187,N_898,N_612);
xnor U1188 (N_1188,N_807,N_290);
or U1189 (N_1189,N_597,N_858);
or U1190 (N_1190,N_215,N_254);
and U1191 (N_1191,N_293,N_574);
or U1192 (N_1192,N_307,N_737);
and U1193 (N_1193,N_914,N_186);
and U1194 (N_1194,N_577,N_433);
nand U1195 (N_1195,N_595,N_981);
nor U1196 (N_1196,N_103,N_557);
nand U1197 (N_1197,N_717,N_974);
xor U1198 (N_1198,N_906,N_345);
nand U1199 (N_1199,N_623,N_328);
xor U1200 (N_1200,N_901,N_302);
and U1201 (N_1201,N_449,N_916);
nand U1202 (N_1202,N_819,N_61);
nand U1203 (N_1203,N_539,N_689);
xnor U1204 (N_1204,N_814,N_723);
nor U1205 (N_1205,N_650,N_448);
nor U1206 (N_1206,N_417,N_359);
xor U1207 (N_1207,N_972,N_225);
or U1208 (N_1208,N_178,N_289);
nand U1209 (N_1209,N_9,N_687);
nand U1210 (N_1210,N_540,N_667);
nand U1211 (N_1211,N_440,N_622);
or U1212 (N_1212,N_190,N_551);
nand U1213 (N_1213,N_930,N_164);
or U1214 (N_1214,N_741,N_351);
nand U1215 (N_1215,N_333,N_960);
and U1216 (N_1216,N_95,N_619);
and U1217 (N_1217,N_14,N_588);
nand U1218 (N_1218,N_608,N_192);
nor U1219 (N_1219,N_472,N_301);
or U1220 (N_1220,N_742,N_309);
nand U1221 (N_1221,N_390,N_441);
nor U1222 (N_1222,N_337,N_660);
and U1223 (N_1223,N_855,N_859);
or U1224 (N_1224,N_208,N_415);
nor U1225 (N_1225,N_816,N_407);
nand U1226 (N_1226,N_527,N_210);
and U1227 (N_1227,N_834,N_421);
and U1228 (N_1228,N_940,N_711);
xnor U1229 (N_1229,N_284,N_691);
nand U1230 (N_1230,N_805,N_151);
nor U1231 (N_1231,N_890,N_124);
or U1232 (N_1232,N_26,N_643);
or U1233 (N_1233,N_714,N_832);
nor U1234 (N_1234,N_553,N_501);
or U1235 (N_1235,N_365,N_729);
nand U1236 (N_1236,N_260,N_159);
xnor U1237 (N_1237,N_698,N_923);
nor U1238 (N_1238,N_262,N_112);
or U1239 (N_1239,N_59,N_809);
and U1240 (N_1240,N_873,N_518);
nor U1241 (N_1241,N_107,N_907);
xor U1242 (N_1242,N_697,N_926);
nand U1243 (N_1243,N_122,N_686);
nor U1244 (N_1244,N_624,N_509);
xnor U1245 (N_1245,N_767,N_211);
nor U1246 (N_1246,N_648,N_33);
xnor U1247 (N_1247,N_490,N_7);
or U1248 (N_1248,N_54,N_123);
xor U1249 (N_1249,N_604,N_384);
or U1250 (N_1250,N_564,N_246);
and U1251 (N_1251,N_55,N_306);
and U1252 (N_1252,N_315,N_826);
xnor U1253 (N_1253,N_715,N_320);
and U1254 (N_1254,N_32,N_989);
or U1255 (N_1255,N_502,N_474);
xor U1256 (N_1256,N_94,N_888);
xor U1257 (N_1257,N_470,N_850);
and U1258 (N_1258,N_258,N_402);
and U1259 (N_1259,N_137,N_310);
and U1260 (N_1260,N_802,N_350);
nor U1261 (N_1261,N_962,N_201);
or U1262 (N_1262,N_31,N_672);
or U1263 (N_1263,N_759,N_499);
and U1264 (N_1264,N_542,N_722);
nor U1265 (N_1265,N_139,N_36);
nor U1266 (N_1266,N_636,N_323);
nand U1267 (N_1267,N_305,N_902);
xor U1268 (N_1268,N_533,N_162);
xor U1269 (N_1269,N_426,N_703);
xor U1270 (N_1270,N_228,N_465);
or U1271 (N_1271,N_546,N_27);
or U1272 (N_1272,N_149,N_854);
nand U1273 (N_1273,N_958,N_247);
or U1274 (N_1274,N_56,N_86);
nor U1275 (N_1275,N_827,N_605);
nor U1276 (N_1276,N_766,N_357);
or U1277 (N_1277,N_44,N_552);
or U1278 (N_1278,N_508,N_115);
and U1279 (N_1279,N_191,N_379);
xor U1280 (N_1280,N_79,N_252);
nand U1281 (N_1281,N_529,N_413);
nor U1282 (N_1282,N_332,N_57);
or U1283 (N_1283,N_919,N_108);
nand U1284 (N_1284,N_792,N_197);
nand U1285 (N_1285,N_657,N_707);
nor U1286 (N_1286,N_675,N_696);
and U1287 (N_1287,N_142,N_545);
nor U1288 (N_1288,N_269,N_806);
or U1289 (N_1289,N_414,N_364);
nor U1290 (N_1290,N_550,N_671);
xnor U1291 (N_1291,N_233,N_537);
and U1292 (N_1292,N_451,N_313);
or U1293 (N_1293,N_899,N_631);
and U1294 (N_1294,N_768,N_24);
and U1295 (N_1295,N_528,N_710);
and U1296 (N_1296,N_654,N_795);
and U1297 (N_1297,N_598,N_443);
nand U1298 (N_1298,N_87,N_680);
xnor U1299 (N_1299,N_764,N_664);
nand U1300 (N_1300,N_295,N_283);
nand U1301 (N_1301,N_953,N_782);
nand U1302 (N_1302,N_2,N_264);
or U1303 (N_1303,N_203,N_88);
or U1304 (N_1304,N_917,N_68);
nor U1305 (N_1305,N_240,N_602);
nor U1306 (N_1306,N_259,N_491);
nor U1307 (N_1307,N_861,N_483);
xor U1308 (N_1308,N_968,N_232);
xor U1309 (N_1309,N_836,N_346);
nor U1310 (N_1310,N_220,N_442);
or U1311 (N_1311,N_360,N_487);
nand U1312 (N_1312,N_733,N_438);
xnor U1313 (N_1313,N_841,N_884);
nand U1314 (N_1314,N_430,N_152);
or U1315 (N_1315,N_53,N_874);
nor U1316 (N_1316,N_213,N_548);
nand U1317 (N_1317,N_885,N_959);
or U1318 (N_1318,N_568,N_67);
or U1319 (N_1319,N_275,N_571);
and U1320 (N_1320,N_684,N_339);
or U1321 (N_1321,N_773,N_637);
or U1322 (N_1322,N_949,N_239);
nor U1323 (N_1323,N_6,N_772);
and U1324 (N_1324,N_205,N_460);
nor U1325 (N_1325,N_839,N_105);
and U1326 (N_1326,N_682,N_311);
xnor U1327 (N_1327,N_730,N_867);
nor U1328 (N_1328,N_217,N_168);
and U1329 (N_1329,N_376,N_567);
or U1330 (N_1330,N_825,N_410);
and U1331 (N_1331,N_63,N_857);
or U1332 (N_1332,N_758,N_788);
or U1333 (N_1333,N_261,N_676);
nand U1334 (N_1334,N_957,N_236);
or U1335 (N_1335,N_757,N_134);
or U1336 (N_1336,N_581,N_154);
nor U1337 (N_1337,N_909,N_478);
and U1338 (N_1338,N_843,N_752);
nor U1339 (N_1339,N_793,N_943);
nand U1340 (N_1340,N_291,N_808);
or U1341 (N_1341,N_356,N_821);
nand U1342 (N_1342,N_231,N_145);
nand U1343 (N_1343,N_569,N_209);
nand U1344 (N_1344,N_77,N_928);
xor U1345 (N_1345,N_147,N_750);
and U1346 (N_1346,N_511,N_175);
or U1347 (N_1347,N_78,N_803);
and U1348 (N_1348,N_640,N_405);
or U1349 (N_1349,N_999,N_982);
xnor U1350 (N_1350,N_219,N_82);
and U1351 (N_1351,N_786,N_746);
and U1352 (N_1352,N_83,N_387);
or U1353 (N_1353,N_187,N_65);
nor U1354 (N_1354,N_343,N_955);
nand U1355 (N_1355,N_995,N_367);
and U1356 (N_1356,N_447,N_91);
xor U1357 (N_1357,N_30,N_120);
xnor U1358 (N_1358,N_167,N_538);
nand U1359 (N_1359,N_589,N_221);
nor U1360 (N_1360,N_678,N_515);
or U1361 (N_1361,N_979,N_493);
or U1362 (N_1362,N_862,N_787);
or U1363 (N_1363,N_179,N_237);
nor U1364 (N_1364,N_936,N_361);
or U1365 (N_1365,N_941,N_694);
or U1366 (N_1366,N_939,N_876);
and U1367 (N_1367,N_942,N_954);
or U1368 (N_1368,N_355,N_583);
or U1369 (N_1369,N_580,N_865);
nor U1370 (N_1370,N_224,N_462);
xnor U1371 (N_1371,N_690,N_565);
and U1372 (N_1372,N_844,N_601);
or U1373 (N_1373,N_659,N_459);
or U1374 (N_1374,N_348,N_755);
nand U1375 (N_1375,N_967,N_389);
nand U1376 (N_1376,N_52,N_845);
and U1377 (N_1377,N_912,N_924);
and U1378 (N_1378,N_661,N_412);
nor U1379 (N_1379,N_875,N_121);
xnor U1380 (N_1380,N_75,N_318);
and U1381 (N_1381,N_984,N_133);
nor U1382 (N_1382,N_281,N_401);
nor U1383 (N_1383,N_804,N_575);
or U1384 (N_1384,N_549,N_774);
nor U1385 (N_1385,N_76,N_287);
xnor U1386 (N_1386,N_408,N_481);
nor U1387 (N_1387,N_646,N_892);
xor U1388 (N_1388,N_986,N_607);
nand U1389 (N_1389,N_344,N_49);
or U1390 (N_1390,N_439,N_883);
nand U1391 (N_1391,N_90,N_234);
nand U1392 (N_1392,N_37,N_496);
nand U1393 (N_1393,N_523,N_937);
xnor U1394 (N_1394,N_140,N_933);
xnor U1395 (N_1395,N_444,N_270);
and U1396 (N_1396,N_543,N_500);
xor U1397 (N_1397,N_110,N_158);
nor U1398 (N_1398,N_404,N_81);
nor U1399 (N_1399,N_777,N_838);
nor U1400 (N_1400,N_482,N_587);
and U1401 (N_1401,N_719,N_966);
or U1402 (N_1402,N_611,N_748);
and U1403 (N_1403,N_223,N_116);
nand U1404 (N_1404,N_62,N_51);
and U1405 (N_1405,N_570,N_424);
nor U1406 (N_1406,N_945,N_794);
nand U1407 (N_1407,N_975,N_138);
xor U1408 (N_1408,N_400,N_200);
nand U1409 (N_1409,N_285,N_473);
xnor U1410 (N_1410,N_248,N_798);
nand U1411 (N_1411,N_951,N_994);
xor U1412 (N_1412,N_815,N_852);
or U1413 (N_1413,N_102,N_615);
and U1414 (N_1414,N_416,N_85);
nand U1415 (N_1415,N_559,N_776);
nand U1416 (N_1416,N_681,N_692);
nand U1417 (N_1417,N_222,N_380);
nor U1418 (N_1418,N_977,N_613);
and U1419 (N_1419,N_889,N_963);
nand U1420 (N_1420,N_749,N_635);
or U1421 (N_1421,N_872,N_505);
nor U1422 (N_1422,N_897,N_176);
and U1423 (N_1423,N_267,N_642);
nor U1424 (N_1424,N_521,N_822);
nor U1425 (N_1425,N_96,N_274);
or U1426 (N_1426,N_485,N_479);
and U1427 (N_1427,N_556,N_560);
nand U1428 (N_1428,N_48,N_395);
and U1429 (N_1429,N_863,N_831);
or U1430 (N_1430,N_498,N_978);
and U1431 (N_1431,N_39,N_811);
xor U1432 (N_1432,N_870,N_298);
nand U1433 (N_1433,N_101,N_514);
and U1434 (N_1434,N_319,N_72);
and U1435 (N_1435,N_987,N_800);
or U1436 (N_1436,N_998,N_245);
nor U1437 (N_1437,N_166,N_297);
and U1438 (N_1438,N_373,N_522);
or U1439 (N_1439,N_726,N_198);
nor U1440 (N_1440,N_971,N_16);
nand U1441 (N_1441,N_312,N_126);
nor U1442 (N_1442,N_182,N_965);
nor U1443 (N_1443,N_18,N_452);
nand U1444 (N_1444,N_835,N_19);
and U1445 (N_1445,N_820,N_429);
xor U1446 (N_1446,N_325,N_881);
and U1447 (N_1447,N_656,N_931);
nor U1448 (N_1448,N_489,N_303);
and U1449 (N_1449,N_621,N_369);
nand U1450 (N_1450,N_721,N_895);
nor U1451 (N_1451,N_702,N_461);
nor U1452 (N_1452,N_632,N_620);
xnor U1453 (N_1453,N_784,N_435);
or U1454 (N_1454,N_111,N_243);
nand U1455 (N_1455,N_372,N_397);
xnor U1456 (N_1456,N_745,N_136);
and U1457 (N_1457,N_662,N_135);
xor U1458 (N_1458,N_823,N_276);
nor U1459 (N_1459,N_317,N_738);
or U1460 (N_1460,N_300,N_946);
nand U1461 (N_1461,N_358,N_630);
nor U1462 (N_1462,N_177,N_436);
xnor U1463 (N_1463,N_371,N_590);
nor U1464 (N_1464,N_282,N_871);
and U1465 (N_1465,N_204,N_628);
and U1466 (N_1466,N_868,N_670);
xor U1467 (N_1467,N_520,N_418);
nor U1468 (N_1468,N_797,N_150);
nor U1469 (N_1469,N_578,N_173);
or U1470 (N_1470,N_882,N_71);
xor U1471 (N_1471,N_352,N_434);
and U1472 (N_1472,N_817,N_185);
and U1473 (N_1473,N_724,N_554);
nand U1474 (N_1474,N_4,N_157);
xor U1475 (N_1475,N_853,N_425);
or U1476 (N_1476,N_98,N_238);
nor U1477 (N_1477,N_29,N_463);
or U1478 (N_1478,N_996,N_453);
nand U1479 (N_1479,N_512,N_918);
nand U1480 (N_1480,N_651,N_988);
or U1481 (N_1481,N_189,N_837);
or U1482 (N_1482,N_561,N_21);
xor U1483 (N_1483,N_880,N_925);
nor U1484 (N_1484,N_349,N_652);
nand U1485 (N_1485,N_740,N_763);
and U1486 (N_1486,N_484,N_263);
nand U1487 (N_1487,N_381,N_956);
or U1488 (N_1488,N_535,N_625);
nand U1489 (N_1489,N_353,N_921);
nand U1490 (N_1490,N_716,N_42);
or U1491 (N_1491,N_20,N_428);
or U1492 (N_1492,N_251,N_674);
xnor U1493 (N_1493,N_718,N_377);
and U1494 (N_1494,N_74,N_706);
or U1495 (N_1495,N_526,N_253);
or U1496 (N_1496,N_1,N_45);
and U1497 (N_1497,N_432,N_922);
xnor U1498 (N_1498,N_80,N_856);
and U1499 (N_1499,N_273,N_476);
nor U1500 (N_1500,N_166,N_936);
xnor U1501 (N_1501,N_758,N_879);
xor U1502 (N_1502,N_498,N_746);
or U1503 (N_1503,N_49,N_476);
nand U1504 (N_1504,N_24,N_692);
nor U1505 (N_1505,N_506,N_644);
and U1506 (N_1506,N_345,N_929);
or U1507 (N_1507,N_61,N_244);
xor U1508 (N_1508,N_315,N_716);
nand U1509 (N_1509,N_839,N_470);
nand U1510 (N_1510,N_875,N_260);
nand U1511 (N_1511,N_460,N_514);
and U1512 (N_1512,N_343,N_900);
or U1513 (N_1513,N_34,N_94);
nor U1514 (N_1514,N_569,N_996);
nor U1515 (N_1515,N_529,N_583);
nor U1516 (N_1516,N_711,N_94);
nor U1517 (N_1517,N_179,N_519);
xnor U1518 (N_1518,N_783,N_716);
nand U1519 (N_1519,N_93,N_41);
xnor U1520 (N_1520,N_403,N_196);
xor U1521 (N_1521,N_446,N_602);
or U1522 (N_1522,N_711,N_417);
or U1523 (N_1523,N_56,N_238);
or U1524 (N_1524,N_160,N_438);
or U1525 (N_1525,N_362,N_433);
or U1526 (N_1526,N_669,N_416);
and U1527 (N_1527,N_483,N_218);
nor U1528 (N_1528,N_436,N_248);
nor U1529 (N_1529,N_521,N_263);
nand U1530 (N_1530,N_793,N_762);
nand U1531 (N_1531,N_341,N_141);
xnor U1532 (N_1532,N_323,N_9);
xnor U1533 (N_1533,N_178,N_978);
nor U1534 (N_1534,N_432,N_251);
and U1535 (N_1535,N_391,N_496);
and U1536 (N_1536,N_752,N_306);
nor U1537 (N_1537,N_778,N_219);
or U1538 (N_1538,N_0,N_737);
nor U1539 (N_1539,N_759,N_619);
nor U1540 (N_1540,N_203,N_232);
nand U1541 (N_1541,N_122,N_824);
and U1542 (N_1542,N_887,N_465);
nand U1543 (N_1543,N_752,N_893);
and U1544 (N_1544,N_902,N_705);
or U1545 (N_1545,N_388,N_632);
nor U1546 (N_1546,N_541,N_336);
or U1547 (N_1547,N_493,N_457);
nor U1548 (N_1548,N_600,N_960);
and U1549 (N_1549,N_289,N_961);
xor U1550 (N_1550,N_390,N_766);
and U1551 (N_1551,N_215,N_134);
and U1552 (N_1552,N_847,N_928);
nand U1553 (N_1553,N_725,N_280);
nand U1554 (N_1554,N_171,N_591);
nor U1555 (N_1555,N_408,N_643);
nand U1556 (N_1556,N_400,N_202);
nor U1557 (N_1557,N_832,N_851);
nand U1558 (N_1558,N_397,N_91);
or U1559 (N_1559,N_387,N_42);
nand U1560 (N_1560,N_472,N_924);
and U1561 (N_1561,N_283,N_806);
xnor U1562 (N_1562,N_845,N_588);
nor U1563 (N_1563,N_596,N_693);
and U1564 (N_1564,N_703,N_462);
xnor U1565 (N_1565,N_421,N_630);
or U1566 (N_1566,N_6,N_442);
and U1567 (N_1567,N_652,N_79);
nor U1568 (N_1568,N_349,N_330);
xor U1569 (N_1569,N_475,N_539);
nor U1570 (N_1570,N_580,N_324);
and U1571 (N_1571,N_896,N_124);
and U1572 (N_1572,N_818,N_527);
and U1573 (N_1573,N_901,N_830);
nor U1574 (N_1574,N_390,N_255);
and U1575 (N_1575,N_735,N_175);
nor U1576 (N_1576,N_915,N_134);
nand U1577 (N_1577,N_307,N_7);
nand U1578 (N_1578,N_874,N_931);
nand U1579 (N_1579,N_723,N_782);
and U1580 (N_1580,N_280,N_739);
or U1581 (N_1581,N_231,N_470);
nand U1582 (N_1582,N_49,N_537);
xor U1583 (N_1583,N_610,N_663);
or U1584 (N_1584,N_331,N_348);
nor U1585 (N_1585,N_636,N_503);
or U1586 (N_1586,N_834,N_671);
nand U1587 (N_1587,N_310,N_660);
xnor U1588 (N_1588,N_242,N_902);
nor U1589 (N_1589,N_230,N_119);
xnor U1590 (N_1590,N_657,N_487);
nor U1591 (N_1591,N_188,N_639);
nor U1592 (N_1592,N_69,N_674);
xnor U1593 (N_1593,N_308,N_921);
xor U1594 (N_1594,N_731,N_905);
and U1595 (N_1595,N_327,N_890);
or U1596 (N_1596,N_422,N_391);
nor U1597 (N_1597,N_984,N_224);
and U1598 (N_1598,N_701,N_842);
nor U1599 (N_1599,N_693,N_644);
xnor U1600 (N_1600,N_286,N_671);
xnor U1601 (N_1601,N_587,N_608);
xnor U1602 (N_1602,N_670,N_477);
nor U1603 (N_1603,N_453,N_488);
or U1604 (N_1604,N_374,N_991);
xnor U1605 (N_1605,N_948,N_914);
nand U1606 (N_1606,N_88,N_826);
and U1607 (N_1607,N_113,N_715);
xor U1608 (N_1608,N_748,N_198);
nor U1609 (N_1609,N_707,N_482);
xor U1610 (N_1610,N_293,N_416);
nor U1611 (N_1611,N_800,N_957);
xnor U1612 (N_1612,N_90,N_811);
nor U1613 (N_1613,N_997,N_712);
nor U1614 (N_1614,N_721,N_880);
nor U1615 (N_1615,N_327,N_610);
or U1616 (N_1616,N_55,N_810);
nand U1617 (N_1617,N_690,N_554);
xnor U1618 (N_1618,N_593,N_943);
nor U1619 (N_1619,N_334,N_348);
and U1620 (N_1620,N_105,N_171);
nand U1621 (N_1621,N_326,N_199);
or U1622 (N_1622,N_601,N_290);
nand U1623 (N_1623,N_558,N_981);
and U1624 (N_1624,N_551,N_125);
and U1625 (N_1625,N_895,N_442);
and U1626 (N_1626,N_257,N_216);
nor U1627 (N_1627,N_127,N_986);
and U1628 (N_1628,N_72,N_142);
nor U1629 (N_1629,N_421,N_149);
nor U1630 (N_1630,N_710,N_651);
nand U1631 (N_1631,N_793,N_416);
or U1632 (N_1632,N_28,N_569);
nor U1633 (N_1633,N_178,N_59);
nor U1634 (N_1634,N_163,N_816);
nor U1635 (N_1635,N_175,N_476);
and U1636 (N_1636,N_964,N_547);
nand U1637 (N_1637,N_193,N_327);
or U1638 (N_1638,N_896,N_718);
nor U1639 (N_1639,N_780,N_956);
xor U1640 (N_1640,N_447,N_742);
xor U1641 (N_1641,N_288,N_952);
or U1642 (N_1642,N_660,N_775);
nand U1643 (N_1643,N_660,N_101);
nand U1644 (N_1644,N_312,N_681);
and U1645 (N_1645,N_408,N_550);
xor U1646 (N_1646,N_825,N_497);
and U1647 (N_1647,N_233,N_169);
and U1648 (N_1648,N_640,N_720);
xor U1649 (N_1649,N_882,N_874);
and U1650 (N_1650,N_760,N_226);
nor U1651 (N_1651,N_441,N_603);
nand U1652 (N_1652,N_967,N_419);
xor U1653 (N_1653,N_190,N_572);
nand U1654 (N_1654,N_406,N_241);
or U1655 (N_1655,N_205,N_990);
xnor U1656 (N_1656,N_895,N_36);
or U1657 (N_1657,N_7,N_825);
xnor U1658 (N_1658,N_68,N_381);
xnor U1659 (N_1659,N_714,N_964);
and U1660 (N_1660,N_449,N_922);
nor U1661 (N_1661,N_473,N_45);
nand U1662 (N_1662,N_624,N_584);
and U1663 (N_1663,N_326,N_751);
and U1664 (N_1664,N_686,N_387);
nand U1665 (N_1665,N_23,N_312);
and U1666 (N_1666,N_779,N_945);
nor U1667 (N_1667,N_86,N_614);
nand U1668 (N_1668,N_730,N_808);
nor U1669 (N_1669,N_537,N_744);
or U1670 (N_1670,N_806,N_183);
or U1671 (N_1671,N_675,N_874);
or U1672 (N_1672,N_45,N_533);
nand U1673 (N_1673,N_915,N_95);
nand U1674 (N_1674,N_542,N_664);
nor U1675 (N_1675,N_730,N_624);
nor U1676 (N_1676,N_103,N_54);
or U1677 (N_1677,N_326,N_49);
nor U1678 (N_1678,N_858,N_333);
or U1679 (N_1679,N_762,N_355);
nor U1680 (N_1680,N_303,N_702);
xor U1681 (N_1681,N_979,N_369);
and U1682 (N_1682,N_389,N_714);
nand U1683 (N_1683,N_480,N_489);
nor U1684 (N_1684,N_66,N_591);
and U1685 (N_1685,N_251,N_721);
nand U1686 (N_1686,N_711,N_523);
nor U1687 (N_1687,N_804,N_951);
xor U1688 (N_1688,N_240,N_805);
nand U1689 (N_1689,N_648,N_780);
or U1690 (N_1690,N_86,N_28);
and U1691 (N_1691,N_246,N_266);
or U1692 (N_1692,N_825,N_41);
nand U1693 (N_1693,N_674,N_370);
xor U1694 (N_1694,N_421,N_769);
xor U1695 (N_1695,N_825,N_137);
or U1696 (N_1696,N_295,N_89);
nor U1697 (N_1697,N_219,N_603);
nor U1698 (N_1698,N_748,N_801);
or U1699 (N_1699,N_413,N_517);
and U1700 (N_1700,N_59,N_18);
xor U1701 (N_1701,N_984,N_678);
or U1702 (N_1702,N_100,N_201);
nand U1703 (N_1703,N_782,N_392);
xor U1704 (N_1704,N_95,N_110);
nand U1705 (N_1705,N_962,N_233);
and U1706 (N_1706,N_714,N_466);
xor U1707 (N_1707,N_859,N_37);
and U1708 (N_1708,N_991,N_64);
nand U1709 (N_1709,N_275,N_613);
nor U1710 (N_1710,N_194,N_961);
or U1711 (N_1711,N_412,N_721);
and U1712 (N_1712,N_283,N_603);
xnor U1713 (N_1713,N_661,N_385);
nand U1714 (N_1714,N_340,N_346);
and U1715 (N_1715,N_203,N_496);
nand U1716 (N_1716,N_893,N_622);
nor U1717 (N_1717,N_295,N_244);
nand U1718 (N_1718,N_114,N_949);
and U1719 (N_1719,N_246,N_960);
or U1720 (N_1720,N_15,N_120);
and U1721 (N_1721,N_148,N_549);
and U1722 (N_1722,N_267,N_406);
nand U1723 (N_1723,N_953,N_25);
xor U1724 (N_1724,N_167,N_240);
xnor U1725 (N_1725,N_301,N_522);
nand U1726 (N_1726,N_197,N_480);
and U1727 (N_1727,N_990,N_394);
nand U1728 (N_1728,N_164,N_261);
nor U1729 (N_1729,N_385,N_5);
xnor U1730 (N_1730,N_984,N_860);
and U1731 (N_1731,N_822,N_652);
or U1732 (N_1732,N_451,N_463);
or U1733 (N_1733,N_772,N_673);
xor U1734 (N_1734,N_277,N_899);
xnor U1735 (N_1735,N_618,N_653);
xnor U1736 (N_1736,N_318,N_634);
xnor U1737 (N_1737,N_428,N_257);
nand U1738 (N_1738,N_652,N_76);
and U1739 (N_1739,N_220,N_130);
nand U1740 (N_1740,N_517,N_399);
or U1741 (N_1741,N_950,N_929);
nor U1742 (N_1742,N_779,N_278);
xor U1743 (N_1743,N_420,N_624);
or U1744 (N_1744,N_424,N_467);
nor U1745 (N_1745,N_484,N_195);
xnor U1746 (N_1746,N_721,N_369);
or U1747 (N_1747,N_327,N_695);
or U1748 (N_1748,N_995,N_141);
nor U1749 (N_1749,N_784,N_550);
xnor U1750 (N_1750,N_156,N_93);
xnor U1751 (N_1751,N_331,N_472);
or U1752 (N_1752,N_420,N_683);
xor U1753 (N_1753,N_122,N_918);
nand U1754 (N_1754,N_496,N_232);
nor U1755 (N_1755,N_84,N_831);
xnor U1756 (N_1756,N_35,N_882);
nand U1757 (N_1757,N_225,N_676);
nand U1758 (N_1758,N_546,N_463);
xor U1759 (N_1759,N_159,N_392);
and U1760 (N_1760,N_601,N_207);
and U1761 (N_1761,N_777,N_752);
xor U1762 (N_1762,N_728,N_497);
xor U1763 (N_1763,N_531,N_666);
and U1764 (N_1764,N_136,N_342);
nand U1765 (N_1765,N_569,N_938);
nor U1766 (N_1766,N_584,N_26);
nor U1767 (N_1767,N_241,N_622);
nor U1768 (N_1768,N_319,N_454);
xnor U1769 (N_1769,N_387,N_427);
and U1770 (N_1770,N_532,N_337);
or U1771 (N_1771,N_951,N_613);
or U1772 (N_1772,N_629,N_631);
and U1773 (N_1773,N_784,N_199);
xnor U1774 (N_1774,N_745,N_332);
nor U1775 (N_1775,N_559,N_274);
and U1776 (N_1776,N_26,N_335);
nor U1777 (N_1777,N_630,N_407);
or U1778 (N_1778,N_669,N_356);
or U1779 (N_1779,N_35,N_599);
and U1780 (N_1780,N_36,N_988);
xor U1781 (N_1781,N_696,N_718);
nand U1782 (N_1782,N_813,N_456);
nand U1783 (N_1783,N_444,N_874);
nand U1784 (N_1784,N_976,N_791);
nor U1785 (N_1785,N_323,N_92);
and U1786 (N_1786,N_69,N_421);
xnor U1787 (N_1787,N_393,N_103);
xor U1788 (N_1788,N_398,N_230);
xor U1789 (N_1789,N_252,N_479);
or U1790 (N_1790,N_967,N_100);
and U1791 (N_1791,N_124,N_948);
xor U1792 (N_1792,N_624,N_936);
and U1793 (N_1793,N_220,N_86);
and U1794 (N_1794,N_766,N_340);
or U1795 (N_1795,N_364,N_178);
or U1796 (N_1796,N_859,N_811);
nand U1797 (N_1797,N_373,N_268);
and U1798 (N_1798,N_58,N_136);
or U1799 (N_1799,N_157,N_741);
nand U1800 (N_1800,N_236,N_99);
nand U1801 (N_1801,N_815,N_867);
xnor U1802 (N_1802,N_194,N_358);
or U1803 (N_1803,N_570,N_181);
xor U1804 (N_1804,N_376,N_692);
or U1805 (N_1805,N_804,N_306);
xnor U1806 (N_1806,N_895,N_777);
nand U1807 (N_1807,N_293,N_746);
and U1808 (N_1808,N_365,N_734);
xor U1809 (N_1809,N_422,N_3);
xor U1810 (N_1810,N_420,N_697);
nand U1811 (N_1811,N_694,N_625);
xor U1812 (N_1812,N_24,N_953);
nor U1813 (N_1813,N_654,N_949);
or U1814 (N_1814,N_64,N_150);
nor U1815 (N_1815,N_889,N_498);
nand U1816 (N_1816,N_559,N_327);
xor U1817 (N_1817,N_638,N_164);
nor U1818 (N_1818,N_182,N_354);
nor U1819 (N_1819,N_511,N_878);
or U1820 (N_1820,N_947,N_888);
nand U1821 (N_1821,N_35,N_937);
nor U1822 (N_1822,N_326,N_650);
nand U1823 (N_1823,N_143,N_587);
nor U1824 (N_1824,N_657,N_936);
nand U1825 (N_1825,N_793,N_692);
nor U1826 (N_1826,N_837,N_341);
nor U1827 (N_1827,N_423,N_218);
nand U1828 (N_1828,N_614,N_867);
nand U1829 (N_1829,N_573,N_504);
or U1830 (N_1830,N_199,N_198);
nor U1831 (N_1831,N_421,N_401);
or U1832 (N_1832,N_115,N_798);
xor U1833 (N_1833,N_201,N_157);
or U1834 (N_1834,N_67,N_420);
nor U1835 (N_1835,N_612,N_440);
or U1836 (N_1836,N_16,N_686);
nor U1837 (N_1837,N_687,N_466);
nor U1838 (N_1838,N_58,N_503);
xnor U1839 (N_1839,N_969,N_681);
xor U1840 (N_1840,N_333,N_417);
and U1841 (N_1841,N_225,N_887);
or U1842 (N_1842,N_610,N_24);
nand U1843 (N_1843,N_383,N_162);
nand U1844 (N_1844,N_750,N_508);
and U1845 (N_1845,N_321,N_188);
and U1846 (N_1846,N_613,N_17);
nand U1847 (N_1847,N_350,N_77);
nand U1848 (N_1848,N_330,N_77);
nand U1849 (N_1849,N_731,N_529);
or U1850 (N_1850,N_579,N_843);
nand U1851 (N_1851,N_269,N_765);
xor U1852 (N_1852,N_254,N_37);
and U1853 (N_1853,N_187,N_310);
nor U1854 (N_1854,N_508,N_298);
xor U1855 (N_1855,N_756,N_629);
xnor U1856 (N_1856,N_468,N_921);
nor U1857 (N_1857,N_546,N_986);
xnor U1858 (N_1858,N_879,N_461);
nand U1859 (N_1859,N_530,N_615);
or U1860 (N_1860,N_38,N_608);
nor U1861 (N_1861,N_578,N_451);
nor U1862 (N_1862,N_322,N_124);
xor U1863 (N_1863,N_925,N_643);
or U1864 (N_1864,N_621,N_109);
nand U1865 (N_1865,N_803,N_881);
or U1866 (N_1866,N_415,N_482);
or U1867 (N_1867,N_134,N_673);
or U1868 (N_1868,N_468,N_806);
nand U1869 (N_1869,N_824,N_774);
nand U1870 (N_1870,N_477,N_927);
xor U1871 (N_1871,N_882,N_481);
and U1872 (N_1872,N_236,N_469);
or U1873 (N_1873,N_764,N_731);
nand U1874 (N_1874,N_372,N_539);
nand U1875 (N_1875,N_568,N_225);
or U1876 (N_1876,N_428,N_70);
nand U1877 (N_1877,N_464,N_497);
xor U1878 (N_1878,N_802,N_20);
or U1879 (N_1879,N_870,N_928);
nor U1880 (N_1880,N_791,N_740);
or U1881 (N_1881,N_507,N_707);
nor U1882 (N_1882,N_167,N_7);
nand U1883 (N_1883,N_386,N_694);
xor U1884 (N_1884,N_205,N_891);
nand U1885 (N_1885,N_231,N_107);
or U1886 (N_1886,N_63,N_550);
nor U1887 (N_1887,N_0,N_250);
and U1888 (N_1888,N_662,N_255);
nor U1889 (N_1889,N_588,N_907);
or U1890 (N_1890,N_122,N_272);
and U1891 (N_1891,N_457,N_299);
nor U1892 (N_1892,N_12,N_756);
xnor U1893 (N_1893,N_199,N_566);
or U1894 (N_1894,N_340,N_211);
nor U1895 (N_1895,N_590,N_608);
or U1896 (N_1896,N_481,N_83);
nand U1897 (N_1897,N_132,N_245);
xnor U1898 (N_1898,N_516,N_645);
xor U1899 (N_1899,N_810,N_310);
nor U1900 (N_1900,N_469,N_619);
or U1901 (N_1901,N_306,N_853);
and U1902 (N_1902,N_55,N_491);
nand U1903 (N_1903,N_897,N_618);
nor U1904 (N_1904,N_192,N_810);
nor U1905 (N_1905,N_309,N_389);
nor U1906 (N_1906,N_487,N_932);
and U1907 (N_1907,N_721,N_390);
nor U1908 (N_1908,N_261,N_199);
nand U1909 (N_1909,N_937,N_586);
xnor U1910 (N_1910,N_135,N_246);
nand U1911 (N_1911,N_520,N_111);
or U1912 (N_1912,N_916,N_485);
nor U1913 (N_1913,N_112,N_982);
nand U1914 (N_1914,N_438,N_802);
nor U1915 (N_1915,N_790,N_463);
and U1916 (N_1916,N_89,N_671);
or U1917 (N_1917,N_60,N_963);
or U1918 (N_1918,N_358,N_770);
nor U1919 (N_1919,N_754,N_541);
and U1920 (N_1920,N_402,N_361);
nand U1921 (N_1921,N_682,N_472);
and U1922 (N_1922,N_813,N_675);
nor U1923 (N_1923,N_137,N_761);
or U1924 (N_1924,N_515,N_546);
nor U1925 (N_1925,N_212,N_691);
nand U1926 (N_1926,N_625,N_166);
xnor U1927 (N_1927,N_269,N_224);
and U1928 (N_1928,N_375,N_945);
or U1929 (N_1929,N_911,N_587);
and U1930 (N_1930,N_98,N_856);
or U1931 (N_1931,N_375,N_885);
nor U1932 (N_1932,N_167,N_459);
and U1933 (N_1933,N_483,N_498);
or U1934 (N_1934,N_993,N_849);
or U1935 (N_1935,N_660,N_461);
or U1936 (N_1936,N_577,N_323);
nand U1937 (N_1937,N_312,N_905);
xnor U1938 (N_1938,N_791,N_664);
nor U1939 (N_1939,N_504,N_347);
nor U1940 (N_1940,N_101,N_419);
nor U1941 (N_1941,N_451,N_699);
xor U1942 (N_1942,N_792,N_304);
and U1943 (N_1943,N_690,N_143);
nor U1944 (N_1944,N_1,N_943);
nand U1945 (N_1945,N_193,N_968);
xor U1946 (N_1946,N_987,N_442);
nand U1947 (N_1947,N_955,N_268);
nor U1948 (N_1948,N_504,N_556);
or U1949 (N_1949,N_711,N_622);
nand U1950 (N_1950,N_86,N_635);
or U1951 (N_1951,N_623,N_552);
and U1952 (N_1952,N_205,N_612);
nor U1953 (N_1953,N_885,N_948);
xor U1954 (N_1954,N_918,N_941);
nor U1955 (N_1955,N_698,N_904);
nor U1956 (N_1956,N_717,N_779);
nor U1957 (N_1957,N_23,N_831);
nor U1958 (N_1958,N_839,N_315);
and U1959 (N_1959,N_138,N_886);
xnor U1960 (N_1960,N_904,N_712);
xnor U1961 (N_1961,N_521,N_626);
xnor U1962 (N_1962,N_116,N_291);
xor U1963 (N_1963,N_535,N_144);
nor U1964 (N_1964,N_974,N_311);
nor U1965 (N_1965,N_869,N_290);
and U1966 (N_1966,N_577,N_436);
nand U1967 (N_1967,N_688,N_677);
and U1968 (N_1968,N_331,N_993);
nor U1969 (N_1969,N_839,N_535);
xnor U1970 (N_1970,N_832,N_889);
nor U1971 (N_1971,N_374,N_200);
nand U1972 (N_1972,N_168,N_88);
and U1973 (N_1973,N_879,N_560);
nand U1974 (N_1974,N_820,N_13);
and U1975 (N_1975,N_3,N_754);
xor U1976 (N_1976,N_302,N_598);
nand U1977 (N_1977,N_480,N_226);
xor U1978 (N_1978,N_941,N_997);
xnor U1979 (N_1979,N_65,N_323);
nand U1980 (N_1980,N_582,N_593);
xor U1981 (N_1981,N_722,N_424);
and U1982 (N_1982,N_389,N_699);
xor U1983 (N_1983,N_230,N_72);
nand U1984 (N_1984,N_160,N_347);
or U1985 (N_1985,N_98,N_225);
nand U1986 (N_1986,N_548,N_209);
nand U1987 (N_1987,N_941,N_176);
nor U1988 (N_1988,N_523,N_264);
and U1989 (N_1989,N_958,N_743);
xor U1990 (N_1990,N_411,N_147);
nand U1991 (N_1991,N_343,N_546);
nand U1992 (N_1992,N_499,N_454);
or U1993 (N_1993,N_150,N_172);
nand U1994 (N_1994,N_228,N_11);
nand U1995 (N_1995,N_79,N_133);
nor U1996 (N_1996,N_920,N_166);
xnor U1997 (N_1997,N_834,N_329);
or U1998 (N_1998,N_93,N_772);
xnor U1999 (N_1999,N_218,N_575);
and U2000 (N_2000,N_1297,N_1768);
and U2001 (N_2001,N_1595,N_1034);
or U2002 (N_2002,N_1889,N_1948);
or U2003 (N_2003,N_1617,N_1782);
nor U2004 (N_2004,N_1578,N_1284);
and U2005 (N_2005,N_1438,N_1465);
or U2006 (N_2006,N_1745,N_1681);
or U2007 (N_2007,N_1237,N_1611);
nand U2008 (N_2008,N_1463,N_1885);
or U2009 (N_2009,N_1644,N_1091);
xor U2010 (N_2010,N_1675,N_1957);
nor U2011 (N_2011,N_1328,N_1335);
nor U2012 (N_2012,N_1464,N_1175);
xnor U2013 (N_2013,N_1567,N_1994);
and U2014 (N_2014,N_1615,N_1873);
or U2015 (N_2015,N_1662,N_1254);
nor U2016 (N_2016,N_1743,N_1565);
nor U2017 (N_2017,N_1120,N_1862);
xnor U2018 (N_2018,N_1387,N_1532);
and U2019 (N_2019,N_1445,N_1262);
xnor U2020 (N_2020,N_1779,N_1864);
and U2021 (N_2021,N_1434,N_1521);
or U2022 (N_2022,N_1389,N_1668);
nor U2023 (N_2023,N_1986,N_1150);
and U2024 (N_2024,N_1451,N_1588);
and U2025 (N_2025,N_1226,N_1934);
nor U2026 (N_2026,N_1817,N_1966);
xnor U2027 (N_2027,N_1173,N_1100);
nor U2028 (N_2028,N_1345,N_1059);
nor U2029 (N_2029,N_1677,N_1625);
nand U2030 (N_2030,N_1912,N_1846);
nand U2031 (N_2031,N_1718,N_1001);
nand U2032 (N_2032,N_1334,N_1865);
nand U2033 (N_2033,N_1703,N_1461);
xor U2034 (N_2034,N_1241,N_1312);
xor U2035 (N_2035,N_1198,N_1057);
or U2036 (N_2036,N_1996,N_1601);
xor U2037 (N_2037,N_1468,N_1989);
or U2038 (N_2038,N_1716,N_1272);
or U2039 (N_2039,N_1110,N_1933);
xor U2040 (N_2040,N_1800,N_1375);
nand U2041 (N_2041,N_1596,N_1115);
xor U2042 (N_2042,N_1095,N_1991);
nor U2043 (N_2043,N_1992,N_1256);
or U2044 (N_2044,N_1664,N_1545);
nor U2045 (N_2045,N_1103,N_1574);
nand U2046 (N_2046,N_1659,N_1166);
and U2047 (N_2047,N_1831,N_1376);
and U2048 (N_2048,N_1024,N_1361);
nor U2049 (N_2049,N_1520,N_1340);
xor U2050 (N_2050,N_1436,N_1242);
nand U2051 (N_2051,N_1357,N_1697);
xnor U2052 (N_2052,N_1177,N_1943);
or U2053 (N_2053,N_1193,N_1129);
nor U2054 (N_2054,N_1495,N_1932);
or U2055 (N_2055,N_1493,N_1701);
xnor U2056 (N_2056,N_1552,N_1987);
nor U2057 (N_2057,N_1896,N_1229);
xor U2058 (N_2058,N_1645,N_1750);
or U2059 (N_2059,N_1952,N_1211);
nand U2060 (N_2060,N_1190,N_1268);
nand U2061 (N_2061,N_1043,N_1795);
and U2062 (N_2062,N_1674,N_1431);
xnor U2063 (N_2063,N_1618,N_1378);
nor U2064 (N_2064,N_1756,N_1806);
and U2065 (N_2065,N_1698,N_1594);
nand U2066 (N_2066,N_1672,N_1926);
nand U2067 (N_2067,N_1972,N_1012);
xnor U2068 (N_2068,N_1801,N_1196);
or U2069 (N_2069,N_1397,N_1139);
or U2070 (N_2070,N_1614,N_1822);
xnor U2071 (N_2071,N_1248,N_1084);
and U2072 (N_2072,N_1810,N_1266);
nand U2073 (N_2073,N_1581,N_1887);
nand U2074 (N_2074,N_1570,N_1878);
nand U2075 (N_2075,N_1286,N_1880);
nand U2076 (N_2076,N_1054,N_1367);
nor U2077 (N_2077,N_1481,N_1789);
and U2078 (N_2078,N_1185,N_1841);
nor U2079 (N_2079,N_1205,N_1065);
xor U2080 (N_2080,N_1542,N_1146);
nand U2081 (N_2081,N_1627,N_1778);
nand U2082 (N_2082,N_1737,N_1606);
nor U2083 (N_2083,N_1148,N_1402);
xor U2084 (N_2084,N_1646,N_1071);
or U2085 (N_2085,N_1206,N_1690);
and U2086 (N_2086,N_1279,N_1304);
xnor U2087 (N_2087,N_1858,N_1311);
and U2088 (N_2088,N_1610,N_1658);
or U2089 (N_2089,N_1489,N_1354);
xnor U2090 (N_2090,N_1187,N_1786);
and U2091 (N_2091,N_1514,N_1920);
or U2092 (N_2092,N_1330,N_1523);
nand U2093 (N_2093,N_1861,N_1723);
xnor U2094 (N_2094,N_1519,N_1787);
xor U2095 (N_2095,N_1970,N_1501);
xor U2096 (N_2096,N_1949,N_1855);
and U2097 (N_2097,N_1360,N_1118);
nor U2098 (N_2098,N_1021,N_1734);
or U2099 (N_2099,N_1751,N_1170);
or U2100 (N_2100,N_1480,N_1998);
nand U2101 (N_2101,N_1530,N_1052);
nand U2102 (N_2102,N_1213,N_1780);
nand U2103 (N_2103,N_1126,N_1356);
xnor U2104 (N_2104,N_1859,N_1791);
nand U2105 (N_2105,N_1713,N_1838);
and U2106 (N_2106,N_1660,N_1769);
nand U2107 (N_2107,N_1484,N_1515);
nor U2108 (N_2108,N_1416,N_1911);
xor U2109 (N_2109,N_1503,N_1881);
and U2110 (N_2110,N_1825,N_1979);
nand U2111 (N_2111,N_1784,N_1066);
or U2112 (N_2112,N_1650,N_1452);
nand U2113 (N_2113,N_1893,N_1852);
or U2114 (N_2114,N_1937,N_1848);
or U2115 (N_2115,N_1669,N_1485);
nand U2116 (N_2116,N_1094,N_1586);
or U2117 (N_2117,N_1764,N_1724);
and U2118 (N_2118,N_1122,N_1260);
or U2119 (N_2119,N_1323,N_1526);
and U2120 (N_2120,N_1337,N_1289);
and U2121 (N_2121,N_1396,N_1826);
nand U2122 (N_2122,N_1137,N_1171);
or U2123 (N_2123,N_1613,N_1068);
nand U2124 (N_2124,N_1679,N_1234);
xor U2125 (N_2125,N_1758,N_1077);
or U2126 (N_2126,N_1028,N_1539);
and U2127 (N_2127,N_1313,N_1113);
and U2128 (N_2128,N_1405,N_1419);
nor U2129 (N_2129,N_1045,N_1412);
xnor U2130 (N_2130,N_1935,N_1712);
xnor U2131 (N_2131,N_1808,N_1104);
nand U2132 (N_2132,N_1217,N_1194);
xor U2133 (N_2133,N_1482,N_1850);
and U2134 (N_2134,N_1781,N_1270);
nor U2135 (N_2135,N_1562,N_1680);
xnor U2136 (N_2136,N_1834,N_1592);
nand U2137 (N_2137,N_1423,N_1144);
nor U2138 (N_2138,N_1127,N_1301);
and U2139 (N_2139,N_1954,N_1264);
or U2140 (N_2140,N_1442,N_1522);
xor U2141 (N_2141,N_1225,N_1741);
nand U2142 (N_2142,N_1003,N_1049);
and U2143 (N_2143,N_1473,N_1212);
or U2144 (N_2144,N_1244,N_1816);
nor U2145 (N_2145,N_1051,N_1796);
nand U2146 (N_2146,N_1271,N_1156);
nor U2147 (N_2147,N_1455,N_1426);
or U2148 (N_2148,N_1710,N_1114);
xnor U2149 (N_2149,N_1776,N_1292);
xor U2150 (N_2150,N_1004,N_1875);
or U2151 (N_2151,N_1929,N_1326);
xor U2152 (N_2152,N_1267,N_1263);
nor U2153 (N_2153,N_1783,N_1706);
nand U2154 (N_2154,N_1060,N_1078);
and U2155 (N_2155,N_1090,N_1568);
xor U2156 (N_2156,N_1287,N_1398);
xor U2157 (N_2157,N_1296,N_1597);
and U2158 (N_2158,N_1392,N_1753);
and U2159 (N_2159,N_1245,N_1535);
nand U2160 (N_2160,N_1319,N_1062);
or U2161 (N_2161,N_1840,N_1874);
nor U2162 (N_2162,N_1812,N_1643);
xor U2163 (N_2163,N_1634,N_1216);
xnor U2164 (N_2164,N_1528,N_1092);
xor U2165 (N_2165,N_1897,N_1269);
nor U2166 (N_2166,N_1981,N_1327);
nor U2167 (N_2167,N_1651,N_1007);
nand U2168 (N_2168,N_1543,N_1457);
xnor U2169 (N_2169,N_1945,N_1676);
or U2170 (N_2170,N_1018,N_1444);
xor U2171 (N_2171,N_1559,N_1491);
or U2172 (N_2172,N_1253,N_1566);
xor U2173 (N_2173,N_1757,N_1720);
nor U2174 (N_2174,N_1409,N_1070);
and U2175 (N_2175,N_1117,N_1030);
or U2176 (N_2176,N_1888,N_1692);
and U2177 (N_2177,N_1362,N_1790);
or U2178 (N_2178,N_1160,N_1999);
or U2179 (N_2179,N_1906,N_1860);
nor U2180 (N_2180,N_1638,N_1908);
xor U2181 (N_2181,N_1797,N_1707);
nand U2182 (N_2182,N_1702,N_1309);
or U2183 (N_2183,N_1938,N_1064);
xnor U2184 (N_2184,N_1971,N_1366);
nand U2185 (N_2185,N_1359,N_1046);
xor U2186 (N_2186,N_1058,N_1133);
nand U2187 (N_2187,N_1635,N_1496);
or U2188 (N_2188,N_1015,N_1694);
or U2189 (N_2189,N_1583,N_1916);
and U2190 (N_2190,N_1995,N_1202);
xor U2191 (N_2191,N_1161,N_1306);
or U2192 (N_2192,N_1714,N_1839);
and U2193 (N_2193,N_1576,N_1733);
or U2194 (N_2194,N_1134,N_1176);
nor U2195 (N_2195,N_1130,N_1890);
and U2196 (N_2196,N_1506,N_1620);
nand U2197 (N_2197,N_1988,N_1179);
nor U2198 (N_2198,N_1023,N_1466);
or U2199 (N_2199,N_1119,N_1830);
xnor U2200 (N_2200,N_1096,N_1564);
nand U2201 (N_2201,N_1305,N_1632);
or U2202 (N_2202,N_1699,N_1538);
nor U2203 (N_2203,N_1494,N_1725);
nand U2204 (N_2204,N_1821,N_1002);
xnor U2205 (N_2205,N_1490,N_1965);
and U2206 (N_2206,N_1766,N_1449);
and U2207 (N_2207,N_1832,N_1338);
nor U2208 (N_2208,N_1794,N_1440);
nor U2209 (N_2209,N_1293,N_1993);
or U2210 (N_2210,N_1197,N_1919);
or U2211 (N_2211,N_1961,N_1549);
or U2212 (N_2212,N_1837,N_1290);
xnor U2213 (N_2213,N_1894,N_1607);
nor U2214 (N_2214,N_1321,N_1901);
and U2215 (N_2215,N_1554,N_1502);
and U2216 (N_2216,N_1792,N_1960);
and U2217 (N_2217,N_1460,N_1022);
xnor U2218 (N_2218,N_1715,N_1738);
nor U2219 (N_2219,N_1772,N_1450);
xor U2220 (N_2220,N_1541,N_1358);
or U2221 (N_2221,N_1163,N_1470);
or U2222 (N_2222,N_1788,N_1191);
nand U2223 (N_2223,N_1879,N_1325);
nor U2224 (N_2224,N_1430,N_1990);
nor U2225 (N_2225,N_1511,N_1555);
nand U2226 (N_2226,N_1384,N_1138);
nor U2227 (N_2227,N_1964,N_1507);
xor U2228 (N_2228,N_1410,N_1136);
and U2229 (N_2229,N_1153,N_1891);
nor U2230 (N_2230,N_1347,N_1391);
and U2231 (N_2231,N_1093,N_1947);
and U2232 (N_2232,N_1900,N_1131);
xor U2233 (N_2233,N_1164,N_1976);
or U2234 (N_2234,N_1320,N_1368);
nand U2235 (N_2235,N_1128,N_1563);
and U2236 (N_2236,N_1422,N_1238);
nand U2237 (N_2237,N_1687,N_1483);
or U2238 (N_2238,N_1278,N_1383);
nand U2239 (N_2239,N_1969,N_1162);
xor U2240 (N_2240,N_1394,N_1414);
xnor U2241 (N_2241,N_1609,N_1582);
nor U2242 (N_2242,N_1400,N_1558);
xnor U2243 (N_2243,N_1343,N_1302);
xor U2244 (N_2244,N_1590,N_1868);
nand U2245 (N_2245,N_1006,N_1529);
xor U2246 (N_2246,N_1039,N_1350);
nand U2247 (N_2247,N_1428,N_1203);
or U2248 (N_2248,N_1275,N_1295);
or U2249 (N_2249,N_1258,N_1172);
or U2250 (N_2250,N_1011,N_1956);
nand U2251 (N_2251,N_1441,N_1845);
or U2252 (N_2252,N_1742,N_1097);
nand U2253 (N_2253,N_1393,N_1629);
nand U2254 (N_2254,N_1116,N_1656);
nor U2255 (N_2255,N_1324,N_1285);
nor U2256 (N_2256,N_1577,N_1793);
or U2257 (N_2257,N_1940,N_1492);
xnor U2258 (N_2258,N_1333,N_1510);
and U2259 (N_2259,N_1322,N_1331);
or U2260 (N_2260,N_1898,N_1804);
xor U2261 (N_2261,N_1849,N_1917);
nand U2262 (N_2262,N_1214,N_1572);
xor U2263 (N_2263,N_1299,N_1499);
or U2264 (N_2264,N_1432,N_1446);
and U2265 (N_2265,N_1017,N_1531);
nand U2266 (N_2266,N_1630,N_1589);
xnor U2267 (N_2267,N_1073,N_1612);
or U2268 (N_2268,N_1199,N_1208);
nor U2269 (N_2269,N_1771,N_1041);
xnor U2270 (N_2270,N_1151,N_1798);
or U2271 (N_2271,N_1958,N_1291);
nor U2272 (N_2272,N_1380,N_1135);
and U2273 (N_2273,N_1184,N_1824);
or U2274 (N_2274,N_1369,N_1277);
and U2275 (N_2275,N_1477,N_1728);
nand U2276 (N_2276,N_1641,N_1833);
nand U2277 (N_2277,N_1882,N_1844);
nor U2278 (N_2278,N_1132,N_1181);
nor U2279 (N_2279,N_1928,N_1722);
and U2280 (N_2280,N_1854,N_1892);
or U2281 (N_2281,N_1765,N_1069);
xnor U2282 (N_2282,N_1421,N_1866);
or U2283 (N_2283,N_1280,N_1719);
or U2284 (N_2284,N_1693,N_1038);
or U2285 (N_2285,N_1063,N_1851);
nor U2286 (N_2286,N_1497,N_1475);
nand U2287 (N_2287,N_1767,N_1747);
nor U2288 (N_2288,N_1186,N_1315);
nor U2289 (N_2289,N_1339,N_1053);
or U2290 (N_2290,N_1918,N_1282);
nor U2291 (N_2291,N_1835,N_1910);
and U2292 (N_2292,N_1142,N_1904);
xnor U2293 (N_2293,N_1726,N_1774);
xnor U2294 (N_2294,N_1036,N_1518);
nor U2295 (N_2295,N_1623,N_1686);
nor U2296 (N_2296,N_1454,N_1561);
and U2297 (N_2297,N_1232,N_1207);
nor U2298 (N_2298,N_1755,N_1385);
nor U2299 (N_2299,N_1700,N_1124);
nor U2300 (N_2300,N_1020,N_1310);
nor U2301 (N_2301,N_1598,N_1717);
nand U2302 (N_2302,N_1476,N_1927);
nand U2303 (N_2303,N_1067,N_1079);
or U2304 (N_2304,N_1209,N_1427);
or U2305 (N_2305,N_1406,N_1649);
xor U2306 (N_2306,N_1671,N_1239);
xor U2307 (N_2307,N_1827,N_1602);
or U2308 (N_2308,N_1599,N_1259);
nor U2309 (N_2309,N_1735,N_1370);
or U2310 (N_2310,N_1283,N_1418);
nand U2311 (N_2311,N_1924,N_1178);
or U2312 (N_2312,N_1803,N_1106);
or U2313 (N_2313,N_1631,N_1955);
nand U2314 (N_2314,N_1504,N_1505);
and U2315 (N_2315,N_1536,N_1294);
nor U2316 (N_2316,N_1642,N_1459);
xnor U2317 (N_2317,N_1210,N_1000);
and U2318 (N_2318,N_1759,N_1773);
xnor U2319 (N_2319,N_1037,N_1950);
or U2320 (N_2320,N_1274,N_1624);
nor U2321 (N_2321,N_1474,N_1219);
or U2322 (N_2322,N_1863,N_1047);
and U2323 (N_2323,N_1195,N_1711);
and U2324 (N_2324,N_1344,N_1364);
and U2325 (N_2325,N_1752,N_1685);
or U2326 (N_2326,N_1963,N_1869);
or U2327 (N_2327,N_1390,N_1029);
nand U2328 (N_2328,N_1647,N_1317);
nand U2329 (N_2329,N_1903,N_1407);
or U2330 (N_2330,N_1843,N_1872);
xnor U2331 (N_2331,N_1637,N_1169);
nand U2332 (N_2332,N_1140,N_1342);
and U2333 (N_2333,N_1967,N_1946);
or U2334 (N_2334,N_1984,N_1867);
xnor U2335 (N_2335,N_1415,N_1551);
xnor U2336 (N_2336,N_1276,N_1667);
and U2337 (N_2337,N_1183,N_1080);
nor U2338 (N_2338,N_1820,N_1513);
xor U2339 (N_2339,N_1019,N_1372);
or U2340 (N_2340,N_1125,N_1828);
xor U2341 (N_2341,N_1533,N_1157);
and U2342 (N_2342,N_1182,N_1168);
nand U2343 (N_2343,N_1013,N_1075);
xor U2344 (N_2344,N_1042,N_1395);
and U2345 (N_2345,N_1154,N_1349);
xnor U2346 (N_2346,N_1557,N_1089);
xor U2347 (N_2347,N_1871,N_1222);
nor U2348 (N_2348,N_1035,N_1224);
nor U2349 (N_2349,N_1524,N_1180);
and U2350 (N_2350,N_1425,N_1925);
xnor U2351 (N_2351,N_1159,N_1997);
xor U2352 (N_2352,N_1158,N_1382);
xnor U2353 (N_2353,N_1404,N_1281);
xnor U2354 (N_2354,N_1775,N_1962);
xor U2355 (N_2355,N_1628,N_1009);
nor U2356 (N_2356,N_1739,N_1227);
nor U2357 (N_2357,N_1678,N_1856);
and U2358 (N_2358,N_1329,N_1108);
or U2359 (N_2359,N_1626,N_1300);
nor U2360 (N_2360,N_1913,N_1760);
xor U2361 (N_2361,N_1048,N_1544);
nor U2362 (N_2362,N_1098,N_1857);
or U2363 (N_2363,N_1525,N_1732);
and U2364 (N_2364,N_1026,N_1569);
or U2365 (N_2365,N_1512,N_1663);
or U2366 (N_2366,N_1941,N_1200);
xnor U2367 (N_2367,N_1240,N_1931);
xor U2368 (N_2368,N_1811,N_1088);
nor U2369 (N_2369,N_1014,N_1785);
and U2370 (N_2370,N_1746,N_1149);
and U2371 (N_2371,N_1978,N_1033);
nand U2372 (N_2372,N_1591,N_1031);
or U2373 (N_2373,N_1167,N_1968);
nand U2374 (N_2374,N_1593,N_1332);
nand U2375 (N_2375,N_1975,N_1192);
or U2376 (N_2376,N_1353,N_1189);
or U2377 (N_2377,N_1303,N_1622);
or U2378 (N_2378,N_1579,N_1654);
nand U2379 (N_2379,N_1705,N_1235);
nor U2380 (N_2380,N_1488,N_1652);
nand U2381 (N_2381,N_1777,N_1408);
or U2382 (N_2382,N_1251,N_1727);
xor U2383 (N_2383,N_1221,N_1346);
xor U2384 (N_2384,N_1255,N_1508);
nor U2385 (N_2385,N_1942,N_1381);
nand U2386 (N_2386,N_1905,N_1223);
and U2387 (N_2387,N_1683,N_1374);
or U2388 (N_2388,N_1616,N_1439);
xnor U2389 (N_2389,N_1684,N_1341);
nor U2390 (N_2390,N_1373,N_1749);
or U2391 (N_2391,N_1744,N_1008);
or U2392 (N_2392,N_1107,N_1983);
nand U2393 (N_2393,N_1704,N_1307);
nand U2394 (N_2394,N_1252,N_1923);
and U2395 (N_2395,N_1799,N_1498);
or U2396 (N_2396,N_1708,N_1980);
nor U2397 (N_2397,N_1636,N_1121);
xor U2398 (N_2398,N_1648,N_1143);
nor U2399 (N_2399,N_1413,N_1853);
nor U2400 (N_2400,N_1695,N_1215);
xor U2401 (N_2401,N_1099,N_1371);
and U2402 (N_2402,N_1471,N_1056);
xor U2403 (N_2403,N_1883,N_1619);
and U2404 (N_2404,N_1761,N_1639);
nand U2405 (N_2405,N_1388,N_1842);
xnor U2406 (N_2406,N_1453,N_1633);
xnor U2407 (N_2407,N_1467,N_1417);
or U2408 (N_2408,N_1936,N_1540);
nand U2409 (N_2409,N_1265,N_1081);
or U2410 (N_2410,N_1573,N_1604);
and U2411 (N_2411,N_1433,N_1657);
or U2412 (N_2412,N_1249,N_1876);
nand U2413 (N_2413,N_1653,N_1086);
nand U2414 (N_2414,N_1500,N_1655);
nand U2415 (N_2415,N_1762,N_1829);
or U2416 (N_2416,N_1915,N_1640);
or U2417 (N_2417,N_1560,N_1584);
or U2418 (N_2418,N_1575,N_1478);
xnor U2419 (N_2419,N_1977,N_1914);
xor U2420 (N_2420,N_1585,N_1236);
nor U2421 (N_2421,N_1072,N_1288);
xnor U2422 (N_2422,N_1101,N_1922);
and U2423 (N_2423,N_1748,N_1201);
nor U2424 (N_2424,N_1959,N_1487);
nand U2425 (N_2425,N_1257,N_1836);
or U2426 (N_2426,N_1813,N_1316);
nand U2427 (N_2427,N_1550,N_1155);
nand U2428 (N_2428,N_1673,N_1082);
xor U2429 (N_2429,N_1895,N_1603);
and U2430 (N_2430,N_1308,N_1246);
nand U2431 (N_2431,N_1469,N_1548);
nand U2432 (N_2432,N_1546,N_1665);
nor U2433 (N_2433,N_1074,N_1102);
and U2434 (N_2434,N_1429,N_1486);
xnor U2435 (N_2435,N_1516,N_1709);
and U2436 (N_2436,N_1016,N_1076);
and U2437 (N_2437,N_1688,N_1886);
or U2438 (N_2438,N_1447,N_1479);
or U2439 (N_2439,N_1435,N_1670);
nor U2440 (N_2440,N_1580,N_1899);
xnor U2441 (N_2441,N_1218,N_1448);
xor U2442 (N_2442,N_1902,N_1005);
nand U2443 (N_2443,N_1721,N_1083);
nand U2444 (N_2444,N_1907,N_1351);
xor U2445 (N_2445,N_1985,N_1689);
nor U2446 (N_2446,N_1025,N_1740);
nand U2447 (N_2447,N_1230,N_1411);
or U2448 (N_2448,N_1420,N_1930);
nor U2449 (N_2449,N_1818,N_1807);
and U2450 (N_2450,N_1809,N_1534);
xor U2451 (N_2451,N_1939,N_1666);
nand U2452 (N_2452,N_1174,N_1401);
nand U2453 (N_2453,N_1087,N_1399);
nand U2454 (N_2454,N_1696,N_1621);
or U2455 (N_2455,N_1953,N_1847);
nor U2456 (N_2456,N_1763,N_1509);
or U2457 (N_2457,N_1085,N_1111);
and U2458 (N_2458,N_1884,N_1691);
and U2459 (N_2459,N_1273,N_1250);
and U2460 (N_2460,N_1352,N_1123);
and U2461 (N_2461,N_1220,N_1571);
or U2462 (N_2462,N_1061,N_1973);
nand U2463 (N_2463,N_1600,N_1032);
and U2464 (N_2464,N_1458,N_1729);
and U2465 (N_2465,N_1877,N_1443);
and U2466 (N_2466,N_1363,N_1517);
nand U2467 (N_2467,N_1261,N_1050);
nor U2468 (N_2468,N_1152,N_1233);
xnor U2469 (N_2469,N_1377,N_1608);
and U2470 (N_2470,N_1228,N_1547);
or U2471 (N_2471,N_1823,N_1736);
nor U2472 (N_2472,N_1437,N_1336);
xor U2473 (N_2473,N_1055,N_1365);
xor U2474 (N_2474,N_1815,N_1105);
nor U2475 (N_2475,N_1188,N_1982);
nand U2476 (N_2476,N_1802,N_1112);
nand U2477 (N_2477,N_1145,N_1147);
xor U2478 (N_2478,N_1424,N_1379);
nor U2479 (N_2479,N_1348,N_1141);
nor U2480 (N_2480,N_1010,N_1682);
nand U2481 (N_2481,N_1109,N_1044);
or U2482 (N_2482,N_1909,N_1165);
xor U2483 (N_2483,N_1231,N_1870);
nor U2484 (N_2484,N_1805,N_1537);
nor U2485 (N_2485,N_1556,N_1386);
and U2486 (N_2486,N_1974,N_1462);
nor U2487 (N_2487,N_1314,N_1472);
nor U2488 (N_2488,N_1770,N_1553);
nor U2489 (N_2489,N_1605,N_1204);
xnor U2490 (N_2490,N_1527,N_1814);
nor U2491 (N_2491,N_1730,N_1944);
nand U2492 (N_2492,N_1355,N_1298);
xor U2493 (N_2493,N_1951,N_1027);
nand U2494 (N_2494,N_1243,N_1456);
nor U2495 (N_2495,N_1661,N_1731);
nor U2496 (N_2496,N_1921,N_1819);
nand U2497 (N_2497,N_1754,N_1318);
xor U2498 (N_2498,N_1587,N_1040);
and U2499 (N_2499,N_1403,N_1247);
nor U2500 (N_2500,N_1090,N_1266);
nand U2501 (N_2501,N_1865,N_1970);
nor U2502 (N_2502,N_1481,N_1642);
nand U2503 (N_2503,N_1587,N_1426);
nor U2504 (N_2504,N_1751,N_1004);
and U2505 (N_2505,N_1060,N_1390);
xor U2506 (N_2506,N_1794,N_1744);
and U2507 (N_2507,N_1270,N_1796);
xor U2508 (N_2508,N_1776,N_1895);
nor U2509 (N_2509,N_1657,N_1675);
and U2510 (N_2510,N_1647,N_1960);
nor U2511 (N_2511,N_1082,N_1424);
nand U2512 (N_2512,N_1820,N_1793);
or U2513 (N_2513,N_1865,N_1803);
and U2514 (N_2514,N_1325,N_1309);
nand U2515 (N_2515,N_1088,N_1375);
or U2516 (N_2516,N_1805,N_1204);
nand U2517 (N_2517,N_1093,N_1547);
nor U2518 (N_2518,N_1967,N_1527);
nor U2519 (N_2519,N_1291,N_1683);
nand U2520 (N_2520,N_1293,N_1217);
nor U2521 (N_2521,N_1181,N_1999);
xnor U2522 (N_2522,N_1762,N_1787);
or U2523 (N_2523,N_1262,N_1979);
nor U2524 (N_2524,N_1228,N_1674);
xor U2525 (N_2525,N_1710,N_1134);
xnor U2526 (N_2526,N_1996,N_1310);
nor U2527 (N_2527,N_1631,N_1834);
nor U2528 (N_2528,N_1774,N_1244);
and U2529 (N_2529,N_1115,N_1963);
xor U2530 (N_2530,N_1714,N_1258);
nand U2531 (N_2531,N_1422,N_1713);
nand U2532 (N_2532,N_1403,N_1048);
xor U2533 (N_2533,N_1799,N_1714);
nand U2534 (N_2534,N_1545,N_1315);
and U2535 (N_2535,N_1531,N_1525);
or U2536 (N_2536,N_1221,N_1183);
xor U2537 (N_2537,N_1575,N_1440);
nand U2538 (N_2538,N_1684,N_1481);
or U2539 (N_2539,N_1131,N_1830);
or U2540 (N_2540,N_1462,N_1761);
nand U2541 (N_2541,N_1876,N_1389);
xor U2542 (N_2542,N_1986,N_1860);
xor U2543 (N_2543,N_1167,N_1525);
and U2544 (N_2544,N_1529,N_1174);
xor U2545 (N_2545,N_1419,N_1828);
nor U2546 (N_2546,N_1983,N_1898);
and U2547 (N_2547,N_1635,N_1662);
or U2548 (N_2548,N_1553,N_1689);
xnor U2549 (N_2549,N_1589,N_1233);
and U2550 (N_2550,N_1172,N_1024);
nor U2551 (N_2551,N_1984,N_1023);
and U2552 (N_2552,N_1797,N_1057);
xnor U2553 (N_2553,N_1638,N_1051);
nand U2554 (N_2554,N_1079,N_1576);
nor U2555 (N_2555,N_1734,N_1964);
xor U2556 (N_2556,N_1073,N_1735);
xnor U2557 (N_2557,N_1192,N_1058);
nand U2558 (N_2558,N_1214,N_1767);
and U2559 (N_2559,N_1063,N_1903);
or U2560 (N_2560,N_1037,N_1867);
or U2561 (N_2561,N_1308,N_1839);
nor U2562 (N_2562,N_1078,N_1583);
xor U2563 (N_2563,N_1607,N_1514);
xnor U2564 (N_2564,N_1447,N_1732);
or U2565 (N_2565,N_1757,N_1311);
nor U2566 (N_2566,N_1386,N_1024);
nand U2567 (N_2567,N_1122,N_1270);
nand U2568 (N_2568,N_1274,N_1760);
xnor U2569 (N_2569,N_1983,N_1142);
nand U2570 (N_2570,N_1318,N_1674);
xor U2571 (N_2571,N_1274,N_1483);
and U2572 (N_2572,N_1999,N_1604);
and U2573 (N_2573,N_1063,N_1248);
xor U2574 (N_2574,N_1239,N_1297);
nand U2575 (N_2575,N_1261,N_1540);
nor U2576 (N_2576,N_1867,N_1439);
nand U2577 (N_2577,N_1615,N_1318);
and U2578 (N_2578,N_1940,N_1002);
or U2579 (N_2579,N_1955,N_1181);
nand U2580 (N_2580,N_1996,N_1720);
nor U2581 (N_2581,N_1657,N_1948);
nand U2582 (N_2582,N_1905,N_1403);
or U2583 (N_2583,N_1382,N_1130);
xnor U2584 (N_2584,N_1396,N_1113);
and U2585 (N_2585,N_1447,N_1209);
nand U2586 (N_2586,N_1400,N_1941);
and U2587 (N_2587,N_1003,N_1969);
nand U2588 (N_2588,N_1599,N_1825);
nor U2589 (N_2589,N_1130,N_1105);
and U2590 (N_2590,N_1688,N_1989);
nand U2591 (N_2591,N_1067,N_1264);
nand U2592 (N_2592,N_1634,N_1545);
xor U2593 (N_2593,N_1017,N_1396);
nand U2594 (N_2594,N_1236,N_1689);
nor U2595 (N_2595,N_1985,N_1056);
xnor U2596 (N_2596,N_1402,N_1303);
xor U2597 (N_2597,N_1273,N_1459);
xor U2598 (N_2598,N_1393,N_1073);
nor U2599 (N_2599,N_1676,N_1549);
or U2600 (N_2600,N_1965,N_1348);
xor U2601 (N_2601,N_1041,N_1988);
or U2602 (N_2602,N_1737,N_1903);
xnor U2603 (N_2603,N_1853,N_1638);
xnor U2604 (N_2604,N_1068,N_1536);
xor U2605 (N_2605,N_1491,N_1394);
nand U2606 (N_2606,N_1713,N_1166);
and U2607 (N_2607,N_1019,N_1665);
xnor U2608 (N_2608,N_1284,N_1848);
or U2609 (N_2609,N_1179,N_1858);
or U2610 (N_2610,N_1157,N_1321);
and U2611 (N_2611,N_1957,N_1164);
or U2612 (N_2612,N_1965,N_1896);
nor U2613 (N_2613,N_1957,N_1829);
nor U2614 (N_2614,N_1951,N_1494);
or U2615 (N_2615,N_1596,N_1056);
nand U2616 (N_2616,N_1777,N_1929);
or U2617 (N_2617,N_1626,N_1413);
and U2618 (N_2618,N_1335,N_1209);
nor U2619 (N_2619,N_1901,N_1931);
and U2620 (N_2620,N_1550,N_1340);
xnor U2621 (N_2621,N_1322,N_1876);
or U2622 (N_2622,N_1951,N_1573);
nand U2623 (N_2623,N_1060,N_1885);
xnor U2624 (N_2624,N_1140,N_1974);
and U2625 (N_2625,N_1865,N_1491);
or U2626 (N_2626,N_1212,N_1389);
xor U2627 (N_2627,N_1766,N_1313);
nand U2628 (N_2628,N_1821,N_1737);
and U2629 (N_2629,N_1040,N_1548);
nor U2630 (N_2630,N_1564,N_1701);
xor U2631 (N_2631,N_1928,N_1126);
or U2632 (N_2632,N_1283,N_1409);
nand U2633 (N_2633,N_1510,N_1604);
xnor U2634 (N_2634,N_1460,N_1749);
or U2635 (N_2635,N_1334,N_1006);
and U2636 (N_2636,N_1294,N_1358);
nor U2637 (N_2637,N_1544,N_1670);
nor U2638 (N_2638,N_1103,N_1948);
nor U2639 (N_2639,N_1283,N_1272);
and U2640 (N_2640,N_1052,N_1987);
nand U2641 (N_2641,N_1903,N_1383);
nand U2642 (N_2642,N_1762,N_1061);
nor U2643 (N_2643,N_1526,N_1924);
nand U2644 (N_2644,N_1701,N_1084);
xnor U2645 (N_2645,N_1307,N_1388);
nand U2646 (N_2646,N_1235,N_1241);
or U2647 (N_2647,N_1614,N_1421);
and U2648 (N_2648,N_1464,N_1343);
nor U2649 (N_2649,N_1125,N_1242);
or U2650 (N_2650,N_1603,N_1049);
xor U2651 (N_2651,N_1885,N_1386);
and U2652 (N_2652,N_1067,N_1534);
and U2653 (N_2653,N_1020,N_1983);
and U2654 (N_2654,N_1878,N_1531);
nor U2655 (N_2655,N_1396,N_1592);
xor U2656 (N_2656,N_1896,N_1911);
nor U2657 (N_2657,N_1304,N_1059);
xor U2658 (N_2658,N_1957,N_1797);
nand U2659 (N_2659,N_1982,N_1580);
xor U2660 (N_2660,N_1091,N_1270);
nand U2661 (N_2661,N_1123,N_1510);
xnor U2662 (N_2662,N_1281,N_1162);
xnor U2663 (N_2663,N_1968,N_1948);
nor U2664 (N_2664,N_1514,N_1557);
nor U2665 (N_2665,N_1477,N_1157);
xor U2666 (N_2666,N_1938,N_1795);
xor U2667 (N_2667,N_1607,N_1331);
nand U2668 (N_2668,N_1474,N_1997);
nand U2669 (N_2669,N_1315,N_1275);
or U2670 (N_2670,N_1877,N_1486);
and U2671 (N_2671,N_1501,N_1155);
and U2672 (N_2672,N_1955,N_1622);
nor U2673 (N_2673,N_1841,N_1593);
nor U2674 (N_2674,N_1930,N_1850);
and U2675 (N_2675,N_1477,N_1856);
xnor U2676 (N_2676,N_1550,N_1980);
nor U2677 (N_2677,N_1181,N_1547);
xor U2678 (N_2678,N_1617,N_1936);
and U2679 (N_2679,N_1604,N_1995);
xor U2680 (N_2680,N_1505,N_1782);
and U2681 (N_2681,N_1542,N_1261);
and U2682 (N_2682,N_1952,N_1805);
or U2683 (N_2683,N_1025,N_1300);
nand U2684 (N_2684,N_1316,N_1832);
or U2685 (N_2685,N_1437,N_1385);
nand U2686 (N_2686,N_1964,N_1762);
and U2687 (N_2687,N_1767,N_1395);
nor U2688 (N_2688,N_1319,N_1915);
or U2689 (N_2689,N_1030,N_1683);
nand U2690 (N_2690,N_1896,N_1691);
nand U2691 (N_2691,N_1586,N_1840);
nand U2692 (N_2692,N_1056,N_1846);
and U2693 (N_2693,N_1315,N_1716);
and U2694 (N_2694,N_1377,N_1208);
nand U2695 (N_2695,N_1315,N_1592);
xnor U2696 (N_2696,N_1886,N_1356);
and U2697 (N_2697,N_1251,N_1123);
nand U2698 (N_2698,N_1533,N_1406);
or U2699 (N_2699,N_1636,N_1488);
and U2700 (N_2700,N_1718,N_1618);
or U2701 (N_2701,N_1019,N_1257);
xnor U2702 (N_2702,N_1474,N_1785);
nor U2703 (N_2703,N_1191,N_1627);
nand U2704 (N_2704,N_1776,N_1728);
xor U2705 (N_2705,N_1212,N_1414);
and U2706 (N_2706,N_1654,N_1110);
nand U2707 (N_2707,N_1771,N_1505);
nand U2708 (N_2708,N_1876,N_1772);
or U2709 (N_2709,N_1215,N_1618);
xnor U2710 (N_2710,N_1983,N_1328);
or U2711 (N_2711,N_1625,N_1719);
nor U2712 (N_2712,N_1335,N_1974);
nand U2713 (N_2713,N_1350,N_1052);
nor U2714 (N_2714,N_1692,N_1167);
and U2715 (N_2715,N_1609,N_1347);
nor U2716 (N_2716,N_1503,N_1839);
or U2717 (N_2717,N_1692,N_1881);
and U2718 (N_2718,N_1542,N_1854);
nand U2719 (N_2719,N_1149,N_1846);
or U2720 (N_2720,N_1988,N_1752);
nor U2721 (N_2721,N_1130,N_1522);
nand U2722 (N_2722,N_1554,N_1597);
or U2723 (N_2723,N_1255,N_1655);
nor U2724 (N_2724,N_1837,N_1174);
nor U2725 (N_2725,N_1907,N_1748);
or U2726 (N_2726,N_1966,N_1421);
xor U2727 (N_2727,N_1505,N_1693);
nand U2728 (N_2728,N_1335,N_1285);
nand U2729 (N_2729,N_1515,N_1768);
xnor U2730 (N_2730,N_1612,N_1038);
nor U2731 (N_2731,N_1242,N_1052);
and U2732 (N_2732,N_1377,N_1165);
nor U2733 (N_2733,N_1911,N_1803);
xnor U2734 (N_2734,N_1202,N_1874);
or U2735 (N_2735,N_1338,N_1327);
nor U2736 (N_2736,N_1719,N_1715);
and U2737 (N_2737,N_1730,N_1298);
nand U2738 (N_2738,N_1541,N_1162);
and U2739 (N_2739,N_1393,N_1215);
nor U2740 (N_2740,N_1033,N_1485);
or U2741 (N_2741,N_1802,N_1657);
xor U2742 (N_2742,N_1454,N_1342);
and U2743 (N_2743,N_1981,N_1003);
or U2744 (N_2744,N_1417,N_1130);
or U2745 (N_2745,N_1420,N_1323);
and U2746 (N_2746,N_1719,N_1414);
nor U2747 (N_2747,N_1553,N_1778);
nor U2748 (N_2748,N_1830,N_1536);
nor U2749 (N_2749,N_1818,N_1416);
xnor U2750 (N_2750,N_1272,N_1046);
xor U2751 (N_2751,N_1309,N_1732);
or U2752 (N_2752,N_1501,N_1750);
xnor U2753 (N_2753,N_1603,N_1314);
nand U2754 (N_2754,N_1473,N_1536);
nor U2755 (N_2755,N_1453,N_1696);
nor U2756 (N_2756,N_1179,N_1581);
or U2757 (N_2757,N_1100,N_1885);
nand U2758 (N_2758,N_1822,N_1185);
or U2759 (N_2759,N_1881,N_1145);
and U2760 (N_2760,N_1514,N_1342);
or U2761 (N_2761,N_1969,N_1118);
nand U2762 (N_2762,N_1748,N_1939);
or U2763 (N_2763,N_1057,N_1838);
xor U2764 (N_2764,N_1068,N_1122);
nor U2765 (N_2765,N_1836,N_1343);
nand U2766 (N_2766,N_1901,N_1366);
and U2767 (N_2767,N_1268,N_1369);
or U2768 (N_2768,N_1020,N_1166);
nand U2769 (N_2769,N_1503,N_1772);
nand U2770 (N_2770,N_1260,N_1818);
or U2771 (N_2771,N_1297,N_1386);
nor U2772 (N_2772,N_1800,N_1113);
nor U2773 (N_2773,N_1484,N_1463);
xor U2774 (N_2774,N_1712,N_1973);
or U2775 (N_2775,N_1733,N_1879);
or U2776 (N_2776,N_1488,N_1845);
nor U2777 (N_2777,N_1470,N_1501);
and U2778 (N_2778,N_1903,N_1003);
or U2779 (N_2779,N_1012,N_1289);
nand U2780 (N_2780,N_1359,N_1184);
nor U2781 (N_2781,N_1566,N_1043);
and U2782 (N_2782,N_1335,N_1495);
or U2783 (N_2783,N_1144,N_1127);
xor U2784 (N_2784,N_1226,N_1532);
and U2785 (N_2785,N_1582,N_1949);
nor U2786 (N_2786,N_1529,N_1517);
nand U2787 (N_2787,N_1449,N_1818);
or U2788 (N_2788,N_1147,N_1818);
nand U2789 (N_2789,N_1153,N_1546);
and U2790 (N_2790,N_1946,N_1344);
or U2791 (N_2791,N_1073,N_1098);
nor U2792 (N_2792,N_1981,N_1191);
xnor U2793 (N_2793,N_1677,N_1328);
and U2794 (N_2794,N_1286,N_1361);
xor U2795 (N_2795,N_1786,N_1255);
or U2796 (N_2796,N_1364,N_1713);
nand U2797 (N_2797,N_1323,N_1633);
nor U2798 (N_2798,N_1080,N_1845);
or U2799 (N_2799,N_1580,N_1006);
nand U2800 (N_2800,N_1927,N_1950);
nor U2801 (N_2801,N_1936,N_1588);
and U2802 (N_2802,N_1232,N_1816);
nor U2803 (N_2803,N_1825,N_1537);
nor U2804 (N_2804,N_1807,N_1592);
and U2805 (N_2805,N_1297,N_1885);
or U2806 (N_2806,N_1923,N_1137);
nand U2807 (N_2807,N_1517,N_1883);
nand U2808 (N_2808,N_1038,N_1857);
xnor U2809 (N_2809,N_1995,N_1000);
nor U2810 (N_2810,N_1243,N_1781);
and U2811 (N_2811,N_1238,N_1269);
xor U2812 (N_2812,N_1400,N_1094);
and U2813 (N_2813,N_1903,N_1110);
xnor U2814 (N_2814,N_1548,N_1855);
nand U2815 (N_2815,N_1902,N_1964);
nor U2816 (N_2816,N_1401,N_1514);
or U2817 (N_2817,N_1180,N_1464);
and U2818 (N_2818,N_1153,N_1704);
xnor U2819 (N_2819,N_1809,N_1324);
nand U2820 (N_2820,N_1591,N_1826);
nor U2821 (N_2821,N_1204,N_1862);
nor U2822 (N_2822,N_1846,N_1635);
nand U2823 (N_2823,N_1205,N_1903);
xnor U2824 (N_2824,N_1151,N_1584);
nor U2825 (N_2825,N_1786,N_1579);
or U2826 (N_2826,N_1628,N_1476);
or U2827 (N_2827,N_1144,N_1475);
or U2828 (N_2828,N_1123,N_1544);
and U2829 (N_2829,N_1061,N_1178);
or U2830 (N_2830,N_1806,N_1620);
nand U2831 (N_2831,N_1331,N_1792);
or U2832 (N_2832,N_1638,N_1046);
xor U2833 (N_2833,N_1792,N_1143);
nand U2834 (N_2834,N_1874,N_1985);
or U2835 (N_2835,N_1717,N_1979);
nand U2836 (N_2836,N_1746,N_1363);
nand U2837 (N_2837,N_1749,N_1479);
xor U2838 (N_2838,N_1619,N_1863);
or U2839 (N_2839,N_1472,N_1930);
xnor U2840 (N_2840,N_1608,N_1906);
xor U2841 (N_2841,N_1235,N_1343);
or U2842 (N_2842,N_1645,N_1850);
nand U2843 (N_2843,N_1176,N_1511);
nor U2844 (N_2844,N_1176,N_1501);
nand U2845 (N_2845,N_1615,N_1569);
nand U2846 (N_2846,N_1070,N_1678);
nand U2847 (N_2847,N_1980,N_1410);
or U2848 (N_2848,N_1563,N_1808);
xnor U2849 (N_2849,N_1197,N_1594);
and U2850 (N_2850,N_1134,N_1221);
or U2851 (N_2851,N_1240,N_1154);
and U2852 (N_2852,N_1304,N_1851);
and U2853 (N_2853,N_1274,N_1873);
xnor U2854 (N_2854,N_1976,N_1325);
or U2855 (N_2855,N_1951,N_1578);
nand U2856 (N_2856,N_1667,N_1062);
nand U2857 (N_2857,N_1268,N_1439);
or U2858 (N_2858,N_1109,N_1912);
or U2859 (N_2859,N_1335,N_1716);
xor U2860 (N_2860,N_1155,N_1679);
nor U2861 (N_2861,N_1591,N_1526);
or U2862 (N_2862,N_1178,N_1352);
xor U2863 (N_2863,N_1510,N_1816);
or U2864 (N_2864,N_1478,N_1821);
nand U2865 (N_2865,N_1348,N_1560);
or U2866 (N_2866,N_1144,N_1974);
nor U2867 (N_2867,N_1923,N_1673);
and U2868 (N_2868,N_1482,N_1867);
xor U2869 (N_2869,N_1427,N_1608);
or U2870 (N_2870,N_1928,N_1352);
nor U2871 (N_2871,N_1994,N_1793);
and U2872 (N_2872,N_1220,N_1139);
nand U2873 (N_2873,N_1235,N_1995);
xor U2874 (N_2874,N_1274,N_1055);
and U2875 (N_2875,N_1387,N_1994);
nand U2876 (N_2876,N_1569,N_1031);
or U2877 (N_2877,N_1704,N_1306);
and U2878 (N_2878,N_1153,N_1460);
nand U2879 (N_2879,N_1230,N_1486);
xor U2880 (N_2880,N_1070,N_1363);
xnor U2881 (N_2881,N_1388,N_1829);
nand U2882 (N_2882,N_1918,N_1563);
nand U2883 (N_2883,N_1457,N_1688);
and U2884 (N_2884,N_1150,N_1087);
or U2885 (N_2885,N_1648,N_1896);
and U2886 (N_2886,N_1639,N_1654);
nor U2887 (N_2887,N_1839,N_1986);
nand U2888 (N_2888,N_1798,N_1868);
or U2889 (N_2889,N_1368,N_1212);
or U2890 (N_2890,N_1468,N_1136);
and U2891 (N_2891,N_1542,N_1363);
nor U2892 (N_2892,N_1397,N_1687);
or U2893 (N_2893,N_1356,N_1428);
nand U2894 (N_2894,N_1828,N_1433);
and U2895 (N_2895,N_1268,N_1449);
or U2896 (N_2896,N_1677,N_1639);
nor U2897 (N_2897,N_1478,N_1692);
xnor U2898 (N_2898,N_1581,N_1616);
or U2899 (N_2899,N_1931,N_1101);
nand U2900 (N_2900,N_1270,N_1874);
or U2901 (N_2901,N_1896,N_1088);
and U2902 (N_2902,N_1776,N_1354);
xnor U2903 (N_2903,N_1255,N_1711);
or U2904 (N_2904,N_1294,N_1770);
and U2905 (N_2905,N_1995,N_1657);
or U2906 (N_2906,N_1503,N_1595);
and U2907 (N_2907,N_1253,N_1236);
xnor U2908 (N_2908,N_1780,N_1852);
nor U2909 (N_2909,N_1651,N_1722);
nor U2910 (N_2910,N_1635,N_1849);
xnor U2911 (N_2911,N_1431,N_1567);
nand U2912 (N_2912,N_1866,N_1180);
nand U2913 (N_2913,N_1709,N_1950);
xor U2914 (N_2914,N_1977,N_1476);
nor U2915 (N_2915,N_1218,N_1523);
nor U2916 (N_2916,N_1896,N_1169);
xor U2917 (N_2917,N_1260,N_1720);
xor U2918 (N_2918,N_1147,N_1638);
nor U2919 (N_2919,N_1604,N_1306);
xor U2920 (N_2920,N_1111,N_1007);
and U2921 (N_2921,N_1096,N_1754);
xor U2922 (N_2922,N_1665,N_1321);
nand U2923 (N_2923,N_1552,N_1290);
xnor U2924 (N_2924,N_1280,N_1331);
xor U2925 (N_2925,N_1798,N_1267);
xor U2926 (N_2926,N_1915,N_1844);
or U2927 (N_2927,N_1277,N_1815);
or U2928 (N_2928,N_1482,N_1279);
xor U2929 (N_2929,N_1908,N_1336);
nor U2930 (N_2930,N_1396,N_1943);
or U2931 (N_2931,N_1192,N_1804);
nor U2932 (N_2932,N_1824,N_1674);
nand U2933 (N_2933,N_1065,N_1176);
xnor U2934 (N_2934,N_1386,N_1101);
nand U2935 (N_2935,N_1724,N_1774);
xnor U2936 (N_2936,N_1364,N_1501);
nor U2937 (N_2937,N_1150,N_1248);
and U2938 (N_2938,N_1766,N_1653);
or U2939 (N_2939,N_1242,N_1709);
xnor U2940 (N_2940,N_1874,N_1214);
nand U2941 (N_2941,N_1713,N_1301);
or U2942 (N_2942,N_1967,N_1293);
xor U2943 (N_2943,N_1478,N_1603);
nor U2944 (N_2944,N_1406,N_1141);
xor U2945 (N_2945,N_1362,N_1062);
and U2946 (N_2946,N_1375,N_1977);
and U2947 (N_2947,N_1099,N_1404);
nand U2948 (N_2948,N_1424,N_1406);
nand U2949 (N_2949,N_1604,N_1795);
nand U2950 (N_2950,N_1497,N_1733);
and U2951 (N_2951,N_1072,N_1892);
nand U2952 (N_2952,N_1328,N_1869);
xnor U2953 (N_2953,N_1029,N_1966);
xor U2954 (N_2954,N_1935,N_1884);
or U2955 (N_2955,N_1161,N_1035);
nor U2956 (N_2956,N_1271,N_1414);
xor U2957 (N_2957,N_1293,N_1484);
xnor U2958 (N_2958,N_1623,N_1640);
nor U2959 (N_2959,N_1017,N_1689);
nor U2960 (N_2960,N_1430,N_1304);
xor U2961 (N_2961,N_1254,N_1923);
nand U2962 (N_2962,N_1079,N_1870);
nand U2963 (N_2963,N_1184,N_1355);
or U2964 (N_2964,N_1158,N_1911);
nand U2965 (N_2965,N_1504,N_1567);
and U2966 (N_2966,N_1459,N_1380);
xor U2967 (N_2967,N_1566,N_1805);
xnor U2968 (N_2968,N_1333,N_1683);
and U2969 (N_2969,N_1159,N_1445);
xnor U2970 (N_2970,N_1682,N_1742);
nor U2971 (N_2971,N_1528,N_1191);
nand U2972 (N_2972,N_1112,N_1213);
xor U2973 (N_2973,N_1353,N_1008);
xor U2974 (N_2974,N_1155,N_1066);
and U2975 (N_2975,N_1890,N_1745);
and U2976 (N_2976,N_1397,N_1403);
nand U2977 (N_2977,N_1860,N_1419);
nand U2978 (N_2978,N_1533,N_1639);
nand U2979 (N_2979,N_1558,N_1987);
xor U2980 (N_2980,N_1598,N_1793);
nor U2981 (N_2981,N_1256,N_1574);
or U2982 (N_2982,N_1186,N_1746);
nor U2983 (N_2983,N_1478,N_1510);
or U2984 (N_2984,N_1844,N_1273);
nand U2985 (N_2985,N_1682,N_1018);
nand U2986 (N_2986,N_1935,N_1155);
or U2987 (N_2987,N_1294,N_1452);
xnor U2988 (N_2988,N_1282,N_1055);
and U2989 (N_2989,N_1417,N_1235);
nand U2990 (N_2990,N_1312,N_1844);
xnor U2991 (N_2991,N_1021,N_1437);
nor U2992 (N_2992,N_1275,N_1768);
xnor U2993 (N_2993,N_1411,N_1043);
xnor U2994 (N_2994,N_1317,N_1189);
nand U2995 (N_2995,N_1723,N_1499);
and U2996 (N_2996,N_1295,N_1556);
nand U2997 (N_2997,N_1861,N_1954);
xnor U2998 (N_2998,N_1968,N_1910);
xnor U2999 (N_2999,N_1247,N_1665);
xor UO_0 (O_0,N_2486,N_2651);
xor UO_1 (O_1,N_2956,N_2169);
and UO_2 (O_2,N_2796,N_2825);
nand UO_3 (O_3,N_2023,N_2259);
and UO_4 (O_4,N_2219,N_2831);
nor UO_5 (O_5,N_2102,N_2257);
and UO_6 (O_6,N_2669,N_2276);
nand UO_7 (O_7,N_2474,N_2761);
nand UO_8 (O_8,N_2741,N_2821);
nand UO_9 (O_9,N_2898,N_2179);
xor UO_10 (O_10,N_2238,N_2093);
nand UO_11 (O_11,N_2841,N_2798);
nand UO_12 (O_12,N_2282,N_2658);
and UO_13 (O_13,N_2014,N_2333);
nand UO_14 (O_14,N_2777,N_2725);
nor UO_15 (O_15,N_2220,N_2789);
and UO_16 (O_16,N_2029,N_2211);
nand UO_17 (O_17,N_2968,N_2731);
or UO_18 (O_18,N_2690,N_2226);
nand UO_19 (O_19,N_2630,N_2908);
nor UO_20 (O_20,N_2168,N_2598);
xor UO_21 (O_21,N_2479,N_2755);
xnor UO_22 (O_22,N_2647,N_2255);
xor UO_23 (O_23,N_2171,N_2880);
xor UO_24 (O_24,N_2028,N_2445);
nor UO_25 (O_25,N_2573,N_2995);
nor UO_26 (O_26,N_2191,N_2672);
xnor UO_27 (O_27,N_2116,N_2495);
or UO_28 (O_28,N_2625,N_2585);
xnor UO_29 (O_29,N_2962,N_2991);
and UO_30 (O_30,N_2198,N_2779);
nand UO_31 (O_31,N_2158,N_2719);
and UO_32 (O_32,N_2215,N_2264);
or UO_33 (O_33,N_2832,N_2683);
nand UO_34 (O_34,N_2764,N_2792);
nor UO_35 (O_35,N_2590,N_2501);
and UO_36 (O_36,N_2963,N_2930);
nor UO_37 (O_37,N_2716,N_2917);
and UO_38 (O_38,N_2132,N_2843);
xnor UO_39 (O_39,N_2752,N_2315);
nand UO_40 (O_40,N_2600,N_2267);
nand UO_41 (O_41,N_2151,N_2355);
and UO_42 (O_42,N_2945,N_2136);
nor UO_43 (O_43,N_2039,N_2975);
nand UO_44 (O_44,N_2998,N_2915);
nand UO_45 (O_45,N_2582,N_2635);
xor UO_46 (O_46,N_2539,N_2130);
xor UO_47 (O_47,N_2839,N_2707);
nor UO_48 (O_48,N_2113,N_2738);
nand UO_49 (O_49,N_2071,N_2184);
nor UO_50 (O_50,N_2813,N_2531);
xor UO_51 (O_51,N_2966,N_2758);
nor UO_52 (O_52,N_2608,N_2393);
nor UO_53 (O_53,N_2233,N_2828);
and UO_54 (O_54,N_2440,N_2468);
xnor UO_55 (O_55,N_2567,N_2718);
nand UO_56 (O_56,N_2304,N_2229);
and UO_57 (O_57,N_2089,N_2555);
nor UO_58 (O_58,N_2463,N_2734);
and UO_59 (O_59,N_2147,N_2927);
or UO_60 (O_60,N_2404,N_2938);
nand UO_61 (O_61,N_2186,N_2854);
xor UO_62 (O_62,N_2162,N_2131);
nand UO_63 (O_63,N_2033,N_2302);
or UO_64 (O_64,N_2876,N_2408);
nor UO_65 (O_65,N_2227,N_2090);
and UO_66 (O_66,N_2403,N_2778);
nor UO_67 (O_67,N_2344,N_2324);
nand UO_68 (O_68,N_2096,N_2670);
and UO_69 (O_69,N_2218,N_2932);
or UO_70 (O_70,N_2252,N_2011);
xnor UO_71 (O_71,N_2989,N_2596);
nand UO_72 (O_72,N_2817,N_2526);
nand UO_73 (O_73,N_2981,N_2959);
nand UO_74 (O_74,N_2699,N_2894);
and UO_75 (O_75,N_2583,N_2756);
nand UO_76 (O_76,N_2307,N_2472);
and UO_77 (O_77,N_2978,N_2656);
and UO_78 (O_78,N_2139,N_2693);
or UO_79 (O_79,N_2339,N_2153);
and UO_80 (O_80,N_2711,N_2970);
or UO_81 (O_81,N_2618,N_2035);
or UO_82 (O_82,N_2691,N_2192);
or UO_83 (O_83,N_2747,N_2914);
or UO_84 (O_84,N_2824,N_2146);
and UO_85 (O_85,N_2059,N_2972);
xor UO_86 (O_86,N_2603,N_2353);
nor UO_87 (O_87,N_2613,N_2819);
nor UO_88 (O_88,N_2532,N_2230);
nand UO_89 (O_89,N_2465,N_2352);
nor UO_90 (O_90,N_2961,N_2543);
nor UO_91 (O_91,N_2835,N_2086);
nor UO_92 (O_92,N_2949,N_2503);
or UO_93 (O_93,N_2629,N_2743);
nand UO_94 (O_94,N_2614,N_2921);
and UO_95 (O_95,N_2510,N_2833);
nor UO_96 (O_96,N_2265,N_2006);
and UO_97 (O_97,N_2548,N_2997);
xnor UO_98 (O_98,N_2143,N_2977);
nor UO_99 (O_99,N_2247,N_2572);
nand UO_100 (O_100,N_2668,N_2281);
and UO_101 (O_101,N_2729,N_2581);
xor UO_102 (O_102,N_2263,N_2421);
or UO_103 (O_103,N_2072,N_2675);
nor UO_104 (O_104,N_2178,N_2291);
nand UO_105 (O_105,N_2564,N_2855);
and UO_106 (O_106,N_2366,N_2918);
and UO_107 (O_107,N_2783,N_2615);
or UO_108 (O_108,N_2957,N_2119);
nand UO_109 (O_109,N_2334,N_2507);
nand UO_110 (O_110,N_2622,N_2657);
or UO_111 (O_111,N_2273,N_2565);
nor UO_112 (O_112,N_2768,N_2958);
xor UO_113 (O_113,N_2266,N_2575);
or UO_114 (O_114,N_2815,N_2104);
xnor UO_115 (O_115,N_2073,N_2884);
or UO_116 (O_116,N_2239,N_2044);
nor UO_117 (O_117,N_2415,N_2636);
xor UO_118 (O_118,N_2713,N_2203);
xnor UO_119 (O_119,N_2368,N_2390);
xor UO_120 (O_120,N_2748,N_2053);
xor UO_121 (O_121,N_2142,N_2409);
xor UO_122 (O_122,N_2504,N_2292);
or UO_123 (O_123,N_2148,N_2015);
xor UO_124 (O_124,N_2907,N_2274);
nand UO_125 (O_125,N_2018,N_2494);
or UO_126 (O_126,N_2427,N_2433);
nand UO_127 (O_127,N_2173,N_2554);
nand UO_128 (O_128,N_2061,N_2296);
or UO_129 (O_129,N_2559,N_2974);
nand UO_130 (O_130,N_2881,N_2842);
xnor UO_131 (O_131,N_2781,N_2330);
and UO_132 (O_132,N_2458,N_2858);
and UO_133 (O_133,N_2709,N_2482);
and UO_134 (O_134,N_2380,N_2641);
nand UO_135 (O_135,N_2473,N_2485);
and UO_136 (O_136,N_2551,N_2346);
xnor UO_137 (O_137,N_2865,N_2523);
nand UO_138 (O_138,N_2318,N_2662);
nand UO_139 (O_139,N_2338,N_2275);
nor UO_140 (O_140,N_2735,N_2935);
xnor UO_141 (O_141,N_2607,N_2969);
xnor UO_142 (O_142,N_2475,N_2952);
xnor UO_143 (O_143,N_2899,N_2677);
or UO_144 (O_144,N_2386,N_2308);
nor UO_145 (O_145,N_2529,N_2224);
nor UO_146 (O_146,N_2426,N_2068);
nand UO_147 (O_147,N_2205,N_2785);
nand UO_148 (O_148,N_2425,N_2754);
nor UO_149 (O_149,N_2262,N_2003);
nor UO_150 (O_150,N_2384,N_2394);
nor UO_151 (O_151,N_2048,N_2484);
nor UO_152 (O_152,N_2721,N_2530);
nor UO_153 (O_153,N_2714,N_2175);
and UO_154 (O_154,N_2528,N_2850);
nor UO_155 (O_155,N_2395,N_2418);
or UO_156 (O_156,N_2517,N_2320);
nor UO_157 (O_157,N_2996,N_2505);
nor UO_158 (O_158,N_2558,N_2182);
or UO_159 (O_159,N_2289,N_2547);
nor UO_160 (O_160,N_2589,N_2836);
nand UO_161 (O_161,N_2631,N_2154);
nor UO_162 (O_162,N_2456,N_2696);
nor UO_163 (O_163,N_2114,N_2809);
and UO_164 (O_164,N_2818,N_2990);
nand UO_165 (O_165,N_2512,N_2419);
and UO_166 (O_166,N_2051,N_2370);
nor UO_167 (O_167,N_2212,N_2834);
nor UO_168 (O_168,N_2207,N_2665);
nor UO_169 (O_169,N_2109,N_2549);
xnor UO_170 (O_170,N_2478,N_2269);
nand UO_171 (O_171,N_2605,N_2084);
and UO_172 (O_172,N_2703,N_2736);
nor UO_173 (O_173,N_2432,N_2745);
and UO_174 (O_174,N_2070,N_2883);
xnor UO_175 (O_175,N_2595,N_2196);
and UO_176 (O_176,N_2038,N_2377);
and UO_177 (O_177,N_2032,N_2910);
nor UO_178 (O_178,N_2284,N_2381);
xnor UO_179 (O_179,N_2980,N_2939);
and UO_180 (O_180,N_2705,N_2452);
xor UO_181 (O_181,N_2137,N_2967);
or UO_182 (O_182,N_2621,N_2133);
and UO_183 (O_183,N_2776,N_2634);
nor UO_184 (O_184,N_2944,N_2112);
and UO_185 (O_185,N_2389,N_2365);
and UO_186 (O_186,N_2862,N_2763);
nand UO_187 (O_187,N_2410,N_2732);
nor UO_188 (O_188,N_2519,N_2050);
and UO_189 (O_189,N_2062,N_2101);
or UO_190 (O_190,N_2655,N_2724);
nor UO_191 (O_191,N_2864,N_2720);
xor UO_192 (O_192,N_2378,N_2188);
xnor UO_193 (O_193,N_2597,N_2242);
or UO_194 (O_194,N_2481,N_2319);
nand UO_195 (O_195,N_2678,N_2871);
nor UO_196 (O_196,N_2730,N_2128);
or UO_197 (O_197,N_2451,N_2666);
nor UO_198 (O_198,N_2054,N_2111);
nor UO_199 (O_199,N_2926,N_2744);
xnor UO_200 (O_200,N_2698,N_2087);
xnor UO_201 (O_201,N_2194,N_2727);
nor UO_202 (O_202,N_2513,N_2826);
or UO_203 (O_203,N_2217,N_2420);
or UO_204 (O_204,N_2213,N_2623);
nand UO_205 (O_205,N_2115,N_2337);
or UO_206 (O_206,N_2594,N_2870);
nand UO_207 (O_207,N_2775,N_2206);
and UO_208 (O_208,N_2953,N_2638);
and UO_209 (O_209,N_2249,N_2679);
and UO_210 (O_210,N_2012,N_2082);
nand UO_211 (O_211,N_2350,N_2568);
nor UO_212 (O_212,N_2470,N_2447);
and UO_213 (O_213,N_2435,N_2492);
nor UO_214 (O_214,N_2847,N_2922);
or UO_215 (O_215,N_2201,N_2804);
nand UO_216 (O_216,N_2022,N_2293);
or UO_217 (O_217,N_2579,N_2988);
nor UO_218 (O_218,N_2488,N_2243);
nor UO_219 (O_219,N_2013,N_2020);
and UO_220 (O_220,N_2611,N_2004);
or UO_221 (O_221,N_2288,N_2042);
nor UO_222 (O_222,N_2412,N_2376);
and UO_223 (O_223,N_2040,N_2477);
or UO_224 (O_224,N_2722,N_2661);
xor UO_225 (O_225,N_2385,N_2450);
nand UO_226 (O_226,N_2570,N_2144);
nand UO_227 (O_227,N_2872,N_2576);
nor UO_228 (O_228,N_2197,N_2041);
nor UO_229 (O_229,N_2449,N_2701);
or UO_230 (O_230,N_2692,N_2545);
nand UO_231 (O_231,N_2106,N_2637);
and UO_232 (O_232,N_2476,N_2000);
xnor UO_233 (O_233,N_2840,N_2626);
xnor UO_234 (O_234,N_2993,N_2016);
nand UO_235 (O_235,N_2897,N_2866);
and UO_236 (O_236,N_2397,N_2571);
nor UO_237 (O_237,N_2329,N_2500);
or UO_238 (O_238,N_2912,N_2909);
xnor UO_239 (O_239,N_2904,N_2103);
nand UO_240 (O_240,N_2309,N_2066);
nand UO_241 (O_241,N_2964,N_2578);
xor UO_242 (O_242,N_2373,N_2080);
or UO_243 (O_243,N_2214,N_2860);
or UO_244 (O_244,N_2960,N_2183);
or UO_245 (O_245,N_2587,N_2441);
or UO_246 (O_246,N_2717,N_2160);
nor UO_247 (O_247,N_2534,N_2660);
nor UO_248 (O_248,N_2108,N_2467);
nand UO_249 (O_249,N_2652,N_2896);
or UO_250 (O_250,N_2499,N_2359);
nor UO_251 (O_251,N_2047,N_2875);
xnor UO_252 (O_252,N_2976,N_2628);
xor UO_253 (O_253,N_2848,N_2455);
and UO_254 (O_254,N_2342,N_2535);
nor UO_255 (O_255,N_2135,N_2873);
or UO_256 (O_256,N_2762,N_2314);
or UO_257 (O_257,N_2712,N_2299);
nand UO_258 (O_258,N_2077,N_2123);
or UO_259 (O_259,N_2794,N_2514);
xnor UO_260 (O_260,N_2934,N_2877);
nor UO_261 (O_261,N_2195,N_2985);
nand UO_262 (O_262,N_2844,N_2820);
nor UO_263 (O_263,N_2055,N_2592);
or UO_264 (O_264,N_2074,N_2092);
and UO_265 (O_265,N_2868,N_2491);
nand UO_266 (O_266,N_2685,N_2317);
nand UO_267 (O_267,N_2673,N_2541);
xnor UO_268 (O_268,N_2795,N_2244);
or UO_269 (O_269,N_2994,N_2616);
and UO_270 (O_270,N_2766,N_2118);
or UO_271 (O_271,N_2936,N_2924);
or UO_272 (O_272,N_2327,N_2489);
and UO_273 (O_273,N_2867,N_2793);
nand UO_274 (O_274,N_2550,N_2733);
nor UO_275 (O_275,N_2246,N_2814);
xor UO_276 (O_276,N_2017,N_2105);
and UO_277 (O_277,N_2286,N_2790);
or UO_278 (O_278,N_2199,N_2094);
or UO_279 (O_279,N_2354,N_2973);
and UO_280 (O_280,N_2237,N_2399);
nand UO_281 (O_281,N_2697,N_2955);
or UO_282 (O_282,N_2913,N_2398);
and UO_283 (O_283,N_2401,N_2911);
and UO_284 (O_284,N_2010,N_2574);
or UO_285 (O_285,N_2297,N_2163);
and UO_286 (O_286,N_2326,N_2786);
nor UO_287 (O_287,N_2429,N_2434);
nand UO_288 (O_288,N_2279,N_2903);
nor UO_289 (O_289,N_2208,N_2391);
xor UO_290 (O_290,N_2671,N_2704);
and UO_291 (O_291,N_2822,N_2803);
or UO_292 (O_292,N_2174,N_2929);
nor UO_293 (O_293,N_2357,N_2599);
nand UO_294 (O_294,N_2537,N_2552);
nor UO_295 (O_295,N_2560,N_2740);
xor UO_296 (O_296,N_2680,N_2739);
or UO_297 (O_297,N_2648,N_2438);
and UO_298 (O_298,N_2088,N_2009);
and UO_299 (O_299,N_2428,N_2874);
and UO_300 (O_300,N_2802,N_2853);
nand UO_301 (O_301,N_2382,N_2954);
xnor UO_302 (O_302,N_2542,N_2210);
nor UO_303 (O_303,N_2430,N_2002);
or UO_304 (O_304,N_2193,N_2250);
nand UO_305 (O_305,N_2161,N_2928);
and UO_306 (O_306,N_2710,N_2480);
and UO_307 (O_307,N_2271,N_2863);
nand UO_308 (O_308,N_2882,N_2063);
xnor UO_309 (O_309,N_2125,N_2240);
nand UO_310 (O_310,N_2774,N_2525);
nand UO_311 (O_311,N_2138,N_2083);
nor UO_312 (O_312,N_2947,N_2800);
and UO_313 (O_313,N_2979,N_2462);
nand UO_314 (O_314,N_2852,N_2737);
nor UO_315 (O_315,N_2684,N_2402);
or UO_316 (O_316,N_2878,N_2971);
nand UO_317 (O_317,N_2037,N_2369);
or UO_318 (O_318,N_2640,N_2965);
or UO_319 (O_319,N_2190,N_2987);
nand UO_320 (O_320,N_2331,N_2005);
and UO_321 (O_321,N_2805,N_2335);
or UO_322 (O_322,N_2624,N_2157);
xor UO_323 (O_323,N_2659,N_2085);
or UO_324 (O_324,N_2388,N_2122);
and UO_325 (O_325,N_2437,N_2688);
and UO_326 (O_326,N_2602,N_2859);
and UO_327 (O_327,N_2466,N_2187);
nor UO_328 (O_328,N_2580,N_2838);
and UO_329 (O_329,N_2769,N_2782);
or UO_330 (O_330,N_2586,N_2770);
and UO_331 (O_331,N_2469,N_2577);
or UO_332 (O_332,N_2305,N_2170);
xor UO_333 (O_333,N_2007,N_2444);
nand UO_334 (O_334,N_2807,N_2164);
xor UO_335 (O_335,N_2019,N_2845);
xnor UO_336 (O_336,N_2411,N_2923);
or UO_337 (O_337,N_2806,N_2676);
nor UO_338 (O_338,N_2172,N_2516);
xnor UO_339 (O_339,N_2361,N_2436);
xnor UO_340 (O_340,N_2941,N_2290);
or UO_341 (O_341,N_2268,N_2498);
xor UO_342 (O_342,N_2540,N_2950);
or UO_343 (O_343,N_2837,N_2442);
and UO_344 (O_344,N_2221,N_2439);
xor UO_345 (O_345,N_2064,N_2356);
and UO_346 (O_346,N_2569,N_2645);
or UO_347 (O_347,N_2791,N_2323);
nor UO_348 (O_348,N_2627,N_2951);
or UO_349 (O_349,N_2021,N_2986);
or UO_350 (O_350,N_2700,N_2856);
nand UO_351 (O_351,N_2364,N_2067);
and UO_352 (O_352,N_2260,N_2076);
nor UO_353 (O_353,N_2490,N_2069);
nand UO_354 (O_354,N_2303,N_2746);
and UO_355 (O_355,N_2316,N_2509);
xnor UO_356 (O_356,N_2563,N_2689);
and UO_357 (O_357,N_2593,N_2827);
xnor UO_358 (O_358,N_2493,N_2277);
and UO_359 (O_359,N_2301,N_2036);
nand UO_360 (O_360,N_2245,N_2797);
and UO_361 (O_361,N_2008,N_2392);
and UO_362 (O_362,N_2508,N_2209);
nand UO_363 (O_363,N_2283,N_2632);
and UO_364 (O_364,N_2232,N_2052);
xor UO_365 (O_365,N_2294,N_2298);
or UO_366 (O_366,N_2236,N_2506);
or UO_367 (O_367,N_2150,N_2757);
or UO_368 (O_368,N_2256,N_2453);
xor UO_369 (O_369,N_2431,N_2533);
xnor UO_370 (O_370,N_2156,N_2780);
and UO_371 (O_371,N_2633,N_2422);
nor UO_372 (O_372,N_2515,N_2706);
xor UO_373 (O_373,N_2846,N_2177);
nor UO_374 (O_374,N_2141,N_2254);
nor UO_375 (O_375,N_2687,N_2120);
nand UO_376 (O_376,N_2321,N_2612);
xnor UO_377 (O_377,N_2332,N_2027);
nand UO_378 (O_378,N_2649,N_2235);
xnor UO_379 (O_379,N_2056,N_2134);
or UO_380 (O_380,N_2345,N_2124);
or UO_381 (O_381,N_2371,N_2916);
and UO_382 (O_382,N_2886,N_2423);
nor UO_383 (O_383,N_2992,N_2811);
xor UO_384 (O_384,N_2241,N_2751);
nor UO_385 (O_385,N_2372,N_2760);
nand UO_386 (O_386,N_2562,N_2667);
nor UO_387 (O_387,N_2749,N_2180);
nor UO_388 (O_388,N_2823,N_2620);
nor UO_389 (O_389,N_2272,N_2261);
nor UO_390 (O_390,N_2152,N_2176);
and UO_391 (O_391,N_2643,N_2584);
xnor UO_392 (O_392,N_2520,N_2400);
xor UO_393 (O_393,N_2065,N_2686);
xor UO_394 (O_394,N_2816,N_2216);
or UO_395 (O_395,N_2285,N_2617);
and UO_396 (O_396,N_2202,N_2695);
xor UO_397 (O_397,N_2937,N_2888);
nor UO_398 (O_398,N_2367,N_2057);
xnor UO_399 (O_399,N_2496,N_2906);
nand UO_400 (O_400,N_2715,N_2098);
and UO_401 (O_401,N_2374,N_2270);
or UO_402 (O_402,N_2681,N_2849);
xor UO_403 (O_403,N_2079,N_2225);
or UO_404 (O_404,N_2604,N_2772);
nand UO_405 (O_405,N_2879,N_2487);
or UO_406 (O_406,N_2248,N_2060);
nand UO_407 (O_407,N_2362,N_2166);
and UO_408 (O_408,N_2149,N_2081);
xor UO_409 (O_409,N_2251,N_2383);
or UO_410 (O_410,N_2295,N_2300);
xor UO_411 (O_411,N_2046,N_2925);
nand UO_412 (O_412,N_2043,N_2413);
nor UO_413 (O_413,N_2946,N_2905);
xor UO_414 (O_414,N_2129,N_2145);
nand UO_415 (O_415,N_2891,N_2810);
nor UO_416 (O_416,N_2030,N_2787);
xnor UO_417 (O_417,N_2322,N_2609);
nand UO_418 (O_418,N_2341,N_2702);
nor UO_419 (O_419,N_2121,N_2049);
nor UO_420 (O_420,N_2566,N_2097);
nand UO_421 (O_421,N_2726,N_2920);
nand UO_422 (O_422,N_2642,N_2471);
and UO_423 (O_423,N_2536,N_2117);
nand UO_424 (O_424,N_2728,N_2078);
nor UO_425 (O_425,N_2406,N_2885);
xor UO_426 (O_426,N_2258,N_2459);
and UO_427 (O_427,N_2784,N_2155);
nor UO_428 (O_428,N_2200,N_2887);
or UO_429 (O_429,N_2405,N_2424);
and UO_430 (O_430,N_2031,N_2464);
nand UO_431 (O_431,N_2663,N_2557);
nand UO_432 (O_432,N_2753,N_2387);
xnor UO_433 (O_433,N_2588,N_2561);
xnor UO_434 (O_434,N_2511,N_2773);
nand UO_435 (O_435,N_2765,N_2407);
nand UO_436 (O_436,N_2933,N_2253);
or UO_437 (O_437,N_2287,N_2610);
nor UO_438 (O_438,N_2140,N_2457);
nor UO_439 (O_439,N_2521,N_2460);
xnor UO_440 (O_440,N_2483,N_2278);
or UO_441 (O_441,N_2351,N_2723);
nand UO_442 (O_442,N_2556,N_2851);
or UO_443 (O_443,N_2416,N_2234);
or UO_444 (O_444,N_2461,N_2280);
nor UO_445 (O_445,N_2310,N_2646);
xnor UO_446 (O_446,N_2982,N_2553);
nand UO_447 (O_447,N_2034,N_2546);
nor UO_448 (O_448,N_2750,N_2808);
and UO_449 (O_449,N_2771,N_2983);
or UO_450 (O_450,N_2340,N_2375);
xnor UO_451 (O_451,N_2674,N_2812);
xor UO_452 (O_452,N_2204,N_2110);
and UO_453 (O_453,N_2830,N_2091);
nand UO_454 (O_454,N_2619,N_2518);
and UO_455 (O_455,N_2606,N_2095);
and UO_456 (O_456,N_2497,N_2448);
nor UO_457 (O_457,N_2892,N_2075);
nor UO_458 (O_458,N_2025,N_2167);
nand UO_459 (O_459,N_2664,N_2379);
and UO_460 (O_460,N_2396,N_2948);
nand UO_461 (O_461,N_2829,N_2524);
nand UO_462 (O_462,N_2919,N_2895);
nor UO_463 (O_463,N_2653,N_2999);
or UO_464 (O_464,N_2650,N_2889);
and UO_465 (O_465,N_2943,N_2328);
nor UO_466 (O_466,N_2024,N_2347);
or UO_467 (O_467,N_2502,N_2189);
or UO_468 (O_468,N_2544,N_2107);
xnor UO_469 (O_469,N_2311,N_2228);
and UO_470 (O_470,N_2185,N_2857);
and UO_471 (O_471,N_2126,N_2358);
nor UO_472 (O_472,N_2306,N_2165);
and UO_473 (O_473,N_2639,N_2313);
or UO_474 (O_474,N_2454,N_2654);
or UO_475 (O_475,N_2901,N_2893);
or UO_476 (O_476,N_2026,N_2001);
and UO_477 (O_477,N_2902,N_2742);
or UO_478 (O_478,N_2446,N_2538);
and UO_479 (O_479,N_2890,N_2527);
and UO_480 (O_480,N_2682,N_2349);
and UO_481 (O_481,N_2900,N_2127);
and UO_482 (O_482,N_2759,N_2591);
and UO_483 (O_483,N_2869,N_2931);
or UO_484 (O_484,N_2767,N_2861);
nand UO_485 (O_485,N_2360,N_2799);
and UO_486 (O_486,N_2336,N_2099);
or UO_487 (O_487,N_2181,N_2801);
or UO_488 (O_488,N_2058,N_2312);
nand UO_489 (O_489,N_2708,N_2363);
and UO_490 (O_490,N_2644,N_2159);
nand UO_491 (O_491,N_2045,N_2343);
nor UO_492 (O_492,N_2414,N_2601);
xor UO_493 (O_493,N_2788,N_2100);
or UO_494 (O_494,N_2222,N_2348);
nor UO_495 (O_495,N_2940,N_2984);
nand UO_496 (O_496,N_2231,N_2223);
or UO_497 (O_497,N_2522,N_2694);
nor UO_498 (O_498,N_2443,N_2942);
nand UO_499 (O_499,N_2325,N_2417);
endmodule