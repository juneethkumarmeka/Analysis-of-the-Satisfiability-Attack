module basic_1000_10000_1500_2_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5002,N_5003,N_5005,N_5006,N_5007,N_5009,N_5011,N_5012,N_5013,N_5015,N_5020,N_5021,N_5024,N_5025,N_5026,N_5029,N_5031,N_5033,N_5034,N_5039,N_5040,N_5041,N_5044,N_5046,N_5048,N_5049,N_5050,N_5052,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5061,N_5062,N_5064,N_5067,N_5068,N_5069,N_5070,N_5072,N_5074,N_5076,N_5077,N_5078,N_5079,N_5081,N_5082,N_5083,N_5084,N_5085,N_5088,N_5091,N_5092,N_5093,N_5096,N_5097,N_5099,N_5102,N_5104,N_5105,N_5106,N_5107,N_5108,N_5110,N_5111,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5122,N_5124,N_5127,N_5128,N_5129,N_5130,N_5137,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5147,N_5148,N_5150,N_5152,N_5155,N_5156,N_5157,N_5159,N_5160,N_5166,N_5169,N_5170,N_5171,N_5172,N_5173,N_5175,N_5176,N_5177,N_5179,N_5180,N_5181,N_5183,N_5184,N_5185,N_5189,N_5190,N_5191,N_5193,N_5194,N_5195,N_5197,N_5199,N_5203,N_5204,N_5205,N_5206,N_5208,N_5209,N_5210,N_5213,N_5214,N_5216,N_5217,N_5219,N_5221,N_5223,N_5224,N_5225,N_5226,N_5227,N_5230,N_5231,N_5232,N_5233,N_5235,N_5237,N_5238,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5250,N_5252,N_5253,N_5255,N_5257,N_5258,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5267,N_5268,N_5269,N_5271,N_5273,N_5274,N_5276,N_5278,N_5279,N_5280,N_5281,N_5283,N_5286,N_5289,N_5290,N_5292,N_5293,N_5294,N_5295,N_5296,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5307,N_5308,N_5309,N_5310,N_5315,N_5316,N_5319,N_5323,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5335,N_5336,N_5337,N_5339,N_5341,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5351,N_5353,N_5354,N_5357,N_5358,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5368,N_5369,N_5370,N_5372,N_5375,N_5376,N_5378,N_5381,N_5382,N_5383,N_5384,N_5386,N_5387,N_5392,N_5396,N_5398,N_5400,N_5402,N_5403,N_5404,N_5406,N_5408,N_5409,N_5410,N_5412,N_5413,N_5414,N_5415,N_5417,N_5418,N_5419,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5429,N_5431,N_5433,N_5434,N_5435,N_5436,N_5439,N_5440,N_5442,N_5444,N_5446,N_5447,N_5448,N_5449,N_5452,N_5454,N_5456,N_5457,N_5458,N_5459,N_5460,N_5462,N_5463,N_5464,N_5466,N_5467,N_5468,N_5469,N_5471,N_5475,N_5476,N_5477,N_5480,N_5481,N_5482,N_5483,N_5485,N_5487,N_5488,N_5489,N_5490,N_5491,N_5495,N_5496,N_5497,N_5498,N_5502,N_5503,N_5505,N_5506,N_5508,N_5511,N_5512,N_5515,N_5516,N_5517,N_5519,N_5522,N_5525,N_5528,N_5529,N_5530,N_5532,N_5533,N_5535,N_5540,N_5542,N_5544,N_5550,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5561,N_5563,N_5565,N_5566,N_5568,N_5570,N_5571,N_5576,N_5580,N_5581,N_5582,N_5583,N_5586,N_5588,N_5590,N_5593,N_5594,N_5595,N_5597,N_5600,N_5601,N_5603,N_5604,N_5605,N_5606,N_5607,N_5610,N_5612,N_5613,N_5614,N_5615,N_5618,N_5620,N_5623,N_5624,N_5626,N_5629,N_5630,N_5631,N_5632,N_5634,N_5635,N_5636,N_5637,N_5638,N_5640,N_5641,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5651,N_5652,N_5653,N_5655,N_5656,N_5658,N_5660,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5670,N_5671,N_5672,N_5675,N_5676,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5688,N_5690,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5703,N_5705,N_5706,N_5708,N_5709,N_5713,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5729,N_5732,N_5734,N_5739,N_5746,N_5747,N_5748,N_5749,N_5751,N_5753,N_5758,N_5759,N_5760,N_5761,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5775,N_5776,N_5777,N_5778,N_5779,N_5781,N_5782,N_5783,N_5786,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5799,N_5800,N_5801,N_5805,N_5808,N_5810,N_5813,N_5814,N_5815,N_5816,N_5817,N_5819,N_5821,N_5822,N_5824,N_5827,N_5828,N_5830,N_5831,N_5833,N_5834,N_5835,N_5836,N_5838,N_5840,N_5841,N_5845,N_5846,N_5850,N_5851,N_5852,N_5854,N_5856,N_5860,N_5861,N_5862,N_5863,N_5869,N_5870,N_5873,N_5874,N_5875,N_5877,N_5880,N_5881,N_5883,N_5885,N_5886,N_5887,N_5888,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5900,N_5902,N_5903,N_5905,N_5908,N_5909,N_5911,N_5913,N_5915,N_5921,N_5922,N_5923,N_5924,N_5926,N_5928,N_5931,N_5935,N_5936,N_5938,N_5939,N_5940,N_5941,N_5943,N_5944,N_5945,N_5946,N_5952,N_5954,N_5955,N_5956,N_5957,N_5959,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5971,N_5972,N_5974,N_5976,N_5977,N_5980,N_5981,N_5982,N_5983,N_5984,N_5986,N_5988,N_5990,N_5991,N_5993,N_5995,N_5996,N_6000,N_6003,N_6004,N_6005,N_6007,N_6009,N_6012,N_6013,N_6015,N_6018,N_6019,N_6020,N_6022,N_6024,N_6026,N_6027,N_6029,N_6032,N_6034,N_6035,N_6036,N_6037,N_6039,N_6040,N_6041,N_6043,N_6044,N_6047,N_6049,N_6050,N_6054,N_6056,N_6057,N_6059,N_6060,N_6061,N_6064,N_6065,N_6067,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6090,N_6091,N_6093,N_6095,N_6096,N_6097,N_6098,N_6100,N_6102,N_6103,N_6104,N_6106,N_6112,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6121,N_6122,N_6124,N_6125,N_6127,N_6128,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6142,N_6143,N_6145,N_6147,N_6148,N_6151,N_6155,N_6156,N_6158,N_6159,N_6160,N_6161,N_6166,N_6167,N_6168,N_6169,N_6173,N_6175,N_6176,N_6177,N_6183,N_6186,N_6187,N_6188,N_6189,N_6191,N_6192,N_6197,N_6198,N_6202,N_6203,N_6205,N_6206,N_6207,N_6209,N_6212,N_6213,N_6215,N_6218,N_6220,N_6222,N_6225,N_6226,N_6229,N_6230,N_6232,N_6233,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6243,N_6244,N_6246,N_6247,N_6249,N_6250,N_6252,N_6254,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6264,N_6265,N_6266,N_6267,N_6268,N_6270,N_6273,N_6276,N_6278,N_6280,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6302,N_6304,N_6306,N_6307,N_6309,N_6310,N_6311,N_6312,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6324,N_6325,N_6327,N_6328,N_6330,N_6331,N_6334,N_6338,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6356,N_6359,N_6360,N_6362,N_6363,N_6366,N_6367,N_6368,N_6370,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6379,N_6382,N_6383,N_6386,N_6388,N_6393,N_6395,N_6396,N_6398,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6414,N_6416,N_6417,N_6418,N_6420,N_6421,N_6424,N_6425,N_6426,N_6427,N_6428,N_6430,N_6434,N_6436,N_6438,N_6439,N_6441,N_6442,N_6443,N_6444,N_6446,N_6447,N_6450,N_6452,N_6453,N_6455,N_6456,N_6458,N_6459,N_6461,N_6462,N_6464,N_6465,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6477,N_6478,N_6481,N_6482,N_6483,N_6487,N_6488,N_6490,N_6491,N_6494,N_6495,N_6497,N_6498,N_6500,N_6501,N_6502,N_6504,N_6505,N_6506,N_6507,N_6509,N_6512,N_6514,N_6516,N_6519,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6534,N_6537,N_6542,N_6543,N_6544,N_6545,N_6550,N_6551,N_6555,N_6556,N_6557,N_6560,N_6561,N_6562,N_6564,N_6568,N_6570,N_6573,N_6574,N_6575,N_6576,N_6577,N_6580,N_6581,N_6582,N_6587,N_6590,N_6592,N_6593,N_6594,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6618,N_6621,N_6622,N_6625,N_6627,N_6628,N_6629,N_6630,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6646,N_6647,N_6648,N_6649,N_6652,N_6654,N_6656,N_6659,N_6662,N_6664,N_6665,N_6669,N_6670,N_6671,N_6672,N_6675,N_6676,N_6677,N_6679,N_6682,N_6683,N_6684,N_6685,N_6686,N_6688,N_6690,N_6691,N_6693,N_6695,N_6696,N_6698,N_6699,N_6700,N_6703,N_6704,N_6705,N_6706,N_6709,N_6711,N_6712,N_6713,N_6715,N_6716,N_6718,N_6719,N_6720,N_6721,N_6723,N_6725,N_6727,N_6730,N_6732,N_6733,N_6735,N_6737,N_6738,N_6740,N_6745,N_6747,N_6748,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6766,N_6768,N_6772,N_6773,N_6774,N_6775,N_6777,N_6778,N_6779,N_6780,N_6782,N_6783,N_6785,N_6787,N_6789,N_6791,N_6793,N_6794,N_6797,N_6798,N_6799,N_6801,N_6802,N_6803,N_6804,N_6805,N_6808,N_6809,N_6810,N_6812,N_6813,N_6814,N_6816,N_6818,N_6820,N_6821,N_6823,N_6824,N_6825,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6837,N_6838,N_6841,N_6843,N_6847,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6858,N_6859,N_6862,N_6863,N_6864,N_6865,N_6866,N_6868,N_6870,N_6873,N_6874,N_6875,N_6876,N_6878,N_6887,N_6888,N_6891,N_6892,N_6893,N_6895,N_6896,N_6900,N_6901,N_6904,N_6906,N_6907,N_6909,N_6913,N_6914,N_6916,N_6917,N_6919,N_6920,N_6922,N_6923,N_6926,N_6927,N_6928,N_6929,N_6933,N_6934,N_6935,N_6936,N_6939,N_6941,N_6945,N_6947,N_6948,N_6949,N_6951,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6972,N_6974,N_6976,N_6977,N_6978,N_6979,N_6982,N_6983,N_6984,N_6986,N_6989,N_6994,N_6996,N_6997,N_7000,N_7001,N_7003,N_7004,N_7006,N_7007,N_7009,N_7010,N_7011,N_7012,N_7016,N_7023,N_7024,N_7025,N_7026,N_7028,N_7029,N_7032,N_7037,N_7038,N_7041,N_7042,N_7044,N_7045,N_7047,N_7048,N_7050,N_7051,N_7052,N_7053,N_7054,N_7057,N_7059,N_7060,N_7061,N_7062,N_7063,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7079,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7091,N_7092,N_7094,N_7095,N_7096,N_7097,N_7099,N_7100,N_7102,N_7103,N_7104,N_7105,N_7109,N_7110,N_7111,N_7113,N_7114,N_7116,N_7117,N_7118,N_7119,N_7121,N_7122,N_7123,N_7124,N_7127,N_7128,N_7129,N_7130,N_7132,N_7133,N_7134,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7143,N_7145,N_7146,N_7149,N_7150,N_7153,N_7154,N_7156,N_7161,N_7162,N_7163,N_7164,N_7165,N_7167,N_7168,N_7169,N_7171,N_7172,N_7173,N_7175,N_7176,N_7179,N_7181,N_7182,N_7183,N_7185,N_7186,N_7187,N_7188,N_7190,N_7191,N_7192,N_7195,N_7196,N_7197,N_7198,N_7204,N_7205,N_7209,N_7210,N_7211,N_7214,N_7215,N_7216,N_7218,N_7219,N_7222,N_7223,N_7224,N_7225,N_7227,N_7228,N_7229,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7241,N_7242,N_7243,N_7244,N_7246,N_7247,N_7248,N_7249,N_7250,N_7252,N_7253,N_7254,N_7256,N_7258,N_7259,N_7260,N_7261,N_7264,N_7265,N_7266,N_7267,N_7269,N_7271,N_7273,N_7276,N_7278,N_7281,N_7282,N_7283,N_7284,N_7285,N_7288,N_7289,N_7290,N_7293,N_7294,N_7296,N_7298,N_7299,N_7303,N_7304,N_7305,N_7306,N_7307,N_7310,N_7311,N_7312,N_7313,N_7315,N_7317,N_7318,N_7319,N_7320,N_7322,N_7323,N_7325,N_7326,N_7331,N_7333,N_7334,N_7335,N_7336,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7352,N_7354,N_7358,N_7360,N_7361,N_7362,N_7363,N_7365,N_7366,N_7367,N_7371,N_7372,N_7373,N_7374,N_7375,N_7379,N_7380,N_7383,N_7385,N_7386,N_7388,N_7389,N_7390,N_7392,N_7393,N_7394,N_7396,N_7397,N_7398,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7415,N_7418,N_7420,N_7424,N_7425,N_7426,N_7427,N_7429,N_7430,N_7433,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7443,N_7445,N_7448,N_7449,N_7450,N_7452,N_7453,N_7454,N_7456,N_7457,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7466,N_7469,N_7471,N_7472,N_7473,N_7474,N_7476,N_7479,N_7480,N_7482,N_7486,N_7488,N_7490,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7501,N_7502,N_7506,N_7507,N_7508,N_7509,N_7511,N_7517,N_7520,N_7521,N_7522,N_7523,N_7527,N_7529,N_7532,N_7534,N_7535,N_7536,N_7539,N_7541,N_7543,N_7545,N_7547,N_7548,N_7549,N_7550,N_7551,N_7553,N_7555,N_7558,N_7560,N_7561,N_7563,N_7564,N_7565,N_7566,N_7567,N_7570,N_7571,N_7575,N_7576,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7590,N_7592,N_7593,N_7594,N_7595,N_7596,N_7598,N_7599,N_7600,N_7601,N_7603,N_7604,N_7605,N_7606,N_7608,N_7609,N_7610,N_7611,N_7614,N_7617,N_7618,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7628,N_7633,N_7636,N_7637,N_7639,N_7640,N_7641,N_7642,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7653,N_7654,N_7655,N_7656,N_7659,N_7660,N_7661,N_7662,N_7667,N_7668,N_7669,N_7671,N_7672,N_7673,N_7674,N_7677,N_7679,N_7681,N_7682,N_7683,N_7684,N_7686,N_7687,N_7688,N_7692,N_7696,N_7697,N_7699,N_7700,N_7701,N_7702,N_7707,N_7708,N_7709,N_7710,N_7711,N_7713,N_7714,N_7715,N_7717,N_7718,N_7719,N_7720,N_7724,N_7728,N_7729,N_7732,N_7734,N_7738,N_7740,N_7742,N_7743,N_7744,N_7747,N_7748,N_7749,N_7751,N_7754,N_7755,N_7757,N_7758,N_7759,N_7761,N_7765,N_7769,N_7770,N_7772,N_7775,N_7776,N_7779,N_7782,N_7783,N_7788,N_7790,N_7793,N_7794,N_7795,N_7796,N_7798,N_7799,N_7801,N_7802,N_7803,N_7805,N_7806,N_7807,N_7809,N_7810,N_7811,N_7812,N_7814,N_7815,N_7822,N_7826,N_7827,N_7829,N_7830,N_7831,N_7833,N_7835,N_7836,N_7837,N_7838,N_7839,N_7841,N_7842,N_7843,N_7846,N_7848,N_7852,N_7853,N_7854,N_7855,N_7861,N_7863,N_7864,N_7865,N_7866,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7876,N_7877,N_7879,N_7880,N_7881,N_7883,N_7885,N_7886,N_7887,N_7889,N_7892,N_7893,N_7894,N_7895,N_7896,N_7898,N_7901,N_7902,N_7904,N_7905,N_7911,N_7912,N_7915,N_7916,N_7919,N_7920,N_7921,N_7922,N_7923,N_7925,N_7926,N_7927,N_7928,N_7932,N_7933,N_7935,N_7942,N_7948,N_7949,N_7950,N_7952,N_7953,N_7957,N_7958,N_7961,N_7962,N_7965,N_7970,N_7972,N_7973,N_7974,N_7975,N_7978,N_7982,N_7983,N_7984,N_7986,N_7987,N_7988,N_7989,N_7990,N_7994,N_7995,N_8000,N_8003,N_8004,N_8005,N_8007,N_8009,N_8010,N_8011,N_8013,N_8014,N_8015,N_8016,N_8018,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8028,N_8029,N_8030,N_8032,N_8033,N_8035,N_8041,N_8044,N_8046,N_8049,N_8051,N_8052,N_8053,N_8054,N_8056,N_8057,N_8061,N_8062,N_8064,N_8065,N_8068,N_8072,N_8074,N_8075,N_8076,N_8078,N_8081,N_8082,N_8083,N_8085,N_8087,N_8090,N_8092,N_8093,N_8094,N_8095,N_8096,N_8099,N_8100,N_8102,N_8103,N_8107,N_8108,N_8109,N_8110,N_8113,N_8114,N_8115,N_8117,N_8121,N_8122,N_8123,N_8124,N_8128,N_8130,N_8131,N_8132,N_8133,N_8135,N_8136,N_8137,N_8138,N_8140,N_8141,N_8142,N_8143,N_8149,N_8150,N_8154,N_8155,N_8158,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8169,N_8170,N_8171,N_8172,N_8175,N_8177,N_8178,N_8180,N_8181,N_8182,N_8184,N_8185,N_8186,N_8189,N_8190,N_8191,N_8192,N_8194,N_8196,N_8197,N_8198,N_8200,N_8201,N_8202,N_8203,N_8205,N_8207,N_8210,N_8211,N_8214,N_8215,N_8217,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8226,N_8227,N_8229,N_8231,N_8232,N_8233,N_8237,N_8241,N_8243,N_8244,N_8245,N_8249,N_8251,N_8252,N_8254,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8263,N_8265,N_8266,N_8267,N_8268,N_8269,N_8271,N_8278,N_8279,N_8280,N_8282,N_8285,N_8286,N_8288,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8314,N_8319,N_8321,N_8322,N_8323,N_8324,N_8326,N_8327,N_8329,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8338,N_8339,N_8341,N_8342,N_8344,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8362,N_8364,N_8365,N_8366,N_8367,N_8368,N_8371,N_8372,N_8374,N_8375,N_8377,N_8379,N_8380,N_8381,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8390,N_8391,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8402,N_8403,N_8405,N_8406,N_8407,N_8408,N_8409,N_8413,N_8414,N_8415,N_8416,N_8418,N_8419,N_8423,N_8426,N_8427,N_8428,N_8429,N_8430,N_8432,N_8434,N_8436,N_8437,N_8438,N_8439,N_8442,N_8444,N_8445,N_8446,N_8447,N_8449,N_8451,N_8452,N_8453,N_8454,N_8455,N_8457,N_8459,N_8465,N_8466,N_8469,N_8474,N_8475,N_8476,N_8478,N_8479,N_8480,N_8484,N_8485,N_8486,N_8487,N_8489,N_8491,N_8492,N_8493,N_8494,N_8495,N_8497,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8507,N_8508,N_8509,N_8511,N_8512,N_8513,N_8514,N_8515,N_8517,N_8519,N_8522,N_8526,N_8528,N_8529,N_8530,N_8532,N_8533,N_8535,N_8536,N_8537,N_8540,N_8543,N_8544,N_8545,N_8547,N_8548,N_8549,N_8550,N_8552,N_8553,N_8554,N_8556,N_8557,N_8559,N_8561,N_8562,N_8563,N_8565,N_8566,N_8568,N_8572,N_8574,N_8575,N_8576,N_8577,N_8578,N_8580,N_8581,N_8582,N_8585,N_8587,N_8588,N_8590,N_8591,N_8594,N_8595,N_8596,N_8597,N_8599,N_8600,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8610,N_8611,N_8612,N_8613,N_8617,N_8618,N_8619,N_8621,N_8623,N_8624,N_8627,N_8628,N_8630,N_8631,N_8634,N_8636,N_8639,N_8640,N_8642,N_8644,N_8645,N_8646,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8656,N_8658,N_8659,N_8660,N_8662,N_8663,N_8666,N_8667,N_8670,N_8672,N_8673,N_8674,N_8675,N_8677,N_8678,N_8682,N_8684,N_8688,N_8689,N_8691,N_8692,N_8696,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8706,N_8708,N_8709,N_8710,N_8712,N_8713,N_8714,N_8716,N_8717,N_8719,N_8720,N_8721,N_8722,N_8724,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8733,N_8736,N_8737,N_8738,N_8740,N_8744,N_8746,N_8747,N_8748,N_8749,N_8750,N_8752,N_8753,N_8755,N_8757,N_8758,N_8761,N_8762,N_8763,N_8765,N_8772,N_8773,N_8777,N_8779,N_8781,N_8782,N_8785,N_8786,N_8789,N_8791,N_8793,N_8794,N_8796,N_8797,N_8798,N_8799,N_8801,N_8802,N_8804,N_8806,N_8807,N_8808,N_8809,N_8810,N_8813,N_8814,N_8815,N_8817,N_8821,N_8822,N_8823,N_8824,N_8825,N_8827,N_8829,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8840,N_8842,N_8843,N_8846,N_8847,N_8848,N_8851,N_8852,N_8853,N_8855,N_8857,N_8861,N_8864,N_8867,N_8868,N_8869,N_8872,N_8874,N_8875,N_8876,N_8877,N_8879,N_8880,N_8881,N_8884,N_8889,N_8890,N_8894,N_8897,N_8898,N_8899,N_8900,N_8901,N_8904,N_8907,N_8908,N_8909,N_8910,N_8912,N_8913,N_8914,N_8915,N_8919,N_8920,N_8922,N_8924,N_8925,N_8926,N_8928,N_8929,N_8931,N_8932,N_8933,N_8934,N_8935,N_8939,N_8940,N_8941,N_8942,N_8944,N_8946,N_8947,N_8950,N_8953,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8963,N_8966,N_8967,N_8970,N_8975,N_8979,N_8980,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8993,N_8994,N_8995,N_8996,N_8999,N_9000,N_9001,N_9002,N_9004,N_9005,N_9006,N_9007,N_9008,N_9011,N_9012,N_9014,N_9016,N_9017,N_9020,N_9021,N_9022,N_9024,N_9025,N_9026,N_9027,N_9029,N_9030,N_9033,N_9034,N_9036,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9047,N_9048,N_9049,N_9050,N_9053,N_9056,N_9058,N_9060,N_9061,N_9062,N_9063,N_9065,N_9066,N_9067,N_9068,N_9071,N_9074,N_9077,N_9078,N_9082,N_9084,N_9085,N_9088,N_9089,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9104,N_9106,N_9107,N_9108,N_9110,N_9112,N_9116,N_9117,N_9118,N_9119,N_9120,N_9125,N_9127,N_9128,N_9129,N_9132,N_9133,N_9134,N_9138,N_9139,N_9140,N_9141,N_9142,N_9144,N_9145,N_9146,N_9148,N_9151,N_9156,N_9157,N_9158,N_9162,N_9164,N_9165,N_9169,N_9172,N_9173,N_9174,N_9175,N_9177,N_9178,N_9180,N_9181,N_9183,N_9186,N_9188,N_9190,N_9191,N_9194,N_9195,N_9196,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9205,N_9206,N_9208,N_9209,N_9210,N_9211,N_9218,N_9219,N_9220,N_9224,N_9226,N_9227,N_9228,N_9231,N_9233,N_9234,N_9235,N_9237,N_9238,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9249,N_9250,N_9251,N_9252,N_9255,N_9256,N_9258,N_9260,N_9261,N_9264,N_9265,N_9267,N_9271,N_9272,N_9273,N_9274,N_9277,N_9280,N_9281,N_9282,N_9286,N_9287,N_9289,N_9293,N_9294,N_9297,N_9298,N_9299,N_9300,N_9301,N_9304,N_9307,N_9308,N_9311,N_9312,N_9317,N_9321,N_9322,N_9323,N_9326,N_9327,N_9328,N_9329,N_9332,N_9336,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9353,N_9354,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9370,N_9372,N_9373,N_9375,N_9376,N_9378,N_9379,N_9381,N_9382,N_9383,N_9385,N_9386,N_9390,N_9392,N_9393,N_9394,N_9396,N_9397,N_9400,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9409,N_9412,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9425,N_9427,N_9428,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9440,N_9441,N_9443,N_9445,N_9447,N_9448,N_9450,N_9451,N_9453,N_9457,N_9458,N_9459,N_9461,N_9463,N_9464,N_9465,N_9466,N_9467,N_9470,N_9471,N_9474,N_9475,N_9476,N_9477,N_9478,N_9483,N_9484,N_9485,N_9487,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9504,N_9506,N_9507,N_9510,N_9511,N_9513,N_9515,N_9516,N_9519,N_9520,N_9521,N_9523,N_9524,N_9526,N_9528,N_9531,N_9532,N_9533,N_9534,N_9536,N_9538,N_9539,N_9540,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9557,N_9559,N_9560,N_9564,N_9565,N_9566,N_9567,N_9568,N_9570,N_9572,N_9573,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9596,N_9597,N_9598,N_9601,N_9602,N_9605,N_9606,N_9607,N_9609,N_9611,N_9613,N_9614,N_9616,N_9619,N_9621,N_9623,N_9624,N_9627,N_9630,N_9631,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9652,N_9653,N_9655,N_9656,N_9657,N_9660,N_9661,N_9662,N_9664,N_9665,N_9666,N_9668,N_9671,N_9673,N_9675,N_9676,N_9677,N_9681,N_9682,N_9684,N_9686,N_9688,N_9689,N_9690,N_9692,N_9693,N_9696,N_9700,N_9703,N_9704,N_9705,N_9706,N_9707,N_9709,N_9713,N_9714,N_9716,N_9717,N_9719,N_9721,N_9724,N_9726,N_9727,N_9728,N_9730,N_9733,N_9734,N_9735,N_9737,N_9742,N_9743,N_9745,N_9746,N_9747,N_9751,N_9753,N_9754,N_9755,N_9756,N_9759,N_9762,N_9765,N_9766,N_9768,N_9770,N_9771,N_9772,N_9773,N_9777,N_9779,N_9783,N_9784,N_9785,N_9792,N_9797,N_9799,N_9800,N_9801,N_9805,N_9806,N_9809,N_9811,N_9813,N_9814,N_9816,N_9817,N_9818,N_9820,N_9821,N_9822,N_9823,N_9825,N_9828,N_9829,N_9832,N_9834,N_9835,N_9836,N_9837,N_9839,N_9841,N_9843,N_9844,N_9846,N_9847,N_9848,N_9849,N_9850,N_9852,N_9853,N_9854,N_9855,N_9857,N_9858,N_9859,N_9862,N_9864,N_9865,N_9868,N_9869,N_9870,N_9873,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9884,N_9888,N_9890,N_9891,N_9892,N_9893,N_9895,N_9896,N_9898,N_9899,N_9901,N_9906,N_9907,N_9909,N_9911,N_9913,N_9914,N_9915,N_9918,N_9919,N_9923,N_9924,N_9925,N_9926,N_9929,N_9930,N_9931,N_9932,N_9933,N_9935,N_9937,N_9938,N_9939,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9951,N_9952,N_9953,N_9955,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9965,N_9968,N_9971,N_9973,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9986,N_9987,N_9988,N_9992,N_9993,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_162,In_509);
xor U1 (N_1,In_885,In_186);
nand U2 (N_2,In_198,In_2);
xnor U3 (N_3,In_788,In_612);
xnor U4 (N_4,In_38,In_778);
xnor U5 (N_5,In_481,In_622);
or U6 (N_6,In_127,In_707);
or U7 (N_7,In_72,In_56);
nand U8 (N_8,In_295,In_462);
and U9 (N_9,In_582,In_3);
xnor U10 (N_10,In_351,In_113);
xor U11 (N_11,In_114,In_247);
xnor U12 (N_12,In_650,In_841);
xor U13 (N_13,In_663,In_907);
or U14 (N_14,In_790,In_855);
nor U15 (N_15,In_456,In_294);
or U16 (N_16,In_987,In_196);
xnor U17 (N_17,In_697,In_20);
nor U18 (N_18,In_129,In_146);
nand U19 (N_19,In_434,In_416);
nand U20 (N_20,In_506,In_637);
or U21 (N_21,In_608,In_693);
xor U22 (N_22,In_976,In_802);
and U23 (N_23,In_255,In_537);
or U24 (N_24,In_237,In_32);
and U25 (N_25,In_743,In_552);
or U26 (N_26,In_577,In_111);
nor U27 (N_27,In_95,In_651);
nand U28 (N_28,In_494,In_503);
and U29 (N_29,In_123,In_380);
xor U30 (N_30,In_632,In_732);
nand U31 (N_31,In_935,In_309);
xnor U32 (N_32,In_461,In_65);
nor U33 (N_33,In_614,In_924);
nor U34 (N_34,In_776,In_31);
nand U35 (N_35,In_216,In_915);
nand U36 (N_36,In_433,In_562);
or U37 (N_37,In_925,In_635);
or U38 (N_38,In_920,In_643);
or U39 (N_39,In_593,In_808);
and U40 (N_40,In_476,In_46);
xnor U41 (N_41,In_443,In_540);
and U42 (N_42,In_278,In_902);
nand U43 (N_43,In_618,In_735);
xnor U44 (N_44,In_166,In_190);
nor U45 (N_45,In_159,In_345);
and U46 (N_46,In_490,In_656);
xnor U47 (N_47,In_686,In_662);
nand U48 (N_48,In_567,In_45);
and U49 (N_49,In_394,In_704);
and U50 (N_50,In_795,In_664);
and U51 (N_51,In_318,In_944);
nand U52 (N_52,In_22,In_782);
nand U53 (N_53,In_457,In_926);
nor U54 (N_54,In_279,In_884);
nor U55 (N_55,In_763,In_454);
and U56 (N_56,In_785,In_269);
nand U57 (N_57,In_135,In_496);
nor U58 (N_58,In_984,In_600);
and U59 (N_59,In_212,In_605);
nand U60 (N_60,In_718,In_849);
nor U61 (N_61,In_224,In_557);
xor U62 (N_62,In_177,In_969);
xor U63 (N_63,In_765,In_185);
xnor U64 (N_64,In_33,In_100);
nand U65 (N_65,In_522,In_489);
and U66 (N_66,In_681,In_909);
nand U67 (N_67,In_303,In_938);
xnor U68 (N_68,In_187,In_756);
nand U69 (N_69,In_375,In_329);
and U70 (N_70,In_19,In_420);
or U71 (N_71,In_170,In_304);
xnor U72 (N_72,In_603,In_449);
nand U73 (N_73,In_535,In_682);
nor U74 (N_74,In_985,In_52);
nand U75 (N_75,In_575,In_759);
nor U76 (N_76,In_228,In_695);
xor U77 (N_77,In_996,In_30);
nand U78 (N_78,In_912,In_940);
nand U79 (N_79,In_820,In_429);
and U80 (N_80,In_721,In_534);
nor U81 (N_81,In_426,In_812);
nor U82 (N_82,In_698,In_836);
or U83 (N_83,In_583,In_156);
nor U84 (N_84,In_236,In_871);
nand U85 (N_85,In_405,In_395);
xor U86 (N_86,In_641,In_222);
nor U87 (N_87,In_565,In_447);
or U88 (N_88,In_676,In_179);
nor U89 (N_89,In_148,In_524);
or U90 (N_90,In_708,In_860);
xor U91 (N_91,In_754,In_898);
and U92 (N_92,In_208,In_328);
nor U93 (N_93,In_629,In_644);
nor U94 (N_94,In_119,In_571);
nor U95 (N_95,In_78,In_850);
xnor U96 (N_96,In_197,In_734);
xnor U97 (N_97,In_899,In_687);
or U98 (N_98,In_134,In_206);
nor U99 (N_99,In_966,In_263);
xnor U100 (N_100,In_178,In_417);
nand U101 (N_101,In_492,In_117);
nand U102 (N_102,In_144,In_515);
nand U103 (N_103,In_883,In_964);
or U104 (N_104,In_872,In_427);
nor U105 (N_105,In_740,In_947);
and U106 (N_106,In_357,In_918);
nor U107 (N_107,In_742,In_432);
and U108 (N_108,In_955,In_320);
nor U109 (N_109,In_268,In_630);
and U110 (N_110,In_659,In_911);
or U111 (N_111,In_54,In_865);
and U112 (N_112,In_974,In_202);
nor U113 (N_113,In_770,In_448);
nor U114 (N_114,In_63,In_726);
and U115 (N_115,In_81,In_842);
or U116 (N_116,In_767,In_978);
and U117 (N_117,In_786,In_339);
nor U118 (N_118,In_270,In_98);
nor U119 (N_119,In_719,In_195);
or U120 (N_120,In_981,In_35);
or U121 (N_121,In_973,In_758);
nor U122 (N_122,In_946,In_407);
nor U123 (N_123,In_590,In_660);
nand U124 (N_124,In_486,In_837);
nand U125 (N_125,In_933,In_150);
xnor U126 (N_126,In_610,In_455);
nand U127 (N_127,In_402,In_854);
xor U128 (N_128,In_10,In_326);
and U129 (N_129,In_665,In_59);
xor U130 (N_130,In_891,In_922);
or U131 (N_131,In_826,In_276);
and U132 (N_132,In_999,In_231);
and U133 (N_133,In_904,In_741);
xnor U134 (N_134,In_755,In_798);
xor U135 (N_135,In_516,In_58);
and U136 (N_136,In_53,In_163);
xnor U137 (N_137,In_803,In_67);
nand U138 (N_138,In_383,In_669);
xor U139 (N_139,In_672,In_221);
xor U140 (N_140,In_281,In_404);
nand U141 (N_141,In_893,In_239);
or U142 (N_142,In_513,In_886);
nand U143 (N_143,In_832,In_439);
nand U144 (N_144,In_271,In_40);
xnor U145 (N_145,In_949,In_988);
xor U146 (N_146,In_518,In_50);
and U147 (N_147,In_131,In_241);
nor U148 (N_148,In_772,In_725);
nand U149 (N_149,In_471,In_728);
xnor U150 (N_150,In_624,In_596);
nor U151 (N_151,In_360,In_792);
nand U152 (N_152,In_544,In_235);
nand U153 (N_153,In_602,In_723);
xor U154 (N_154,In_61,In_232);
and U155 (N_155,In_678,In_809);
or U156 (N_156,In_415,In_777);
or U157 (N_157,In_959,In_253);
xnor U158 (N_158,In_8,In_274);
or U159 (N_159,In_108,In_149);
nand U160 (N_160,In_892,In_807);
nand U161 (N_161,In_342,In_673);
xor U162 (N_162,In_962,In_843);
nor U163 (N_163,In_352,In_376);
xnor U164 (N_164,In_474,In_386);
nand U165 (N_165,In_161,In_227);
or U166 (N_166,In_485,In_675);
nand U167 (N_167,In_667,In_140);
or U168 (N_168,In_514,In_688);
nor U169 (N_169,In_536,In_958);
nand U170 (N_170,In_573,In_153);
and U171 (N_171,In_184,In_0);
and U172 (N_172,In_287,In_469);
nor U173 (N_173,In_685,In_240);
nor U174 (N_174,In_219,In_753);
and U175 (N_175,In_9,In_746);
nor U176 (N_176,In_312,In_7);
or U177 (N_177,In_257,In_314);
and U178 (N_178,In_505,In_873);
or U179 (N_179,In_530,In_181);
or U180 (N_180,In_679,In_680);
or U181 (N_181,In_406,In_211);
xnor U182 (N_182,In_588,In_289);
or U183 (N_183,In_254,In_69);
nand U184 (N_184,In_623,In_830);
nand U185 (N_185,In_835,In_256);
xor U186 (N_186,In_613,In_482);
nor U187 (N_187,In_397,In_929);
and U188 (N_188,In_442,In_878);
and U189 (N_189,In_852,In_388);
and U190 (N_190,In_863,In_817);
nand U191 (N_191,In_639,In_79);
xnor U192 (N_192,In_880,In_501);
or U193 (N_193,In_994,In_599);
nor U194 (N_194,In_587,In_561);
nand U195 (N_195,In_607,In_259);
nor U196 (N_196,In_604,In_344);
nor U197 (N_197,In_658,In_337);
xor U198 (N_198,In_497,In_652);
nor U199 (N_199,In_244,In_191);
and U200 (N_200,In_422,In_645);
nor U201 (N_201,In_617,In_99);
nand U202 (N_202,In_960,In_372);
xnor U203 (N_203,In_327,In_220);
nand U204 (N_204,In_277,In_369);
and U205 (N_205,In_34,In_288);
nor U206 (N_206,In_945,In_701);
nor U207 (N_207,In_670,In_889);
nand U208 (N_208,In_47,In_74);
or U209 (N_209,In_390,In_616);
nand U210 (N_210,In_97,In_138);
and U211 (N_211,In_581,In_176);
and U212 (N_212,In_273,In_814);
nor U213 (N_213,In_174,In_297);
or U214 (N_214,In_125,In_18);
and U215 (N_215,In_5,In_91);
or U216 (N_216,In_638,In_619);
and U217 (N_217,In_655,In_818);
and U218 (N_218,In_779,In_750);
xor U219 (N_219,In_261,In_167);
xor U220 (N_220,In_316,In_706);
nor U221 (N_221,In_943,In_82);
xor U222 (N_222,In_296,In_49);
or U223 (N_223,In_175,In_549);
nor U224 (N_224,In_789,In_6);
nor U225 (N_225,In_711,In_311);
nand U226 (N_226,In_106,In_868);
or U227 (N_227,In_80,In_477);
or U228 (N_228,In_410,In_358);
nand U229 (N_229,In_346,In_931);
xnor U230 (N_230,In_242,In_661);
and U231 (N_231,In_142,In_188);
xor U232 (N_232,In_411,In_745);
xor U233 (N_233,In_139,In_511);
xor U234 (N_234,In_396,In_528);
xnor U235 (N_235,In_887,In_363);
and U236 (N_236,In_862,In_570);
and U237 (N_237,In_709,In_264);
nor U238 (N_238,In_951,In_169);
or U239 (N_239,In_507,In_995);
and U240 (N_240,In_229,In_724);
or U241 (N_241,In_475,In_611);
nand U242 (N_242,In_594,In_574);
and U243 (N_243,In_260,In_94);
nor U244 (N_244,In_234,In_634);
nand U245 (N_245,In_677,In_737);
and U246 (N_246,In_601,In_165);
xnor U247 (N_247,In_425,In_452);
xnor U248 (N_248,In_546,In_251);
or U249 (N_249,In_356,In_648);
xnor U250 (N_250,In_822,In_160);
nor U251 (N_251,In_293,In_298);
nand U252 (N_252,In_334,In_824);
and U253 (N_253,In_285,In_823);
nor U254 (N_254,In_838,In_858);
nand U255 (N_255,In_831,In_580);
nor U256 (N_256,In_730,In_751);
nor U257 (N_257,In_980,In_547);
and U258 (N_258,In_903,In_896);
and U259 (N_259,In_781,In_428);
xor U260 (N_260,In_834,In_464);
and U261 (N_261,In_523,In_401);
xor U262 (N_262,In_15,In_403);
nand U263 (N_263,In_983,In_136);
nor U264 (N_264,In_440,In_102);
nor U265 (N_265,In_280,In_498);
nor U266 (N_266,In_952,In_816);
xor U267 (N_267,In_705,In_615);
nand U268 (N_268,In_488,In_101);
and U269 (N_269,In_654,In_459);
nand U270 (N_270,In_313,In_716);
or U271 (N_271,In_73,In_76);
nor U272 (N_272,In_888,In_867);
and U273 (N_273,In_200,In_180);
or U274 (N_274,In_783,In_870);
nor U275 (N_275,In_90,In_364);
nor U276 (N_276,In_172,In_928);
or U277 (N_277,In_700,In_545);
or U278 (N_278,In_609,In_936);
nand U279 (N_279,In_963,In_93);
nor U280 (N_280,In_466,In_393);
nor U281 (N_281,In_225,In_265);
xnor U282 (N_282,In_121,In_155);
xnor U283 (N_283,In_720,In_764);
or U284 (N_284,In_541,In_133);
nor U285 (N_285,In_747,In_950);
nor U286 (N_286,In_866,In_532);
and U287 (N_287,In_591,In_444);
or U288 (N_288,In_463,In_894);
nor U289 (N_289,In_302,In_927);
nor U290 (N_290,In_733,In_727);
nor U291 (N_291,In_631,In_189);
nand U292 (N_292,In_436,In_961);
xnor U293 (N_293,In_453,In_939);
xnor U294 (N_294,In_301,In_173);
and U295 (N_295,In_17,In_702);
and U296 (N_296,In_578,In_649);
nand U297 (N_297,In_520,In_209);
nand U298 (N_298,In_306,In_762);
nand U299 (N_299,In_768,In_16);
nand U300 (N_300,In_62,In_744);
nor U301 (N_301,In_563,In_692);
or U302 (N_302,In_122,In_840);
or U303 (N_303,In_343,In_282);
xnor U304 (N_304,In_671,In_585);
or U305 (N_305,In_527,In_479);
xor U306 (N_306,In_4,In_458);
xnor U307 (N_307,In_771,In_627);
or U308 (N_308,In_666,In_684);
nor U309 (N_309,In_472,In_572);
or U310 (N_310,In_24,In_699);
xnor U311 (N_311,In_749,In_598);
nand U312 (N_312,In_584,In_908);
and U313 (N_313,In_86,In_991);
nor U314 (N_314,In_731,In_215);
nand U315 (N_315,In_857,In_874);
nor U316 (N_316,In_330,In_853);
or U317 (N_317,In_48,In_194);
xor U318 (N_318,In_223,In_780);
xor U319 (N_319,In_333,In_606);
xor U320 (N_320,In_531,In_761);
nand U321 (N_321,In_468,In_27);
nand U322 (N_322,In_154,In_272);
xnor U323 (N_323,In_968,In_451);
nor U324 (N_324,In_266,In_130);
xor U325 (N_325,In_152,In_145);
and U326 (N_326,In_512,In_900);
nor U327 (N_327,In_491,In_207);
nor U328 (N_328,In_92,In_819);
or U329 (N_329,In_193,In_729);
or U330 (N_330,In_797,In_923);
and U331 (N_331,In_362,In_151);
and U332 (N_332,In_470,In_934);
or U333 (N_333,In_322,In_794);
nor U334 (N_334,In_799,In_847);
nand U335 (N_335,In_942,In_977);
or U336 (N_336,In_460,In_529);
nand U337 (N_337,In_954,In_877);
xnor U338 (N_338,In_307,In_539);
and U339 (N_339,In_483,In_14);
xnor U340 (N_340,In_965,In_210);
or U341 (N_341,In_331,In_290);
and U342 (N_342,In_787,In_332);
nor U343 (N_343,In_238,In_398);
nor U344 (N_344,In_864,In_249);
or U345 (N_345,In_876,In_41);
xor U346 (N_346,In_89,In_217);
xor U347 (N_347,In_784,In_431);
and U348 (N_348,In_11,In_29);
xnor U349 (N_349,In_203,In_245);
xnor U350 (N_350,In_226,In_848);
or U351 (N_351,In_810,In_930);
nor U352 (N_352,In_646,In_748);
nand U353 (N_353,In_275,In_109);
or U354 (N_354,In_205,In_694);
xor U355 (N_355,In_418,In_502);
or U356 (N_356,In_553,In_164);
and U357 (N_357,In_478,In_589);
nand U358 (N_358,In_430,In_910);
nand U359 (N_359,In_710,In_104);
xor U360 (N_360,In_495,In_901);
xnor U361 (N_361,In_657,In_424);
nand U362 (N_362,In_806,In_391);
nand U363 (N_363,In_120,In_218);
nand U364 (N_364,In_250,In_653);
nor U365 (N_365,In_246,In_696);
and U366 (N_366,In_308,In_538);
and U367 (N_367,In_284,In_989);
nand U368 (N_368,In_559,In_465);
nor U369 (N_369,In_44,In_42);
nand U370 (N_370,In_993,In_569);
nor U371 (N_371,In_480,In_856);
xor U372 (N_372,In_445,In_201);
nand U373 (N_373,In_508,In_592);
xor U374 (N_374,In_997,In_674);
nor U375 (N_375,In_689,In_640);
or U376 (N_376,In_917,In_714);
nand U377 (N_377,In_752,In_568);
or U378 (N_378,In_126,In_57);
and U379 (N_379,In_365,In_551);
or U380 (N_380,In_839,In_875);
and U381 (N_381,In_555,In_642);
xnor U382 (N_382,In_213,In_595);
or U383 (N_383,In_37,In_628);
nor U384 (N_384,In_116,In_804);
nor U385 (N_385,In_336,In_636);
or U386 (N_386,In_811,In_982);
and U387 (N_387,In_846,In_370);
or U388 (N_388,In_319,In_967);
nor U389 (N_389,In_906,In_387);
nor U390 (N_390,In_813,In_542);
nor U391 (N_391,In_828,In_199);
xnor U392 (N_392,In_77,In_132);
or U393 (N_393,In_550,In_377);
xnor U394 (N_394,In_739,In_521);
nand U395 (N_395,In_341,In_510);
nor U396 (N_396,In_554,In_315);
nor U397 (N_397,In_408,In_349);
nand U398 (N_398,In_992,In_438);
nor U399 (N_399,In_283,In_413);
and U400 (N_400,In_441,In_805);
or U401 (N_401,In_399,In_353);
xor U402 (N_402,In_325,In_183);
and U403 (N_403,In_558,In_374);
and U404 (N_404,In_1,In_712);
xnor U405 (N_405,In_367,In_300);
xnor U406 (N_406,In_378,In_21);
and U407 (N_407,In_171,In_919);
nand U408 (N_408,In_347,In_948);
nand U409 (N_409,In_791,In_467);
and U410 (N_410,In_586,In_499);
or U411 (N_411,In_833,In_321);
or U412 (N_412,In_621,In_350);
xor U413 (N_413,In_310,In_446);
nand U414 (N_414,In_392,In_233);
and U415 (N_415,In_112,In_158);
and U416 (N_416,In_774,In_827);
xor U417 (N_417,In_703,In_533);
and U418 (N_418,In_103,In_286);
nand U419 (N_419,In_147,In_317);
xnor U420 (N_420,In_579,In_26);
nor U421 (N_421,In_389,In_690);
and U422 (N_422,In_971,In_916);
or U423 (N_423,In_576,In_400);
nor U424 (N_424,In_775,In_55);
or U425 (N_425,In_423,In_39);
xor U426 (N_426,In_597,In_937);
nor U427 (N_427,In_861,In_548);
nand U428 (N_428,In_487,In_85);
and U429 (N_429,In_970,In_525);
or U430 (N_430,In_115,In_738);
nand U431 (N_431,In_473,In_986);
or U432 (N_432,In_182,In_157);
nor U433 (N_433,In_291,In_879);
or U434 (N_434,In_248,In_760);
xnor U435 (N_435,In_437,In_230);
and U436 (N_436,In_825,In_36);
xor U437 (N_437,In_715,In_371);
and U438 (N_438,In_801,In_414);
xnor U439 (N_439,In_373,In_60);
or U440 (N_440,In_564,In_668);
or U441 (N_441,In_626,In_88);
or U442 (N_442,In_168,In_897);
xnor U443 (N_443,In_381,In_543);
or U444 (N_444,In_13,In_348);
xor U445 (N_445,In_869,In_829);
nor U446 (N_446,In_204,In_335);
nor U447 (N_447,In_137,In_258);
nor U448 (N_448,In_299,In_815);
nor U449 (N_449,In_267,In_379);
or U450 (N_450,In_66,In_214);
or U451 (N_451,In_107,In_262);
and U452 (N_452,In_647,In_713);
nand U453 (N_453,In_324,In_105);
nand U454 (N_454,In_800,In_796);
and U455 (N_455,In_368,In_517);
xnor U456 (N_456,In_354,In_355);
or U457 (N_457,In_359,In_83);
or U458 (N_458,In_450,In_717);
xor U459 (N_459,In_70,In_736);
nor U460 (N_460,In_504,In_292);
or U461 (N_461,In_914,In_252);
xnor U462 (N_462,In_124,In_773);
and U463 (N_463,In_128,In_998);
or U464 (N_464,In_382,In_882);
and U465 (N_465,In_972,In_691);
nand U466 (N_466,In_881,In_23);
or U467 (N_467,In_941,In_519);
nand U468 (N_468,In_366,In_560);
nor U469 (N_469,In_921,In_722);
xor U470 (N_470,In_566,In_956);
and U471 (N_471,In_769,In_323);
and U472 (N_472,In_75,In_84);
nor U473 (N_473,In_757,In_953);
or U474 (N_474,In_851,In_143);
and U475 (N_475,In_338,In_385);
and U476 (N_476,In_384,In_419);
or U477 (N_477,In_932,In_361);
and U478 (N_478,In_110,In_890);
and U479 (N_479,In_957,In_913);
xor U480 (N_480,In_412,In_68);
and U481 (N_481,In_64,In_500);
nor U482 (N_482,In_633,In_859);
or U483 (N_483,In_141,In_620);
and U484 (N_484,In_793,In_975);
nand U485 (N_485,In_895,In_192);
xnor U486 (N_486,In_28,In_305);
nand U487 (N_487,In_625,In_421);
and U488 (N_488,In_43,In_340);
and U489 (N_489,In_905,In_683);
xor U490 (N_490,In_96,In_71);
xnor U491 (N_491,In_51,In_493);
xor U492 (N_492,In_526,In_821);
xor U493 (N_493,In_844,In_979);
and U494 (N_494,In_484,In_556);
xor U495 (N_495,In_243,In_118);
nand U496 (N_496,In_25,In_409);
xor U497 (N_497,In_766,In_990);
or U498 (N_498,In_12,In_87);
nand U499 (N_499,In_845,In_435);
nor U500 (N_500,In_642,In_781);
nand U501 (N_501,In_421,In_642);
xor U502 (N_502,In_315,In_430);
and U503 (N_503,In_492,In_845);
xnor U504 (N_504,In_350,In_190);
nand U505 (N_505,In_104,In_804);
xor U506 (N_506,In_482,In_852);
nand U507 (N_507,In_653,In_824);
and U508 (N_508,In_801,In_646);
xnor U509 (N_509,In_909,In_376);
xor U510 (N_510,In_527,In_128);
or U511 (N_511,In_740,In_93);
nand U512 (N_512,In_410,In_281);
or U513 (N_513,In_728,In_299);
xnor U514 (N_514,In_94,In_689);
nor U515 (N_515,In_865,In_676);
nand U516 (N_516,In_233,In_821);
xnor U517 (N_517,In_581,In_253);
nand U518 (N_518,In_780,In_171);
or U519 (N_519,In_715,In_757);
or U520 (N_520,In_680,In_272);
nand U521 (N_521,In_465,In_941);
and U522 (N_522,In_30,In_157);
or U523 (N_523,In_11,In_517);
or U524 (N_524,In_964,In_875);
nor U525 (N_525,In_901,In_466);
xnor U526 (N_526,In_378,In_44);
or U527 (N_527,In_634,In_332);
or U528 (N_528,In_754,In_694);
and U529 (N_529,In_924,In_280);
nor U530 (N_530,In_701,In_465);
and U531 (N_531,In_100,In_468);
or U532 (N_532,In_789,In_176);
xor U533 (N_533,In_382,In_912);
xnor U534 (N_534,In_804,In_86);
nand U535 (N_535,In_277,In_574);
or U536 (N_536,In_286,In_929);
and U537 (N_537,In_324,In_919);
nand U538 (N_538,In_967,In_696);
xor U539 (N_539,In_615,In_994);
or U540 (N_540,In_664,In_374);
nand U541 (N_541,In_746,In_872);
nand U542 (N_542,In_531,In_703);
or U543 (N_543,In_740,In_364);
or U544 (N_544,In_805,In_204);
and U545 (N_545,In_691,In_284);
and U546 (N_546,In_553,In_632);
nor U547 (N_547,In_382,In_355);
and U548 (N_548,In_524,In_159);
nand U549 (N_549,In_745,In_515);
and U550 (N_550,In_295,In_647);
nor U551 (N_551,In_498,In_852);
nand U552 (N_552,In_147,In_268);
xor U553 (N_553,In_822,In_171);
and U554 (N_554,In_807,In_211);
and U555 (N_555,In_145,In_559);
nand U556 (N_556,In_499,In_308);
or U557 (N_557,In_925,In_46);
or U558 (N_558,In_461,In_11);
nand U559 (N_559,In_846,In_982);
and U560 (N_560,In_998,In_210);
nor U561 (N_561,In_470,In_707);
or U562 (N_562,In_387,In_22);
nor U563 (N_563,In_656,In_593);
or U564 (N_564,In_192,In_145);
nand U565 (N_565,In_125,In_915);
nand U566 (N_566,In_469,In_900);
nand U567 (N_567,In_992,In_457);
nand U568 (N_568,In_345,In_315);
xor U569 (N_569,In_566,In_969);
nand U570 (N_570,In_758,In_451);
and U571 (N_571,In_617,In_573);
and U572 (N_572,In_10,In_253);
and U573 (N_573,In_390,In_179);
and U574 (N_574,In_83,In_917);
xor U575 (N_575,In_797,In_4);
and U576 (N_576,In_394,In_227);
nor U577 (N_577,In_961,In_286);
nor U578 (N_578,In_991,In_613);
nand U579 (N_579,In_258,In_602);
nor U580 (N_580,In_836,In_18);
or U581 (N_581,In_399,In_939);
nand U582 (N_582,In_626,In_874);
xor U583 (N_583,In_52,In_359);
nor U584 (N_584,In_294,In_748);
and U585 (N_585,In_324,In_266);
and U586 (N_586,In_890,In_261);
and U587 (N_587,In_607,In_336);
xnor U588 (N_588,In_991,In_810);
nand U589 (N_589,In_131,In_546);
nor U590 (N_590,In_989,In_937);
and U591 (N_591,In_413,In_198);
nand U592 (N_592,In_659,In_804);
xnor U593 (N_593,In_907,In_757);
nand U594 (N_594,In_781,In_65);
or U595 (N_595,In_895,In_704);
or U596 (N_596,In_755,In_369);
and U597 (N_597,In_822,In_688);
and U598 (N_598,In_822,In_133);
xnor U599 (N_599,In_720,In_599);
or U600 (N_600,In_789,In_461);
nand U601 (N_601,In_37,In_229);
and U602 (N_602,In_945,In_357);
xor U603 (N_603,In_156,In_358);
nor U604 (N_604,In_904,In_649);
nand U605 (N_605,In_108,In_33);
or U606 (N_606,In_947,In_658);
nor U607 (N_607,In_739,In_254);
nor U608 (N_608,In_797,In_462);
and U609 (N_609,In_707,In_302);
xnor U610 (N_610,In_592,In_31);
xnor U611 (N_611,In_18,In_918);
nand U612 (N_612,In_441,In_782);
and U613 (N_613,In_482,In_955);
nor U614 (N_614,In_160,In_721);
and U615 (N_615,In_889,In_689);
and U616 (N_616,In_774,In_130);
xor U617 (N_617,In_383,In_614);
or U618 (N_618,In_173,In_285);
nand U619 (N_619,In_431,In_906);
and U620 (N_620,In_569,In_669);
and U621 (N_621,In_694,In_981);
nand U622 (N_622,In_209,In_514);
xnor U623 (N_623,In_495,In_355);
nand U624 (N_624,In_111,In_278);
xnor U625 (N_625,In_196,In_586);
or U626 (N_626,In_585,In_153);
and U627 (N_627,In_122,In_213);
xor U628 (N_628,In_760,In_25);
or U629 (N_629,In_949,In_648);
xor U630 (N_630,In_521,In_947);
nand U631 (N_631,In_974,In_430);
and U632 (N_632,In_780,In_992);
xor U633 (N_633,In_162,In_99);
nand U634 (N_634,In_985,In_189);
or U635 (N_635,In_128,In_340);
nand U636 (N_636,In_472,In_450);
nor U637 (N_637,In_530,In_87);
or U638 (N_638,In_456,In_577);
nor U639 (N_639,In_928,In_968);
nor U640 (N_640,In_992,In_856);
xnor U641 (N_641,In_361,In_458);
and U642 (N_642,In_130,In_818);
and U643 (N_643,In_811,In_552);
nor U644 (N_644,In_24,In_990);
xor U645 (N_645,In_556,In_983);
nand U646 (N_646,In_700,In_82);
nand U647 (N_647,In_269,In_12);
nand U648 (N_648,In_618,In_220);
and U649 (N_649,In_775,In_52);
nand U650 (N_650,In_184,In_582);
xor U651 (N_651,In_41,In_472);
or U652 (N_652,In_45,In_655);
xor U653 (N_653,In_363,In_918);
xor U654 (N_654,In_74,In_929);
or U655 (N_655,In_955,In_933);
and U656 (N_656,In_174,In_548);
nor U657 (N_657,In_75,In_748);
nor U658 (N_658,In_611,In_379);
xnor U659 (N_659,In_488,In_770);
and U660 (N_660,In_582,In_547);
or U661 (N_661,In_455,In_817);
nor U662 (N_662,In_638,In_602);
nor U663 (N_663,In_882,In_338);
nor U664 (N_664,In_930,In_284);
xor U665 (N_665,In_65,In_930);
xor U666 (N_666,In_408,In_62);
xor U667 (N_667,In_629,In_532);
or U668 (N_668,In_500,In_893);
nor U669 (N_669,In_183,In_456);
and U670 (N_670,In_583,In_553);
nor U671 (N_671,In_267,In_438);
nand U672 (N_672,In_481,In_185);
nand U673 (N_673,In_827,In_239);
xnor U674 (N_674,In_518,In_919);
nand U675 (N_675,In_802,In_700);
xnor U676 (N_676,In_282,In_274);
nand U677 (N_677,In_123,In_940);
or U678 (N_678,In_739,In_987);
nand U679 (N_679,In_605,In_582);
nand U680 (N_680,In_620,In_401);
nor U681 (N_681,In_31,In_154);
nand U682 (N_682,In_4,In_317);
nand U683 (N_683,In_78,In_225);
or U684 (N_684,In_36,In_777);
nand U685 (N_685,In_979,In_591);
nand U686 (N_686,In_416,In_326);
nor U687 (N_687,In_447,In_90);
nor U688 (N_688,In_854,In_535);
or U689 (N_689,In_292,In_572);
xor U690 (N_690,In_392,In_562);
and U691 (N_691,In_912,In_877);
and U692 (N_692,In_95,In_374);
and U693 (N_693,In_656,In_574);
nor U694 (N_694,In_525,In_198);
nor U695 (N_695,In_379,In_932);
and U696 (N_696,In_235,In_112);
or U697 (N_697,In_440,In_396);
nor U698 (N_698,In_764,In_765);
and U699 (N_699,In_201,In_537);
nand U700 (N_700,In_147,In_924);
and U701 (N_701,In_751,In_649);
and U702 (N_702,In_947,In_794);
or U703 (N_703,In_681,In_515);
xor U704 (N_704,In_780,In_253);
and U705 (N_705,In_326,In_164);
nor U706 (N_706,In_295,In_824);
nor U707 (N_707,In_899,In_47);
nand U708 (N_708,In_21,In_792);
or U709 (N_709,In_835,In_444);
nor U710 (N_710,In_79,In_35);
xor U711 (N_711,In_18,In_715);
or U712 (N_712,In_410,In_599);
and U713 (N_713,In_918,In_286);
nand U714 (N_714,In_508,In_699);
and U715 (N_715,In_907,In_512);
nor U716 (N_716,In_655,In_896);
and U717 (N_717,In_921,In_784);
nand U718 (N_718,In_332,In_419);
nand U719 (N_719,In_539,In_645);
nor U720 (N_720,In_434,In_102);
or U721 (N_721,In_244,In_176);
and U722 (N_722,In_386,In_23);
xor U723 (N_723,In_364,In_273);
or U724 (N_724,In_393,In_162);
and U725 (N_725,In_577,In_302);
or U726 (N_726,In_459,In_620);
nand U727 (N_727,In_636,In_285);
nor U728 (N_728,In_994,In_334);
nor U729 (N_729,In_445,In_51);
and U730 (N_730,In_510,In_286);
and U731 (N_731,In_304,In_19);
nand U732 (N_732,In_292,In_419);
and U733 (N_733,In_878,In_385);
nor U734 (N_734,In_456,In_160);
nand U735 (N_735,In_422,In_888);
and U736 (N_736,In_264,In_284);
or U737 (N_737,In_781,In_124);
xnor U738 (N_738,In_243,In_604);
and U739 (N_739,In_966,In_290);
or U740 (N_740,In_641,In_972);
xor U741 (N_741,In_564,In_5);
xnor U742 (N_742,In_982,In_672);
and U743 (N_743,In_268,In_830);
nand U744 (N_744,In_533,In_792);
xnor U745 (N_745,In_595,In_235);
nor U746 (N_746,In_137,In_403);
xor U747 (N_747,In_32,In_81);
and U748 (N_748,In_322,In_943);
nor U749 (N_749,In_319,In_496);
or U750 (N_750,In_306,In_838);
nand U751 (N_751,In_259,In_341);
nand U752 (N_752,In_486,In_399);
nand U753 (N_753,In_117,In_494);
nor U754 (N_754,In_807,In_187);
and U755 (N_755,In_199,In_181);
nor U756 (N_756,In_483,In_559);
nor U757 (N_757,In_427,In_692);
xnor U758 (N_758,In_475,In_556);
or U759 (N_759,In_598,In_408);
and U760 (N_760,In_155,In_401);
and U761 (N_761,In_608,In_127);
xnor U762 (N_762,In_305,In_656);
xnor U763 (N_763,In_377,In_445);
nor U764 (N_764,In_184,In_110);
or U765 (N_765,In_477,In_778);
and U766 (N_766,In_573,In_9);
nand U767 (N_767,In_701,In_169);
or U768 (N_768,In_8,In_778);
nor U769 (N_769,In_827,In_619);
nand U770 (N_770,In_535,In_577);
or U771 (N_771,In_826,In_138);
xor U772 (N_772,In_992,In_313);
or U773 (N_773,In_220,In_907);
or U774 (N_774,In_127,In_451);
nand U775 (N_775,In_147,In_113);
or U776 (N_776,In_984,In_521);
and U777 (N_777,In_326,In_49);
xor U778 (N_778,In_390,In_880);
or U779 (N_779,In_974,In_268);
or U780 (N_780,In_289,In_84);
and U781 (N_781,In_521,In_818);
nor U782 (N_782,In_817,In_564);
or U783 (N_783,In_762,In_849);
xnor U784 (N_784,In_933,In_210);
nor U785 (N_785,In_370,In_620);
nand U786 (N_786,In_497,In_601);
or U787 (N_787,In_281,In_776);
or U788 (N_788,In_181,In_762);
nor U789 (N_789,In_426,In_620);
nand U790 (N_790,In_308,In_171);
and U791 (N_791,In_751,In_181);
and U792 (N_792,In_487,In_922);
or U793 (N_793,In_437,In_441);
and U794 (N_794,In_654,In_806);
nand U795 (N_795,In_509,In_512);
or U796 (N_796,In_92,In_567);
or U797 (N_797,In_649,In_281);
nand U798 (N_798,In_260,In_760);
or U799 (N_799,In_828,In_90);
or U800 (N_800,In_804,In_779);
nand U801 (N_801,In_28,In_358);
nand U802 (N_802,In_975,In_920);
nor U803 (N_803,In_933,In_932);
or U804 (N_804,In_692,In_962);
xor U805 (N_805,In_66,In_476);
nor U806 (N_806,In_420,In_559);
xnor U807 (N_807,In_61,In_188);
or U808 (N_808,In_57,In_818);
or U809 (N_809,In_395,In_380);
nor U810 (N_810,In_328,In_640);
nor U811 (N_811,In_519,In_983);
and U812 (N_812,In_952,In_551);
and U813 (N_813,In_502,In_365);
or U814 (N_814,In_370,In_853);
and U815 (N_815,In_161,In_60);
nand U816 (N_816,In_985,In_839);
xnor U817 (N_817,In_521,In_157);
or U818 (N_818,In_104,In_248);
xor U819 (N_819,In_812,In_429);
or U820 (N_820,In_607,In_185);
xor U821 (N_821,In_107,In_869);
or U822 (N_822,In_468,In_377);
and U823 (N_823,In_145,In_156);
nor U824 (N_824,In_820,In_246);
and U825 (N_825,In_674,In_225);
or U826 (N_826,In_993,In_738);
nor U827 (N_827,In_862,In_222);
nor U828 (N_828,In_163,In_502);
or U829 (N_829,In_492,In_379);
xnor U830 (N_830,In_624,In_748);
and U831 (N_831,In_204,In_119);
or U832 (N_832,In_906,In_641);
or U833 (N_833,In_17,In_65);
and U834 (N_834,In_594,In_58);
and U835 (N_835,In_739,In_713);
nand U836 (N_836,In_159,In_876);
nor U837 (N_837,In_406,In_480);
and U838 (N_838,In_736,In_211);
nor U839 (N_839,In_727,In_242);
and U840 (N_840,In_389,In_569);
xor U841 (N_841,In_993,In_174);
nor U842 (N_842,In_482,In_591);
xor U843 (N_843,In_194,In_26);
or U844 (N_844,In_176,In_35);
nor U845 (N_845,In_340,In_276);
or U846 (N_846,In_825,In_922);
nor U847 (N_847,In_953,In_71);
xnor U848 (N_848,In_896,In_847);
xnor U849 (N_849,In_698,In_89);
xor U850 (N_850,In_721,In_729);
or U851 (N_851,In_893,In_722);
xor U852 (N_852,In_52,In_335);
or U853 (N_853,In_798,In_511);
or U854 (N_854,In_916,In_725);
nor U855 (N_855,In_474,In_855);
or U856 (N_856,In_662,In_567);
and U857 (N_857,In_203,In_14);
nand U858 (N_858,In_575,In_216);
or U859 (N_859,In_187,In_423);
and U860 (N_860,In_171,In_395);
nor U861 (N_861,In_988,In_575);
nor U862 (N_862,In_843,In_929);
nand U863 (N_863,In_29,In_982);
nor U864 (N_864,In_546,In_617);
or U865 (N_865,In_797,In_706);
nor U866 (N_866,In_930,In_266);
nor U867 (N_867,In_254,In_386);
and U868 (N_868,In_48,In_751);
xnor U869 (N_869,In_382,In_602);
nand U870 (N_870,In_601,In_636);
or U871 (N_871,In_432,In_656);
nand U872 (N_872,In_400,In_307);
nand U873 (N_873,In_51,In_505);
xnor U874 (N_874,In_809,In_932);
nand U875 (N_875,In_879,In_312);
or U876 (N_876,In_497,In_647);
nand U877 (N_877,In_192,In_874);
xor U878 (N_878,In_553,In_287);
or U879 (N_879,In_126,In_318);
nor U880 (N_880,In_225,In_779);
nor U881 (N_881,In_506,In_25);
nand U882 (N_882,In_503,In_127);
nand U883 (N_883,In_392,In_584);
nand U884 (N_884,In_675,In_191);
nand U885 (N_885,In_296,In_477);
xor U886 (N_886,In_180,In_322);
and U887 (N_887,In_583,In_82);
or U888 (N_888,In_242,In_190);
nand U889 (N_889,In_951,In_145);
nor U890 (N_890,In_177,In_220);
and U891 (N_891,In_869,In_635);
or U892 (N_892,In_252,In_113);
nand U893 (N_893,In_115,In_213);
xor U894 (N_894,In_617,In_614);
and U895 (N_895,In_151,In_70);
or U896 (N_896,In_423,In_981);
xnor U897 (N_897,In_843,In_544);
xnor U898 (N_898,In_99,In_326);
and U899 (N_899,In_892,In_74);
or U900 (N_900,In_665,In_905);
and U901 (N_901,In_452,In_5);
xor U902 (N_902,In_469,In_485);
or U903 (N_903,In_209,In_148);
nand U904 (N_904,In_757,In_974);
nand U905 (N_905,In_252,In_917);
xor U906 (N_906,In_306,In_468);
or U907 (N_907,In_119,In_713);
xnor U908 (N_908,In_385,In_997);
nand U909 (N_909,In_564,In_129);
nand U910 (N_910,In_753,In_631);
nand U911 (N_911,In_668,In_22);
nor U912 (N_912,In_660,In_333);
or U913 (N_913,In_310,In_186);
and U914 (N_914,In_482,In_12);
nand U915 (N_915,In_643,In_345);
or U916 (N_916,In_732,In_285);
xnor U917 (N_917,In_98,In_896);
nor U918 (N_918,In_260,In_502);
or U919 (N_919,In_388,In_166);
nand U920 (N_920,In_776,In_11);
or U921 (N_921,In_89,In_794);
nand U922 (N_922,In_925,In_219);
or U923 (N_923,In_849,In_154);
or U924 (N_924,In_509,In_666);
nand U925 (N_925,In_82,In_798);
and U926 (N_926,In_761,In_925);
and U927 (N_927,In_735,In_294);
xnor U928 (N_928,In_520,In_805);
and U929 (N_929,In_141,In_708);
xnor U930 (N_930,In_26,In_610);
xor U931 (N_931,In_741,In_798);
nor U932 (N_932,In_546,In_912);
or U933 (N_933,In_681,In_208);
and U934 (N_934,In_406,In_374);
nor U935 (N_935,In_466,In_362);
xnor U936 (N_936,In_611,In_858);
and U937 (N_937,In_840,In_344);
and U938 (N_938,In_620,In_284);
nor U939 (N_939,In_841,In_578);
xor U940 (N_940,In_631,In_840);
nand U941 (N_941,In_243,In_753);
nand U942 (N_942,In_590,In_2);
xnor U943 (N_943,In_579,In_279);
or U944 (N_944,In_322,In_427);
and U945 (N_945,In_48,In_348);
nand U946 (N_946,In_311,In_942);
and U947 (N_947,In_466,In_88);
and U948 (N_948,In_780,In_665);
xor U949 (N_949,In_64,In_515);
nor U950 (N_950,In_867,In_20);
and U951 (N_951,In_688,In_702);
and U952 (N_952,In_358,In_616);
nor U953 (N_953,In_9,In_427);
nor U954 (N_954,In_561,In_908);
or U955 (N_955,In_414,In_184);
nor U956 (N_956,In_309,In_898);
and U957 (N_957,In_649,In_22);
and U958 (N_958,In_715,In_586);
xnor U959 (N_959,In_715,In_15);
and U960 (N_960,In_330,In_285);
xnor U961 (N_961,In_657,In_734);
or U962 (N_962,In_425,In_565);
xor U963 (N_963,In_575,In_183);
nand U964 (N_964,In_742,In_458);
nor U965 (N_965,In_666,In_384);
nand U966 (N_966,In_432,In_797);
and U967 (N_967,In_235,In_29);
and U968 (N_968,In_274,In_715);
and U969 (N_969,In_881,In_125);
or U970 (N_970,In_381,In_907);
and U971 (N_971,In_110,In_903);
nor U972 (N_972,In_622,In_630);
and U973 (N_973,In_347,In_118);
or U974 (N_974,In_894,In_365);
nor U975 (N_975,In_26,In_452);
nor U976 (N_976,In_682,In_162);
nand U977 (N_977,In_418,In_723);
xnor U978 (N_978,In_403,In_959);
nand U979 (N_979,In_198,In_812);
or U980 (N_980,In_990,In_249);
nand U981 (N_981,In_775,In_419);
nand U982 (N_982,In_347,In_805);
xnor U983 (N_983,In_35,In_336);
and U984 (N_984,In_885,In_295);
or U985 (N_985,In_583,In_30);
nor U986 (N_986,In_102,In_894);
nor U987 (N_987,In_331,In_259);
or U988 (N_988,In_768,In_83);
nand U989 (N_989,In_790,In_468);
xnor U990 (N_990,In_652,In_233);
xnor U991 (N_991,In_276,In_582);
nor U992 (N_992,In_492,In_644);
nand U993 (N_993,In_835,In_363);
nand U994 (N_994,In_412,In_657);
nand U995 (N_995,In_198,In_59);
xnor U996 (N_996,In_360,In_310);
nand U997 (N_997,In_398,In_464);
or U998 (N_998,In_447,In_672);
or U999 (N_999,In_769,In_346);
nand U1000 (N_1000,In_189,In_526);
xnor U1001 (N_1001,In_255,In_504);
and U1002 (N_1002,In_376,In_246);
and U1003 (N_1003,In_989,In_539);
nor U1004 (N_1004,In_191,In_553);
and U1005 (N_1005,In_796,In_477);
nor U1006 (N_1006,In_919,In_911);
and U1007 (N_1007,In_890,In_152);
nand U1008 (N_1008,In_650,In_753);
or U1009 (N_1009,In_219,In_10);
or U1010 (N_1010,In_66,In_434);
xnor U1011 (N_1011,In_632,In_707);
and U1012 (N_1012,In_833,In_104);
nor U1013 (N_1013,In_880,In_97);
nor U1014 (N_1014,In_616,In_573);
nor U1015 (N_1015,In_623,In_350);
nor U1016 (N_1016,In_235,In_713);
and U1017 (N_1017,In_323,In_445);
xor U1018 (N_1018,In_804,In_74);
xnor U1019 (N_1019,In_840,In_190);
or U1020 (N_1020,In_843,In_480);
xnor U1021 (N_1021,In_488,In_270);
and U1022 (N_1022,In_284,In_306);
or U1023 (N_1023,In_42,In_253);
nand U1024 (N_1024,In_511,In_829);
nand U1025 (N_1025,In_317,In_156);
nor U1026 (N_1026,In_195,In_807);
nand U1027 (N_1027,In_999,In_977);
xnor U1028 (N_1028,In_800,In_903);
xnor U1029 (N_1029,In_605,In_722);
xnor U1030 (N_1030,In_664,In_595);
xnor U1031 (N_1031,In_424,In_324);
nand U1032 (N_1032,In_587,In_188);
nand U1033 (N_1033,In_777,In_605);
xor U1034 (N_1034,In_775,In_74);
xnor U1035 (N_1035,In_789,In_35);
xor U1036 (N_1036,In_677,In_183);
and U1037 (N_1037,In_946,In_552);
xor U1038 (N_1038,In_581,In_363);
nand U1039 (N_1039,In_569,In_991);
and U1040 (N_1040,In_574,In_886);
or U1041 (N_1041,In_384,In_810);
or U1042 (N_1042,In_584,In_138);
and U1043 (N_1043,In_5,In_915);
xnor U1044 (N_1044,In_445,In_603);
nand U1045 (N_1045,In_507,In_873);
and U1046 (N_1046,In_738,In_780);
nor U1047 (N_1047,In_422,In_248);
and U1048 (N_1048,In_61,In_229);
nand U1049 (N_1049,In_423,In_881);
nand U1050 (N_1050,In_498,In_913);
or U1051 (N_1051,In_221,In_266);
nand U1052 (N_1052,In_563,In_272);
xor U1053 (N_1053,In_353,In_29);
nor U1054 (N_1054,In_70,In_719);
nand U1055 (N_1055,In_596,In_957);
and U1056 (N_1056,In_110,In_121);
xor U1057 (N_1057,In_146,In_420);
nand U1058 (N_1058,In_527,In_981);
and U1059 (N_1059,In_981,In_597);
nand U1060 (N_1060,In_670,In_745);
nor U1061 (N_1061,In_822,In_970);
nand U1062 (N_1062,In_18,In_422);
nand U1063 (N_1063,In_986,In_917);
xnor U1064 (N_1064,In_881,In_945);
xor U1065 (N_1065,In_215,In_769);
xnor U1066 (N_1066,In_301,In_378);
or U1067 (N_1067,In_894,In_641);
xor U1068 (N_1068,In_456,In_147);
nand U1069 (N_1069,In_860,In_749);
xnor U1070 (N_1070,In_207,In_73);
xnor U1071 (N_1071,In_689,In_500);
or U1072 (N_1072,In_468,In_614);
xnor U1073 (N_1073,In_204,In_583);
xor U1074 (N_1074,In_657,In_116);
nand U1075 (N_1075,In_233,In_340);
or U1076 (N_1076,In_299,In_293);
nor U1077 (N_1077,In_411,In_427);
or U1078 (N_1078,In_510,In_576);
nor U1079 (N_1079,In_545,In_842);
nand U1080 (N_1080,In_846,In_583);
or U1081 (N_1081,In_592,In_584);
and U1082 (N_1082,In_182,In_291);
or U1083 (N_1083,In_725,In_623);
and U1084 (N_1084,In_380,In_874);
or U1085 (N_1085,In_872,In_946);
xnor U1086 (N_1086,In_342,In_726);
nor U1087 (N_1087,In_887,In_393);
xor U1088 (N_1088,In_11,In_424);
nand U1089 (N_1089,In_40,In_455);
or U1090 (N_1090,In_147,In_697);
and U1091 (N_1091,In_868,In_840);
xnor U1092 (N_1092,In_773,In_8);
or U1093 (N_1093,In_447,In_781);
nor U1094 (N_1094,In_753,In_652);
nand U1095 (N_1095,In_662,In_708);
and U1096 (N_1096,In_406,In_806);
and U1097 (N_1097,In_845,In_591);
xnor U1098 (N_1098,In_761,In_889);
or U1099 (N_1099,In_139,In_73);
or U1100 (N_1100,In_162,In_283);
xor U1101 (N_1101,In_728,In_872);
xnor U1102 (N_1102,In_139,In_58);
and U1103 (N_1103,In_246,In_22);
xnor U1104 (N_1104,In_53,In_407);
nand U1105 (N_1105,In_250,In_422);
xor U1106 (N_1106,In_273,In_607);
or U1107 (N_1107,In_312,In_876);
or U1108 (N_1108,In_318,In_145);
nor U1109 (N_1109,In_536,In_748);
nor U1110 (N_1110,In_448,In_461);
nor U1111 (N_1111,In_458,In_882);
nand U1112 (N_1112,In_617,In_963);
nand U1113 (N_1113,In_390,In_445);
nand U1114 (N_1114,In_268,In_22);
nor U1115 (N_1115,In_229,In_118);
nand U1116 (N_1116,In_6,In_43);
nand U1117 (N_1117,In_981,In_446);
and U1118 (N_1118,In_140,In_639);
xor U1119 (N_1119,In_947,In_510);
nor U1120 (N_1120,In_871,In_997);
nor U1121 (N_1121,In_434,In_747);
xnor U1122 (N_1122,In_923,In_834);
or U1123 (N_1123,In_859,In_783);
nor U1124 (N_1124,In_232,In_752);
or U1125 (N_1125,In_923,In_633);
xnor U1126 (N_1126,In_727,In_784);
or U1127 (N_1127,In_235,In_975);
or U1128 (N_1128,In_872,In_285);
or U1129 (N_1129,In_60,In_763);
nor U1130 (N_1130,In_523,In_570);
nor U1131 (N_1131,In_892,In_806);
nor U1132 (N_1132,In_845,In_85);
nand U1133 (N_1133,In_665,In_388);
xor U1134 (N_1134,In_15,In_755);
xnor U1135 (N_1135,In_523,In_111);
and U1136 (N_1136,In_922,In_360);
nor U1137 (N_1137,In_901,In_260);
nor U1138 (N_1138,In_659,In_482);
or U1139 (N_1139,In_604,In_775);
or U1140 (N_1140,In_565,In_694);
or U1141 (N_1141,In_894,In_119);
and U1142 (N_1142,In_536,In_53);
nand U1143 (N_1143,In_185,In_758);
nand U1144 (N_1144,In_943,In_810);
xnor U1145 (N_1145,In_573,In_292);
nand U1146 (N_1146,In_96,In_834);
xnor U1147 (N_1147,In_96,In_513);
nor U1148 (N_1148,In_345,In_958);
or U1149 (N_1149,In_958,In_63);
or U1150 (N_1150,In_573,In_160);
nor U1151 (N_1151,In_295,In_889);
nor U1152 (N_1152,In_895,In_403);
and U1153 (N_1153,In_632,In_476);
or U1154 (N_1154,In_473,In_1);
or U1155 (N_1155,In_414,In_715);
or U1156 (N_1156,In_123,In_581);
nand U1157 (N_1157,In_255,In_361);
and U1158 (N_1158,In_782,In_262);
xor U1159 (N_1159,In_128,In_485);
and U1160 (N_1160,In_195,In_262);
nand U1161 (N_1161,In_433,In_768);
and U1162 (N_1162,In_728,In_145);
nor U1163 (N_1163,In_37,In_609);
xor U1164 (N_1164,In_904,In_552);
nand U1165 (N_1165,In_673,In_134);
xnor U1166 (N_1166,In_7,In_986);
or U1167 (N_1167,In_513,In_395);
nor U1168 (N_1168,In_103,In_86);
xnor U1169 (N_1169,In_211,In_627);
xor U1170 (N_1170,In_29,In_7);
or U1171 (N_1171,In_706,In_650);
and U1172 (N_1172,In_424,In_292);
nand U1173 (N_1173,In_407,In_900);
nor U1174 (N_1174,In_925,In_855);
nand U1175 (N_1175,In_365,In_542);
and U1176 (N_1176,In_988,In_146);
or U1177 (N_1177,In_884,In_862);
or U1178 (N_1178,In_196,In_744);
nand U1179 (N_1179,In_26,In_303);
or U1180 (N_1180,In_209,In_300);
or U1181 (N_1181,In_425,In_4);
nor U1182 (N_1182,In_709,In_122);
or U1183 (N_1183,In_169,In_487);
or U1184 (N_1184,In_464,In_427);
xor U1185 (N_1185,In_543,In_41);
xor U1186 (N_1186,In_192,In_958);
and U1187 (N_1187,In_687,In_270);
nor U1188 (N_1188,In_4,In_1);
nor U1189 (N_1189,In_917,In_584);
and U1190 (N_1190,In_267,In_447);
and U1191 (N_1191,In_635,In_606);
xnor U1192 (N_1192,In_452,In_190);
and U1193 (N_1193,In_659,In_206);
xor U1194 (N_1194,In_415,In_144);
xor U1195 (N_1195,In_242,In_956);
or U1196 (N_1196,In_934,In_275);
nor U1197 (N_1197,In_572,In_38);
nor U1198 (N_1198,In_216,In_573);
xnor U1199 (N_1199,In_146,In_409);
or U1200 (N_1200,In_518,In_753);
nor U1201 (N_1201,In_432,In_623);
nor U1202 (N_1202,In_990,In_540);
xor U1203 (N_1203,In_716,In_303);
and U1204 (N_1204,In_711,In_731);
or U1205 (N_1205,In_391,In_186);
nand U1206 (N_1206,In_227,In_134);
xor U1207 (N_1207,In_954,In_980);
nand U1208 (N_1208,In_201,In_668);
or U1209 (N_1209,In_641,In_317);
xor U1210 (N_1210,In_416,In_248);
nor U1211 (N_1211,In_176,In_980);
and U1212 (N_1212,In_135,In_645);
and U1213 (N_1213,In_740,In_870);
xnor U1214 (N_1214,In_460,In_652);
xor U1215 (N_1215,In_16,In_287);
or U1216 (N_1216,In_7,In_972);
nand U1217 (N_1217,In_631,In_88);
or U1218 (N_1218,In_398,In_684);
or U1219 (N_1219,In_432,In_687);
or U1220 (N_1220,In_137,In_104);
and U1221 (N_1221,In_316,In_545);
nand U1222 (N_1222,In_334,In_772);
nand U1223 (N_1223,In_25,In_645);
xor U1224 (N_1224,In_916,In_999);
and U1225 (N_1225,In_209,In_47);
xnor U1226 (N_1226,In_291,In_707);
nor U1227 (N_1227,In_581,In_867);
nand U1228 (N_1228,In_470,In_13);
or U1229 (N_1229,In_665,In_484);
nand U1230 (N_1230,In_673,In_945);
and U1231 (N_1231,In_521,In_750);
nor U1232 (N_1232,In_788,In_360);
and U1233 (N_1233,In_148,In_850);
and U1234 (N_1234,In_715,In_819);
nand U1235 (N_1235,In_45,In_541);
xor U1236 (N_1236,In_521,In_870);
nor U1237 (N_1237,In_968,In_648);
nor U1238 (N_1238,In_989,In_733);
or U1239 (N_1239,In_441,In_828);
and U1240 (N_1240,In_535,In_623);
nand U1241 (N_1241,In_957,In_90);
xor U1242 (N_1242,In_678,In_187);
and U1243 (N_1243,In_813,In_709);
or U1244 (N_1244,In_243,In_294);
and U1245 (N_1245,In_849,In_884);
nand U1246 (N_1246,In_621,In_990);
xnor U1247 (N_1247,In_980,In_987);
xnor U1248 (N_1248,In_494,In_253);
and U1249 (N_1249,In_874,In_106);
xor U1250 (N_1250,In_736,In_528);
nor U1251 (N_1251,In_679,In_414);
or U1252 (N_1252,In_194,In_260);
nand U1253 (N_1253,In_698,In_899);
nor U1254 (N_1254,In_346,In_581);
nor U1255 (N_1255,In_220,In_815);
xor U1256 (N_1256,In_457,In_282);
nor U1257 (N_1257,In_518,In_375);
or U1258 (N_1258,In_615,In_544);
or U1259 (N_1259,In_624,In_583);
xor U1260 (N_1260,In_474,In_528);
or U1261 (N_1261,In_274,In_200);
and U1262 (N_1262,In_981,In_721);
or U1263 (N_1263,In_66,In_193);
or U1264 (N_1264,In_888,In_994);
or U1265 (N_1265,In_142,In_389);
nor U1266 (N_1266,In_410,In_464);
nand U1267 (N_1267,In_858,In_13);
nand U1268 (N_1268,In_647,In_93);
nand U1269 (N_1269,In_872,In_356);
and U1270 (N_1270,In_470,In_648);
and U1271 (N_1271,In_623,In_220);
xnor U1272 (N_1272,In_357,In_459);
nor U1273 (N_1273,In_542,In_196);
or U1274 (N_1274,In_642,In_560);
or U1275 (N_1275,In_425,In_759);
nor U1276 (N_1276,In_288,In_615);
and U1277 (N_1277,In_370,In_177);
nor U1278 (N_1278,In_723,In_619);
xor U1279 (N_1279,In_456,In_530);
or U1280 (N_1280,In_123,In_766);
xnor U1281 (N_1281,In_602,In_87);
and U1282 (N_1282,In_279,In_373);
or U1283 (N_1283,In_30,In_916);
and U1284 (N_1284,In_154,In_49);
or U1285 (N_1285,In_486,In_429);
nand U1286 (N_1286,In_308,In_531);
or U1287 (N_1287,In_870,In_435);
nor U1288 (N_1288,In_547,In_272);
nor U1289 (N_1289,In_936,In_989);
and U1290 (N_1290,In_591,In_261);
and U1291 (N_1291,In_524,In_35);
nor U1292 (N_1292,In_301,In_144);
nor U1293 (N_1293,In_591,In_765);
nand U1294 (N_1294,In_840,In_805);
xnor U1295 (N_1295,In_490,In_13);
or U1296 (N_1296,In_24,In_426);
or U1297 (N_1297,In_815,In_439);
and U1298 (N_1298,In_329,In_70);
nand U1299 (N_1299,In_509,In_388);
nand U1300 (N_1300,In_203,In_944);
nor U1301 (N_1301,In_550,In_35);
or U1302 (N_1302,In_323,In_529);
and U1303 (N_1303,In_786,In_365);
nand U1304 (N_1304,In_392,In_699);
or U1305 (N_1305,In_728,In_265);
and U1306 (N_1306,In_901,In_184);
nand U1307 (N_1307,In_211,In_839);
or U1308 (N_1308,In_338,In_312);
and U1309 (N_1309,In_975,In_386);
nand U1310 (N_1310,In_763,In_945);
or U1311 (N_1311,In_736,In_32);
xnor U1312 (N_1312,In_166,In_773);
nor U1313 (N_1313,In_266,In_137);
nor U1314 (N_1314,In_856,In_343);
xor U1315 (N_1315,In_564,In_928);
nand U1316 (N_1316,In_572,In_823);
and U1317 (N_1317,In_966,In_397);
or U1318 (N_1318,In_452,In_807);
nor U1319 (N_1319,In_632,In_846);
and U1320 (N_1320,In_16,In_989);
and U1321 (N_1321,In_188,In_318);
nor U1322 (N_1322,In_553,In_739);
xor U1323 (N_1323,In_729,In_17);
and U1324 (N_1324,In_693,In_766);
or U1325 (N_1325,In_543,In_507);
and U1326 (N_1326,In_143,In_298);
or U1327 (N_1327,In_727,In_603);
nor U1328 (N_1328,In_499,In_739);
xnor U1329 (N_1329,In_772,In_930);
xnor U1330 (N_1330,In_69,In_910);
or U1331 (N_1331,In_162,In_845);
nor U1332 (N_1332,In_231,In_32);
xnor U1333 (N_1333,In_303,In_840);
xor U1334 (N_1334,In_921,In_134);
or U1335 (N_1335,In_458,In_164);
or U1336 (N_1336,In_182,In_616);
nor U1337 (N_1337,In_269,In_133);
xor U1338 (N_1338,In_190,In_745);
and U1339 (N_1339,In_523,In_600);
nor U1340 (N_1340,In_256,In_562);
or U1341 (N_1341,In_80,In_821);
and U1342 (N_1342,In_736,In_702);
xnor U1343 (N_1343,In_752,In_445);
or U1344 (N_1344,In_518,In_202);
xnor U1345 (N_1345,In_422,In_227);
nor U1346 (N_1346,In_264,In_0);
nor U1347 (N_1347,In_936,In_455);
nor U1348 (N_1348,In_764,In_191);
nand U1349 (N_1349,In_394,In_229);
xor U1350 (N_1350,In_977,In_397);
or U1351 (N_1351,In_130,In_333);
nand U1352 (N_1352,In_70,In_770);
xnor U1353 (N_1353,In_499,In_227);
nor U1354 (N_1354,In_674,In_93);
xnor U1355 (N_1355,In_7,In_645);
and U1356 (N_1356,In_390,In_320);
or U1357 (N_1357,In_799,In_747);
nand U1358 (N_1358,In_415,In_101);
or U1359 (N_1359,In_813,In_889);
xor U1360 (N_1360,In_646,In_599);
nor U1361 (N_1361,In_114,In_111);
or U1362 (N_1362,In_752,In_527);
xnor U1363 (N_1363,In_195,In_394);
and U1364 (N_1364,In_237,In_715);
and U1365 (N_1365,In_202,In_980);
or U1366 (N_1366,In_984,In_265);
or U1367 (N_1367,In_116,In_157);
and U1368 (N_1368,In_664,In_967);
xor U1369 (N_1369,In_119,In_425);
or U1370 (N_1370,In_400,In_366);
and U1371 (N_1371,In_769,In_368);
xor U1372 (N_1372,In_207,In_46);
nand U1373 (N_1373,In_260,In_763);
xor U1374 (N_1374,In_51,In_191);
nand U1375 (N_1375,In_887,In_620);
or U1376 (N_1376,In_661,In_222);
or U1377 (N_1377,In_653,In_85);
nor U1378 (N_1378,In_139,In_696);
or U1379 (N_1379,In_804,In_238);
or U1380 (N_1380,In_277,In_532);
xor U1381 (N_1381,In_486,In_958);
nand U1382 (N_1382,In_737,In_748);
nor U1383 (N_1383,In_276,In_139);
nor U1384 (N_1384,In_156,In_540);
nor U1385 (N_1385,In_731,In_724);
nand U1386 (N_1386,In_698,In_292);
xnor U1387 (N_1387,In_504,In_402);
nand U1388 (N_1388,In_284,In_631);
or U1389 (N_1389,In_833,In_115);
nand U1390 (N_1390,In_944,In_176);
or U1391 (N_1391,In_861,In_24);
and U1392 (N_1392,In_134,In_626);
nor U1393 (N_1393,In_171,In_167);
xor U1394 (N_1394,In_558,In_257);
and U1395 (N_1395,In_874,In_741);
nand U1396 (N_1396,In_45,In_898);
nor U1397 (N_1397,In_573,In_605);
xor U1398 (N_1398,In_484,In_501);
nor U1399 (N_1399,In_591,In_194);
nor U1400 (N_1400,In_463,In_730);
xor U1401 (N_1401,In_210,In_386);
or U1402 (N_1402,In_571,In_848);
and U1403 (N_1403,In_698,In_773);
and U1404 (N_1404,In_471,In_373);
or U1405 (N_1405,In_572,In_279);
xor U1406 (N_1406,In_400,In_573);
nand U1407 (N_1407,In_498,In_806);
nor U1408 (N_1408,In_992,In_634);
and U1409 (N_1409,In_782,In_774);
or U1410 (N_1410,In_107,In_50);
nor U1411 (N_1411,In_613,In_961);
xnor U1412 (N_1412,In_253,In_116);
nor U1413 (N_1413,In_465,In_824);
nand U1414 (N_1414,In_114,In_539);
and U1415 (N_1415,In_114,In_778);
nand U1416 (N_1416,In_348,In_606);
or U1417 (N_1417,In_384,In_536);
and U1418 (N_1418,In_108,In_934);
nor U1419 (N_1419,In_306,In_532);
nor U1420 (N_1420,In_851,In_134);
nand U1421 (N_1421,In_675,In_135);
or U1422 (N_1422,In_305,In_990);
and U1423 (N_1423,In_332,In_808);
nor U1424 (N_1424,In_345,In_375);
xor U1425 (N_1425,In_703,In_864);
and U1426 (N_1426,In_84,In_575);
nor U1427 (N_1427,In_831,In_376);
and U1428 (N_1428,In_959,In_615);
and U1429 (N_1429,In_278,In_14);
nand U1430 (N_1430,In_713,In_138);
and U1431 (N_1431,In_772,In_688);
nand U1432 (N_1432,In_866,In_327);
or U1433 (N_1433,In_281,In_803);
and U1434 (N_1434,In_402,In_257);
nor U1435 (N_1435,In_675,In_849);
nand U1436 (N_1436,In_671,In_756);
xnor U1437 (N_1437,In_756,In_827);
and U1438 (N_1438,In_716,In_261);
xnor U1439 (N_1439,In_17,In_553);
xor U1440 (N_1440,In_447,In_527);
or U1441 (N_1441,In_139,In_902);
xnor U1442 (N_1442,In_446,In_612);
or U1443 (N_1443,In_502,In_392);
nor U1444 (N_1444,In_982,In_553);
xor U1445 (N_1445,In_914,In_508);
xor U1446 (N_1446,In_681,In_534);
and U1447 (N_1447,In_374,In_146);
xor U1448 (N_1448,In_430,In_368);
nand U1449 (N_1449,In_160,In_155);
and U1450 (N_1450,In_831,In_654);
and U1451 (N_1451,In_763,In_163);
xnor U1452 (N_1452,In_744,In_965);
xnor U1453 (N_1453,In_916,In_218);
and U1454 (N_1454,In_635,In_424);
and U1455 (N_1455,In_634,In_377);
xnor U1456 (N_1456,In_23,In_166);
xnor U1457 (N_1457,In_910,In_668);
nand U1458 (N_1458,In_515,In_178);
xor U1459 (N_1459,In_354,In_434);
xor U1460 (N_1460,In_804,In_98);
xnor U1461 (N_1461,In_984,In_76);
xor U1462 (N_1462,In_745,In_826);
or U1463 (N_1463,In_679,In_75);
or U1464 (N_1464,In_229,In_28);
nand U1465 (N_1465,In_746,In_959);
xor U1466 (N_1466,In_457,In_360);
or U1467 (N_1467,In_852,In_846);
or U1468 (N_1468,In_653,In_422);
and U1469 (N_1469,In_235,In_256);
xor U1470 (N_1470,In_297,In_124);
or U1471 (N_1471,In_161,In_175);
xor U1472 (N_1472,In_944,In_839);
xnor U1473 (N_1473,In_463,In_965);
nand U1474 (N_1474,In_837,In_574);
and U1475 (N_1475,In_39,In_920);
xor U1476 (N_1476,In_196,In_600);
and U1477 (N_1477,In_653,In_197);
nand U1478 (N_1478,In_238,In_177);
nand U1479 (N_1479,In_100,In_858);
nand U1480 (N_1480,In_728,In_688);
or U1481 (N_1481,In_173,In_263);
xnor U1482 (N_1482,In_782,In_969);
and U1483 (N_1483,In_63,In_753);
nand U1484 (N_1484,In_81,In_500);
nand U1485 (N_1485,In_270,In_328);
nand U1486 (N_1486,In_168,In_398);
and U1487 (N_1487,In_166,In_5);
xor U1488 (N_1488,In_356,In_143);
nor U1489 (N_1489,In_286,In_96);
or U1490 (N_1490,In_402,In_564);
or U1491 (N_1491,In_668,In_511);
nor U1492 (N_1492,In_365,In_249);
nand U1493 (N_1493,In_771,In_730);
nand U1494 (N_1494,In_357,In_785);
nand U1495 (N_1495,In_162,In_918);
nor U1496 (N_1496,In_471,In_372);
xor U1497 (N_1497,In_9,In_6);
nor U1498 (N_1498,In_912,In_329);
xnor U1499 (N_1499,In_177,In_31);
xnor U1500 (N_1500,In_119,In_411);
xnor U1501 (N_1501,In_433,In_38);
xor U1502 (N_1502,In_19,In_201);
or U1503 (N_1503,In_432,In_988);
xor U1504 (N_1504,In_688,In_653);
nand U1505 (N_1505,In_258,In_904);
nand U1506 (N_1506,In_293,In_147);
nor U1507 (N_1507,In_901,In_464);
nor U1508 (N_1508,In_45,In_23);
xor U1509 (N_1509,In_742,In_292);
nor U1510 (N_1510,In_241,In_749);
or U1511 (N_1511,In_859,In_501);
xor U1512 (N_1512,In_442,In_788);
xor U1513 (N_1513,In_170,In_879);
nand U1514 (N_1514,In_515,In_965);
or U1515 (N_1515,In_220,In_189);
and U1516 (N_1516,In_215,In_994);
nor U1517 (N_1517,In_542,In_228);
xnor U1518 (N_1518,In_364,In_939);
or U1519 (N_1519,In_589,In_461);
and U1520 (N_1520,In_251,In_108);
xor U1521 (N_1521,In_317,In_708);
nand U1522 (N_1522,In_923,In_775);
and U1523 (N_1523,In_5,In_561);
nor U1524 (N_1524,In_492,In_454);
or U1525 (N_1525,In_564,In_271);
nand U1526 (N_1526,In_79,In_705);
nor U1527 (N_1527,In_208,In_83);
xor U1528 (N_1528,In_472,In_468);
or U1529 (N_1529,In_337,In_926);
nor U1530 (N_1530,In_946,In_87);
nor U1531 (N_1531,In_18,In_483);
xnor U1532 (N_1532,In_291,In_574);
nor U1533 (N_1533,In_934,In_639);
and U1534 (N_1534,In_533,In_419);
xor U1535 (N_1535,In_919,In_230);
or U1536 (N_1536,In_99,In_985);
xor U1537 (N_1537,In_377,In_810);
and U1538 (N_1538,In_936,In_94);
nor U1539 (N_1539,In_649,In_910);
xor U1540 (N_1540,In_552,In_128);
and U1541 (N_1541,In_402,In_333);
nor U1542 (N_1542,In_36,In_162);
and U1543 (N_1543,In_459,In_819);
nor U1544 (N_1544,In_712,In_121);
and U1545 (N_1545,In_668,In_380);
nor U1546 (N_1546,In_459,In_515);
nor U1547 (N_1547,In_488,In_796);
and U1548 (N_1548,In_908,In_755);
nand U1549 (N_1549,In_832,In_568);
and U1550 (N_1550,In_845,In_787);
nand U1551 (N_1551,In_890,In_676);
or U1552 (N_1552,In_682,In_815);
nor U1553 (N_1553,In_346,In_444);
and U1554 (N_1554,In_767,In_5);
nor U1555 (N_1555,In_909,In_925);
xnor U1556 (N_1556,In_553,In_72);
or U1557 (N_1557,In_474,In_655);
nor U1558 (N_1558,In_410,In_930);
or U1559 (N_1559,In_388,In_347);
and U1560 (N_1560,In_747,In_256);
or U1561 (N_1561,In_26,In_601);
and U1562 (N_1562,In_301,In_563);
nor U1563 (N_1563,In_106,In_695);
nand U1564 (N_1564,In_758,In_623);
nand U1565 (N_1565,In_753,In_164);
nand U1566 (N_1566,In_932,In_270);
or U1567 (N_1567,In_104,In_471);
nor U1568 (N_1568,In_873,In_899);
nor U1569 (N_1569,In_862,In_914);
xor U1570 (N_1570,In_668,In_971);
and U1571 (N_1571,In_659,In_745);
nand U1572 (N_1572,In_329,In_203);
or U1573 (N_1573,In_438,In_214);
nor U1574 (N_1574,In_518,In_676);
nor U1575 (N_1575,In_601,In_331);
nor U1576 (N_1576,In_154,In_645);
nand U1577 (N_1577,In_429,In_493);
and U1578 (N_1578,In_190,In_732);
nand U1579 (N_1579,In_42,In_784);
or U1580 (N_1580,In_807,In_675);
and U1581 (N_1581,In_609,In_264);
and U1582 (N_1582,In_196,In_194);
nor U1583 (N_1583,In_646,In_818);
xnor U1584 (N_1584,In_626,In_766);
xnor U1585 (N_1585,In_307,In_904);
nand U1586 (N_1586,In_227,In_363);
nand U1587 (N_1587,In_528,In_5);
nor U1588 (N_1588,In_393,In_12);
or U1589 (N_1589,In_370,In_775);
xor U1590 (N_1590,In_866,In_924);
xnor U1591 (N_1591,In_777,In_39);
and U1592 (N_1592,In_72,In_101);
or U1593 (N_1593,In_77,In_857);
and U1594 (N_1594,In_258,In_149);
xnor U1595 (N_1595,In_906,In_17);
xnor U1596 (N_1596,In_697,In_998);
xor U1597 (N_1597,In_428,In_34);
xor U1598 (N_1598,In_815,In_174);
and U1599 (N_1599,In_729,In_712);
xor U1600 (N_1600,In_94,In_893);
and U1601 (N_1601,In_430,In_302);
nand U1602 (N_1602,In_347,In_121);
and U1603 (N_1603,In_316,In_288);
nor U1604 (N_1604,In_835,In_890);
nor U1605 (N_1605,In_846,In_178);
nand U1606 (N_1606,In_580,In_589);
xor U1607 (N_1607,In_21,In_511);
and U1608 (N_1608,In_898,In_596);
or U1609 (N_1609,In_803,In_599);
xnor U1610 (N_1610,In_335,In_412);
nor U1611 (N_1611,In_913,In_859);
nor U1612 (N_1612,In_426,In_63);
nor U1613 (N_1613,In_921,In_350);
xor U1614 (N_1614,In_381,In_174);
xnor U1615 (N_1615,In_876,In_951);
nand U1616 (N_1616,In_462,In_912);
or U1617 (N_1617,In_462,In_332);
xor U1618 (N_1618,In_650,In_948);
xor U1619 (N_1619,In_974,In_23);
nor U1620 (N_1620,In_643,In_314);
xnor U1621 (N_1621,In_490,In_863);
nor U1622 (N_1622,In_84,In_700);
xnor U1623 (N_1623,In_411,In_580);
and U1624 (N_1624,In_336,In_896);
xnor U1625 (N_1625,In_571,In_970);
nand U1626 (N_1626,In_512,In_146);
nand U1627 (N_1627,In_508,In_623);
xnor U1628 (N_1628,In_152,In_767);
xnor U1629 (N_1629,In_24,In_52);
nor U1630 (N_1630,In_407,In_225);
nand U1631 (N_1631,In_291,In_184);
xor U1632 (N_1632,In_496,In_843);
nor U1633 (N_1633,In_666,In_457);
nand U1634 (N_1634,In_253,In_223);
and U1635 (N_1635,In_808,In_575);
or U1636 (N_1636,In_822,In_9);
nor U1637 (N_1637,In_70,In_586);
and U1638 (N_1638,In_282,In_640);
nor U1639 (N_1639,In_356,In_845);
xor U1640 (N_1640,In_259,In_662);
xnor U1641 (N_1641,In_395,In_318);
nand U1642 (N_1642,In_310,In_125);
nand U1643 (N_1643,In_236,In_896);
xor U1644 (N_1644,In_330,In_406);
xnor U1645 (N_1645,In_400,In_603);
nand U1646 (N_1646,In_694,In_381);
xnor U1647 (N_1647,In_229,In_181);
nor U1648 (N_1648,In_615,In_31);
or U1649 (N_1649,In_470,In_835);
and U1650 (N_1650,In_980,In_94);
nor U1651 (N_1651,In_828,In_978);
nand U1652 (N_1652,In_624,In_369);
and U1653 (N_1653,In_47,In_256);
and U1654 (N_1654,In_472,In_32);
or U1655 (N_1655,In_833,In_693);
and U1656 (N_1656,In_138,In_819);
nor U1657 (N_1657,In_121,In_307);
nand U1658 (N_1658,In_386,In_559);
xor U1659 (N_1659,In_15,In_806);
xor U1660 (N_1660,In_354,In_126);
and U1661 (N_1661,In_332,In_385);
or U1662 (N_1662,In_715,In_920);
and U1663 (N_1663,In_536,In_206);
nor U1664 (N_1664,In_372,In_666);
nor U1665 (N_1665,In_27,In_19);
and U1666 (N_1666,In_398,In_795);
or U1667 (N_1667,In_549,In_515);
or U1668 (N_1668,In_74,In_678);
or U1669 (N_1669,In_653,In_903);
and U1670 (N_1670,In_478,In_860);
nor U1671 (N_1671,In_503,In_185);
nor U1672 (N_1672,In_359,In_540);
and U1673 (N_1673,In_626,In_152);
nand U1674 (N_1674,In_998,In_658);
nand U1675 (N_1675,In_473,In_111);
xnor U1676 (N_1676,In_763,In_529);
or U1677 (N_1677,In_772,In_875);
and U1678 (N_1678,In_827,In_144);
nand U1679 (N_1679,In_393,In_666);
nand U1680 (N_1680,In_791,In_318);
and U1681 (N_1681,In_136,In_394);
nand U1682 (N_1682,In_149,In_529);
xnor U1683 (N_1683,In_565,In_753);
and U1684 (N_1684,In_495,In_341);
xor U1685 (N_1685,In_268,In_866);
nand U1686 (N_1686,In_442,In_962);
and U1687 (N_1687,In_970,In_265);
nand U1688 (N_1688,In_510,In_462);
or U1689 (N_1689,In_333,In_767);
or U1690 (N_1690,In_811,In_955);
or U1691 (N_1691,In_858,In_827);
nand U1692 (N_1692,In_823,In_552);
nor U1693 (N_1693,In_952,In_296);
or U1694 (N_1694,In_312,In_274);
and U1695 (N_1695,In_312,In_432);
and U1696 (N_1696,In_669,In_294);
nand U1697 (N_1697,In_233,In_308);
nand U1698 (N_1698,In_973,In_464);
or U1699 (N_1699,In_62,In_220);
and U1700 (N_1700,In_475,In_187);
nor U1701 (N_1701,In_327,In_972);
nor U1702 (N_1702,In_400,In_805);
and U1703 (N_1703,In_975,In_296);
nand U1704 (N_1704,In_519,In_307);
nor U1705 (N_1705,In_285,In_736);
nand U1706 (N_1706,In_960,In_774);
or U1707 (N_1707,In_291,In_616);
xnor U1708 (N_1708,In_962,In_165);
and U1709 (N_1709,In_262,In_939);
and U1710 (N_1710,In_341,In_551);
nand U1711 (N_1711,In_598,In_259);
nor U1712 (N_1712,In_599,In_199);
nand U1713 (N_1713,In_880,In_395);
nand U1714 (N_1714,In_449,In_303);
and U1715 (N_1715,In_334,In_798);
xnor U1716 (N_1716,In_451,In_846);
or U1717 (N_1717,In_199,In_108);
nand U1718 (N_1718,In_430,In_919);
nand U1719 (N_1719,In_865,In_867);
or U1720 (N_1720,In_6,In_69);
or U1721 (N_1721,In_912,In_358);
or U1722 (N_1722,In_513,In_329);
xnor U1723 (N_1723,In_449,In_919);
or U1724 (N_1724,In_215,In_958);
nor U1725 (N_1725,In_155,In_479);
xor U1726 (N_1726,In_19,In_429);
xor U1727 (N_1727,In_636,In_838);
nand U1728 (N_1728,In_775,In_544);
nand U1729 (N_1729,In_486,In_225);
nand U1730 (N_1730,In_662,In_266);
and U1731 (N_1731,In_833,In_197);
and U1732 (N_1732,In_334,In_767);
nand U1733 (N_1733,In_308,In_707);
and U1734 (N_1734,In_246,In_658);
xnor U1735 (N_1735,In_810,In_706);
nor U1736 (N_1736,In_65,In_394);
and U1737 (N_1737,In_259,In_553);
xor U1738 (N_1738,In_787,In_342);
nand U1739 (N_1739,In_288,In_934);
or U1740 (N_1740,In_856,In_631);
nor U1741 (N_1741,In_550,In_720);
and U1742 (N_1742,In_5,In_48);
and U1743 (N_1743,In_924,In_18);
and U1744 (N_1744,In_627,In_501);
xor U1745 (N_1745,In_803,In_846);
xor U1746 (N_1746,In_344,In_322);
nand U1747 (N_1747,In_635,In_983);
or U1748 (N_1748,In_953,In_191);
xnor U1749 (N_1749,In_182,In_236);
nand U1750 (N_1750,In_944,In_464);
or U1751 (N_1751,In_172,In_574);
nor U1752 (N_1752,In_330,In_633);
nand U1753 (N_1753,In_124,In_685);
or U1754 (N_1754,In_279,In_679);
nand U1755 (N_1755,In_263,In_812);
and U1756 (N_1756,In_394,In_446);
nor U1757 (N_1757,In_194,In_17);
nand U1758 (N_1758,In_64,In_545);
xor U1759 (N_1759,In_441,In_481);
or U1760 (N_1760,In_829,In_762);
and U1761 (N_1761,In_534,In_332);
xnor U1762 (N_1762,In_947,In_227);
xor U1763 (N_1763,In_427,In_294);
or U1764 (N_1764,In_154,In_250);
nand U1765 (N_1765,In_511,In_915);
and U1766 (N_1766,In_94,In_677);
and U1767 (N_1767,In_302,In_215);
nor U1768 (N_1768,In_685,In_58);
nor U1769 (N_1769,In_695,In_956);
nor U1770 (N_1770,In_742,In_352);
nand U1771 (N_1771,In_878,In_136);
nor U1772 (N_1772,In_447,In_190);
and U1773 (N_1773,In_737,In_372);
nand U1774 (N_1774,In_715,In_566);
nand U1775 (N_1775,In_403,In_105);
xnor U1776 (N_1776,In_271,In_979);
xor U1777 (N_1777,In_19,In_698);
xnor U1778 (N_1778,In_913,In_806);
and U1779 (N_1779,In_90,In_171);
nand U1780 (N_1780,In_59,In_690);
or U1781 (N_1781,In_233,In_526);
xnor U1782 (N_1782,In_981,In_248);
or U1783 (N_1783,In_552,In_851);
xor U1784 (N_1784,In_961,In_845);
nand U1785 (N_1785,In_401,In_94);
and U1786 (N_1786,In_655,In_880);
and U1787 (N_1787,In_102,In_436);
nor U1788 (N_1788,In_246,In_728);
or U1789 (N_1789,In_789,In_637);
nor U1790 (N_1790,In_715,In_791);
nand U1791 (N_1791,In_393,In_711);
nor U1792 (N_1792,In_194,In_408);
nand U1793 (N_1793,In_833,In_866);
and U1794 (N_1794,In_857,In_20);
nand U1795 (N_1795,In_575,In_788);
xor U1796 (N_1796,In_180,In_437);
xor U1797 (N_1797,In_57,In_939);
xor U1798 (N_1798,In_781,In_945);
nor U1799 (N_1799,In_103,In_780);
and U1800 (N_1800,In_287,In_364);
nand U1801 (N_1801,In_78,In_445);
and U1802 (N_1802,In_684,In_473);
or U1803 (N_1803,In_630,In_472);
nor U1804 (N_1804,In_195,In_671);
and U1805 (N_1805,In_321,In_699);
and U1806 (N_1806,In_836,In_165);
nor U1807 (N_1807,In_559,In_321);
nor U1808 (N_1808,In_940,In_165);
or U1809 (N_1809,In_776,In_408);
xor U1810 (N_1810,In_379,In_571);
xnor U1811 (N_1811,In_579,In_359);
nor U1812 (N_1812,In_442,In_677);
and U1813 (N_1813,In_801,In_375);
nor U1814 (N_1814,In_950,In_405);
nand U1815 (N_1815,In_734,In_912);
and U1816 (N_1816,In_852,In_226);
xor U1817 (N_1817,In_858,In_468);
and U1818 (N_1818,In_157,In_292);
nor U1819 (N_1819,In_553,In_593);
or U1820 (N_1820,In_347,In_1);
or U1821 (N_1821,In_445,In_493);
and U1822 (N_1822,In_426,In_635);
nor U1823 (N_1823,In_500,In_79);
or U1824 (N_1824,In_127,In_582);
xor U1825 (N_1825,In_540,In_822);
and U1826 (N_1826,In_379,In_349);
nor U1827 (N_1827,In_920,In_533);
and U1828 (N_1828,In_65,In_276);
and U1829 (N_1829,In_644,In_754);
or U1830 (N_1830,In_659,In_17);
and U1831 (N_1831,In_131,In_653);
xor U1832 (N_1832,In_506,In_762);
and U1833 (N_1833,In_359,In_239);
xor U1834 (N_1834,In_593,In_789);
nand U1835 (N_1835,In_825,In_994);
nand U1836 (N_1836,In_769,In_712);
and U1837 (N_1837,In_484,In_716);
nor U1838 (N_1838,In_634,In_704);
or U1839 (N_1839,In_642,In_335);
xor U1840 (N_1840,In_593,In_458);
nand U1841 (N_1841,In_599,In_763);
nand U1842 (N_1842,In_402,In_53);
nand U1843 (N_1843,In_2,In_337);
xor U1844 (N_1844,In_251,In_902);
xor U1845 (N_1845,In_664,In_916);
or U1846 (N_1846,In_805,In_633);
nand U1847 (N_1847,In_510,In_606);
nand U1848 (N_1848,In_744,In_653);
or U1849 (N_1849,In_945,In_733);
and U1850 (N_1850,In_512,In_258);
xor U1851 (N_1851,In_939,In_846);
nand U1852 (N_1852,In_635,In_849);
nand U1853 (N_1853,In_100,In_149);
nand U1854 (N_1854,In_989,In_104);
nor U1855 (N_1855,In_127,In_477);
nand U1856 (N_1856,In_36,In_402);
nor U1857 (N_1857,In_40,In_936);
xnor U1858 (N_1858,In_407,In_167);
and U1859 (N_1859,In_191,In_125);
nor U1860 (N_1860,In_976,In_815);
xnor U1861 (N_1861,In_232,In_632);
or U1862 (N_1862,In_536,In_397);
nand U1863 (N_1863,In_849,In_614);
nand U1864 (N_1864,In_887,In_247);
nand U1865 (N_1865,In_320,In_563);
nor U1866 (N_1866,In_34,In_155);
nand U1867 (N_1867,In_709,In_130);
nor U1868 (N_1868,In_460,In_695);
nand U1869 (N_1869,In_226,In_626);
and U1870 (N_1870,In_846,In_886);
nand U1871 (N_1871,In_491,In_591);
or U1872 (N_1872,In_303,In_586);
nand U1873 (N_1873,In_656,In_395);
nand U1874 (N_1874,In_190,In_278);
or U1875 (N_1875,In_701,In_67);
xnor U1876 (N_1876,In_652,In_837);
nor U1877 (N_1877,In_562,In_788);
and U1878 (N_1878,In_465,In_871);
and U1879 (N_1879,In_419,In_658);
and U1880 (N_1880,In_451,In_259);
and U1881 (N_1881,In_726,In_181);
nand U1882 (N_1882,In_408,In_225);
nor U1883 (N_1883,In_802,In_248);
nor U1884 (N_1884,In_681,In_296);
and U1885 (N_1885,In_746,In_980);
nand U1886 (N_1886,In_54,In_832);
nor U1887 (N_1887,In_511,In_937);
or U1888 (N_1888,In_379,In_614);
or U1889 (N_1889,In_840,In_584);
nand U1890 (N_1890,In_896,In_842);
and U1891 (N_1891,In_216,In_366);
nand U1892 (N_1892,In_829,In_884);
or U1893 (N_1893,In_429,In_253);
nand U1894 (N_1894,In_250,In_857);
nor U1895 (N_1895,In_100,In_447);
xnor U1896 (N_1896,In_546,In_292);
and U1897 (N_1897,In_668,In_333);
and U1898 (N_1898,In_877,In_20);
or U1899 (N_1899,In_954,In_862);
nand U1900 (N_1900,In_38,In_884);
nor U1901 (N_1901,In_735,In_456);
xnor U1902 (N_1902,In_598,In_124);
xnor U1903 (N_1903,In_116,In_941);
or U1904 (N_1904,In_381,In_841);
and U1905 (N_1905,In_540,In_676);
nor U1906 (N_1906,In_12,In_919);
and U1907 (N_1907,In_569,In_896);
nor U1908 (N_1908,In_367,In_114);
nor U1909 (N_1909,In_675,In_198);
or U1910 (N_1910,In_645,In_73);
or U1911 (N_1911,In_396,In_947);
xor U1912 (N_1912,In_617,In_77);
xnor U1913 (N_1913,In_71,In_359);
and U1914 (N_1914,In_600,In_653);
or U1915 (N_1915,In_735,In_184);
nand U1916 (N_1916,In_533,In_352);
xnor U1917 (N_1917,In_554,In_368);
xor U1918 (N_1918,In_383,In_712);
nand U1919 (N_1919,In_807,In_479);
and U1920 (N_1920,In_822,In_76);
or U1921 (N_1921,In_384,In_382);
nand U1922 (N_1922,In_932,In_223);
nor U1923 (N_1923,In_675,In_368);
nand U1924 (N_1924,In_414,In_301);
nor U1925 (N_1925,In_117,In_563);
nor U1926 (N_1926,In_337,In_622);
xor U1927 (N_1927,In_420,In_278);
or U1928 (N_1928,In_928,In_197);
nand U1929 (N_1929,In_518,In_782);
nor U1930 (N_1930,In_575,In_755);
or U1931 (N_1931,In_799,In_235);
xnor U1932 (N_1932,In_189,In_38);
nand U1933 (N_1933,In_549,In_608);
and U1934 (N_1934,In_419,In_243);
or U1935 (N_1935,In_589,In_992);
xnor U1936 (N_1936,In_227,In_340);
and U1937 (N_1937,In_561,In_827);
nand U1938 (N_1938,In_583,In_896);
and U1939 (N_1939,In_668,In_104);
nand U1940 (N_1940,In_126,In_138);
and U1941 (N_1941,In_595,In_69);
and U1942 (N_1942,In_137,In_550);
and U1943 (N_1943,In_293,In_595);
xnor U1944 (N_1944,In_854,In_693);
or U1945 (N_1945,In_399,In_227);
or U1946 (N_1946,In_261,In_24);
or U1947 (N_1947,In_251,In_758);
nor U1948 (N_1948,In_465,In_512);
xor U1949 (N_1949,In_507,In_687);
nor U1950 (N_1950,In_465,In_951);
xor U1951 (N_1951,In_949,In_936);
nor U1952 (N_1952,In_123,In_35);
xnor U1953 (N_1953,In_19,In_388);
and U1954 (N_1954,In_252,In_77);
nor U1955 (N_1955,In_710,In_10);
or U1956 (N_1956,In_79,In_784);
nor U1957 (N_1957,In_843,In_553);
or U1958 (N_1958,In_692,In_597);
and U1959 (N_1959,In_738,In_352);
and U1960 (N_1960,In_743,In_793);
and U1961 (N_1961,In_381,In_622);
nor U1962 (N_1962,In_658,In_444);
xnor U1963 (N_1963,In_422,In_40);
nand U1964 (N_1964,In_860,In_761);
nor U1965 (N_1965,In_585,In_89);
or U1966 (N_1966,In_715,In_44);
and U1967 (N_1967,In_632,In_541);
xor U1968 (N_1968,In_277,In_221);
nor U1969 (N_1969,In_611,In_319);
xor U1970 (N_1970,In_298,In_769);
and U1971 (N_1971,In_924,In_843);
nand U1972 (N_1972,In_796,In_100);
and U1973 (N_1973,In_782,In_547);
nand U1974 (N_1974,In_767,In_928);
xnor U1975 (N_1975,In_418,In_611);
xor U1976 (N_1976,In_699,In_227);
nor U1977 (N_1977,In_187,In_661);
nand U1978 (N_1978,In_905,In_104);
or U1979 (N_1979,In_821,In_413);
xor U1980 (N_1980,In_149,In_194);
or U1981 (N_1981,In_250,In_969);
and U1982 (N_1982,In_460,In_401);
nand U1983 (N_1983,In_780,In_802);
nand U1984 (N_1984,In_531,In_136);
nor U1985 (N_1985,In_181,In_436);
nor U1986 (N_1986,In_612,In_843);
and U1987 (N_1987,In_332,In_632);
nand U1988 (N_1988,In_661,In_468);
nand U1989 (N_1989,In_344,In_862);
nand U1990 (N_1990,In_264,In_94);
xor U1991 (N_1991,In_322,In_85);
xor U1992 (N_1992,In_756,In_470);
nand U1993 (N_1993,In_832,In_371);
and U1994 (N_1994,In_969,In_859);
nor U1995 (N_1995,In_40,In_235);
xnor U1996 (N_1996,In_276,In_696);
nor U1997 (N_1997,In_936,In_758);
or U1998 (N_1998,In_192,In_832);
nand U1999 (N_1999,In_315,In_83);
nand U2000 (N_2000,In_790,In_6);
and U2001 (N_2001,In_322,In_786);
or U2002 (N_2002,In_667,In_886);
nor U2003 (N_2003,In_619,In_574);
nor U2004 (N_2004,In_426,In_549);
or U2005 (N_2005,In_727,In_502);
xor U2006 (N_2006,In_345,In_823);
nor U2007 (N_2007,In_177,In_225);
nor U2008 (N_2008,In_157,In_198);
or U2009 (N_2009,In_739,In_737);
or U2010 (N_2010,In_949,In_368);
and U2011 (N_2011,In_536,In_610);
nand U2012 (N_2012,In_330,In_905);
or U2013 (N_2013,In_571,In_450);
xor U2014 (N_2014,In_85,In_235);
nand U2015 (N_2015,In_180,In_845);
and U2016 (N_2016,In_575,In_647);
or U2017 (N_2017,In_862,In_941);
xor U2018 (N_2018,In_490,In_138);
nor U2019 (N_2019,In_151,In_721);
and U2020 (N_2020,In_326,In_61);
or U2021 (N_2021,In_494,In_352);
and U2022 (N_2022,In_74,In_568);
and U2023 (N_2023,In_375,In_476);
nand U2024 (N_2024,In_565,In_30);
nand U2025 (N_2025,In_889,In_331);
xnor U2026 (N_2026,In_437,In_907);
or U2027 (N_2027,In_682,In_934);
and U2028 (N_2028,In_661,In_349);
nand U2029 (N_2029,In_504,In_73);
xnor U2030 (N_2030,In_719,In_208);
xnor U2031 (N_2031,In_339,In_235);
and U2032 (N_2032,In_60,In_854);
nor U2033 (N_2033,In_624,In_514);
nand U2034 (N_2034,In_410,In_919);
or U2035 (N_2035,In_191,In_690);
nand U2036 (N_2036,In_402,In_674);
and U2037 (N_2037,In_345,In_99);
nor U2038 (N_2038,In_803,In_694);
xor U2039 (N_2039,In_579,In_533);
xnor U2040 (N_2040,In_812,In_14);
nand U2041 (N_2041,In_425,In_468);
and U2042 (N_2042,In_665,In_416);
nand U2043 (N_2043,In_141,In_693);
nor U2044 (N_2044,In_542,In_711);
nor U2045 (N_2045,In_213,In_942);
or U2046 (N_2046,In_606,In_413);
nor U2047 (N_2047,In_30,In_944);
or U2048 (N_2048,In_636,In_976);
xor U2049 (N_2049,In_534,In_42);
xor U2050 (N_2050,In_245,In_131);
nand U2051 (N_2051,In_624,In_520);
nand U2052 (N_2052,In_444,In_964);
nand U2053 (N_2053,In_301,In_844);
nor U2054 (N_2054,In_876,In_992);
xnor U2055 (N_2055,In_535,In_869);
or U2056 (N_2056,In_809,In_389);
xnor U2057 (N_2057,In_473,In_293);
nand U2058 (N_2058,In_152,In_244);
nor U2059 (N_2059,In_115,In_567);
or U2060 (N_2060,In_405,In_911);
or U2061 (N_2061,In_775,In_488);
or U2062 (N_2062,In_327,In_621);
nand U2063 (N_2063,In_328,In_313);
or U2064 (N_2064,In_621,In_747);
nand U2065 (N_2065,In_330,In_274);
xnor U2066 (N_2066,In_699,In_790);
nand U2067 (N_2067,In_675,In_832);
or U2068 (N_2068,In_440,In_119);
or U2069 (N_2069,In_170,In_794);
and U2070 (N_2070,In_610,In_664);
and U2071 (N_2071,In_50,In_527);
xor U2072 (N_2072,In_683,In_160);
nor U2073 (N_2073,In_38,In_610);
nor U2074 (N_2074,In_188,In_59);
xnor U2075 (N_2075,In_506,In_64);
nor U2076 (N_2076,In_9,In_76);
and U2077 (N_2077,In_377,In_542);
nand U2078 (N_2078,In_755,In_50);
and U2079 (N_2079,In_293,In_837);
and U2080 (N_2080,In_261,In_988);
nand U2081 (N_2081,In_361,In_673);
or U2082 (N_2082,In_520,In_895);
nand U2083 (N_2083,In_525,In_27);
nor U2084 (N_2084,In_477,In_379);
or U2085 (N_2085,In_506,In_995);
nand U2086 (N_2086,In_98,In_65);
nand U2087 (N_2087,In_175,In_409);
and U2088 (N_2088,In_332,In_422);
or U2089 (N_2089,In_571,In_865);
nor U2090 (N_2090,In_693,In_707);
or U2091 (N_2091,In_840,In_270);
or U2092 (N_2092,In_847,In_92);
or U2093 (N_2093,In_845,In_107);
nand U2094 (N_2094,In_739,In_126);
nand U2095 (N_2095,In_38,In_944);
nor U2096 (N_2096,In_285,In_641);
or U2097 (N_2097,In_62,In_785);
nand U2098 (N_2098,In_692,In_101);
nand U2099 (N_2099,In_603,In_296);
nor U2100 (N_2100,In_970,In_447);
nor U2101 (N_2101,In_54,In_0);
xnor U2102 (N_2102,In_790,In_526);
and U2103 (N_2103,In_812,In_56);
xnor U2104 (N_2104,In_165,In_67);
nand U2105 (N_2105,In_181,In_268);
and U2106 (N_2106,In_38,In_945);
or U2107 (N_2107,In_380,In_390);
nor U2108 (N_2108,In_590,In_199);
and U2109 (N_2109,In_340,In_790);
nand U2110 (N_2110,In_378,In_504);
or U2111 (N_2111,In_300,In_498);
xor U2112 (N_2112,In_58,In_710);
xnor U2113 (N_2113,In_665,In_724);
nand U2114 (N_2114,In_899,In_594);
xnor U2115 (N_2115,In_520,In_229);
and U2116 (N_2116,In_2,In_235);
or U2117 (N_2117,In_419,In_704);
or U2118 (N_2118,In_506,In_66);
nor U2119 (N_2119,In_556,In_373);
nor U2120 (N_2120,In_684,In_19);
and U2121 (N_2121,In_386,In_840);
and U2122 (N_2122,In_874,In_634);
or U2123 (N_2123,In_963,In_597);
xnor U2124 (N_2124,In_529,In_226);
and U2125 (N_2125,In_493,In_855);
and U2126 (N_2126,In_231,In_281);
nor U2127 (N_2127,In_239,In_388);
nor U2128 (N_2128,In_740,In_245);
nor U2129 (N_2129,In_412,In_600);
nand U2130 (N_2130,In_518,In_803);
nor U2131 (N_2131,In_697,In_457);
nand U2132 (N_2132,In_806,In_537);
nand U2133 (N_2133,In_926,In_427);
nand U2134 (N_2134,In_986,In_652);
and U2135 (N_2135,In_407,In_758);
nor U2136 (N_2136,In_247,In_297);
and U2137 (N_2137,In_403,In_204);
xnor U2138 (N_2138,In_186,In_478);
nor U2139 (N_2139,In_444,In_343);
nand U2140 (N_2140,In_473,In_197);
nand U2141 (N_2141,In_460,In_760);
and U2142 (N_2142,In_949,In_68);
and U2143 (N_2143,In_577,In_572);
nor U2144 (N_2144,In_242,In_383);
nand U2145 (N_2145,In_452,In_944);
nand U2146 (N_2146,In_473,In_985);
and U2147 (N_2147,In_175,In_350);
nor U2148 (N_2148,In_996,In_450);
and U2149 (N_2149,In_864,In_452);
nand U2150 (N_2150,In_689,In_448);
and U2151 (N_2151,In_229,In_406);
and U2152 (N_2152,In_318,In_817);
nor U2153 (N_2153,In_460,In_615);
nand U2154 (N_2154,In_635,In_721);
nand U2155 (N_2155,In_444,In_395);
or U2156 (N_2156,In_720,In_836);
or U2157 (N_2157,In_999,In_516);
nand U2158 (N_2158,In_986,In_750);
and U2159 (N_2159,In_123,In_971);
and U2160 (N_2160,In_627,In_511);
or U2161 (N_2161,In_994,In_542);
xor U2162 (N_2162,In_550,In_203);
or U2163 (N_2163,In_447,In_916);
xor U2164 (N_2164,In_416,In_506);
and U2165 (N_2165,In_611,In_334);
nand U2166 (N_2166,In_98,In_92);
or U2167 (N_2167,In_837,In_715);
nor U2168 (N_2168,In_700,In_360);
and U2169 (N_2169,In_973,In_219);
and U2170 (N_2170,In_48,In_774);
and U2171 (N_2171,In_616,In_270);
or U2172 (N_2172,In_445,In_372);
xnor U2173 (N_2173,In_701,In_633);
nor U2174 (N_2174,In_333,In_958);
nor U2175 (N_2175,In_52,In_609);
nand U2176 (N_2176,In_826,In_363);
nor U2177 (N_2177,In_88,In_20);
nor U2178 (N_2178,In_943,In_799);
or U2179 (N_2179,In_418,In_387);
or U2180 (N_2180,In_827,In_536);
xor U2181 (N_2181,In_784,In_863);
or U2182 (N_2182,In_711,In_628);
nor U2183 (N_2183,In_281,In_814);
and U2184 (N_2184,In_459,In_318);
nor U2185 (N_2185,In_683,In_838);
nor U2186 (N_2186,In_57,In_851);
nor U2187 (N_2187,In_730,In_259);
xor U2188 (N_2188,In_967,In_444);
or U2189 (N_2189,In_797,In_37);
and U2190 (N_2190,In_722,In_177);
nor U2191 (N_2191,In_938,In_613);
or U2192 (N_2192,In_352,In_195);
nor U2193 (N_2193,In_722,In_37);
nor U2194 (N_2194,In_637,In_800);
nor U2195 (N_2195,In_124,In_483);
and U2196 (N_2196,In_207,In_794);
nand U2197 (N_2197,In_46,In_822);
or U2198 (N_2198,In_840,In_572);
or U2199 (N_2199,In_168,In_324);
xnor U2200 (N_2200,In_906,In_8);
nand U2201 (N_2201,In_357,In_863);
nor U2202 (N_2202,In_130,In_463);
nor U2203 (N_2203,In_262,In_998);
xor U2204 (N_2204,In_707,In_802);
xnor U2205 (N_2205,In_515,In_0);
xnor U2206 (N_2206,In_462,In_813);
and U2207 (N_2207,In_861,In_953);
xor U2208 (N_2208,In_547,In_650);
or U2209 (N_2209,In_206,In_86);
xnor U2210 (N_2210,In_26,In_957);
nand U2211 (N_2211,In_988,In_249);
and U2212 (N_2212,In_202,In_986);
and U2213 (N_2213,In_21,In_545);
nor U2214 (N_2214,In_637,In_312);
nor U2215 (N_2215,In_961,In_614);
nor U2216 (N_2216,In_660,In_128);
and U2217 (N_2217,In_648,In_707);
nand U2218 (N_2218,In_9,In_880);
nor U2219 (N_2219,In_187,In_207);
xnor U2220 (N_2220,In_202,In_237);
and U2221 (N_2221,In_29,In_172);
nand U2222 (N_2222,In_786,In_307);
xor U2223 (N_2223,In_175,In_293);
xnor U2224 (N_2224,In_660,In_599);
xnor U2225 (N_2225,In_894,In_262);
or U2226 (N_2226,In_159,In_350);
nand U2227 (N_2227,In_948,In_690);
nand U2228 (N_2228,In_928,In_695);
nand U2229 (N_2229,In_44,In_930);
and U2230 (N_2230,In_493,In_928);
nand U2231 (N_2231,In_444,In_338);
xnor U2232 (N_2232,In_440,In_735);
nand U2233 (N_2233,In_264,In_327);
nor U2234 (N_2234,In_847,In_55);
or U2235 (N_2235,In_504,In_180);
xor U2236 (N_2236,In_634,In_128);
and U2237 (N_2237,In_327,In_572);
xor U2238 (N_2238,In_259,In_947);
nand U2239 (N_2239,In_257,In_214);
and U2240 (N_2240,In_198,In_816);
or U2241 (N_2241,In_603,In_563);
xnor U2242 (N_2242,In_292,In_993);
and U2243 (N_2243,In_738,In_879);
and U2244 (N_2244,In_503,In_516);
or U2245 (N_2245,In_70,In_143);
nor U2246 (N_2246,In_418,In_114);
nor U2247 (N_2247,In_123,In_395);
xnor U2248 (N_2248,In_638,In_468);
and U2249 (N_2249,In_825,In_830);
nor U2250 (N_2250,In_166,In_154);
and U2251 (N_2251,In_267,In_326);
or U2252 (N_2252,In_653,In_664);
and U2253 (N_2253,In_906,In_506);
nand U2254 (N_2254,In_631,In_614);
nor U2255 (N_2255,In_59,In_744);
and U2256 (N_2256,In_579,In_475);
nand U2257 (N_2257,In_809,In_595);
nor U2258 (N_2258,In_700,In_221);
nor U2259 (N_2259,In_517,In_143);
nand U2260 (N_2260,In_124,In_485);
xor U2261 (N_2261,In_109,In_447);
and U2262 (N_2262,In_46,In_440);
nor U2263 (N_2263,In_837,In_196);
or U2264 (N_2264,In_671,In_896);
nand U2265 (N_2265,In_113,In_102);
nand U2266 (N_2266,In_523,In_99);
or U2267 (N_2267,In_915,In_867);
and U2268 (N_2268,In_24,In_914);
and U2269 (N_2269,In_270,In_798);
or U2270 (N_2270,In_98,In_978);
and U2271 (N_2271,In_469,In_343);
nor U2272 (N_2272,In_191,In_116);
nor U2273 (N_2273,In_572,In_157);
nor U2274 (N_2274,In_682,In_553);
or U2275 (N_2275,In_556,In_661);
xnor U2276 (N_2276,In_968,In_428);
or U2277 (N_2277,In_346,In_313);
xnor U2278 (N_2278,In_609,In_544);
nand U2279 (N_2279,In_660,In_624);
nand U2280 (N_2280,In_213,In_504);
or U2281 (N_2281,In_523,In_472);
xnor U2282 (N_2282,In_563,In_713);
xnor U2283 (N_2283,In_368,In_247);
nand U2284 (N_2284,In_273,In_930);
nand U2285 (N_2285,In_467,In_290);
nand U2286 (N_2286,In_332,In_440);
and U2287 (N_2287,In_796,In_204);
xnor U2288 (N_2288,In_49,In_33);
and U2289 (N_2289,In_336,In_376);
nor U2290 (N_2290,In_158,In_308);
xor U2291 (N_2291,In_465,In_578);
nand U2292 (N_2292,In_346,In_789);
nand U2293 (N_2293,In_607,In_774);
nand U2294 (N_2294,In_298,In_428);
nor U2295 (N_2295,In_274,In_364);
nand U2296 (N_2296,In_204,In_334);
xnor U2297 (N_2297,In_903,In_977);
nand U2298 (N_2298,In_613,In_875);
and U2299 (N_2299,In_931,In_923);
nand U2300 (N_2300,In_956,In_129);
and U2301 (N_2301,In_366,In_597);
xor U2302 (N_2302,In_217,In_648);
or U2303 (N_2303,In_412,In_448);
xnor U2304 (N_2304,In_286,In_61);
or U2305 (N_2305,In_377,In_533);
nand U2306 (N_2306,In_609,In_503);
and U2307 (N_2307,In_464,In_602);
nand U2308 (N_2308,In_45,In_947);
nand U2309 (N_2309,In_348,In_925);
or U2310 (N_2310,In_154,In_391);
xnor U2311 (N_2311,In_137,In_483);
or U2312 (N_2312,In_166,In_669);
nor U2313 (N_2313,In_121,In_973);
or U2314 (N_2314,In_448,In_65);
or U2315 (N_2315,In_664,In_382);
nand U2316 (N_2316,In_374,In_677);
xor U2317 (N_2317,In_908,In_657);
and U2318 (N_2318,In_172,In_199);
nand U2319 (N_2319,In_304,In_526);
and U2320 (N_2320,In_686,In_292);
or U2321 (N_2321,In_298,In_205);
nor U2322 (N_2322,In_251,In_444);
nand U2323 (N_2323,In_92,In_322);
xnor U2324 (N_2324,In_114,In_146);
nand U2325 (N_2325,In_781,In_647);
nor U2326 (N_2326,In_484,In_159);
nand U2327 (N_2327,In_235,In_596);
and U2328 (N_2328,In_792,In_484);
and U2329 (N_2329,In_857,In_186);
and U2330 (N_2330,In_22,In_21);
or U2331 (N_2331,In_658,In_316);
or U2332 (N_2332,In_560,In_639);
or U2333 (N_2333,In_282,In_182);
xnor U2334 (N_2334,In_221,In_578);
or U2335 (N_2335,In_735,In_773);
nor U2336 (N_2336,In_512,In_479);
and U2337 (N_2337,In_267,In_995);
and U2338 (N_2338,In_284,In_202);
nand U2339 (N_2339,In_360,In_866);
or U2340 (N_2340,In_234,In_920);
xnor U2341 (N_2341,In_636,In_621);
nand U2342 (N_2342,In_552,In_473);
xnor U2343 (N_2343,In_255,In_157);
and U2344 (N_2344,In_981,In_117);
nor U2345 (N_2345,In_395,In_324);
and U2346 (N_2346,In_615,In_722);
xnor U2347 (N_2347,In_437,In_407);
nor U2348 (N_2348,In_835,In_316);
nand U2349 (N_2349,In_653,In_875);
nand U2350 (N_2350,In_859,In_697);
nand U2351 (N_2351,In_686,In_11);
nor U2352 (N_2352,In_702,In_53);
or U2353 (N_2353,In_315,In_584);
nand U2354 (N_2354,In_764,In_679);
and U2355 (N_2355,In_146,In_936);
xnor U2356 (N_2356,In_882,In_205);
nand U2357 (N_2357,In_586,In_836);
and U2358 (N_2358,In_444,In_493);
xnor U2359 (N_2359,In_229,In_726);
nor U2360 (N_2360,In_150,In_345);
xnor U2361 (N_2361,In_708,In_427);
or U2362 (N_2362,In_793,In_411);
xor U2363 (N_2363,In_754,In_604);
or U2364 (N_2364,In_600,In_116);
or U2365 (N_2365,In_10,In_766);
xnor U2366 (N_2366,In_760,In_413);
xor U2367 (N_2367,In_706,In_447);
nand U2368 (N_2368,In_269,In_175);
nand U2369 (N_2369,In_686,In_491);
nand U2370 (N_2370,In_951,In_314);
or U2371 (N_2371,In_247,In_31);
nand U2372 (N_2372,In_404,In_386);
or U2373 (N_2373,In_228,In_316);
xor U2374 (N_2374,In_105,In_41);
xnor U2375 (N_2375,In_317,In_49);
nor U2376 (N_2376,In_447,In_59);
nor U2377 (N_2377,In_706,In_928);
and U2378 (N_2378,In_124,In_746);
nor U2379 (N_2379,In_172,In_616);
nor U2380 (N_2380,In_7,In_147);
or U2381 (N_2381,In_977,In_337);
or U2382 (N_2382,In_736,In_173);
xnor U2383 (N_2383,In_484,In_908);
or U2384 (N_2384,In_151,In_179);
nand U2385 (N_2385,In_162,In_395);
and U2386 (N_2386,In_997,In_514);
or U2387 (N_2387,In_584,In_119);
nand U2388 (N_2388,In_993,In_46);
nor U2389 (N_2389,In_803,In_87);
xnor U2390 (N_2390,In_41,In_729);
and U2391 (N_2391,In_493,In_328);
or U2392 (N_2392,In_762,In_773);
or U2393 (N_2393,In_781,In_596);
nand U2394 (N_2394,In_500,In_675);
and U2395 (N_2395,In_213,In_427);
nand U2396 (N_2396,In_776,In_373);
nor U2397 (N_2397,In_164,In_934);
and U2398 (N_2398,In_591,In_824);
nand U2399 (N_2399,In_833,In_497);
nor U2400 (N_2400,In_577,In_897);
nor U2401 (N_2401,In_850,In_6);
xor U2402 (N_2402,In_256,In_561);
or U2403 (N_2403,In_598,In_975);
xor U2404 (N_2404,In_850,In_250);
nor U2405 (N_2405,In_360,In_832);
nor U2406 (N_2406,In_575,In_675);
or U2407 (N_2407,In_715,In_258);
xor U2408 (N_2408,In_682,In_895);
nand U2409 (N_2409,In_662,In_942);
or U2410 (N_2410,In_63,In_74);
nor U2411 (N_2411,In_80,In_618);
xnor U2412 (N_2412,In_736,In_549);
and U2413 (N_2413,In_490,In_715);
and U2414 (N_2414,In_598,In_252);
nand U2415 (N_2415,In_89,In_348);
or U2416 (N_2416,In_54,In_74);
or U2417 (N_2417,In_863,In_713);
nor U2418 (N_2418,In_773,In_138);
and U2419 (N_2419,In_576,In_717);
and U2420 (N_2420,In_659,In_953);
xor U2421 (N_2421,In_313,In_971);
nand U2422 (N_2422,In_328,In_900);
or U2423 (N_2423,In_966,In_639);
xnor U2424 (N_2424,In_184,In_647);
xor U2425 (N_2425,In_602,In_424);
nor U2426 (N_2426,In_84,In_401);
nor U2427 (N_2427,In_998,In_673);
xor U2428 (N_2428,In_568,In_830);
nor U2429 (N_2429,In_174,In_583);
or U2430 (N_2430,In_632,In_368);
nor U2431 (N_2431,In_41,In_944);
and U2432 (N_2432,In_513,In_789);
nor U2433 (N_2433,In_999,In_665);
nand U2434 (N_2434,In_971,In_34);
or U2435 (N_2435,In_819,In_372);
and U2436 (N_2436,In_11,In_882);
xnor U2437 (N_2437,In_239,In_677);
or U2438 (N_2438,In_717,In_818);
and U2439 (N_2439,In_620,In_140);
nand U2440 (N_2440,In_951,In_358);
or U2441 (N_2441,In_970,In_904);
or U2442 (N_2442,In_85,In_527);
xnor U2443 (N_2443,In_439,In_212);
nor U2444 (N_2444,In_413,In_673);
nor U2445 (N_2445,In_556,In_47);
nor U2446 (N_2446,In_339,In_279);
nand U2447 (N_2447,In_865,In_429);
nand U2448 (N_2448,In_670,In_633);
nand U2449 (N_2449,In_630,In_367);
xor U2450 (N_2450,In_664,In_484);
or U2451 (N_2451,In_768,In_749);
and U2452 (N_2452,In_824,In_84);
xnor U2453 (N_2453,In_696,In_863);
and U2454 (N_2454,In_546,In_576);
xor U2455 (N_2455,In_205,In_278);
nand U2456 (N_2456,In_685,In_429);
or U2457 (N_2457,In_306,In_287);
and U2458 (N_2458,In_961,In_601);
xnor U2459 (N_2459,In_205,In_875);
nor U2460 (N_2460,In_224,In_24);
nand U2461 (N_2461,In_373,In_618);
nor U2462 (N_2462,In_569,In_246);
nor U2463 (N_2463,In_450,In_338);
nand U2464 (N_2464,In_817,In_7);
or U2465 (N_2465,In_437,In_450);
xor U2466 (N_2466,In_722,In_793);
xor U2467 (N_2467,In_417,In_598);
xor U2468 (N_2468,In_839,In_869);
nor U2469 (N_2469,In_814,In_872);
xnor U2470 (N_2470,In_309,In_191);
xnor U2471 (N_2471,In_892,In_715);
nand U2472 (N_2472,In_239,In_343);
nor U2473 (N_2473,In_299,In_920);
nor U2474 (N_2474,In_368,In_176);
xnor U2475 (N_2475,In_198,In_615);
xor U2476 (N_2476,In_114,In_175);
or U2477 (N_2477,In_822,In_908);
or U2478 (N_2478,In_100,In_671);
nand U2479 (N_2479,In_693,In_858);
and U2480 (N_2480,In_187,In_103);
nor U2481 (N_2481,In_508,In_496);
xnor U2482 (N_2482,In_998,In_921);
or U2483 (N_2483,In_120,In_856);
and U2484 (N_2484,In_945,In_93);
nor U2485 (N_2485,In_756,In_516);
nor U2486 (N_2486,In_363,In_194);
nand U2487 (N_2487,In_581,In_351);
or U2488 (N_2488,In_660,In_253);
nor U2489 (N_2489,In_937,In_298);
nor U2490 (N_2490,In_373,In_26);
nor U2491 (N_2491,In_137,In_375);
and U2492 (N_2492,In_239,In_971);
nand U2493 (N_2493,In_680,In_103);
nand U2494 (N_2494,In_884,In_34);
or U2495 (N_2495,In_122,In_321);
xor U2496 (N_2496,In_802,In_483);
nor U2497 (N_2497,In_637,In_308);
or U2498 (N_2498,In_886,In_95);
xor U2499 (N_2499,In_83,In_758);
nor U2500 (N_2500,In_222,In_612);
xor U2501 (N_2501,In_331,In_221);
nor U2502 (N_2502,In_853,In_94);
xnor U2503 (N_2503,In_360,In_372);
nand U2504 (N_2504,In_572,In_546);
xor U2505 (N_2505,In_981,In_257);
nand U2506 (N_2506,In_955,In_499);
or U2507 (N_2507,In_403,In_110);
and U2508 (N_2508,In_85,In_804);
xnor U2509 (N_2509,In_548,In_60);
nor U2510 (N_2510,In_360,In_636);
nand U2511 (N_2511,In_487,In_172);
or U2512 (N_2512,In_856,In_718);
nor U2513 (N_2513,In_702,In_812);
or U2514 (N_2514,In_718,In_525);
nor U2515 (N_2515,In_493,In_829);
nor U2516 (N_2516,In_654,In_172);
or U2517 (N_2517,In_482,In_585);
xnor U2518 (N_2518,In_202,In_43);
nor U2519 (N_2519,In_318,In_342);
or U2520 (N_2520,In_744,In_561);
and U2521 (N_2521,In_190,In_928);
xor U2522 (N_2522,In_680,In_515);
nor U2523 (N_2523,In_619,In_883);
and U2524 (N_2524,In_111,In_418);
nor U2525 (N_2525,In_633,In_246);
nand U2526 (N_2526,In_906,In_379);
xor U2527 (N_2527,In_528,In_51);
or U2528 (N_2528,In_411,In_716);
nand U2529 (N_2529,In_39,In_304);
nor U2530 (N_2530,In_517,In_237);
nor U2531 (N_2531,In_73,In_990);
and U2532 (N_2532,In_628,In_677);
nor U2533 (N_2533,In_110,In_138);
nand U2534 (N_2534,In_945,In_335);
or U2535 (N_2535,In_637,In_995);
nand U2536 (N_2536,In_88,In_771);
xnor U2537 (N_2537,In_557,In_402);
nand U2538 (N_2538,In_88,In_803);
and U2539 (N_2539,In_219,In_774);
or U2540 (N_2540,In_412,In_302);
nor U2541 (N_2541,In_389,In_846);
and U2542 (N_2542,In_446,In_717);
nor U2543 (N_2543,In_218,In_492);
nand U2544 (N_2544,In_328,In_16);
xnor U2545 (N_2545,In_376,In_862);
xor U2546 (N_2546,In_416,In_779);
nor U2547 (N_2547,In_845,In_710);
nor U2548 (N_2548,In_125,In_446);
xor U2549 (N_2549,In_438,In_607);
or U2550 (N_2550,In_506,In_486);
nand U2551 (N_2551,In_714,In_923);
nand U2552 (N_2552,In_161,In_208);
or U2553 (N_2553,In_386,In_79);
xor U2554 (N_2554,In_982,In_207);
nor U2555 (N_2555,In_405,In_37);
xnor U2556 (N_2556,In_200,In_563);
and U2557 (N_2557,In_78,In_73);
or U2558 (N_2558,In_304,In_982);
nand U2559 (N_2559,In_353,In_909);
nand U2560 (N_2560,In_801,In_389);
xnor U2561 (N_2561,In_884,In_280);
xor U2562 (N_2562,In_433,In_158);
or U2563 (N_2563,In_421,In_749);
and U2564 (N_2564,In_768,In_850);
and U2565 (N_2565,In_45,In_261);
or U2566 (N_2566,In_270,In_124);
nor U2567 (N_2567,In_289,In_362);
and U2568 (N_2568,In_442,In_467);
xnor U2569 (N_2569,In_399,In_320);
or U2570 (N_2570,In_844,In_848);
nor U2571 (N_2571,In_515,In_84);
nor U2572 (N_2572,In_476,In_680);
or U2573 (N_2573,In_325,In_435);
or U2574 (N_2574,In_874,In_454);
nor U2575 (N_2575,In_762,In_72);
nand U2576 (N_2576,In_362,In_992);
nand U2577 (N_2577,In_524,In_543);
nand U2578 (N_2578,In_115,In_347);
or U2579 (N_2579,In_902,In_962);
nor U2580 (N_2580,In_757,In_121);
and U2581 (N_2581,In_304,In_644);
nor U2582 (N_2582,In_146,In_656);
nor U2583 (N_2583,In_813,In_930);
nand U2584 (N_2584,In_648,In_93);
or U2585 (N_2585,In_600,In_594);
and U2586 (N_2586,In_24,In_127);
xnor U2587 (N_2587,In_559,In_812);
and U2588 (N_2588,In_264,In_782);
nand U2589 (N_2589,In_827,In_672);
xor U2590 (N_2590,In_642,In_168);
nand U2591 (N_2591,In_693,In_23);
or U2592 (N_2592,In_828,In_413);
or U2593 (N_2593,In_746,In_825);
or U2594 (N_2594,In_597,In_719);
and U2595 (N_2595,In_509,In_514);
xor U2596 (N_2596,In_838,In_76);
xnor U2597 (N_2597,In_41,In_14);
or U2598 (N_2598,In_702,In_961);
nand U2599 (N_2599,In_693,In_423);
or U2600 (N_2600,In_182,In_240);
xor U2601 (N_2601,In_962,In_467);
or U2602 (N_2602,In_149,In_165);
nand U2603 (N_2603,In_988,In_55);
and U2604 (N_2604,In_308,In_749);
nand U2605 (N_2605,In_377,In_207);
nand U2606 (N_2606,In_492,In_670);
nand U2607 (N_2607,In_591,In_252);
nor U2608 (N_2608,In_142,In_496);
nand U2609 (N_2609,In_80,In_788);
nor U2610 (N_2610,In_196,In_272);
and U2611 (N_2611,In_662,In_19);
or U2612 (N_2612,In_994,In_693);
nand U2613 (N_2613,In_253,In_436);
nor U2614 (N_2614,In_579,In_45);
or U2615 (N_2615,In_63,In_746);
nand U2616 (N_2616,In_135,In_490);
xor U2617 (N_2617,In_824,In_635);
nand U2618 (N_2618,In_566,In_666);
and U2619 (N_2619,In_611,In_492);
or U2620 (N_2620,In_371,In_337);
xor U2621 (N_2621,In_22,In_785);
and U2622 (N_2622,In_457,In_682);
xor U2623 (N_2623,In_978,In_328);
xor U2624 (N_2624,In_73,In_960);
xnor U2625 (N_2625,In_419,In_75);
xor U2626 (N_2626,In_890,In_302);
nand U2627 (N_2627,In_370,In_15);
xnor U2628 (N_2628,In_757,In_74);
nor U2629 (N_2629,In_440,In_794);
xor U2630 (N_2630,In_829,In_284);
and U2631 (N_2631,In_259,In_644);
or U2632 (N_2632,In_50,In_358);
nand U2633 (N_2633,In_647,In_669);
xor U2634 (N_2634,In_914,In_184);
xnor U2635 (N_2635,In_992,In_314);
nand U2636 (N_2636,In_897,In_258);
nand U2637 (N_2637,In_966,In_784);
or U2638 (N_2638,In_46,In_782);
nor U2639 (N_2639,In_198,In_291);
and U2640 (N_2640,In_31,In_681);
nor U2641 (N_2641,In_173,In_576);
and U2642 (N_2642,In_687,In_656);
nor U2643 (N_2643,In_70,In_545);
or U2644 (N_2644,In_101,In_998);
xnor U2645 (N_2645,In_816,In_679);
nand U2646 (N_2646,In_971,In_344);
nand U2647 (N_2647,In_466,In_141);
or U2648 (N_2648,In_736,In_275);
xor U2649 (N_2649,In_511,In_980);
xor U2650 (N_2650,In_430,In_161);
or U2651 (N_2651,In_591,In_124);
nor U2652 (N_2652,In_984,In_71);
nand U2653 (N_2653,In_788,In_807);
nor U2654 (N_2654,In_455,In_551);
nand U2655 (N_2655,In_176,In_878);
nand U2656 (N_2656,In_223,In_241);
or U2657 (N_2657,In_8,In_485);
nand U2658 (N_2658,In_927,In_346);
or U2659 (N_2659,In_280,In_978);
nand U2660 (N_2660,In_676,In_614);
nand U2661 (N_2661,In_779,In_8);
nand U2662 (N_2662,In_792,In_500);
and U2663 (N_2663,In_192,In_755);
and U2664 (N_2664,In_625,In_522);
nand U2665 (N_2665,In_953,In_232);
or U2666 (N_2666,In_822,In_409);
and U2667 (N_2667,In_811,In_778);
nor U2668 (N_2668,In_477,In_998);
nor U2669 (N_2669,In_580,In_501);
nand U2670 (N_2670,In_672,In_353);
and U2671 (N_2671,In_268,In_262);
or U2672 (N_2672,In_419,In_304);
nor U2673 (N_2673,In_924,In_365);
nor U2674 (N_2674,In_725,In_988);
nor U2675 (N_2675,In_747,In_777);
xor U2676 (N_2676,In_620,In_462);
and U2677 (N_2677,In_74,In_801);
nand U2678 (N_2678,In_439,In_409);
and U2679 (N_2679,In_303,In_13);
xnor U2680 (N_2680,In_691,In_563);
xnor U2681 (N_2681,In_671,In_878);
and U2682 (N_2682,In_14,In_325);
and U2683 (N_2683,In_561,In_247);
or U2684 (N_2684,In_574,In_70);
nand U2685 (N_2685,In_179,In_164);
or U2686 (N_2686,In_368,In_425);
nand U2687 (N_2687,In_757,In_733);
and U2688 (N_2688,In_299,In_840);
xor U2689 (N_2689,In_155,In_491);
and U2690 (N_2690,In_847,In_161);
or U2691 (N_2691,In_519,In_991);
or U2692 (N_2692,In_633,In_868);
nor U2693 (N_2693,In_466,In_717);
and U2694 (N_2694,In_112,In_204);
nand U2695 (N_2695,In_285,In_972);
nand U2696 (N_2696,In_893,In_566);
and U2697 (N_2697,In_534,In_570);
nor U2698 (N_2698,In_82,In_46);
and U2699 (N_2699,In_719,In_316);
or U2700 (N_2700,In_708,In_420);
or U2701 (N_2701,In_971,In_320);
nand U2702 (N_2702,In_593,In_299);
nor U2703 (N_2703,In_506,In_630);
or U2704 (N_2704,In_338,In_133);
nand U2705 (N_2705,In_494,In_601);
and U2706 (N_2706,In_507,In_70);
or U2707 (N_2707,In_722,In_208);
xnor U2708 (N_2708,In_657,In_982);
nand U2709 (N_2709,In_995,In_82);
nor U2710 (N_2710,In_159,In_722);
xor U2711 (N_2711,In_135,In_174);
xnor U2712 (N_2712,In_213,In_75);
xnor U2713 (N_2713,In_925,In_605);
nor U2714 (N_2714,In_393,In_688);
and U2715 (N_2715,In_167,In_717);
nand U2716 (N_2716,In_712,In_506);
or U2717 (N_2717,In_749,In_140);
or U2718 (N_2718,In_309,In_810);
nor U2719 (N_2719,In_552,In_844);
nor U2720 (N_2720,In_174,In_375);
nand U2721 (N_2721,In_536,In_166);
and U2722 (N_2722,In_159,In_587);
nand U2723 (N_2723,In_9,In_601);
or U2724 (N_2724,In_100,In_664);
and U2725 (N_2725,In_481,In_775);
nor U2726 (N_2726,In_68,In_715);
nor U2727 (N_2727,In_920,In_954);
nor U2728 (N_2728,In_845,In_115);
nor U2729 (N_2729,In_993,In_997);
xor U2730 (N_2730,In_319,In_65);
nor U2731 (N_2731,In_444,In_908);
nor U2732 (N_2732,In_510,In_257);
and U2733 (N_2733,In_656,In_473);
and U2734 (N_2734,In_75,In_318);
or U2735 (N_2735,In_566,In_109);
nand U2736 (N_2736,In_104,In_464);
nor U2737 (N_2737,In_609,In_24);
and U2738 (N_2738,In_4,In_721);
nor U2739 (N_2739,In_362,In_367);
and U2740 (N_2740,In_31,In_127);
or U2741 (N_2741,In_832,In_450);
and U2742 (N_2742,In_329,In_217);
xnor U2743 (N_2743,In_728,In_807);
nand U2744 (N_2744,In_202,In_557);
xor U2745 (N_2745,In_732,In_107);
and U2746 (N_2746,In_552,In_461);
nor U2747 (N_2747,In_966,In_633);
and U2748 (N_2748,In_477,In_978);
nor U2749 (N_2749,In_342,In_368);
or U2750 (N_2750,In_875,In_337);
nand U2751 (N_2751,In_664,In_855);
xor U2752 (N_2752,In_328,In_834);
and U2753 (N_2753,In_214,In_79);
or U2754 (N_2754,In_932,In_83);
xnor U2755 (N_2755,In_382,In_189);
xor U2756 (N_2756,In_685,In_892);
xor U2757 (N_2757,In_194,In_781);
or U2758 (N_2758,In_298,In_162);
xor U2759 (N_2759,In_642,In_774);
nand U2760 (N_2760,In_913,In_967);
and U2761 (N_2761,In_43,In_267);
xor U2762 (N_2762,In_803,In_763);
or U2763 (N_2763,In_987,In_588);
or U2764 (N_2764,In_745,In_540);
or U2765 (N_2765,In_95,In_897);
and U2766 (N_2766,In_564,In_216);
xnor U2767 (N_2767,In_697,In_80);
nor U2768 (N_2768,In_743,In_794);
xor U2769 (N_2769,In_118,In_948);
and U2770 (N_2770,In_71,In_270);
and U2771 (N_2771,In_621,In_701);
nand U2772 (N_2772,In_86,In_783);
or U2773 (N_2773,In_510,In_277);
xor U2774 (N_2774,In_105,In_210);
and U2775 (N_2775,In_749,In_322);
xnor U2776 (N_2776,In_73,In_571);
xor U2777 (N_2777,In_410,In_237);
nand U2778 (N_2778,In_863,In_463);
nand U2779 (N_2779,In_349,In_184);
and U2780 (N_2780,In_574,In_917);
nor U2781 (N_2781,In_17,In_434);
and U2782 (N_2782,In_512,In_177);
or U2783 (N_2783,In_2,In_192);
or U2784 (N_2784,In_818,In_785);
and U2785 (N_2785,In_8,In_638);
and U2786 (N_2786,In_548,In_829);
xor U2787 (N_2787,In_600,In_652);
nand U2788 (N_2788,In_102,In_814);
nand U2789 (N_2789,In_355,In_480);
and U2790 (N_2790,In_310,In_808);
nor U2791 (N_2791,In_421,In_589);
nor U2792 (N_2792,In_801,In_214);
or U2793 (N_2793,In_341,In_638);
nand U2794 (N_2794,In_186,In_837);
nor U2795 (N_2795,In_834,In_277);
nand U2796 (N_2796,In_387,In_333);
nand U2797 (N_2797,In_550,In_918);
and U2798 (N_2798,In_897,In_233);
nand U2799 (N_2799,In_225,In_354);
nor U2800 (N_2800,In_672,In_159);
and U2801 (N_2801,In_601,In_224);
xnor U2802 (N_2802,In_800,In_229);
nand U2803 (N_2803,In_644,In_375);
nor U2804 (N_2804,In_76,In_520);
or U2805 (N_2805,In_596,In_750);
xor U2806 (N_2806,In_638,In_591);
nand U2807 (N_2807,In_16,In_683);
nor U2808 (N_2808,In_110,In_432);
and U2809 (N_2809,In_682,In_109);
nor U2810 (N_2810,In_791,In_561);
nor U2811 (N_2811,In_128,In_853);
and U2812 (N_2812,In_705,In_147);
nand U2813 (N_2813,In_361,In_814);
xor U2814 (N_2814,In_515,In_964);
xnor U2815 (N_2815,In_394,In_498);
or U2816 (N_2816,In_81,In_380);
xor U2817 (N_2817,In_100,In_911);
nor U2818 (N_2818,In_904,In_187);
nor U2819 (N_2819,In_352,In_685);
and U2820 (N_2820,In_334,In_484);
nor U2821 (N_2821,In_906,In_220);
nand U2822 (N_2822,In_905,In_758);
nor U2823 (N_2823,In_377,In_459);
and U2824 (N_2824,In_493,In_412);
xnor U2825 (N_2825,In_787,In_890);
nor U2826 (N_2826,In_896,In_904);
and U2827 (N_2827,In_95,In_827);
and U2828 (N_2828,In_290,In_268);
nor U2829 (N_2829,In_486,In_33);
or U2830 (N_2830,In_394,In_628);
or U2831 (N_2831,In_943,In_53);
or U2832 (N_2832,In_325,In_978);
nand U2833 (N_2833,In_7,In_152);
xnor U2834 (N_2834,In_500,In_255);
nor U2835 (N_2835,In_10,In_518);
nor U2836 (N_2836,In_281,In_598);
nand U2837 (N_2837,In_462,In_608);
xnor U2838 (N_2838,In_329,In_854);
xor U2839 (N_2839,In_22,In_140);
xor U2840 (N_2840,In_683,In_943);
nand U2841 (N_2841,In_358,In_45);
nor U2842 (N_2842,In_407,In_164);
and U2843 (N_2843,In_545,In_0);
nand U2844 (N_2844,In_485,In_446);
or U2845 (N_2845,In_752,In_14);
xor U2846 (N_2846,In_846,In_189);
nand U2847 (N_2847,In_538,In_849);
xnor U2848 (N_2848,In_716,In_900);
and U2849 (N_2849,In_5,In_573);
or U2850 (N_2850,In_0,In_687);
nor U2851 (N_2851,In_480,In_58);
xnor U2852 (N_2852,In_368,In_367);
or U2853 (N_2853,In_53,In_475);
nor U2854 (N_2854,In_764,In_328);
nand U2855 (N_2855,In_332,In_765);
and U2856 (N_2856,In_725,In_49);
xnor U2857 (N_2857,In_505,In_916);
or U2858 (N_2858,In_154,In_399);
or U2859 (N_2859,In_522,In_563);
and U2860 (N_2860,In_979,In_511);
or U2861 (N_2861,In_456,In_916);
xor U2862 (N_2862,In_664,In_416);
nor U2863 (N_2863,In_662,In_690);
or U2864 (N_2864,In_866,In_138);
or U2865 (N_2865,In_304,In_730);
nor U2866 (N_2866,In_115,In_426);
nand U2867 (N_2867,In_592,In_22);
or U2868 (N_2868,In_440,In_374);
and U2869 (N_2869,In_507,In_673);
nor U2870 (N_2870,In_591,In_273);
nand U2871 (N_2871,In_922,In_876);
nand U2872 (N_2872,In_393,In_891);
xor U2873 (N_2873,In_930,In_27);
nor U2874 (N_2874,In_8,In_456);
nor U2875 (N_2875,In_392,In_711);
or U2876 (N_2876,In_842,In_748);
nand U2877 (N_2877,In_309,In_590);
xor U2878 (N_2878,In_366,In_70);
nor U2879 (N_2879,In_178,In_818);
nand U2880 (N_2880,In_521,In_698);
or U2881 (N_2881,In_363,In_357);
xor U2882 (N_2882,In_48,In_814);
xor U2883 (N_2883,In_601,In_901);
nand U2884 (N_2884,In_268,In_588);
nor U2885 (N_2885,In_792,In_264);
xnor U2886 (N_2886,In_737,In_385);
xnor U2887 (N_2887,In_397,In_390);
nor U2888 (N_2888,In_533,In_13);
or U2889 (N_2889,In_275,In_607);
and U2890 (N_2890,In_945,In_67);
nand U2891 (N_2891,In_338,In_620);
and U2892 (N_2892,In_664,In_429);
or U2893 (N_2893,In_42,In_288);
nand U2894 (N_2894,In_939,In_457);
nor U2895 (N_2895,In_76,In_734);
nor U2896 (N_2896,In_775,In_765);
and U2897 (N_2897,In_497,In_857);
nand U2898 (N_2898,In_721,In_776);
nand U2899 (N_2899,In_849,In_583);
xnor U2900 (N_2900,In_435,In_946);
xor U2901 (N_2901,In_898,In_833);
or U2902 (N_2902,In_301,In_324);
and U2903 (N_2903,In_20,In_595);
and U2904 (N_2904,In_615,In_20);
nor U2905 (N_2905,In_162,In_163);
nor U2906 (N_2906,In_184,In_287);
nor U2907 (N_2907,In_773,In_3);
nor U2908 (N_2908,In_794,In_984);
or U2909 (N_2909,In_397,In_309);
xnor U2910 (N_2910,In_192,In_805);
and U2911 (N_2911,In_474,In_200);
and U2912 (N_2912,In_663,In_247);
and U2913 (N_2913,In_730,In_785);
and U2914 (N_2914,In_967,In_162);
xor U2915 (N_2915,In_605,In_337);
and U2916 (N_2916,In_427,In_133);
xnor U2917 (N_2917,In_546,In_630);
or U2918 (N_2918,In_295,In_441);
xor U2919 (N_2919,In_64,In_141);
nand U2920 (N_2920,In_845,In_877);
or U2921 (N_2921,In_228,In_952);
nand U2922 (N_2922,In_71,In_488);
xor U2923 (N_2923,In_538,In_206);
nor U2924 (N_2924,In_170,In_627);
or U2925 (N_2925,In_202,In_779);
nand U2926 (N_2926,In_802,In_919);
or U2927 (N_2927,In_134,In_12);
or U2928 (N_2928,In_22,In_558);
or U2929 (N_2929,In_824,In_895);
and U2930 (N_2930,In_930,In_269);
nand U2931 (N_2931,In_456,In_290);
nor U2932 (N_2932,In_87,In_414);
nor U2933 (N_2933,In_354,In_481);
nand U2934 (N_2934,In_387,In_688);
nor U2935 (N_2935,In_653,In_206);
nor U2936 (N_2936,In_585,In_379);
nor U2937 (N_2937,In_87,In_684);
or U2938 (N_2938,In_342,In_354);
nor U2939 (N_2939,In_530,In_99);
xnor U2940 (N_2940,In_580,In_353);
xnor U2941 (N_2941,In_490,In_502);
or U2942 (N_2942,In_315,In_324);
or U2943 (N_2943,In_302,In_691);
or U2944 (N_2944,In_303,In_514);
nor U2945 (N_2945,In_98,In_49);
and U2946 (N_2946,In_113,In_865);
xnor U2947 (N_2947,In_985,In_529);
nor U2948 (N_2948,In_183,In_928);
and U2949 (N_2949,In_887,In_39);
and U2950 (N_2950,In_160,In_20);
and U2951 (N_2951,In_796,In_301);
or U2952 (N_2952,In_835,In_534);
xor U2953 (N_2953,In_654,In_363);
and U2954 (N_2954,In_17,In_108);
or U2955 (N_2955,In_479,In_85);
or U2956 (N_2956,In_258,In_752);
nor U2957 (N_2957,In_162,In_584);
or U2958 (N_2958,In_376,In_87);
xor U2959 (N_2959,In_601,In_302);
nor U2960 (N_2960,In_263,In_532);
xor U2961 (N_2961,In_303,In_682);
nor U2962 (N_2962,In_299,In_253);
xor U2963 (N_2963,In_865,In_413);
or U2964 (N_2964,In_670,In_746);
and U2965 (N_2965,In_993,In_310);
nor U2966 (N_2966,In_146,In_876);
nand U2967 (N_2967,In_434,In_223);
xnor U2968 (N_2968,In_559,In_480);
and U2969 (N_2969,In_235,In_461);
or U2970 (N_2970,In_309,In_196);
xnor U2971 (N_2971,In_268,In_639);
nor U2972 (N_2972,In_530,In_882);
nor U2973 (N_2973,In_477,In_821);
nand U2974 (N_2974,In_972,In_565);
and U2975 (N_2975,In_391,In_58);
or U2976 (N_2976,In_93,In_922);
xnor U2977 (N_2977,In_859,In_657);
and U2978 (N_2978,In_763,In_77);
and U2979 (N_2979,In_12,In_256);
or U2980 (N_2980,In_228,In_768);
and U2981 (N_2981,In_674,In_202);
or U2982 (N_2982,In_293,In_979);
and U2983 (N_2983,In_843,In_486);
nor U2984 (N_2984,In_515,In_528);
xnor U2985 (N_2985,In_58,In_733);
and U2986 (N_2986,In_456,In_510);
xnor U2987 (N_2987,In_422,In_782);
nand U2988 (N_2988,In_6,In_815);
xor U2989 (N_2989,In_381,In_427);
nor U2990 (N_2990,In_298,In_514);
and U2991 (N_2991,In_764,In_33);
nor U2992 (N_2992,In_750,In_770);
and U2993 (N_2993,In_842,In_27);
nor U2994 (N_2994,In_542,In_787);
nor U2995 (N_2995,In_492,In_184);
xor U2996 (N_2996,In_466,In_500);
xnor U2997 (N_2997,In_31,In_957);
nand U2998 (N_2998,In_72,In_532);
nor U2999 (N_2999,In_768,In_246);
xnor U3000 (N_3000,In_625,In_773);
nor U3001 (N_3001,In_104,In_940);
and U3002 (N_3002,In_267,In_381);
and U3003 (N_3003,In_412,In_825);
and U3004 (N_3004,In_812,In_636);
or U3005 (N_3005,In_870,In_702);
and U3006 (N_3006,In_74,In_184);
xnor U3007 (N_3007,In_784,In_832);
or U3008 (N_3008,In_711,In_553);
and U3009 (N_3009,In_615,In_955);
nand U3010 (N_3010,In_217,In_162);
nor U3011 (N_3011,In_421,In_216);
nor U3012 (N_3012,In_882,In_185);
nor U3013 (N_3013,In_672,In_899);
xnor U3014 (N_3014,In_401,In_650);
or U3015 (N_3015,In_723,In_879);
nand U3016 (N_3016,In_467,In_692);
nor U3017 (N_3017,In_58,In_783);
or U3018 (N_3018,In_707,In_51);
or U3019 (N_3019,In_228,In_559);
nand U3020 (N_3020,In_951,In_319);
or U3021 (N_3021,In_247,In_333);
or U3022 (N_3022,In_427,In_490);
and U3023 (N_3023,In_300,In_729);
nor U3024 (N_3024,In_826,In_205);
nor U3025 (N_3025,In_651,In_108);
or U3026 (N_3026,In_438,In_995);
and U3027 (N_3027,In_717,In_220);
or U3028 (N_3028,In_675,In_998);
xnor U3029 (N_3029,In_490,In_806);
and U3030 (N_3030,In_315,In_68);
nor U3031 (N_3031,In_787,In_733);
and U3032 (N_3032,In_862,In_462);
and U3033 (N_3033,In_595,In_187);
nor U3034 (N_3034,In_659,In_778);
xor U3035 (N_3035,In_424,In_404);
nand U3036 (N_3036,In_115,In_41);
nand U3037 (N_3037,In_31,In_15);
xnor U3038 (N_3038,In_821,In_744);
nor U3039 (N_3039,In_378,In_317);
nor U3040 (N_3040,In_68,In_196);
nand U3041 (N_3041,In_995,In_263);
xor U3042 (N_3042,In_871,In_617);
xnor U3043 (N_3043,In_142,In_485);
or U3044 (N_3044,In_90,In_486);
and U3045 (N_3045,In_136,In_402);
nor U3046 (N_3046,In_768,In_931);
or U3047 (N_3047,In_376,In_222);
or U3048 (N_3048,In_69,In_826);
xor U3049 (N_3049,In_362,In_134);
and U3050 (N_3050,In_156,In_288);
and U3051 (N_3051,In_333,In_474);
nor U3052 (N_3052,In_829,In_226);
xnor U3053 (N_3053,In_334,In_199);
nand U3054 (N_3054,In_645,In_248);
or U3055 (N_3055,In_53,In_730);
or U3056 (N_3056,In_131,In_647);
or U3057 (N_3057,In_479,In_511);
nand U3058 (N_3058,In_411,In_27);
or U3059 (N_3059,In_728,In_499);
or U3060 (N_3060,In_742,In_331);
and U3061 (N_3061,In_419,In_3);
and U3062 (N_3062,In_300,In_495);
or U3063 (N_3063,In_213,In_514);
nor U3064 (N_3064,In_268,In_463);
xnor U3065 (N_3065,In_401,In_702);
or U3066 (N_3066,In_47,In_732);
and U3067 (N_3067,In_406,In_648);
or U3068 (N_3068,In_236,In_246);
xor U3069 (N_3069,In_253,In_679);
nand U3070 (N_3070,In_102,In_245);
or U3071 (N_3071,In_745,In_732);
nor U3072 (N_3072,In_209,In_485);
nand U3073 (N_3073,In_587,In_347);
nand U3074 (N_3074,In_249,In_200);
nor U3075 (N_3075,In_519,In_274);
and U3076 (N_3076,In_572,In_366);
and U3077 (N_3077,In_488,In_110);
or U3078 (N_3078,In_164,In_615);
or U3079 (N_3079,In_61,In_358);
and U3080 (N_3080,In_38,In_793);
or U3081 (N_3081,In_748,In_184);
and U3082 (N_3082,In_11,In_54);
nor U3083 (N_3083,In_814,In_247);
and U3084 (N_3084,In_10,In_810);
and U3085 (N_3085,In_25,In_743);
and U3086 (N_3086,In_995,In_426);
nand U3087 (N_3087,In_356,In_651);
and U3088 (N_3088,In_645,In_287);
and U3089 (N_3089,In_51,In_200);
xor U3090 (N_3090,In_493,In_290);
or U3091 (N_3091,In_256,In_752);
or U3092 (N_3092,In_798,In_640);
and U3093 (N_3093,In_982,In_279);
or U3094 (N_3094,In_371,In_320);
xnor U3095 (N_3095,In_664,In_131);
xor U3096 (N_3096,In_320,In_558);
xor U3097 (N_3097,In_73,In_222);
nand U3098 (N_3098,In_682,In_65);
or U3099 (N_3099,In_836,In_905);
nor U3100 (N_3100,In_898,In_824);
xor U3101 (N_3101,In_918,In_633);
nor U3102 (N_3102,In_6,In_273);
nand U3103 (N_3103,In_833,In_390);
nand U3104 (N_3104,In_985,In_173);
and U3105 (N_3105,In_611,In_942);
xor U3106 (N_3106,In_470,In_711);
xnor U3107 (N_3107,In_974,In_323);
nand U3108 (N_3108,In_931,In_302);
nor U3109 (N_3109,In_438,In_675);
nand U3110 (N_3110,In_738,In_872);
and U3111 (N_3111,In_830,In_771);
or U3112 (N_3112,In_405,In_586);
and U3113 (N_3113,In_380,In_761);
xnor U3114 (N_3114,In_394,In_975);
nor U3115 (N_3115,In_795,In_796);
nand U3116 (N_3116,In_778,In_351);
and U3117 (N_3117,In_850,In_946);
xnor U3118 (N_3118,In_56,In_733);
nand U3119 (N_3119,In_396,In_486);
and U3120 (N_3120,In_973,In_831);
and U3121 (N_3121,In_426,In_460);
xnor U3122 (N_3122,In_448,In_759);
and U3123 (N_3123,In_777,In_470);
or U3124 (N_3124,In_317,In_45);
or U3125 (N_3125,In_99,In_881);
xnor U3126 (N_3126,In_409,In_967);
or U3127 (N_3127,In_304,In_435);
nand U3128 (N_3128,In_563,In_281);
nand U3129 (N_3129,In_585,In_453);
nand U3130 (N_3130,In_0,In_902);
nor U3131 (N_3131,In_599,In_974);
and U3132 (N_3132,In_280,In_694);
nor U3133 (N_3133,In_186,In_501);
and U3134 (N_3134,In_715,In_966);
and U3135 (N_3135,In_922,In_547);
nand U3136 (N_3136,In_224,In_688);
and U3137 (N_3137,In_471,In_409);
or U3138 (N_3138,In_447,In_429);
and U3139 (N_3139,In_753,In_141);
nand U3140 (N_3140,In_360,In_628);
or U3141 (N_3141,In_436,In_133);
nand U3142 (N_3142,In_394,In_169);
or U3143 (N_3143,In_775,In_148);
nor U3144 (N_3144,In_979,In_405);
and U3145 (N_3145,In_35,In_814);
xnor U3146 (N_3146,In_882,In_573);
xnor U3147 (N_3147,In_620,In_513);
or U3148 (N_3148,In_140,In_525);
and U3149 (N_3149,In_688,In_55);
nor U3150 (N_3150,In_430,In_450);
or U3151 (N_3151,In_656,In_779);
xnor U3152 (N_3152,In_200,In_380);
and U3153 (N_3153,In_876,In_164);
nor U3154 (N_3154,In_808,In_124);
xnor U3155 (N_3155,In_750,In_133);
nor U3156 (N_3156,In_311,In_216);
nand U3157 (N_3157,In_710,In_8);
nor U3158 (N_3158,In_698,In_924);
nor U3159 (N_3159,In_790,In_883);
nand U3160 (N_3160,In_396,In_441);
xnor U3161 (N_3161,In_732,In_233);
or U3162 (N_3162,In_148,In_165);
and U3163 (N_3163,In_752,In_393);
nor U3164 (N_3164,In_350,In_424);
nor U3165 (N_3165,In_429,In_629);
or U3166 (N_3166,In_578,In_613);
or U3167 (N_3167,In_872,In_890);
xor U3168 (N_3168,In_655,In_737);
or U3169 (N_3169,In_215,In_20);
nor U3170 (N_3170,In_930,In_54);
xnor U3171 (N_3171,In_319,In_709);
or U3172 (N_3172,In_293,In_917);
or U3173 (N_3173,In_213,In_1);
nand U3174 (N_3174,In_331,In_161);
nand U3175 (N_3175,In_138,In_635);
xor U3176 (N_3176,In_364,In_391);
or U3177 (N_3177,In_245,In_75);
nor U3178 (N_3178,In_674,In_769);
nor U3179 (N_3179,In_297,In_716);
or U3180 (N_3180,In_851,In_983);
nor U3181 (N_3181,In_13,In_257);
xnor U3182 (N_3182,In_225,In_304);
and U3183 (N_3183,In_444,In_664);
nand U3184 (N_3184,In_620,In_810);
and U3185 (N_3185,In_329,In_920);
and U3186 (N_3186,In_911,In_190);
and U3187 (N_3187,In_958,In_276);
or U3188 (N_3188,In_583,In_422);
and U3189 (N_3189,In_430,In_199);
nor U3190 (N_3190,In_370,In_407);
nand U3191 (N_3191,In_888,In_965);
or U3192 (N_3192,In_38,In_664);
and U3193 (N_3193,In_782,In_335);
nand U3194 (N_3194,In_327,In_520);
nand U3195 (N_3195,In_780,In_415);
nand U3196 (N_3196,In_786,In_672);
nor U3197 (N_3197,In_828,In_644);
xnor U3198 (N_3198,In_482,In_103);
and U3199 (N_3199,In_94,In_863);
xnor U3200 (N_3200,In_145,In_126);
xnor U3201 (N_3201,In_751,In_763);
or U3202 (N_3202,In_236,In_61);
and U3203 (N_3203,In_129,In_116);
or U3204 (N_3204,In_48,In_140);
nand U3205 (N_3205,In_544,In_714);
xor U3206 (N_3206,In_850,In_357);
xnor U3207 (N_3207,In_916,In_104);
nand U3208 (N_3208,In_350,In_492);
or U3209 (N_3209,In_40,In_243);
or U3210 (N_3210,In_673,In_883);
xor U3211 (N_3211,In_794,In_523);
nand U3212 (N_3212,In_392,In_630);
or U3213 (N_3213,In_636,In_923);
nand U3214 (N_3214,In_124,In_252);
and U3215 (N_3215,In_518,In_196);
or U3216 (N_3216,In_419,In_445);
xnor U3217 (N_3217,In_518,In_249);
or U3218 (N_3218,In_797,In_504);
nor U3219 (N_3219,In_757,In_133);
xor U3220 (N_3220,In_345,In_312);
or U3221 (N_3221,In_346,In_864);
nand U3222 (N_3222,In_857,In_615);
and U3223 (N_3223,In_715,In_285);
nand U3224 (N_3224,In_803,In_799);
nor U3225 (N_3225,In_372,In_697);
and U3226 (N_3226,In_918,In_53);
or U3227 (N_3227,In_678,In_656);
xnor U3228 (N_3228,In_581,In_105);
or U3229 (N_3229,In_298,In_93);
xor U3230 (N_3230,In_421,In_285);
xnor U3231 (N_3231,In_840,In_249);
nand U3232 (N_3232,In_132,In_105);
nor U3233 (N_3233,In_48,In_68);
nand U3234 (N_3234,In_896,In_807);
nand U3235 (N_3235,In_598,In_452);
and U3236 (N_3236,In_235,In_714);
nor U3237 (N_3237,In_424,In_691);
or U3238 (N_3238,In_141,In_507);
xor U3239 (N_3239,In_844,In_439);
nand U3240 (N_3240,In_174,In_875);
nand U3241 (N_3241,In_365,In_142);
and U3242 (N_3242,In_817,In_748);
nor U3243 (N_3243,In_684,In_62);
nand U3244 (N_3244,In_100,In_373);
nor U3245 (N_3245,In_312,In_168);
nor U3246 (N_3246,In_71,In_651);
xor U3247 (N_3247,In_692,In_90);
nor U3248 (N_3248,In_497,In_16);
nor U3249 (N_3249,In_772,In_138);
or U3250 (N_3250,In_986,In_646);
xnor U3251 (N_3251,In_238,In_377);
and U3252 (N_3252,In_752,In_99);
nor U3253 (N_3253,In_72,In_443);
nor U3254 (N_3254,In_354,In_169);
nand U3255 (N_3255,In_781,In_163);
nand U3256 (N_3256,In_428,In_623);
xnor U3257 (N_3257,In_170,In_727);
nand U3258 (N_3258,In_681,In_61);
nand U3259 (N_3259,In_922,In_134);
and U3260 (N_3260,In_786,In_471);
nor U3261 (N_3261,In_308,In_698);
and U3262 (N_3262,In_798,In_534);
nand U3263 (N_3263,In_442,In_663);
or U3264 (N_3264,In_535,In_951);
xor U3265 (N_3265,In_883,In_975);
xor U3266 (N_3266,In_238,In_973);
or U3267 (N_3267,In_585,In_637);
xor U3268 (N_3268,In_115,In_909);
or U3269 (N_3269,In_633,In_21);
and U3270 (N_3270,In_779,In_628);
nor U3271 (N_3271,In_227,In_140);
or U3272 (N_3272,In_800,In_771);
nand U3273 (N_3273,In_456,In_101);
and U3274 (N_3274,In_781,In_605);
nor U3275 (N_3275,In_118,In_794);
or U3276 (N_3276,In_879,In_331);
nand U3277 (N_3277,In_250,In_770);
nand U3278 (N_3278,In_112,In_576);
or U3279 (N_3279,In_655,In_753);
or U3280 (N_3280,In_577,In_846);
and U3281 (N_3281,In_359,In_59);
or U3282 (N_3282,In_234,In_959);
xnor U3283 (N_3283,In_592,In_375);
nor U3284 (N_3284,In_418,In_164);
nand U3285 (N_3285,In_338,In_842);
nand U3286 (N_3286,In_990,In_973);
or U3287 (N_3287,In_689,In_948);
xor U3288 (N_3288,In_391,In_990);
xor U3289 (N_3289,In_55,In_200);
and U3290 (N_3290,In_795,In_778);
or U3291 (N_3291,In_148,In_399);
or U3292 (N_3292,In_168,In_631);
or U3293 (N_3293,In_408,In_113);
and U3294 (N_3294,In_323,In_76);
nor U3295 (N_3295,In_931,In_766);
nand U3296 (N_3296,In_261,In_403);
and U3297 (N_3297,In_644,In_799);
xor U3298 (N_3298,In_467,In_810);
nand U3299 (N_3299,In_270,In_466);
nor U3300 (N_3300,In_214,In_713);
nor U3301 (N_3301,In_820,In_595);
xor U3302 (N_3302,In_672,In_395);
nand U3303 (N_3303,In_575,In_430);
and U3304 (N_3304,In_627,In_126);
nor U3305 (N_3305,In_931,In_33);
xnor U3306 (N_3306,In_73,In_503);
nor U3307 (N_3307,In_457,In_72);
nor U3308 (N_3308,In_420,In_927);
or U3309 (N_3309,In_252,In_96);
and U3310 (N_3310,In_197,In_459);
or U3311 (N_3311,In_557,In_20);
and U3312 (N_3312,In_211,In_907);
nor U3313 (N_3313,In_847,In_377);
nor U3314 (N_3314,In_116,In_637);
and U3315 (N_3315,In_649,In_840);
and U3316 (N_3316,In_600,In_994);
nor U3317 (N_3317,In_517,In_631);
or U3318 (N_3318,In_285,In_260);
and U3319 (N_3319,In_239,In_7);
nor U3320 (N_3320,In_895,In_17);
or U3321 (N_3321,In_850,In_637);
nor U3322 (N_3322,In_704,In_961);
xnor U3323 (N_3323,In_372,In_596);
nor U3324 (N_3324,In_764,In_722);
nor U3325 (N_3325,In_378,In_633);
nor U3326 (N_3326,In_639,In_408);
or U3327 (N_3327,In_178,In_49);
xor U3328 (N_3328,In_554,In_197);
xor U3329 (N_3329,In_56,In_822);
nor U3330 (N_3330,In_406,In_94);
nor U3331 (N_3331,In_161,In_696);
or U3332 (N_3332,In_653,In_975);
and U3333 (N_3333,In_905,In_392);
xnor U3334 (N_3334,In_891,In_950);
and U3335 (N_3335,In_819,In_361);
and U3336 (N_3336,In_332,In_387);
and U3337 (N_3337,In_999,In_976);
xor U3338 (N_3338,In_145,In_162);
and U3339 (N_3339,In_36,In_104);
xor U3340 (N_3340,In_849,In_787);
xor U3341 (N_3341,In_534,In_215);
nand U3342 (N_3342,In_61,In_897);
xnor U3343 (N_3343,In_204,In_52);
or U3344 (N_3344,In_33,In_515);
xor U3345 (N_3345,In_945,In_304);
and U3346 (N_3346,In_772,In_444);
and U3347 (N_3347,In_202,In_401);
and U3348 (N_3348,In_351,In_934);
and U3349 (N_3349,In_943,In_869);
xnor U3350 (N_3350,In_101,In_363);
and U3351 (N_3351,In_845,In_206);
nand U3352 (N_3352,In_57,In_257);
nor U3353 (N_3353,In_458,In_481);
nand U3354 (N_3354,In_111,In_70);
xnor U3355 (N_3355,In_81,In_855);
or U3356 (N_3356,In_815,In_191);
nor U3357 (N_3357,In_184,In_24);
or U3358 (N_3358,In_900,In_298);
nor U3359 (N_3359,In_860,In_292);
and U3360 (N_3360,In_824,In_137);
xnor U3361 (N_3361,In_432,In_972);
or U3362 (N_3362,In_463,In_159);
or U3363 (N_3363,In_34,In_461);
xnor U3364 (N_3364,In_44,In_487);
or U3365 (N_3365,In_220,In_668);
and U3366 (N_3366,In_512,In_598);
nand U3367 (N_3367,In_145,In_514);
xor U3368 (N_3368,In_806,In_233);
and U3369 (N_3369,In_675,In_40);
and U3370 (N_3370,In_538,In_391);
xor U3371 (N_3371,In_731,In_721);
and U3372 (N_3372,In_141,In_208);
nor U3373 (N_3373,In_721,In_40);
nor U3374 (N_3374,In_357,In_101);
nor U3375 (N_3375,In_564,In_543);
or U3376 (N_3376,In_437,In_877);
or U3377 (N_3377,In_19,In_169);
xnor U3378 (N_3378,In_650,In_695);
or U3379 (N_3379,In_289,In_659);
or U3380 (N_3380,In_485,In_930);
xor U3381 (N_3381,In_903,In_245);
xor U3382 (N_3382,In_42,In_460);
xor U3383 (N_3383,In_160,In_24);
xnor U3384 (N_3384,In_76,In_361);
nand U3385 (N_3385,In_93,In_185);
xor U3386 (N_3386,In_717,In_304);
nand U3387 (N_3387,In_261,In_382);
nand U3388 (N_3388,In_548,In_615);
xnor U3389 (N_3389,In_660,In_298);
xor U3390 (N_3390,In_750,In_696);
nand U3391 (N_3391,In_737,In_902);
and U3392 (N_3392,In_441,In_825);
nand U3393 (N_3393,In_254,In_983);
nand U3394 (N_3394,In_754,In_766);
and U3395 (N_3395,In_780,In_860);
xor U3396 (N_3396,In_229,In_489);
nand U3397 (N_3397,In_470,In_213);
nor U3398 (N_3398,In_554,In_918);
or U3399 (N_3399,In_384,In_895);
or U3400 (N_3400,In_458,In_480);
xor U3401 (N_3401,In_195,In_309);
xor U3402 (N_3402,In_461,In_535);
or U3403 (N_3403,In_690,In_279);
xor U3404 (N_3404,In_279,In_684);
or U3405 (N_3405,In_716,In_990);
nand U3406 (N_3406,In_22,In_511);
nand U3407 (N_3407,In_312,In_812);
nand U3408 (N_3408,In_377,In_721);
nand U3409 (N_3409,In_133,In_262);
nor U3410 (N_3410,In_456,In_654);
nand U3411 (N_3411,In_990,In_610);
and U3412 (N_3412,In_22,In_274);
nor U3413 (N_3413,In_746,In_161);
or U3414 (N_3414,In_739,In_963);
and U3415 (N_3415,In_312,In_509);
nor U3416 (N_3416,In_404,In_361);
nor U3417 (N_3417,In_826,In_869);
and U3418 (N_3418,In_348,In_179);
and U3419 (N_3419,In_905,In_929);
and U3420 (N_3420,In_255,In_353);
or U3421 (N_3421,In_569,In_439);
and U3422 (N_3422,In_584,In_413);
and U3423 (N_3423,In_540,In_673);
or U3424 (N_3424,In_196,In_915);
nor U3425 (N_3425,In_736,In_486);
nand U3426 (N_3426,In_641,In_178);
nor U3427 (N_3427,In_451,In_108);
nor U3428 (N_3428,In_874,In_718);
or U3429 (N_3429,In_553,In_96);
nor U3430 (N_3430,In_665,In_631);
xnor U3431 (N_3431,In_681,In_904);
xor U3432 (N_3432,In_319,In_624);
xnor U3433 (N_3433,In_711,In_679);
or U3434 (N_3434,In_739,In_439);
or U3435 (N_3435,In_434,In_984);
nor U3436 (N_3436,In_748,In_785);
xor U3437 (N_3437,In_505,In_79);
and U3438 (N_3438,In_424,In_63);
and U3439 (N_3439,In_260,In_529);
nand U3440 (N_3440,In_508,In_890);
or U3441 (N_3441,In_243,In_875);
nor U3442 (N_3442,In_411,In_899);
xor U3443 (N_3443,In_136,In_823);
nand U3444 (N_3444,In_157,In_448);
and U3445 (N_3445,In_239,In_968);
xnor U3446 (N_3446,In_144,In_117);
nor U3447 (N_3447,In_52,In_758);
and U3448 (N_3448,In_307,In_505);
nor U3449 (N_3449,In_823,In_140);
xor U3450 (N_3450,In_451,In_20);
nor U3451 (N_3451,In_624,In_467);
or U3452 (N_3452,In_659,In_934);
nand U3453 (N_3453,In_705,In_687);
and U3454 (N_3454,In_664,In_152);
nand U3455 (N_3455,In_150,In_320);
xnor U3456 (N_3456,In_93,In_942);
and U3457 (N_3457,In_626,In_247);
xnor U3458 (N_3458,In_525,In_469);
nor U3459 (N_3459,In_775,In_474);
xnor U3460 (N_3460,In_557,In_408);
and U3461 (N_3461,In_442,In_382);
xnor U3462 (N_3462,In_645,In_922);
or U3463 (N_3463,In_143,In_73);
nand U3464 (N_3464,In_388,In_403);
or U3465 (N_3465,In_734,In_603);
nand U3466 (N_3466,In_574,In_52);
or U3467 (N_3467,In_920,In_450);
nor U3468 (N_3468,In_787,In_945);
nor U3469 (N_3469,In_683,In_576);
and U3470 (N_3470,In_709,In_589);
nor U3471 (N_3471,In_60,In_659);
or U3472 (N_3472,In_446,In_131);
nor U3473 (N_3473,In_47,In_255);
nor U3474 (N_3474,In_151,In_497);
and U3475 (N_3475,In_985,In_536);
and U3476 (N_3476,In_244,In_816);
and U3477 (N_3477,In_18,In_571);
and U3478 (N_3478,In_26,In_843);
xor U3479 (N_3479,In_359,In_501);
and U3480 (N_3480,In_577,In_942);
nor U3481 (N_3481,In_133,In_138);
nand U3482 (N_3482,In_45,In_673);
and U3483 (N_3483,In_31,In_217);
nor U3484 (N_3484,In_330,In_45);
nand U3485 (N_3485,In_470,In_257);
nor U3486 (N_3486,In_427,In_107);
xor U3487 (N_3487,In_297,In_270);
and U3488 (N_3488,In_282,In_229);
xor U3489 (N_3489,In_628,In_69);
nor U3490 (N_3490,In_146,In_134);
or U3491 (N_3491,In_353,In_851);
nand U3492 (N_3492,In_47,In_382);
nor U3493 (N_3493,In_815,In_877);
nor U3494 (N_3494,In_245,In_977);
xnor U3495 (N_3495,In_698,In_441);
xor U3496 (N_3496,In_700,In_94);
xnor U3497 (N_3497,In_922,In_786);
and U3498 (N_3498,In_805,In_19);
and U3499 (N_3499,In_456,In_776);
or U3500 (N_3500,In_119,In_49);
nand U3501 (N_3501,In_42,In_206);
or U3502 (N_3502,In_877,In_940);
or U3503 (N_3503,In_387,In_666);
and U3504 (N_3504,In_248,In_823);
xor U3505 (N_3505,In_768,In_321);
nor U3506 (N_3506,In_23,In_252);
xor U3507 (N_3507,In_720,In_388);
or U3508 (N_3508,In_662,In_589);
nand U3509 (N_3509,In_837,In_221);
and U3510 (N_3510,In_236,In_78);
and U3511 (N_3511,In_660,In_519);
or U3512 (N_3512,In_197,In_427);
nor U3513 (N_3513,In_442,In_941);
and U3514 (N_3514,In_261,In_760);
nand U3515 (N_3515,In_569,In_979);
and U3516 (N_3516,In_188,In_476);
xnor U3517 (N_3517,In_681,In_586);
xor U3518 (N_3518,In_524,In_446);
or U3519 (N_3519,In_941,In_185);
and U3520 (N_3520,In_337,In_454);
xor U3521 (N_3521,In_701,In_281);
xnor U3522 (N_3522,In_901,In_60);
xnor U3523 (N_3523,In_337,In_802);
xor U3524 (N_3524,In_641,In_916);
nand U3525 (N_3525,In_196,In_512);
xnor U3526 (N_3526,In_374,In_441);
nand U3527 (N_3527,In_508,In_449);
nand U3528 (N_3528,In_587,In_320);
xor U3529 (N_3529,In_80,In_484);
nor U3530 (N_3530,In_471,In_682);
nand U3531 (N_3531,In_790,In_958);
nor U3532 (N_3532,In_400,In_494);
xnor U3533 (N_3533,In_860,In_25);
xnor U3534 (N_3534,In_389,In_817);
and U3535 (N_3535,In_172,In_906);
xor U3536 (N_3536,In_102,In_220);
or U3537 (N_3537,In_834,In_729);
nand U3538 (N_3538,In_30,In_312);
xor U3539 (N_3539,In_526,In_199);
and U3540 (N_3540,In_369,In_397);
nand U3541 (N_3541,In_894,In_470);
xor U3542 (N_3542,In_798,In_997);
and U3543 (N_3543,In_149,In_182);
and U3544 (N_3544,In_281,In_420);
nand U3545 (N_3545,In_689,In_584);
or U3546 (N_3546,In_273,In_53);
xor U3547 (N_3547,In_3,In_225);
and U3548 (N_3548,In_958,In_107);
xor U3549 (N_3549,In_886,In_324);
and U3550 (N_3550,In_139,In_444);
or U3551 (N_3551,In_755,In_996);
nor U3552 (N_3552,In_959,In_219);
or U3553 (N_3553,In_143,In_767);
nand U3554 (N_3554,In_408,In_468);
or U3555 (N_3555,In_364,In_989);
and U3556 (N_3556,In_626,In_675);
and U3557 (N_3557,In_98,In_313);
nand U3558 (N_3558,In_249,In_643);
nor U3559 (N_3559,In_926,In_958);
nor U3560 (N_3560,In_802,In_593);
and U3561 (N_3561,In_132,In_729);
or U3562 (N_3562,In_616,In_587);
or U3563 (N_3563,In_767,In_954);
nand U3564 (N_3564,In_820,In_887);
or U3565 (N_3565,In_195,In_207);
nand U3566 (N_3566,In_161,In_993);
or U3567 (N_3567,In_319,In_753);
nand U3568 (N_3568,In_248,In_113);
nand U3569 (N_3569,In_765,In_908);
and U3570 (N_3570,In_115,In_707);
or U3571 (N_3571,In_151,In_398);
nand U3572 (N_3572,In_35,In_330);
nand U3573 (N_3573,In_793,In_565);
nor U3574 (N_3574,In_908,In_430);
nand U3575 (N_3575,In_341,In_521);
nor U3576 (N_3576,In_455,In_90);
or U3577 (N_3577,In_897,In_889);
nor U3578 (N_3578,In_573,In_348);
nand U3579 (N_3579,In_602,In_118);
nand U3580 (N_3580,In_957,In_618);
xor U3581 (N_3581,In_8,In_744);
xor U3582 (N_3582,In_793,In_210);
and U3583 (N_3583,In_628,In_791);
or U3584 (N_3584,In_749,In_35);
or U3585 (N_3585,In_664,In_495);
nor U3586 (N_3586,In_474,In_589);
or U3587 (N_3587,In_380,In_614);
nand U3588 (N_3588,In_980,In_100);
or U3589 (N_3589,In_663,In_804);
nand U3590 (N_3590,In_632,In_103);
nor U3591 (N_3591,In_179,In_962);
xnor U3592 (N_3592,In_105,In_217);
xor U3593 (N_3593,In_358,In_159);
nand U3594 (N_3594,In_479,In_340);
xor U3595 (N_3595,In_486,In_735);
nand U3596 (N_3596,In_606,In_127);
nand U3597 (N_3597,In_506,In_686);
nor U3598 (N_3598,In_409,In_843);
nand U3599 (N_3599,In_653,In_388);
xor U3600 (N_3600,In_593,In_71);
and U3601 (N_3601,In_720,In_840);
xnor U3602 (N_3602,In_280,In_450);
or U3603 (N_3603,In_465,In_948);
and U3604 (N_3604,In_32,In_915);
or U3605 (N_3605,In_754,In_249);
xor U3606 (N_3606,In_397,In_894);
nor U3607 (N_3607,In_313,In_101);
and U3608 (N_3608,In_740,In_486);
or U3609 (N_3609,In_11,In_98);
and U3610 (N_3610,In_53,In_900);
or U3611 (N_3611,In_967,In_857);
or U3612 (N_3612,In_53,In_815);
or U3613 (N_3613,In_317,In_770);
nor U3614 (N_3614,In_493,In_260);
and U3615 (N_3615,In_17,In_919);
and U3616 (N_3616,In_987,In_90);
xnor U3617 (N_3617,In_959,In_815);
nand U3618 (N_3618,In_166,In_475);
nand U3619 (N_3619,In_195,In_869);
and U3620 (N_3620,In_94,In_398);
nor U3621 (N_3621,In_177,In_485);
and U3622 (N_3622,In_310,In_432);
and U3623 (N_3623,In_404,In_463);
nor U3624 (N_3624,In_499,In_544);
or U3625 (N_3625,In_717,In_567);
xor U3626 (N_3626,In_706,In_806);
nor U3627 (N_3627,In_104,In_400);
or U3628 (N_3628,In_47,In_806);
xor U3629 (N_3629,In_966,In_70);
nor U3630 (N_3630,In_52,In_98);
and U3631 (N_3631,In_883,In_623);
nor U3632 (N_3632,In_461,In_242);
nand U3633 (N_3633,In_526,In_914);
and U3634 (N_3634,In_128,In_817);
nand U3635 (N_3635,In_988,In_661);
or U3636 (N_3636,In_157,In_129);
or U3637 (N_3637,In_853,In_322);
xnor U3638 (N_3638,In_674,In_511);
or U3639 (N_3639,In_945,In_717);
nand U3640 (N_3640,In_29,In_561);
nor U3641 (N_3641,In_586,In_278);
nor U3642 (N_3642,In_179,In_130);
or U3643 (N_3643,In_8,In_372);
nor U3644 (N_3644,In_288,In_884);
nor U3645 (N_3645,In_324,In_261);
and U3646 (N_3646,In_12,In_363);
nor U3647 (N_3647,In_284,In_96);
or U3648 (N_3648,In_557,In_134);
or U3649 (N_3649,In_790,In_236);
nor U3650 (N_3650,In_739,In_409);
nor U3651 (N_3651,In_940,In_29);
or U3652 (N_3652,In_85,In_292);
nor U3653 (N_3653,In_788,In_969);
nand U3654 (N_3654,In_477,In_120);
or U3655 (N_3655,In_102,In_327);
nor U3656 (N_3656,In_177,In_410);
xnor U3657 (N_3657,In_97,In_201);
and U3658 (N_3658,In_339,In_584);
nor U3659 (N_3659,In_629,In_356);
nor U3660 (N_3660,In_341,In_262);
nor U3661 (N_3661,In_130,In_412);
nand U3662 (N_3662,In_528,In_895);
and U3663 (N_3663,In_330,In_788);
nand U3664 (N_3664,In_743,In_742);
and U3665 (N_3665,In_84,In_328);
nor U3666 (N_3666,In_652,In_144);
or U3667 (N_3667,In_814,In_6);
and U3668 (N_3668,In_754,In_334);
and U3669 (N_3669,In_145,In_747);
and U3670 (N_3670,In_820,In_218);
xnor U3671 (N_3671,In_667,In_879);
and U3672 (N_3672,In_934,In_240);
nand U3673 (N_3673,In_378,In_324);
nand U3674 (N_3674,In_232,In_623);
or U3675 (N_3675,In_899,In_840);
nor U3676 (N_3676,In_288,In_358);
nor U3677 (N_3677,In_128,In_907);
and U3678 (N_3678,In_10,In_646);
xor U3679 (N_3679,In_853,In_426);
and U3680 (N_3680,In_618,In_641);
xor U3681 (N_3681,In_791,In_906);
and U3682 (N_3682,In_310,In_338);
or U3683 (N_3683,In_957,In_736);
and U3684 (N_3684,In_605,In_297);
nor U3685 (N_3685,In_900,In_817);
nor U3686 (N_3686,In_948,In_991);
or U3687 (N_3687,In_387,In_493);
and U3688 (N_3688,In_64,In_702);
or U3689 (N_3689,In_906,In_263);
or U3690 (N_3690,In_747,In_31);
nor U3691 (N_3691,In_617,In_238);
nand U3692 (N_3692,In_655,In_517);
and U3693 (N_3693,In_104,In_650);
nor U3694 (N_3694,In_677,In_184);
or U3695 (N_3695,In_286,In_291);
or U3696 (N_3696,In_364,In_164);
nor U3697 (N_3697,In_573,In_655);
nor U3698 (N_3698,In_576,In_348);
nand U3699 (N_3699,In_136,In_565);
nor U3700 (N_3700,In_472,In_75);
nand U3701 (N_3701,In_665,In_554);
nand U3702 (N_3702,In_722,In_359);
nand U3703 (N_3703,In_765,In_54);
and U3704 (N_3704,In_643,In_163);
or U3705 (N_3705,In_255,In_772);
and U3706 (N_3706,In_226,In_52);
nand U3707 (N_3707,In_98,In_863);
or U3708 (N_3708,In_556,In_277);
xnor U3709 (N_3709,In_16,In_121);
xor U3710 (N_3710,In_745,In_350);
and U3711 (N_3711,In_146,In_517);
and U3712 (N_3712,In_559,In_865);
and U3713 (N_3713,In_34,In_248);
nor U3714 (N_3714,In_985,In_240);
and U3715 (N_3715,In_904,In_888);
xor U3716 (N_3716,In_951,In_23);
and U3717 (N_3717,In_978,In_557);
and U3718 (N_3718,In_742,In_66);
xnor U3719 (N_3719,In_160,In_23);
nand U3720 (N_3720,In_393,In_217);
nand U3721 (N_3721,In_370,In_213);
or U3722 (N_3722,In_78,In_688);
nand U3723 (N_3723,In_745,In_860);
and U3724 (N_3724,In_358,In_57);
nor U3725 (N_3725,In_174,In_243);
nand U3726 (N_3726,In_438,In_554);
xor U3727 (N_3727,In_241,In_521);
nor U3728 (N_3728,In_552,In_67);
xnor U3729 (N_3729,In_253,In_182);
xnor U3730 (N_3730,In_906,In_541);
or U3731 (N_3731,In_952,In_662);
or U3732 (N_3732,In_356,In_731);
and U3733 (N_3733,In_159,In_199);
nor U3734 (N_3734,In_573,In_835);
or U3735 (N_3735,In_739,In_490);
or U3736 (N_3736,In_926,In_207);
nand U3737 (N_3737,In_352,In_445);
nand U3738 (N_3738,In_813,In_652);
or U3739 (N_3739,In_105,In_162);
nor U3740 (N_3740,In_682,In_630);
xor U3741 (N_3741,In_137,In_180);
or U3742 (N_3742,In_109,In_207);
nor U3743 (N_3743,In_744,In_954);
or U3744 (N_3744,In_433,In_753);
nand U3745 (N_3745,In_991,In_787);
and U3746 (N_3746,In_708,In_489);
xor U3747 (N_3747,In_127,In_965);
and U3748 (N_3748,In_991,In_397);
or U3749 (N_3749,In_910,In_641);
or U3750 (N_3750,In_221,In_178);
nor U3751 (N_3751,In_670,In_503);
nor U3752 (N_3752,In_868,In_27);
or U3753 (N_3753,In_969,In_978);
or U3754 (N_3754,In_822,In_789);
nand U3755 (N_3755,In_682,In_35);
and U3756 (N_3756,In_957,In_634);
nand U3757 (N_3757,In_415,In_868);
xnor U3758 (N_3758,In_481,In_35);
nand U3759 (N_3759,In_180,In_818);
or U3760 (N_3760,In_512,In_306);
and U3761 (N_3761,In_892,In_262);
xor U3762 (N_3762,In_548,In_998);
or U3763 (N_3763,In_810,In_341);
or U3764 (N_3764,In_434,In_445);
nand U3765 (N_3765,In_803,In_665);
and U3766 (N_3766,In_335,In_981);
or U3767 (N_3767,In_241,In_722);
nor U3768 (N_3768,In_98,In_853);
and U3769 (N_3769,In_597,In_467);
nand U3770 (N_3770,In_871,In_650);
nor U3771 (N_3771,In_416,In_891);
and U3772 (N_3772,In_162,In_33);
nand U3773 (N_3773,In_75,In_666);
or U3774 (N_3774,In_716,In_229);
xor U3775 (N_3775,In_86,In_113);
nand U3776 (N_3776,In_696,In_950);
xnor U3777 (N_3777,In_635,In_375);
nand U3778 (N_3778,In_807,In_941);
nor U3779 (N_3779,In_257,In_720);
nor U3780 (N_3780,In_77,In_840);
and U3781 (N_3781,In_61,In_471);
xnor U3782 (N_3782,In_781,In_751);
nor U3783 (N_3783,In_583,In_203);
and U3784 (N_3784,In_458,In_862);
nand U3785 (N_3785,In_431,In_583);
and U3786 (N_3786,In_88,In_399);
nor U3787 (N_3787,In_69,In_458);
or U3788 (N_3788,In_923,In_191);
nand U3789 (N_3789,In_305,In_549);
nand U3790 (N_3790,In_769,In_249);
nor U3791 (N_3791,In_667,In_833);
nand U3792 (N_3792,In_678,In_881);
nand U3793 (N_3793,In_851,In_563);
nor U3794 (N_3794,In_59,In_430);
nand U3795 (N_3795,In_133,In_561);
nand U3796 (N_3796,In_259,In_661);
or U3797 (N_3797,In_931,In_233);
and U3798 (N_3798,In_248,In_935);
or U3799 (N_3799,In_806,In_216);
nor U3800 (N_3800,In_674,In_967);
nor U3801 (N_3801,In_257,In_843);
nor U3802 (N_3802,In_101,In_535);
and U3803 (N_3803,In_924,In_482);
and U3804 (N_3804,In_380,In_977);
xnor U3805 (N_3805,In_516,In_843);
and U3806 (N_3806,In_933,In_230);
nor U3807 (N_3807,In_802,In_755);
nor U3808 (N_3808,In_354,In_299);
and U3809 (N_3809,In_624,In_756);
and U3810 (N_3810,In_549,In_297);
nand U3811 (N_3811,In_840,In_169);
nand U3812 (N_3812,In_100,In_164);
and U3813 (N_3813,In_168,In_824);
nand U3814 (N_3814,In_68,In_807);
and U3815 (N_3815,In_269,In_791);
or U3816 (N_3816,In_41,In_150);
xor U3817 (N_3817,In_582,In_675);
nor U3818 (N_3818,In_777,In_274);
xor U3819 (N_3819,In_255,In_19);
xnor U3820 (N_3820,In_46,In_787);
or U3821 (N_3821,In_362,In_785);
nand U3822 (N_3822,In_150,In_508);
xor U3823 (N_3823,In_409,In_586);
nor U3824 (N_3824,In_475,In_872);
or U3825 (N_3825,In_496,In_88);
nand U3826 (N_3826,In_88,In_624);
or U3827 (N_3827,In_579,In_228);
xnor U3828 (N_3828,In_748,In_720);
xor U3829 (N_3829,In_849,In_609);
nand U3830 (N_3830,In_31,In_865);
or U3831 (N_3831,In_616,In_30);
nor U3832 (N_3832,In_469,In_611);
nand U3833 (N_3833,In_235,In_335);
xnor U3834 (N_3834,In_598,In_190);
xnor U3835 (N_3835,In_288,In_866);
and U3836 (N_3836,In_5,In_318);
nor U3837 (N_3837,In_860,In_947);
nand U3838 (N_3838,In_388,In_193);
or U3839 (N_3839,In_690,In_800);
xnor U3840 (N_3840,In_914,In_843);
nand U3841 (N_3841,In_893,In_278);
or U3842 (N_3842,In_202,In_448);
nor U3843 (N_3843,In_299,In_363);
xnor U3844 (N_3844,In_204,In_736);
nor U3845 (N_3845,In_549,In_492);
or U3846 (N_3846,In_402,In_198);
nand U3847 (N_3847,In_461,In_136);
xor U3848 (N_3848,In_107,In_918);
and U3849 (N_3849,In_487,In_324);
and U3850 (N_3850,In_815,In_680);
nor U3851 (N_3851,In_163,In_165);
or U3852 (N_3852,In_54,In_208);
nor U3853 (N_3853,In_914,In_947);
xor U3854 (N_3854,In_348,In_819);
and U3855 (N_3855,In_837,In_766);
xnor U3856 (N_3856,In_677,In_715);
nand U3857 (N_3857,In_405,In_693);
nor U3858 (N_3858,In_351,In_142);
xnor U3859 (N_3859,In_29,In_374);
xnor U3860 (N_3860,In_858,In_834);
and U3861 (N_3861,In_600,In_920);
or U3862 (N_3862,In_486,In_3);
nor U3863 (N_3863,In_77,In_986);
nor U3864 (N_3864,In_25,In_752);
nand U3865 (N_3865,In_40,In_561);
or U3866 (N_3866,In_621,In_782);
nor U3867 (N_3867,In_741,In_824);
or U3868 (N_3868,In_463,In_822);
nand U3869 (N_3869,In_920,In_708);
or U3870 (N_3870,In_766,In_783);
or U3871 (N_3871,In_734,In_137);
xor U3872 (N_3872,In_402,In_834);
nand U3873 (N_3873,In_712,In_591);
xnor U3874 (N_3874,In_495,In_510);
nand U3875 (N_3875,In_674,In_228);
nand U3876 (N_3876,In_400,In_345);
or U3877 (N_3877,In_390,In_439);
and U3878 (N_3878,In_287,In_371);
and U3879 (N_3879,In_879,In_499);
or U3880 (N_3880,In_445,In_969);
xnor U3881 (N_3881,In_533,In_537);
nor U3882 (N_3882,In_236,In_113);
nor U3883 (N_3883,In_741,In_918);
nor U3884 (N_3884,In_500,In_402);
nand U3885 (N_3885,In_803,In_69);
nor U3886 (N_3886,In_352,In_50);
nand U3887 (N_3887,In_437,In_248);
xnor U3888 (N_3888,In_36,In_268);
or U3889 (N_3889,In_103,In_175);
and U3890 (N_3890,In_718,In_441);
nand U3891 (N_3891,In_621,In_225);
or U3892 (N_3892,In_495,In_888);
or U3893 (N_3893,In_680,In_275);
or U3894 (N_3894,In_937,In_949);
nand U3895 (N_3895,In_351,In_960);
or U3896 (N_3896,In_878,In_130);
and U3897 (N_3897,In_757,In_104);
and U3898 (N_3898,In_881,In_71);
nor U3899 (N_3899,In_981,In_801);
xor U3900 (N_3900,In_745,In_119);
and U3901 (N_3901,In_75,In_977);
nor U3902 (N_3902,In_443,In_970);
xor U3903 (N_3903,In_869,In_128);
or U3904 (N_3904,In_252,In_374);
and U3905 (N_3905,In_74,In_289);
nand U3906 (N_3906,In_175,In_612);
or U3907 (N_3907,In_302,In_818);
xor U3908 (N_3908,In_427,In_396);
or U3909 (N_3909,In_428,In_50);
or U3910 (N_3910,In_9,In_927);
nand U3911 (N_3911,In_427,In_963);
or U3912 (N_3912,In_851,In_310);
xor U3913 (N_3913,In_410,In_590);
nand U3914 (N_3914,In_99,In_820);
xor U3915 (N_3915,In_972,In_628);
and U3916 (N_3916,In_982,In_226);
or U3917 (N_3917,In_365,In_230);
xor U3918 (N_3918,In_178,In_955);
nand U3919 (N_3919,In_314,In_725);
nor U3920 (N_3920,In_53,In_827);
or U3921 (N_3921,In_713,In_832);
or U3922 (N_3922,In_797,In_936);
nor U3923 (N_3923,In_937,In_59);
nor U3924 (N_3924,In_784,In_100);
nand U3925 (N_3925,In_579,In_33);
xnor U3926 (N_3926,In_214,In_198);
xnor U3927 (N_3927,In_770,In_531);
nor U3928 (N_3928,In_727,In_698);
nand U3929 (N_3929,In_311,In_176);
nand U3930 (N_3930,In_377,In_322);
xnor U3931 (N_3931,In_392,In_954);
xor U3932 (N_3932,In_179,In_364);
or U3933 (N_3933,In_249,In_112);
or U3934 (N_3934,In_29,In_81);
and U3935 (N_3935,In_425,In_263);
or U3936 (N_3936,In_773,In_279);
and U3937 (N_3937,In_443,In_154);
and U3938 (N_3938,In_576,In_530);
or U3939 (N_3939,In_374,In_229);
nor U3940 (N_3940,In_140,In_891);
nand U3941 (N_3941,In_231,In_1);
and U3942 (N_3942,In_699,In_207);
xnor U3943 (N_3943,In_530,In_9);
nor U3944 (N_3944,In_939,In_51);
and U3945 (N_3945,In_95,In_579);
nor U3946 (N_3946,In_947,In_979);
xnor U3947 (N_3947,In_755,In_460);
or U3948 (N_3948,In_397,In_987);
and U3949 (N_3949,In_663,In_839);
or U3950 (N_3950,In_570,In_80);
xnor U3951 (N_3951,In_142,In_197);
nand U3952 (N_3952,In_872,In_982);
and U3953 (N_3953,In_360,In_72);
or U3954 (N_3954,In_16,In_421);
and U3955 (N_3955,In_322,In_588);
and U3956 (N_3956,In_803,In_974);
nor U3957 (N_3957,In_121,In_749);
and U3958 (N_3958,In_359,In_892);
nand U3959 (N_3959,In_610,In_741);
xnor U3960 (N_3960,In_78,In_474);
nor U3961 (N_3961,In_169,In_537);
nor U3962 (N_3962,In_706,In_262);
xor U3963 (N_3963,In_943,In_936);
and U3964 (N_3964,In_451,In_328);
nand U3965 (N_3965,In_104,In_474);
nor U3966 (N_3966,In_122,In_163);
nand U3967 (N_3967,In_857,In_853);
xnor U3968 (N_3968,In_480,In_202);
xnor U3969 (N_3969,In_429,In_594);
nand U3970 (N_3970,In_236,In_968);
nand U3971 (N_3971,In_157,In_449);
nor U3972 (N_3972,In_583,In_279);
nand U3973 (N_3973,In_589,In_124);
xor U3974 (N_3974,In_202,In_147);
nand U3975 (N_3975,In_995,In_748);
nand U3976 (N_3976,In_690,In_520);
and U3977 (N_3977,In_723,In_102);
nor U3978 (N_3978,In_1,In_25);
and U3979 (N_3979,In_862,In_269);
nand U3980 (N_3980,In_45,In_843);
xor U3981 (N_3981,In_614,In_669);
and U3982 (N_3982,In_440,In_884);
or U3983 (N_3983,In_498,In_615);
or U3984 (N_3984,In_66,In_310);
or U3985 (N_3985,In_607,In_428);
xnor U3986 (N_3986,In_397,In_5);
and U3987 (N_3987,In_725,In_499);
xor U3988 (N_3988,In_519,In_208);
and U3989 (N_3989,In_305,In_160);
nand U3990 (N_3990,In_359,In_361);
nand U3991 (N_3991,In_88,In_336);
and U3992 (N_3992,In_373,In_971);
nand U3993 (N_3993,In_683,In_358);
nor U3994 (N_3994,In_75,In_361);
nand U3995 (N_3995,In_637,In_407);
and U3996 (N_3996,In_794,In_74);
nand U3997 (N_3997,In_901,In_322);
xor U3998 (N_3998,In_170,In_797);
nor U3999 (N_3999,In_28,In_749);
or U4000 (N_4000,In_4,In_669);
or U4001 (N_4001,In_712,In_98);
and U4002 (N_4002,In_939,In_556);
xnor U4003 (N_4003,In_451,In_484);
xor U4004 (N_4004,In_605,In_63);
nor U4005 (N_4005,In_535,In_663);
nor U4006 (N_4006,In_828,In_729);
nand U4007 (N_4007,In_889,In_51);
nor U4008 (N_4008,In_330,In_478);
nor U4009 (N_4009,In_880,In_87);
and U4010 (N_4010,In_956,In_853);
and U4011 (N_4011,In_881,In_850);
and U4012 (N_4012,In_744,In_817);
nand U4013 (N_4013,In_317,In_691);
or U4014 (N_4014,In_36,In_976);
nand U4015 (N_4015,In_276,In_901);
nand U4016 (N_4016,In_814,In_950);
xnor U4017 (N_4017,In_283,In_892);
and U4018 (N_4018,In_274,In_91);
nor U4019 (N_4019,In_898,In_112);
nor U4020 (N_4020,In_84,In_339);
and U4021 (N_4021,In_925,In_351);
xnor U4022 (N_4022,In_960,In_243);
nor U4023 (N_4023,In_195,In_870);
nand U4024 (N_4024,In_523,In_691);
and U4025 (N_4025,In_473,In_170);
nor U4026 (N_4026,In_903,In_999);
xnor U4027 (N_4027,In_988,In_939);
or U4028 (N_4028,In_483,In_722);
or U4029 (N_4029,In_166,In_947);
or U4030 (N_4030,In_698,In_967);
or U4031 (N_4031,In_107,In_683);
and U4032 (N_4032,In_359,In_15);
xnor U4033 (N_4033,In_485,In_384);
nand U4034 (N_4034,In_37,In_126);
nand U4035 (N_4035,In_687,In_798);
and U4036 (N_4036,In_993,In_251);
xor U4037 (N_4037,In_906,In_811);
xor U4038 (N_4038,In_599,In_869);
and U4039 (N_4039,In_679,In_451);
nor U4040 (N_4040,In_167,In_61);
nor U4041 (N_4041,In_942,In_441);
nand U4042 (N_4042,In_7,In_876);
nor U4043 (N_4043,In_990,In_906);
and U4044 (N_4044,In_290,In_312);
nand U4045 (N_4045,In_564,In_775);
and U4046 (N_4046,In_350,In_952);
and U4047 (N_4047,In_382,In_22);
nand U4048 (N_4048,In_828,In_61);
nor U4049 (N_4049,In_716,In_747);
or U4050 (N_4050,In_822,In_273);
or U4051 (N_4051,In_277,In_147);
xor U4052 (N_4052,In_591,In_15);
nand U4053 (N_4053,In_909,In_928);
xnor U4054 (N_4054,In_396,In_684);
nand U4055 (N_4055,In_539,In_843);
xor U4056 (N_4056,In_92,In_24);
nor U4057 (N_4057,In_65,In_535);
nor U4058 (N_4058,In_799,In_65);
xnor U4059 (N_4059,In_266,In_898);
xor U4060 (N_4060,In_615,In_322);
or U4061 (N_4061,In_389,In_693);
and U4062 (N_4062,In_990,In_291);
nand U4063 (N_4063,In_808,In_804);
nand U4064 (N_4064,In_771,In_716);
xnor U4065 (N_4065,In_174,In_427);
nand U4066 (N_4066,In_251,In_336);
nor U4067 (N_4067,In_669,In_584);
xnor U4068 (N_4068,In_263,In_481);
nor U4069 (N_4069,In_915,In_82);
nand U4070 (N_4070,In_231,In_614);
xnor U4071 (N_4071,In_476,In_415);
nand U4072 (N_4072,In_924,In_383);
nand U4073 (N_4073,In_565,In_229);
nand U4074 (N_4074,In_42,In_797);
nor U4075 (N_4075,In_740,In_815);
and U4076 (N_4076,In_246,In_379);
or U4077 (N_4077,In_347,In_251);
nand U4078 (N_4078,In_155,In_889);
nor U4079 (N_4079,In_708,In_498);
or U4080 (N_4080,In_408,In_805);
and U4081 (N_4081,In_732,In_914);
or U4082 (N_4082,In_30,In_63);
and U4083 (N_4083,In_42,In_195);
nor U4084 (N_4084,In_418,In_389);
nor U4085 (N_4085,In_782,In_399);
nand U4086 (N_4086,In_66,In_490);
or U4087 (N_4087,In_501,In_533);
xnor U4088 (N_4088,In_838,In_303);
nand U4089 (N_4089,In_352,In_125);
xnor U4090 (N_4090,In_711,In_273);
and U4091 (N_4091,In_403,In_564);
and U4092 (N_4092,In_561,In_149);
xor U4093 (N_4093,In_460,In_961);
or U4094 (N_4094,In_412,In_830);
nor U4095 (N_4095,In_96,In_271);
xor U4096 (N_4096,In_673,In_723);
and U4097 (N_4097,In_959,In_311);
nor U4098 (N_4098,In_427,In_838);
or U4099 (N_4099,In_598,In_610);
nand U4100 (N_4100,In_151,In_206);
xnor U4101 (N_4101,In_395,In_505);
nor U4102 (N_4102,In_436,In_692);
or U4103 (N_4103,In_761,In_807);
nand U4104 (N_4104,In_339,In_831);
nand U4105 (N_4105,In_958,In_865);
and U4106 (N_4106,In_12,In_728);
or U4107 (N_4107,In_917,In_739);
nor U4108 (N_4108,In_531,In_724);
or U4109 (N_4109,In_678,In_489);
and U4110 (N_4110,In_561,In_946);
nand U4111 (N_4111,In_892,In_284);
and U4112 (N_4112,In_765,In_63);
and U4113 (N_4113,In_108,In_305);
nor U4114 (N_4114,In_24,In_9);
nor U4115 (N_4115,In_103,In_77);
and U4116 (N_4116,In_621,In_841);
nand U4117 (N_4117,In_807,In_287);
xor U4118 (N_4118,In_943,In_977);
nor U4119 (N_4119,In_181,In_385);
or U4120 (N_4120,In_473,In_245);
nand U4121 (N_4121,In_580,In_884);
xnor U4122 (N_4122,In_817,In_218);
nor U4123 (N_4123,In_989,In_288);
xnor U4124 (N_4124,In_851,In_743);
nor U4125 (N_4125,In_233,In_755);
or U4126 (N_4126,In_803,In_405);
xor U4127 (N_4127,In_30,In_536);
nor U4128 (N_4128,In_663,In_671);
and U4129 (N_4129,In_565,In_612);
nand U4130 (N_4130,In_49,In_305);
xor U4131 (N_4131,In_217,In_310);
xor U4132 (N_4132,In_19,In_331);
or U4133 (N_4133,In_189,In_162);
or U4134 (N_4134,In_555,In_543);
nand U4135 (N_4135,In_657,In_176);
xnor U4136 (N_4136,In_801,In_588);
xnor U4137 (N_4137,In_296,In_167);
xnor U4138 (N_4138,In_630,In_935);
xnor U4139 (N_4139,In_290,In_856);
nor U4140 (N_4140,In_207,In_541);
and U4141 (N_4141,In_953,In_450);
or U4142 (N_4142,In_800,In_30);
nand U4143 (N_4143,In_399,In_787);
nand U4144 (N_4144,In_993,In_383);
and U4145 (N_4145,In_793,In_949);
or U4146 (N_4146,In_747,In_476);
and U4147 (N_4147,In_401,In_957);
xnor U4148 (N_4148,In_530,In_270);
xnor U4149 (N_4149,In_896,In_195);
nand U4150 (N_4150,In_146,In_185);
nor U4151 (N_4151,In_105,In_257);
xor U4152 (N_4152,In_440,In_73);
nand U4153 (N_4153,In_760,In_572);
xnor U4154 (N_4154,In_91,In_514);
or U4155 (N_4155,In_326,In_698);
and U4156 (N_4156,In_814,In_425);
nand U4157 (N_4157,In_486,In_870);
and U4158 (N_4158,In_744,In_159);
or U4159 (N_4159,In_355,In_99);
nor U4160 (N_4160,In_763,In_328);
or U4161 (N_4161,In_611,In_714);
xnor U4162 (N_4162,In_790,In_127);
and U4163 (N_4163,In_66,In_154);
and U4164 (N_4164,In_767,In_321);
nand U4165 (N_4165,In_645,In_909);
or U4166 (N_4166,In_484,In_871);
xor U4167 (N_4167,In_624,In_401);
nand U4168 (N_4168,In_999,In_211);
nor U4169 (N_4169,In_668,In_744);
nor U4170 (N_4170,In_723,In_720);
and U4171 (N_4171,In_608,In_683);
or U4172 (N_4172,In_319,In_350);
or U4173 (N_4173,In_657,In_281);
and U4174 (N_4174,In_553,In_483);
xnor U4175 (N_4175,In_323,In_775);
and U4176 (N_4176,In_246,In_514);
nand U4177 (N_4177,In_879,In_426);
or U4178 (N_4178,In_577,In_949);
and U4179 (N_4179,In_75,In_928);
xor U4180 (N_4180,In_546,In_136);
nor U4181 (N_4181,In_802,In_242);
xor U4182 (N_4182,In_937,In_254);
or U4183 (N_4183,In_812,In_188);
xor U4184 (N_4184,In_417,In_491);
nor U4185 (N_4185,In_988,In_490);
nand U4186 (N_4186,In_320,In_656);
or U4187 (N_4187,In_457,In_522);
or U4188 (N_4188,In_949,In_619);
or U4189 (N_4189,In_149,In_192);
and U4190 (N_4190,In_810,In_306);
nand U4191 (N_4191,In_618,In_178);
or U4192 (N_4192,In_982,In_89);
or U4193 (N_4193,In_133,In_260);
and U4194 (N_4194,In_420,In_581);
and U4195 (N_4195,In_784,In_414);
nor U4196 (N_4196,In_798,In_424);
or U4197 (N_4197,In_626,In_133);
and U4198 (N_4198,In_468,In_415);
xor U4199 (N_4199,In_702,In_764);
xor U4200 (N_4200,In_759,In_99);
nor U4201 (N_4201,In_956,In_150);
xnor U4202 (N_4202,In_480,In_698);
and U4203 (N_4203,In_942,In_808);
xor U4204 (N_4204,In_438,In_646);
and U4205 (N_4205,In_878,In_309);
or U4206 (N_4206,In_168,In_237);
xnor U4207 (N_4207,In_248,In_294);
nor U4208 (N_4208,In_694,In_817);
xnor U4209 (N_4209,In_442,In_450);
xor U4210 (N_4210,In_386,In_433);
nor U4211 (N_4211,In_790,In_351);
xor U4212 (N_4212,In_151,In_99);
and U4213 (N_4213,In_606,In_396);
xnor U4214 (N_4214,In_799,In_413);
nand U4215 (N_4215,In_204,In_957);
and U4216 (N_4216,In_763,In_911);
xor U4217 (N_4217,In_941,In_90);
xor U4218 (N_4218,In_338,In_203);
nor U4219 (N_4219,In_916,In_122);
nor U4220 (N_4220,In_367,In_400);
nand U4221 (N_4221,In_5,In_938);
and U4222 (N_4222,In_947,In_587);
nand U4223 (N_4223,In_903,In_210);
xnor U4224 (N_4224,In_86,In_202);
and U4225 (N_4225,In_857,In_640);
nand U4226 (N_4226,In_437,In_886);
xor U4227 (N_4227,In_313,In_739);
nor U4228 (N_4228,In_877,In_904);
nor U4229 (N_4229,In_421,In_325);
or U4230 (N_4230,In_359,In_654);
nand U4231 (N_4231,In_661,In_54);
nand U4232 (N_4232,In_949,In_687);
or U4233 (N_4233,In_91,In_689);
nand U4234 (N_4234,In_413,In_461);
nor U4235 (N_4235,In_699,In_916);
xor U4236 (N_4236,In_115,In_422);
nor U4237 (N_4237,In_690,In_485);
nand U4238 (N_4238,In_668,In_941);
nand U4239 (N_4239,In_710,In_518);
and U4240 (N_4240,In_595,In_370);
xnor U4241 (N_4241,In_741,In_31);
and U4242 (N_4242,In_961,In_508);
and U4243 (N_4243,In_521,In_503);
nand U4244 (N_4244,In_977,In_114);
and U4245 (N_4245,In_773,In_578);
nand U4246 (N_4246,In_372,In_826);
xor U4247 (N_4247,In_594,In_673);
nand U4248 (N_4248,In_747,In_188);
or U4249 (N_4249,In_681,In_627);
or U4250 (N_4250,In_970,In_413);
and U4251 (N_4251,In_833,In_786);
and U4252 (N_4252,In_325,In_221);
xnor U4253 (N_4253,In_81,In_921);
nand U4254 (N_4254,In_54,In_158);
and U4255 (N_4255,In_521,In_998);
nor U4256 (N_4256,In_986,In_384);
and U4257 (N_4257,In_177,In_433);
nand U4258 (N_4258,In_229,In_497);
nor U4259 (N_4259,In_974,In_787);
nor U4260 (N_4260,In_30,In_812);
nor U4261 (N_4261,In_45,In_679);
and U4262 (N_4262,In_825,In_730);
xor U4263 (N_4263,In_850,In_150);
and U4264 (N_4264,In_307,In_207);
or U4265 (N_4265,In_68,In_90);
and U4266 (N_4266,In_854,In_189);
nand U4267 (N_4267,In_716,In_419);
xnor U4268 (N_4268,In_974,In_242);
and U4269 (N_4269,In_446,In_903);
nand U4270 (N_4270,In_664,In_688);
nand U4271 (N_4271,In_447,In_523);
nor U4272 (N_4272,In_246,In_333);
nand U4273 (N_4273,In_728,In_295);
xor U4274 (N_4274,In_343,In_409);
nor U4275 (N_4275,In_977,In_266);
nor U4276 (N_4276,In_857,In_807);
xnor U4277 (N_4277,In_359,In_709);
nor U4278 (N_4278,In_666,In_214);
and U4279 (N_4279,In_95,In_160);
nor U4280 (N_4280,In_98,In_879);
or U4281 (N_4281,In_561,In_351);
xor U4282 (N_4282,In_499,In_170);
or U4283 (N_4283,In_27,In_423);
or U4284 (N_4284,In_780,In_281);
xnor U4285 (N_4285,In_869,In_973);
or U4286 (N_4286,In_160,In_436);
nor U4287 (N_4287,In_578,In_326);
xnor U4288 (N_4288,In_625,In_304);
nand U4289 (N_4289,In_673,In_362);
nand U4290 (N_4290,In_639,In_955);
nand U4291 (N_4291,In_136,In_543);
and U4292 (N_4292,In_49,In_947);
nand U4293 (N_4293,In_61,In_293);
and U4294 (N_4294,In_125,In_270);
nand U4295 (N_4295,In_111,In_799);
or U4296 (N_4296,In_714,In_327);
nand U4297 (N_4297,In_819,In_37);
and U4298 (N_4298,In_680,In_466);
nand U4299 (N_4299,In_839,In_39);
nand U4300 (N_4300,In_733,In_215);
nor U4301 (N_4301,In_540,In_526);
and U4302 (N_4302,In_512,In_433);
nand U4303 (N_4303,In_243,In_204);
nor U4304 (N_4304,In_121,In_997);
nand U4305 (N_4305,In_714,In_747);
and U4306 (N_4306,In_275,In_270);
nor U4307 (N_4307,In_719,In_471);
and U4308 (N_4308,In_655,In_861);
nand U4309 (N_4309,In_87,In_328);
and U4310 (N_4310,In_638,In_202);
xor U4311 (N_4311,In_235,In_292);
and U4312 (N_4312,In_724,In_556);
nand U4313 (N_4313,In_617,In_283);
xor U4314 (N_4314,In_232,In_996);
nor U4315 (N_4315,In_620,In_93);
nand U4316 (N_4316,In_953,In_567);
nor U4317 (N_4317,In_76,In_647);
and U4318 (N_4318,In_503,In_536);
nand U4319 (N_4319,In_65,In_507);
nor U4320 (N_4320,In_626,In_994);
nor U4321 (N_4321,In_991,In_139);
and U4322 (N_4322,In_826,In_467);
xor U4323 (N_4323,In_928,In_311);
nor U4324 (N_4324,In_685,In_607);
and U4325 (N_4325,In_253,In_730);
nor U4326 (N_4326,In_498,In_146);
nor U4327 (N_4327,In_452,In_830);
nor U4328 (N_4328,In_176,In_202);
and U4329 (N_4329,In_744,In_809);
nor U4330 (N_4330,In_29,In_901);
or U4331 (N_4331,In_756,In_537);
and U4332 (N_4332,In_279,In_145);
nor U4333 (N_4333,In_441,In_587);
nor U4334 (N_4334,In_285,In_392);
or U4335 (N_4335,In_664,In_308);
and U4336 (N_4336,In_287,In_11);
nor U4337 (N_4337,In_642,In_899);
and U4338 (N_4338,In_808,In_564);
nor U4339 (N_4339,In_575,In_321);
and U4340 (N_4340,In_611,In_491);
and U4341 (N_4341,In_779,In_200);
and U4342 (N_4342,In_554,In_925);
nor U4343 (N_4343,In_734,In_925);
nand U4344 (N_4344,In_377,In_623);
and U4345 (N_4345,In_733,In_10);
nand U4346 (N_4346,In_848,In_918);
xnor U4347 (N_4347,In_932,In_736);
and U4348 (N_4348,In_500,In_258);
nand U4349 (N_4349,In_461,In_701);
xor U4350 (N_4350,In_906,In_612);
nor U4351 (N_4351,In_664,In_690);
or U4352 (N_4352,In_262,In_875);
nor U4353 (N_4353,In_771,In_997);
and U4354 (N_4354,In_38,In_472);
xor U4355 (N_4355,In_669,In_660);
nor U4356 (N_4356,In_922,In_838);
nand U4357 (N_4357,In_797,In_556);
nand U4358 (N_4358,In_679,In_868);
or U4359 (N_4359,In_410,In_461);
nand U4360 (N_4360,In_913,In_702);
nand U4361 (N_4361,In_747,In_229);
nor U4362 (N_4362,In_697,In_894);
xnor U4363 (N_4363,In_71,In_963);
xor U4364 (N_4364,In_766,In_346);
nand U4365 (N_4365,In_526,In_402);
xnor U4366 (N_4366,In_573,In_756);
or U4367 (N_4367,In_757,In_938);
nand U4368 (N_4368,In_521,In_936);
xnor U4369 (N_4369,In_154,In_340);
and U4370 (N_4370,In_895,In_893);
nor U4371 (N_4371,In_982,In_551);
and U4372 (N_4372,In_77,In_432);
xor U4373 (N_4373,In_770,In_683);
or U4374 (N_4374,In_403,In_937);
nor U4375 (N_4375,In_130,In_594);
nor U4376 (N_4376,In_831,In_704);
nand U4377 (N_4377,In_274,In_396);
xor U4378 (N_4378,In_361,In_40);
nor U4379 (N_4379,In_375,In_856);
xor U4380 (N_4380,In_159,In_107);
and U4381 (N_4381,In_215,In_65);
xor U4382 (N_4382,In_29,In_257);
nand U4383 (N_4383,In_921,In_564);
or U4384 (N_4384,In_829,In_648);
nor U4385 (N_4385,In_614,In_915);
and U4386 (N_4386,In_32,In_972);
and U4387 (N_4387,In_371,In_19);
or U4388 (N_4388,In_457,In_615);
nand U4389 (N_4389,In_408,In_482);
nand U4390 (N_4390,In_407,In_539);
and U4391 (N_4391,In_404,In_139);
or U4392 (N_4392,In_728,In_962);
xnor U4393 (N_4393,In_0,In_280);
nand U4394 (N_4394,In_83,In_828);
nand U4395 (N_4395,In_897,In_252);
xor U4396 (N_4396,In_78,In_268);
nand U4397 (N_4397,In_447,In_899);
and U4398 (N_4398,In_107,In_993);
xor U4399 (N_4399,In_316,In_405);
and U4400 (N_4400,In_483,In_236);
and U4401 (N_4401,In_340,In_332);
or U4402 (N_4402,In_674,In_145);
and U4403 (N_4403,In_422,In_446);
nand U4404 (N_4404,In_675,In_903);
nand U4405 (N_4405,In_617,In_197);
or U4406 (N_4406,In_825,In_644);
and U4407 (N_4407,In_615,In_352);
or U4408 (N_4408,In_451,In_736);
and U4409 (N_4409,In_210,In_346);
and U4410 (N_4410,In_865,In_154);
nand U4411 (N_4411,In_279,In_156);
xor U4412 (N_4412,In_793,In_157);
or U4413 (N_4413,In_882,In_405);
nand U4414 (N_4414,In_88,In_768);
nand U4415 (N_4415,In_331,In_241);
nand U4416 (N_4416,In_548,In_815);
xnor U4417 (N_4417,In_825,In_651);
nor U4418 (N_4418,In_5,In_239);
nor U4419 (N_4419,In_972,In_806);
nand U4420 (N_4420,In_364,In_947);
and U4421 (N_4421,In_700,In_677);
and U4422 (N_4422,In_900,In_561);
xnor U4423 (N_4423,In_963,In_906);
nor U4424 (N_4424,In_518,In_816);
or U4425 (N_4425,In_839,In_820);
and U4426 (N_4426,In_915,In_239);
or U4427 (N_4427,In_736,In_523);
nand U4428 (N_4428,In_894,In_63);
xor U4429 (N_4429,In_166,In_603);
xor U4430 (N_4430,In_850,In_55);
nor U4431 (N_4431,In_626,In_28);
xor U4432 (N_4432,In_460,In_411);
xor U4433 (N_4433,In_343,In_842);
nand U4434 (N_4434,In_771,In_172);
xnor U4435 (N_4435,In_490,In_604);
or U4436 (N_4436,In_963,In_606);
xor U4437 (N_4437,In_349,In_598);
xor U4438 (N_4438,In_169,In_292);
nor U4439 (N_4439,In_494,In_959);
nand U4440 (N_4440,In_14,In_870);
nor U4441 (N_4441,In_716,In_144);
nand U4442 (N_4442,In_550,In_163);
or U4443 (N_4443,In_131,In_304);
and U4444 (N_4444,In_438,In_375);
nor U4445 (N_4445,In_926,In_344);
xnor U4446 (N_4446,In_819,In_352);
nand U4447 (N_4447,In_832,In_6);
or U4448 (N_4448,In_541,In_804);
nand U4449 (N_4449,In_566,In_676);
or U4450 (N_4450,In_158,In_288);
xor U4451 (N_4451,In_169,In_778);
nor U4452 (N_4452,In_689,In_971);
or U4453 (N_4453,In_181,In_270);
nor U4454 (N_4454,In_965,In_491);
or U4455 (N_4455,In_521,In_717);
or U4456 (N_4456,In_927,In_860);
nor U4457 (N_4457,In_378,In_153);
nor U4458 (N_4458,In_100,In_459);
nand U4459 (N_4459,In_846,In_591);
or U4460 (N_4460,In_630,In_143);
nand U4461 (N_4461,In_29,In_615);
nor U4462 (N_4462,In_922,In_449);
and U4463 (N_4463,In_958,In_907);
xor U4464 (N_4464,In_997,In_363);
or U4465 (N_4465,In_503,In_5);
nand U4466 (N_4466,In_17,In_207);
and U4467 (N_4467,In_263,In_908);
nor U4468 (N_4468,In_663,In_917);
xor U4469 (N_4469,In_254,In_621);
or U4470 (N_4470,In_954,In_254);
or U4471 (N_4471,In_62,In_832);
nand U4472 (N_4472,In_428,In_834);
xor U4473 (N_4473,In_691,In_358);
nand U4474 (N_4474,In_218,In_256);
nor U4475 (N_4475,In_774,In_872);
nor U4476 (N_4476,In_158,In_754);
or U4477 (N_4477,In_94,In_567);
nor U4478 (N_4478,In_328,In_137);
nor U4479 (N_4479,In_121,In_419);
xor U4480 (N_4480,In_12,In_44);
xnor U4481 (N_4481,In_145,In_32);
or U4482 (N_4482,In_29,In_978);
xor U4483 (N_4483,In_217,In_398);
xnor U4484 (N_4484,In_900,In_177);
and U4485 (N_4485,In_965,In_696);
nor U4486 (N_4486,In_38,In_460);
or U4487 (N_4487,In_605,In_727);
nor U4488 (N_4488,In_542,In_371);
xor U4489 (N_4489,In_319,In_490);
xor U4490 (N_4490,In_284,In_574);
xor U4491 (N_4491,In_598,In_747);
xor U4492 (N_4492,In_719,In_415);
and U4493 (N_4493,In_539,In_94);
nor U4494 (N_4494,In_387,In_850);
nor U4495 (N_4495,In_814,In_303);
or U4496 (N_4496,In_207,In_688);
and U4497 (N_4497,In_79,In_975);
or U4498 (N_4498,In_47,In_242);
or U4499 (N_4499,In_564,In_440);
nand U4500 (N_4500,In_514,In_440);
xnor U4501 (N_4501,In_925,In_23);
or U4502 (N_4502,In_645,In_509);
xor U4503 (N_4503,In_235,In_117);
xor U4504 (N_4504,In_901,In_798);
or U4505 (N_4505,In_542,In_241);
or U4506 (N_4506,In_345,In_367);
or U4507 (N_4507,In_64,In_409);
or U4508 (N_4508,In_808,In_832);
or U4509 (N_4509,In_793,In_507);
nor U4510 (N_4510,In_210,In_456);
nand U4511 (N_4511,In_588,In_297);
xnor U4512 (N_4512,In_383,In_453);
nor U4513 (N_4513,In_401,In_408);
nand U4514 (N_4514,In_840,In_964);
and U4515 (N_4515,In_554,In_868);
or U4516 (N_4516,In_877,In_779);
xor U4517 (N_4517,In_515,In_431);
nand U4518 (N_4518,In_336,In_61);
and U4519 (N_4519,In_102,In_194);
and U4520 (N_4520,In_599,In_791);
nor U4521 (N_4521,In_190,In_127);
nor U4522 (N_4522,In_870,In_948);
or U4523 (N_4523,In_94,In_3);
nor U4524 (N_4524,In_210,In_448);
or U4525 (N_4525,In_243,In_186);
nor U4526 (N_4526,In_312,In_837);
nand U4527 (N_4527,In_744,In_583);
and U4528 (N_4528,In_23,In_401);
nor U4529 (N_4529,In_443,In_982);
nor U4530 (N_4530,In_846,In_893);
nor U4531 (N_4531,In_707,In_313);
nand U4532 (N_4532,In_81,In_642);
nor U4533 (N_4533,In_126,In_615);
nor U4534 (N_4534,In_922,In_526);
xnor U4535 (N_4535,In_994,In_42);
and U4536 (N_4536,In_63,In_135);
nand U4537 (N_4537,In_840,In_148);
xnor U4538 (N_4538,In_739,In_189);
nand U4539 (N_4539,In_434,In_549);
nor U4540 (N_4540,In_603,In_922);
and U4541 (N_4541,In_615,In_280);
nor U4542 (N_4542,In_51,In_631);
nor U4543 (N_4543,In_863,In_916);
nor U4544 (N_4544,In_555,In_134);
or U4545 (N_4545,In_250,In_310);
xnor U4546 (N_4546,In_807,In_663);
and U4547 (N_4547,In_314,In_73);
nand U4548 (N_4548,In_594,In_487);
nand U4549 (N_4549,In_344,In_883);
nand U4550 (N_4550,In_60,In_733);
xnor U4551 (N_4551,In_446,In_961);
nor U4552 (N_4552,In_496,In_827);
nor U4553 (N_4553,In_770,In_674);
xor U4554 (N_4554,In_493,In_432);
xnor U4555 (N_4555,In_54,In_551);
and U4556 (N_4556,In_862,In_605);
and U4557 (N_4557,In_573,In_708);
xor U4558 (N_4558,In_903,In_31);
nor U4559 (N_4559,In_410,In_518);
nand U4560 (N_4560,In_192,In_520);
or U4561 (N_4561,In_495,In_967);
nand U4562 (N_4562,In_474,In_709);
or U4563 (N_4563,In_674,In_325);
nor U4564 (N_4564,In_660,In_563);
and U4565 (N_4565,In_827,In_485);
nand U4566 (N_4566,In_260,In_210);
nor U4567 (N_4567,In_289,In_258);
nand U4568 (N_4568,In_94,In_988);
nor U4569 (N_4569,In_120,In_870);
nand U4570 (N_4570,In_123,In_482);
nand U4571 (N_4571,In_984,In_745);
and U4572 (N_4572,In_242,In_375);
xor U4573 (N_4573,In_640,In_667);
xnor U4574 (N_4574,In_938,In_552);
nor U4575 (N_4575,In_837,In_200);
nand U4576 (N_4576,In_794,In_813);
or U4577 (N_4577,In_821,In_505);
nand U4578 (N_4578,In_566,In_835);
or U4579 (N_4579,In_459,In_503);
nand U4580 (N_4580,In_902,In_621);
xnor U4581 (N_4581,In_738,In_511);
and U4582 (N_4582,In_537,In_411);
nor U4583 (N_4583,In_137,In_595);
nor U4584 (N_4584,In_18,In_474);
xnor U4585 (N_4585,In_198,In_614);
nand U4586 (N_4586,In_921,In_627);
nand U4587 (N_4587,In_404,In_487);
and U4588 (N_4588,In_38,In_885);
and U4589 (N_4589,In_468,In_348);
xor U4590 (N_4590,In_647,In_736);
nand U4591 (N_4591,In_692,In_177);
and U4592 (N_4592,In_418,In_815);
nor U4593 (N_4593,In_47,In_788);
nand U4594 (N_4594,In_387,In_579);
nand U4595 (N_4595,In_356,In_663);
nand U4596 (N_4596,In_749,In_819);
nor U4597 (N_4597,In_733,In_965);
nand U4598 (N_4598,In_354,In_669);
nand U4599 (N_4599,In_552,In_746);
nand U4600 (N_4600,In_809,In_548);
or U4601 (N_4601,In_969,In_208);
nand U4602 (N_4602,In_520,In_124);
xnor U4603 (N_4603,In_15,In_958);
and U4604 (N_4604,In_241,In_413);
xnor U4605 (N_4605,In_322,In_990);
or U4606 (N_4606,In_73,In_850);
or U4607 (N_4607,In_281,In_714);
or U4608 (N_4608,In_929,In_586);
and U4609 (N_4609,In_127,In_824);
nand U4610 (N_4610,In_142,In_203);
nand U4611 (N_4611,In_857,In_390);
xnor U4612 (N_4612,In_101,In_983);
xnor U4613 (N_4613,In_723,In_646);
nor U4614 (N_4614,In_868,In_874);
nand U4615 (N_4615,In_325,In_311);
xnor U4616 (N_4616,In_984,In_317);
xnor U4617 (N_4617,In_570,In_83);
or U4618 (N_4618,In_425,In_50);
nor U4619 (N_4619,In_596,In_461);
nand U4620 (N_4620,In_359,In_218);
xnor U4621 (N_4621,In_688,In_378);
nand U4622 (N_4622,In_44,In_482);
nand U4623 (N_4623,In_975,In_880);
nand U4624 (N_4624,In_511,In_657);
and U4625 (N_4625,In_917,In_338);
or U4626 (N_4626,In_232,In_168);
or U4627 (N_4627,In_992,In_363);
and U4628 (N_4628,In_750,In_272);
nor U4629 (N_4629,In_933,In_702);
and U4630 (N_4630,In_60,In_482);
or U4631 (N_4631,In_897,In_18);
nor U4632 (N_4632,In_105,In_449);
and U4633 (N_4633,In_381,In_476);
or U4634 (N_4634,In_511,In_923);
nor U4635 (N_4635,In_672,In_34);
nor U4636 (N_4636,In_794,In_394);
and U4637 (N_4637,In_915,In_651);
xnor U4638 (N_4638,In_693,In_203);
nor U4639 (N_4639,In_999,In_122);
and U4640 (N_4640,In_811,In_68);
and U4641 (N_4641,In_284,In_800);
and U4642 (N_4642,In_88,In_579);
and U4643 (N_4643,In_437,In_808);
or U4644 (N_4644,In_629,In_848);
and U4645 (N_4645,In_754,In_43);
or U4646 (N_4646,In_784,In_826);
or U4647 (N_4647,In_775,In_89);
and U4648 (N_4648,In_747,In_78);
and U4649 (N_4649,In_626,In_89);
nor U4650 (N_4650,In_801,In_819);
or U4651 (N_4651,In_989,In_781);
and U4652 (N_4652,In_498,In_145);
nor U4653 (N_4653,In_169,In_755);
or U4654 (N_4654,In_74,In_967);
or U4655 (N_4655,In_319,In_926);
or U4656 (N_4656,In_33,In_307);
xor U4657 (N_4657,In_239,In_71);
and U4658 (N_4658,In_272,In_522);
nand U4659 (N_4659,In_381,In_711);
and U4660 (N_4660,In_559,In_196);
or U4661 (N_4661,In_189,In_688);
or U4662 (N_4662,In_869,In_214);
nand U4663 (N_4663,In_273,In_226);
or U4664 (N_4664,In_213,In_271);
or U4665 (N_4665,In_56,In_481);
nor U4666 (N_4666,In_125,In_670);
nand U4667 (N_4667,In_229,In_463);
and U4668 (N_4668,In_178,In_470);
xnor U4669 (N_4669,In_962,In_987);
or U4670 (N_4670,In_964,In_644);
or U4671 (N_4671,In_464,In_318);
nand U4672 (N_4672,In_244,In_639);
nor U4673 (N_4673,In_121,In_490);
nor U4674 (N_4674,In_779,In_378);
nand U4675 (N_4675,In_385,In_735);
xor U4676 (N_4676,In_278,In_197);
nor U4677 (N_4677,In_700,In_95);
and U4678 (N_4678,In_610,In_162);
nor U4679 (N_4679,In_732,In_121);
nand U4680 (N_4680,In_352,In_906);
or U4681 (N_4681,In_877,In_332);
nor U4682 (N_4682,In_886,In_125);
nand U4683 (N_4683,In_277,In_535);
or U4684 (N_4684,In_935,In_27);
nand U4685 (N_4685,In_684,In_580);
xor U4686 (N_4686,In_418,In_638);
nand U4687 (N_4687,In_970,In_9);
and U4688 (N_4688,In_917,In_346);
xor U4689 (N_4689,In_855,In_651);
and U4690 (N_4690,In_696,In_61);
nand U4691 (N_4691,In_8,In_393);
nor U4692 (N_4692,In_597,In_814);
or U4693 (N_4693,In_511,In_733);
or U4694 (N_4694,In_347,In_908);
and U4695 (N_4695,In_423,In_509);
and U4696 (N_4696,In_215,In_691);
xnor U4697 (N_4697,In_740,In_57);
or U4698 (N_4698,In_477,In_432);
nand U4699 (N_4699,In_733,In_148);
xnor U4700 (N_4700,In_721,In_404);
xnor U4701 (N_4701,In_159,In_228);
nor U4702 (N_4702,In_442,In_344);
or U4703 (N_4703,In_537,In_731);
and U4704 (N_4704,In_887,In_984);
and U4705 (N_4705,In_885,In_929);
and U4706 (N_4706,In_905,In_533);
nor U4707 (N_4707,In_577,In_699);
nor U4708 (N_4708,In_933,In_846);
nand U4709 (N_4709,In_266,In_459);
and U4710 (N_4710,In_648,In_480);
xnor U4711 (N_4711,In_390,In_634);
and U4712 (N_4712,In_193,In_209);
nand U4713 (N_4713,In_188,In_739);
nand U4714 (N_4714,In_500,In_537);
and U4715 (N_4715,In_830,In_379);
nor U4716 (N_4716,In_833,In_71);
or U4717 (N_4717,In_897,In_820);
and U4718 (N_4718,In_964,In_571);
nor U4719 (N_4719,In_256,In_862);
and U4720 (N_4720,In_802,In_283);
or U4721 (N_4721,In_168,In_81);
or U4722 (N_4722,In_352,In_286);
nand U4723 (N_4723,In_248,In_429);
nand U4724 (N_4724,In_167,In_346);
nor U4725 (N_4725,In_196,In_97);
and U4726 (N_4726,In_43,In_211);
nand U4727 (N_4727,In_454,In_227);
nand U4728 (N_4728,In_424,In_288);
or U4729 (N_4729,In_333,In_252);
and U4730 (N_4730,In_502,In_434);
xnor U4731 (N_4731,In_425,In_501);
or U4732 (N_4732,In_325,In_428);
nor U4733 (N_4733,In_526,In_84);
nand U4734 (N_4734,In_879,In_531);
nor U4735 (N_4735,In_76,In_567);
xnor U4736 (N_4736,In_541,In_245);
nand U4737 (N_4737,In_548,In_987);
or U4738 (N_4738,In_89,In_299);
xnor U4739 (N_4739,In_392,In_949);
or U4740 (N_4740,In_775,In_568);
and U4741 (N_4741,In_270,In_165);
xor U4742 (N_4742,In_772,In_448);
and U4743 (N_4743,In_306,In_866);
or U4744 (N_4744,In_653,In_292);
xor U4745 (N_4745,In_704,In_442);
nor U4746 (N_4746,In_246,In_183);
xnor U4747 (N_4747,In_403,In_149);
nor U4748 (N_4748,In_962,In_67);
or U4749 (N_4749,In_957,In_97);
xnor U4750 (N_4750,In_7,In_94);
nand U4751 (N_4751,In_549,In_646);
and U4752 (N_4752,In_589,In_592);
nand U4753 (N_4753,In_602,In_641);
and U4754 (N_4754,In_678,In_693);
or U4755 (N_4755,In_0,In_222);
or U4756 (N_4756,In_758,In_636);
xor U4757 (N_4757,In_847,In_63);
nor U4758 (N_4758,In_137,In_704);
nand U4759 (N_4759,In_268,In_613);
and U4760 (N_4760,In_828,In_655);
and U4761 (N_4761,In_775,In_237);
and U4762 (N_4762,In_566,In_357);
or U4763 (N_4763,In_895,In_18);
xor U4764 (N_4764,In_891,In_173);
nand U4765 (N_4765,In_663,In_643);
and U4766 (N_4766,In_951,In_494);
xnor U4767 (N_4767,In_627,In_908);
nand U4768 (N_4768,In_420,In_737);
or U4769 (N_4769,In_265,In_773);
nor U4770 (N_4770,In_684,In_56);
xor U4771 (N_4771,In_502,In_435);
nand U4772 (N_4772,In_866,In_451);
nor U4773 (N_4773,In_304,In_387);
or U4774 (N_4774,In_885,In_587);
nand U4775 (N_4775,In_113,In_65);
nand U4776 (N_4776,In_871,In_231);
nor U4777 (N_4777,In_648,In_14);
and U4778 (N_4778,In_295,In_259);
nor U4779 (N_4779,In_889,In_6);
nor U4780 (N_4780,In_164,In_651);
and U4781 (N_4781,In_879,In_530);
or U4782 (N_4782,In_620,In_536);
nor U4783 (N_4783,In_972,In_449);
xnor U4784 (N_4784,In_562,In_595);
xnor U4785 (N_4785,In_434,In_96);
nand U4786 (N_4786,In_202,In_345);
and U4787 (N_4787,In_611,In_285);
and U4788 (N_4788,In_118,In_640);
and U4789 (N_4789,In_394,In_48);
and U4790 (N_4790,In_654,In_127);
xnor U4791 (N_4791,In_729,In_888);
nand U4792 (N_4792,In_915,In_816);
or U4793 (N_4793,In_634,In_960);
nand U4794 (N_4794,In_158,In_693);
nor U4795 (N_4795,In_522,In_206);
nor U4796 (N_4796,In_597,In_474);
nor U4797 (N_4797,In_688,In_467);
xnor U4798 (N_4798,In_539,In_347);
and U4799 (N_4799,In_61,In_395);
nor U4800 (N_4800,In_255,In_176);
xnor U4801 (N_4801,In_487,In_148);
nand U4802 (N_4802,In_221,In_808);
xor U4803 (N_4803,In_742,In_134);
nor U4804 (N_4804,In_817,In_64);
nand U4805 (N_4805,In_529,In_735);
or U4806 (N_4806,In_156,In_282);
and U4807 (N_4807,In_704,In_954);
nand U4808 (N_4808,In_9,In_886);
nand U4809 (N_4809,In_888,In_323);
or U4810 (N_4810,In_696,In_582);
or U4811 (N_4811,In_567,In_321);
and U4812 (N_4812,In_266,In_119);
xor U4813 (N_4813,In_759,In_52);
nand U4814 (N_4814,In_530,In_520);
xnor U4815 (N_4815,In_380,In_447);
xor U4816 (N_4816,In_823,In_683);
or U4817 (N_4817,In_655,In_590);
nor U4818 (N_4818,In_159,In_239);
nor U4819 (N_4819,In_510,In_966);
or U4820 (N_4820,In_828,In_721);
nor U4821 (N_4821,In_113,In_311);
xnor U4822 (N_4822,In_923,In_271);
xnor U4823 (N_4823,In_5,In_357);
nand U4824 (N_4824,In_191,In_291);
nand U4825 (N_4825,In_946,In_204);
and U4826 (N_4826,In_858,In_371);
nor U4827 (N_4827,In_825,In_101);
xnor U4828 (N_4828,In_721,In_762);
nand U4829 (N_4829,In_498,In_867);
or U4830 (N_4830,In_323,In_9);
or U4831 (N_4831,In_909,In_538);
and U4832 (N_4832,In_915,In_88);
nor U4833 (N_4833,In_535,In_955);
nand U4834 (N_4834,In_738,In_777);
and U4835 (N_4835,In_389,In_631);
or U4836 (N_4836,In_377,In_512);
xor U4837 (N_4837,In_535,In_746);
and U4838 (N_4838,In_467,In_947);
nor U4839 (N_4839,In_675,In_562);
and U4840 (N_4840,In_381,In_398);
xnor U4841 (N_4841,In_268,In_752);
or U4842 (N_4842,In_102,In_297);
and U4843 (N_4843,In_894,In_661);
or U4844 (N_4844,In_966,In_691);
and U4845 (N_4845,In_246,In_478);
nand U4846 (N_4846,In_321,In_800);
xor U4847 (N_4847,In_375,In_711);
or U4848 (N_4848,In_878,In_679);
and U4849 (N_4849,In_330,In_101);
and U4850 (N_4850,In_425,In_331);
or U4851 (N_4851,In_276,In_644);
or U4852 (N_4852,In_291,In_108);
or U4853 (N_4853,In_476,In_228);
xnor U4854 (N_4854,In_983,In_405);
nor U4855 (N_4855,In_125,In_799);
nand U4856 (N_4856,In_460,In_633);
nand U4857 (N_4857,In_439,In_264);
nor U4858 (N_4858,In_481,In_113);
nand U4859 (N_4859,In_505,In_476);
and U4860 (N_4860,In_394,In_181);
nor U4861 (N_4861,In_291,In_200);
and U4862 (N_4862,In_750,In_330);
or U4863 (N_4863,In_85,In_685);
xor U4864 (N_4864,In_909,In_631);
nor U4865 (N_4865,In_718,In_479);
xnor U4866 (N_4866,In_455,In_365);
xnor U4867 (N_4867,In_886,In_825);
or U4868 (N_4868,In_730,In_680);
xnor U4869 (N_4869,In_772,In_221);
xnor U4870 (N_4870,In_153,In_870);
nor U4871 (N_4871,In_433,In_491);
xor U4872 (N_4872,In_411,In_847);
xnor U4873 (N_4873,In_118,In_356);
nor U4874 (N_4874,In_611,In_168);
xnor U4875 (N_4875,In_90,In_669);
xnor U4876 (N_4876,In_246,In_870);
and U4877 (N_4877,In_655,In_976);
nand U4878 (N_4878,In_612,In_365);
nor U4879 (N_4879,In_545,In_544);
and U4880 (N_4880,In_594,In_797);
or U4881 (N_4881,In_607,In_998);
nor U4882 (N_4882,In_148,In_598);
and U4883 (N_4883,In_61,In_922);
nor U4884 (N_4884,In_319,In_902);
and U4885 (N_4885,In_635,In_537);
xor U4886 (N_4886,In_111,In_124);
xnor U4887 (N_4887,In_224,In_323);
nand U4888 (N_4888,In_786,In_505);
xnor U4889 (N_4889,In_153,In_646);
xor U4890 (N_4890,In_852,In_923);
nand U4891 (N_4891,In_511,In_87);
xnor U4892 (N_4892,In_114,In_94);
nand U4893 (N_4893,In_564,In_445);
or U4894 (N_4894,In_597,In_38);
or U4895 (N_4895,In_72,In_143);
or U4896 (N_4896,In_135,In_563);
and U4897 (N_4897,In_199,In_965);
xnor U4898 (N_4898,In_538,In_369);
nor U4899 (N_4899,In_876,In_433);
xor U4900 (N_4900,In_145,In_767);
nand U4901 (N_4901,In_990,In_869);
and U4902 (N_4902,In_357,In_576);
nand U4903 (N_4903,In_499,In_370);
nor U4904 (N_4904,In_627,In_541);
xnor U4905 (N_4905,In_805,In_563);
xnor U4906 (N_4906,In_717,In_31);
xnor U4907 (N_4907,In_884,In_998);
xnor U4908 (N_4908,In_252,In_822);
xnor U4909 (N_4909,In_460,In_404);
or U4910 (N_4910,In_904,In_843);
xor U4911 (N_4911,In_130,In_359);
nor U4912 (N_4912,In_583,In_731);
or U4913 (N_4913,In_191,In_484);
xor U4914 (N_4914,In_205,In_658);
xnor U4915 (N_4915,In_417,In_410);
nor U4916 (N_4916,In_404,In_433);
nor U4917 (N_4917,In_796,In_557);
xnor U4918 (N_4918,In_992,In_551);
or U4919 (N_4919,In_380,In_381);
xor U4920 (N_4920,In_33,In_791);
or U4921 (N_4921,In_378,In_916);
nand U4922 (N_4922,In_228,In_685);
or U4923 (N_4923,In_371,In_349);
and U4924 (N_4924,In_119,In_260);
and U4925 (N_4925,In_815,In_539);
nand U4926 (N_4926,In_188,In_822);
or U4927 (N_4927,In_464,In_713);
and U4928 (N_4928,In_365,In_428);
nand U4929 (N_4929,In_680,In_121);
and U4930 (N_4930,In_238,In_495);
and U4931 (N_4931,In_963,In_138);
and U4932 (N_4932,In_944,In_813);
nor U4933 (N_4933,In_192,In_421);
nand U4934 (N_4934,In_570,In_303);
nor U4935 (N_4935,In_361,In_731);
and U4936 (N_4936,In_44,In_142);
and U4937 (N_4937,In_99,In_904);
nand U4938 (N_4938,In_601,In_51);
or U4939 (N_4939,In_966,In_133);
nand U4940 (N_4940,In_103,In_354);
nor U4941 (N_4941,In_963,In_151);
or U4942 (N_4942,In_776,In_522);
nand U4943 (N_4943,In_81,In_839);
and U4944 (N_4944,In_460,In_63);
and U4945 (N_4945,In_504,In_856);
and U4946 (N_4946,In_842,In_952);
and U4947 (N_4947,In_164,In_886);
and U4948 (N_4948,In_230,In_457);
nand U4949 (N_4949,In_750,In_278);
nand U4950 (N_4950,In_819,In_220);
nor U4951 (N_4951,In_615,In_494);
xnor U4952 (N_4952,In_713,In_655);
nor U4953 (N_4953,In_834,In_340);
and U4954 (N_4954,In_434,In_547);
xnor U4955 (N_4955,In_683,In_911);
or U4956 (N_4956,In_381,In_831);
xor U4957 (N_4957,In_403,In_515);
or U4958 (N_4958,In_244,In_632);
and U4959 (N_4959,In_268,In_239);
xor U4960 (N_4960,In_56,In_527);
xor U4961 (N_4961,In_804,In_983);
and U4962 (N_4962,In_270,In_893);
nor U4963 (N_4963,In_851,In_460);
xor U4964 (N_4964,In_430,In_729);
nand U4965 (N_4965,In_606,In_37);
nand U4966 (N_4966,In_116,In_669);
and U4967 (N_4967,In_254,In_715);
and U4968 (N_4968,In_189,In_45);
nor U4969 (N_4969,In_879,In_810);
or U4970 (N_4970,In_706,In_537);
nand U4971 (N_4971,In_488,In_199);
and U4972 (N_4972,In_414,In_605);
or U4973 (N_4973,In_292,In_569);
or U4974 (N_4974,In_417,In_384);
or U4975 (N_4975,In_353,In_229);
xor U4976 (N_4976,In_767,In_245);
and U4977 (N_4977,In_652,In_912);
nand U4978 (N_4978,In_827,In_550);
nand U4979 (N_4979,In_33,In_216);
nand U4980 (N_4980,In_424,In_556);
or U4981 (N_4981,In_643,In_466);
nand U4982 (N_4982,In_180,In_713);
nor U4983 (N_4983,In_836,In_581);
xor U4984 (N_4984,In_70,In_211);
nor U4985 (N_4985,In_869,In_500);
nor U4986 (N_4986,In_40,In_894);
and U4987 (N_4987,In_283,In_321);
or U4988 (N_4988,In_936,In_985);
nor U4989 (N_4989,In_189,In_605);
or U4990 (N_4990,In_449,In_456);
and U4991 (N_4991,In_776,In_661);
xnor U4992 (N_4992,In_123,In_575);
nand U4993 (N_4993,In_465,In_256);
or U4994 (N_4994,In_732,In_842);
nand U4995 (N_4995,In_268,In_320);
or U4996 (N_4996,In_989,In_350);
xor U4997 (N_4997,In_496,In_327);
or U4998 (N_4998,In_581,In_816);
or U4999 (N_4999,In_219,In_256);
or U5000 (N_5000,N_2073,N_1880);
and U5001 (N_5001,N_4159,N_3546);
nor U5002 (N_5002,N_2726,N_4783);
nor U5003 (N_5003,N_1172,N_4083);
nand U5004 (N_5004,N_864,N_1430);
and U5005 (N_5005,N_3132,N_2525);
xor U5006 (N_5006,N_2124,N_1257);
or U5007 (N_5007,N_4796,N_281);
nor U5008 (N_5008,N_194,N_4516);
and U5009 (N_5009,N_345,N_1514);
xor U5010 (N_5010,N_3828,N_2428);
and U5011 (N_5011,N_390,N_3939);
nor U5012 (N_5012,N_2328,N_4471);
or U5013 (N_5013,N_4726,N_1958);
or U5014 (N_5014,N_4180,N_4333);
nand U5015 (N_5015,N_3443,N_1326);
and U5016 (N_5016,N_346,N_1397);
nand U5017 (N_5017,N_1106,N_18);
xnor U5018 (N_5018,N_4293,N_3517);
or U5019 (N_5019,N_4661,N_485);
nand U5020 (N_5020,N_420,N_1310);
xor U5021 (N_5021,N_1267,N_4272);
and U5022 (N_5022,N_1584,N_2893);
or U5023 (N_5023,N_2481,N_3583);
nor U5024 (N_5024,N_476,N_1893);
xnor U5025 (N_5025,N_1329,N_222);
or U5026 (N_5026,N_4693,N_442);
nor U5027 (N_5027,N_545,N_3129);
xnor U5028 (N_5028,N_3815,N_3559);
or U5029 (N_5029,N_2998,N_1647);
or U5030 (N_5030,N_2942,N_4678);
xor U5031 (N_5031,N_976,N_975);
nor U5032 (N_5032,N_338,N_4908);
and U5033 (N_5033,N_2440,N_3216);
nor U5034 (N_5034,N_1130,N_3104);
nand U5035 (N_5035,N_4244,N_3072);
xnor U5036 (N_5036,N_2925,N_3777);
nand U5037 (N_5037,N_1420,N_3200);
or U5038 (N_5038,N_2196,N_3719);
xor U5039 (N_5039,N_3958,N_683);
or U5040 (N_5040,N_2444,N_2483);
and U5041 (N_5041,N_1571,N_326);
nor U5042 (N_5042,N_182,N_1645);
nand U5043 (N_5043,N_788,N_4292);
xor U5044 (N_5044,N_3512,N_943);
nand U5045 (N_5045,N_4323,N_4288);
nor U5046 (N_5046,N_2050,N_4216);
nand U5047 (N_5047,N_4325,N_3511);
or U5048 (N_5048,N_4703,N_718);
nand U5049 (N_5049,N_2777,N_1205);
nor U5050 (N_5050,N_1650,N_144);
xnor U5051 (N_5051,N_2195,N_1895);
xor U5052 (N_5052,N_463,N_664);
xnor U5053 (N_5053,N_4403,N_4740);
xor U5054 (N_5054,N_4009,N_2297);
or U5055 (N_5055,N_2907,N_3769);
nand U5056 (N_5056,N_334,N_758);
nor U5057 (N_5057,N_1460,N_4566);
nand U5058 (N_5058,N_1371,N_4968);
and U5059 (N_5059,N_2127,N_3331);
nand U5060 (N_5060,N_1194,N_806);
nand U5061 (N_5061,N_982,N_1635);
nor U5062 (N_5062,N_777,N_3797);
and U5063 (N_5063,N_698,N_2789);
nor U5064 (N_5064,N_195,N_4922);
and U5065 (N_5065,N_499,N_1579);
xnor U5066 (N_5066,N_2864,N_1742);
and U5067 (N_5067,N_761,N_1570);
xor U5068 (N_5068,N_3606,N_1922);
and U5069 (N_5069,N_2953,N_837);
nor U5070 (N_5070,N_302,N_3526);
and U5071 (N_5071,N_4575,N_79);
nor U5072 (N_5072,N_2778,N_1466);
nand U5073 (N_5073,N_647,N_2429);
xor U5074 (N_5074,N_2075,N_298);
xnor U5075 (N_5075,N_4670,N_2947);
and U5076 (N_5076,N_3148,N_4601);
nor U5077 (N_5077,N_2140,N_2850);
and U5078 (N_5078,N_2593,N_2496);
nor U5079 (N_5079,N_4376,N_4609);
or U5080 (N_5080,N_2467,N_12);
nor U5081 (N_5081,N_3738,N_1015);
nand U5082 (N_5082,N_1588,N_635);
and U5083 (N_5083,N_4849,N_2624);
and U5084 (N_5084,N_3354,N_3370);
or U5085 (N_5085,N_3663,N_2388);
nand U5086 (N_5086,N_4467,N_1608);
nand U5087 (N_5087,N_3409,N_2586);
nand U5088 (N_5088,N_348,N_494);
nand U5089 (N_5089,N_3808,N_2455);
nor U5090 (N_5090,N_4553,N_2457);
nand U5091 (N_5091,N_4161,N_2674);
and U5092 (N_5092,N_2311,N_4058);
nor U5093 (N_5093,N_204,N_1692);
or U5094 (N_5094,N_4195,N_3593);
xnor U5095 (N_5095,N_4228,N_3976);
xor U5096 (N_5096,N_2431,N_3996);
nand U5097 (N_5097,N_3700,N_3854);
xor U5098 (N_5098,N_1667,N_2938);
nand U5099 (N_5099,N_3016,N_4816);
and U5100 (N_5100,N_2543,N_4734);
and U5101 (N_5101,N_4818,N_4565);
and U5102 (N_5102,N_1903,N_3472);
nor U5103 (N_5103,N_1639,N_4508);
nor U5104 (N_5104,N_2748,N_3914);
and U5105 (N_5105,N_2937,N_419);
nor U5106 (N_5106,N_2619,N_1464);
and U5107 (N_5107,N_952,N_2539);
nand U5108 (N_5108,N_1998,N_2280);
or U5109 (N_5109,N_2815,N_1538);
xnor U5110 (N_5110,N_55,N_4128);
nand U5111 (N_5111,N_4250,N_189);
nor U5112 (N_5112,N_3498,N_1687);
and U5113 (N_5113,N_537,N_2693);
nor U5114 (N_5114,N_4976,N_4502);
nor U5115 (N_5115,N_381,N_2191);
or U5116 (N_5116,N_1821,N_4141);
and U5117 (N_5117,N_3225,N_4921);
and U5118 (N_5118,N_4539,N_2057);
or U5119 (N_5119,N_2519,N_2324);
nor U5120 (N_5120,N_944,N_2498);
xnor U5121 (N_5121,N_40,N_1259);
nand U5122 (N_5122,N_2225,N_3131);
xnor U5123 (N_5123,N_3675,N_3991);
or U5124 (N_5124,N_3164,N_1099);
nor U5125 (N_5125,N_4275,N_1127);
xor U5126 (N_5126,N_162,N_4738);
nand U5127 (N_5127,N_1402,N_3199);
nand U5128 (N_5128,N_241,N_388);
or U5129 (N_5129,N_3007,N_532);
nor U5130 (N_5130,N_106,N_1951);
nand U5131 (N_5131,N_4366,N_3144);
nor U5132 (N_5132,N_4540,N_1613);
and U5133 (N_5133,N_4654,N_1715);
or U5134 (N_5134,N_4016,N_3625);
and U5135 (N_5135,N_3706,N_3725);
nor U5136 (N_5136,N_4302,N_3591);
nor U5137 (N_5137,N_4820,N_3403);
and U5138 (N_5138,N_3448,N_4782);
nor U5139 (N_5139,N_2829,N_2474);
nor U5140 (N_5140,N_556,N_4353);
nor U5141 (N_5141,N_3181,N_4551);
xor U5142 (N_5142,N_1707,N_3324);
nand U5143 (N_5143,N_2290,N_3188);
nand U5144 (N_5144,N_4231,N_4252);
xor U5145 (N_5145,N_3080,N_3014);
nor U5146 (N_5146,N_2736,N_921);
nor U5147 (N_5147,N_565,N_2422);
nor U5148 (N_5148,N_876,N_2058);
nand U5149 (N_5149,N_2318,N_1452);
or U5150 (N_5150,N_425,N_2765);
or U5151 (N_5151,N_892,N_2548);
and U5152 (N_5152,N_2838,N_2718);
nor U5153 (N_5153,N_3787,N_1062);
nand U5154 (N_5154,N_1118,N_1000);
xor U5155 (N_5155,N_640,N_2803);
xor U5156 (N_5156,N_4345,N_1449);
nand U5157 (N_5157,N_2197,N_4615);
nand U5158 (N_5158,N_2788,N_626);
nand U5159 (N_5159,N_649,N_2480);
nand U5160 (N_5160,N_2346,N_1197);
nand U5161 (N_5161,N_430,N_1818);
or U5162 (N_5162,N_956,N_437);
and U5163 (N_5163,N_2355,N_1090);
and U5164 (N_5164,N_1658,N_4884);
nand U5165 (N_5165,N_3340,N_109);
or U5166 (N_5166,N_779,N_404);
nor U5167 (N_5167,N_2326,N_2048);
xnor U5168 (N_5168,N_1626,N_1989);
and U5169 (N_5169,N_1427,N_3390);
nand U5170 (N_5170,N_3266,N_2161);
and U5171 (N_5171,N_4148,N_3849);
and U5172 (N_5172,N_3605,N_4057);
nand U5173 (N_5173,N_1157,N_4452);
and U5174 (N_5174,N_4249,N_2147);
nor U5175 (N_5175,N_1132,N_712);
or U5176 (N_5176,N_2226,N_1915);
or U5177 (N_5177,N_3252,N_4567);
nand U5178 (N_5178,N_4001,N_2895);
nand U5179 (N_5179,N_28,N_468);
nor U5180 (N_5180,N_4752,N_2275);
nand U5181 (N_5181,N_1287,N_2700);
xnor U5182 (N_5182,N_4179,N_2660);
nor U5183 (N_5183,N_2514,N_1597);
and U5184 (N_5184,N_1374,N_4318);
nand U5185 (N_5185,N_518,N_96);
nand U5186 (N_5186,N_2308,N_2627);
xor U5187 (N_5187,N_1407,N_2955);
or U5188 (N_5188,N_3649,N_2950);
nand U5189 (N_5189,N_844,N_71);
nor U5190 (N_5190,N_3141,N_3102);
or U5191 (N_5191,N_3933,N_928);
nor U5192 (N_5192,N_399,N_2019);
xnor U5193 (N_5193,N_1731,N_1540);
nor U5194 (N_5194,N_544,N_2361);
xor U5195 (N_5195,N_3342,N_2639);
nand U5196 (N_5196,N_4227,N_1975);
or U5197 (N_5197,N_4483,N_1999);
nand U5198 (N_5198,N_4097,N_1121);
or U5199 (N_5199,N_3088,N_4966);
or U5200 (N_5200,N_321,N_4084);
nand U5201 (N_5201,N_2997,N_2785);
and U5202 (N_5202,N_1049,N_4432);
nand U5203 (N_5203,N_1004,N_4115);
xnor U5204 (N_5204,N_2065,N_2592);
and U5205 (N_5205,N_2042,N_1887);
or U5206 (N_5206,N_2899,N_2077);
nor U5207 (N_5207,N_4264,N_1288);
nand U5208 (N_5208,N_274,N_3634);
or U5209 (N_5209,N_947,N_862);
or U5210 (N_5210,N_3945,N_4929);
or U5211 (N_5211,N_1864,N_1394);
and U5212 (N_5212,N_4205,N_2367);
nor U5213 (N_5213,N_2461,N_3528);
xor U5214 (N_5214,N_2671,N_292);
xnor U5215 (N_5215,N_2745,N_827);
nand U5216 (N_5216,N_4715,N_2632);
nor U5217 (N_5217,N_245,N_1468);
nand U5218 (N_5218,N_583,N_1344);
and U5219 (N_5219,N_3733,N_3315);
or U5220 (N_5220,N_2452,N_4330);
or U5221 (N_5221,N_2106,N_1798);
nand U5222 (N_5222,N_4630,N_4759);
nand U5223 (N_5223,N_3338,N_4639);
or U5224 (N_5224,N_2824,N_3819);
nand U5225 (N_5225,N_2131,N_4582);
nor U5226 (N_5226,N_1438,N_171);
nand U5227 (N_5227,N_2577,N_4418);
and U5228 (N_5228,N_4449,N_695);
and U5229 (N_5229,N_1070,N_3867);
nor U5230 (N_5230,N_3684,N_4979);
and U5231 (N_5231,N_1439,N_838);
and U5232 (N_5232,N_1128,N_475);
xnor U5233 (N_5233,N_8,N_2793);
or U5234 (N_5234,N_4101,N_2049);
nor U5235 (N_5235,N_2951,N_4913);
nor U5236 (N_5236,N_2250,N_873);
nor U5237 (N_5237,N_3516,N_3710);
xnor U5238 (N_5238,N_2218,N_1303);
and U5239 (N_5239,N_193,N_2672);
nor U5240 (N_5240,N_2331,N_2764);
xnor U5241 (N_5241,N_3683,N_2210);
and U5242 (N_5242,N_2766,N_3839);
and U5243 (N_5243,N_3881,N_1446);
nor U5244 (N_5244,N_832,N_1741);
or U5245 (N_5245,N_282,N_3665);
or U5246 (N_5246,N_3647,N_3310);
and U5247 (N_5247,N_3946,N_3553);
and U5248 (N_5248,N_3964,N_1551);
and U5249 (N_5249,N_1255,N_3470);
xor U5250 (N_5250,N_3021,N_4108);
or U5251 (N_5251,N_680,N_2737);
and U5252 (N_5252,N_720,N_402);
and U5253 (N_5253,N_3704,N_4486);
xnor U5254 (N_5254,N_724,N_4380);
nor U5255 (N_5255,N_180,N_3176);
xor U5256 (N_5256,N_2233,N_2258);
and U5257 (N_5257,N_3543,N_2756);
or U5258 (N_5258,N_1227,N_3929);
xnor U5259 (N_5259,N_2060,N_1828);
nor U5260 (N_5260,N_1115,N_347);
nand U5261 (N_5261,N_612,N_1734);
and U5262 (N_5262,N_4812,N_2842);
or U5263 (N_5263,N_2236,N_410);
nand U5264 (N_5264,N_2087,N_660);
and U5265 (N_5265,N_4618,N_3061);
nor U5266 (N_5266,N_3380,N_1523);
nand U5267 (N_5267,N_4807,N_1577);
xnor U5268 (N_5268,N_4861,N_2809);
and U5269 (N_5269,N_1252,N_2387);
nor U5270 (N_5270,N_636,N_14);
or U5271 (N_5271,N_880,N_97);
or U5272 (N_5272,N_3499,N_3573);
nand U5273 (N_5273,N_1988,N_2614);
nor U5274 (N_5274,N_133,N_939);
and U5275 (N_5275,N_4136,N_434);
xor U5276 (N_5276,N_3918,N_901);
xnor U5277 (N_5277,N_479,N_172);
nand U5278 (N_5278,N_3792,N_3533);
xor U5279 (N_5279,N_1116,N_2362);
nor U5280 (N_5280,N_303,N_4521);
and U5281 (N_5281,N_4920,N_2239);
xnor U5282 (N_5282,N_4758,N_4993);
and U5283 (N_5283,N_2634,N_86);
nor U5284 (N_5284,N_4282,N_2464);
xor U5285 (N_5285,N_361,N_2816);
and U5286 (N_5286,N_3239,N_3105);
and U5287 (N_5287,N_3651,N_4623);
and U5288 (N_5288,N_1890,N_4583);
xor U5289 (N_5289,N_2112,N_2611);
or U5290 (N_5290,N_2596,N_3026);
or U5291 (N_5291,N_4204,N_610);
nand U5292 (N_5292,N_4073,N_3008);
and U5293 (N_5293,N_3905,N_1079);
xnor U5294 (N_5294,N_3648,N_4160);
nor U5295 (N_5295,N_673,N_4580);
and U5296 (N_5296,N_2405,N_729);
and U5297 (N_5297,N_696,N_4684);
and U5298 (N_5298,N_3741,N_2932);
or U5299 (N_5299,N_3662,N_3095);
and U5300 (N_5300,N_2980,N_634);
nand U5301 (N_5301,N_2744,N_2890);
nand U5302 (N_5302,N_534,N_4594);
nand U5303 (N_5303,N_2495,N_2635);
xnor U5304 (N_5304,N_4699,N_929);
and U5305 (N_5305,N_161,N_3155);
xnor U5306 (N_5306,N_722,N_159);
xnor U5307 (N_5307,N_1594,N_4042);
nor U5308 (N_5308,N_3742,N_1387);
nand U5309 (N_5309,N_2013,N_3562);
nor U5310 (N_5310,N_4225,N_3465);
nor U5311 (N_5311,N_2833,N_4370);
nor U5312 (N_5312,N_4342,N_3628);
nor U5313 (N_5313,N_3536,N_890);
nand U5314 (N_5314,N_3885,N_3588);
or U5315 (N_5315,N_48,N_2007);
and U5316 (N_5316,N_4835,N_351);
nor U5317 (N_5317,N_4387,N_2101);
and U5318 (N_5318,N_3904,N_3123);
nor U5319 (N_5319,N_4593,N_1307);
xor U5320 (N_5320,N_2409,N_619);
xnor U5321 (N_5321,N_76,N_360);
xor U5322 (N_5322,N_123,N_3635);
or U5323 (N_5323,N_2914,N_887);
xnor U5324 (N_5324,N_503,N_3241);
nand U5325 (N_5325,N_2653,N_1910);
and U5326 (N_5326,N_3373,N_1776);
or U5327 (N_5327,N_820,N_2291);
xor U5328 (N_5328,N_1040,N_869);
xnor U5329 (N_5329,N_4436,N_3408);
nor U5330 (N_5330,N_4197,N_4645);
nand U5331 (N_5331,N_3049,N_176);
xnor U5332 (N_5332,N_396,N_871);
nor U5333 (N_5333,N_459,N_4421);
nor U5334 (N_5334,N_460,N_4675);
xor U5335 (N_5335,N_529,N_3869);
and U5336 (N_5336,N_1974,N_1874);
nand U5337 (N_5337,N_1269,N_694);
xnor U5338 (N_5338,N_4468,N_452);
xor U5339 (N_5339,N_2156,N_4459);
xnor U5340 (N_5340,N_4605,N_3232);
nor U5341 (N_5341,N_1114,N_3886);
and U5342 (N_5342,N_3180,N_386);
or U5343 (N_5343,N_3714,N_4040);
xnor U5344 (N_5344,N_1833,N_1163);
and U5345 (N_5345,N_2000,N_186);
xor U5346 (N_5346,N_1202,N_3735);
or U5347 (N_5347,N_4953,N_4688);
nor U5348 (N_5348,N_157,N_4038);
or U5349 (N_5349,N_1976,N_661);
or U5350 (N_5350,N_4191,N_3427);
and U5351 (N_5351,N_2800,N_3350);
nor U5352 (N_5352,N_1965,N_4182);
nand U5353 (N_5353,N_998,N_4087);
and U5354 (N_5354,N_2348,N_1515);
nand U5355 (N_5355,N_4023,N_1785);
and U5356 (N_5356,N_991,N_2507);
xor U5357 (N_5357,N_3218,N_2926);
nand U5358 (N_5358,N_441,N_2316);
nor U5359 (N_5359,N_2551,N_3842);
or U5360 (N_5360,N_3768,N_598);
and U5361 (N_5361,N_2782,N_3410);
nor U5362 (N_5362,N_4017,N_2654);
xnor U5363 (N_5363,N_294,N_1005);
or U5364 (N_5364,N_3560,N_469);
xor U5365 (N_5365,N_2874,N_3149);
and U5366 (N_5366,N_2434,N_4124);
nor U5367 (N_5367,N_981,N_21);
nor U5368 (N_5368,N_877,N_4927);
or U5369 (N_5369,N_1192,N_1251);
or U5370 (N_5370,N_3280,N_3988);
and U5371 (N_5371,N_2668,N_1018);
nor U5372 (N_5372,N_4672,N_961);
nor U5373 (N_5373,N_4397,N_848);
nand U5374 (N_5374,N_286,N_1531);
nand U5375 (N_5375,N_4668,N_3321);
xor U5376 (N_5376,N_4006,N_3173);
and U5377 (N_5377,N_1559,N_4980);
nor U5378 (N_5378,N_2265,N_125);
xor U5379 (N_5379,N_3316,N_3345);
and U5380 (N_5380,N_2557,N_2511);
and U5381 (N_5381,N_4229,N_2699);
nor U5382 (N_5382,N_628,N_1492);
nand U5383 (N_5383,N_1124,N_514);
and U5384 (N_5384,N_2345,N_2695);
nor U5385 (N_5385,N_2056,N_429);
xnor U5386 (N_5386,N_4100,N_523);
xor U5387 (N_5387,N_4928,N_4352);
nor U5388 (N_5388,N_4030,N_658);
xor U5389 (N_5389,N_3279,N_4842);
nand U5390 (N_5390,N_2830,N_2747);
and U5391 (N_5391,N_1292,N_1794);
and U5392 (N_5392,N_1176,N_260);
and U5393 (N_5393,N_3040,N_3237);
xor U5394 (N_5394,N_3391,N_903);
or U5395 (N_5395,N_1110,N_3860);
nand U5396 (N_5396,N_1926,N_4748);
and U5397 (N_5397,N_4813,N_1892);
and U5398 (N_5398,N_3071,N_811);
or U5399 (N_5399,N_1939,N_336);
or U5400 (N_5400,N_3602,N_4608);
and U5401 (N_5401,N_1912,N_2563);
and U5402 (N_5402,N_1444,N_1582);
nor U5403 (N_5403,N_3576,N_1053);
nor U5404 (N_5404,N_1954,N_2567);
nor U5405 (N_5405,N_993,N_3035);
xor U5406 (N_5406,N_780,N_0);
and U5407 (N_5407,N_2575,N_3680);
nand U5408 (N_5408,N_4299,N_917);
or U5409 (N_5409,N_4354,N_4236);
nor U5410 (N_5410,N_173,N_1749);
or U5411 (N_5411,N_3766,N_1195);
nand U5412 (N_5412,N_860,N_4711);
nor U5413 (N_5413,N_150,N_4846);
and U5414 (N_5414,N_1323,N_2924);
xor U5415 (N_5415,N_3389,N_1750);
or U5416 (N_5416,N_4771,N_2792);
xor U5417 (N_5417,N_630,N_2527);
nor U5418 (N_5418,N_2703,N_3287);
xnor U5419 (N_5419,N_415,N_3940);
and U5420 (N_5420,N_4202,N_4984);
xnor U5421 (N_5421,N_1152,N_201);
or U5422 (N_5422,N_2532,N_2451);
nand U5423 (N_5423,N_4455,N_1960);
nand U5424 (N_5424,N_322,N_3466);
xnor U5425 (N_5425,N_4315,N_4443);
and U5426 (N_5426,N_4127,N_4021);
and U5427 (N_5427,N_2176,N_3335);
or U5428 (N_5428,N_3798,N_4558);
or U5429 (N_5429,N_4142,N_3112);
xnor U5430 (N_5430,N_4561,N_4157);
nand U5431 (N_5431,N_2424,N_1600);
xor U5432 (N_5432,N_4200,N_1373);
nand U5433 (N_5433,N_3404,N_3729);
or U5434 (N_5434,N_4674,N_4062);
or U5435 (N_5435,N_3814,N_706);
xor U5436 (N_5436,N_3669,N_4401);
and U5437 (N_5437,N_4390,N_3208);
nor U5438 (N_5438,N_828,N_4722);
nor U5439 (N_5439,N_3853,N_2351);
xor U5440 (N_5440,N_384,N_1472);
or U5441 (N_5441,N_4116,N_725);
nand U5442 (N_5442,N_2292,N_1813);
nand U5443 (N_5443,N_139,N_4707);
and U5444 (N_5444,N_4689,N_4186);
or U5445 (N_5445,N_1834,N_1806);
or U5446 (N_5446,N_1800,N_3312);
nor U5447 (N_5447,N_1386,N_750);
xor U5448 (N_5448,N_4836,N_3348);
nand U5449 (N_5449,N_1333,N_398);
nand U5450 (N_5450,N_3009,N_3406);
xor U5451 (N_5451,N_393,N_3152);
or U5452 (N_5452,N_3695,N_3657);
and U5453 (N_5453,N_3726,N_1990);
nor U5454 (N_5454,N_716,N_270);
nor U5455 (N_5455,N_786,N_2039);
and U5456 (N_5456,N_4067,N_4795);
and U5457 (N_5457,N_236,N_4651);
nand U5458 (N_5458,N_3460,N_1724);
nand U5459 (N_5459,N_611,N_521);
xnor U5460 (N_5460,N_2965,N_1657);
nor U5461 (N_5461,N_1761,N_3962);
nor U5462 (N_5462,N_4776,N_2515);
xnor U5463 (N_5463,N_1869,N_153);
xor U5464 (N_5464,N_3545,N_4978);
and U5465 (N_5465,N_488,N_538);
nor U5466 (N_5466,N_1408,N_4469);
xor U5467 (N_5467,N_3166,N_3245);
or U5468 (N_5468,N_3626,N_4472);
or U5469 (N_5469,N_1179,N_4346);
or U5470 (N_5470,N_1718,N_483);
and U5471 (N_5471,N_47,N_3267);
or U5472 (N_5472,N_618,N_42);
or U5473 (N_5473,N_3196,N_3643);
nor U5474 (N_5474,N_3568,N_1883);
or U5475 (N_5475,N_3844,N_3228);
and U5476 (N_5476,N_767,N_799);
xnor U5477 (N_5477,N_2794,N_688);
and U5478 (N_5478,N_1236,N_685);
and U5479 (N_5479,N_1823,N_2871);
xor U5480 (N_5480,N_1348,N_3036);
xor U5481 (N_5481,N_2781,N_4717);
and U5482 (N_5482,N_3539,N_4173);
and U5483 (N_5483,N_1173,N_117);
xnor U5484 (N_5484,N_2394,N_4033);
nand U5485 (N_5485,N_3262,N_4305);
nand U5486 (N_5486,N_2246,N_4012);
nor U5487 (N_5487,N_3450,N_4951);
nor U5488 (N_5488,N_3302,N_1896);
nor U5489 (N_5489,N_3066,N_2649);
and U5490 (N_5490,N_4695,N_4356);
nor U5491 (N_5491,N_771,N_379);
and U5492 (N_5492,N_4014,N_4158);
nor U5493 (N_5493,N_2194,N_3231);
and U5494 (N_5494,N_4576,N_208);
and U5495 (N_5495,N_4649,N_3915);
xnor U5496 (N_5496,N_1491,N_2574);
nand U5497 (N_5497,N_1359,N_4297);
and U5498 (N_5498,N_315,N_3277);
nand U5499 (N_5499,N_1662,N_4788);
nand U5500 (N_5500,N_4456,N_81);
or U5501 (N_5501,N_2329,N_2274);
and U5502 (N_5502,N_515,N_4607);
xor U5503 (N_5503,N_88,N_44);
xor U5504 (N_5504,N_588,N_3595);
or U5505 (N_5505,N_1494,N_2350);
and U5506 (N_5506,N_3718,N_3575);
xor U5507 (N_5507,N_500,N_4278);
xor U5508 (N_5508,N_3047,N_637);
nand U5509 (N_5509,N_4629,N_2491);
nor U5510 (N_5510,N_4408,N_2560);
nor U5511 (N_5511,N_3953,N_3025);
xnor U5512 (N_5512,N_4015,N_38);
nand U5513 (N_5513,N_2325,N_4242);
or U5514 (N_5514,N_3122,N_4744);
nand U5515 (N_5515,N_644,N_3999);
and U5516 (N_5516,N_4270,N_2608);
or U5517 (N_5517,N_843,N_2638);
and U5518 (N_5518,N_3346,N_2271);
or U5519 (N_5519,N_614,N_1530);
nand U5520 (N_5520,N_4389,N_4730);
and U5521 (N_5521,N_285,N_2701);
nand U5522 (N_5522,N_2206,N_3187);
xnor U5523 (N_5523,N_2183,N_516);
and U5524 (N_5524,N_3508,N_530);
and U5525 (N_5525,N_2379,N_1544);
nor U5526 (N_5526,N_4102,N_2028);
nor U5527 (N_5527,N_4780,N_1162);
or U5528 (N_5528,N_3476,N_3170);
nand U5529 (N_5529,N_3554,N_405);
or U5530 (N_5530,N_2041,N_2011);
nand U5531 (N_5531,N_1228,N_4739);
and U5532 (N_5532,N_3361,N_1983);
and U5533 (N_5533,N_2779,N_2650);
and U5534 (N_5534,N_2397,N_3524);
nor U5535 (N_5535,N_1308,N_3418);
or U5536 (N_5536,N_4805,N_4736);
and U5537 (N_5537,N_513,N_231);
xor U5538 (N_5538,N_1147,N_1332);
and U5539 (N_5539,N_3195,N_2733);
nand U5540 (N_5540,N_2360,N_701);
nor U5541 (N_5541,N_3273,N_2015);
or U5542 (N_5542,N_1760,N_1768);
or U5543 (N_5543,N_1671,N_2863);
nor U5544 (N_5544,N_3771,N_4701);
nand U5545 (N_5545,N_4291,N_3674);
or U5546 (N_5546,N_397,N_2180);
or U5547 (N_5547,N_337,N_4473);
and U5548 (N_5548,N_4276,N_970);
nor U5549 (N_5549,N_4634,N_3870);
nand U5550 (N_5550,N_4451,N_4218);
nor U5551 (N_5551,N_3561,N_1720);
xor U5552 (N_5552,N_4902,N_3687);
xnor U5553 (N_5553,N_152,N_1092);
xor U5554 (N_5554,N_299,N_3320);
or U5555 (N_5555,N_3630,N_4749);
nand U5556 (N_5556,N_1772,N_2356);
xnor U5557 (N_5557,N_4187,N_4865);
or U5558 (N_5558,N_4422,N_2807);
or U5559 (N_5559,N_4411,N_1217);
and U5560 (N_5560,N_3456,N_2097);
and U5561 (N_5561,N_1263,N_3207);
and U5562 (N_5562,N_1076,N_2837);
nor U5563 (N_5563,N_3487,N_3134);
nor U5564 (N_5564,N_2198,N_4714);
and U5565 (N_5565,N_2199,N_3801);
or U5566 (N_5566,N_3793,N_3271);
xnor U5567 (N_5567,N_2396,N_1738);
and U5568 (N_5568,N_652,N_266);
or U5569 (N_5569,N_4822,N_3479);
or U5570 (N_5570,N_1666,N_2134);
and U5571 (N_5571,N_2805,N_4904);
or U5572 (N_5572,N_2999,N_2003);
nand U5573 (N_5573,N_1403,N_2878);
and U5574 (N_5574,N_3433,N_3243);
xor U5575 (N_5575,N_560,N_3783);
nand U5576 (N_5576,N_522,N_1271);
nor U5577 (N_5577,N_4918,N_4706);
xnor U5578 (N_5578,N_2812,N_3774);
or U5579 (N_5579,N_3054,N_850);
nand U5580 (N_5580,N_4437,N_1961);
nand U5581 (N_5581,N_4107,N_2122);
nand U5582 (N_5582,N_226,N_1942);
nand U5583 (N_5583,N_3486,N_354);
xnor U5584 (N_5584,N_3172,N_1498);
and U5585 (N_5585,N_824,N_2982);
and U5586 (N_5586,N_2963,N_567);
nand U5587 (N_5587,N_3610,N_4153);
xor U5588 (N_5588,N_4535,N_462);
nor U5589 (N_5589,N_1506,N_1247);
nand U5590 (N_5590,N_4144,N_3949);
xnor U5591 (N_5591,N_1396,N_1169);
xor U5592 (N_5592,N_3446,N_2763);
nor U5593 (N_5593,N_4942,N_641);
nand U5594 (N_5594,N_4814,N_427);
nand U5595 (N_5595,N_2256,N_535);
nand U5596 (N_5596,N_859,N_2868);
and U5597 (N_5597,N_3168,N_1680);
xnor U5598 (N_5598,N_2392,N_916);
and U5599 (N_5599,N_268,N_1919);
and U5600 (N_5600,N_1822,N_3260);
xnor U5601 (N_5601,N_1009,N_1681);
xnor U5602 (N_5602,N_1024,N_4384);
nand U5603 (N_5603,N_61,N_1946);
and U5604 (N_5604,N_2027,N_349);
nand U5605 (N_5605,N_1889,N_4696);
xnor U5606 (N_5606,N_656,N_3889);
or U5607 (N_5607,N_2283,N_1501);
or U5608 (N_5608,N_3809,N_4857);
xor U5609 (N_5609,N_101,N_4475);
nand U5610 (N_5610,N_505,N_3341);
nand U5611 (N_5611,N_2179,N_2107);
nor U5612 (N_5612,N_4429,N_1304);
and U5613 (N_5613,N_4059,N_3178);
xor U5614 (N_5614,N_165,N_631);
xnor U5615 (N_5615,N_2637,N_4586);
nor U5616 (N_5616,N_2849,N_3197);
xnor U5617 (N_5617,N_4199,N_3850);
nor U5618 (N_5618,N_3387,N_4492);
xnor U5619 (N_5619,N_1495,N_2071);
and U5620 (N_5620,N_4666,N_391);
and U5621 (N_5621,N_75,N_1283);
nand U5622 (N_5622,N_3018,N_287);
nor U5623 (N_5623,N_4151,N_2113);
and U5624 (N_5624,N_1784,N_3960);
nand U5625 (N_5625,N_1572,N_1134);
nand U5626 (N_5626,N_4234,N_3162);
nand U5627 (N_5627,N_1968,N_1112);
and U5628 (N_5628,N_2968,N_470);
xnor U5629 (N_5629,N_4724,N_622);
nand U5630 (N_5630,N_973,N_2721);
or U5631 (N_5631,N_1331,N_3761);
and U5632 (N_5632,N_2493,N_1268);
xnor U5633 (N_5633,N_1780,N_775);
and U5634 (N_5634,N_1609,N_4099);
or U5635 (N_5635,N_4719,N_19);
nor U5636 (N_5636,N_50,N_3485);
nor U5637 (N_5637,N_137,N_971);
xor U5638 (N_5638,N_3217,N_1921);
and U5639 (N_5639,N_3494,N_4369);
or U5640 (N_5640,N_1712,N_4497);
nor U5641 (N_5641,N_2051,N_4332);
or U5642 (N_5642,N_57,N_1413);
nand U5643 (N_5643,N_566,N_1622);
and U5644 (N_5644,N_1792,N_2581);
nand U5645 (N_5645,N_3156,N_3070);
and U5646 (N_5646,N_80,N_504);
and U5647 (N_5647,N_2299,N_2433);
xor U5648 (N_5648,N_3519,N_2835);
nand U5649 (N_5649,N_1555,N_3656);
and U5650 (N_5650,N_677,N_2712);
nand U5651 (N_5651,N_2617,N_3795);
nor U5652 (N_5652,N_3917,N_115);
and U5653 (N_5653,N_1863,N_1161);
nor U5654 (N_5654,N_4716,N_1419);
nand U5655 (N_5655,N_4360,N_3412);
nor U5656 (N_5656,N_1755,N_2941);
nand U5657 (N_5657,N_2979,N_1432);
nor U5658 (N_5658,N_1679,N_909);
xnor U5659 (N_5659,N_1502,N_528);
xor U5660 (N_5660,N_70,N_3747);
and U5661 (N_5661,N_4269,N_3401);
and U5662 (N_5662,N_252,N_2182);
xnor U5663 (N_5663,N_4029,N_4945);
xnor U5664 (N_5664,N_3086,N_1624);
or U5665 (N_5665,N_4961,N_3579);
or U5666 (N_5666,N_881,N_3691);
and U5667 (N_5667,N_1708,N_2459);
nand U5668 (N_5668,N_819,N_2372);
or U5669 (N_5669,N_1223,N_4398);
nand U5670 (N_5670,N_3694,N_872);
or U5671 (N_5671,N_2972,N_4374);
and U5672 (N_5672,N_965,N_829);
xor U5673 (N_5673,N_3242,N_432);
nor U5674 (N_5674,N_3491,N_3004);
and U5675 (N_5675,N_3587,N_4962);
and U5676 (N_5676,N_2300,N_1135);
nor U5677 (N_5677,N_4680,N_737);
nand U5678 (N_5678,N_894,N_2);
or U5679 (N_5679,N_2204,N_3283);
or U5680 (N_5680,N_234,N_3257);
or U5681 (N_5681,N_913,N_3343);
and U5682 (N_5682,N_2784,N_818);
nor U5683 (N_5683,N_4453,N_2804);
nand U5684 (N_5684,N_1668,N_620);
xor U5685 (N_5685,N_2002,N_2090);
or U5686 (N_5686,N_3882,N_1994);
and U5687 (N_5687,N_4139,N_3351);
xnor U5688 (N_5688,N_3206,N_1418);
or U5689 (N_5689,N_4306,N_2099);
nand U5690 (N_5690,N_1897,N_4167);
nor U5691 (N_5691,N_320,N_1325);
and U5692 (N_5692,N_4890,N_3843);
xnor U5693 (N_5693,N_2173,N_132);
nand U5694 (N_5694,N_2673,N_1014);
xnor U5695 (N_5695,N_3806,N_2055);
nor U5696 (N_5696,N_3468,N_60);
xnor U5697 (N_5697,N_1576,N_1804);
nand U5698 (N_5698,N_2450,N_4937);
nor U5699 (N_5699,N_2544,N_3829);
or U5700 (N_5700,N_2309,N_2436);
nand U5701 (N_5701,N_4131,N_4697);
or U5702 (N_5702,N_3416,N_3308);
and U5703 (N_5703,N_2368,N_1278);
nor U5704 (N_5704,N_1428,N_754);
nand U5705 (N_5705,N_366,N_4893);
or U5706 (N_5706,N_1026,N_94);
nor U5707 (N_5707,N_957,N_4114);
xor U5708 (N_5708,N_3420,N_3226);
xnor U5709 (N_5709,N_2036,N_3926);
xnor U5710 (N_5710,N_3142,N_3250);
xnor U5711 (N_5711,N_1131,N_3530);
or U5712 (N_5712,N_3421,N_3705);
nor U5713 (N_5713,N_2234,N_230);
or U5714 (N_5714,N_4767,N_1095);
xnor U5715 (N_5715,N_4597,N_1496);
or U5716 (N_5716,N_4905,N_4511);
or U5717 (N_5717,N_4393,N_2796);
and U5718 (N_5718,N_1781,N_465);
xor U5719 (N_5719,N_98,N_1216);
nand U5720 (N_5720,N_428,N_4223);
or U5721 (N_5721,N_13,N_2958);
and U5722 (N_5722,N_264,N_3833);
xor U5723 (N_5723,N_2583,N_3087);
or U5724 (N_5724,N_847,N_1819);
or U5725 (N_5725,N_4350,N_3816);
xor U5726 (N_5726,N_3,N_1187);
nand U5727 (N_5727,N_679,N_2488);
nor U5728 (N_5728,N_918,N_2839);
nand U5729 (N_5729,N_3229,N_1918);
xor U5730 (N_5730,N_942,N_912);
xnor U5731 (N_5731,N_1035,N_2074);
xor U5732 (N_5732,N_657,N_1797);
nand U5733 (N_5733,N_3110,N_1739);
nor U5734 (N_5734,N_2139,N_4930);
xor U5735 (N_5735,N_1208,N_4690);
xor U5736 (N_5736,N_4407,N_4125);
xnor U5737 (N_5737,N_280,N_3884);
xor U5738 (N_5738,N_30,N_1069);
xnor U5739 (N_5739,N_1330,N_2985);
xor U5740 (N_5740,N_1605,N_4321);
nor U5741 (N_5741,N_1604,N_3264);
nand U5742 (N_5742,N_2319,N_4564);
nor U5743 (N_5743,N_3139,N_72);
or U5744 (N_5744,N_1928,N_2882);
nor U5745 (N_5745,N_732,N_2908);
xor U5746 (N_5746,N_4995,N_3616);
nor U5747 (N_5747,N_3596,N_3322);
and U5748 (N_5748,N_4869,N_2217);
xor U5749 (N_5749,N_2605,N_3764);
and U5750 (N_5750,N_1803,N_2059);
xnor U5751 (N_5751,N_3859,N_301);
xnor U5752 (N_5752,N_3093,N_587);
and U5753 (N_5753,N_3862,N_187);
nor U5754 (N_5754,N_3221,N_633);
and U5755 (N_5755,N_2321,N_4406);
nor U5756 (N_5756,N_2043,N_2471);
and U5757 (N_5757,N_4755,N_4120);
nor U5758 (N_5758,N_2255,N_2940);
xor U5759 (N_5759,N_3659,N_2786);
and U5760 (N_5760,N_3836,N_291);
and U5761 (N_5761,N_1039,N_4434);
or U5762 (N_5762,N_4510,N_2473);
nor U5763 (N_5763,N_2714,N_251);
or U5764 (N_5764,N_1091,N_1795);
xor U5765 (N_5765,N_339,N_781);
xor U5766 (N_5766,N_3682,N_4481);
nor U5767 (N_5767,N_3863,N_3325);
nand U5768 (N_5768,N_3582,N_2165);
and U5769 (N_5769,N_1229,N_4261);
and U5770 (N_5770,N_2146,N_1050);
xnor U5771 (N_5771,N_1453,N_1703);
xnor U5772 (N_5772,N_305,N_2909);
or U5773 (N_5773,N_3902,N_1701);
or U5774 (N_5774,N_4165,N_3147);
xor U5775 (N_5775,N_4357,N_2505);
nand U5776 (N_5776,N_2380,N_3437);
nor U5777 (N_5777,N_3301,N_2089);
and U5778 (N_5778,N_1378,N_3538);
or U5779 (N_5779,N_1935,N_3056);
xnor U5780 (N_5780,N_1546,N_4769);
or U5781 (N_5781,N_1101,N_1356);
xor U5782 (N_5782,N_1198,N_546);
or U5783 (N_5783,N_4212,N_2594);
and U5784 (N_5784,N_4194,N_3065);
or U5785 (N_5785,N_1473,N_645);
nand U5786 (N_5786,N_4958,N_2219);
nand U5787 (N_5787,N_2395,N_2426);
or U5788 (N_5788,N_922,N_1773);
or U5789 (N_5789,N_3807,N_1002);
and U5790 (N_5790,N_2983,N_2568);
or U5791 (N_5791,N_1636,N_4126);
or U5792 (N_5792,N_4447,N_1526);
nor U5793 (N_5793,N_2825,N_4074);
nand U5794 (N_5794,N_4003,N_803);
nand U5795 (N_5795,N_2876,N_1690);
nand U5796 (N_5796,N_2339,N_211);
nor U5797 (N_5797,N_1298,N_2386);
xnor U5798 (N_5798,N_1023,N_1274);
nor U5799 (N_5799,N_1119,N_1726);
and U5800 (N_5800,N_2376,N_1848);
or U5801 (N_5801,N_2656,N_3078);
and U5802 (N_5802,N_4111,N_1315);
xor U5803 (N_5803,N_1997,N_4924);
nand U5804 (N_5804,N_1455,N_3372);
or U5805 (N_5805,N_378,N_2956);
and U5806 (N_5806,N_1158,N_51);
nand U5807 (N_5807,N_341,N_2602);
nand U5808 (N_5808,N_1232,N_785);
xor U5809 (N_5809,N_297,N_755);
and U5810 (N_5810,N_2631,N_3749);
nor U5811 (N_5811,N_4880,N_3333);
nor U5812 (N_5812,N_166,N_4652);
or U5813 (N_5813,N_4154,N_512);
nand U5814 (N_5814,N_736,N_3615);
or U5815 (N_5815,N_4671,N_3002);
nor U5816 (N_5816,N_4515,N_1044);
and U5817 (N_5817,N_1102,N_2332);
nand U5818 (N_5818,N_1607,N_1993);
nand U5819 (N_5819,N_573,N_39);
nor U5820 (N_5820,N_1743,N_3818);
or U5821 (N_5821,N_1878,N_1266);
or U5822 (N_5822,N_3838,N_2753);
and U5823 (N_5823,N_1104,N_4851);
or U5824 (N_5824,N_2819,N_3383);
or U5825 (N_5825,N_2911,N_4046);
and U5826 (N_5826,N_2260,N_4987);
nor U5827 (N_5827,N_2307,N_179);
and U5828 (N_5828,N_2076,N_1249);
or U5829 (N_5829,N_4065,N_2900);
nor U5830 (N_5830,N_2774,N_1409);
and U5831 (N_5831,N_3557,N_1835);
nor U5832 (N_5832,N_2160,N_4513);
nor U5833 (N_5833,N_4156,N_1156);
xnor U5834 (N_5834,N_569,N_3246);
nor U5835 (N_5835,N_2946,N_327);
nand U5836 (N_5836,N_1038,N_2231);
nor U5837 (N_5837,N_4243,N_1185);
or U5838 (N_5838,N_2641,N_3115);
or U5839 (N_5839,N_3564,N_4343);
xor U5840 (N_5840,N_4495,N_930);
nand U5841 (N_5841,N_4143,N_1700);
and U5842 (N_5842,N_83,N_2528);
xnor U5843 (N_5843,N_2991,N_1401);
nand U5844 (N_5844,N_3664,N_1809);
nand U5845 (N_5845,N_2373,N_408);
or U5846 (N_5846,N_1805,N_4901);
or U5847 (N_5847,N_4002,N_67);
xor U5848 (N_5848,N_1390,N_1108);
or U5849 (N_5849,N_3558,N_4579);
and U5850 (N_5850,N_218,N_4066);
nor U5851 (N_5851,N_4727,N_4879);
xor U5852 (N_5852,N_4681,N_4590);
nor U5853 (N_5853,N_4840,N_4911);
and U5854 (N_5854,N_4631,N_104);
nand U5855 (N_5855,N_3145,N_689);
nand U5856 (N_5856,N_4728,N_4400);
nand U5857 (N_5857,N_3817,N_3980);
and U5858 (N_5858,N_4047,N_3282);
nand U5859 (N_5859,N_3238,N_1234);
and U5860 (N_5860,N_1599,N_4079);
nor U5861 (N_5861,N_3012,N_3594);
nor U5862 (N_5862,N_210,N_2681);
or U5863 (N_5863,N_4992,N_2790);
nand U5864 (N_5864,N_1380,N_4417);
and U5865 (N_5865,N_1684,N_884);
and U5866 (N_5866,N_2208,N_709);
and U5867 (N_5867,N_784,N_4022);
xor U5868 (N_5868,N_3360,N_2393);
nand U5869 (N_5869,N_2462,N_1876);
and U5870 (N_5870,N_1847,N_4906);
or U5871 (N_5871,N_213,N_1981);
nor U5872 (N_5872,N_4176,N_1820);
xor U5873 (N_5873,N_4965,N_796);
nor U5874 (N_5874,N_4514,N_4013);
xnor U5875 (N_5875,N_1193,N_1456);
nand U5876 (N_5876,N_2771,N_2203);
or U5877 (N_5877,N_3633,N_1788);
or U5878 (N_5878,N_1886,N_4643);
and U5879 (N_5879,N_4479,N_3971);
nor U5880 (N_5880,N_3309,N_1500);
nand U5881 (N_5881,N_4106,N_885);
nand U5882 (N_5882,N_2661,N_4391);
or U5883 (N_5883,N_790,N_3329);
xnor U5884 (N_5884,N_2181,N_406);
xnor U5885 (N_5885,N_1068,N_105);
nor U5886 (N_5886,N_2276,N_26);
and U5887 (N_5887,N_3827,N_4460);
xnor U5888 (N_5888,N_2288,N_896);
and U5889 (N_5889,N_4610,N_1089);
nand U5890 (N_5890,N_2364,N_4655);
xnor U5891 (N_5891,N_2419,N_1120);
or U5892 (N_5892,N_4878,N_3966);
nor U5893 (N_5893,N_3092,N_1757);
or U5894 (N_5894,N_3169,N_63);
nand U5895 (N_5895,N_3417,N_4091);
nand U5896 (N_5896,N_3876,N_629);
nor U5897 (N_5897,N_2966,N_3258);
nand U5898 (N_5898,N_243,N_4573);
or U5899 (N_5899,N_3547,N_2920);
and U5900 (N_5900,N_3090,N_2740);
and U5901 (N_5901,N_3213,N_1711);
or U5902 (N_5902,N_2865,N_148);
xnor U5903 (N_5903,N_3748,N_1745);
nor U5904 (N_5904,N_902,N_1256);
and U5905 (N_5905,N_3024,N_2391);
or U5906 (N_5906,N_2371,N_3812);
or U5907 (N_5907,N_1843,N_580);
nand U5908 (N_5908,N_1884,N_4439);
nor U5909 (N_5909,N_4008,N_4052);
and U5910 (N_5910,N_3369,N_4055);
xnor U5911 (N_5911,N_304,N_1071);
and U5912 (N_5912,N_3438,N_3703);
xor U5913 (N_5913,N_4997,N_2303);
or U5914 (N_5914,N_2171,N_978);
or U5915 (N_5915,N_1587,N_1482);
or U5916 (N_5916,N_2559,N_870);
xnor U5917 (N_5917,N_735,N_1618);
xor U5918 (N_5918,N_1166,N_188);
nand U5919 (N_5919,N_2472,N_3916);
or U5920 (N_5920,N_1900,N_4998);
or U5921 (N_5921,N_2150,N_1085);
and U5922 (N_5922,N_4338,N_2847);
nand U5923 (N_5923,N_2145,N_4347);
and U5924 (N_5924,N_3388,N_4578);
nor U5925 (N_5925,N_4232,N_4174);
xnor U5926 (N_5926,N_2857,N_615);
or U5927 (N_5927,N_2655,N_3678);
and U5928 (N_5928,N_2677,N_114);
nand U5929 (N_5929,N_4326,N_2682);
nor U5930 (N_5930,N_4541,N_3030);
nor U5931 (N_5931,N_1966,N_4068);
xor U5932 (N_5932,N_1702,N_4110);
nand U5933 (N_5933,N_746,N_3463);
and U5934 (N_5934,N_711,N_1318);
xor U5935 (N_5935,N_3534,N_4837);
and U5936 (N_5936,N_2530,N_308);
and U5937 (N_5937,N_203,N_2977);
or U5938 (N_5938,N_2104,N_3290);
nor U5939 (N_5939,N_3732,N_4899);
xnor U5940 (N_5940,N_4745,N_2466);
xor U5941 (N_5941,N_3136,N_2652);
and U5942 (N_5942,N_774,N_3268);
and U5943 (N_5943,N_262,N_2836);
or U5944 (N_5944,N_4656,N_865);
nand U5945 (N_5945,N_2663,N_4378);
and U5946 (N_5946,N_4622,N_2420);
or U5947 (N_5947,N_1279,N_2531);
or U5948 (N_5948,N_492,N_1617);
and U5949 (N_5949,N_4877,N_3001);
or U5950 (N_5950,N_1282,N_1592);
or U5951 (N_5951,N_306,N_1901);
xnor U5952 (N_5952,N_4663,N_3866);
and U5953 (N_5953,N_3010,N_3994);
nor U5954 (N_5954,N_457,N_1436);
xor U5955 (N_5955,N_2435,N_1995);
or U5956 (N_5956,N_2168,N_842);
nor U5957 (N_5957,N_4555,N_4316);
nand U5958 (N_5958,N_4800,N_3868);
nand U5959 (N_5959,N_2035,N_3567);
nand U5960 (N_5960,N_261,N_3731);
nor U5961 (N_5961,N_778,N_4433);
and U5962 (N_5962,N_3992,N_2590);
nor U5963 (N_5963,N_3034,N_3255);
nand U5964 (N_5964,N_3708,N_1037);
nand U5965 (N_5965,N_3702,N_1637);
and U5966 (N_5966,N_2713,N_3191);
nor U5967 (N_5967,N_1137,N_4123);
xnor U5968 (N_5968,N_809,N_2945);
and U5969 (N_5969,N_2533,N_723);
nor U5970 (N_5970,N_3650,N_1669);
or U5971 (N_5971,N_3439,N_1242);
nand U5972 (N_5972,N_3165,N_550);
xnor U5973 (N_5973,N_3919,N_2915);
or U5974 (N_5974,N_3481,N_2791);
xor U5975 (N_5975,N_2352,N_4894);
or U5976 (N_5976,N_6,N_3826);
xnor U5977 (N_5977,N_2192,N_4604);
or U5978 (N_5978,N_4485,N_749);
or U5979 (N_5979,N_2636,N_3215);
and U5980 (N_5980,N_517,N_2642);
xnor U5981 (N_5981,N_3051,N_1593);
and U5982 (N_5982,N_2163,N_3318);
or U5983 (N_5983,N_2750,N_2534);
nor U5984 (N_5984,N_2026,N_1412);
or U5985 (N_5985,N_3622,N_3529);
and U5986 (N_5986,N_4841,N_702);
nand U5987 (N_5987,N_1882,N_4859);
nor U5988 (N_5988,N_3845,N_2828);
or U5989 (N_5989,N_1938,N_273);
or U5990 (N_5990,N_926,N_1846);
or U5991 (N_5991,N_2347,N_1875);
xnor U5992 (N_5992,N_835,N_4919);
and U5993 (N_5993,N_1029,N_11);
or U5994 (N_5994,N_4088,N_4952);
xnor U5995 (N_5995,N_714,N_2957);
nand U5996 (N_5996,N_760,N_3205);
or U5997 (N_5997,N_2024,N_4294);
xnor U5998 (N_5998,N_2040,N_3824);
nor U5999 (N_5999,N_1377,N_403);
or U6000 (N_6000,N_3328,N_707);
and U6001 (N_6001,N_183,N_2662);
and U6002 (N_6002,N_1561,N_4348);
nor U6003 (N_6003,N_914,N_1159);
and U6004 (N_6004,N_4895,N_3174);
xor U6005 (N_6005,N_1638,N_3652);
or U6006 (N_6006,N_4527,N_4897);
xor U6007 (N_6007,N_3640,N_3744);
nand U6008 (N_6008,N_1751,N_27);
nand U6009 (N_6009,N_164,N_4265);
nand U6010 (N_6010,N_205,N_1335);
xnor U6011 (N_6011,N_542,N_1598);
and U6012 (N_6012,N_1602,N_4613);
xor U6013 (N_6013,N_1728,N_3822);
xnor U6014 (N_6014,N_2912,N_3323);
or U6015 (N_6015,N_1209,N_174);
and U6016 (N_6016,N_3375,N_2538);
nand U6017 (N_6017,N_1929,N_58);
xnor U6018 (N_6018,N_2418,N_2981);
and U6019 (N_6019,N_3382,N_2761);
nor U6020 (N_6020,N_4602,N_794);
nand U6021 (N_6021,N_4589,N_3803);
nor U6022 (N_6022,N_2783,N_4912);
or U6023 (N_6023,N_4239,N_4458);
nor U6024 (N_6024,N_663,N_3796);
nor U6025 (N_6025,N_3483,N_4056);
xnor U6026 (N_6026,N_1967,N_3978);
nor U6027 (N_6027,N_3097,N_667);
and U6028 (N_6028,N_1885,N_1756);
nor U6029 (N_6029,N_4092,N_4830);
nand U6030 (N_6030,N_4596,N_607);
xor U6031 (N_6031,N_1518,N_1016);
and U6032 (N_6032,N_1574,N_3039);
nor U6033 (N_6033,N_2413,N_1086);
or U6034 (N_6034,N_3077,N_4164);
nor U6035 (N_6035,N_3864,N_3423);
and U6036 (N_6036,N_4898,N_3540);
or U6037 (N_6037,N_4379,N_3500);
and U6038 (N_6038,N_2363,N_3052);
and U6039 (N_6039,N_2322,N_682);
nor U6040 (N_6040,N_3805,N_1450);
xor U6041 (N_6041,N_4799,N_2667);
nand U6042 (N_6042,N_2341,N_670);
nor U6043 (N_6043,N_687,N_1285);
nor U6044 (N_6044,N_1917,N_249);
xnor U6045 (N_6045,N_582,N_577);
xnor U6046 (N_6046,N_290,N_3293);
nand U6047 (N_6047,N_4170,N_1143);
or U6048 (N_6048,N_1509,N_4635);
nor U6049 (N_6049,N_2902,N_1493);
or U6050 (N_6050,N_875,N_1894);
xnor U6051 (N_6051,N_4644,N_1270);
and U6052 (N_6052,N_2320,N_1769);
nand U6053 (N_6053,N_168,N_4687);
or U6054 (N_6054,N_272,N_1034);
or U6055 (N_6055,N_1689,N_4450);
nand U6056 (N_6056,N_375,N_1590);
nor U6057 (N_6057,N_4870,N_4349);
or U6058 (N_6058,N_3542,N_935);
or U6059 (N_6059,N_2153,N_3851);
nand U6060 (N_6060,N_974,N_906);
and U6061 (N_6061,N_3082,N_248);
and U6062 (N_6062,N_733,N_2017);
nand U6063 (N_6063,N_867,N_364);
or U6064 (N_6064,N_1048,N_4563);
nor U6065 (N_6065,N_3288,N_2685);
nor U6066 (N_6066,N_1317,N_2151);
nor U6067 (N_6067,N_269,N_129);
xor U6068 (N_6068,N_713,N_3811);
xnor U6069 (N_6069,N_2133,N_4274);
xnor U6070 (N_6070,N_2494,N_3154);
xnor U6071 (N_6071,N_4284,N_4351);
and U6072 (N_6072,N_3475,N_2044);
and U6073 (N_6073,N_2975,N_3760);
and U6074 (N_6074,N_4320,N_1296);
or U6075 (N_6075,N_4936,N_4119);
nand U6076 (N_6076,N_1877,N_1614);
xor U6077 (N_6077,N_490,N_2284);
and U6078 (N_6078,N_3194,N_4557);
and U6079 (N_6079,N_2358,N_46);
and U6080 (N_6080,N_4290,N_1814);
nand U6081 (N_6081,N_2399,N_4075);
nand U6082 (N_6082,N_1991,N_2092);
nor U6083 (N_6083,N_455,N_131);
and U6084 (N_6084,N_814,N_4874);
or U6085 (N_6085,N_2185,N_3364);
and U6086 (N_6086,N_1686,N_2293);
nand U6087 (N_6087,N_4983,N_557);
or U6088 (N_6088,N_4885,N_2599);
or U6089 (N_6089,N_2270,N_1475);
nor U6090 (N_6090,N_559,N_1425);
xnor U6091 (N_6091,N_2053,N_3848);
nor U6092 (N_6092,N_4442,N_1653);
nand U6093 (N_6093,N_2158,N_1293);
nand U6094 (N_6094,N_3544,N_4664);
nand U6095 (N_6095,N_2688,N_2881);
xnor U6096 (N_6096,N_394,N_293);
or U6097 (N_6097,N_2263,N_1294);
and U6098 (N_6098,N_4220,N_3471);
and U6099 (N_6099,N_552,N_932);
nand U6100 (N_6100,N_1844,N_4647);
or U6101 (N_6101,N_3908,N_946);
and U6102 (N_6102,N_1534,N_4792);
and U6103 (N_6103,N_4064,N_2359);
and U6104 (N_6104,N_3745,N_4947);
xor U6105 (N_6105,N_2078,N_4944);
or U6106 (N_6106,N_2135,N_2064);
and U6107 (N_6107,N_62,N_4364);
and U6108 (N_6108,N_920,N_3895);
xnor U6109 (N_6109,N_3928,N_3522);
nand U6110 (N_6110,N_547,N_1567);
nor U6111 (N_6111,N_2207,N_768);
xnor U6112 (N_6112,N_4794,N_4018);
nor U6113 (N_6113,N_1872,N_4373);
nor U6114 (N_6114,N_2477,N_4815);
or U6115 (N_6115,N_310,N_116);
or U6116 (N_6116,N_4889,N_2167);
and U6117 (N_6117,N_4549,N_3823);
nand U6118 (N_6118,N_3079,N_937);
nand U6119 (N_6119,N_350,N_2018);
or U6120 (N_6120,N_1569,N_3269);
or U6121 (N_6121,N_1366,N_3825);
nor U6122 (N_6122,N_4781,N_1164);
nand U6123 (N_6123,N_2159,N_4640);
nand U6124 (N_6124,N_2012,N_2994);
xor U6125 (N_6125,N_1827,N_571);
xnor U6126 (N_6126,N_363,N_2929);
nor U6127 (N_6127,N_438,N_2506);
nor U6128 (N_6128,N_192,N_855);
nor U6129 (N_6129,N_330,N_3942);
or U6130 (N_6130,N_868,N_721);
nor U6131 (N_6131,N_4611,N_4534);
and U6132 (N_6132,N_4914,N_1963);
and U6133 (N_6133,N_3204,N_1870);
or U6134 (N_6134,N_3645,N_185);
xor U6135 (N_6135,N_1888,N_177);
or U6136 (N_6136,N_4667,N_15);
xor U6137 (N_6137,N_1443,N_487);
xor U6138 (N_6138,N_3236,N_1153);
nand U6139 (N_6139,N_3501,N_1678);
xnor U6140 (N_6140,N_4181,N_2827);
or U6141 (N_6141,N_4041,N_1543);
nand U6142 (N_6142,N_2354,N_2866);
nand U6143 (N_6143,N_3160,N_4581);
or U6144 (N_6144,N_3455,N_1685);
nor U6145 (N_6145,N_4496,N_2928);
nor U6146 (N_6146,N_4552,N_155);
and U6147 (N_6147,N_1097,N_3453);
nand U6148 (N_6148,N_2240,N_4676);
nor U6149 (N_6149,N_217,N_4705);
xor U6150 (N_6150,N_389,N_2840);
xor U6151 (N_6151,N_1691,N_883);
nand U6152 (N_6152,N_4839,N_163);
nand U6153 (N_6153,N_335,N_2248);
nand U6154 (N_6154,N_4414,N_2903);
nand U6155 (N_6155,N_126,N_3937);
nand U6156 (N_6156,N_4855,N_3941);
and U6157 (N_6157,N_2047,N_2813);
or U6158 (N_6158,N_1654,N_1856);
nand U6159 (N_6159,N_1174,N_2894);
or U6160 (N_6160,N_2725,N_2442);
and U6161 (N_6161,N_1696,N_4026);
or U6162 (N_6162,N_1184,N_3489);
and U6163 (N_6163,N_2425,N_357);
or U6164 (N_6164,N_1324,N_2612);
or U6165 (N_6165,N_325,N_491);
nor U6166 (N_6166,N_2509,N_2174);
xnor U6167 (N_6167,N_2580,N_4028);
xor U6168 (N_6168,N_2546,N_4184);
and U6169 (N_6169,N_4208,N_1352);
or U6170 (N_6170,N_672,N_540);
and U6171 (N_6171,N_3620,N_1012);
nor U6172 (N_6172,N_4189,N_3901);
nand U6173 (N_6173,N_726,N_477);
or U6174 (N_6174,N_2556,N_1829);
xnor U6175 (N_6175,N_823,N_740);
and U6176 (N_6176,N_2697,N_450);
or U6177 (N_6177,N_3775,N_2769);
xnor U6178 (N_6178,N_4692,N_1340);
xnor U6179 (N_6179,N_3993,N_77);
or U6180 (N_6180,N_1956,N_2898);
or U6181 (N_6181,N_3304,N_1640);
or U6182 (N_6182,N_4289,N_3570);
or U6183 (N_6183,N_4977,N_2802);
xor U6184 (N_6184,N_836,N_2555);
and U6185 (N_6185,N_1213,N_4628);
and U6186 (N_6186,N_1125,N_1665);
xnor U6187 (N_6187,N_553,N_987);
and U6188 (N_6188,N_2184,N_1058);
nor U6189 (N_6189,N_3607,N_3985);
and U6190 (N_6190,N_3297,N_4569);
nor U6191 (N_6191,N_1499,N_1341);
xnor U6192 (N_6192,N_1239,N_2884);
xor U6193 (N_6193,N_2453,N_400);
or U6194 (N_6194,N_1527,N_4424);
or U6195 (N_6195,N_1461,N_501);
and U6196 (N_6196,N_4683,N_4025);
and U6197 (N_6197,N_3847,N_3060);
or U6198 (N_6198,N_3782,N_1336);
and U6199 (N_6199,N_2243,N_118);
xor U6200 (N_6200,N_3482,N_1953);
and U6201 (N_6201,N_1180,N_4854);
or U6202 (N_6202,N_3031,N_2357);
or U6203 (N_6203,N_244,N_2564);
or U6204 (N_6204,N_312,N_3064);
xnor U6205 (N_6205,N_2119,N_196);
and U6206 (N_6206,N_3970,N_3444);
or U6207 (N_6207,N_3449,N_1557);
or U6208 (N_6208,N_949,N_385);
nor U6209 (N_6209,N_3989,N_1437);
or U6210 (N_6210,N_2205,N_3084);
xor U6211 (N_6211,N_3124,N_1245);
nand U6212 (N_6212,N_1451,N_854);
xnor U6213 (N_6213,N_383,N_4135);
nand U6214 (N_6214,N_704,N_4773);
nand U6215 (N_6215,N_3074,N_3707);
nand U6216 (N_6216,N_3831,N_1284);
and U6217 (N_6217,N_3632,N_3344);
or U6218 (N_6218,N_4385,N_20);
and U6219 (N_6219,N_3219,N_4821);
nor U6220 (N_6220,N_1706,N_4856);
nor U6221 (N_6221,N_3712,N_3395);
and U6222 (N_6222,N_2843,N_4402);
nand U6223 (N_6223,N_2080,N_3858);
xor U6224 (N_6224,N_409,N_874);
nor U6225 (N_6225,N_1096,N_493);
nand U6226 (N_6226,N_3767,N_1621);
nand U6227 (N_6227,N_4503,N_1774);
nor U6228 (N_6228,N_1710,N_3029);
xor U6229 (N_6229,N_1463,N_1947);
xnor U6230 (N_6230,N_3424,N_2417);
nand U6231 (N_6231,N_1230,N_3923);
and U6232 (N_6232,N_984,N_4766);
nand U6233 (N_6233,N_370,N_143);
nor U6234 (N_6234,N_4095,N_4617);
and U6235 (N_6235,N_2415,N_2626);
nor U6236 (N_6236,N_4036,N_804);
nand U6237 (N_6237,N_4844,N_1791);
xnor U6238 (N_6238,N_3877,N_4509);
and U6239 (N_6239,N_3757,N_2091);
xnor U6240 (N_6240,N_3063,N_3921);
or U6241 (N_6241,N_1150,N_3314);
or U6242 (N_6242,N_2072,N_2918);
xor U6243 (N_6243,N_3167,N_4638);
xnor U6244 (N_6244,N_56,N_1334);
nor U6245 (N_6245,N_2875,N_617);
or U6246 (N_6246,N_4105,N_581);
nor U6247 (N_6247,N_2743,N_3126);
xnor U6248 (N_6248,N_3464,N_3585);
nand U6249 (N_6249,N_3135,N_2582);
nand U6250 (N_6250,N_934,N_2432);
xor U6251 (N_6251,N_365,N_1191);
nor U6252 (N_6252,N_1370,N_1224);
nor U6253 (N_6253,N_3906,N_605);
or U6254 (N_6254,N_33,N_1295);
nand U6255 (N_6255,N_2456,N_323);
nand U6256 (N_6256,N_2954,N_2403);
or U6257 (N_6257,N_3274,N_4007);
nor U6258 (N_6258,N_3182,N_3381);
xnor U6259 (N_6259,N_3284,N_2022);
or U6260 (N_6260,N_3800,N_36);
nor U6261 (N_6261,N_3763,N_3100);
xnor U6262 (N_6262,N_3713,N_254);
nand U6263 (N_6263,N_4731,N_446);
and U6264 (N_6264,N_3349,N_3378);
nor U6265 (N_6265,N_1508,N_795);
nand U6266 (N_6266,N_3577,N_989);
xnor U6267 (N_6267,N_3770,N_4301);
and U6268 (N_6268,N_3119,N_1984);
nor U6269 (N_6269,N_453,N_4327);
nand U6270 (N_6270,N_3488,N_3613);
nor U6271 (N_6271,N_506,N_2959);
or U6272 (N_6272,N_4753,N_359);
nand U6273 (N_6273,N_29,N_151);
and U6274 (N_6274,N_4650,N_3185);
nor U6275 (N_6275,N_1389,N_4262);
nand U6276 (N_6276,N_2571,N_3184);
nand U6277 (N_6277,N_3549,N_3518);
nor U6278 (N_6278,N_1519,N_1328);
or U6279 (N_6279,N_2984,N_2689);
or U6280 (N_6280,N_4828,N_2416);
xor U6281 (N_6281,N_3601,N_3855);
or U6282 (N_6282,N_2268,N_2990);
nand U6283 (N_6283,N_1619,N_84);
nor U6284 (N_6284,N_4824,N_1729);
or U6285 (N_6285,N_4245,N_2821);
or U6286 (N_6286,N_507,N_4512);
nor U6287 (N_6287,N_4210,N_4355);
nand U6288 (N_6288,N_2370,N_4568);
nand U6289 (N_6289,N_3893,N_3875);
nand U6290 (N_6290,N_1481,N_3393);
nand U6291 (N_6291,N_648,N_2707);
and U6292 (N_6292,N_1077,N_1512);
or U6293 (N_6293,N_1949,N_2630);
nand U6294 (N_6294,N_710,N_2944);
nand U6295 (N_6295,N_2023,N_333);
nor U6296 (N_6296,N_1911,N_473);
nor U6297 (N_6297,N_4071,N_4659);
xor U6298 (N_6298,N_1351,N_1525);
or U6299 (N_6299,N_128,N_2856);
or U6300 (N_6300,N_3513,N_2501);
and U6301 (N_6301,N_2616,N_130);
and U6302 (N_6302,N_2342,N_2421);
nand U6303 (N_6303,N_4826,N_3983);
xor U6304 (N_6304,N_2323,N_1941);
xnor U6305 (N_6305,N_4872,N_1986);
nand U6306 (N_6306,N_4381,N_2123);
nor U6307 (N_6307,N_2969,N_4438);
xnor U6308 (N_6308,N_4871,N_4574);
nor U6309 (N_6309,N_3473,N_810);
xor U6310 (N_6310,N_2014,N_2213);
or U6311 (N_6311,N_220,N_2499);
and U6312 (N_6312,N_4522,N_382);
and U6313 (N_6313,N_3820,N_4335);
nand U6314 (N_6314,N_996,N_861);
nand U6315 (N_6315,N_3523,N_3617);
nor U6316 (N_6316,N_1231,N_2267);
and U6317 (N_6317,N_4775,N_3352);
or U6318 (N_6318,N_4285,N_3419);
and U6319 (N_6319,N_3532,N_592);
nand U6320 (N_6320,N_1873,N_4482);
and U6321 (N_6321,N_3357,N_3728);
xnor U6322 (N_6322,N_3614,N_4412);
nand U6323 (N_6323,N_995,N_531);
xnor U6324 (N_6324,N_4273,N_2896);
nor U6325 (N_6325,N_1346,N_2935);
xor U6326 (N_6326,N_2235,N_1054);
nand U6327 (N_6327,N_4876,N_953);
nand U6328 (N_6328,N_4113,N_3913);
nand U6329 (N_6329,N_2304,N_1218);
or U6330 (N_6330,N_4147,N_1758);
xor U6331 (N_6331,N_4933,N_4259);
and U6332 (N_6332,N_1007,N_2172);
nand U6333 (N_6333,N_1521,N_4192);
nor U6334 (N_6334,N_1431,N_3138);
xor U6335 (N_6335,N_2029,N_4253);
nand U6336 (N_6336,N_3337,N_4883);
and U6337 (N_6337,N_2921,N_2098);
nand U6338 (N_6338,N_1063,N_2562);
nand U6339 (N_6339,N_4867,N_32);
xor U6340 (N_6340,N_2540,N_2880);
nor U6341 (N_6341,N_3572,N_4910);
and U6342 (N_6342,N_4506,N_2337);
xor U6343 (N_6343,N_1849,N_787);
nor U6344 (N_6344,N_4037,N_2005);
nand U6345 (N_6345,N_2822,N_16);
or U6346 (N_6346,N_1717,N_2389);
nor U6347 (N_6347,N_3265,N_910);
and U6348 (N_6348,N_2033,N_4049);
nor U6349 (N_6349,N_960,N_3688);
nor U6350 (N_6350,N_966,N_3028);
and U6351 (N_6351,N_638,N_2561);
xnor U6352 (N_6352,N_2109,N_4950);
nor U6353 (N_6353,N_1003,N_816);
nand U6354 (N_6354,N_4507,N_1183);
nor U6355 (N_6355,N_1705,N_4177);
or U6356 (N_6356,N_2879,N_2643);
nand U6357 (N_6357,N_4193,N_1796);
or U6358 (N_6358,N_1601,N_4925);
and U6359 (N_6359,N_3430,N_2478);
nand U6360 (N_6360,N_3192,N_4741);
xor U6361 (N_6361,N_3804,N_2762);
nor U6362 (N_6362,N_2411,N_3397);
and U6363 (N_6363,N_1982,N_632);
or U6364 (N_6364,N_4531,N_1841);
xnor U6365 (N_6365,N_4939,N_3890);
nor U6366 (N_6366,N_2943,N_4283);
nand U6367 (N_6367,N_1719,N_209);
nor U6368 (N_6368,N_2591,N_4132);
or U6369 (N_6369,N_3900,N_866);
and U6370 (N_6370,N_4051,N_2193);
and U6371 (N_6371,N_1379,N_4708);
nor U6372 (N_6372,N_2620,N_411);
xor U6373 (N_6373,N_3888,N_1358);
nor U6374 (N_6374,N_968,N_1881);
nand U6375 (N_6375,N_2034,N_1047);
nor U6376 (N_6376,N_1082,N_1845);
xnor U6377 (N_6377,N_275,N_753);
nor U6378 (N_6378,N_4550,N_314);
nor U6379 (N_6379,N_3541,N_2085);
and U6380 (N_6380,N_807,N_4712);
xor U6381 (N_6381,N_3955,N_1652);
or U6382 (N_6382,N_1237,N_915);
xnor U6383 (N_6383,N_2214,N_2129);
xnor U6384 (N_6384,N_107,N_1275);
and U6385 (N_6385,N_2732,N_3434);
nand U6386 (N_6386,N_1775,N_2948);
or U6387 (N_6387,N_1196,N_3436);
and U6388 (N_6388,N_1059,N_539);
and U6389 (N_6389,N_1168,N_1355);
and U6390 (N_6390,N_3355,N_1633);
or U6391 (N_6391,N_2759,N_2238);
nor U6392 (N_6392,N_454,N_2008);
and U6393 (N_6393,N_1503,N_1766);
xor U6394 (N_6394,N_2269,N_1782);
xnor U6395 (N_6395,N_3377,N_2799);
or U6396 (N_6396,N_73,N_2273);
xnor U6397 (N_6397,N_4489,N_4525);
or U6398 (N_6398,N_1553,N_3636);
and U6399 (N_6399,N_3555,N_110);
or U6400 (N_6400,N_1342,N_2992);
xor U6401 (N_6401,N_3256,N_4303);
or U6402 (N_6402,N_2675,N_4875);
nand U6403 (N_6403,N_2524,N_1931);
nor U6404 (N_6404,N_4255,N_2987);
xor U6405 (N_6405,N_3597,N_1145);
nor U6406 (N_6406,N_2045,N_1094);
nor U6407 (N_6407,N_4211,N_3609);
nand U6408 (N_6408,N_3106,N_95);
nor U6409 (N_6409,N_3429,N_1629);
and U6410 (N_6410,N_2860,N_2423);
and U6411 (N_6411,N_1562,N_65);
nor U6412 (N_6412,N_3835,N_856);
xor U6413 (N_6413,N_2232,N_3259);
nor U6414 (N_6414,N_2690,N_3932);
xnor U6415 (N_6415,N_69,N_1583);
or U6416 (N_6416,N_770,N_1001);
and U6417 (N_6417,N_1513,N_122);
and U6418 (N_6418,N_4090,N_324);
nand U6419 (N_6419,N_1098,N_3272);
or U6420 (N_6420,N_7,N_4591);
or U6421 (N_6421,N_904,N_3667);
nor U6422 (N_6422,N_671,N_4827);
and U6423 (N_6423,N_4718,N_2449);
or U6424 (N_6424,N_2680,N_1753);
xnor U6425 (N_6425,N_1122,N_1246);
xnor U6426 (N_6426,N_1233,N_1977);
xor U6427 (N_6427,N_4570,N_3099);
nand U6428 (N_6428,N_3458,N_1859);
and U6429 (N_6429,N_2604,N_558);
and U6430 (N_6430,N_2826,N_574);
nand U6431 (N_6431,N_2930,N_1563);
xor U6432 (N_6432,N_1017,N_4060);
xnor U6433 (N_6433,N_4957,N_4614);
or U6434 (N_6434,N_4886,N_4169);
nor U6435 (N_6435,N_2727,N_4464);
nand U6436 (N_6436,N_730,N_1426);
nand U6437 (N_6437,N_3611,N_4168);
nor U6438 (N_6438,N_447,N_4793);
or U6439 (N_6439,N_1478,N_4226);
or U6440 (N_6440,N_748,N_1388);
xor U6441 (N_6441,N_2855,N_2823);
nor U6442 (N_6442,N_4454,N_2961);
and U6443 (N_6443,N_1510,N_458);
or U6444 (N_6444,N_3679,N_4490);
nor U6445 (N_6445,N_3177,N_4404);
nor U6446 (N_6446,N_639,N_919);
and U6447 (N_6447,N_3697,N_4868);
nor U6448 (N_6448,N_2497,N_3920);
xnor U6449 (N_6449,N_283,N_533);
nor U6450 (N_6450,N_2020,N_2585);
or U6451 (N_6451,N_4085,N_3303);
nand U6452 (N_6452,N_568,N_907);
or U6453 (N_6453,N_2385,N_692);
nand U6454 (N_6454,N_4096,N_4985);
nand U6455 (N_6455,N_4619,N_1253);
nor U6456 (N_6456,N_23,N_2646);
nor U6457 (N_6457,N_825,N_2310);
and U6458 (N_6458,N_3263,N_1474);
nor U6459 (N_6459,N_4461,N_4394);
nand U6460 (N_6460,N_4094,N_3785);
xnor U6461 (N_6461,N_1025,N_87);
nor U6462 (N_6462,N_4825,N_2475);
nor U6463 (N_6463,N_659,N_4544);
xor U6464 (N_6464,N_3311,N_4171);
nand U6465 (N_6465,N_4658,N_2254);
nand U6466 (N_6466,N_4832,N_4823);
nor U6467 (N_6467,N_2760,N_2869);
nor U6468 (N_6468,N_951,N_2084);
xor U6469 (N_6469,N_4476,N_1511);
and U6470 (N_6470,N_990,N_2817);
and U6471 (N_6471,N_2887,N_256);
and U6472 (N_6472,N_1262,N_1838);
xor U6473 (N_6473,N_3644,N_708);
and U6474 (N_6474,N_2407,N_2717);
and U6475 (N_6475,N_3362,N_1644);
nor U6476 (N_6476,N_2148,N_1046);
nand U6477 (N_6477,N_4967,N_2486);
and U6478 (N_6478,N_1136,N_4248);
or U6479 (N_6479,N_3598,N_2082);
nor U6480 (N_6480,N_2349,N_2295);
and U6481 (N_6481,N_1433,N_1485);
xor U6482 (N_6482,N_2031,N_2220);
and U6483 (N_6483,N_3951,N_2872);
nand U6484 (N_6484,N_812,N_2522);
nor U6485 (N_6485,N_684,N_3780);
xnor U6486 (N_6486,N_3754,N_4263);
nor U6487 (N_6487,N_4819,N_3681);
and U6488 (N_6488,N_2702,N_1030);
or U6489 (N_6489,N_2190,N_2110);
and U6490 (N_6490,N_2676,N_2888);
nor U6491 (N_6491,N_3067,N_1171);
and U6492 (N_6492,N_496,N_2917);
nand U6493 (N_6493,N_374,N_4946);
and U6494 (N_6494,N_2818,N_1469);
nand U6495 (N_6495,N_3756,N_4887);
or U6496 (N_6496,N_4529,N_4698);
xnor U6497 (N_6497,N_863,N_1793);
or U6498 (N_6498,N_4224,N_1200);
xnor U6499 (N_6499,N_4104,N_2787);
xnor U6500 (N_6500,N_1532,N_37);
and U6501 (N_6501,N_1280,N_3840);
and U6502 (N_6502,N_1363,N_2378);
nand U6503 (N_6503,N_1862,N_1309);
nand U6504 (N_6504,N_3581,N_232);
nand U6505 (N_6505,N_4743,N_3091);
or U6506 (N_6506,N_1631,N_791);
and U6507 (N_6507,N_1189,N_703);
and U6508 (N_6508,N_4909,N_2313);
nor U6509 (N_6509,N_3050,N_135);
nand U6510 (N_6510,N_2978,N_3927);
or U6511 (N_6511,N_1021,N_1060);
nand U6512 (N_6512,N_3107,N_2936);
or U6513 (N_6513,N_4520,N_1596);
nand U6514 (N_6514,N_4994,N_4341);
or U6515 (N_6515,N_697,N_3629);
xnor U6516 (N_6516,N_839,N_623);
and U6517 (N_6517,N_2279,N_1861);
or U6518 (N_6518,N_1817,N_368);
or U6519 (N_6519,N_4011,N_2460);
xnor U6520 (N_6520,N_1969,N_3211);
and U6521 (N_6521,N_3580,N_2729);
nor U6522 (N_6522,N_2569,N_3505);
or U6523 (N_6523,N_4466,N_4377);
or U6524 (N_6524,N_2584,N_4336);
nor U6525 (N_6525,N_235,N_3552);
and U6526 (N_6526,N_3612,N_3631);
nor U6527 (N_6527,N_1971,N_1414);
or U6528 (N_6528,N_933,N_10);
nand U6529 (N_6529,N_1950,N_4686);
xnor U6530 (N_6530,N_1808,N_1764);
or U6531 (N_6531,N_3158,N_1723);
nand U6532 (N_6532,N_3183,N_3779);
nor U6533 (N_6533,N_2974,N_979);
nand U6534 (N_6534,N_591,N_2704);
and U6535 (N_6535,N_2537,N_4237);
or U6536 (N_6536,N_2032,N_3660);
and U6537 (N_6537,N_2492,N_4457);
and U6538 (N_6538,N_1611,N_4599);
and U6539 (N_6539,N_3356,N_1361);
and U6540 (N_6540,N_1625,N_1290);
nand U6541 (N_6541,N_102,N_751);
xor U6542 (N_6542,N_202,N_948);
nand U6543 (N_6543,N_4448,N_2601);
and U6544 (N_6544,N_3950,N_2251);
xor U6545 (N_6545,N_3059,N_2062);
or U6546 (N_6546,N_4847,N_3190);
and U6547 (N_6547,N_2541,N_2201);
nor U6548 (N_6548,N_1714,N_4592);
and U6549 (N_6549,N_1866,N_2259);
or U6550 (N_6550,N_3053,N_4103);
or U6551 (N_6551,N_1930,N_4537);
nor U6552 (N_6552,N_2739,N_2242);
xnor U6553 (N_6553,N_2773,N_4219);
or U6554 (N_6554,N_2623,N_3758);
nand U6555 (N_6555,N_342,N_64);
nand U6556 (N_6556,N_2720,N_1857);
and U6557 (N_6557,N_2665,N_4133);
nor U6558 (N_6558,N_3043,N_3531);
nand U6559 (N_6559,N_4314,N_1524);
and U6560 (N_6560,N_3944,N_1727);
and U6561 (N_6561,N_4600,N_830);
or U6562 (N_6562,N_782,N_2149);
xor U6563 (N_6563,N_2305,N_525);
or U6564 (N_6564,N_4519,N_3445);
and U6565 (N_6565,N_24,N_3214);
nand U6566 (N_6566,N_3285,N_451);
and U6567 (N_6567,N_2069,N_3685);
nor U6568 (N_6568,N_600,N_2030);
nand U6569 (N_6569,N_593,N_4215);
nor U6570 (N_6570,N_2375,N_1207);
nand U6571 (N_6571,N_1545,N_3359);
nand U6572 (N_6572,N_4626,N_2841);
xnor U6573 (N_6573,N_1313,N_1367);
nor U6574 (N_6574,N_1815,N_4463);
and U6575 (N_6575,N_4505,N_481);
or U6576 (N_6576,N_4386,N_2610);
or U6577 (N_6577,N_3925,N_1343);
and U6578 (N_6578,N_2598,N_1286);
nor U6579 (N_6579,N_4388,N_4873);
xnor U6580 (N_6580,N_4963,N_34);
or U6581 (N_6581,N_3405,N_3128);
nand U6582 (N_6582,N_4641,N_4627);
and U6583 (N_6583,N_2382,N_3967);
or U6584 (N_6584,N_1151,N_3935);
or U6585 (N_6585,N_813,N_3592);
and U6586 (N_6586,N_1036,N_90);
and U6587 (N_6587,N_2227,N_3762);
nor U6588 (N_6588,N_3413,N_4556);
and U6589 (N_6589,N_2698,N_4543);
or U6590 (N_6590,N_2301,N_3947);
xnor U6591 (N_6591,N_456,N_4733);
or U6592 (N_6592,N_1316,N_2079);
nand U6593 (N_6593,N_2520,N_3305);
nor U6594 (N_6594,N_108,N_1146);
nand U6595 (N_6595,N_2102,N_2327);
nor U6596 (N_6596,N_1973,N_4493);
nor U6597 (N_6597,N_4682,N_674);
nand U6598 (N_6598,N_2986,N_2108);
nor U6599 (N_6599,N_1297,N_1471);
nand U6600 (N_6600,N_4317,N_742);
and U6601 (N_6601,N_2247,N_3556);
nand U6602 (N_6602,N_3894,N_3452);
nor U6603 (N_6603,N_3716,N_423);
and U6604 (N_6604,N_1302,N_3794);
nand U6605 (N_6605,N_1830,N_2613);
nand U6606 (N_6606,N_4642,N_206);
and U6607 (N_6607,N_3326,N_668);
or U6608 (N_6608,N_1867,N_3755);
nand U6609 (N_6609,N_149,N_1623);
xor U6610 (N_6610,N_2916,N_4488);
xnor U6611 (N_6611,N_3730,N_4559);
and U6612 (N_6612,N_2716,N_4657);
xnor U6613 (N_6613,N_3296,N_1467);
and U6614 (N_6614,N_2365,N_200);
nand U6615 (N_6615,N_4093,N_4833);
and U6616 (N_6616,N_3641,N_4328);
xor U6617 (N_6617,N_841,N_4710);
nor U6618 (N_6618,N_3846,N_184);
or U6619 (N_6619,N_170,N_4122);
and U6620 (N_6620,N_3289,N_4117);
nor U6621 (N_6621,N_237,N_1504);
or U6622 (N_6622,N_3227,N_655);
or U6623 (N_6623,N_4304,N_4196);
nand U6624 (N_6624,N_585,N_2410);
or U6625 (N_6625,N_1013,N_3085);
xnor U6626 (N_6626,N_4585,N_4415);
or U6627 (N_6627,N_3006,N_214);
nor U6628 (N_6628,N_4742,N_2314);
nand U6629 (N_6629,N_2001,N_4949);
nor U6630 (N_6630,N_4145,N_3968);
and U6631 (N_6631,N_2272,N_1778);
and U6632 (N_6632,N_4811,N_879);
xor U6633 (N_6633,N_91,N_1084);
and U6634 (N_6634,N_1181,N_4691);
nand U6635 (N_6635,N_1347,N_2366);
and U6636 (N_6636,N_3878,N_4277);
and U6637 (N_6637,N_92,N_4050);
nand U6638 (N_6638,N_1241,N_124);
or U6639 (N_6639,N_924,N_4287);
nor U6640 (N_6640,N_700,N_2118);
or U6641 (N_6641,N_1201,N_1210);
nand U6642 (N_6642,N_1105,N_604);
and U6643 (N_6643,N_2960,N_3379);
and U6644 (N_6644,N_2448,N_3752);
or U6645 (N_6645,N_1927,N_1078);
nand U6646 (N_6646,N_2683,N_265);
and U6647 (N_6647,N_3723,N_3143);
nor U6648 (N_6648,N_878,N_103);
xnor U6649 (N_6649,N_1260,N_2465);
and U6650 (N_6650,N_3670,N_2728);
or U6651 (N_6651,N_4694,N_2484);
nand U6652 (N_6652,N_3909,N_3637);
or U6653 (N_6653,N_747,N_4431);
xor U6654 (N_6654,N_625,N_1477);
or U6655 (N_6655,N_4530,N_3193);
nand U6656 (N_6656,N_4789,N_3699);
nand U6657 (N_6657,N_3186,N_2883);
and U6658 (N_6658,N_2096,N_1219);
or U6659 (N_6659,N_4770,N_772);
or U6660 (N_6660,N_1199,N_983);
or U6661 (N_6661,N_1904,N_1520);
and U6662 (N_6662,N_1660,N_4203);
xnor U6663 (N_6663,N_4737,N_1033);
nand U6664 (N_6664,N_4802,N_2508);
nand U6665 (N_6665,N_4,N_1673);
or U6666 (N_6666,N_2414,N_3248);
and U6667 (N_6667,N_2095,N_2266);
or U6668 (N_6668,N_4162,N_3089);
xnor U6669 (N_6669,N_3041,N_554);
xor U6670 (N_6670,N_905,N_4423);
xor U6671 (N_6671,N_1541,N_849);
nand U6672 (N_6672,N_1575,N_728);
and U6673 (N_6673,N_3759,N_4251);
nand U6674 (N_6674,N_4140,N_1041);
and U6675 (N_6675,N_2264,N_199);
nand U6676 (N_6676,N_963,N_4045);
xor U6677 (N_6677,N_2132,N_1064);
and U6678 (N_6678,N_2162,N_3298);
or U6679 (N_6679,N_3240,N_3973);
or U6680 (N_6680,N_2454,N_1490);
and U6681 (N_6681,N_464,N_3566);
nand U6682 (N_6682,N_1322,N_1957);
or U6683 (N_6683,N_2870,N_756);
nand U6684 (N_6684,N_113,N_2742);
or U6685 (N_6685,N_4598,N_1214);
or U6686 (N_6686,N_3365,N_4786);
nand U6687 (N_6687,N_2529,N_4858);
or U6688 (N_6688,N_3673,N_1235);
nor U6689 (N_6689,N_89,N_1339);
xor U6690 (N_6690,N_449,N_443);
and U6691 (N_6691,N_4653,N_3023);
xor U6692 (N_6692,N_3722,N_4480);
and U6693 (N_6693,N_650,N_1138);
xnor U6694 (N_6694,N_1087,N_4300);
nand U6695 (N_6695,N_4637,N_2854);
xor U6696 (N_6696,N_3563,N_3415);
or U6697 (N_6697,N_4938,N_3117);
nor U6698 (N_6698,N_1672,N_597);
xor U6699 (N_6699,N_263,N_4572);
and U6700 (N_6700,N_599,N_2795);
nand U6701 (N_6701,N_3270,N_2576);
and U6702 (N_6702,N_1149,N_4217);
nand U6703 (N_6703,N_4943,N_3638);
nand U6704 (N_6704,N_765,N_1952);
or U6705 (N_6705,N_2772,N_3912);
or U6706 (N_6706,N_1327,N_1694);
or U6707 (N_6707,N_4185,N_3130);
and U6708 (N_6708,N_2906,N_3852);
xnor U6709 (N_6709,N_1345,N_4935);
nor U6710 (N_6710,N_1220,N_3431);
nor U6711 (N_6711,N_891,N_1111);
nand U6712 (N_6712,N_3943,N_4425);
nor U6713 (N_6713,N_426,N_1182);
and U6714 (N_6714,N_3872,N_4971);
nand U6715 (N_6715,N_4470,N_3469);
xor U6716 (N_6716,N_145,N_3727);
nor U6717 (N_6717,N_3358,N_4679);
or U6718 (N_6718,N_3203,N_4747);
nand U6719 (N_6719,N_3751,N_3784);
xnor U6720 (N_6720,N_3646,N_1682);
nand U6721 (N_6721,N_3027,N_1923);
nor U6722 (N_6722,N_2052,N_1117);
nor U6723 (N_6723,N_4784,N_2200);
and U6724 (N_6724,N_1075,N_3936);
nor U6725 (N_6725,N_219,N_3319);
or U6726 (N_6726,N_1955,N_1457);
or U6727 (N_6727,N_1368,N_1865);
or U6728 (N_6728,N_1920,N_4024);
nand U6729 (N_6729,N_1392,N_1141);
and U6730 (N_6730,N_1747,N_3623);
nand U6731 (N_6731,N_4934,N_1393);
nor U6732 (N_6732,N_2070,N_3253);
and U6733 (N_6733,N_3435,N_2579);
and U6734 (N_6734,N_2517,N_2905);
nand U6735 (N_6735,N_1907,N_3979);
nand U6736 (N_6736,N_2170,N_2687);
xnor U6737 (N_6737,N_1320,N_2545);
and U6738 (N_6738,N_3535,N_1627);
nand U6739 (N_6739,N_207,N_2229);
or U6740 (N_6740,N_967,N_461);
or U6741 (N_6741,N_1299,N_888);
and U6742 (N_6742,N_2315,N_2211);
or U6743 (N_6743,N_4329,N_1381);
nand U6744 (N_6744,N_1655,N_1364);
xor U6745 (N_6745,N_246,N_1400);
nand U6746 (N_6746,N_851,N_4054);
nor U6747 (N_6747,N_1,N_2178);
xnor U6748 (N_6748,N_4233,N_4081);
xor U6749 (N_6749,N_4322,N_4361);
and U6750 (N_6750,N_2891,N_4940);
nand U6751 (N_6751,N_2892,N_586);
nand U6752 (N_6752,N_2606,N_2504);
or U6753 (N_6753,N_783,N_509);
or U6754 (N_6754,N_1964,N_3721);
nor U6755 (N_6755,N_4238,N_3451);
and U6756 (N_6756,N_908,N_727);
xor U6757 (N_6757,N_355,N_4307);
nor U6758 (N_6758,N_1031,N_4621);
xor U6759 (N_6759,N_2446,N_3907);
nand U6760 (N_6760,N_4334,N_3874);
or U6761 (N_6761,N_25,N_1462);
nor U6762 (N_6762,N_440,N_3480);
and U6763 (N_6763,N_1704,N_1736);
or U6764 (N_6764,N_2216,N_3677);
xnor U6765 (N_6765,N_2885,N_4440);
and U6766 (N_6766,N_1067,N_845);
nor U6767 (N_6767,N_3931,N_666);
nor U6768 (N_6768,N_4633,N_4375);
and U6769 (N_6769,N_4533,N_1709);
or U6770 (N_6770,N_2067,N_3019);
xnor U6771 (N_6771,N_1301,N_738);
or U6772 (N_6772,N_606,N_3952);
nand U6773 (N_6773,N_1962,N_448);
nor U6774 (N_6774,N_416,N_2202);
and U6775 (N_6775,N_570,N_2066);
or U6776 (N_6776,N_4632,N_309);
and U6777 (N_6777,N_808,N_4955);
and U6778 (N_6778,N_1447,N_376);
and U6779 (N_6779,N_4900,N_2412);
or U6780 (N_6780,N_4183,N_1123);
or U6781 (N_6781,N_1902,N_1006);
nor U6782 (N_6782,N_4487,N_2377);
xor U6783 (N_6783,N_3810,N_3514);
nor U6784 (N_6784,N_4843,N_353);
xnor U6785 (N_6785,N_300,N_2105);
and U6786 (N_6786,N_284,N_1190);
xnor U6787 (N_6787,N_549,N_3385);
nand U6788 (N_6788,N_2487,N_3042);
nand U6789 (N_6789,N_717,N_2046);
and U6790 (N_6790,N_1721,N_2572);
xor U6791 (N_6791,N_147,N_1916);
xor U6792 (N_6792,N_4445,N_889);
or U6793 (N_6793,N_3157,N_4720);
and U6794 (N_6794,N_1391,N_964);
nor U6795 (N_6795,N_1659,N_4296);
and U6796 (N_6796,N_1051,N_424);
nand U6797 (N_6797,N_3589,N_1441);
and U6798 (N_6798,N_1338,N_3038);
and U6799 (N_6799,N_3608,N_3503);
xnor U6800 (N_6800,N_3426,N_4892);
nand U6801 (N_6801,N_358,N_1807);
and U6802 (N_6802,N_3891,N_4258);
xnor U6803 (N_6803,N_3261,N_2927);
nand U6804 (N_6804,N_662,N_4761);
nor U6805 (N_6805,N_1871,N_4048);
nand U6806 (N_6806,N_3977,N_4222);
nand U6807 (N_6807,N_643,N_1754);
or U6808 (N_6808,N_4838,N_3081);
nand U6809 (N_6809,N_1698,N_4295);
or U6810 (N_6810,N_2640,N_2664);
nand U6811 (N_6811,N_3281,N_2061);
nor U6812 (N_6812,N_1027,N_1628);
or U6813 (N_6813,N_3327,N_2115);
nor U6814 (N_6814,N_572,N_2858);
nor U6815 (N_6815,N_2021,N_3959);
and U6816 (N_6816,N_678,N_2758);
nor U6817 (N_6817,N_2188,N_595);
nor U6818 (N_6818,N_4311,N_2724);
xnor U6819 (N_6819,N_3972,N_2621);
or U6820 (N_6820,N_1786,N_4010);
or U6821 (N_6821,N_4685,N_3015);
xnor U6822 (N_6822,N_2933,N_3832);
xnor U6823 (N_6823,N_3083,N_367);
nor U6824 (N_6824,N_2390,N_3462);
nand U6825 (N_6825,N_1277,N_3527);
or U6826 (N_6826,N_1573,N_2996);
or U6827 (N_6827,N_1578,N_1586);
or U6828 (N_6828,N_4757,N_3055);
nand U6829 (N_6829,N_3244,N_798);
nand U6830 (N_6830,N_603,N_4954);
nand U6831 (N_6831,N_3020,N_3515);
or U6832 (N_6832,N_4750,N_624);
nand U6833 (N_6833,N_240,N_1996);
and U6834 (N_6834,N_1906,N_969);
nor U6835 (N_6835,N_4713,N_2186);
nand U6836 (N_6836,N_510,N_524);
nor U6837 (N_6837,N_840,N_4034);
nor U6838 (N_6838,N_316,N_2798);
xnor U6839 (N_6839,N_1763,N_616);
or U6840 (N_6840,N_1656,N_4624);
or U6841 (N_6841,N_3671,N_2709);
and U6842 (N_6842,N_2086,N_4260);
xnor U6843 (N_6843,N_4266,N_4428);
nor U6844 (N_6844,N_2964,N_2995);
nor U6845 (N_6845,N_2679,N_734);
or U6846 (N_6846,N_994,N_1291);
and U6847 (N_6847,N_1435,N_4972);
nor U6848 (N_6848,N_802,N_1568);
or U6849 (N_6849,N_3692,N_4548);
xor U6850 (N_6850,N_377,N_1061);
xnor U6851 (N_6851,N_2989,N_3294);
nand U6852 (N_6852,N_2281,N_3222);
xor U6853 (N_6853,N_2164,N_4175);
and U6854 (N_6854,N_1547,N_4474);
and U6855 (N_6855,N_980,N_3984);
and U6856 (N_6856,N_2861,N_1088);
nand U6857 (N_6857,N_2244,N_175);
nor U6858 (N_6858,N_2121,N_3299);
nor U6859 (N_6859,N_3003,N_435);
xnor U6860 (N_6860,N_1357,N_2962);
and U6861 (N_6861,N_1186,N_3422);
or U6862 (N_6862,N_4246,N_745);
and U6863 (N_6863,N_433,N_2340);
xnor U6864 (N_6864,N_4662,N_4112);
and U6865 (N_6865,N_1057,N_140);
or U6866 (N_6866,N_1019,N_238);
xnor U6867 (N_6867,N_940,N_4207);
and U6868 (N_6868,N_2400,N_3618);
nor U6869 (N_6869,N_1992,N_1314);
xor U6870 (N_6870,N_1799,N_412);
xnor U6871 (N_6871,N_276,N_1272);
xnor U6872 (N_6872,N_3586,N_2971);
xnor U6873 (N_6873,N_484,N_1222);
nor U6874 (N_6874,N_1980,N_380);
or U6875 (N_6875,N_1759,N_422);
nand U6876 (N_6876,N_4538,N_1399);
nor U6877 (N_6877,N_3163,N_3210);
and U6878 (N_6878,N_822,N_2846);
nand U6879 (N_6879,N_4383,N_1240);
nand U6880 (N_6880,N_1032,N_4546);
nand U6881 (N_6881,N_227,N_191);
nand U6882 (N_6882,N_1832,N_579);
nand U6883 (N_6883,N_4494,N_2221);
and U6884 (N_6884,N_2844,N_167);
nor U6885 (N_6885,N_2489,N_4700);
nor U6886 (N_6886,N_3118,N_2157);
nand U6887 (N_6887,N_563,N_4309);
nand U6888 (N_6888,N_897,N_4709);
and U6889 (N_6889,N_4372,N_4031);
and U6890 (N_6890,N_2490,N_2088);
nand U6891 (N_6891,N_3223,N_2542);
nand U6892 (N_6892,N_4484,N_3661);
xnor U6893 (N_6893,N_3068,N_3394);
nor U6894 (N_6894,N_1107,N_578);
or U6895 (N_6895,N_2651,N_2754);
nand U6896 (N_6896,N_3504,N_3497);
or U6897 (N_6897,N_2144,N_1664);
or U6898 (N_6898,N_4362,N_489);
xnor U6899 (N_6899,N_4547,N_4382);
xnor U6900 (N_6900,N_2647,N_3276);
and U6901 (N_6901,N_4864,N_3033);
nor U6902 (N_6902,N_3642,N_1258);
xor U6903 (N_6903,N_1080,N_4808);
or U6904 (N_6904,N_1612,N_3734);
nand U6905 (N_6905,N_4214,N_1065);
nand U6906 (N_6906,N_4061,N_4721);
and U6907 (N_6907,N_1522,N_3292);
xor U6908 (N_6908,N_621,N_3834);
nor U6909 (N_6909,N_100,N_4665);
nand U6910 (N_6910,N_1959,N_2873);
and U6911 (N_6911,N_2705,N_4004);
xnor U6912 (N_6912,N_2808,N_817);
and U6913 (N_6913,N_2404,N_4560);
or U6914 (N_6914,N_2554,N_344);
and U6915 (N_6915,N_1972,N_3813);
and U6916 (N_6916,N_3114,N_3094);
xor U6917 (N_6917,N_1581,N_4991);
nand U6918 (N_6918,N_3521,N_3189);
nor U6919 (N_6919,N_4797,N_1826);
or U6920 (N_6920,N_3461,N_1454);
xor U6921 (N_6921,N_2142,N_4677);
nand U6922 (N_6922,N_4416,N_4941);
nand U6923 (N_6923,N_4478,N_2853);
nor U6924 (N_6924,N_4206,N_4044);
nand U6925 (N_6925,N_3509,N_4098);
and U6926 (N_6926,N_675,N_1165);
or U6927 (N_6927,N_1011,N_1459);
xor U6928 (N_6928,N_1649,N_2336);
nand U6929 (N_6929,N_4152,N_142);
and U6930 (N_6930,N_3291,N_1752);
xor U6931 (N_6931,N_3746,N_4528);
or U6932 (N_6932,N_2780,N_1353);
and U6933 (N_6933,N_584,N_1693);
or U6934 (N_6934,N_1528,N_93);
nor U6935 (N_6935,N_898,N_2093);
and U6936 (N_6936,N_3781,N_2468);
xnor U6937 (N_6937,N_1486,N_2482);
nor U6938 (N_6938,N_3000,N_2566);
or U6939 (N_6939,N_3655,N_3150);
xnor U6940 (N_6940,N_2516,N_1771);
or U6941 (N_6941,N_3045,N_1858);
xnor U6942 (N_6942,N_821,N_4339);
or U6943 (N_6943,N_4213,N_296);
xnor U6944 (N_6944,N_3963,N_3017);
nor U6945 (N_6945,N_1073,N_764);
or U6946 (N_6946,N_1365,N_3022);
and U6947 (N_6947,N_815,N_2976);
xnor U6948 (N_6948,N_52,N_2731);
or U6949 (N_6949,N_1855,N_1909);
nor U6950 (N_6950,N_1226,N_2618);
nor U6951 (N_6951,N_1595,N_4430);
and U6952 (N_6952,N_4166,N_1160);
and U6953 (N_6953,N_1816,N_328);
xor U6954 (N_6954,N_2228,N_4523);
and U6955 (N_6955,N_1480,N_4756);
xor U6956 (N_6956,N_2130,N_2374);
nor U6957 (N_6957,N_3402,N_3220);
nand U6958 (N_6958,N_3571,N_3786);
nand U6959 (N_6959,N_4595,N_3212);
xor U6960 (N_6960,N_1215,N_601);
nand U6961 (N_6961,N_3856,N_4279);
nand U6962 (N_6962,N_999,N_1558);
nand U6963 (N_6963,N_1725,N_2734);
xor U6964 (N_6964,N_911,N_1936);
xnor U6965 (N_6965,N_45,N_3300);
or U6966 (N_6966,N_4444,N_1022);
or U6967 (N_6967,N_4337,N_1940);
and U6968 (N_6968,N_4324,N_1404);
nand U6969 (N_6969,N_1406,N_4358);
nand U6970 (N_6970,N_4462,N_1616);
and U6971 (N_6971,N_4089,N_1699);
nor U6972 (N_6972,N_156,N_1440);
or U6973 (N_6973,N_3161,N_1560);
nand U6974 (N_6974,N_267,N_1170);
nand U6975 (N_6975,N_54,N_1497);
nor U6976 (N_6976,N_4086,N_1305);
nand U6977 (N_6977,N_2128,N_4053);
and U6978 (N_6978,N_2137,N_112);
xnor U6979 (N_6979,N_2768,N_1306);
nand U6980 (N_6980,N_2587,N_4969);
nand U6981 (N_6981,N_3753,N_2277);
nor U6982 (N_6982,N_3990,N_4020);
or U6983 (N_6983,N_1177,N_1405);
xor U6984 (N_6984,N_2988,N_676);
nand U6985 (N_6985,N_3934,N_2852);
nand U6986 (N_6986,N_3502,N_1737);
nor U6987 (N_6987,N_1188,N_2406);
or U6988 (N_6988,N_4917,N_1566);
nand U6989 (N_6989,N_3922,N_800);
and U6990 (N_6990,N_596,N_4725);
nor U6991 (N_6991,N_4916,N_2749);
nor U6992 (N_6992,N_2479,N_669);
and U6993 (N_6993,N_858,N_3140);
and U6994 (N_6994,N_17,N_562);
nand U6995 (N_6995,N_766,N_319);
nand U6996 (N_6996,N_2155,N_1221);
xnor U6997 (N_6997,N_797,N_4221);
nor U6998 (N_6998,N_1376,N_41);
nand U6999 (N_6999,N_3073,N_4804);
or U7000 (N_7000,N_3788,N_3111);
nor U7001 (N_7001,N_3791,N_2025);
or U7002 (N_7002,N_2565,N_3654);
and U7003 (N_7003,N_1384,N_4072);
and U7004 (N_7004,N_1580,N_1642);
nand U7005 (N_7005,N_895,N_1337);
nand U7006 (N_7006,N_4526,N_3484);
or U7007 (N_7007,N_2010,N_1056);
xnor U7008 (N_7008,N_3736,N_4926);
or U7009 (N_7009,N_4499,N_511);
xor U7010 (N_7010,N_4230,N_3133);
nor U7011 (N_7011,N_2810,N_5);
nand U7012 (N_7012,N_2103,N_653);
or U7013 (N_7013,N_1289,N_3428);
nor U7014 (N_7014,N_3275,N_2006);
xnor U7015 (N_7015,N_743,N_3058);
and U7016 (N_7016,N_1746,N_3981);
nor U7017 (N_7017,N_3765,N_1424);
nor U7018 (N_7018,N_882,N_1676);
and U7019 (N_7019,N_4973,N_3447);
or U7020 (N_7020,N_955,N_3371);
xor U7021 (N_7021,N_3709,N_4190);
and U7022 (N_7022,N_1722,N_1697);
xnor U7023 (N_7023,N_1924,N_4999);
and U7024 (N_7024,N_2169,N_3739);
and U7025 (N_7025,N_744,N_2447);
or U7026 (N_7026,N_4280,N_4209);
or U7027 (N_7027,N_4981,N_3249);
nor U7028 (N_7028,N_4446,N_3376);
and U7029 (N_7029,N_923,N_2715);
or U7030 (N_7030,N_239,N_497);
nor U7031 (N_7031,N_1634,N_1860);
xor U7032 (N_7032,N_3841,N_4932);
or U7033 (N_7033,N_1789,N_2553);
nor U7034 (N_7034,N_2886,N_3873);
xnor U7035 (N_7035,N_3821,N_228);
and U7036 (N_7036,N_2670,N_3278);
or U7037 (N_7037,N_229,N_576);
and U7038 (N_7038,N_3653,N_4729);
nand U7039 (N_7039,N_1113,N_2848);
nand U7040 (N_7040,N_3098,N_613);
and U7041 (N_7041,N_3799,N_4907);
xnor U7042 (N_7042,N_4078,N_1470);
nor U7043 (N_7043,N_2889,N_2730);
nor U7044 (N_7044,N_387,N_4256);
nor U7045 (N_7045,N_444,N_3565);
nor U7046 (N_7046,N_3386,N_4518);
or U7047 (N_7047,N_2503,N_2136);
or U7048 (N_7048,N_589,N_4134);
nor U7049 (N_7049,N_1978,N_543);
nor U7050 (N_7050,N_3101,N_4760);
xnor U7051 (N_7051,N_2597,N_2706);
xnor U7052 (N_7052,N_4989,N_223);
or U7053 (N_7053,N_1074,N_4298);
nor U7054 (N_7054,N_3334,N_1539);
nand U7055 (N_7055,N_9,N_1465);
or U7056 (N_7056,N_1535,N_3896);
nor U7057 (N_7057,N_225,N_3569);
nand U7058 (N_7058,N_4860,N_834);
xnor U7059 (N_7059,N_1777,N_1853);
nand U7060 (N_7060,N_4188,N_3113);
and U7061 (N_7061,N_2249,N_1484);
nor U7062 (N_7062,N_3120,N_3398);
or U7063 (N_7063,N_2381,N_2224);
and U7064 (N_7064,N_1093,N_1281);
and U7065 (N_7065,N_4150,N_3496);
and U7066 (N_7066,N_654,N_3400);
nor U7067 (N_7067,N_1416,N_2286);
and U7068 (N_7068,N_988,N_3525);
nand U7069 (N_7069,N_2746,N_2037);
or U7070 (N_7070,N_719,N_3127);
nand U7071 (N_7071,N_1369,N_1052);
nor U7072 (N_7072,N_1505,N_2383);
and U7073 (N_7073,N_997,N_3151);
and U7074 (N_7074,N_2438,N_1043);
and U7075 (N_7075,N_4831,N_4603);
and U7076 (N_7076,N_1748,N_369);
xor U7077 (N_7077,N_1300,N_1811);
xnor U7078 (N_7078,N_731,N_3666);
or U7079 (N_7079,N_1641,N_4286);
nand U7080 (N_7080,N_977,N_1020);
nor U7081 (N_7081,N_1779,N_1042);
or U7082 (N_7082,N_1382,N_2437);
or U7083 (N_7083,N_1350,N_2253);
nor U7084 (N_7084,N_4313,N_519);
xnor U7085 (N_7085,N_395,N_4616);
nor U7086 (N_7086,N_2867,N_1905);
or U7087 (N_7087,N_3969,N_311);
xnor U7088 (N_7088,N_2257,N_3103);
xnor U7089 (N_7089,N_564,N_3363);
nand U7090 (N_7090,N_4118,N_4562);
and U7091 (N_7091,N_2401,N_2189);
xnor U7092 (N_7092,N_3837,N_3235);
nand U7093 (N_7093,N_2939,N_4465);
nor U7094 (N_7094,N_3965,N_1311);
and U7095 (N_7095,N_2615,N_2710);
xnor U7096 (N_7096,N_1630,N_4673);
or U7097 (N_7097,N_759,N_136);
nand U7098 (N_7098,N_4109,N_4850);
nand U7099 (N_7099,N_3772,N_3057);
xnor U7100 (N_7100,N_1362,N_4032);
and U7101 (N_7101,N_2904,N_4852);
xnor U7102 (N_7102,N_3224,N_277);
nand U7103 (N_7103,N_2152,N_4891);
or U7104 (N_7104,N_852,N_4882);
and U7105 (N_7105,N_4319,N_945);
nand U7106 (N_7106,N_4834,N_482);
xnor U7107 (N_7107,N_2333,N_2578);
and U7108 (N_7108,N_1126,N_1066);
xor U7109 (N_7109,N_2931,N_3830);
nand U7110 (N_7110,N_4774,N_2262);
xnor U7111 (N_7111,N_3603,N_1429);
nand U7112 (N_7112,N_257,N_439);
and U7113 (N_7113,N_1483,N_2500);
nand U7114 (N_7114,N_431,N_1349);
nand U7115 (N_7115,N_2469,N_373);
and U7116 (N_7116,N_2312,N_931);
or U7117 (N_7117,N_3957,N_4426);
xor U7118 (N_7118,N_190,N_2919);
and U7119 (N_7119,N_472,N_4798);
or U7120 (N_7120,N_3407,N_762);
or U7121 (N_7121,N_3548,N_1554);
nand U7122 (N_7122,N_3880,N_686);
nor U7123 (N_7123,N_4982,N_4069);
and U7124 (N_7124,N_1854,N_2820);
xnor U7125 (N_7125,N_2317,N_295);
nand U7126 (N_7126,N_2439,N_4625);
or U7127 (N_7127,N_3997,N_478);
nor U7128 (N_7128,N_4791,N_2344);
nand U7129 (N_7129,N_3011,N_4931);
and U7130 (N_7130,N_43,N_2285);
nor U7131 (N_7131,N_3474,N_3865);
nor U7132 (N_7132,N_2550,N_3995);
and U7133 (N_7133,N_3658,N_801);
or U7134 (N_7134,N_2806,N_414);
nor U7135 (N_7135,N_486,N_4790);
nor U7136 (N_7136,N_2973,N_4866);
and U7137 (N_7137,N_1244,N_4735);
nor U7138 (N_7138,N_2536,N_1948);
or U7139 (N_7139,N_154,N_1868);
nand U7140 (N_7140,N_962,N_1516);
nor U7141 (N_7141,N_831,N_66);
nor U7142 (N_7142,N_4777,N_2282);
xnor U7143 (N_7143,N_3306,N_1620);
or U7144 (N_7144,N_3861,N_4853);
or U7145 (N_7145,N_2521,N_2859);
and U7146 (N_7146,N_3392,N_2408);
or U7147 (N_7147,N_4809,N_1677);
xor U7148 (N_7148,N_4410,N_2245);
nor U7149 (N_7149,N_699,N_2384);
xor U7150 (N_7150,N_2752,N_1716);
or U7151 (N_7151,N_3062,N_1733);
nand U7152 (N_7152,N_1448,N_4178);
nand U7153 (N_7153,N_4138,N_705);
xnor U7154 (N_7154,N_4915,N_1238);
or U7155 (N_7155,N_3013,N_3317);
or U7156 (N_7156,N_2335,N_85);
xor U7157 (N_7157,N_22,N_4163);
and U7158 (N_7158,N_3551,N_4076);
xor U7159 (N_7159,N_1932,N_121);
and U7160 (N_7160,N_215,N_1129);
or U7161 (N_7161,N_2083,N_4801);
and U7162 (N_7162,N_4996,N_356);
nor U7163 (N_7163,N_3459,N_1445);
nor U7164 (N_7164,N_2949,N_418);
nand U7165 (N_7165,N_2510,N_2686);
xor U7166 (N_7166,N_2696,N_3790);
or U7167 (N_7167,N_2657,N_480);
or U7168 (N_7168,N_1836,N_2678);
nor U7169 (N_7169,N_3414,N_2669);
xnor U7170 (N_7170,N_2877,N_1139);
nor U7171 (N_7171,N_74,N_2767);
nor U7172 (N_7172,N_3857,N_3627);
or U7173 (N_7173,N_3368,N_1250);
xnor U7174 (N_7174,N_4785,N_4764);
nand U7175 (N_7175,N_715,N_3584);
xor U7176 (N_7176,N_1385,N_4732);
and U7177 (N_7177,N_3159,N_4923);
and U7178 (N_7178,N_1398,N_4201);
or U7179 (N_7179,N_1175,N_3961);
nand U7180 (N_7180,N_1243,N_1937);
xor U7181 (N_7181,N_3672,N_2125);
or U7182 (N_7182,N_1879,N_4271);
xor U7183 (N_7183,N_1648,N_4427);
nand U7184 (N_7184,N_146,N_1851);
nor U7185 (N_7185,N_3044,N_665);
and U7186 (N_7186,N_2607,N_3442);
nand U7187 (N_7187,N_4536,N_3330);
nor U7188 (N_7188,N_4368,N_216);
nand U7189 (N_7189,N_1913,N_3975);
and U7190 (N_7190,N_1790,N_1415);
or U7191 (N_7191,N_4365,N_769);
and U7192 (N_7192,N_899,N_392);
or U7193 (N_7193,N_4005,N_1744);
nand U7194 (N_7194,N_4312,N_3802);
xor U7195 (N_7195,N_2287,N_1225);
or U7196 (N_7196,N_4606,N_548);
and U7197 (N_7197,N_3701,N_2741);
xnor U7198 (N_7198,N_3776,N_3075);
nor U7199 (N_7199,N_3574,N_1144);
xor U7200 (N_7200,N_2552,N_2512);
nand U7201 (N_7201,N_1321,N_1945);
xor U7202 (N_7202,N_2441,N_371);
nand U7203 (N_7203,N_3690,N_4803);
and U7204 (N_7204,N_255,N_3639);
nor U7205 (N_7205,N_4588,N_2845);
or U7206 (N_7206,N_4420,N_2302);
nor U7207 (N_7207,N_1565,N_3624);
nand U7208 (N_7208,N_3109,N_1081);
nand U7209 (N_7209,N_2934,N_3032);
or U7210 (N_7210,N_2757,N_4964);
or U7211 (N_7211,N_4829,N_259);
nor U7212 (N_7212,N_2518,N_691);
nand U7213 (N_7213,N_313,N_2138);
or U7214 (N_7214,N_1178,N_3454);
or U7215 (N_7215,N_2068,N_3871);
nand U7216 (N_7216,N_1103,N_141);
or U7217 (N_7217,N_372,N_279);
nor U7218 (N_7218,N_2776,N_4810);
or U7219 (N_7219,N_4772,N_3743);
nor U7220 (N_7220,N_3737,N_1683);
and U7221 (N_7221,N_1970,N_1603);
or U7222 (N_7222,N_763,N_1140);
nand U7223 (N_7223,N_1383,N_1550);
nor U7224 (N_7224,N_1028,N_1372);
nor U7225 (N_7225,N_197,N_1010);
nand U7226 (N_7226,N_4545,N_4477);
nand U7227 (N_7227,N_2209,N_627);
and U7228 (N_7228,N_2402,N_826);
nor U7229 (N_7229,N_221,N_536);
nor U7230 (N_7230,N_4863,N_886);
xor U7231 (N_7231,N_1943,N_2343);
or U7232 (N_7232,N_1375,N_3599);
and U7233 (N_7233,N_35,N_1908);
xnor U7234 (N_7234,N_2353,N_2222);
and U7235 (N_7235,N_340,N_1529);
nand U7236 (N_7236,N_3037,N_329);
or U7237 (N_7237,N_3492,N_4392);
and U7238 (N_7238,N_3619,N_2967);
nor U7239 (N_7239,N_3198,N_1762);
nand U7240 (N_7240,N_4751,N_2558);
xnor U7241 (N_7241,N_4554,N_2923);
and U7242 (N_7242,N_59,N_3493);
xor U7243 (N_7243,N_160,N_739);
nor U7244 (N_7244,N_608,N_1767);
xnor U7245 (N_7245,N_4063,N_1812);
xor U7246 (N_7246,N_2166,N_4371);
or U7247 (N_7247,N_1072,N_2625);
nand U7248 (N_7248,N_1083,N_3209);
nor U7249 (N_7249,N_401,N_1695);
or U7250 (N_7250,N_2711,N_1564);
nor U7251 (N_7251,N_2694,N_2589);
and U7252 (N_7252,N_3307,N_4517);
nand U7253 (N_7253,N_1899,N_247);
and U7254 (N_7254,N_1206,N_2294);
or U7255 (N_7255,N_954,N_1979);
nand U7256 (N_7256,N_2573,N_1850);
and U7257 (N_7257,N_278,N_1801);
nor U7258 (N_7258,N_1254,N_1148);
nand U7259 (N_7259,N_1556,N_3506);
and U7260 (N_7260,N_4806,N_992);
xnor U7261 (N_7261,N_3384,N_4587);
or U7262 (N_7262,N_466,N_4660);
and U7263 (N_7263,N_3153,N_3046);
nor U7264 (N_7264,N_224,N_3930);
xnor U7265 (N_7265,N_3313,N_4235);
xor U7266 (N_7266,N_4577,N_1458);
and U7267 (N_7267,N_2111,N_1925);
nand U7268 (N_7268,N_752,N_4405);
xor U7269 (N_7269,N_520,N_4620);
nand U7270 (N_7270,N_4082,N_1421);
xor U7271 (N_7271,N_2126,N_2427);
and U7272 (N_7272,N_4848,N_2910);
nor U7273 (N_7273,N_4121,N_3048);
and U7274 (N_7274,N_792,N_49);
and U7275 (N_7275,N_1824,N_3510);
nand U7276 (N_7276,N_2252,N_3399);
nand U7277 (N_7277,N_53,N_1770);
and U7278 (N_7278,N_2770,N_413);
xor U7279 (N_7279,N_3887,N_343);
xor U7280 (N_7280,N_2644,N_3924);
nand U7281 (N_7281,N_2298,N_331);
xnor U7282 (N_7282,N_3108,N_3899);
xor U7283 (N_7283,N_2603,N_2175);
xnor U7284 (N_7284,N_4862,N_307);
or U7285 (N_7285,N_2645,N_646);
nand U7286 (N_7286,N_3233,N_3490);
nand U7287 (N_7287,N_3956,N_3911);
or U7288 (N_7288,N_288,N_1411);
and U7289 (N_7289,N_1934,N_250);
xnor U7290 (N_7290,N_2223,N_3898);
or U7291 (N_7291,N_4504,N_4817);
and U7292 (N_7292,N_4077,N_690);
nand U7293 (N_7293,N_2278,N_3374);
nand U7294 (N_7294,N_4779,N_3171);
xor U7295 (N_7295,N_1670,N_3230);
nand U7296 (N_7296,N_609,N_4669);
nor U7297 (N_7297,N_1831,N_3938);
xor U7298 (N_7298,N_4257,N_2570);
nand U7299 (N_7299,N_551,N_2600);
and U7300 (N_7300,N_2230,N_2398);
and U7301 (N_7301,N_4765,N_1261);
or U7302 (N_7302,N_4723,N_3715);
nor U7303 (N_7303,N_4241,N_4000);
nor U7304 (N_7304,N_508,N_4881);
or U7305 (N_7305,N_1434,N_495);
or U7306 (N_7306,N_3411,N_3425);
nor U7307 (N_7307,N_2622,N_3696);
xor U7308 (N_7308,N_332,N_2289);
xnor U7309 (N_7309,N_3982,N_4331);
nor U7310 (N_7310,N_927,N_3998);
or U7311 (N_7311,N_4903,N_3954);
and U7312 (N_7312,N_4395,N_1591);
nor U7313 (N_7313,N_2719,N_3457);
xor U7314 (N_7314,N_3689,N_3125);
xnor U7315 (N_7315,N_4986,N_3740);
nand U7316 (N_7316,N_2470,N_1802);
xnor U7317 (N_7317,N_4130,N_4702);
nor U7318 (N_7318,N_3604,N_1517);
or U7319 (N_7319,N_271,N_1045);
or U7320 (N_7320,N_2369,N_1898);
or U7321 (N_7321,N_134,N_3711);
nor U7322 (N_7322,N_4500,N_900);
nor U7323 (N_7323,N_2177,N_2100);
xor U7324 (N_7324,N_498,N_4359);
nor U7325 (N_7325,N_2811,N_4367);
nand U7326 (N_7326,N_4990,N_2708);
and U7327 (N_7327,N_4035,N_2897);
or U7328 (N_7328,N_2094,N_4155);
or U7329 (N_7329,N_1479,N_3879);
and U7330 (N_7330,N_1476,N_651);
xor U7331 (N_7331,N_31,N_857);
xor U7332 (N_7332,N_773,N_3686);
xor U7333 (N_7333,N_4762,N_3720);
xor U7334 (N_7334,N_4491,N_2735);
and U7335 (N_7335,N_4845,N_2629);
nand U7336 (N_7336,N_3396,N_4648);
nor U7337 (N_7337,N_1914,N_1422);
nand U7338 (N_7338,N_4268,N_4308);
and U7339 (N_7339,N_1442,N_2513);
and U7340 (N_7340,N_590,N_2004);
xor U7341 (N_7341,N_2187,N_2237);
and U7342 (N_7342,N_2648,N_4584);
nand U7343 (N_7343,N_1842,N_1487);
nand U7344 (N_7344,N_2016,N_1765);
nand U7345 (N_7345,N_1840,N_1212);
xor U7346 (N_7346,N_4441,N_1825);
nor U7347 (N_7347,N_119,N_853);
nor U7348 (N_7348,N_4501,N_2692);
nor U7349 (N_7349,N_4763,N_555);
nor U7350 (N_7350,N_1154,N_4409);
and U7351 (N_7351,N_2901,N_4959);
nand U7352 (N_7352,N_2154,N_3234);
nor U7353 (N_7353,N_3202,N_1552);
nand U7354 (N_7354,N_941,N_417);
xnor U7355 (N_7355,N_1891,N_2241);
nand U7356 (N_7356,N_1155,N_1987);
xnor U7357 (N_7357,N_2751,N_1944);
or U7358 (N_7358,N_3668,N_2801);
nand U7359 (N_7359,N_2038,N_1651);
nor U7360 (N_7360,N_362,N_1410);
or U7361 (N_7361,N_4435,N_2081);
nand U7362 (N_7362,N_2775,N_3750);
xnor U7363 (N_7363,N_181,N_4646);
and U7364 (N_7364,N_541,N_2659);
xor U7365 (N_7365,N_1167,N_1839);
or U7366 (N_7366,N_1732,N_2535);
xor U7367 (N_7367,N_3478,N_3987);
or U7368 (N_7368,N_2330,N_789);
nor U7369 (N_7369,N_3336,N_253);
nor U7370 (N_7370,N_2458,N_4960);
and U7371 (N_7371,N_4571,N_1507);
xnor U7372 (N_7372,N_938,N_352);
nand U7373 (N_7373,N_99,N_1810);
xor U7374 (N_7374,N_111,N_2755);
and U7375 (N_7375,N_1533,N_681);
and U7376 (N_7376,N_1488,N_3175);
nor U7377 (N_7377,N_2831,N_3974);
or U7378 (N_7378,N_2306,N_4281);
nand U7379 (N_7379,N_2063,N_4754);
or U7380 (N_7380,N_3201,N_959);
and U7381 (N_7381,N_2595,N_846);
nor U7382 (N_7382,N_82,N_2814);
or U7383 (N_7383,N_2502,N_1319);
and U7384 (N_7384,N_2476,N_198);
xnor U7385 (N_7385,N_242,N_4080);
xor U7386 (N_7386,N_3621,N_2723);
nor U7387 (N_7387,N_1985,N_2970);
xnor U7388 (N_7388,N_474,N_1055);
xor U7389 (N_7389,N_4363,N_1109);
nand U7390 (N_7390,N_1273,N_2738);
nor U7391 (N_7391,N_3116,N_3332);
and U7392 (N_7392,N_4524,N_3883);
nand U7393 (N_7393,N_2797,N_3590);
nor U7394 (N_7394,N_1735,N_1730);
nor U7395 (N_7395,N_471,N_2633);
and U7396 (N_7396,N_2588,N_4896);
xor U7397 (N_7397,N_2463,N_4532);
nor U7398 (N_7398,N_1423,N_4970);
xor U7399 (N_7399,N_4778,N_3069);
xnor U7400 (N_7400,N_2009,N_4240);
xor U7401 (N_7401,N_1675,N_1713);
or U7402 (N_7402,N_1548,N_4146);
nand U7403 (N_7403,N_2722,N_120);
nor U7404 (N_7404,N_212,N_741);
and U7405 (N_7405,N_4267,N_4247);
and U7406 (N_7406,N_2445,N_4419);
nor U7407 (N_7407,N_3286,N_1264);
or U7408 (N_7408,N_1395,N_1615);
nor U7409 (N_7409,N_4498,N_3724);
nand U7410 (N_7410,N_2609,N_2261);
xor U7411 (N_7411,N_3495,N_4027);
or U7412 (N_7412,N_2666,N_3693);
or U7413 (N_7413,N_4254,N_3295);
xor U7414 (N_7414,N_2549,N_1632);
and U7415 (N_7415,N_3467,N_805);
xor U7416 (N_7416,N_986,N_4070);
and U7417 (N_7417,N_1606,N_4974);
nand U7418 (N_7418,N_3005,N_3948);
nor U7419 (N_7419,N_3698,N_3076);
or U7420 (N_7420,N_4019,N_317);
nand U7421 (N_7421,N_4956,N_1852);
xor U7422 (N_7422,N_4413,N_2658);
nor U7423 (N_7423,N_4768,N_467);
xor U7424 (N_7424,N_3247,N_3137);
nor U7425 (N_7425,N_3339,N_407);
nand U7426 (N_7426,N_833,N_2547);
xnor U7427 (N_7427,N_1537,N_4975);
nor U7428 (N_7428,N_4888,N_1837);
nand U7429 (N_7429,N_3910,N_4039);
or U7430 (N_7430,N_138,N_4988);
nor U7431 (N_7431,N_2691,N_2628);
nand U7432 (N_7432,N_693,N_1674);
nand U7433 (N_7433,N_2215,N_1589);
nand U7434 (N_7434,N_1688,N_1740);
nand U7435 (N_7435,N_3550,N_2141);
nand U7436 (N_7436,N_3778,N_4948);
xor U7437 (N_7437,N_1783,N_2120);
nand U7438 (N_7438,N_1933,N_2338);
nand U7439 (N_7439,N_1265,N_2114);
nand U7440 (N_7440,N_642,N_4636);
xor U7441 (N_7441,N_3477,N_4704);
nor U7442 (N_7442,N_3676,N_2526);
xnor U7443 (N_7443,N_1542,N_4396);
xnor U7444 (N_7444,N_2523,N_1646);
nor U7445 (N_7445,N_3897,N_1133);
and U7446 (N_7446,N_936,N_3986);
and U7447 (N_7447,N_1312,N_2834);
nor U7448 (N_7448,N_1354,N_1248);
or U7449 (N_7449,N_3578,N_3537);
nand U7450 (N_7450,N_2117,N_3367);
xnor U7451 (N_7451,N_602,N_2443);
nor U7452 (N_7452,N_2054,N_2212);
or U7453 (N_7453,N_893,N_2430);
or U7454 (N_7454,N_4787,N_445);
or U7455 (N_7455,N_127,N_1643);
nor U7456 (N_7456,N_1142,N_2485);
or U7457 (N_7457,N_3121,N_2116);
nor U7458 (N_7458,N_793,N_4172);
xor U7459 (N_7459,N_4198,N_3179);
xnor U7460 (N_7460,N_318,N_2993);
nor U7461 (N_7461,N_4612,N_757);
nor U7462 (N_7462,N_2862,N_1661);
and U7463 (N_7463,N_2334,N_1787);
and U7464 (N_7464,N_2684,N_527);
nor U7465 (N_7465,N_2913,N_158);
or U7466 (N_7466,N_1204,N_3717);
xor U7467 (N_7467,N_289,N_1100);
or U7468 (N_7468,N_1489,N_1585);
nand U7469 (N_7469,N_3347,N_526);
or U7470 (N_7470,N_925,N_3441);
nand U7471 (N_7471,N_4137,N_3773);
and U7472 (N_7472,N_169,N_3353);
and U7473 (N_7473,N_3520,N_502);
xnor U7474 (N_7474,N_1417,N_3096);
or U7475 (N_7475,N_2832,N_3146);
nand U7476 (N_7476,N_178,N_561);
nand U7477 (N_7477,N_2922,N_68);
and U7478 (N_7478,N_3432,N_3254);
or U7479 (N_7479,N_958,N_594);
or U7480 (N_7480,N_2296,N_2952);
nor U7481 (N_7481,N_233,N_1663);
and U7482 (N_7482,N_3903,N_1610);
nor U7483 (N_7483,N_4746,N_3366);
xnor U7484 (N_7484,N_436,N_3600);
nand U7485 (N_7485,N_985,N_2143);
or U7486 (N_7486,N_950,N_258);
xor U7487 (N_7487,N_4340,N_1211);
nand U7488 (N_7488,N_3440,N_1203);
and U7489 (N_7489,N_4344,N_3892);
nand U7490 (N_7490,N_1360,N_776);
nor U7491 (N_7491,N_3507,N_1536);
or U7492 (N_7492,N_4149,N_421);
xnor U7493 (N_7493,N_3789,N_1549);
or U7494 (N_7494,N_4542,N_4043);
and U7495 (N_7495,N_3251,N_575);
nor U7496 (N_7496,N_4129,N_1008);
or U7497 (N_7497,N_972,N_2851);
or U7498 (N_7498,N_78,N_4310);
and U7499 (N_7499,N_4399,N_1276);
nand U7500 (N_7500,N_765,N_4318);
nor U7501 (N_7501,N_2597,N_750);
nor U7502 (N_7502,N_2444,N_2156);
nor U7503 (N_7503,N_1616,N_1595);
nand U7504 (N_7504,N_4097,N_3544);
or U7505 (N_7505,N_2739,N_1338);
or U7506 (N_7506,N_2646,N_3996);
or U7507 (N_7507,N_3892,N_2440);
and U7508 (N_7508,N_1161,N_427);
nand U7509 (N_7509,N_1578,N_1901);
xor U7510 (N_7510,N_1337,N_3687);
nand U7511 (N_7511,N_1583,N_512);
nand U7512 (N_7512,N_2448,N_3221);
or U7513 (N_7513,N_2446,N_4241);
nor U7514 (N_7514,N_1966,N_1473);
and U7515 (N_7515,N_1159,N_3022);
nor U7516 (N_7516,N_4920,N_1383);
nor U7517 (N_7517,N_4200,N_1457);
nand U7518 (N_7518,N_3549,N_2056);
nand U7519 (N_7519,N_4258,N_2837);
xor U7520 (N_7520,N_2987,N_4461);
nor U7521 (N_7521,N_3314,N_1668);
or U7522 (N_7522,N_448,N_3558);
nand U7523 (N_7523,N_1252,N_1158);
or U7524 (N_7524,N_4021,N_997);
and U7525 (N_7525,N_1246,N_3018);
or U7526 (N_7526,N_216,N_341);
nor U7527 (N_7527,N_3211,N_3634);
xnor U7528 (N_7528,N_4090,N_4033);
or U7529 (N_7529,N_1006,N_4217);
and U7530 (N_7530,N_440,N_1357);
nor U7531 (N_7531,N_2820,N_4840);
and U7532 (N_7532,N_2230,N_2191);
or U7533 (N_7533,N_3430,N_4815);
or U7534 (N_7534,N_4692,N_3505);
and U7535 (N_7535,N_1108,N_3387);
or U7536 (N_7536,N_906,N_3057);
or U7537 (N_7537,N_3260,N_1748);
nand U7538 (N_7538,N_3907,N_557);
and U7539 (N_7539,N_4493,N_4762);
and U7540 (N_7540,N_4904,N_2391);
xor U7541 (N_7541,N_3913,N_2082);
and U7542 (N_7542,N_668,N_1386);
nand U7543 (N_7543,N_1995,N_4391);
nor U7544 (N_7544,N_3811,N_2496);
nand U7545 (N_7545,N_2588,N_2668);
nor U7546 (N_7546,N_3602,N_3162);
nand U7547 (N_7547,N_4353,N_4714);
xnor U7548 (N_7548,N_973,N_806);
nor U7549 (N_7549,N_4520,N_1580);
xor U7550 (N_7550,N_347,N_2841);
nand U7551 (N_7551,N_3850,N_2644);
nand U7552 (N_7552,N_407,N_3839);
nand U7553 (N_7553,N_3686,N_279);
or U7554 (N_7554,N_342,N_4318);
and U7555 (N_7555,N_2650,N_3298);
and U7556 (N_7556,N_4053,N_4691);
nor U7557 (N_7557,N_4759,N_3161);
nor U7558 (N_7558,N_2980,N_2189);
xor U7559 (N_7559,N_330,N_2102);
and U7560 (N_7560,N_3733,N_1819);
and U7561 (N_7561,N_452,N_3566);
and U7562 (N_7562,N_529,N_1726);
or U7563 (N_7563,N_2811,N_2939);
nand U7564 (N_7564,N_3200,N_2842);
nand U7565 (N_7565,N_2033,N_292);
and U7566 (N_7566,N_3615,N_4129);
nor U7567 (N_7567,N_2924,N_3115);
xor U7568 (N_7568,N_449,N_4769);
or U7569 (N_7569,N_1143,N_4209);
xnor U7570 (N_7570,N_4919,N_3629);
or U7571 (N_7571,N_1004,N_1893);
nor U7572 (N_7572,N_1677,N_3351);
nor U7573 (N_7573,N_1035,N_4178);
nand U7574 (N_7574,N_2762,N_290);
xor U7575 (N_7575,N_2099,N_2073);
xnor U7576 (N_7576,N_3071,N_1914);
xor U7577 (N_7577,N_3917,N_4849);
or U7578 (N_7578,N_1519,N_2235);
nand U7579 (N_7579,N_923,N_2402);
xor U7580 (N_7580,N_3468,N_3492);
nand U7581 (N_7581,N_1178,N_117);
xnor U7582 (N_7582,N_3438,N_509);
or U7583 (N_7583,N_3637,N_3769);
nand U7584 (N_7584,N_439,N_1040);
and U7585 (N_7585,N_866,N_119);
nor U7586 (N_7586,N_2004,N_2669);
nor U7587 (N_7587,N_4766,N_4295);
or U7588 (N_7588,N_2085,N_2861);
or U7589 (N_7589,N_1927,N_3874);
or U7590 (N_7590,N_1932,N_1056);
nand U7591 (N_7591,N_816,N_3132);
xnor U7592 (N_7592,N_275,N_4809);
nor U7593 (N_7593,N_3449,N_3740);
xor U7594 (N_7594,N_2194,N_3426);
or U7595 (N_7595,N_1459,N_4141);
and U7596 (N_7596,N_2373,N_3531);
xor U7597 (N_7597,N_1307,N_4420);
or U7598 (N_7598,N_3507,N_3453);
xnor U7599 (N_7599,N_4013,N_3797);
nand U7600 (N_7600,N_1411,N_3167);
nor U7601 (N_7601,N_1692,N_3876);
and U7602 (N_7602,N_1671,N_2727);
nand U7603 (N_7603,N_1446,N_977);
or U7604 (N_7604,N_149,N_582);
nor U7605 (N_7605,N_2987,N_616);
nand U7606 (N_7606,N_1535,N_4472);
and U7607 (N_7607,N_4509,N_820);
or U7608 (N_7608,N_3927,N_1442);
or U7609 (N_7609,N_4311,N_2579);
nand U7610 (N_7610,N_2874,N_3851);
nor U7611 (N_7611,N_1532,N_111);
and U7612 (N_7612,N_1308,N_1325);
or U7613 (N_7613,N_3084,N_3132);
nor U7614 (N_7614,N_972,N_3044);
nor U7615 (N_7615,N_1346,N_3750);
nor U7616 (N_7616,N_1728,N_3167);
nor U7617 (N_7617,N_4940,N_383);
and U7618 (N_7618,N_1935,N_237);
and U7619 (N_7619,N_3237,N_3803);
or U7620 (N_7620,N_1976,N_2363);
nor U7621 (N_7621,N_4232,N_2784);
nor U7622 (N_7622,N_2658,N_2512);
and U7623 (N_7623,N_1879,N_4354);
or U7624 (N_7624,N_4801,N_3982);
and U7625 (N_7625,N_158,N_652);
nor U7626 (N_7626,N_2532,N_4649);
nor U7627 (N_7627,N_2018,N_2341);
and U7628 (N_7628,N_671,N_4011);
nand U7629 (N_7629,N_1188,N_1530);
nor U7630 (N_7630,N_2118,N_2599);
nand U7631 (N_7631,N_814,N_3848);
and U7632 (N_7632,N_1701,N_4969);
nor U7633 (N_7633,N_3535,N_4555);
nand U7634 (N_7634,N_805,N_1483);
or U7635 (N_7635,N_2998,N_3073);
or U7636 (N_7636,N_973,N_3429);
nor U7637 (N_7637,N_66,N_4340);
and U7638 (N_7638,N_4959,N_4695);
nand U7639 (N_7639,N_2445,N_1749);
nand U7640 (N_7640,N_2253,N_2161);
and U7641 (N_7641,N_3160,N_174);
nor U7642 (N_7642,N_3977,N_2743);
xnor U7643 (N_7643,N_2707,N_3142);
or U7644 (N_7644,N_219,N_2687);
nor U7645 (N_7645,N_3322,N_4713);
or U7646 (N_7646,N_4253,N_2339);
and U7647 (N_7647,N_165,N_1107);
xor U7648 (N_7648,N_716,N_1751);
nand U7649 (N_7649,N_114,N_2294);
nand U7650 (N_7650,N_175,N_2197);
nand U7651 (N_7651,N_3137,N_2037);
nand U7652 (N_7652,N_2186,N_3386);
nand U7653 (N_7653,N_2294,N_1635);
nor U7654 (N_7654,N_1460,N_2933);
xnor U7655 (N_7655,N_4112,N_601);
or U7656 (N_7656,N_3760,N_2357);
or U7657 (N_7657,N_4038,N_4678);
and U7658 (N_7658,N_1476,N_118);
nand U7659 (N_7659,N_1220,N_3695);
or U7660 (N_7660,N_1489,N_1251);
nor U7661 (N_7661,N_517,N_1968);
nand U7662 (N_7662,N_27,N_3999);
and U7663 (N_7663,N_2445,N_787);
xor U7664 (N_7664,N_268,N_2056);
and U7665 (N_7665,N_4915,N_999);
or U7666 (N_7666,N_3819,N_650);
and U7667 (N_7667,N_3859,N_4643);
or U7668 (N_7668,N_3105,N_4075);
xnor U7669 (N_7669,N_1308,N_3376);
xnor U7670 (N_7670,N_3386,N_4217);
and U7671 (N_7671,N_2018,N_4010);
and U7672 (N_7672,N_3738,N_3317);
or U7673 (N_7673,N_2367,N_684);
nor U7674 (N_7674,N_280,N_3172);
xnor U7675 (N_7675,N_1569,N_4980);
xnor U7676 (N_7676,N_213,N_1617);
or U7677 (N_7677,N_2834,N_3053);
nor U7678 (N_7678,N_3777,N_2582);
or U7679 (N_7679,N_3334,N_1502);
and U7680 (N_7680,N_238,N_1932);
nor U7681 (N_7681,N_1056,N_3210);
xor U7682 (N_7682,N_4864,N_4727);
nor U7683 (N_7683,N_1553,N_1612);
or U7684 (N_7684,N_1307,N_2130);
nand U7685 (N_7685,N_611,N_1346);
and U7686 (N_7686,N_476,N_146);
nor U7687 (N_7687,N_484,N_1926);
or U7688 (N_7688,N_3302,N_4950);
xnor U7689 (N_7689,N_692,N_2879);
or U7690 (N_7690,N_3298,N_4229);
nand U7691 (N_7691,N_3799,N_4479);
and U7692 (N_7692,N_2125,N_320);
and U7693 (N_7693,N_3975,N_4766);
xor U7694 (N_7694,N_4710,N_470);
or U7695 (N_7695,N_1303,N_3065);
and U7696 (N_7696,N_778,N_2802);
nand U7697 (N_7697,N_2599,N_899);
nor U7698 (N_7698,N_4043,N_1749);
or U7699 (N_7699,N_4196,N_4443);
nor U7700 (N_7700,N_4575,N_4339);
nor U7701 (N_7701,N_4208,N_684);
xor U7702 (N_7702,N_916,N_2156);
xnor U7703 (N_7703,N_367,N_3497);
or U7704 (N_7704,N_3048,N_3506);
nand U7705 (N_7705,N_3531,N_1394);
and U7706 (N_7706,N_1463,N_2446);
nor U7707 (N_7707,N_2875,N_3323);
or U7708 (N_7708,N_1689,N_2011);
xnor U7709 (N_7709,N_1689,N_4770);
xor U7710 (N_7710,N_1943,N_392);
nand U7711 (N_7711,N_1261,N_209);
nand U7712 (N_7712,N_2446,N_3443);
xor U7713 (N_7713,N_4184,N_3468);
xor U7714 (N_7714,N_750,N_4969);
or U7715 (N_7715,N_2470,N_403);
and U7716 (N_7716,N_3772,N_2434);
and U7717 (N_7717,N_1735,N_4928);
nand U7718 (N_7718,N_3358,N_891);
nand U7719 (N_7719,N_134,N_4764);
nor U7720 (N_7720,N_3925,N_2299);
xor U7721 (N_7721,N_1096,N_3571);
or U7722 (N_7722,N_1245,N_1074);
or U7723 (N_7723,N_2083,N_2636);
and U7724 (N_7724,N_3631,N_1982);
and U7725 (N_7725,N_4565,N_1441);
nand U7726 (N_7726,N_1491,N_2298);
nand U7727 (N_7727,N_3088,N_2640);
nand U7728 (N_7728,N_522,N_905);
xor U7729 (N_7729,N_406,N_1119);
and U7730 (N_7730,N_1893,N_1344);
and U7731 (N_7731,N_3451,N_2694);
nor U7732 (N_7732,N_77,N_2386);
or U7733 (N_7733,N_1610,N_1811);
and U7734 (N_7734,N_4581,N_4118);
or U7735 (N_7735,N_1186,N_3810);
nand U7736 (N_7736,N_3150,N_4715);
and U7737 (N_7737,N_4265,N_4109);
and U7738 (N_7738,N_782,N_1705);
xnor U7739 (N_7739,N_2161,N_3357);
xnor U7740 (N_7740,N_1064,N_584);
xor U7741 (N_7741,N_2256,N_1768);
xnor U7742 (N_7742,N_4290,N_398);
and U7743 (N_7743,N_4452,N_2294);
or U7744 (N_7744,N_4624,N_1436);
nand U7745 (N_7745,N_4191,N_2972);
nor U7746 (N_7746,N_2743,N_3148);
xnor U7747 (N_7747,N_1428,N_3058);
xnor U7748 (N_7748,N_616,N_3293);
or U7749 (N_7749,N_417,N_1751);
nand U7750 (N_7750,N_1511,N_3189);
nor U7751 (N_7751,N_4885,N_204);
nor U7752 (N_7752,N_203,N_1554);
or U7753 (N_7753,N_3131,N_1787);
nor U7754 (N_7754,N_3217,N_2987);
xor U7755 (N_7755,N_1673,N_4579);
and U7756 (N_7756,N_1038,N_3091);
xnor U7757 (N_7757,N_477,N_4520);
xnor U7758 (N_7758,N_1370,N_4836);
nand U7759 (N_7759,N_3352,N_2573);
or U7760 (N_7760,N_1362,N_2655);
nor U7761 (N_7761,N_3635,N_2523);
and U7762 (N_7762,N_2185,N_3326);
and U7763 (N_7763,N_2148,N_2943);
nand U7764 (N_7764,N_3286,N_168);
or U7765 (N_7765,N_4648,N_2105);
nand U7766 (N_7766,N_3152,N_2702);
or U7767 (N_7767,N_3658,N_3260);
nand U7768 (N_7768,N_968,N_451);
nor U7769 (N_7769,N_454,N_3972);
or U7770 (N_7770,N_1069,N_2718);
xnor U7771 (N_7771,N_3851,N_829);
or U7772 (N_7772,N_4001,N_1732);
nor U7773 (N_7773,N_1439,N_2933);
nand U7774 (N_7774,N_1507,N_4931);
and U7775 (N_7775,N_2823,N_3925);
and U7776 (N_7776,N_2959,N_2562);
or U7777 (N_7777,N_3867,N_1004);
nand U7778 (N_7778,N_4932,N_1066);
nand U7779 (N_7779,N_2059,N_3075);
nor U7780 (N_7780,N_3685,N_1565);
xor U7781 (N_7781,N_1566,N_1572);
nor U7782 (N_7782,N_1741,N_918);
or U7783 (N_7783,N_481,N_3121);
nor U7784 (N_7784,N_4266,N_3330);
nor U7785 (N_7785,N_4876,N_4772);
and U7786 (N_7786,N_2248,N_4207);
nand U7787 (N_7787,N_2884,N_709);
nor U7788 (N_7788,N_1643,N_4072);
nor U7789 (N_7789,N_3414,N_3154);
nor U7790 (N_7790,N_4131,N_3344);
or U7791 (N_7791,N_3489,N_4958);
nand U7792 (N_7792,N_1879,N_3685);
and U7793 (N_7793,N_4873,N_622);
and U7794 (N_7794,N_4019,N_1724);
or U7795 (N_7795,N_28,N_3681);
nor U7796 (N_7796,N_3547,N_2185);
xor U7797 (N_7797,N_4293,N_639);
and U7798 (N_7798,N_407,N_1216);
or U7799 (N_7799,N_2463,N_77);
nor U7800 (N_7800,N_2402,N_704);
or U7801 (N_7801,N_1057,N_2585);
or U7802 (N_7802,N_1984,N_4458);
and U7803 (N_7803,N_4604,N_4533);
and U7804 (N_7804,N_4861,N_89);
nand U7805 (N_7805,N_3091,N_4434);
nor U7806 (N_7806,N_1140,N_1959);
nor U7807 (N_7807,N_4593,N_3428);
xnor U7808 (N_7808,N_2337,N_1607);
or U7809 (N_7809,N_2106,N_4260);
nor U7810 (N_7810,N_2410,N_1546);
nor U7811 (N_7811,N_4936,N_2482);
and U7812 (N_7812,N_3777,N_4785);
and U7813 (N_7813,N_3447,N_4845);
and U7814 (N_7814,N_3741,N_2020);
or U7815 (N_7815,N_3469,N_3279);
nor U7816 (N_7816,N_2064,N_3465);
and U7817 (N_7817,N_2212,N_534);
xor U7818 (N_7818,N_4225,N_4691);
and U7819 (N_7819,N_99,N_4123);
or U7820 (N_7820,N_3655,N_3824);
xnor U7821 (N_7821,N_507,N_4798);
xnor U7822 (N_7822,N_3567,N_344);
nand U7823 (N_7823,N_2319,N_1593);
and U7824 (N_7824,N_1439,N_1306);
nand U7825 (N_7825,N_2496,N_4538);
or U7826 (N_7826,N_127,N_3167);
xor U7827 (N_7827,N_1853,N_1314);
xnor U7828 (N_7828,N_1940,N_3062);
xor U7829 (N_7829,N_568,N_2173);
or U7830 (N_7830,N_1343,N_3277);
nor U7831 (N_7831,N_3290,N_942);
nand U7832 (N_7832,N_376,N_2773);
xor U7833 (N_7833,N_4284,N_2497);
xnor U7834 (N_7834,N_3910,N_3117);
xor U7835 (N_7835,N_1234,N_1341);
or U7836 (N_7836,N_2676,N_290);
xnor U7837 (N_7837,N_1467,N_3274);
nand U7838 (N_7838,N_3025,N_672);
xnor U7839 (N_7839,N_3600,N_1782);
or U7840 (N_7840,N_1641,N_1936);
nand U7841 (N_7841,N_2958,N_2288);
nor U7842 (N_7842,N_2226,N_4209);
and U7843 (N_7843,N_4795,N_611);
xnor U7844 (N_7844,N_267,N_3215);
and U7845 (N_7845,N_961,N_3823);
and U7846 (N_7846,N_3231,N_1305);
and U7847 (N_7847,N_4866,N_3551);
nand U7848 (N_7848,N_4964,N_1659);
nor U7849 (N_7849,N_217,N_4025);
nor U7850 (N_7850,N_3055,N_3238);
nand U7851 (N_7851,N_3539,N_1733);
nand U7852 (N_7852,N_433,N_3544);
or U7853 (N_7853,N_3058,N_4156);
xor U7854 (N_7854,N_3704,N_621);
nand U7855 (N_7855,N_1183,N_3243);
nor U7856 (N_7856,N_3578,N_2471);
and U7857 (N_7857,N_1628,N_2200);
nand U7858 (N_7858,N_4456,N_4820);
nor U7859 (N_7859,N_3287,N_4442);
and U7860 (N_7860,N_93,N_1749);
and U7861 (N_7861,N_3429,N_473);
or U7862 (N_7862,N_2704,N_445);
and U7863 (N_7863,N_254,N_4995);
and U7864 (N_7864,N_855,N_371);
nand U7865 (N_7865,N_4953,N_4998);
xnor U7866 (N_7866,N_434,N_3040);
nor U7867 (N_7867,N_651,N_823);
or U7868 (N_7868,N_3771,N_2847);
nand U7869 (N_7869,N_2301,N_4128);
nand U7870 (N_7870,N_1927,N_2298);
or U7871 (N_7871,N_1681,N_1603);
nand U7872 (N_7872,N_751,N_3982);
nand U7873 (N_7873,N_4298,N_1178);
nor U7874 (N_7874,N_881,N_3909);
xor U7875 (N_7875,N_3126,N_109);
nand U7876 (N_7876,N_1951,N_3603);
nand U7877 (N_7877,N_4452,N_1592);
xor U7878 (N_7878,N_4903,N_3729);
nor U7879 (N_7879,N_4940,N_4753);
nand U7880 (N_7880,N_2522,N_2452);
or U7881 (N_7881,N_2487,N_1382);
nor U7882 (N_7882,N_2656,N_1867);
or U7883 (N_7883,N_3779,N_2494);
and U7884 (N_7884,N_389,N_3547);
or U7885 (N_7885,N_3489,N_2857);
or U7886 (N_7886,N_1545,N_3701);
or U7887 (N_7887,N_907,N_3383);
xor U7888 (N_7888,N_4971,N_4193);
nand U7889 (N_7889,N_2779,N_816);
and U7890 (N_7890,N_4696,N_4513);
or U7891 (N_7891,N_1891,N_4144);
nor U7892 (N_7892,N_4973,N_1368);
nand U7893 (N_7893,N_3127,N_4504);
or U7894 (N_7894,N_2670,N_1986);
and U7895 (N_7895,N_1519,N_2739);
nand U7896 (N_7896,N_2295,N_3479);
nor U7897 (N_7897,N_38,N_2971);
nor U7898 (N_7898,N_2344,N_3856);
or U7899 (N_7899,N_280,N_3885);
nor U7900 (N_7900,N_4928,N_468);
xor U7901 (N_7901,N_1194,N_564);
or U7902 (N_7902,N_4198,N_551);
and U7903 (N_7903,N_527,N_4514);
and U7904 (N_7904,N_4970,N_3573);
and U7905 (N_7905,N_4587,N_950);
and U7906 (N_7906,N_4971,N_2917);
nand U7907 (N_7907,N_57,N_363);
nor U7908 (N_7908,N_3622,N_2032);
xor U7909 (N_7909,N_1826,N_2160);
xor U7910 (N_7910,N_683,N_2677);
or U7911 (N_7911,N_2071,N_3171);
and U7912 (N_7912,N_698,N_3060);
and U7913 (N_7913,N_4161,N_4582);
and U7914 (N_7914,N_721,N_4374);
or U7915 (N_7915,N_2317,N_4814);
xor U7916 (N_7916,N_3680,N_4507);
nand U7917 (N_7917,N_2227,N_2236);
or U7918 (N_7918,N_149,N_1854);
xnor U7919 (N_7919,N_2550,N_281);
xor U7920 (N_7920,N_1731,N_365);
or U7921 (N_7921,N_3446,N_2899);
or U7922 (N_7922,N_843,N_4901);
xor U7923 (N_7923,N_3028,N_4028);
or U7924 (N_7924,N_3966,N_2119);
xnor U7925 (N_7925,N_1027,N_1937);
xor U7926 (N_7926,N_467,N_2134);
xnor U7927 (N_7927,N_2140,N_1170);
and U7928 (N_7928,N_2002,N_3237);
nand U7929 (N_7929,N_152,N_3726);
and U7930 (N_7930,N_1758,N_4256);
and U7931 (N_7931,N_3956,N_2518);
and U7932 (N_7932,N_4309,N_3512);
nor U7933 (N_7933,N_4194,N_2223);
nor U7934 (N_7934,N_3450,N_1413);
xor U7935 (N_7935,N_3693,N_2916);
xor U7936 (N_7936,N_4810,N_3466);
xnor U7937 (N_7937,N_129,N_2842);
nor U7938 (N_7938,N_2826,N_3869);
nand U7939 (N_7939,N_18,N_3347);
or U7940 (N_7940,N_4992,N_4338);
and U7941 (N_7941,N_4886,N_195);
nand U7942 (N_7942,N_3999,N_4401);
or U7943 (N_7943,N_4553,N_655);
nand U7944 (N_7944,N_440,N_4528);
xnor U7945 (N_7945,N_1283,N_4713);
or U7946 (N_7946,N_1075,N_4274);
nor U7947 (N_7947,N_3598,N_3037);
or U7948 (N_7948,N_4172,N_129);
and U7949 (N_7949,N_4929,N_2970);
xor U7950 (N_7950,N_4323,N_1842);
nor U7951 (N_7951,N_2537,N_3363);
nor U7952 (N_7952,N_1298,N_2114);
nor U7953 (N_7953,N_338,N_4296);
xor U7954 (N_7954,N_2042,N_3525);
nand U7955 (N_7955,N_4556,N_1997);
or U7956 (N_7956,N_3811,N_3548);
and U7957 (N_7957,N_3792,N_3622);
and U7958 (N_7958,N_631,N_414);
or U7959 (N_7959,N_1745,N_3228);
and U7960 (N_7960,N_448,N_806);
nand U7961 (N_7961,N_184,N_2445);
nand U7962 (N_7962,N_2194,N_3562);
nor U7963 (N_7963,N_4570,N_1905);
nor U7964 (N_7964,N_3360,N_1358);
nand U7965 (N_7965,N_2733,N_4022);
nand U7966 (N_7966,N_4171,N_846);
xnor U7967 (N_7967,N_3234,N_1281);
xnor U7968 (N_7968,N_1946,N_3310);
nor U7969 (N_7969,N_1870,N_1576);
nand U7970 (N_7970,N_3606,N_4283);
nor U7971 (N_7971,N_1699,N_558);
and U7972 (N_7972,N_3441,N_1826);
nand U7973 (N_7973,N_3309,N_1345);
nand U7974 (N_7974,N_1661,N_4224);
or U7975 (N_7975,N_4899,N_4020);
xor U7976 (N_7976,N_2742,N_4785);
xnor U7977 (N_7977,N_2120,N_483);
or U7978 (N_7978,N_4135,N_3134);
and U7979 (N_7979,N_1154,N_4443);
nor U7980 (N_7980,N_3962,N_3729);
and U7981 (N_7981,N_2293,N_3836);
nand U7982 (N_7982,N_1596,N_4970);
xnor U7983 (N_7983,N_480,N_2638);
or U7984 (N_7984,N_1956,N_112);
nor U7985 (N_7985,N_1914,N_3959);
nand U7986 (N_7986,N_3806,N_1919);
and U7987 (N_7987,N_3878,N_2264);
and U7988 (N_7988,N_1728,N_4427);
nand U7989 (N_7989,N_1060,N_4963);
nor U7990 (N_7990,N_614,N_1469);
nor U7991 (N_7991,N_306,N_4910);
nand U7992 (N_7992,N_2475,N_451);
or U7993 (N_7993,N_1678,N_130);
nor U7994 (N_7994,N_1571,N_3899);
nor U7995 (N_7995,N_1027,N_3716);
or U7996 (N_7996,N_2441,N_487);
nand U7997 (N_7997,N_1392,N_2387);
xnor U7998 (N_7998,N_4857,N_1483);
and U7999 (N_7999,N_1678,N_2041);
nor U8000 (N_8000,N_2807,N_2210);
nor U8001 (N_8001,N_1434,N_4156);
or U8002 (N_8002,N_2087,N_113);
and U8003 (N_8003,N_3364,N_4798);
and U8004 (N_8004,N_2326,N_3989);
and U8005 (N_8005,N_4009,N_4377);
nand U8006 (N_8006,N_4711,N_4628);
and U8007 (N_8007,N_1851,N_4551);
or U8008 (N_8008,N_28,N_1388);
nand U8009 (N_8009,N_3222,N_3400);
or U8010 (N_8010,N_2824,N_3253);
xor U8011 (N_8011,N_3210,N_3978);
nor U8012 (N_8012,N_1206,N_715);
nor U8013 (N_8013,N_4776,N_1322);
or U8014 (N_8014,N_1365,N_266);
nand U8015 (N_8015,N_1227,N_2082);
xnor U8016 (N_8016,N_3611,N_4874);
xnor U8017 (N_8017,N_3370,N_479);
nand U8018 (N_8018,N_2160,N_441);
and U8019 (N_8019,N_1727,N_3432);
nand U8020 (N_8020,N_4584,N_3961);
nor U8021 (N_8021,N_3067,N_3854);
nand U8022 (N_8022,N_671,N_1116);
nand U8023 (N_8023,N_3684,N_3386);
and U8024 (N_8024,N_1839,N_2069);
nand U8025 (N_8025,N_1721,N_4169);
nand U8026 (N_8026,N_3020,N_2174);
nand U8027 (N_8027,N_1075,N_301);
and U8028 (N_8028,N_1262,N_2934);
and U8029 (N_8029,N_917,N_3730);
or U8030 (N_8030,N_1560,N_3530);
nand U8031 (N_8031,N_2190,N_3420);
nor U8032 (N_8032,N_2368,N_4155);
nand U8033 (N_8033,N_10,N_3857);
or U8034 (N_8034,N_1961,N_3285);
xor U8035 (N_8035,N_4831,N_1320);
and U8036 (N_8036,N_1855,N_2515);
or U8037 (N_8037,N_3347,N_3568);
xor U8038 (N_8038,N_2959,N_2659);
nor U8039 (N_8039,N_2104,N_1315);
or U8040 (N_8040,N_616,N_329);
nor U8041 (N_8041,N_3216,N_2117);
nand U8042 (N_8042,N_678,N_2895);
nor U8043 (N_8043,N_2003,N_2752);
or U8044 (N_8044,N_2394,N_1634);
nand U8045 (N_8045,N_1719,N_2497);
nor U8046 (N_8046,N_4275,N_2607);
nor U8047 (N_8047,N_2651,N_1955);
or U8048 (N_8048,N_54,N_3985);
nand U8049 (N_8049,N_4815,N_2919);
and U8050 (N_8050,N_4014,N_2550);
or U8051 (N_8051,N_1539,N_4575);
nor U8052 (N_8052,N_1467,N_2175);
nand U8053 (N_8053,N_1792,N_856);
nor U8054 (N_8054,N_4714,N_4800);
nand U8055 (N_8055,N_3807,N_3850);
nor U8056 (N_8056,N_4893,N_3970);
xor U8057 (N_8057,N_2866,N_3573);
nand U8058 (N_8058,N_1498,N_3072);
or U8059 (N_8059,N_1042,N_2431);
xnor U8060 (N_8060,N_3134,N_4168);
xor U8061 (N_8061,N_3268,N_1636);
xnor U8062 (N_8062,N_84,N_2263);
or U8063 (N_8063,N_764,N_1590);
nand U8064 (N_8064,N_4128,N_1320);
or U8065 (N_8065,N_4712,N_3484);
nor U8066 (N_8066,N_2343,N_16);
and U8067 (N_8067,N_4,N_2104);
and U8068 (N_8068,N_1930,N_173);
nand U8069 (N_8069,N_3815,N_2898);
and U8070 (N_8070,N_1933,N_1955);
and U8071 (N_8071,N_3208,N_1159);
nand U8072 (N_8072,N_2983,N_1707);
nand U8073 (N_8073,N_4390,N_4626);
nor U8074 (N_8074,N_1880,N_3526);
nor U8075 (N_8075,N_171,N_2676);
or U8076 (N_8076,N_3114,N_4827);
nand U8077 (N_8077,N_3480,N_1217);
nor U8078 (N_8078,N_4529,N_4135);
nor U8079 (N_8079,N_189,N_1124);
nor U8080 (N_8080,N_1752,N_3099);
nor U8081 (N_8081,N_775,N_598);
or U8082 (N_8082,N_1612,N_2588);
and U8083 (N_8083,N_2597,N_636);
nand U8084 (N_8084,N_4388,N_2511);
and U8085 (N_8085,N_2539,N_959);
and U8086 (N_8086,N_4214,N_3188);
or U8087 (N_8087,N_2838,N_2595);
xor U8088 (N_8088,N_3608,N_204);
nand U8089 (N_8089,N_1642,N_1746);
and U8090 (N_8090,N_2335,N_4675);
and U8091 (N_8091,N_3576,N_1778);
or U8092 (N_8092,N_4853,N_4138);
xor U8093 (N_8093,N_398,N_4922);
and U8094 (N_8094,N_1243,N_160);
nand U8095 (N_8095,N_1641,N_788);
or U8096 (N_8096,N_2545,N_3510);
xnor U8097 (N_8097,N_3034,N_4643);
xor U8098 (N_8098,N_929,N_4357);
and U8099 (N_8099,N_4181,N_3537);
nand U8100 (N_8100,N_600,N_3552);
xnor U8101 (N_8101,N_3941,N_3874);
nand U8102 (N_8102,N_420,N_2214);
and U8103 (N_8103,N_3822,N_2168);
or U8104 (N_8104,N_1480,N_2127);
xnor U8105 (N_8105,N_1323,N_1102);
or U8106 (N_8106,N_2194,N_4624);
nand U8107 (N_8107,N_3414,N_2905);
xnor U8108 (N_8108,N_731,N_1050);
nor U8109 (N_8109,N_2610,N_3713);
and U8110 (N_8110,N_781,N_1531);
nand U8111 (N_8111,N_3675,N_3795);
nor U8112 (N_8112,N_4639,N_3514);
and U8113 (N_8113,N_3817,N_1007);
and U8114 (N_8114,N_3897,N_3940);
xnor U8115 (N_8115,N_1516,N_4660);
xor U8116 (N_8116,N_2450,N_726);
and U8117 (N_8117,N_2759,N_1279);
nand U8118 (N_8118,N_1749,N_945);
or U8119 (N_8119,N_3349,N_1142);
nor U8120 (N_8120,N_2844,N_3669);
nor U8121 (N_8121,N_476,N_1126);
nand U8122 (N_8122,N_690,N_2892);
nand U8123 (N_8123,N_4801,N_3924);
xor U8124 (N_8124,N_3644,N_35);
xor U8125 (N_8125,N_48,N_3918);
xor U8126 (N_8126,N_4258,N_1712);
nor U8127 (N_8127,N_1842,N_1601);
and U8128 (N_8128,N_1968,N_1753);
or U8129 (N_8129,N_193,N_4735);
and U8130 (N_8130,N_944,N_2443);
or U8131 (N_8131,N_4929,N_4554);
and U8132 (N_8132,N_1634,N_2487);
xor U8133 (N_8133,N_462,N_4031);
nor U8134 (N_8134,N_887,N_3046);
nor U8135 (N_8135,N_3948,N_332);
and U8136 (N_8136,N_1679,N_2988);
or U8137 (N_8137,N_4827,N_3127);
and U8138 (N_8138,N_1373,N_281);
or U8139 (N_8139,N_1932,N_3487);
or U8140 (N_8140,N_199,N_1606);
xor U8141 (N_8141,N_3271,N_4598);
nand U8142 (N_8142,N_4585,N_4900);
nand U8143 (N_8143,N_666,N_1708);
or U8144 (N_8144,N_2084,N_2833);
nand U8145 (N_8145,N_3050,N_1058);
or U8146 (N_8146,N_149,N_2513);
nor U8147 (N_8147,N_3339,N_3442);
or U8148 (N_8148,N_2125,N_2645);
nand U8149 (N_8149,N_783,N_3399);
nand U8150 (N_8150,N_2618,N_1503);
nor U8151 (N_8151,N_4294,N_606);
or U8152 (N_8152,N_147,N_3490);
nand U8153 (N_8153,N_4763,N_3306);
nand U8154 (N_8154,N_2561,N_2804);
and U8155 (N_8155,N_2314,N_1334);
nand U8156 (N_8156,N_4989,N_4378);
xnor U8157 (N_8157,N_3539,N_1600);
nand U8158 (N_8158,N_3480,N_580);
and U8159 (N_8159,N_865,N_967);
and U8160 (N_8160,N_4614,N_4117);
nand U8161 (N_8161,N_2319,N_3891);
and U8162 (N_8162,N_1092,N_3535);
xnor U8163 (N_8163,N_1584,N_249);
xnor U8164 (N_8164,N_4448,N_2183);
nor U8165 (N_8165,N_4874,N_2355);
nor U8166 (N_8166,N_978,N_1016);
or U8167 (N_8167,N_3766,N_671);
and U8168 (N_8168,N_3635,N_588);
xor U8169 (N_8169,N_1876,N_4645);
xor U8170 (N_8170,N_1739,N_671);
and U8171 (N_8171,N_68,N_1259);
nand U8172 (N_8172,N_2831,N_4255);
and U8173 (N_8173,N_2841,N_4826);
and U8174 (N_8174,N_3464,N_174);
and U8175 (N_8175,N_501,N_349);
nand U8176 (N_8176,N_2086,N_1770);
xor U8177 (N_8177,N_3529,N_568);
and U8178 (N_8178,N_1187,N_3168);
nor U8179 (N_8179,N_1148,N_2690);
nor U8180 (N_8180,N_205,N_2012);
and U8181 (N_8181,N_4290,N_2406);
or U8182 (N_8182,N_1375,N_2163);
or U8183 (N_8183,N_3445,N_4067);
or U8184 (N_8184,N_567,N_1451);
and U8185 (N_8185,N_1277,N_866);
or U8186 (N_8186,N_647,N_3441);
nand U8187 (N_8187,N_915,N_380);
nor U8188 (N_8188,N_4143,N_3953);
nor U8189 (N_8189,N_4074,N_508);
nand U8190 (N_8190,N_3043,N_907);
and U8191 (N_8191,N_2766,N_1003);
xnor U8192 (N_8192,N_201,N_2689);
and U8193 (N_8193,N_455,N_2992);
nor U8194 (N_8194,N_4606,N_4422);
or U8195 (N_8195,N_312,N_4749);
nor U8196 (N_8196,N_4877,N_4229);
nor U8197 (N_8197,N_3237,N_288);
nand U8198 (N_8198,N_1757,N_3822);
and U8199 (N_8199,N_3058,N_2471);
nand U8200 (N_8200,N_42,N_2753);
xnor U8201 (N_8201,N_30,N_4134);
nand U8202 (N_8202,N_426,N_4800);
nand U8203 (N_8203,N_3017,N_1530);
nor U8204 (N_8204,N_451,N_4337);
or U8205 (N_8205,N_626,N_4046);
and U8206 (N_8206,N_1278,N_1641);
nand U8207 (N_8207,N_3408,N_3316);
nor U8208 (N_8208,N_1896,N_3814);
and U8209 (N_8209,N_2535,N_3487);
or U8210 (N_8210,N_3410,N_3385);
nor U8211 (N_8211,N_2597,N_3529);
nor U8212 (N_8212,N_3572,N_3397);
nor U8213 (N_8213,N_4926,N_2561);
nand U8214 (N_8214,N_3368,N_711);
nor U8215 (N_8215,N_955,N_2051);
or U8216 (N_8216,N_1666,N_560);
and U8217 (N_8217,N_102,N_3867);
nor U8218 (N_8218,N_2976,N_4098);
xnor U8219 (N_8219,N_4800,N_915);
nand U8220 (N_8220,N_4250,N_4579);
and U8221 (N_8221,N_2188,N_8);
and U8222 (N_8222,N_4584,N_161);
or U8223 (N_8223,N_355,N_2556);
or U8224 (N_8224,N_2990,N_4991);
nor U8225 (N_8225,N_422,N_4507);
xor U8226 (N_8226,N_3966,N_2457);
nand U8227 (N_8227,N_2190,N_486);
or U8228 (N_8228,N_1351,N_4923);
or U8229 (N_8229,N_3699,N_1340);
or U8230 (N_8230,N_4701,N_2166);
or U8231 (N_8231,N_3707,N_3663);
nand U8232 (N_8232,N_1665,N_2150);
xor U8233 (N_8233,N_3760,N_3768);
nor U8234 (N_8234,N_1770,N_1093);
or U8235 (N_8235,N_2021,N_26);
or U8236 (N_8236,N_2704,N_3496);
xnor U8237 (N_8237,N_1240,N_1530);
and U8238 (N_8238,N_4532,N_4613);
nand U8239 (N_8239,N_3699,N_654);
nor U8240 (N_8240,N_2920,N_1217);
or U8241 (N_8241,N_3910,N_1955);
or U8242 (N_8242,N_3113,N_2298);
nor U8243 (N_8243,N_4464,N_1715);
and U8244 (N_8244,N_4093,N_4587);
nor U8245 (N_8245,N_4453,N_4210);
nor U8246 (N_8246,N_1351,N_2671);
and U8247 (N_8247,N_3708,N_2232);
xor U8248 (N_8248,N_4713,N_1724);
xnor U8249 (N_8249,N_4954,N_1120);
nand U8250 (N_8250,N_885,N_4237);
xor U8251 (N_8251,N_2144,N_3380);
xor U8252 (N_8252,N_1241,N_4306);
nand U8253 (N_8253,N_410,N_2663);
nor U8254 (N_8254,N_4927,N_4616);
nand U8255 (N_8255,N_3132,N_3905);
or U8256 (N_8256,N_4131,N_2844);
and U8257 (N_8257,N_955,N_4593);
or U8258 (N_8258,N_1169,N_541);
nor U8259 (N_8259,N_2936,N_3331);
nand U8260 (N_8260,N_3246,N_658);
nand U8261 (N_8261,N_1451,N_1883);
xnor U8262 (N_8262,N_839,N_2230);
or U8263 (N_8263,N_3680,N_2514);
xnor U8264 (N_8264,N_2919,N_2089);
nand U8265 (N_8265,N_988,N_1182);
or U8266 (N_8266,N_3245,N_3914);
nand U8267 (N_8267,N_2932,N_2900);
or U8268 (N_8268,N_2887,N_3192);
nand U8269 (N_8269,N_2477,N_2669);
nand U8270 (N_8270,N_3580,N_3999);
xor U8271 (N_8271,N_2332,N_2014);
nor U8272 (N_8272,N_3944,N_3684);
or U8273 (N_8273,N_2301,N_2191);
xor U8274 (N_8274,N_2171,N_2225);
nor U8275 (N_8275,N_2011,N_1892);
xor U8276 (N_8276,N_487,N_3628);
or U8277 (N_8277,N_384,N_2653);
nand U8278 (N_8278,N_4357,N_3851);
nand U8279 (N_8279,N_2777,N_1722);
and U8280 (N_8280,N_3916,N_601);
nor U8281 (N_8281,N_2933,N_3560);
nor U8282 (N_8282,N_2508,N_4689);
or U8283 (N_8283,N_3928,N_4038);
or U8284 (N_8284,N_3167,N_702);
or U8285 (N_8285,N_3278,N_4130);
nand U8286 (N_8286,N_720,N_2210);
nand U8287 (N_8287,N_709,N_330);
or U8288 (N_8288,N_1737,N_1614);
xnor U8289 (N_8289,N_1134,N_2757);
or U8290 (N_8290,N_2167,N_222);
nor U8291 (N_8291,N_4251,N_423);
or U8292 (N_8292,N_633,N_726);
and U8293 (N_8293,N_1352,N_3451);
or U8294 (N_8294,N_4223,N_1478);
and U8295 (N_8295,N_3624,N_1639);
nand U8296 (N_8296,N_3494,N_4868);
nor U8297 (N_8297,N_2720,N_4574);
and U8298 (N_8298,N_1858,N_3892);
nand U8299 (N_8299,N_714,N_4747);
or U8300 (N_8300,N_2775,N_3905);
or U8301 (N_8301,N_4731,N_136);
or U8302 (N_8302,N_1256,N_222);
and U8303 (N_8303,N_1435,N_4082);
nor U8304 (N_8304,N_2307,N_3195);
nor U8305 (N_8305,N_1385,N_932);
and U8306 (N_8306,N_1391,N_3198);
nand U8307 (N_8307,N_1850,N_768);
and U8308 (N_8308,N_3593,N_1241);
nand U8309 (N_8309,N_2708,N_1415);
and U8310 (N_8310,N_557,N_1656);
xor U8311 (N_8311,N_3877,N_2270);
nand U8312 (N_8312,N_2971,N_284);
or U8313 (N_8313,N_526,N_1296);
or U8314 (N_8314,N_473,N_3526);
nor U8315 (N_8315,N_2707,N_4257);
nor U8316 (N_8316,N_3009,N_4867);
or U8317 (N_8317,N_453,N_2167);
or U8318 (N_8318,N_2798,N_1353);
and U8319 (N_8319,N_3275,N_1206);
or U8320 (N_8320,N_3499,N_1587);
and U8321 (N_8321,N_1774,N_1108);
nand U8322 (N_8322,N_3541,N_39);
xor U8323 (N_8323,N_1956,N_139);
xnor U8324 (N_8324,N_731,N_3533);
nand U8325 (N_8325,N_806,N_422);
and U8326 (N_8326,N_4667,N_1901);
nor U8327 (N_8327,N_4321,N_4944);
or U8328 (N_8328,N_2396,N_1235);
nand U8329 (N_8329,N_166,N_2279);
and U8330 (N_8330,N_502,N_2561);
and U8331 (N_8331,N_1160,N_2537);
nand U8332 (N_8332,N_2456,N_3152);
or U8333 (N_8333,N_3021,N_1130);
and U8334 (N_8334,N_1229,N_829);
nor U8335 (N_8335,N_4762,N_2840);
or U8336 (N_8336,N_1709,N_4859);
xor U8337 (N_8337,N_1794,N_174);
xor U8338 (N_8338,N_4646,N_1456);
xor U8339 (N_8339,N_2748,N_2872);
xor U8340 (N_8340,N_4096,N_1593);
nor U8341 (N_8341,N_2399,N_3815);
and U8342 (N_8342,N_3938,N_1956);
and U8343 (N_8343,N_2486,N_2901);
nor U8344 (N_8344,N_3244,N_4904);
nor U8345 (N_8345,N_3867,N_1569);
and U8346 (N_8346,N_2769,N_4120);
nor U8347 (N_8347,N_1683,N_3371);
nand U8348 (N_8348,N_1868,N_747);
xnor U8349 (N_8349,N_624,N_3730);
xor U8350 (N_8350,N_4257,N_4898);
and U8351 (N_8351,N_1998,N_2);
xnor U8352 (N_8352,N_1249,N_3481);
and U8353 (N_8353,N_3824,N_2943);
or U8354 (N_8354,N_4404,N_687);
or U8355 (N_8355,N_3686,N_4342);
xnor U8356 (N_8356,N_3914,N_4641);
nor U8357 (N_8357,N_2869,N_1489);
nand U8358 (N_8358,N_566,N_4805);
or U8359 (N_8359,N_3063,N_2761);
and U8360 (N_8360,N_1727,N_103);
and U8361 (N_8361,N_3350,N_1216);
and U8362 (N_8362,N_3997,N_4294);
xnor U8363 (N_8363,N_826,N_807);
and U8364 (N_8364,N_1972,N_3085);
xnor U8365 (N_8365,N_1513,N_993);
and U8366 (N_8366,N_3640,N_4412);
nand U8367 (N_8367,N_376,N_3772);
xnor U8368 (N_8368,N_680,N_1961);
and U8369 (N_8369,N_1171,N_4320);
nor U8370 (N_8370,N_378,N_879);
nor U8371 (N_8371,N_2871,N_1930);
or U8372 (N_8372,N_1498,N_3132);
nand U8373 (N_8373,N_3647,N_3738);
xor U8374 (N_8374,N_4962,N_1681);
nand U8375 (N_8375,N_91,N_4772);
xor U8376 (N_8376,N_4279,N_2971);
or U8377 (N_8377,N_3436,N_1287);
or U8378 (N_8378,N_3696,N_1476);
nor U8379 (N_8379,N_2568,N_3420);
nand U8380 (N_8380,N_334,N_10);
xnor U8381 (N_8381,N_2070,N_2287);
nor U8382 (N_8382,N_2472,N_3081);
or U8383 (N_8383,N_312,N_1168);
or U8384 (N_8384,N_2666,N_4944);
xor U8385 (N_8385,N_17,N_1401);
nand U8386 (N_8386,N_2743,N_4076);
and U8387 (N_8387,N_1922,N_2970);
xor U8388 (N_8388,N_577,N_330);
xnor U8389 (N_8389,N_4678,N_143);
and U8390 (N_8390,N_4819,N_217);
nor U8391 (N_8391,N_3761,N_2530);
and U8392 (N_8392,N_1749,N_4851);
or U8393 (N_8393,N_3017,N_4523);
nand U8394 (N_8394,N_397,N_1203);
and U8395 (N_8395,N_4656,N_4716);
nand U8396 (N_8396,N_266,N_2729);
nand U8397 (N_8397,N_2317,N_467);
nor U8398 (N_8398,N_4286,N_2772);
or U8399 (N_8399,N_862,N_4394);
nor U8400 (N_8400,N_3204,N_918);
or U8401 (N_8401,N_3609,N_786);
and U8402 (N_8402,N_164,N_764);
nor U8403 (N_8403,N_1535,N_4101);
and U8404 (N_8404,N_683,N_4905);
nor U8405 (N_8405,N_1776,N_4892);
or U8406 (N_8406,N_548,N_2053);
xor U8407 (N_8407,N_1582,N_3810);
xor U8408 (N_8408,N_1508,N_1325);
and U8409 (N_8409,N_1510,N_1289);
xor U8410 (N_8410,N_3723,N_4905);
nor U8411 (N_8411,N_3209,N_4149);
nor U8412 (N_8412,N_1905,N_2732);
or U8413 (N_8413,N_3147,N_551);
nor U8414 (N_8414,N_4235,N_4335);
nor U8415 (N_8415,N_330,N_1948);
nand U8416 (N_8416,N_984,N_1764);
nor U8417 (N_8417,N_1886,N_2373);
and U8418 (N_8418,N_2608,N_4864);
nand U8419 (N_8419,N_3516,N_4842);
and U8420 (N_8420,N_819,N_1479);
and U8421 (N_8421,N_1125,N_1680);
and U8422 (N_8422,N_1239,N_1089);
xnor U8423 (N_8423,N_3858,N_727);
nand U8424 (N_8424,N_2773,N_610);
and U8425 (N_8425,N_3893,N_4836);
xnor U8426 (N_8426,N_3226,N_249);
nor U8427 (N_8427,N_1985,N_2540);
and U8428 (N_8428,N_2134,N_796);
nor U8429 (N_8429,N_2807,N_805);
or U8430 (N_8430,N_4558,N_1129);
nor U8431 (N_8431,N_196,N_409);
or U8432 (N_8432,N_704,N_382);
nor U8433 (N_8433,N_4323,N_925);
nor U8434 (N_8434,N_3602,N_2831);
and U8435 (N_8435,N_4893,N_1963);
xor U8436 (N_8436,N_2723,N_2089);
and U8437 (N_8437,N_4180,N_1142);
and U8438 (N_8438,N_4693,N_2705);
nor U8439 (N_8439,N_4885,N_668);
nand U8440 (N_8440,N_1693,N_4786);
nor U8441 (N_8441,N_4012,N_450);
nand U8442 (N_8442,N_1941,N_3282);
and U8443 (N_8443,N_3036,N_777);
xor U8444 (N_8444,N_4705,N_4526);
and U8445 (N_8445,N_788,N_4940);
or U8446 (N_8446,N_4030,N_1988);
nand U8447 (N_8447,N_2092,N_3052);
nor U8448 (N_8448,N_3591,N_538);
and U8449 (N_8449,N_3273,N_3373);
xor U8450 (N_8450,N_346,N_2555);
and U8451 (N_8451,N_330,N_2771);
nor U8452 (N_8452,N_1213,N_1652);
xor U8453 (N_8453,N_4003,N_3888);
and U8454 (N_8454,N_1404,N_1220);
and U8455 (N_8455,N_878,N_1512);
xnor U8456 (N_8456,N_3523,N_508);
xor U8457 (N_8457,N_55,N_963);
nor U8458 (N_8458,N_517,N_2491);
and U8459 (N_8459,N_3639,N_2179);
and U8460 (N_8460,N_107,N_1682);
nor U8461 (N_8461,N_2749,N_3943);
nand U8462 (N_8462,N_1864,N_4209);
and U8463 (N_8463,N_1326,N_3787);
nor U8464 (N_8464,N_4697,N_2582);
xor U8465 (N_8465,N_397,N_231);
or U8466 (N_8466,N_555,N_1444);
and U8467 (N_8467,N_2611,N_3847);
xnor U8468 (N_8468,N_4643,N_928);
nor U8469 (N_8469,N_3338,N_1899);
nor U8470 (N_8470,N_3094,N_2343);
or U8471 (N_8471,N_3093,N_302);
xnor U8472 (N_8472,N_677,N_3836);
nand U8473 (N_8473,N_4952,N_3447);
nor U8474 (N_8474,N_1211,N_407);
nor U8475 (N_8475,N_4462,N_4935);
and U8476 (N_8476,N_3369,N_1071);
nand U8477 (N_8477,N_4009,N_4264);
or U8478 (N_8478,N_184,N_744);
nor U8479 (N_8479,N_3261,N_4930);
and U8480 (N_8480,N_3649,N_4263);
nor U8481 (N_8481,N_673,N_1199);
or U8482 (N_8482,N_1218,N_3602);
or U8483 (N_8483,N_4727,N_4587);
or U8484 (N_8484,N_3881,N_1696);
or U8485 (N_8485,N_3267,N_4474);
xor U8486 (N_8486,N_3574,N_1732);
nor U8487 (N_8487,N_2451,N_1705);
or U8488 (N_8488,N_308,N_2836);
and U8489 (N_8489,N_697,N_1070);
nand U8490 (N_8490,N_1897,N_2061);
xor U8491 (N_8491,N_3305,N_637);
xnor U8492 (N_8492,N_2611,N_1699);
or U8493 (N_8493,N_3870,N_2328);
or U8494 (N_8494,N_2063,N_101);
xor U8495 (N_8495,N_699,N_1041);
or U8496 (N_8496,N_3451,N_3798);
nand U8497 (N_8497,N_921,N_1692);
nor U8498 (N_8498,N_3171,N_1573);
xnor U8499 (N_8499,N_4211,N_4476);
and U8500 (N_8500,N_2228,N_2112);
xor U8501 (N_8501,N_258,N_2035);
and U8502 (N_8502,N_2933,N_2579);
nand U8503 (N_8503,N_2269,N_2313);
and U8504 (N_8504,N_4534,N_2957);
or U8505 (N_8505,N_4712,N_1249);
or U8506 (N_8506,N_1114,N_3803);
nand U8507 (N_8507,N_4841,N_974);
and U8508 (N_8508,N_505,N_1151);
xnor U8509 (N_8509,N_2457,N_476);
xor U8510 (N_8510,N_1143,N_4705);
nor U8511 (N_8511,N_767,N_4507);
xnor U8512 (N_8512,N_3266,N_1935);
xor U8513 (N_8513,N_649,N_335);
xor U8514 (N_8514,N_2515,N_1653);
and U8515 (N_8515,N_2968,N_1845);
nor U8516 (N_8516,N_797,N_4564);
and U8517 (N_8517,N_1468,N_280);
nor U8518 (N_8518,N_771,N_872);
and U8519 (N_8519,N_1059,N_3844);
xnor U8520 (N_8520,N_2580,N_1973);
nand U8521 (N_8521,N_589,N_3898);
and U8522 (N_8522,N_3260,N_3333);
nand U8523 (N_8523,N_1856,N_3588);
or U8524 (N_8524,N_3125,N_4770);
nor U8525 (N_8525,N_1811,N_1294);
nor U8526 (N_8526,N_4156,N_862);
nor U8527 (N_8527,N_2313,N_1862);
and U8528 (N_8528,N_1658,N_4233);
xnor U8529 (N_8529,N_4884,N_623);
or U8530 (N_8530,N_2411,N_398);
and U8531 (N_8531,N_4557,N_930);
and U8532 (N_8532,N_864,N_3469);
and U8533 (N_8533,N_3356,N_92);
or U8534 (N_8534,N_1153,N_3021);
nand U8535 (N_8535,N_4185,N_422);
nor U8536 (N_8536,N_3396,N_4003);
or U8537 (N_8537,N_3311,N_347);
nor U8538 (N_8538,N_4820,N_3967);
and U8539 (N_8539,N_3613,N_4054);
nor U8540 (N_8540,N_1805,N_3408);
nor U8541 (N_8541,N_222,N_1074);
and U8542 (N_8542,N_3149,N_52);
and U8543 (N_8543,N_2841,N_4014);
xnor U8544 (N_8544,N_3499,N_2754);
or U8545 (N_8545,N_4698,N_160);
nand U8546 (N_8546,N_3629,N_2023);
nand U8547 (N_8547,N_2243,N_3774);
xor U8548 (N_8548,N_4879,N_907);
nand U8549 (N_8549,N_4712,N_1143);
nand U8550 (N_8550,N_1633,N_3987);
and U8551 (N_8551,N_929,N_4155);
or U8552 (N_8552,N_3070,N_4187);
nor U8553 (N_8553,N_3390,N_3544);
and U8554 (N_8554,N_4298,N_3452);
or U8555 (N_8555,N_2244,N_812);
nor U8556 (N_8556,N_4455,N_4703);
nor U8557 (N_8557,N_1505,N_3005);
xnor U8558 (N_8558,N_169,N_898);
nor U8559 (N_8559,N_3023,N_3485);
xnor U8560 (N_8560,N_3791,N_4154);
and U8561 (N_8561,N_3105,N_3345);
xnor U8562 (N_8562,N_1478,N_779);
nand U8563 (N_8563,N_228,N_3474);
nor U8564 (N_8564,N_3416,N_4503);
or U8565 (N_8565,N_1743,N_4244);
nor U8566 (N_8566,N_2972,N_1577);
nor U8567 (N_8567,N_3883,N_4305);
nor U8568 (N_8568,N_2864,N_1056);
xnor U8569 (N_8569,N_4196,N_869);
xor U8570 (N_8570,N_1898,N_286);
nand U8571 (N_8571,N_3617,N_1058);
xor U8572 (N_8572,N_2467,N_207);
and U8573 (N_8573,N_4113,N_1544);
nand U8574 (N_8574,N_4612,N_4418);
nor U8575 (N_8575,N_164,N_3887);
xor U8576 (N_8576,N_455,N_4752);
nand U8577 (N_8577,N_3416,N_4999);
nor U8578 (N_8578,N_246,N_1607);
nor U8579 (N_8579,N_2421,N_4342);
xor U8580 (N_8580,N_4767,N_2487);
nor U8581 (N_8581,N_4261,N_3873);
or U8582 (N_8582,N_1418,N_3967);
or U8583 (N_8583,N_1622,N_2410);
or U8584 (N_8584,N_2436,N_2989);
and U8585 (N_8585,N_128,N_2953);
and U8586 (N_8586,N_494,N_4027);
xor U8587 (N_8587,N_406,N_3671);
xnor U8588 (N_8588,N_2135,N_4673);
xnor U8589 (N_8589,N_333,N_4809);
or U8590 (N_8590,N_918,N_3585);
and U8591 (N_8591,N_767,N_1884);
xor U8592 (N_8592,N_2972,N_4280);
nand U8593 (N_8593,N_1473,N_2989);
and U8594 (N_8594,N_2290,N_4599);
xnor U8595 (N_8595,N_513,N_1791);
or U8596 (N_8596,N_628,N_2442);
nor U8597 (N_8597,N_4611,N_3510);
nor U8598 (N_8598,N_3969,N_191);
or U8599 (N_8599,N_4184,N_2011);
xor U8600 (N_8600,N_516,N_1898);
nor U8601 (N_8601,N_4728,N_841);
nand U8602 (N_8602,N_2183,N_2936);
and U8603 (N_8603,N_1470,N_3079);
or U8604 (N_8604,N_4077,N_4133);
or U8605 (N_8605,N_4841,N_3571);
nand U8606 (N_8606,N_3506,N_23);
nand U8607 (N_8607,N_4217,N_2450);
nor U8608 (N_8608,N_914,N_4598);
nand U8609 (N_8609,N_4391,N_971);
nor U8610 (N_8610,N_777,N_2823);
xor U8611 (N_8611,N_2309,N_4483);
nand U8612 (N_8612,N_2477,N_4980);
and U8613 (N_8613,N_4864,N_768);
and U8614 (N_8614,N_2504,N_3619);
xor U8615 (N_8615,N_1995,N_4008);
and U8616 (N_8616,N_1801,N_3857);
or U8617 (N_8617,N_3021,N_2471);
and U8618 (N_8618,N_3684,N_1939);
and U8619 (N_8619,N_2909,N_397);
nor U8620 (N_8620,N_2969,N_1392);
or U8621 (N_8621,N_1604,N_1886);
nor U8622 (N_8622,N_3560,N_1430);
xor U8623 (N_8623,N_2472,N_3758);
and U8624 (N_8624,N_595,N_3438);
and U8625 (N_8625,N_2647,N_170);
nor U8626 (N_8626,N_2576,N_33);
and U8627 (N_8627,N_4538,N_3434);
nand U8628 (N_8628,N_92,N_2090);
or U8629 (N_8629,N_4237,N_2301);
nand U8630 (N_8630,N_2337,N_2576);
xor U8631 (N_8631,N_1925,N_451);
xor U8632 (N_8632,N_876,N_2251);
xor U8633 (N_8633,N_521,N_622);
nand U8634 (N_8634,N_2573,N_2235);
or U8635 (N_8635,N_901,N_2591);
nor U8636 (N_8636,N_4515,N_831);
and U8637 (N_8637,N_3882,N_3817);
xor U8638 (N_8638,N_808,N_4922);
and U8639 (N_8639,N_1681,N_3531);
nor U8640 (N_8640,N_1350,N_3687);
nor U8641 (N_8641,N_3113,N_2782);
nor U8642 (N_8642,N_4190,N_2941);
xnor U8643 (N_8643,N_3194,N_286);
or U8644 (N_8644,N_1723,N_1849);
or U8645 (N_8645,N_1392,N_4188);
or U8646 (N_8646,N_522,N_1691);
or U8647 (N_8647,N_3569,N_3382);
nand U8648 (N_8648,N_4487,N_3860);
or U8649 (N_8649,N_4943,N_2032);
xnor U8650 (N_8650,N_3750,N_3636);
or U8651 (N_8651,N_2043,N_3778);
nor U8652 (N_8652,N_3901,N_3931);
xnor U8653 (N_8653,N_3112,N_2907);
or U8654 (N_8654,N_3457,N_3685);
xnor U8655 (N_8655,N_3664,N_4639);
nand U8656 (N_8656,N_1260,N_4666);
nand U8657 (N_8657,N_3725,N_3598);
nand U8658 (N_8658,N_1986,N_2100);
and U8659 (N_8659,N_1395,N_4700);
nor U8660 (N_8660,N_1943,N_3478);
or U8661 (N_8661,N_1557,N_280);
or U8662 (N_8662,N_3093,N_860);
xor U8663 (N_8663,N_4909,N_3065);
nand U8664 (N_8664,N_2531,N_3974);
or U8665 (N_8665,N_3467,N_4372);
and U8666 (N_8666,N_4284,N_3015);
and U8667 (N_8667,N_1167,N_382);
xnor U8668 (N_8668,N_834,N_3828);
nor U8669 (N_8669,N_4915,N_4835);
nor U8670 (N_8670,N_1815,N_161);
or U8671 (N_8671,N_523,N_108);
nand U8672 (N_8672,N_2452,N_1722);
nand U8673 (N_8673,N_3283,N_807);
nor U8674 (N_8674,N_3777,N_2899);
or U8675 (N_8675,N_263,N_3711);
nor U8676 (N_8676,N_3639,N_4727);
nand U8677 (N_8677,N_269,N_4512);
and U8678 (N_8678,N_2204,N_3288);
and U8679 (N_8679,N_2915,N_1960);
and U8680 (N_8680,N_273,N_4265);
and U8681 (N_8681,N_4882,N_3083);
nand U8682 (N_8682,N_976,N_2065);
and U8683 (N_8683,N_3293,N_567);
xnor U8684 (N_8684,N_691,N_1837);
or U8685 (N_8685,N_1872,N_3321);
or U8686 (N_8686,N_572,N_455);
nor U8687 (N_8687,N_2628,N_1046);
nor U8688 (N_8688,N_3258,N_1365);
xnor U8689 (N_8689,N_24,N_442);
nand U8690 (N_8690,N_1274,N_1243);
and U8691 (N_8691,N_4028,N_511);
xor U8692 (N_8692,N_3037,N_4551);
nor U8693 (N_8693,N_1345,N_2758);
nor U8694 (N_8694,N_4185,N_3623);
nand U8695 (N_8695,N_2066,N_3947);
nor U8696 (N_8696,N_2271,N_1832);
xor U8697 (N_8697,N_2220,N_3257);
nor U8698 (N_8698,N_3311,N_299);
and U8699 (N_8699,N_1096,N_2935);
xnor U8700 (N_8700,N_645,N_4570);
or U8701 (N_8701,N_1482,N_431);
xnor U8702 (N_8702,N_4184,N_4194);
nand U8703 (N_8703,N_896,N_1955);
and U8704 (N_8704,N_3983,N_2406);
nand U8705 (N_8705,N_544,N_4009);
or U8706 (N_8706,N_103,N_4065);
nand U8707 (N_8707,N_4575,N_2452);
nor U8708 (N_8708,N_1574,N_2024);
nand U8709 (N_8709,N_4751,N_576);
or U8710 (N_8710,N_2800,N_4899);
nor U8711 (N_8711,N_3781,N_1934);
nor U8712 (N_8712,N_1248,N_4192);
and U8713 (N_8713,N_4840,N_4758);
nand U8714 (N_8714,N_1751,N_4144);
nand U8715 (N_8715,N_2423,N_4926);
nor U8716 (N_8716,N_696,N_4676);
or U8717 (N_8717,N_499,N_3216);
xnor U8718 (N_8718,N_4631,N_2924);
xor U8719 (N_8719,N_2757,N_4803);
and U8720 (N_8720,N_3822,N_3451);
or U8721 (N_8721,N_669,N_259);
xnor U8722 (N_8722,N_3276,N_934);
or U8723 (N_8723,N_4755,N_3175);
and U8724 (N_8724,N_3201,N_3371);
and U8725 (N_8725,N_2054,N_231);
nor U8726 (N_8726,N_2943,N_524);
or U8727 (N_8727,N_1082,N_1137);
nor U8728 (N_8728,N_1975,N_998);
and U8729 (N_8729,N_1172,N_1590);
nand U8730 (N_8730,N_2630,N_1047);
nand U8731 (N_8731,N_3387,N_1812);
nand U8732 (N_8732,N_2239,N_2999);
nor U8733 (N_8733,N_4221,N_2057);
and U8734 (N_8734,N_3046,N_2867);
and U8735 (N_8735,N_4119,N_1573);
nand U8736 (N_8736,N_3063,N_742);
and U8737 (N_8737,N_4917,N_3837);
nand U8738 (N_8738,N_4879,N_746);
nor U8739 (N_8739,N_2438,N_2248);
and U8740 (N_8740,N_539,N_1096);
or U8741 (N_8741,N_3192,N_4212);
nor U8742 (N_8742,N_3245,N_400);
nor U8743 (N_8743,N_1578,N_122);
xor U8744 (N_8744,N_3732,N_2165);
or U8745 (N_8745,N_2245,N_2447);
nand U8746 (N_8746,N_694,N_3830);
xnor U8747 (N_8747,N_961,N_3600);
xnor U8748 (N_8748,N_3867,N_1207);
nor U8749 (N_8749,N_3488,N_273);
and U8750 (N_8750,N_456,N_2638);
and U8751 (N_8751,N_1592,N_2708);
nand U8752 (N_8752,N_3135,N_2092);
or U8753 (N_8753,N_4425,N_4218);
or U8754 (N_8754,N_134,N_1514);
xor U8755 (N_8755,N_4770,N_1373);
nor U8756 (N_8756,N_3474,N_3883);
nor U8757 (N_8757,N_1857,N_537);
and U8758 (N_8758,N_384,N_4536);
and U8759 (N_8759,N_2756,N_1665);
and U8760 (N_8760,N_1234,N_211);
nand U8761 (N_8761,N_696,N_1829);
xnor U8762 (N_8762,N_4599,N_2706);
or U8763 (N_8763,N_2651,N_48);
nor U8764 (N_8764,N_751,N_2472);
xor U8765 (N_8765,N_345,N_1176);
or U8766 (N_8766,N_3516,N_3514);
xnor U8767 (N_8767,N_1982,N_1098);
and U8768 (N_8768,N_1720,N_3882);
xor U8769 (N_8769,N_4752,N_1370);
and U8770 (N_8770,N_8,N_732);
xnor U8771 (N_8771,N_662,N_1932);
xnor U8772 (N_8772,N_1696,N_225);
nor U8773 (N_8773,N_3179,N_566);
or U8774 (N_8774,N_399,N_3141);
or U8775 (N_8775,N_3666,N_3885);
xnor U8776 (N_8776,N_324,N_4944);
and U8777 (N_8777,N_3799,N_1064);
and U8778 (N_8778,N_2868,N_4049);
nor U8779 (N_8779,N_4198,N_2106);
nor U8780 (N_8780,N_4030,N_1876);
and U8781 (N_8781,N_1746,N_4005);
nor U8782 (N_8782,N_87,N_3918);
xor U8783 (N_8783,N_4100,N_4064);
and U8784 (N_8784,N_3193,N_3351);
nor U8785 (N_8785,N_3772,N_4768);
or U8786 (N_8786,N_2603,N_1866);
nor U8787 (N_8787,N_3831,N_918);
and U8788 (N_8788,N_2641,N_499);
nand U8789 (N_8789,N_2301,N_373);
nand U8790 (N_8790,N_4730,N_1811);
or U8791 (N_8791,N_1487,N_937);
and U8792 (N_8792,N_4878,N_3508);
or U8793 (N_8793,N_1200,N_421);
and U8794 (N_8794,N_1315,N_234);
nand U8795 (N_8795,N_3570,N_847);
and U8796 (N_8796,N_1124,N_1094);
or U8797 (N_8797,N_706,N_109);
or U8798 (N_8798,N_3699,N_3640);
nand U8799 (N_8799,N_4653,N_1510);
and U8800 (N_8800,N_2068,N_1562);
and U8801 (N_8801,N_659,N_1892);
xor U8802 (N_8802,N_2513,N_1976);
and U8803 (N_8803,N_859,N_886);
nand U8804 (N_8804,N_2991,N_3907);
and U8805 (N_8805,N_790,N_4372);
nor U8806 (N_8806,N_3701,N_2251);
nor U8807 (N_8807,N_215,N_3953);
and U8808 (N_8808,N_3723,N_3404);
xor U8809 (N_8809,N_4590,N_411);
xnor U8810 (N_8810,N_1794,N_4108);
xor U8811 (N_8811,N_882,N_4892);
nor U8812 (N_8812,N_1918,N_87);
and U8813 (N_8813,N_2454,N_897);
xor U8814 (N_8814,N_1934,N_1011);
nand U8815 (N_8815,N_2590,N_3452);
nor U8816 (N_8816,N_1370,N_1153);
nor U8817 (N_8817,N_459,N_2926);
or U8818 (N_8818,N_1619,N_1886);
or U8819 (N_8819,N_1333,N_405);
or U8820 (N_8820,N_2417,N_1277);
nand U8821 (N_8821,N_1389,N_2912);
and U8822 (N_8822,N_1212,N_4723);
nor U8823 (N_8823,N_2775,N_2458);
or U8824 (N_8824,N_4771,N_2844);
nor U8825 (N_8825,N_4404,N_929);
nor U8826 (N_8826,N_1540,N_3669);
nand U8827 (N_8827,N_1864,N_1439);
xnor U8828 (N_8828,N_2925,N_1418);
nor U8829 (N_8829,N_2334,N_2781);
and U8830 (N_8830,N_2084,N_1827);
and U8831 (N_8831,N_5,N_2196);
nor U8832 (N_8832,N_495,N_2193);
and U8833 (N_8833,N_790,N_2241);
xor U8834 (N_8834,N_1325,N_356);
nor U8835 (N_8835,N_2022,N_953);
nor U8836 (N_8836,N_4410,N_4130);
and U8837 (N_8837,N_271,N_204);
xnor U8838 (N_8838,N_743,N_4861);
or U8839 (N_8839,N_3632,N_2899);
xor U8840 (N_8840,N_3932,N_978);
nand U8841 (N_8841,N_3245,N_1128);
nand U8842 (N_8842,N_143,N_3377);
nand U8843 (N_8843,N_4055,N_557);
and U8844 (N_8844,N_714,N_1817);
or U8845 (N_8845,N_4724,N_707);
or U8846 (N_8846,N_4567,N_3950);
or U8847 (N_8847,N_3654,N_4774);
nand U8848 (N_8848,N_1862,N_4644);
xnor U8849 (N_8849,N_3346,N_4246);
nand U8850 (N_8850,N_1734,N_1828);
and U8851 (N_8851,N_1823,N_4680);
xor U8852 (N_8852,N_4787,N_221);
xor U8853 (N_8853,N_2881,N_4791);
xor U8854 (N_8854,N_1735,N_1406);
or U8855 (N_8855,N_432,N_973);
nand U8856 (N_8856,N_3641,N_1747);
and U8857 (N_8857,N_1917,N_148);
nor U8858 (N_8858,N_815,N_1535);
nand U8859 (N_8859,N_2295,N_2434);
or U8860 (N_8860,N_960,N_322);
or U8861 (N_8861,N_751,N_1249);
nand U8862 (N_8862,N_4632,N_1517);
and U8863 (N_8863,N_118,N_3250);
xnor U8864 (N_8864,N_3430,N_4787);
and U8865 (N_8865,N_2983,N_2345);
and U8866 (N_8866,N_224,N_1798);
xnor U8867 (N_8867,N_4535,N_295);
or U8868 (N_8868,N_2913,N_1981);
xor U8869 (N_8869,N_1665,N_3765);
or U8870 (N_8870,N_632,N_1723);
xnor U8871 (N_8871,N_137,N_544);
or U8872 (N_8872,N_4914,N_3301);
and U8873 (N_8873,N_4451,N_4304);
nor U8874 (N_8874,N_3657,N_420);
nor U8875 (N_8875,N_3193,N_2331);
xnor U8876 (N_8876,N_4520,N_66);
and U8877 (N_8877,N_123,N_4156);
and U8878 (N_8878,N_18,N_3941);
nand U8879 (N_8879,N_3760,N_4022);
and U8880 (N_8880,N_3935,N_3683);
nand U8881 (N_8881,N_1031,N_3731);
and U8882 (N_8882,N_3813,N_3260);
or U8883 (N_8883,N_4718,N_4039);
and U8884 (N_8884,N_3668,N_3724);
nand U8885 (N_8885,N_365,N_4247);
nand U8886 (N_8886,N_4278,N_3957);
nor U8887 (N_8887,N_2639,N_1828);
nand U8888 (N_8888,N_519,N_1478);
and U8889 (N_8889,N_1046,N_2279);
nor U8890 (N_8890,N_4905,N_591);
or U8891 (N_8891,N_1955,N_4956);
nor U8892 (N_8892,N_2720,N_2695);
nand U8893 (N_8893,N_3777,N_2830);
or U8894 (N_8894,N_4172,N_462);
nand U8895 (N_8895,N_116,N_4170);
nor U8896 (N_8896,N_1122,N_933);
and U8897 (N_8897,N_4858,N_3801);
and U8898 (N_8898,N_3579,N_2182);
and U8899 (N_8899,N_3905,N_3871);
nor U8900 (N_8900,N_3947,N_1867);
or U8901 (N_8901,N_4247,N_4210);
nor U8902 (N_8902,N_3224,N_2558);
xnor U8903 (N_8903,N_1152,N_1237);
xor U8904 (N_8904,N_1776,N_4816);
and U8905 (N_8905,N_4535,N_2680);
nand U8906 (N_8906,N_1301,N_1479);
and U8907 (N_8907,N_246,N_3809);
or U8908 (N_8908,N_4054,N_167);
xnor U8909 (N_8909,N_668,N_3173);
or U8910 (N_8910,N_532,N_2886);
and U8911 (N_8911,N_3431,N_996);
xnor U8912 (N_8912,N_2820,N_158);
or U8913 (N_8913,N_3365,N_4072);
or U8914 (N_8914,N_2694,N_329);
nand U8915 (N_8915,N_2758,N_3362);
or U8916 (N_8916,N_1758,N_3809);
nor U8917 (N_8917,N_4855,N_3092);
nand U8918 (N_8918,N_2454,N_1919);
nor U8919 (N_8919,N_4725,N_1595);
and U8920 (N_8920,N_2671,N_66);
nand U8921 (N_8921,N_849,N_4786);
xnor U8922 (N_8922,N_3847,N_4808);
or U8923 (N_8923,N_4753,N_3149);
and U8924 (N_8924,N_3295,N_4040);
xnor U8925 (N_8925,N_198,N_2166);
or U8926 (N_8926,N_3506,N_2627);
xnor U8927 (N_8927,N_3036,N_102);
nor U8928 (N_8928,N_1503,N_1592);
nand U8929 (N_8929,N_3706,N_576);
xor U8930 (N_8930,N_3659,N_633);
xor U8931 (N_8931,N_1573,N_2939);
or U8932 (N_8932,N_178,N_49);
and U8933 (N_8933,N_2800,N_3096);
xor U8934 (N_8934,N_2158,N_3101);
and U8935 (N_8935,N_246,N_4356);
and U8936 (N_8936,N_2035,N_1447);
or U8937 (N_8937,N_1050,N_3203);
and U8938 (N_8938,N_1217,N_1856);
nor U8939 (N_8939,N_2238,N_4109);
xnor U8940 (N_8940,N_4494,N_2480);
or U8941 (N_8941,N_2621,N_588);
or U8942 (N_8942,N_4096,N_2664);
and U8943 (N_8943,N_1738,N_3303);
nand U8944 (N_8944,N_964,N_1789);
and U8945 (N_8945,N_3478,N_2391);
and U8946 (N_8946,N_2065,N_3883);
nand U8947 (N_8947,N_2842,N_1560);
or U8948 (N_8948,N_2435,N_1692);
nand U8949 (N_8949,N_4025,N_4350);
or U8950 (N_8950,N_54,N_3037);
nor U8951 (N_8951,N_4804,N_2599);
and U8952 (N_8952,N_2244,N_4371);
xor U8953 (N_8953,N_4976,N_3363);
xnor U8954 (N_8954,N_3527,N_1802);
or U8955 (N_8955,N_2147,N_1947);
nand U8956 (N_8956,N_391,N_3957);
and U8957 (N_8957,N_1232,N_2226);
nor U8958 (N_8958,N_2129,N_4427);
nand U8959 (N_8959,N_2829,N_2287);
nand U8960 (N_8960,N_3389,N_1286);
or U8961 (N_8961,N_3879,N_529);
xnor U8962 (N_8962,N_4743,N_1431);
nor U8963 (N_8963,N_3911,N_561);
or U8964 (N_8964,N_3681,N_3420);
and U8965 (N_8965,N_4281,N_4908);
or U8966 (N_8966,N_4293,N_1354);
nand U8967 (N_8967,N_2736,N_3511);
nor U8968 (N_8968,N_2140,N_1453);
and U8969 (N_8969,N_4482,N_1898);
nor U8970 (N_8970,N_1632,N_3203);
nor U8971 (N_8971,N_1075,N_4178);
nand U8972 (N_8972,N_1736,N_1680);
nand U8973 (N_8973,N_751,N_2867);
nor U8974 (N_8974,N_3696,N_1154);
nand U8975 (N_8975,N_410,N_101);
or U8976 (N_8976,N_1840,N_4046);
xnor U8977 (N_8977,N_3514,N_4108);
or U8978 (N_8978,N_723,N_4034);
or U8979 (N_8979,N_1205,N_1578);
or U8980 (N_8980,N_435,N_4728);
or U8981 (N_8981,N_3260,N_1010);
and U8982 (N_8982,N_1258,N_1825);
xor U8983 (N_8983,N_3166,N_3650);
nand U8984 (N_8984,N_4434,N_4598);
or U8985 (N_8985,N_64,N_2809);
xnor U8986 (N_8986,N_3298,N_2300);
or U8987 (N_8987,N_4594,N_37);
nand U8988 (N_8988,N_2810,N_1549);
xnor U8989 (N_8989,N_2822,N_1362);
and U8990 (N_8990,N_632,N_3360);
nand U8991 (N_8991,N_4529,N_2128);
and U8992 (N_8992,N_4009,N_1376);
and U8993 (N_8993,N_2546,N_1540);
and U8994 (N_8994,N_4088,N_451);
nand U8995 (N_8995,N_925,N_4195);
or U8996 (N_8996,N_4309,N_1871);
nand U8997 (N_8997,N_2923,N_962);
nand U8998 (N_8998,N_3122,N_3451);
or U8999 (N_8999,N_2841,N_3426);
nand U9000 (N_9000,N_1864,N_1976);
or U9001 (N_9001,N_1555,N_1392);
nor U9002 (N_9002,N_2888,N_4137);
or U9003 (N_9003,N_4649,N_4195);
xnor U9004 (N_9004,N_2181,N_1522);
xor U9005 (N_9005,N_58,N_3854);
and U9006 (N_9006,N_4264,N_4883);
and U9007 (N_9007,N_675,N_1499);
nor U9008 (N_9008,N_1956,N_1217);
and U9009 (N_9009,N_3435,N_2783);
or U9010 (N_9010,N_781,N_35);
nand U9011 (N_9011,N_1985,N_1473);
nand U9012 (N_9012,N_4120,N_4302);
and U9013 (N_9013,N_1283,N_3809);
xnor U9014 (N_9014,N_2003,N_1041);
and U9015 (N_9015,N_1614,N_985);
xnor U9016 (N_9016,N_4777,N_4008);
nor U9017 (N_9017,N_1314,N_3077);
and U9018 (N_9018,N_4783,N_126);
nand U9019 (N_9019,N_699,N_3119);
xnor U9020 (N_9020,N_2814,N_4014);
or U9021 (N_9021,N_849,N_421);
or U9022 (N_9022,N_2601,N_4866);
xor U9023 (N_9023,N_1212,N_37);
and U9024 (N_9024,N_1157,N_3325);
or U9025 (N_9025,N_2335,N_3271);
nand U9026 (N_9026,N_1554,N_3302);
or U9027 (N_9027,N_4329,N_2616);
nand U9028 (N_9028,N_4440,N_1132);
or U9029 (N_9029,N_1394,N_1415);
nand U9030 (N_9030,N_1207,N_4306);
or U9031 (N_9031,N_2158,N_2740);
xor U9032 (N_9032,N_1814,N_721);
or U9033 (N_9033,N_1208,N_3830);
nor U9034 (N_9034,N_1369,N_3047);
or U9035 (N_9035,N_1882,N_2871);
nand U9036 (N_9036,N_3658,N_3720);
or U9037 (N_9037,N_1242,N_790);
nand U9038 (N_9038,N_2824,N_3259);
nor U9039 (N_9039,N_1942,N_2950);
or U9040 (N_9040,N_4218,N_4331);
or U9041 (N_9041,N_859,N_4232);
nor U9042 (N_9042,N_1853,N_3119);
nor U9043 (N_9043,N_3707,N_3535);
nor U9044 (N_9044,N_1963,N_4678);
and U9045 (N_9045,N_1576,N_4034);
and U9046 (N_9046,N_108,N_3393);
nor U9047 (N_9047,N_1904,N_2500);
nor U9048 (N_9048,N_1390,N_3736);
and U9049 (N_9049,N_2272,N_1303);
nor U9050 (N_9050,N_4634,N_3999);
nor U9051 (N_9051,N_3018,N_2260);
nor U9052 (N_9052,N_152,N_1427);
nor U9053 (N_9053,N_1402,N_4762);
and U9054 (N_9054,N_1599,N_1618);
or U9055 (N_9055,N_491,N_502);
nand U9056 (N_9056,N_4480,N_3248);
nor U9057 (N_9057,N_2167,N_158);
and U9058 (N_9058,N_3410,N_567);
nor U9059 (N_9059,N_910,N_1995);
nand U9060 (N_9060,N_2690,N_599);
or U9061 (N_9061,N_1526,N_2095);
xor U9062 (N_9062,N_2120,N_2647);
and U9063 (N_9063,N_1612,N_1172);
nor U9064 (N_9064,N_2271,N_2827);
and U9065 (N_9065,N_2796,N_2579);
nand U9066 (N_9066,N_22,N_1404);
or U9067 (N_9067,N_883,N_4853);
xor U9068 (N_9068,N_3588,N_3266);
or U9069 (N_9069,N_1123,N_262);
or U9070 (N_9070,N_4737,N_2364);
and U9071 (N_9071,N_4996,N_2033);
nor U9072 (N_9072,N_597,N_4575);
nand U9073 (N_9073,N_4510,N_4149);
and U9074 (N_9074,N_2562,N_3353);
and U9075 (N_9075,N_2317,N_3618);
nor U9076 (N_9076,N_2452,N_3459);
or U9077 (N_9077,N_2211,N_164);
nor U9078 (N_9078,N_2188,N_317);
or U9079 (N_9079,N_2076,N_3433);
xor U9080 (N_9080,N_402,N_3960);
xor U9081 (N_9081,N_4717,N_132);
or U9082 (N_9082,N_3312,N_4066);
nor U9083 (N_9083,N_4996,N_1211);
nand U9084 (N_9084,N_3228,N_1487);
nor U9085 (N_9085,N_731,N_2410);
or U9086 (N_9086,N_3820,N_3779);
or U9087 (N_9087,N_2330,N_3441);
nand U9088 (N_9088,N_3193,N_3604);
or U9089 (N_9089,N_151,N_4244);
and U9090 (N_9090,N_2201,N_1528);
xnor U9091 (N_9091,N_1447,N_4255);
nand U9092 (N_9092,N_2113,N_4416);
xor U9093 (N_9093,N_3446,N_2923);
and U9094 (N_9094,N_1683,N_3920);
and U9095 (N_9095,N_4906,N_4049);
and U9096 (N_9096,N_530,N_1457);
and U9097 (N_9097,N_430,N_1673);
and U9098 (N_9098,N_2968,N_2052);
or U9099 (N_9099,N_3330,N_2427);
nor U9100 (N_9100,N_3579,N_781);
and U9101 (N_9101,N_2789,N_34);
nor U9102 (N_9102,N_307,N_1469);
or U9103 (N_9103,N_1137,N_2239);
and U9104 (N_9104,N_2877,N_3608);
or U9105 (N_9105,N_1456,N_3413);
or U9106 (N_9106,N_1345,N_3311);
and U9107 (N_9107,N_2040,N_3702);
nor U9108 (N_9108,N_1789,N_2152);
xnor U9109 (N_9109,N_4079,N_1013);
xor U9110 (N_9110,N_3801,N_3886);
nor U9111 (N_9111,N_2789,N_3381);
nor U9112 (N_9112,N_4258,N_952);
xnor U9113 (N_9113,N_384,N_309);
and U9114 (N_9114,N_1806,N_4013);
or U9115 (N_9115,N_483,N_970);
nor U9116 (N_9116,N_4902,N_4510);
and U9117 (N_9117,N_793,N_1952);
nor U9118 (N_9118,N_4309,N_820);
nand U9119 (N_9119,N_2444,N_1633);
nand U9120 (N_9120,N_3231,N_2102);
nor U9121 (N_9121,N_1673,N_1460);
and U9122 (N_9122,N_1117,N_2081);
nor U9123 (N_9123,N_1159,N_4720);
or U9124 (N_9124,N_3713,N_2983);
or U9125 (N_9125,N_1575,N_3814);
and U9126 (N_9126,N_3877,N_4353);
xor U9127 (N_9127,N_1446,N_4198);
nor U9128 (N_9128,N_907,N_829);
or U9129 (N_9129,N_2543,N_4379);
nor U9130 (N_9130,N_3642,N_447);
nor U9131 (N_9131,N_4451,N_940);
xor U9132 (N_9132,N_4394,N_373);
and U9133 (N_9133,N_24,N_4574);
nand U9134 (N_9134,N_4082,N_4744);
nand U9135 (N_9135,N_3733,N_2100);
nand U9136 (N_9136,N_2338,N_2989);
or U9137 (N_9137,N_660,N_1784);
nand U9138 (N_9138,N_214,N_1050);
xnor U9139 (N_9139,N_807,N_1818);
nand U9140 (N_9140,N_4177,N_1333);
xor U9141 (N_9141,N_564,N_170);
nor U9142 (N_9142,N_3902,N_940);
nand U9143 (N_9143,N_4856,N_2809);
or U9144 (N_9144,N_1397,N_3488);
nor U9145 (N_9145,N_1257,N_2442);
or U9146 (N_9146,N_2019,N_2023);
xnor U9147 (N_9147,N_3948,N_4505);
or U9148 (N_9148,N_2663,N_1223);
xor U9149 (N_9149,N_3661,N_652);
nand U9150 (N_9150,N_500,N_1574);
nand U9151 (N_9151,N_2360,N_1178);
nor U9152 (N_9152,N_3420,N_2405);
nor U9153 (N_9153,N_4013,N_3714);
nor U9154 (N_9154,N_4247,N_2436);
xnor U9155 (N_9155,N_3100,N_3526);
or U9156 (N_9156,N_1967,N_4700);
xnor U9157 (N_9157,N_631,N_3798);
and U9158 (N_9158,N_944,N_4674);
and U9159 (N_9159,N_3683,N_4591);
xnor U9160 (N_9160,N_2927,N_48);
and U9161 (N_9161,N_4695,N_2784);
or U9162 (N_9162,N_716,N_4029);
nor U9163 (N_9163,N_4267,N_4011);
nand U9164 (N_9164,N_251,N_4861);
or U9165 (N_9165,N_3383,N_3821);
xnor U9166 (N_9166,N_4640,N_1176);
xnor U9167 (N_9167,N_4237,N_264);
xor U9168 (N_9168,N_2957,N_1951);
and U9169 (N_9169,N_2368,N_1140);
xor U9170 (N_9170,N_4601,N_438);
or U9171 (N_9171,N_2457,N_4373);
nand U9172 (N_9172,N_3179,N_2205);
nor U9173 (N_9173,N_1059,N_1610);
nand U9174 (N_9174,N_4481,N_1593);
and U9175 (N_9175,N_3470,N_355);
nor U9176 (N_9176,N_188,N_238);
xor U9177 (N_9177,N_49,N_1894);
or U9178 (N_9178,N_4623,N_2482);
and U9179 (N_9179,N_2278,N_1539);
nand U9180 (N_9180,N_533,N_3188);
or U9181 (N_9181,N_4005,N_3550);
nor U9182 (N_9182,N_2865,N_4012);
nor U9183 (N_9183,N_1018,N_3906);
nand U9184 (N_9184,N_1534,N_2643);
nand U9185 (N_9185,N_516,N_2880);
nand U9186 (N_9186,N_3025,N_1673);
nor U9187 (N_9187,N_2304,N_51);
and U9188 (N_9188,N_3387,N_3021);
or U9189 (N_9189,N_2851,N_4919);
and U9190 (N_9190,N_3207,N_4481);
nand U9191 (N_9191,N_4648,N_2970);
or U9192 (N_9192,N_1127,N_4939);
nand U9193 (N_9193,N_1518,N_3345);
or U9194 (N_9194,N_3437,N_1674);
nor U9195 (N_9195,N_3365,N_2934);
nor U9196 (N_9196,N_3259,N_725);
or U9197 (N_9197,N_4292,N_2243);
or U9198 (N_9198,N_2511,N_176);
nand U9199 (N_9199,N_4537,N_4915);
and U9200 (N_9200,N_512,N_528);
nand U9201 (N_9201,N_4732,N_4890);
nor U9202 (N_9202,N_2891,N_3529);
xor U9203 (N_9203,N_1010,N_1906);
nand U9204 (N_9204,N_3767,N_2475);
nand U9205 (N_9205,N_673,N_3397);
and U9206 (N_9206,N_2278,N_670);
nor U9207 (N_9207,N_1985,N_3124);
nor U9208 (N_9208,N_2892,N_410);
nor U9209 (N_9209,N_2159,N_2807);
nand U9210 (N_9210,N_4609,N_4436);
or U9211 (N_9211,N_2630,N_2048);
xor U9212 (N_9212,N_4385,N_3532);
nand U9213 (N_9213,N_2843,N_255);
and U9214 (N_9214,N_3008,N_3987);
and U9215 (N_9215,N_1445,N_2935);
nor U9216 (N_9216,N_2124,N_4397);
and U9217 (N_9217,N_1474,N_3276);
or U9218 (N_9218,N_2306,N_110);
xnor U9219 (N_9219,N_2560,N_1891);
and U9220 (N_9220,N_4201,N_2100);
or U9221 (N_9221,N_4838,N_3560);
nand U9222 (N_9222,N_2779,N_1988);
nor U9223 (N_9223,N_3945,N_2123);
nor U9224 (N_9224,N_4709,N_2260);
xor U9225 (N_9225,N_777,N_220);
nor U9226 (N_9226,N_356,N_731);
xor U9227 (N_9227,N_4875,N_3758);
nand U9228 (N_9228,N_654,N_4166);
and U9229 (N_9229,N_4638,N_1867);
nor U9230 (N_9230,N_3866,N_1415);
nor U9231 (N_9231,N_3836,N_377);
or U9232 (N_9232,N_1797,N_782);
and U9233 (N_9233,N_3705,N_876);
nor U9234 (N_9234,N_4567,N_2040);
nor U9235 (N_9235,N_2421,N_3532);
xor U9236 (N_9236,N_2596,N_1159);
nand U9237 (N_9237,N_3284,N_2773);
and U9238 (N_9238,N_1458,N_3750);
and U9239 (N_9239,N_2492,N_1038);
nor U9240 (N_9240,N_3955,N_2347);
nor U9241 (N_9241,N_2899,N_3217);
and U9242 (N_9242,N_1020,N_456);
nand U9243 (N_9243,N_3731,N_747);
nor U9244 (N_9244,N_4269,N_2017);
and U9245 (N_9245,N_4046,N_4892);
and U9246 (N_9246,N_343,N_1557);
and U9247 (N_9247,N_3807,N_3975);
or U9248 (N_9248,N_1748,N_1449);
xnor U9249 (N_9249,N_683,N_3398);
nand U9250 (N_9250,N_3527,N_713);
and U9251 (N_9251,N_988,N_2909);
xor U9252 (N_9252,N_791,N_1122);
or U9253 (N_9253,N_3067,N_1252);
xnor U9254 (N_9254,N_1163,N_4809);
or U9255 (N_9255,N_1363,N_89);
or U9256 (N_9256,N_2960,N_4138);
xnor U9257 (N_9257,N_1116,N_883);
or U9258 (N_9258,N_2273,N_2219);
xor U9259 (N_9259,N_1519,N_4588);
xnor U9260 (N_9260,N_4326,N_3430);
nor U9261 (N_9261,N_4758,N_3433);
nor U9262 (N_9262,N_1155,N_4494);
xor U9263 (N_9263,N_4591,N_1780);
xnor U9264 (N_9264,N_3389,N_4926);
or U9265 (N_9265,N_2516,N_1994);
nand U9266 (N_9266,N_2865,N_2331);
nand U9267 (N_9267,N_3317,N_4286);
nand U9268 (N_9268,N_3416,N_1891);
nor U9269 (N_9269,N_3382,N_1310);
nor U9270 (N_9270,N_3537,N_1511);
nor U9271 (N_9271,N_2978,N_1353);
or U9272 (N_9272,N_4054,N_2849);
xor U9273 (N_9273,N_1716,N_16);
and U9274 (N_9274,N_19,N_4724);
nand U9275 (N_9275,N_1475,N_3225);
xor U9276 (N_9276,N_3044,N_4036);
and U9277 (N_9277,N_3996,N_751);
nor U9278 (N_9278,N_1628,N_1372);
nand U9279 (N_9279,N_1022,N_4096);
or U9280 (N_9280,N_942,N_3134);
xor U9281 (N_9281,N_1980,N_1266);
and U9282 (N_9282,N_4736,N_4359);
nand U9283 (N_9283,N_1814,N_1134);
or U9284 (N_9284,N_1622,N_2681);
nand U9285 (N_9285,N_2105,N_421);
nand U9286 (N_9286,N_4866,N_3791);
and U9287 (N_9287,N_4368,N_4883);
xnor U9288 (N_9288,N_3987,N_4685);
xor U9289 (N_9289,N_2378,N_1314);
xnor U9290 (N_9290,N_2608,N_2798);
and U9291 (N_9291,N_163,N_839);
nand U9292 (N_9292,N_345,N_1782);
nand U9293 (N_9293,N_632,N_1381);
nand U9294 (N_9294,N_4834,N_4145);
nand U9295 (N_9295,N_4997,N_2637);
or U9296 (N_9296,N_3700,N_2425);
nor U9297 (N_9297,N_4974,N_3582);
and U9298 (N_9298,N_3523,N_196);
xnor U9299 (N_9299,N_1211,N_1713);
nor U9300 (N_9300,N_2595,N_4708);
or U9301 (N_9301,N_976,N_4901);
nand U9302 (N_9302,N_3917,N_3940);
xor U9303 (N_9303,N_1538,N_1118);
nor U9304 (N_9304,N_331,N_2692);
nor U9305 (N_9305,N_3029,N_2652);
or U9306 (N_9306,N_3740,N_4661);
nor U9307 (N_9307,N_3418,N_3181);
and U9308 (N_9308,N_1706,N_1530);
nor U9309 (N_9309,N_3383,N_4684);
nand U9310 (N_9310,N_3692,N_2741);
or U9311 (N_9311,N_1676,N_2022);
nand U9312 (N_9312,N_750,N_2277);
xnor U9313 (N_9313,N_1949,N_3014);
and U9314 (N_9314,N_4588,N_352);
nor U9315 (N_9315,N_2458,N_1799);
and U9316 (N_9316,N_1744,N_3428);
and U9317 (N_9317,N_821,N_1389);
nor U9318 (N_9318,N_3703,N_727);
or U9319 (N_9319,N_766,N_1657);
xor U9320 (N_9320,N_4832,N_1639);
xnor U9321 (N_9321,N_3218,N_1869);
nand U9322 (N_9322,N_358,N_1261);
or U9323 (N_9323,N_2765,N_1603);
nand U9324 (N_9324,N_3445,N_4344);
or U9325 (N_9325,N_1536,N_4227);
xor U9326 (N_9326,N_4713,N_2127);
or U9327 (N_9327,N_1479,N_4065);
and U9328 (N_9328,N_2018,N_3139);
and U9329 (N_9329,N_53,N_3041);
and U9330 (N_9330,N_2174,N_4080);
xnor U9331 (N_9331,N_529,N_4765);
nor U9332 (N_9332,N_3140,N_4836);
nand U9333 (N_9333,N_1715,N_4981);
xnor U9334 (N_9334,N_1030,N_3750);
nor U9335 (N_9335,N_4371,N_2444);
xnor U9336 (N_9336,N_2784,N_1030);
nand U9337 (N_9337,N_4525,N_2976);
and U9338 (N_9338,N_1936,N_3088);
nand U9339 (N_9339,N_1336,N_2117);
nor U9340 (N_9340,N_1066,N_4411);
nor U9341 (N_9341,N_4868,N_4055);
nand U9342 (N_9342,N_320,N_4396);
and U9343 (N_9343,N_1382,N_3653);
and U9344 (N_9344,N_2686,N_56);
nor U9345 (N_9345,N_1049,N_2875);
nor U9346 (N_9346,N_79,N_3487);
and U9347 (N_9347,N_3574,N_3342);
or U9348 (N_9348,N_688,N_1308);
xnor U9349 (N_9349,N_4390,N_1105);
nand U9350 (N_9350,N_3022,N_4478);
or U9351 (N_9351,N_4346,N_3217);
nand U9352 (N_9352,N_3976,N_4809);
or U9353 (N_9353,N_4671,N_2951);
xor U9354 (N_9354,N_3297,N_1491);
nor U9355 (N_9355,N_3032,N_214);
and U9356 (N_9356,N_1864,N_3787);
or U9357 (N_9357,N_4333,N_472);
nor U9358 (N_9358,N_3315,N_1575);
and U9359 (N_9359,N_4167,N_3153);
or U9360 (N_9360,N_1007,N_1719);
and U9361 (N_9361,N_4036,N_190);
or U9362 (N_9362,N_422,N_2827);
xor U9363 (N_9363,N_892,N_2676);
nor U9364 (N_9364,N_3417,N_4704);
xor U9365 (N_9365,N_3526,N_758);
nor U9366 (N_9366,N_2946,N_2809);
nor U9367 (N_9367,N_4928,N_2252);
nand U9368 (N_9368,N_475,N_327);
or U9369 (N_9369,N_3199,N_3038);
nand U9370 (N_9370,N_1201,N_1134);
nor U9371 (N_9371,N_3271,N_3757);
nand U9372 (N_9372,N_3734,N_2383);
nor U9373 (N_9373,N_4535,N_4211);
nand U9374 (N_9374,N_3909,N_3831);
xnor U9375 (N_9375,N_550,N_1351);
nand U9376 (N_9376,N_3190,N_1999);
or U9377 (N_9377,N_3805,N_1271);
xnor U9378 (N_9378,N_4215,N_3725);
and U9379 (N_9379,N_1405,N_2937);
and U9380 (N_9380,N_3925,N_3101);
and U9381 (N_9381,N_1789,N_319);
xnor U9382 (N_9382,N_3887,N_3946);
and U9383 (N_9383,N_592,N_4483);
and U9384 (N_9384,N_3530,N_4848);
nor U9385 (N_9385,N_1850,N_1481);
nand U9386 (N_9386,N_2658,N_232);
xor U9387 (N_9387,N_2109,N_2724);
xor U9388 (N_9388,N_816,N_1939);
and U9389 (N_9389,N_1125,N_520);
xnor U9390 (N_9390,N_2320,N_3393);
and U9391 (N_9391,N_4482,N_3047);
nand U9392 (N_9392,N_1342,N_4407);
and U9393 (N_9393,N_2163,N_3790);
or U9394 (N_9394,N_2582,N_4395);
xnor U9395 (N_9395,N_2287,N_4005);
nor U9396 (N_9396,N_244,N_3154);
or U9397 (N_9397,N_3933,N_3527);
and U9398 (N_9398,N_4275,N_3949);
nand U9399 (N_9399,N_1682,N_4438);
or U9400 (N_9400,N_4911,N_3586);
and U9401 (N_9401,N_1184,N_1390);
nand U9402 (N_9402,N_2203,N_4422);
nand U9403 (N_9403,N_1541,N_4452);
nand U9404 (N_9404,N_2830,N_3741);
xnor U9405 (N_9405,N_1091,N_3299);
and U9406 (N_9406,N_586,N_2017);
or U9407 (N_9407,N_60,N_4626);
nor U9408 (N_9408,N_1984,N_1503);
or U9409 (N_9409,N_4616,N_2777);
nand U9410 (N_9410,N_3856,N_236);
or U9411 (N_9411,N_3837,N_4853);
or U9412 (N_9412,N_2734,N_3304);
or U9413 (N_9413,N_1243,N_4291);
nor U9414 (N_9414,N_3916,N_4626);
xor U9415 (N_9415,N_3132,N_4403);
or U9416 (N_9416,N_89,N_4760);
nor U9417 (N_9417,N_1875,N_4439);
or U9418 (N_9418,N_1706,N_3471);
and U9419 (N_9419,N_2929,N_4954);
xnor U9420 (N_9420,N_1124,N_126);
nand U9421 (N_9421,N_3456,N_3590);
and U9422 (N_9422,N_803,N_3427);
nand U9423 (N_9423,N_1863,N_73);
nand U9424 (N_9424,N_519,N_256);
and U9425 (N_9425,N_4457,N_444);
and U9426 (N_9426,N_555,N_2291);
nor U9427 (N_9427,N_3444,N_2403);
xor U9428 (N_9428,N_3811,N_2373);
nor U9429 (N_9429,N_238,N_741);
nor U9430 (N_9430,N_1668,N_2140);
xor U9431 (N_9431,N_3937,N_743);
nor U9432 (N_9432,N_4946,N_2230);
nand U9433 (N_9433,N_1658,N_331);
nor U9434 (N_9434,N_970,N_4096);
and U9435 (N_9435,N_4133,N_102);
nor U9436 (N_9436,N_2558,N_4627);
xor U9437 (N_9437,N_57,N_4301);
nor U9438 (N_9438,N_1539,N_4914);
nand U9439 (N_9439,N_3583,N_2577);
and U9440 (N_9440,N_3666,N_4931);
nand U9441 (N_9441,N_3288,N_587);
nand U9442 (N_9442,N_923,N_4477);
nor U9443 (N_9443,N_2789,N_3173);
and U9444 (N_9444,N_2470,N_1357);
and U9445 (N_9445,N_3312,N_1309);
xor U9446 (N_9446,N_1426,N_185);
nor U9447 (N_9447,N_123,N_2662);
nand U9448 (N_9448,N_852,N_1617);
or U9449 (N_9449,N_4842,N_463);
xor U9450 (N_9450,N_47,N_2955);
xnor U9451 (N_9451,N_2875,N_728);
or U9452 (N_9452,N_2286,N_1096);
nor U9453 (N_9453,N_2542,N_4873);
and U9454 (N_9454,N_1441,N_4448);
or U9455 (N_9455,N_2061,N_3123);
nand U9456 (N_9456,N_2195,N_3460);
xor U9457 (N_9457,N_3311,N_3930);
or U9458 (N_9458,N_3303,N_2998);
and U9459 (N_9459,N_4128,N_3686);
and U9460 (N_9460,N_2627,N_1650);
nand U9461 (N_9461,N_2827,N_4621);
nand U9462 (N_9462,N_2761,N_4533);
nand U9463 (N_9463,N_1186,N_3676);
or U9464 (N_9464,N_3835,N_1393);
and U9465 (N_9465,N_3320,N_3370);
nand U9466 (N_9466,N_1273,N_1565);
and U9467 (N_9467,N_4514,N_3667);
and U9468 (N_9468,N_1950,N_508);
and U9469 (N_9469,N_748,N_837);
and U9470 (N_9470,N_1493,N_4481);
or U9471 (N_9471,N_1891,N_291);
nor U9472 (N_9472,N_1623,N_1172);
or U9473 (N_9473,N_3183,N_3978);
xor U9474 (N_9474,N_2219,N_3703);
nand U9475 (N_9475,N_1370,N_199);
xor U9476 (N_9476,N_1497,N_4078);
and U9477 (N_9477,N_1317,N_4890);
or U9478 (N_9478,N_2262,N_3432);
nand U9479 (N_9479,N_3081,N_327);
nor U9480 (N_9480,N_1342,N_2026);
and U9481 (N_9481,N_1217,N_239);
nor U9482 (N_9482,N_1023,N_4374);
or U9483 (N_9483,N_1395,N_2478);
and U9484 (N_9484,N_3818,N_4653);
xnor U9485 (N_9485,N_3826,N_3233);
nand U9486 (N_9486,N_3837,N_307);
xor U9487 (N_9487,N_1135,N_2301);
nor U9488 (N_9488,N_3409,N_3550);
nor U9489 (N_9489,N_1307,N_4555);
nor U9490 (N_9490,N_1099,N_1602);
xnor U9491 (N_9491,N_2946,N_431);
nand U9492 (N_9492,N_933,N_1489);
nand U9493 (N_9493,N_3128,N_2642);
or U9494 (N_9494,N_1879,N_3500);
and U9495 (N_9495,N_3618,N_2949);
and U9496 (N_9496,N_2775,N_1871);
xor U9497 (N_9497,N_4626,N_2784);
nand U9498 (N_9498,N_1824,N_4934);
xor U9499 (N_9499,N_3782,N_590);
or U9500 (N_9500,N_56,N_26);
xnor U9501 (N_9501,N_3248,N_3908);
xor U9502 (N_9502,N_2512,N_2156);
and U9503 (N_9503,N_1514,N_2243);
xor U9504 (N_9504,N_4476,N_998);
and U9505 (N_9505,N_1728,N_2624);
nand U9506 (N_9506,N_3559,N_4872);
nor U9507 (N_9507,N_2740,N_1993);
and U9508 (N_9508,N_2949,N_2983);
xor U9509 (N_9509,N_455,N_3341);
nand U9510 (N_9510,N_3996,N_919);
nor U9511 (N_9511,N_1232,N_2616);
and U9512 (N_9512,N_4935,N_1325);
or U9513 (N_9513,N_3848,N_2374);
or U9514 (N_9514,N_2928,N_4429);
and U9515 (N_9515,N_1920,N_2248);
or U9516 (N_9516,N_2741,N_186);
and U9517 (N_9517,N_3132,N_3798);
or U9518 (N_9518,N_2227,N_4513);
xnor U9519 (N_9519,N_3116,N_4430);
nor U9520 (N_9520,N_4529,N_3691);
nor U9521 (N_9521,N_199,N_575);
or U9522 (N_9522,N_1628,N_3476);
nand U9523 (N_9523,N_1075,N_993);
xor U9524 (N_9524,N_2156,N_4007);
and U9525 (N_9525,N_2168,N_4842);
xnor U9526 (N_9526,N_2919,N_4179);
nand U9527 (N_9527,N_1375,N_890);
nand U9528 (N_9528,N_3257,N_1440);
xor U9529 (N_9529,N_3114,N_1589);
or U9530 (N_9530,N_1453,N_4970);
nand U9531 (N_9531,N_3875,N_769);
and U9532 (N_9532,N_47,N_3166);
nand U9533 (N_9533,N_4520,N_2254);
or U9534 (N_9534,N_1547,N_4859);
nor U9535 (N_9535,N_2290,N_2606);
nand U9536 (N_9536,N_1945,N_4722);
xor U9537 (N_9537,N_4851,N_3576);
xor U9538 (N_9538,N_4999,N_4463);
or U9539 (N_9539,N_920,N_2876);
and U9540 (N_9540,N_4792,N_1932);
nand U9541 (N_9541,N_2413,N_2515);
nand U9542 (N_9542,N_4676,N_3865);
nand U9543 (N_9543,N_4752,N_546);
nand U9544 (N_9544,N_1269,N_1463);
or U9545 (N_9545,N_1642,N_841);
nand U9546 (N_9546,N_97,N_4240);
and U9547 (N_9547,N_3119,N_686);
xnor U9548 (N_9548,N_941,N_4428);
and U9549 (N_9549,N_1087,N_2572);
nand U9550 (N_9550,N_2670,N_2486);
and U9551 (N_9551,N_2722,N_292);
xor U9552 (N_9552,N_1680,N_392);
nor U9553 (N_9553,N_2553,N_3374);
xnor U9554 (N_9554,N_1265,N_4178);
or U9555 (N_9555,N_1782,N_2747);
xnor U9556 (N_9556,N_1498,N_770);
or U9557 (N_9557,N_4611,N_4878);
or U9558 (N_9558,N_1823,N_4727);
or U9559 (N_9559,N_3375,N_4343);
xor U9560 (N_9560,N_2285,N_3219);
nor U9561 (N_9561,N_713,N_106);
and U9562 (N_9562,N_2694,N_4790);
nand U9563 (N_9563,N_3657,N_531);
nor U9564 (N_9564,N_155,N_128);
xor U9565 (N_9565,N_2227,N_2324);
nor U9566 (N_9566,N_2125,N_103);
and U9567 (N_9567,N_1042,N_1146);
or U9568 (N_9568,N_1716,N_2032);
nand U9569 (N_9569,N_2243,N_2599);
or U9570 (N_9570,N_2137,N_2384);
or U9571 (N_9571,N_3947,N_2531);
and U9572 (N_9572,N_4378,N_1828);
or U9573 (N_9573,N_1303,N_2579);
and U9574 (N_9574,N_2881,N_3897);
nand U9575 (N_9575,N_3967,N_2927);
xor U9576 (N_9576,N_2995,N_3945);
or U9577 (N_9577,N_2393,N_1814);
and U9578 (N_9578,N_4291,N_4285);
nor U9579 (N_9579,N_3944,N_4587);
nor U9580 (N_9580,N_1274,N_717);
xor U9581 (N_9581,N_4179,N_3019);
or U9582 (N_9582,N_3042,N_2087);
or U9583 (N_9583,N_2905,N_2888);
or U9584 (N_9584,N_811,N_1108);
nand U9585 (N_9585,N_844,N_4203);
nor U9586 (N_9586,N_563,N_2514);
nor U9587 (N_9587,N_1512,N_2695);
nor U9588 (N_9588,N_97,N_4302);
nor U9589 (N_9589,N_2728,N_2747);
nor U9590 (N_9590,N_3550,N_3887);
xor U9591 (N_9591,N_918,N_154);
or U9592 (N_9592,N_3488,N_507);
nor U9593 (N_9593,N_3152,N_787);
and U9594 (N_9594,N_2559,N_2658);
nand U9595 (N_9595,N_3809,N_1646);
xnor U9596 (N_9596,N_2668,N_4402);
and U9597 (N_9597,N_234,N_3206);
and U9598 (N_9598,N_4332,N_3356);
or U9599 (N_9599,N_619,N_155);
nor U9600 (N_9600,N_2103,N_4360);
nor U9601 (N_9601,N_593,N_2859);
nor U9602 (N_9602,N_499,N_3950);
nand U9603 (N_9603,N_1110,N_2844);
xor U9604 (N_9604,N_2702,N_1417);
nand U9605 (N_9605,N_1683,N_312);
and U9606 (N_9606,N_3923,N_4051);
xnor U9607 (N_9607,N_1249,N_1260);
nor U9608 (N_9608,N_1445,N_3570);
or U9609 (N_9609,N_1334,N_2262);
xor U9610 (N_9610,N_3191,N_2765);
nand U9611 (N_9611,N_1759,N_1037);
and U9612 (N_9612,N_3432,N_3810);
xor U9613 (N_9613,N_3415,N_2321);
nand U9614 (N_9614,N_3600,N_4250);
nand U9615 (N_9615,N_3008,N_255);
nand U9616 (N_9616,N_4368,N_3464);
and U9617 (N_9617,N_2409,N_2341);
nand U9618 (N_9618,N_145,N_3719);
nor U9619 (N_9619,N_523,N_1793);
nand U9620 (N_9620,N_4868,N_4623);
nand U9621 (N_9621,N_2974,N_3978);
nor U9622 (N_9622,N_4626,N_3536);
and U9623 (N_9623,N_2103,N_3616);
and U9624 (N_9624,N_641,N_4262);
or U9625 (N_9625,N_4245,N_530);
nor U9626 (N_9626,N_1068,N_2977);
nor U9627 (N_9627,N_4132,N_216);
nor U9628 (N_9628,N_441,N_2121);
xnor U9629 (N_9629,N_1034,N_2764);
or U9630 (N_9630,N_4665,N_4609);
or U9631 (N_9631,N_4333,N_1972);
or U9632 (N_9632,N_4563,N_820);
or U9633 (N_9633,N_1881,N_2722);
xnor U9634 (N_9634,N_1190,N_3799);
and U9635 (N_9635,N_3715,N_3413);
or U9636 (N_9636,N_4845,N_801);
or U9637 (N_9637,N_2815,N_3247);
nor U9638 (N_9638,N_4665,N_2776);
nor U9639 (N_9639,N_4781,N_4030);
or U9640 (N_9640,N_339,N_345);
nand U9641 (N_9641,N_3996,N_1196);
or U9642 (N_9642,N_4878,N_1710);
xnor U9643 (N_9643,N_2912,N_3779);
and U9644 (N_9644,N_2541,N_4240);
nor U9645 (N_9645,N_2916,N_2773);
nand U9646 (N_9646,N_3887,N_4128);
nand U9647 (N_9647,N_1696,N_1493);
nor U9648 (N_9648,N_3419,N_404);
nor U9649 (N_9649,N_353,N_4456);
xnor U9650 (N_9650,N_2372,N_4479);
or U9651 (N_9651,N_3505,N_2725);
nor U9652 (N_9652,N_4632,N_1588);
nor U9653 (N_9653,N_3525,N_4311);
and U9654 (N_9654,N_1048,N_3346);
nor U9655 (N_9655,N_1734,N_1);
and U9656 (N_9656,N_3257,N_3469);
and U9657 (N_9657,N_337,N_1196);
xnor U9658 (N_9658,N_1340,N_180);
or U9659 (N_9659,N_4808,N_3784);
and U9660 (N_9660,N_624,N_1998);
or U9661 (N_9661,N_4554,N_2426);
xor U9662 (N_9662,N_1352,N_2332);
and U9663 (N_9663,N_2895,N_2372);
and U9664 (N_9664,N_1522,N_1822);
or U9665 (N_9665,N_3452,N_4236);
xnor U9666 (N_9666,N_1276,N_4339);
nor U9667 (N_9667,N_213,N_4400);
and U9668 (N_9668,N_2500,N_2921);
xnor U9669 (N_9669,N_1923,N_355);
or U9670 (N_9670,N_1366,N_3269);
nor U9671 (N_9671,N_2670,N_116);
nor U9672 (N_9672,N_1806,N_531);
nand U9673 (N_9673,N_956,N_1471);
and U9674 (N_9674,N_3548,N_4516);
xnor U9675 (N_9675,N_4258,N_4358);
and U9676 (N_9676,N_3553,N_4938);
nand U9677 (N_9677,N_1773,N_1829);
or U9678 (N_9678,N_2562,N_2106);
nand U9679 (N_9679,N_1368,N_705);
nor U9680 (N_9680,N_1521,N_3041);
xnor U9681 (N_9681,N_2266,N_213);
nand U9682 (N_9682,N_3601,N_3617);
and U9683 (N_9683,N_4740,N_2241);
xor U9684 (N_9684,N_1526,N_352);
nor U9685 (N_9685,N_3608,N_1120);
nand U9686 (N_9686,N_9,N_4319);
and U9687 (N_9687,N_3176,N_3270);
nand U9688 (N_9688,N_1360,N_2081);
nand U9689 (N_9689,N_4560,N_3962);
or U9690 (N_9690,N_496,N_1583);
xnor U9691 (N_9691,N_2364,N_364);
or U9692 (N_9692,N_4824,N_4697);
xnor U9693 (N_9693,N_2376,N_4893);
or U9694 (N_9694,N_1654,N_3583);
nand U9695 (N_9695,N_3495,N_3292);
nand U9696 (N_9696,N_2739,N_2376);
nand U9697 (N_9697,N_1200,N_1556);
nor U9698 (N_9698,N_2055,N_4957);
or U9699 (N_9699,N_2846,N_4125);
xnor U9700 (N_9700,N_3639,N_3134);
and U9701 (N_9701,N_507,N_3586);
and U9702 (N_9702,N_550,N_1515);
xnor U9703 (N_9703,N_4685,N_827);
and U9704 (N_9704,N_2872,N_3934);
nor U9705 (N_9705,N_4557,N_427);
nand U9706 (N_9706,N_3852,N_3601);
or U9707 (N_9707,N_1776,N_4963);
nor U9708 (N_9708,N_2132,N_3405);
and U9709 (N_9709,N_4956,N_4952);
nor U9710 (N_9710,N_1657,N_2793);
xnor U9711 (N_9711,N_648,N_4725);
or U9712 (N_9712,N_1246,N_503);
or U9713 (N_9713,N_2690,N_828);
and U9714 (N_9714,N_3869,N_2504);
and U9715 (N_9715,N_3168,N_1873);
nand U9716 (N_9716,N_1672,N_960);
nor U9717 (N_9717,N_2425,N_3256);
nand U9718 (N_9718,N_660,N_4939);
or U9719 (N_9719,N_3576,N_5);
nor U9720 (N_9720,N_929,N_4064);
and U9721 (N_9721,N_3671,N_2657);
nand U9722 (N_9722,N_4005,N_3348);
nor U9723 (N_9723,N_482,N_4845);
nor U9724 (N_9724,N_1779,N_3950);
and U9725 (N_9725,N_370,N_3494);
nor U9726 (N_9726,N_3470,N_4212);
and U9727 (N_9727,N_1685,N_2500);
nor U9728 (N_9728,N_2413,N_3735);
or U9729 (N_9729,N_3306,N_1283);
xnor U9730 (N_9730,N_2153,N_3534);
or U9731 (N_9731,N_3468,N_987);
nand U9732 (N_9732,N_2887,N_3036);
and U9733 (N_9733,N_1046,N_2759);
nor U9734 (N_9734,N_3044,N_4442);
nor U9735 (N_9735,N_901,N_4395);
or U9736 (N_9736,N_4621,N_4143);
xnor U9737 (N_9737,N_2768,N_2112);
xor U9738 (N_9738,N_4216,N_2925);
and U9739 (N_9739,N_4230,N_2946);
nand U9740 (N_9740,N_3233,N_782);
xor U9741 (N_9741,N_1531,N_1730);
xnor U9742 (N_9742,N_823,N_1163);
and U9743 (N_9743,N_597,N_666);
and U9744 (N_9744,N_3186,N_3842);
nand U9745 (N_9745,N_2880,N_2227);
and U9746 (N_9746,N_4409,N_3835);
nand U9747 (N_9747,N_4087,N_3494);
and U9748 (N_9748,N_1654,N_1081);
or U9749 (N_9749,N_3938,N_1432);
xnor U9750 (N_9750,N_219,N_4436);
and U9751 (N_9751,N_3388,N_4565);
or U9752 (N_9752,N_422,N_1901);
nand U9753 (N_9753,N_3508,N_990);
or U9754 (N_9754,N_3563,N_1241);
nand U9755 (N_9755,N_4596,N_1990);
xor U9756 (N_9756,N_3801,N_4766);
and U9757 (N_9757,N_273,N_1414);
nand U9758 (N_9758,N_798,N_214);
nor U9759 (N_9759,N_1732,N_2591);
xor U9760 (N_9760,N_243,N_4984);
nor U9761 (N_9761,N_3415,N_4361);
xnor U9762 (N_9762,N_3939,N_1517);
nand U9763 (N_9763,N_4663,N_50);
and U9764 (N_9764,N_3591,N_4792);
or U9765 (N_9765,N_4522,N_673);
nand U9766 (N_9766,N_1444,N_205);
nor U9767 (N_9767,N_3590,N_3747);
xor U9768 (N_9768,N_3045,N_802);
nor U9769 (N_9769,N_4693,N_2708);
nand U9770 (N_9770,N_1592,N_4853);
xnor U9771 (N_9771,N_4879,N_2721);
or U9772 (N_9772,N_649,N_3588);
nand U9773 (N_9773,N_4160,N_3347);
nor U9774 (N_9774,N_2714,N_2654);
nor U9775 (N_9775,N_4,N_195);
nor U9776 (N_9776,N_4168,N_1657);
xor U9777 (N_9777,N_1290,N_4789);
nor U9778 (N_9778,N_1050,N_484);
xor U9779 (N_9779,N_1985,N_1795);
or U9780 (N_9780,N_902,N_1084);
xnor U9781 (N_9781,N_2206,N_4112);
xor U9782 (N_9782,N_83,N_3102);
nand U9783 (N_9783,N_1354,N_319);
xor U9784 (N_9784,N_1536,N_820);
or U9785 (N_9785,N_2095,N_3601);
nor U9786 (N_9786,N_4753,N_3008);
nand U9787 (N_9787,N_1756,N_2831);
or U9788 (N_9788,N_2602,N_1578);
nor U9789 (N_9789,N_3956,N_4857);
and U9790 (N_9790,N_4191,N_2909);
and U9791 (N_9791,N_1398,N_1999);
or U9792 (N_9792,N_134,N_870);
xnor U9793 (N_9793,N_2883,N_3550);
and U9794 (N_9794,N_1084,N_1028);
nor U9795 (N_9795,N_4377,N_1109);
nor U9796 (N_9796,N_225,N_1949);
xnor U9797 (N_9797,N_3315,N_35);
and U9798 (N_9798,N_4686,N_2564);
nor U9799 (N_9799,N_1753,N_1599);
and U9800 (N_9800,N_447,N_399);
nor U9801 (N_9801,N_762,N_4304);
xnor U9802 (N_9802,N_3753,N_1675);
nand U9803 (N_9803,N_3193,N_738);
and U9804 (N_9804,N_3785,N_4705);
and U9805 (N_9805,N_172,N_3875);
xor U9806 (N_9806,N_3118,N_4163);
or U9807 (N_9807,N_4610,N_1283);
nor U9808 (N_9808,N_4243,N_122);
and U9809 (N_9809,N_1977,N_2003);
nor U9810 (N_9810,N_2794,N_2372);
nor U9811 (N_9811,N_1511,N_3541);
and U9812 (N_9812,N_226,N_1563);
or U9813 (N_9813,N_60,N_686);
nand U9814 (N_9814,N_63,N_3515);
nand U9815 (N_9815,N_3347,N_4951);
nand U9816 (N_9816,N_3148,N_1495);
nor U9817 (N_9817,N_4044,N_4255);
nand U9818 (N_9818,N_522,N_1532);
and U9819 (N_9819,N_1897,N_4125);
xnor U9820 (N_9820,N_143,N_529);
xor U9821 (N_9821,N_1648,N_3648);
or U9822 (N_9822,N_1600,N_2559);
nand U9823 (N_9823,N_169,N_2931);
nor U9824 (N_9824,N_4376,N_4297);
or U9825 (N_9825,N_1463,N_173);
nand U9826 (N_9826,N_1328,N_3196);
nand U9827 (N_9827,N_759,N_851);
and U9828 (N_9828,N_2004,N_3587);
nor U9829 (N_9829,N_3329,N_50);
or U9830 (N_9830,N_1994,N_2300);
nor U9831 (N_9831,N_3017,N_730);
or U9832 (N_9832,N_2408,N_4236);
nor U9833 (N_9833,N_742,N_2160);
nand U9834 (N_9834,N_1824,N_1744);
and U9835 (N_9835,N_4139,N_2034);
and U9836 (N_9836,N_1039,N_1193);
and U9837 (N_9837,N_3764,N_2131);
nor U9838 (N_9838,N_2146,N_2308);
nand U9839 (N_9839,N_1783,N_4691);
xor U9840 (N_9840,N_277,N_393);
nor U9841 (N_9841,N_3726,N_1667);
and U9842 (N_9842,N_1686,N_268);
or U9843 (N_9843,N_626,N_614);
nand U9844 (N_9844,N_546,N_1055);
and U9845 (N_9845,N_4567,N_2695);
nor U9846 (N_9846,N_4321,N_199);
nor U9847 (N_9847,N_2046,N_3620);
xnor U9848 (N_9848,N_2159,N_2224);
or U9849 (N_9849,N_4750,N_4882);
xnor U9850 (N_9850,N_1878,N_2920);
nand U9851 (N_9851,N_4846,N_1283);
nand U9852 (N_9852,N_3950,N_1876);
or U9853 (N_9853,N_3883,N_208);
and U9854 (N_9854,N_3887,N_3589);
or U9855 (N_9855,N_1595,N_3410);
xor U9856 (N_9856,N_1533,N_2179);
nor U9857 (N_9857,N_1336,N_3823);
nand U9858 (N_9858,N_4685,N_4776);
and U9859 (N_9859,N_1698,N_1940);
xor U9860 (N_9860,N_2568,N_4555);
xor U9861 (N_9861,N_1079,N_579);
or U9862 (N_9862,N_3433,N_2909);
nand U9863 (N_9863,N_4108,N_4717);
or U9864 (N_9864,N_918,N_829);
nor U9865 (N_9865,N_3564,N_4458);
nand U9866 (N_9866,N_3591,N_3794);
nor U9867 (N_9867,N_835,N_4360);
nor U9868 (N_9868,N_2005,N_4716);
nand U9869 (N_9869,N_1116,N_3356);
nor U9870 (N_9870,N_2281,N_4078);
xor U9871 (N_9871,N_3151,N_2936);
nand U9872 (N_9872,N_226,N_2779);
xor U9873 (N_9873,N_4107,N_1304);
nor U9874 (N_9874,N_1836,N_324);
nor U9875 (N_9875,N_4899,N_4941);
nand U9876 (N_9876,N_2916,N_2625);
and U9877 (N_9877,N_4090,N_589);
and U9878 (N_9878,N_4012,N_1446);
and U9879 (N_9879,N_182,N_4660);
or U9880 (N_9880,N_4175,N_2022);
nor U9881 (N_9881,N_1328,N_566);
nor U9882 (N_9882,N_3820,N_1899);
xnor U9883 (N_9883,N_4377,N_2565);
and U9884 (N_9884,N_2750,N_97);
nor U9885 (N_9885,N_947,N_538);
and U9886 (N_9886,N_549,N_3468);
nand U9887 (N_9887,N_1086,N_457);
and U9888 (N_9888,N_2667,N_633);
xnor U9889 (N_9889,N_4009,N_1234);
and U9890 (N_9890,N_2651,N_1186);
and U9891 (N_9891,N_2335,N_4217);
and U9892 (N_9892,N_4310,N_1286);
xnor U9893 (N_9893,N_1378,N_657);
xnor U9894 (N_9894,N_743,N_1056);
nand U9895 (N_9895,N_4172,N_4607);
or U9896 (N_9896,N_4528,N_3721);
and U9897 (N_9897,N_3448,N_84);
or U9898 (N_9898,N_254,N_1215);
nand U9899 (N_9899,N_4253,N_4944);
xnor U9900 (N_9900,N_918,N_728);
nor U9901 (N_9901,N_281,N_2735);
and U9902 (N_9902,N_1186,N_1950);
nor U9903 (N_9903,N_4070,N_4533);
or U9904 (N_9904,N_2373,N_2457);
and U9905 (N_9905,N_882,N_531);
xnor U9906 (N_9906,N_2392,N_1335);
or U9907 (N_9907,N_4798,N_3976);
xor U9908 (N_9908,N_4457,N_836);
or U9909 (N_9909,N_3438,N_2269);
and U9910 (N_9910,N_4409,N_656);
nand U9911 (N_9911,N_3862,N_2855);
nand U9912 (N_9912,N_2913,N_2662);
xor U9913 (N_9913,N_3381,N_1846);
and U9914 (N_9914,N_3626,N_651);
and U9915 (N_9915,N_2619,N_3265);
nand U9916 (N_9916,N_4277,N_1840);
nor U9917 (N_9917,N_1952,N_4654);
nor U9918 (N_9918,N_3755,N_4063);
nand U9919 (N_9919,N_1714,N_1197);
xnor U9920 (N_9920,N_3141,N_3455);
and U9921 (N_9921,N_3375,N_391);
nor U9922 (N_9922,N_2154,N_723);
xor U9923 (N_9923,N_1572,N_2348);
or U9924 (N_9924,N_1442,N_2818);
nand U9925 (N_9925,N_462,N_1504);
xnor U9926 (N_9926,N_673,N_1155);
or U9927 (N_9927,N_2864,N_2430);
nor U9928 (N_9928,N_61,N_3412);
xor U9929 (N_9929,N_2293,N_3154);
xnor U9930 (N_9930,N_3022,N_1262);
or U9931 (N_9931,N_4987,N_1556);
xnor U9932 (N_9932,N_1603,N_3511);
and U9933 (N_9933,N_1489,N_2997);
nand U9934 (N_9934,N_421,N_205);
and U9935 (N_9935,N_2578,N_2387);
xor U9936 (N_9936,N_2099,N_1706);
nor U9937 (N_9937,N_3546,N_2796);
nor U9938 (N_9938,N_2498,N_2133);
xnor U9939 (N_9939,N_1531,N_1788);
and U9940 (N_9940,N_230,N_271);
nand U9941 (N_9941,N_3614,N_4059);
or U9942 (N_9942,N_2850,N_4802);
and U9943 (N_9943,N_4170,N_1114);
xor U9944 (N_9944,N_169,N_4422);
nor U9945 (N_9945,N_654,N_3647);
nand U9946 (N_9946,N_2511,N_2855);
xnor U9947 (N_9947,N_1974,N_1482);
nand U9948 (N_9948,N_4212,N_1755);
xnor U9949 (N_9949,N_846,N_1217);
nor U9950 (N_9950,N_1495,N_4158);
nor U9951 (N_9951,N_3928,N_3563);
or U9952 (N_9952,N_2941,N_3903);
xnor U9953 (N_9953,N_2869,N_1546);
xor U9954 (N_9954,N_1444,N_1835);
nand U9955 (N_9955,N_1333,N_4425);
or U9956 (N_9956,N_1603,N_1463);
and U9957 (N_9957,N_752,N_378);
nor U9958 (N_9958,N_798,N_2991);
nand U9959 (N_9959,N_4575,N_2957);
nor U9960 (N_9960,N_887,N_1406);
nor U9961 (N_9961,N_4611,N_3680);
nand U9962 (N_9962,N_3161,N_347);
nor U9963 (N_9963,N_2389,N_4980);
and U9964 (N_9964,N_2096,N_4642);
xnor U9965 (N_9965,N_3151,N_971);
or U9966 (N_9966,N_1013,N_3903);
xnor U9967 (N_9967,N_3026,N_576);
and U9968 (N_9968,N_133,N_3399);
xnor U9969 (N_9969,N_2911,N_4794);
and U9970 (N_9970,N_4754,N_3628);
nor U9971 (N_9971,N_827,N_1186);
nand U9972 (N_9972,N_2413,N_1345);
or U9973 (N_9973,N_4579,N_2944);
xnor U9974 (N_9974,N_2760,N_4443);
or U9975 (N_9975,N_4959,N_3170);
or U9976 (N_9976,N_693,N_586);
xor U9977 (N_9977,N_2549,N_4206);
and U9978 (N_9978,N_356,N_4340);
nand U9979 (N_9979,N_171,N_4201);
and U9980 (N_9980,N_4090,N_4461);
nor U9981 (N_9981,N_94,N_3706);
nor U9982 (N_9982,N_4589,N_1514);
xnor U9983 (N_9983,N_2089,N_1832);
and U9984 (N_9984,N_4730,N_863);
nand U9985 (N_9985,N_4935,N_4416);
nor U9986 (N_9986,N_1834,N_1022);
nor U9987 (N_9987,N_1555,N_2753);
xnor U9988 (N_9988,N_4781,N_1147);
xnor U9989 (N_9989,N_741,N_4590);
nor U9990 (N_9990,N_2065,N_2474);
or U9991 (N_9991,N_4458,N_4486);
nand U9992 (N_9992,N_2643,N_2268);
nand U9993 (N_9993,N_3004,N_1726);
nor U9994 (N_9994,N_2609,N_1973);
and U9995 (N_9995,N_3599,N_3418);
nand U9996 (N_9996,N_1448,N_2503);
nor U9997 (N_9997,N_1983,N_987);
nor U9998 (N_9998,N_2930,N_2781);
nor U9999 (N_9999,N_3054,N_3803);
nand UO_0 (O_0,N_7558,N_8603);
or UO_1 (O_1,N_8556,N_9915);
nand UO_2 (O_2,N_7545,N_6407);
and UO_3 (O_3,N_5971,N_9125);
nor UO_4 (O_4,N_7457,N_9783);
nand UO_5 (O_5,N_7283,N_6434);
and UO_6 (O_6,N_7003,N_6258);
or UO_7 (O_7,N_6756,N_7293);
or UO_8 (O_8,N_9538,N_7168);
nor UO_9 (O_9,N_5316,N_6737);
nand UO_10 (O_10,N_7284,N_5800);
or UO_11 (O_11,N_6202,N_9093);
or UO_12 (O_12,N_6793,N_6075);
nor UO_13 (O_13,N_7744,N_9818);
nand UO_14 (O_14,N_5348,N_5955);
nand UO_15 (O_15,N_8779,N_6529);
and UO_16 (O_16,N_5718,N_6965);
and UO_17 (O_17,N_7644,N_6521);
and UO_18 (O_18,N_9261,N_7677);
xor UO_19 (O_19,N_9858,N_9657);
or UO_20 (O_20,N_9630,N_6505);
nor UO_21 (O_21,N_9881,N_8503);
xnor UO_22 (O_22,N_7134,N_7932);
nand UO_23 (O_23,N_6106,N_5717);
and UO_24 (O_24,N_6036,N_6244);
nor UO_25 (O_25,N_7204,N_6283);
or UO_26 (O_26,N_8232,N_7456);
xor UO_27 (O_27,N_9515,N_7734);
nor UO_28 (O_28,N_5183,N_9181);
nor UO_29 (O_29,N_9343,N_9859);
and UO_30 (O_30,N_7305,N_6024);
nor UO_31 (O_31,N_7345,N_7935);
xnor UO_32 (O_32,N_7375,N_7026);
nor UO_33 (O_33,N_9432,N_5227);
xnor UO_34 (O_34,N_6555,N_8958);
nand UO_35 (O_35,N_6963,N_7660);
xnor UO_36 (O_36,N_7443,N_7523);
and UO_37 (O_37,N_6859,N_5831);
nand UO_38 (O_38,N_6494,N_9577);
xor UO_39 (O_39,N_6895,N_5456);
xor UO_40 (O_40,N_6575,N_5968);
xor UO_41 (O_41,N_5378,N_8349);
and UO_42 (O_42,N_5861,N_6550);
and UO_43 (O_43,N_6875,N_5808);
and UO_44 (O_44,N_9542,N_9836);
or UO_45 (O_45,N_9211,N_8263);
xnor UO_46 (O_46,N_6676,N_8827);
and UO_47 (O_47,N_7242,N_5337);
or UO_48 (O_48,N_8607,N_9942);
nand UO_49 (O_49,N_6459,N_6304);
or UO_50 (O_50,N_5477,N_7367);
nand UO_51 (O_51,N_7624,N_5763);
or UO_52 (O_52,N_6376,N_8164);
nor UO_53 (O_53,N_5240,N_6138);
xor UO_54 (O_54,N_5068,N_5106);
and UO_55 (O_55,N_9583,N_5233);
or UO_56 (O_56,N_8505,N_7499);
nand UO_57 (O_57,N_6087,N_5375);
xor UO_58 (O_58,N_6047,N_7276);
nor UO_59 (O_59,N_6983,N_6268);
and UO_60 (O_60,N_9418,N_6296);
or UO_61 (O_61,N_5362,N_9987);
nor UO_62 (O_62,N_8359,N_8203);
or UO_63 (O_63,N_7234,N_6705);
and UO_64 (O_64,N_6966,N_7060);
and UO_65 (O_65,N_6804,N_5141);
or UO_66 (O_66,N_9024,N_9914);
or UO_67 (O_67,N_6082,N_5952);
nand UO_68 (O_68,N_5671,N_8942);
nand UO_69 (O_69,N_7550,N_8544);
nor UO_70 (O_70,N_9084,N_9250);
nand UO_71 (O_71,N_6627,N_7172);
and UO_72 (O_72,N_7697,N_5117);
nor UO_73 (O_73,N_7877,N_9719);
and UO_74 (O_74,N_6071,N_8700);
and UO_75 (O_75,N_6226,N_9027);
nor UO_76 (O_76,N_9471,N_5515);
nand UO_77 (O_77,N_6443,N_7822);
nor UO_78 (O_78,N_6158,N_5021);
nor UO_79 (O_79,N_9422,N_6207);
and UO_80 (O_80,N_8636,N_5209);
nand UO_81 (O_81,N_8644,N_6235);
xnor UO_82 (O_82,N_9580,N_7463);
nand UO_83 (O_83,N_7179,N_5653);
or UO_84 (O_84,N_6102,N_9463);
xor UO_85 (O_85,N_9546,N_8864);
nor UO_86 (O_86,N_7974,N_7232);
nand UO_87 (O_87,N_7672,N_9382);
and UO_88 (O_88,N_7622,N_9762);
xnor UO_89 (O_89,N_6372,N_7621);
xor UO_90 (O_90,N_8083,N_9363);
nor UO_91 (O_91,N_5344,N_8385);
nand UO_92 (O_92,N_5751,N_8511);
nor UO_93 (O_93,N_9636,N_9174);
nand UO_94 (O_94,N_5911,N_5343);
nand UO_95 (O_95,N_7696,N_8491);
and UO_96 (O_96,N_5353,N_9681);
and UO_97 (O_97,N_6703,N_7958);
or UO_98 (O_98,N_5255,N_8237);
xnor UO_99 (O_99,N_5903,N_8606);
xnor UO_100 (O_100,N_7640,N_5268);
xor UO_101 (O_101,N_8550,N_6896);
nand UO_102 (O_102,N_5727,N_5184);
nand UO_103 (O_103,N_7175,N_8557);
nand UO_104 (O_104,N_5096,N_9039);
nor UO_105 (O_105,N_8227,N_9133);
xnor UO_106 (O_106,N_9841,N_7404);
and UO_107 (O_107,N_9613,N_7835);
xor UO_108 (O_108,N_7892,N_5230);
or UO_109 (O_109,N_7335,N_5497);
and UO_110 (O_110,N_9145,N_5444);
xnor UO_111 (O_111,N_5140,N_5828);
nand UO_112 (O_112,N_7839,N_8646);
xor UO_113 (O_113,N_5732,N_8535);
or UO_114 (O_114,N_9682,N_6752);
or UO_115 (O_115,N_5246,N_5460);
or UO_116 (O_116,N_5721,N_5894);
and UO_117 (O_117,N_6719,N_5724);
and UO_118 (O_118,N_5495,N_5088);
or UO_119 (O_119,N_9095,N_5790);
nor UO_120 (O_120,N_8726,N_7709);
xnor UO_121 (O_121,N_8185,N_8744);
nor UO_122 (O_122,N_6691,N_6720);
nand UO_123 (O_123,N_9264,N_9869);
nand UO_124 (O_124,N_9609,N_9425);
and UO_125 (O_125,N_8057,N_6284);
or UO_126 (O_126,N_7474,N_8847);
or UO_127 (O_127,N_7011,N_8375);
and UO_128 (O_128,N_6192,N_6103);
nor UO_129 (O_129,N_6753,N_8909);
and UO_130 (O_130,N_9202,N_8436);
and UO_131 (O_131,N_8529,N_5506);
xor UO_132 (O_132,N_8501,N_8920);
and UO_133 (O_133,N_6282,N_5252);
nand UO_134 (O_134,N_6363,N_6344);
or UO_135 (O_135,N_5289,N_5062);
or UO_136 (O_136,N_7799,N_5286);
and UO_137 (O_137,N_8804,N_7140);
nor UO_138 (O_138,N_8515,N_8081);
nor UO_139 (O_139,N_5295,N_8704);
nor UO_140 (O_140,N_5552,N_8386);
nor UO_141 (O_141,N_5758,N_5956);
or UO_142 (O_142,N_8128,N_9431);
and UO_143 (O_143,N_6526,N_5166);
xnor UO_144 (O_144,N_7623,N_8032);
xnor UO_145 (O_145,N_8706,N_7407);
and UO_146 (O_146,N_5779,N_5706);
and UO_147 (O_147,N_7580,N_8985);
or UO_148 (O_148,N_6319,N_6482);
nor UO_149 (O_149,N_9882,N_5725);
xnor UO_150 (O_150,N_8109,N_7586);
and UO_151 (O_151,N_7511,N_8449);
nor UO_152 (O_152,N_9138,N_7092);
xor UO_153 (O_153,N_5984,N_9896);
nand UO_154 (O_154,N_8114,N_5694);
or UO_155 (O_155,N_8536,N_8801);
nand UO_156 (O_156,N_6122,N_5310);
nor UO_157 (O_157,N_5583,N_6923);
xnor UO_158 (O_158,N_9893,N_6311);
or UO_159 (O_159,N_5483,N_9164);
nor UO_160 (O_160,N_7692,N_8599);
xor UO_161 (O_161,N_9777,N_7430);
and UO_162 (O_162,N_7278,N_5195);
xor UO_163 (O_163,N_5652,N_9570);
nand UO_164 (O_164,N_6863,N_8415);
nor UO_165 (O_165,N_9047,N_9077);
nand UO_166 (O_166,N_8200,N_5217);
nand UO_167 (O_167,N_7853,N_6057);
nor UO_168 (O_168,N_6473,N_8568);
nand UO_169 (O_169,N_5294,N_9293);
or UO_170 (O_170,N_7087,N_9224);
nor UO_171 (O_171,N_5990,N_9977);
nor UO_172 (O_172,N_8121,N_6373);
nand UO_173 (O_173,N_9498,N_5681);
xor UO_174 (O_174,N_7567,N_6604);
nor UO_175 (O_175,N_8852,N_6964);
and UO_176 (O_176,N_8082,N_7614);
nand UO_177 (O_177,N_5064,N_8670);
nor UO_178 (O_178,N_6294,N_5816);
xnor UO_179 (O_179,N_5965,N_8444);
xor UO_180 (O_180,N_7553,N_9568);
nor UO_181 (O_181,N_7325,N_5302);
nand UO_182 (O_182,N_9784,N_9409);
or UO_183 (O_183,N_6730,N_6396);
or UO_184 (O_184,N_8475,N_8959);
xor UO_185 (O_185,N_7054,N_8406);
nor UO_186 (O_186,N_5347,N_9140);
nand UO_187 (O_187,N_7450,N_6778);
or UO_188 (O_188,N_9396,N_7669);
or UO_189 (O_189,N_5801,N_8466);
or UO_190 (O_190,N_9287,N_6893);
nor UO_191 (O_191,N_7250,N_7810);
nor UO_192 (O_192,N_7016,N_6325);
nor UO_193 (O_193,N_7532,N_9106);
xor UO_194 (O_194,N_8428,N_6267);
nor UO_195 (O_195,N_9092,N_8149);
nand UO_196 (O_196,N_8350,N_6772);
or UO_197 (O_197,N_8773,N_7044);
or UO_198 (O_198,N_7312,N_5361);
xnor UO_199 (O_199,N_6405,N_9226);
or UO_200 (O_200,N_7682,N_5403);
or UO_201 (O_201,N_9342,N_8970);
nor UO_202 (O_202,N_6647,N_8653);
or UO_203 (O_203,N_6870,N_6779);
or UO_204 (O_204,N_9545,N_5454);
and UO_205 (O_205,N_8565,N_8170);
nor UO_206 (O_206,N_9484,N_5749);
or UO_207 (O_207,N_9800,N_5369);
nor UO_208 (O_208,N_8924,N_5768);
and UO_209 (O_209,N_9497,N_5024);
nor UO_210 (O_210,N_9260,N_8426);
nor UO_211 (O_211,N_7413,N_7362);
nor UO_212 (O_212,N_6040,N_8396);
or UO_213 (O_213,N_7410,N_9427);
and UO_214 (O_214,N_7639,N_7565);
nand UO_215 (O_215,N_5082,N_9237);
or UO_216 (O_216,N_8469,N_5638);
or UO_217 (O_217,N_8727,N_8590);
nand UO_218 (O_218,N_7137,N_9531);
nand UO_219 (O_219,N_7265,N_6404);
nand UO_220 (O_220,N_7593,N_8941);
nor UO_221 (O_221,N_7445,N_9012);
xor UO_222 (O_222,N_6816,N_8492);
nor UO_223 (O_223,N_7793,N_5003);
xnor UO_224 (O_224,N_5983,N_7104);
and UO_225 (O_225,N_8362,N_5323);
xor UO_226 (O_226,N_5623,N_6751);
and UO_227 (O_227,N_9361,N_9816);
xnor UO_228 (O_228,N_5382,N_5013);
and UO_229 (O_229,N_7116,N_9968);
nand UO_230 (O_230,N_7405,N_9117);
xor UO_231 (O_231,N_5224,N_5433);
nor UO_232 (O_232,N_8786,N_8720);
and UO_233 (O_233,N_5381,N_9560);
or UO_234 (O_234,N_9108,N_5469);
xor UO_235 (O_235,N_9627,N_6232);
nand UO_236 (O_236,N_6507,N_5115);
and UO_237 (O_237,N_5969,N_5191);
xnor UO_238 (O_238,N_7679,N_7517);
and UO_239 (O_239,N_5447,N_7957);
nand UO_240 (O_240,N_9973,N_8834);
nor UO_241 (O_241,N_9909,N_7603);
xor UO_242 (O_242,N_7388,N_9519);
nor UO_243 (O_243,N_7315,N_9420);
nand UO_244 (O_244,N_8371,N_7079);
and UO_245 (O_245,N_8662,N_7989);
xnor UO_246 (O_246,N_6116,N_8332);
nor UO_247 (O_247,N_9235,N_9228);
or UO_248 (O_248,N_6672,N_6114);
xor UO_249 (O_249,N_5076,N_9042);
or UO_250 (O_250,N_9258,N_9601);
nor UO_251 (O_251,N_9186,N_8857);
nor UO_252 (O_252,N_9564,N_7149);
or UO_253 (O_253,N_8631,N_9960);
nand UO_254 (O_254,N_8714,N_8269);
xor UO_255 (O_255,N_9240,N_6977);
and UO_256 (O_256,N_5535,N_6320);
xor UO_257 (O_257,N_8889,N_6427);
nor UO_258 (O_258,N_5508,N_8054);
and UO_259 (O_259,N_8004,N_5632);
nor UO_260 (O_260,N_9870,N_6852);
nand UO_261 (O_261,N_9689,N_5054);
and UO_262 (O_262,N_7427,N_6257);
or UO_263 (O_263,N_8302,N_7601);
nor UO_264 (O_264,N_7887,N_6222);
or UO_265 (O_265,N_9862,N_9459);
nor UO_266 (O_266,N_8322,N_6901);
and UO_267 (O_267,N_7409,N_9056);
nor UO_268 (O_268,N_6446,N_6322);
nor UO_269 (O_269,N_7904,N_7566);
nand UO_270 (O_270,N_6805,N_8575);
and UO_271 (O_271,N_9465,N_8880);
nor UO_272 (O_272,N_7326,N_6948);
nand UO_273 (O_273,N_7711,N_5668);
xnor UO_274 (O_274,N_5683,N_9906);
nor UO_275 (O_275,N_7502,N_8453);
nor UO_276 (O_276,N_8329,N_5980);
nand UO_277 (O_277,N_5078,N_9407);
or UO_278 (O_278,N_7902,N_7392);
and UO_279 (O_279,N_6472,N_6261);
and UO_280 (O_280,N_9007,N_7266);
nor UO_281 (O_281,N_8791,N_8497);
and UO_282 (O_282,N_8957,N_8474);
nand UO_283 (O_283,N_7371,N_6408);
nor UO_284 (O_284,N_9304,N_7687);
or UO_285 (O_285,N_7896,N_5185);
and UO_286 (O_286,N_7590,N_8451);
and UO_287 (O_287,N_5452,N_5429);
xor UO_288 (O_288,N_9227,N_5415);
nand UO_289 (O_289,N_9511,N_9175);
xnor UO_290 (O_290,N_9879,N_7770);
or UO_291 (O_291,N_8023,N_6733);
xnor UO_292 (O_292,N_9825,N_8418);
nand UO_293 (O_293,N_5593,N_6783);
xor UO_294 (O_294,N_9899,N_5026);
xnor UO_295 (O_295,N_8947,N_7815);
nor UO_296 (O_296,N_9050,N_5607);
or UO_297 (O_297,N_6740,N_8261);
nand UO_298 (O_298,N_5693,N_7122);
nand UO_299 (O_299,N_9089,N_7438);
nand UO_300 (O_300,N_8611,N_8733);
xor UO_301 (O_301,N_7100,N_7535);
or UO_302 (O_302,N_6142,N_9521);
nor UO_303 (O_303,N_8698,N_9058);
or UO_304 (O_304,N_9925,N_8678);
and UO_305 (O_305,N_9127,N_9004);
xnor UO_306 (O_306,N_9450,N_6287);
xor UO_307 (O_307,N_7806,N_7006);
and UO_308 (O_308,N_9944,N_5085);
nor UO_309 (O_309,N_9219,N_7331);
nor UO_310 (O_310,N_7950,N_6097);
and UO_311 (O_311,N_6072,N_8305);
xnor UO_312 (O_312,N_8117,N_5170);
nor UO_313 (O_313,N_5007,N_7396);
xnor UO_314 (O_314,N_7509,N_9773);
and UO_315 (O_315,N_8602,N_9806);
nand UO_316 (O_316,N_7494,N_7224);
xnor UO_317 (O_317,N_7740,N_5346);
or UO_318 (O_318,N_9085,N_6984);
xor UO_319 (O_319,N_7609,N_6198);
xnor UO_320 (O_320,N_5852,N_7662);
nor UO_321 (O_321,N_6713,N_8110);
nand UO_322 (O_322,N_9540,N_8309);
nand UO_323 (O_323,N_9703,N_6646);
nor UO_324 (O_324,N_5893,N_7563);
or UO_325 (O_325,N_8553,N_5993);
nand UO_326 (O_326,N_8000,N_5863);
and UO_327 (O_327,N_7454,N_5954);
xnor UO_328 (O_328,N_8092,N_9404);
nor UO_329 (O_329,N_5891,N_8682);
and UO_330 (O_330,N_8868,N_6967);
xnor UO_331 (O_331,N_9435,N_9638);
xnor UO_332 (O_332,N_6310,N_5488);
nor UO_333 (O_333,N_8899,N_6468);
and UO_334 (O_334,N_8666,N_7749);
and UO_335 (O_335,N_5487,N_9365);
nand UO_336 (O_336,N_8910,N_8932);
nor UO_337 (O_337,N_8691,N_7024);
nand UO_338 (O_338,N_6490,N_9417);
nand UO_339 (O_339,N_5935,N_8738);
and UO_340 (O_340,N_9743,N_7508);
and UO_341 (O_341,N_5778,N_6280);
and UO_342 (O_342,N_8367,N_7214);
and UO_343 (O_343,N_7169,N_9552);
nor UO_344 (O_344,N_7894,N_8231);
xnor UO_345 (O_345,N_5102,N_9029);
nor UO_346 (O_346,N_6834,N_9464);
nor UO_347 (O_347,N_5280,N_5155);
or UO_348 (O_348,N_6259,N_7598);
xnor UO_349 (O_349,N_9372,N_9754);
xnor UO_350 (O_350,N_7258,N_8245);
and UO_351 (O_351,N_7050,N_9648);
nor UO_352 (O_352,N_5850,N_9895);
xor UO_353 (O_353,N_5145,N_6383);
or UO_354 (O_354,N_5922,N_7285);
xor UO_355 (O_355,N_9852,N_9939);
or UO_356 (O_356,N_5226,N_8326);
xor UO_357 (O_357,N_5216,N_7471);
or UO_358 (O_358,N_9533,N_7606);
or UO_359 (O_359,N_6039,N_6237);
and UO_360 (O_360,N_5719,N_8554);
and UO_361 (O_361,N_8413,N_9478);
nor UO_362 (O_362,N_5074,N_7260);
nor UO_363 (O_363,N_7656,N_9194);
nand UO_364 (O_364,N_5655,N_5159);
or UO_365 (O_365,N_9082,N_5410);
nor UO_366 (O_366,N_6542,N_8095);
or UO_367 (O_367,N_7238,N_9146);
or UO_368 (O_368,N_7647,N_7244);
or UO_369 (O_369,N_5304,N_9709);
xnor UO_370 (O_370,N_9327,N_9930);
xnor UO_371 (O_371,N_5613,N_5776);
nand UO_372 (O_372,N_8838,N_9843);
and UO_373 (O_373,N_6374,N_7383);
nor UO_374 (O_374,N_7397,N_9733);
xnor UO_375 (O_375,N_7648,N_5777);
nor UO_376 (O_376,N_5449,N_6506);
or UO_377 (O_377,N_7714,N_6439);
and UO_378 (O_378,N_8201,N_5962);
or UO_379 (O_379,N_8085,N_6866);
or UO_380 (O_380,N_6458,N_5888);
or UO_381 (O_381,N_9461,N_9584);
or UO_382 (O_382,N_5597,N_7123);
or UO_383 (O_383,N_5210,N_6327);
xor UO_384 (O_384,N_5715,N_8494);
xnor UO_385 (O_385,N_5061,N_5791);
nand UO_386 (O_386,N_9107,N_5782);
nor UO_387 (O_387,N_9634,N_6229);
xor UO_388 (O_388,N_5122,N_6958);
and UO_389 (O_389,N_6519,N_8605);
or UO_390 (O_390,N_5988,N_8132);
nand UO_391 (O_391,N_7372,N_9005);
xor UO_392 (O_392,N_6307,N_7190);
and UO_393 (O_393,N_9926,N_9506);
or UO_394 (O_394,N_7948,N_6791);
or UO_395 (O_395,N_9848,N_7009);
and UO_396 (O_396,N_7757,N_7534);
nand UO_397 (O_397,N_7066,N_9656);
nor UO_398 (O_398,N_5237,N_7222);
xnor UO_399 (O_399,N_9362,N_8835);
nand UO_400 (O_400,N_5635,N_6652);
or UO_401 (O_401,N_6828,N_7448);
nor UO_402 (O_402,N_5656,N_7747);
nor UO_403 (O_403,N_6137,N_5697);
xnor UO_404 (O_404,N_6455,N_8171);
nor UO_405 (O_405,N_9707,N_9751);
or UO_406 (O_406,N_7097,N_6044);
and UO_407 (O_407,N_6346,N_6079);
nand UO_408 (O_408,N_5580,N_5396);
or UO_409 (O_409,N_5817,N_9466);
nor UO_410 (O_410,N_6509,N_6941);
or UO_411 (O_411,N_7529,N_5463);
nor UO_412 (O_412,N_5603,N_7281);
nor UO_413 (O_413,N_5890,N_9713);
and UO_414 (O_414,N_6127,N_5376);
nor UO_415 (O_415,N_6350,N_8102);
and UO_416 (O_416,N_9157,N_7798);
nand UO_417 (O_417,N_6370,N_9026);
nor UO_418 (O_418,N_7683,N_8182);
xor UO_419 (O_419,N_9485,N_7086);
xor UO_420 (O_420,N_6803,N_7181);
nor UO_421 (O_421,N_8650,N_9332);
or UO_422 (O_422,N_7012,N_5957);
nor UO_423 (O_423,N_6820,N_9513);
and UO_424 (O_424,N_7642,N_6491);
and UO_425 (O_425,N_8377,N_5498);
nand UO_426 (O_426,N_7288,N_5908);
xor UO_427 (O_427,N_5046,N_6512);
or UO_428 (O_428,N_6292,N_7488);
and UO_429 (O_429,N_8851,N_7843);
nor UO_430 (O_430,N_7318,N_6418);
and UO_431 (O_431,N_8627,N_6077);
nand UO_432 (O_432,N_9172,N_9000);
or UO_433 (O_433,N_9999,N_5909);
xor UO_434 (O_434,N_6868,N_9724);
nand UO_435 (O_435,N_8198,N_6438);
nor UO_436 (O_436,N_7282,N_5540);
nor UO_437 (O_437,N_6080,N_5242);
nor UO_438 (O_438,N_9112,N_9440);
nor UO_439 (O_439,N_5641,N_9400);
nor UO_440 (O_440,N_5996,N_7072);
xnor UO_441 (O_441,N_5176,N_8380);
xor UO_442 (O_442,N_7869,N_7710);
xor UO_443 (O_443,N_9855,N_8897);
nand UO_444 (O_444,N_6798,N_5009);
nor UO_445 (O_445,N_7490,N_6628);
or UO_446 (O_446,N_8809,N_6019);
xnor UO_447 (O_447,N_6243,N_8832);
and UO_448 (O_448,N_8010,N_9347);
nand UO_449 (O_449,N_9416,N_6933);
xor UO_450 (O_450,N_9982,N_6994);
xnor UO_451 (O_451,N_7889,N_8640);
xnor UO_452 (O_452,N_7029,N_6504);
or UO_453 (O_453,N_6821,N_6096);
xnor UO_454 (O_454,N_7854,N_7241);
nor UO_455 (O_455,N_8630,N_7154);
and UO_456 (O_456,N_5841,N_6525);
or UO_457 (O_457,N_6986,N_7167);
or UO_458 (O_458,N_5199,N_6641);
or UO_459 (O_459,N_5946,N_6135);
nand UO_460 (O_460,N_9201,N_7139);
xor UO_461 (O_461,N_6501,N_5357);
xnor UO_462 (O_462,N_8808,N_6050);
xnor UO_463 (O_463,N_5398,N_8190);
xnor UO_464 (O_464,N_7256,N_7755);
and UO_465 (O_465,N_7068,N_9500);
xnor UO_466 (O_466,N_5005,N_8900);
and UO_467 (O_467,N_9120,N_8452);
xnor UO_468 (O_468,N_7743,N_6007);
and UO_469 (O_469,N_8041,N_9282);
or UO_470 (O_470,N_5854,N_5292);
xor UO_471 (O_471,N_7340,N_9063);
or UO_472 (O_472,N_7215,N_5278);
and UO_473 (O_473,N_6643,N_7758);
and UO_474 (O_474,N_9017,N_7965);
or UO_475 (O_475,N_9814,N_9367);
nand UO_476 (O_476,N_9436,N_7344);
nand UO_477 (O_477,N_7390,N_9673);
xnor UO_478 (O_478,N_8181,N_5358);
xor UO_479 (O_479,N_8915,N_9649);
or UO_480 (O_480,N_6763,N_6581);
and UO_481 (O_481,N_6183,N_6131);
or UO_482 (O_482,N_9065,N_8267);
or UO_483 (O_483,N_9241,N_8712);
and UO_484 (O_484,N_5360,N_8867);
xor UO_485 (O_485,N_9394,N_9156);
and UO_486 (O_486,N_9428,N_5423);
and UO_487 (O_487,N_9520,N_8099);
nand UO_488 (O_488,N_6236,N_8879);
nor UO_489 (O_489,N_5943,N_6379);
or UO_490 (O_490,N_5900,N_8414);
or UO_491 (O_491,N_7401,N_9062);
and UO_492 (O_492,N_5862,N_6864);
xor UO_493 (O_493,N_9932,N_9616);
or UO_494 (O_494,N_6926,N_7916);
or UO_495 (O_495,N_7394,N_8003);
xnor UO_496 (O_496,N_5529,N_5156);
nand UO_497 (O_497,N_8677,N_7129);
or UO_498 (O_498,N_7855,N_7653);
or UO_499 (O_499,N_6785,N_5002);
and UO_500 (O_500,N_5544,N_9765);
nand UO_501 (O_501,N_6649,N_7389);
nor UO_502 (O_502,N_9745,N_9864);
xnor UO_503 (O_503,N_6709,N_7062);
xnor UO_504 (O_504,N_6590,N_9737);
nand UO_505 (O_505,N_9742,N_6343);
nand UO_506 (O_506,N_5814,N_6188);
xor UO_507 (O_507,N_6475,N_6004);
or UO_508 (O_508,N_5491,N_8323);
nor UO_509 (O_509,N_5945,N_9946);
xnor UO_510 (O_510,N_5300,N_5069);
xor UO_511 (O_511,N_6148,N_8746);
xnor UO_512 (O_512,N_9602,N_6599);
xnor UO_513 (O_513,N_9614,N_5703);
xnor UO_514 (O_514,N_7570,N_6238);
nor UO_515 (O_515,N_7551,N_7299);
nand UO_516 (O_516,N_8612,N_5206);
nand UO_517 (O_517,N_8710,N_5431);
and UO_518 (O_518,N_5179,N_9665);
xnor UO_519 (O_519,N_6605,N_5244);
nand UO_520 (O_520,N_7088,N_8719);
xor UO_521 (O_521,N_6000,N_9650);
nand UO_522 (O_522,N_5605,N_8660);
xor UO_523 (O_523,N_5386,N_9104);
or UO_524 (O_524,N_8243,N_8353);
xnor UO_525 (O_525,N_9664,N_7143);
and UO_526 (O_526,N_5025,N_8446);
xor UO_527 (O_527,N_8308,N_5476);
xor UO_528 (O_528,N_6483,N_8280);
nand UO_529 (O_529,N_8366,N_6128);
nand UO_530 (O_530,N_8688,N_8999);
xnor UO_531 (O_531,N_6832,N_8388);
nand UO_532 (O_532,N_5550,N_8150);
and UO_533 (O_533,N_6220,N_7317);
nand UO_534 (O_534,N_9662,N_8140);
and UO_535 (O_535,N_6115,N_5404);
and UO_536 (O_536,N_8675,N_5480);
or UO_537 (O_537,N_8137,N_5896);
xor UO_538 (O_538,N_7987,N_6091);
and UO_539 (O_539,N_9277,N_5519);
nand UO_540 (O_540,N_8352,N_5615);
xnor UO_541 (O_541,N_5824,N_6945);
nor UO_542 (O_542,N_7650,N_7788);
nor UO_543 (O_543,N_7807,N_5688);
xor UO_544 (O_544,N_9061,N_7671);
nand UO_545 (O_545,N_9988,N_6887);
and UO_546 (O_546,N_7866,N_6629);
nand UO_547 (O_547,N_7604,N_8304);
or UO_548 (O_548,N_5496,N_9953);
or UO_549 (O_549,N_6888,N_9596);
nor UO_550 (O_550,N_5915,N_6873);
and UO_551 (O_551,N_9034,N_7360);
nor UO_552 (O_552,N_6732,N_9354);
and UO_553 (O_553,N_5760,N_6161);
or UO_554 (O_554,N_9376,N_7247);
nor UO_555 (O_555,N_6189,N_8513);
and UO_556 (O_556,N_5739,N_6683);
nand UO_557 (O_557,N_5363,N_9317);
xnor UO_558 (O_558,N_7699,N_7103);
nor UO_559 (O_559,N_7795,N_9177);
or UO_560 (O_560,N_8577,N_8158);
or UO_561 (O_561,N_5055,N_5040);
nand UO_562 (O_562,N_6203,N_8314);
nor UO_563 (O_563,N_7975,N_8508);
and UO_564 (O_564,N_6130,N_9847);
and UO_565 (O_565,N_7995,N_7479);
xnor UO_566 (O_566,N_9688,N_9898);
xnor UO_567 (O_567,N_6602,N_7596);
and UO_568 (O_568,N_5475,N_5329);
nand UO_569 (O_569,N_9041,N_6855);
xor UO_570 (O_570,N_6069,N_6829);
xnor UO_571 (O_571,N_9183,N_5031);
and UO_572 (O_572,N_9014,N_6240);
nor UO_573 (O_573,N_7880,N_7579);
or UO_574 (O_574,N_9647,N_7000);
and UO_575 (O_575,N_9487,N_5081);
or UO_576 (O_576,N_9644,N_7186);
nand UO_577 (O_577,N_9828,N_6939);
xor UO_578 (O_578,N_6700,N_8430);
nand UO_579 (O_579,N_5175,N_8890);
nand UO_580 (O_580,N_5516,N_7264);
and UO_581 (O_581,N_8582,N_8215);
or UO_582 (O_582,N_6754,N_5419);
nor UO_583 (O_583,N_5033,N_7582);
nor UO_584 (O_584,N_9299,N_8504);
or UO_585 (O_585,N_9496,N_5644);
xnor UO_586 (O_586,N_6715,N_7901);
nor UO_587 (O_587,N_8806,N_5425);
xnor UO_588 (O_588,N_7059,N_9198);
nand UO_589 (O_589,N_8763,N_8324);
xnor UO_590 (O_590,N_7617,N_6360);
nand UO_591 (O_591,N_6487,N_8836);
nor UO_592 (O_592,N_8254,N_8405);
or UO_593 (O_593,N_9470,N_9245);
and UO_594 (O_594,N_5836,N_5079);
and UO_595 (O_595,N_7912,N_9025);
nand UO_596 (O_596,N_5557,N_6375);
or UO_597 (O_597,N_7436,N_7411);
or UO_598 (O_598,N_7920,N_8142);
or UO_599 (O_599,N_8026,N_8252);
nand UO_600 (O_600,N_5336,N_8271);
xnor UO_601 (O_601,N_8044,N_7393);
nand UO_602 (O_602,N_9929,N_8333);
and UO_603 (O_603,N_9251,N_8233);
nor UO_604 (O_604,N_8716,N_5913);
nor UO_605 (O_605,N_6095,N_6789);
or UO_606 (O_606,N_7047,N_8355);
nand UO_607 (O_607,N_8528,N_5250);
nor UO_608 (O_608,N_9414,N_6324);
or UO_609 (O_609,N_8619,N_9706);
or UO_610 (O_610,N_6801,N_9099);
nand UO_611 (O_611,N_5786,N_8434);
xnor UO_612 (O_612,N_9965,N_9415);
nand UO_613 (O_613,N_9865,N_6213);
nor UO_614 (O_614,N_7584,N_6671);
and UO_615 (O_615,N_5874,N_8509);
xor UO_616 (O_616,N_9801,N_7437);
nand UO_617 (O_617,N_9348,N_9406);
nand UO_618 (O_618,N_9980,N_5421);
xnor UO_619 (O_619,N_6347,N_7246);
or UO_620 (O_620,N_5049,N_6462);
and UO_621 (O_621,N_9957,N_9811);
nor UO_622 (O_622,N_8319,N_5245);
and UO_623 (O_623,N_6706,N_5505);
nor UO_624 (O_624,N_5400,N_5372);
xor UO_625 (O_625,N_6766,N_5462);
nor UO_626 (O_626,N_7402,N_5568);
nor UO_627 (O_627,N_6639,N_6083);
or UO_628 (O_628,N_7626,N_6495);
nor UO_629 (O_629,N_8580,N_6934);
nor UO_630 (O_630,N_7826,N_8107);
or UO_631 (O_631,N_5636,N_5684);
nand UO_632 (O_632,N_7001,N_8928);
or UO_633 (O_633,N_5335,N_5424);
and UO_634 (O_634,N_8939,N_7196);
nor UO_635 (O_635,N_7296,N_7441);
and UO_636 (O_636,N_7133,N_9433);
and UO_637 (O_637,N_8740,N_9747);
nand UO_638 (O_638,N_7585,N_6787);
and UO_639 (O_639,N_8306,N_5877);
and UO_640 (O_640,N_7841,N_6699);
nor UO_641 (O_641,N_7461,N_5364);
nand UO_642 (O_642,N_6904,N_5273);
nand UO_643 (O_643,N_7633,N_5522);
nor UO_644 (O_644,N_6498,N_8667);
xor UO_645 (O_645,N_9494,N_8755);
xnor UO_646 (O_646,N_9890,N_5793);
and UO_647 (O_647,N_6972,N_9071);
nor UO_648 (O_648,N_7121,N_5309);
or UO_649 (O_649,N_7829,N_9397);
nor UO_650 (O_650,N_6354,N_6151);
or UO_651 (O_651,N_9995,N_7497);
xor UO_652 (O_652,N_5172,N_5880);
nor UO_653 (O_653,N_9476,N_7185);
nand UO_654 (O_654,N_9646,N_7794);
or UO_655 (O_655,N_8729,N_6393);
or UO_656 (O_656,N_7953,N_8934);
and UO_657 (O_657,N_5875,N_9854);
or UO_658 (O_658,N_8094,N_9792);
nand UO_659 (O_659,N_8984,N_8223);
or UO_660 (O_660,N_5333,N_9607);
and UO_661 (O_661,N_6761,N_5869);
nand UO_662 (O_662,N_8439,N_6725);
xnor UO_663 (O_663,N_6293,N_5670);
nor UO_664 (O_664,N_7162,N_6056);
or UO_665 (O_665,N_8061,N_5241);
nor UO_666 (O_666,N_5118,N_7057);
or UO_667 (O_667,N_7205,N_6686);
xnor UO_668 (O_668,N_8588,N_8848);
nor UO_669 (O_669,N_5177,N_9098);
xor UO_670 (O_670,N_8211,N_7249);
nand UO_671 (O_671,N_9639,N_5264);
or UO_672 (O_672,N_8901,N_9022);
and UO_673 (O_673,N_7304,N_8265);
or UO_674 (O_674,N_9381,N_5402);
nand UO_675 (O_675,N_8351,N_9730);
xor UO_676 (O_676,N_9267,N_9375);
and UO_677 (O_677,N_5734,N_6854);
nor UO_678 (O_678,N_8495,N_6367);
nand UO_679 (O_679,N_8814,N_9243);
nand UO_680 (O_680,N_5663,N_6982);
and UO_681 (O_681,N_6398,N_9233);
nand UO_682 (O_682,N_5640,N_5783);
or UO_683 (O_683,N_5723,N_8933);
and UO_684 (O_684,N_5190,N_8663);
or UO_685 (O_685,N_6613,N_9611);
xor UO_686 (O_686,N_6065,N_6260);
nor UO_687 (O_687,N_9402,N_7988);
or UO_688 (O_688,N_8597,N_8093);
and UO_689 (O_689,N_8708,N_5279);
and UO_690 (O_690,N_6086,N_9386);
or UO_691 (O_691,N_6084,N_6922);
xor UO_692 (O_692,N_5293,N_5059);
nand UO_693 (O_693,N_9907,N_8338);
nand UO_694 (O_694,N_9312,N_7102);
xor UO_695 (O_695,N_6831,N_8046);
xor UO_696 (O_696,N_6824,N_8432);
or UO_697 (O_697,N_9323,N_8074);
xnor UO_698 (O_698,N_9249,N_8674);
nand UO_699 (O_699,N_8135,N_9573);
xnor UO_700 (O_700,N_5765,N_8282);
xor UO_701 (O_701,N_8387,N_5370);
or UO_702 (O_702,N_8295,N_6362);
or UO_703 (O_703,N_5753,N_8221);
and UO_704 (O_704,N_7659,N_5467);
and UO_705 (O_705,N_8645,N_7472);
nor UO_706 (O_706,N_8722,N_9011);
nor UO_707 (O_707,N_6841,N_8840);
xnor UO_708 (O_708,N_8078,N_8457);
nand UO_709 (O_709,N_7130,N_5892);
xor UO_710 (O_710,N_9588,N_6206);
and UO_711 (O_711,N_8757,N_6270);
nand UO_712 (O_712,N_9271,N_6835);
or UO_713 (O_713,N_9575,N_5471);
xnor UO_714 (O_714,N_7684,N_6334);
or UO_715 (O_715,N_9144,N_9234);
nor UO_716 (O_716,N_6470,N_6523);
nor UO_717 (O_717,N_7192,N_7010);
xor UO_718 (O_718,N_9244,N_5039);
nand UO_719 (O_719,N_8956,N_6176);
and UO_720 (O_720,N_8736,N_9892);
and UO_721 (O_721,N_8454,N_9265);
or UO_722 (O_722,N_8618,N_5525);
nor UO_723 (O_723,N_9385,N_8825);
xor UO_724 (O_724,N_5116,N_7608);
or UO_725 (O_725,N_9955,N_7182);
or UO_726 (O_726,N_5676,N_6825);
or UO_727 (O_727,N_8166,N_9242);
or UO_728 (O_728,N_9252,N_7198);
and UO_729 (O_729,N_8772,N_6291);
xor UO_730 (O_730,N_6061,N_6997);
nor UO_731 (O_731,N_6777,N_6516);
nand UO_732 (O_732,N_9727,N_5647);
or UO_733 (O_733,N_6100,N_9516);
or UO_734 (O_734,N_9246,N_6927);
or UO_735 (O_735,N_6015,N_8013);
nand UO_736 (O_736,N_7952,N_9308);
nand UO_737 (O_737,N_5413,N_7765);
nor UO_738 (O_738,N_5365,N_6837);
or UO_739 (O_739,N_9997,N_8205);
xnor UO_740 (O_740,N_5189,N_6246);
xnor UO_741 (O_741,N_9578,N_8226);
and UO_742 (O_742,N_5944,N_5555);
nor UO_743 (O_743,N_7576,N_5157);
nand UO_744 (O_744,N_6537,N_7673);
and UO_745 (O_745,N_8395,N_7336);
xor UO_746 (O_746,N_7197,N_5111);
or UO_747 (O_747,N_8876,N_6799);
nor UO_748 (O_748,N_5705,N_7374);
nor UO_749 (O_749,N_8229,N_7191);
nor UO_750 (O_750,N_7809,N_6136);
nor UO_751 (O_751,N_6794,N_9971);
or UO_752 (O_752,N_6768,N_9849);
xor UO_753 (O_753,N_8989,N_7984);
nand UO_754 (O_754,N_6696,N_6878);
nor UO_755 (O_755,N_8202,N_5368);
nor UO_756 (O_756,N_6656,N_6143);
nor UO_757 (O_757,N_5503,N_9162);
and UO_758 (O_758,N_6366,N_6250);
xor UO_759 (O_759,N_8649,N_9621);
nand UO_760 (O_760,N_5764,N_5517);
nor UO_761 (O_761,N_6570,N_5281);
nand UO_762 (O_762,N_9839,N_9370);
and UO_763 (O_763,N_7439,N_9043);
or UO_764 (O_764,N_8507,N_5991);
nor UO_765 (O_765,N_8853,N_5110);
nor UO_766 (O_766,N_6955,N_8419);
and UO_767 (O_767,N_5205,N_7594);
nor UO_768 (O_768,N_8256,N_7261);
nand UO_769 (O_769,N_7459,N_9006);
or UO_770 (O_770,N_7842,N_7994);
and UO_771 (O_771,N_8241,N_6078);
nor UO_772 (O_772,N_9272,N_8642);
nand UO_773 (O_773,N_8455,N_9097);
xnor UO_774 (O_774,N_9785,N_8165);
xnor UO_775 (O_775,N_7732,N_7833);
xnor UO_776 (O_776,N_5838,N_6755);
xnor UO_777 (O_777,N_8178,N_5695);
and UO_778 (O_778,N_5269,N_5964);
nand UO_779 (O_779,N_7373,N_6481);
nor UO_780 (O_780,N_6478,N_5091);
and UO_781 (O_781,N_7520,N_7379);
or UO_782 (O_782,N_6630,N_5698);
and UO_783 (O_783,N_5129,N_6544);
and UO_784 (O_784,N_8358,N_5243);
and UO_785 (O_785,N_6074,N_6530);
nand UO_786 (O_786,N_9548,N_9458);
and UO_787 (O_787,N_7306,N_7236);
xor UO_788 (O_788,N_7754,N_9586);
nor UO_789 (O_789,N_9390,N_8823);
xnor UO_790 (O_790,N_6191,N_7161);
nand UO_791 (O_791,N_7366,N_5099);
xor UO_792 (O_792,N_9209,N_6125);
xor UO_793 (O_793,N_6022,N_6853);
xnor UO_794 (O_794,N_6441,N_8068);
and UO_795 (O_795,N_5796,N_8480);
and UO_796 (O_796,N_5821,N_8368);
or UO_797 (O_797,N_8782,N_9756);
nor UO_798 (O_798,N_8713,N_6574);
and UO_799 (O_799,N_7923,N_5648);
nand UO_800 (O_800,N_8356,N_7209);
or UO_801 (O_801,N_9060,N_5173);
and UO_802 (O_802,N_5262,N_6173);
xnor UO_803 (O_803,N_9118,N_8517);
xor UO_804 (O_804,N_8979,N_6577);
or UO_805 (O_805,N_9598,N_5482);
nor UO_806 (O_806,N_6957,N_8391);
and UO_807 (O_807,N_7195,N_7082);
or UO_808 (O_808,N_6865,N_9148);
nand UO_809 (O_809,N_7476,N_8296);
nand UO_810 (O_810,N_5626,N_9030);
nor UO_811 (O_811,N_7681,N_8163);
nand UO_812 (O_812,N_6698,N_8703);
xnor UO_813 (O_813,N_8908,N_7495);
nand UO_814 (O_814,N_9693,N_9655);
nor UO_815 (O_815,N_9923,N_8931);
or UO_816 (O_816,N_5766,N_6018);
or UO_817 (O_817,N_5928,N_7462);
and UO_818 (O_818,N_8512,N_5354);
nor UO_819 (O_819,N_9191,N_8950);
nand UO_820 (O_820,N_9820,N_7717);
and UO_821 (O_821,N_9579,N_7334);
xnor UO_822 (O_822,N_6159,N_8489);
or UO_823 (O_823,N_7176,N_8143);
or UO_824 (O_824,N_6133,N_8621);
nand UO_825 (O_825,N_6118,N_5665);
or UO_826 (O_826,N_9447,N_9696);
nor UO_827 (O_827,N_8214,N_5267);
nor UO_828 (O_828,N_6935,N_5614);
or UO_829 (O_829,N_8297,N_8753);
nor UO_830 (O_830,N_8364,N_8547);
xor UO_831 (O_831,N_8087,N_6012);
nor UO_832 (O_832,N_8342,N_7051);
nor UO_833 (O_833,N_5097,N_5601);
nor UO_834 (O_834,N_7248,N_8303);
and UO_835 (O_835,N_7227,N_6818);
and UO_836 (O_836,N_5967,N_7480);
or UO_837 (O_837,N_8610,N_8278);
or UO_838 (O_838,N_6514,N_6782);
nor UO_839 (O_839,N_6005,N_9993);
and UO_840 (O_840,N_8327,N_8673);
xor UO_841 (O_841,N_6266,N_6230);
or UO_842 (O_842,N_6060,N_6090);
or UO_843 (O_843,N_7339,N_9532);
nand UO_844 (O_844,N_6353,N_7171);
xnor UO_845 (O_845,N_8113,N_8532);
and UO_846 (O_846,N_9597,N_8522);
or UO_847 (O_847,N_5860,N_8381);
or UO_848 (O_848,N_7310,N_6850);
nor UO_849 (O_849,N_8986,N_8994);
nand UO_850 (O_850,N_5422,N_5263);
and UO_851 (O_851,N_8052,N_6085);
nand UO_852 (O_852,N_5214,N_9349);
xnor UO_853 (O_853,N_8191,N_6345);
nand UO_854 (O_854,N_6338,N_9918);
nand UO_855 (O_855,N_8794,N_7473);
nand UO_856 (O_856,N_9631,N_8861);
or UO_857 (O_857,N_7893,N_7023);
and UO_858 (O_858,N_6606,N_8021);
or UO_859 (O_859,N_8035,N_8549);
and UO_860 (O_860,N_7646,N_7094);
nand UO_861 (O_861,N_8022,N_5435);
or UO_862 (O_862,N_7708,N_7124);
xor UO_863 (O_863,N_6662,N_6064);
or UO_864 (O_864,N_8194,N_5283);
and UO_865 (O_865,N_6612,N_8286);
nor UO_866 (O_866,N_7081,N_8029);
or UO_867 (O_867,N_7109,N_8341);
nand UO_868 (O_868,N_6139,N_6474);
xnor UO_869 (O_869,N_8831,N_6670);
xor UO_870 (O_870,N_9676,N_8141);
and UO_871 (O_871,N_5675,N_7830);
nor UO_872 (O_872,N_8294,N_8717);
nand UO_873 (O_873,N_6049,N_5700);
or UO_874 (O_874,N_8244,N_7775);
xnor UO_875 (O_875,N_6891,N_5332);
or UO_876 (O_876,N_8124,N_5797);
nand UO_877 (O_877,N_7641,N_6949);
or UO_878 (O_878,N_7385,N_8561);
xnor UO_879 (O_879,N_6978,N_8136);
and UO_880 (O_880,N_5012,N_7728);
xor UO_881 (O_881,N_8438,N_5412);
or UO_882 (O_882,N_9423,N_7307);
or UO_883 (O_883,N_6465,N_6969);
xor UO_884 (O_884,N_8268,N_5319);
xnor UO_885 (O_885,N_5265,N_6757);
or UO_886 (O_886,N_7761,N_6561);
and UO_887 (O_887,N_6309,N_8154);
nor UO_888 (O_888,N_5885,N_7571);
or UO_889 (O_889,N_7961,N_7482);
or UO_890 (O_890,N_8548,N_9048);
nand UO_891 (O_891,N_7188,N_9913);
nor UO_892 (O_892,N_6534,N_9799);
and UO_893 (O_893,N_5015,N_7038);
xor UO_894 (O_894,N_5827,N_9078);
and UO_895 (O_895,N_6711,N_8186);
and UO_896 (O_896,N_7564,N_8005);
nand UO_897 (O_897,N_8459,N_5408);
nand UO_898 (O_898,N_8922,N_6669);
nand UO_899 (O_899,N_7225,N_8913);
xnor UO_900 (O_900,N_9419,N_8572);
and UO_901 (O_901,N_9067,N_9231);
nor UO_902 (O_902,N_9771,N_9992);
nand UO_903 (O_903,N_7117,N_9523);
nor UO_904 (O_904,N_5448,N_8131);
nor UO_905 (O_905,N_5446,N_8987);
nand UO_906 (O_906,N_8881,N_6906);
nand UO_907 (O_907,N_8354,N_9714);
xnor UO_908 (O_908,N_5351,N_5972);
xor UO_909 (O_909,N_9986,N_7667);
nor UO_910 (O_910,N_6928,N_8162);
nand UO_911 (O_911,N_9094,N_6919);
nand UO_912 (O_912,N_6780,N_5795);
and UO_913 (O_913,N_7812,N_8407);
or UO_914 (O_914,N_9300,N_8429);
nor UO_915 (O_915,N_9274,N_6611);
xor UO_916 (O_916,N_8689,N_5630);
nand UO_917 (O_917,N_9165,N_6979);
nand UO_918 (O_918,N_6659,N_8100);
or UO_919 (O_919,N_6197,N_5604);
xnor UO_920 (O_920,N_8752,N_5387);
and UO_921 (O_921,N_8846,N_6610);
xor UO_922 (O_922,N_6070,N_8545);
xnor UO_923 (O_923,N_6723,N_9453);
and UO_924 (O_924,N_5938,N_5223);
nand UO_925 (O_925,N_9360,N_8299);
and UO_926 (O_926,N_6331,N_5846);
nor UO_927 (O_927,N_5296,N_6564);
nor UO_928 (O_928,N_5464,N_8781);
nand UO_929 (O_929,N_6020,N_8293);
nand UO_930 (O_930,N_7836,N_9199);
and UO_931 (O_931,N_5148,N_5588);
xnor UO_932 (O_932,N_6573,N_5274);
nor UO_933 (O_933,N_8526,N_7702);
or UO_934 (O_934,N_8559,N_6330);
or UO_935 (O_935,N_9206,N_7911);
xor UO_936 (O_936,N_5542,N_6665);
or UO_937 (O_937,N_6368,N_9931);
xnor UO_938 (O_938,N_9353,N_7522);
nor UO_939 (O_939,N_7252,N_6067);
xor UO_940 (O_940,N_5819,N_5643);
and UO_941 (O_941,N_7216,N_6421);
nor UO_942 (O_942,N_8874,N_5345);
and UO_943 (O_943,N_6395,N_9998);
or UO_944 (O_944,N_8651,N_6166);
and UO_945 (O_945,N_9477,N_5886);
nand UO_946 (O_946,N_5759,N_8398);
nand UO_947 (O_947,N_5466,N_9040);
and UO_948 (O_948,N_8096,N_6034);
and UO_949 (O_949,N_8821,N_7045);
nor UO_950 (O_950,N_5299,N_6037);
xor UO_951 (O_951,N_9677,N_9467);
or UO_952 (O_952,N_7536,N_6442);
nand UO_953 (O_953,N_5761,N_8822);
nor UO_954 (O_954,N_9359,N_5169);
nand UO_955 (O_955,N_9139,N_7772);
and UO_956 (O_956,N_7595,N_7864);
or UO_957 (O_957,N_6155,N_5556);
nor UO_958 (O_958,N_7319,N_5384);
xor UO_959 (O_959,N_7111,N_7645);
nor UO_960 (O_960,N_5056,N_7527);
and UO_961 (O_961,N_5072,N_6909);
xnor UO_962 (O_962,N_7876,N_5624);
or UO_963 (O_963,N_9322,N_5995);
or UO_964 (O_964,N_9307,N_5561);
xor UO_965 (O_965,N_8180,N_5181);
nand UO_966 (O_966,N_6543,N_7403);
and UO_967 (O_967,N_7986,N_6140);
xnor UO_968 (O_968,N_6119,N_9684);
xnor UO_969 (O_969,N_7861,N_7398);
and UO_970 (O_970,N_8033,N_8197);
or UO_971 (O_971,N_7827,N_5276);
or UO_972 (O_972,N_6112,N_9220);
or UO_973 (O_973,N_6858,N_8484);
nor UO_974 (O_974,N_7701,N_7871);
and UO_975 (O_975,N_5020,N_7365);
nand UO_976 (O_976,N_8837,N_7128);
or UO_977 (O_977,N_5225,N_6175);
nand UO_978 (O_978,N_5092,N_6013);
nor UO_979 (O_979,N_6598,N_8926);
or UO_980 (O_980,N_8747,N_9344);
xor UO_981 (O_981,N_5966,N_7041);
and UO_982 (O_982,N_5610,N_9180);
and UO_983 (O_983,N_9873,N_5897);
xnor UO_984 (O_984,N_9483,N_6342);
and UO_985 (O_985,N_6704,N_6654);
and UO_986 (O_986,N_7400,N_8684);
nand UO_987 (O_987,N_6916,N_5620);
nor UO_988 (O_988,N_8730,N_9624);
xor UO_989 (O_989,N_7163,N_9978);
nor UO_990 (O_990,N_9008,N_5058);
nor UO_991 (O_991,N_6677,N_9759);
and UO_992 (O_992,N_8613,N_6297);
xnor UO_993 (O_993,N_8798,N_7661);
xnor UO_994 (O_994,N_7688,N_6551);
nor UO_995 (O_995,N_8196,N_6762);
and UO_996 (O_996,N_7521,N_5417);
and UO_997 (O_997,N_9951,N_6233);
nor UO_998 (O_998,N_7235,N_9565);
xor UO_999 (O_999,N_5936,N_9033);
nor UO_1000 (O_1000,N_7233,N_8072);
xor UO_1001 (O_1001,N_9158,N_6187);
or UO_1002 (O_1002,N_7132,N_6167);
or UO_1003 (O_1003,N_5150,N_5873);
xnor UO_1004 (O_1004,N_8940,N_6621);
nand UO_1005 (O_1005,N_9544,N_8416);
nor UO_1006 (O_1006,N_7724,N_9366);
xor UO_1007 (O_1007,N_8884,N_8016);
and UO_1008 (O_1008,N_9868,N_8177);
nor UO_1009 (O_1009,N_5193,N_9876);
nand UO_1010 (O_1010,N_8793,N_8437);
nor UO_1011 (O_1011,N_8946,N_6603);
nor UO_1012 (O_1012,N_8207,N_7779);
and UO_1013 (O_1013,N_8217,N_8761);
or UO_1014 (O_1014,N_5709,N_8311);
xor UO_1015 (O_1015,N_6073,N_7700);
and UO_1016 (O_1016,N_8802,N_6738);
or UO_1017 (O_1017,N_8797,N_5974);
and UO_1018 (O_1018,N_9947,N_9770);
or UO_1019 (O_1019,N_5301,N_5582);
or UO_1020 (O_1020,N_6849,N_5923);
xor UO_1021 (O_1021,N_7611,N_6874);
nand UO_1022 (O_1022,N_5815,N_9358);
or UO_1023 (O_1023,N_9499,N_6560);
and UO_1024 (O_1024,N_8251,N_5590);
nor UO_1025 (O_1025,N_7253,N_6386);
nor UO_1026 (O_1026,N_7156,N_7067);
and UO_1027 (O_1027,N_5634,N_8562);
nand UO_1028 (O_1028,N_8259,N_8133);
nand UO_1029 (O_1029,N_9661,N_9543);
or UO_1030 (O_1030,N_6273,N_9492);
xor UO_1031 (O_1031,N_9392,N_9591);
nor UO_1032 (O_1032,N_9581,N_8357);
and UO_1033 (O_1033,N_6814,N_7313);
nor UO_1034 (O_1034,N_9704,N_6298);
or UO_1035 (O_1035,N_7805,N_6685);
and UO_1036 (O_1036,N_9559,N_9772);
or UO_1037 (O_1037,N_6970,N_9943);
and UO_1038 (O_1038,N_7605,N_6527);
nand UO_1039 (O_1039,N_8654,N_7555);
nand UO_1040 (O_1040,N_6688,N_7425);
xor UO_1041 (O_1041,N_8502,N_9196);
xnor UO_1042 (O_1042,N_8699,N_6444);
xnor UO_1043 (O_1043,N_8115,N_9766);
xor UO_1044 (O_1044,N_9553,N_6265);
or UO_1045 (O_1045,N_9526,N_8810);
xor UO_1046 (O_1046,N_7114,N_9134);
or UO_1047 (O_1047,N_8172,N_7320);
xor UO_1048 (O_1048,N_8258,N_6452);
xor UO_1049 (O_1049,N_8596,N_7243);
nand UO_1050 (O_1050,N_5682,N_5830);
or UO_1051 (O_1051,N_8090,N_7575);
nand UO_1052 (O_1052,N_5532,N_6760);
nor UO_1053 (O_1053,N_5271,N_7972);
nand UO_1054 (O_1054,N_8595,N_6156);
xnor UO_1055 (O_1055,N_7915,N_8030);
or UO_1056 (O_1056,N_7452,N_7561);
nor UO_1057 (O_1057,N_8701,N_9495);
and UO_1058 (O_1058,N_5108,N_6356);
nor UO_1059 (O_1059,N_8634,N_6951);
or UO_1060 (O_1060,N_5667,N_7719);
and UO_1061 (O_1061,N_7668,N_7091);
or UO_1062 (O_1062,N_9768,N_6638);
and UO_1063 (O_1063,N_6278,N_6134);
or UO_1064 (O_1064,N_7358,N_9280);
and UO_1065 (O_1065,N_8953,N_9690);
nand UO_1066 (O_1066,N_8656,N_5231);
xor UO_1067 (O_1067,N_5130,N_5553);
or UO_1068 (O_1068,N_9911,N_8639);
nor UO_1069 (O_1069,N_8402,N_9717);
xor UO_1070 (O_1070,N_7259,N_7863);
nand UO_1071 (O_1071,N_9001,N_9850);
nand UO_1072 (O_1072,N_7742,N_8765);
and UO_1073 (O_1073,N_7982,N_9635);
and UO_1074 (O_1074,N_9020,N_5767);
or UO_1075 (O_1075,N_7110,N_6907);
nor UO_1076 (O_1076,N_9735,N_5442);
nand UO_1077 (O_1077,N_8672,N_5565);
xor UO_1078 (O_1078,N_8750,N_5114);
nand UO_1079 (O_1079,N_8210,N_5594);
or UO_1080 (O_1080,N_8372,N_7466);
or UO_1081 (O_1081,N_7342,N_6675);
and UO_1082 (O_1082,N_7290,N_5747);
or UO_1083 (O_1083,N_8980,N_9475);
nand UO_1084 (O_1084,N_9329,N_8617);
and UO_1085 (O_1085,N_7811,N_6851);
and UO_1086 (O_1086,N_9119,N_5696);
and UO_1087 (O_1087,N_7429,N_6802);
nor UO_1088 (O_1088,N_9547,N_6186);
or UO_1089 (O_1089,N_8344,N_5746);
nand UO_1090 (O_1090,N_5142,N_8331);
and UO_1091 (O_1091,N_7921,N_7386);
nor UO_1092 (O_1092,N_9734,N_8960);
or UO_1093 (O_1093,N_9846,N_6913);
and UO_1094 (O_1094,N_7150,N_6812);
and UO_1095 (O_1095,N_9686,N_9572);
nor UO_1096 (O_1096,N_7543,N_5845);
or UO_1097 (O_1097,N_9566,N_9822);
and UO_1098 (O_1098,N_6808,N_6968);
and UO_1099 (O_1099,N_7581,N_7424);
or UO_1100 (O_1100,N_8049,N_5034);
nor UO_1101 (O_1101,N_8585,N_6735);
xor UO_1102 (O_1102,N_7707,N_5290);
xnor UO_1103 (O_1103,N_5981,N_9273);
nand UO_1104 (O_1104,N_6477,N_8184);
xnor UO_1105 (O_1105,N_7879,N_5418);
or UO_1106 (O_1106,N_7973,N_9021);
nor UO_1107 (O_1107,N_9891,N_9238);
nor UO_1108 (O_1108,N_6615,N_6592);
or UO_1109 (O_1109,N_9653,N_6695);
or UO_1110 (O_1110,N_8155,N_5512);
or UO_1111 (O_1111,N_7269,N_6748);
or UO_1112 (O_1112,N_6321,N_7547);
xor UO_1113 (O_1113,N_6664,N_6954);
nor UO_1114 (O_1114,N_9675,N_5940);
xor UO_1115 (O_1115,N_9834,N_6996);
nor UO_1116 (O_1116,N_6377,N_7549);
nand UO_1117 (O_1117,N_7865,N_5666);
xnor UO_1118 (O_1118,N_5258,N_7803);
nor UO_1119 (O_1119,N_5883,N_6225);
xor UO_1120 (O_1120,N_8935,N_7501);
nor UO_1121 (O_1121,N_5976,N_9068);
xnor UO_1122 (O_1122,N_6409,N_5485);
xnor UO_1123 (O_1123,N_8390,N_7426);
xnor UO_1124 (O_1124,N_7113,N_8025);
nor UO_1125 (O_1125,N_8996,N_5898);
and UO_1126 (O_1126,N_9346,N_9116);
and UO_1127 (O_1127,N_6286,N_7145);
nand UO_1128 (O_1128,N_8279,N_9311);
and UO_1129 (O_1129,N_5084,N_9844);
xor UO_1130 (O_1130,N_8393,N_9294);
and UO_1131 (O_1131,N_6642,N_5618);
nor UO_1132 (O_1132,N_9536,N_7105);
xor UO_1133 (O_1133,N_9728,N_9959);
or UO_1134 (O_1134,N_5713,N_6847);
nor UO_1135 (O_1135,N_7990,N_9493);
nor UO_1136 (O_1136,N_5612,N_8748);
and UO_1137 (O_1137,N_8988,N_6249);
nor UO_1138 (O_1138,N_9200,N_9357);
nor UO_1139 (O_1139,N_8904,N_7084);
nand UO_1140 (O_1140,N_7838,N_7254);
xnor UO_1141 (O_1141,N_5982,N_7095);
and UO_1142 (O_1142,N_5905,N_9383);
or UO_1143 (O_1143,N_6562,N_5219);
nor UO_1144 (O_1144,N_8963,N_7229);
and UO_1145 (O_1145,N_7449,N_7790);
or UO_1146 (O_1146,N_9557,N_7333);
and UO_1147 (O_1147,N_5144,N_8724);
xor UO_1148 (O_1148,N_9405,N_6838);
and UO_1149 (O_1149,N_6989,N_9528);
nand UO_1150 (O_1150,N_6420,N_9721);
nand UO_1151 (O_1151,N_5257,N_5921);
nand UO_1152 (O_1152,N_9671,N_6545);
nor UO_1153 (O_1153,N_5680,N_7363);
or UO_1154 (O_1154,N_5119,N_5308);
nor UO_1155 (O_1155,N_6727,N_5490);
xnor UO_1156 (O_1156,N_6306,N_9208);
xor UO_1157 (O_1157,N_9141,N_9880);
and UO_1158 (O_1158,N_9016,N_9326);
nor UO_1159 (O_1159,N_6823,N_9705);
nand UO_1160 (O_1160,N_9716,N_5692);
xnor UO_1161 (O_1161,N_6349,N_9491);
nand UO_1162 (O_1162,N_7048,N_7783);
or UO_1163 (O_1163,N_9101,N_6593);
nor UO_1164 (O_1164,N_5383,N_5716);
xor UO_1165 (O_1165,N_7592,N_8064);
nor UO_1166 (O_1166,N_6117,N_6215);
and UO_1167 (O_1167,N_6625,N_5057);
xor UO_1168 (O_1168,N_5902,N_6359);
nand UO_1169 (O_1169,N_5048,N_6568);
nor UO_1170 (O_1170,N_8519,N_5856);
xor UO_1171 (O_1171,N_7498,N_9809);
and UO_1172 (O_1172,N_9412,N_5011);
and UO_1173 (O_1173,N_5459,N_6471);
nand UO_1174 (O_1174,N_8855,N_6956);
or UO_1175 (O_1175,N_6009,N_7837);
nand UO_1176 (O_1176,N_5232,N_8537);
or UO_1177 (O_1177,N_5672,N_9592);
nand UO_1178 (O_1178,N_8758,N_7433);
and UO_1179 (O_1179,N_5571,N_8383);
nor UO_1180 (O_1180,N_7187,N_6959);
nor UO_1181 (O_1181,N_5699,N_8062);
and UO_1182 (O_1182,N_6093,N_7759);
nand UO_1183 (O_1183,N_7380,N_8709);
nor UO_1184 (O_1184,N_5941,N_8993);
nor UO_1185 (O_1185,N_7718,N_9096);
nand UO_1186 (O_1186,N_8465,N_5489);
or UO_1187 (O_1187,N_5799,N_7099);
nand UO_1188 (O_1188,N_9590,N_7352);
nand UO_1189 (O_1189,N_7925,N_9066);
nor UO_1190 (O_1190,N_6594,N_6424);
nor UO_1191 (O_1191,N_8307,N_9507);
nand UO_1192 (O_1192,N_5658,N_5203);
xor UO_1193 (O_1193,N_9393,N_5931);
nand UO_1194 (O_1194,N_6721,N_5708);
or UO_1195 (O_1195,N_8807,N_6582);
xor UO_1196 (O_1196,N_5805,N_5792);
nor UO_1197 (O_1197,N_9933,N_5581);
and UO_1198 (O_1198,N_8872,N_7942);
nand UO_1199 (O_1199,N_6833,N_7218);
xnor UO_1200 (O_1200,N_6745,N_6862);
nor UO_1201 (O_1201,N_6775,N_5963);
nor UO_1202 (O_1202,N_8445,N_8493);
nand UO_1203 (O_1203,N_6764,N_9203);
nand UO_1204 (O_1204,N_6043,N_9434);
and UO_1205 (O_1205,N_7769,N_8658);
or UO_1206 (O_1206,N_8894,N_9888);
or UO_1207 (O_1207,N_8257,N_6081);
or UO_1208 (O_1208,N_5341,N_9457);
and UO_1209 (O_1209,N_7600,N_9128);
and UO_1210 (O_1210,N_6351,N_5813);
nand UO_1211 (O_1211,N_6502,N_5631);
xor UO_1212 (O_1212,N_7237,N_7541);
nor UO_1213 (O_1213,N_6461,N_5660);
nand UO_1214 (O_1214,N_8623,N_6456);
xnor UO_1215 (O_1215,N_9437,N_7219);
nand UO_1216 (O_1216,N_8815,N_6601);
or UO_1217 (O_1217,N_9100,N_9829);
and UO_1218 (O_1218,N_6428,N_8007);
xor UO_1219 (O_1219,N_7846,N_7962);
and UO_1220 (O_1220,N_9619,N_9289);
nor UO_1221 (O_1221,N_8220,N_9132);
nand UO_1222 (O_1222,N_7464,N_7042);
xor UO_1223 (O_1223,N_7883,N_9606);
or UO_1224 (O_1224,N_5436,N_9036);
and UO_1225 (O_1225,N_8394,N_7037);
or UO_1226 (O_1226,N_7164,N_7223);
and UO_1227 (O_1227,N_6316,N_6712);
xor UO_1228 (O_1228,N_5067,N_5104);
nand UO_1229 (O_1229,N_5563,N_8785);
and UO_1230 (O_1230,N_5939,N_8409);
nor UO_1231 (O_1231,N_9551,N_8447);
nor UO_1232 (O_1232,N_8442,N_9298);
xnor UO_1233 (O_1233,N_8604,N_5406);
xnor UO_1234 (O_1234,N_7610,N_6239);
xor UO_1235 (O_1235,N_8499,N_7983);
xor UO_1236 (O_1236,N_5409,N_8731);
nand UO_1237 (O_1237,N_9053,N_5458);
nand UO_1238 (O_1238,N_6417,N_9539);
and UO_1239 (O_1239,N_8829,N_5870);
nand UO_1240 (O_1240,N_6168,N_6587);
xnor UO_1241 (O_1241,N_7440,N_6947);
nor UO_1242 (O_1242,N_6027,N_8843);
xnor UO_1243 (O_1243,N_9878,N_9038);
nor UO_1244 (O_1244,N_7905,N_8009);
or UO_1245 (O_1245,N_8966,N_6416);
or UO_1246 (O_1246,N_5986,N_5160);
nor UO_1247 (O_1247,N_8310,N_6328);
or UO_1248 (O_1248,N_9049,N_6522);
or UO_1249 (O_1249,N_6104,N_5235);
xnor UO_1250 (O_1250,N_7294,N_7926);
xnor UO_1251 (O_1251,N_6352,N_9151);
xor UO_1252 (O_1252,N_9218,N_8961);
nand UO_1253 (O_1253,N_8728,N_8877);
and UO_1254 (O_1254,N_5105,N_5851);
xnor UO_1255 (O_1255,N_7063,N_8224);
and UO_1256 (O_1256,N_9823,N_9129);
xor UO_1257 (O_1257,N_7949,N_8777);
xnor UO_1258 (O_1258,N_9832,N_7738);
and UO_1259 (O_1259,N_7802,N_7118);
nor UO_1260 (O_1260,N_9589,N_5530);
xor UO_1261 (O_1261,N_7211,N_8384);
or UO_1262 (O_1262,N_8219,N_8967);
nor UO_1263 (O_1263,N_5833,N_8530);
nand UO_1264 (O_1264,N_6430,N_6447);
nor UO_1265 (O_1265,N_8335,N_5139);
nor UO_1266 (O_1266,N_9173,N_5414);
or UO_1267 (O_1267,N_6876,N_9379);
xnor UO_1268 (O_1268,N_8563,N_7361);
and UO_1269 (O_1269,N_8581,N_9637);
xnor UO_1270 (O_1270,N_9142,N_9321);
nor UO_1271 (O_1271,N_7933,N_6212);
or UO_1272 (O_1272,N_6218,N_6618);
and UO_1273 (O_1273,N_5595,N_9286);
xnor UO_1274 (O_1274,N_6124,N_5208);
nand UO_1275 (O_1275,N_5926,N_8875);
and UO_1276 (O_1276,N_7408,N_7873);
xor UO_1277 (O_1277,N_5152,N_5468);
xor UO_1278 (O_1278,N_7298,N_5330);
or UO_1279 (O_1279,N_9524,N_5924);
xor UO_1280 (O_1280,N_5511,N_7412);
xor UO_1281 (O_1281,N_8053,N_9962);
nand UO_1282 (O_1282,N_5248,N_7928);
or UO_1283 (O_1283,N_7096,N_7927);
and UO_1284 (O_1284,N_9726,N_8702);
xor UO_1285 (O_1285,N_8983,N_7028);
xnor UO_1286 (O_1286,N_9582,N_5637);
nor UO_1287 (O_1287,N_5959,N_8552);
or UO_1288 (O_1288,N_7922,N_5887);
or UO_1289 (O_1289,N_9660,N_5328);
and UO_1290 (O_1290,N_6026,N_7654);
nand UO_1291 (O_1291,N_5834,N_8024);
nand UO_1292 (O_1292,N_7210,N_6035);
nand UO_1293 (O_1293,N_7173,N_8587);
nor UO_1294 (O_1294,N_7271,N_8103);
nand UO_1295 (O_1295,N_8692,N_6098);
or UO_1296 (O_1296,N_8486,N_6640);
nor UO_1297 (O_1297,N_9443,N_7599);
nor UO_1298 (O_1298,N_7886,N_6648);
nand UO_1299 (O_1299,N_9421,N_9884);
nand UO_1300 (O_1300,N_8789,N_9937);
nor UO_1301 (O_1301,N_9853,N_6032);
nor UO_1302 (O_1302,N_6276,N_8624);
xor UO_1303 (O_1303,N_5260,N_8813);
nand UO_1304 (O_1304,N_9169,N_9700);
xor UO_1305 (O_1305,N_8500,N_8065);
nor UO_1306 (O_1306,N_6614,N_9445);
and UO_1307 (O_1307,N_7343,N_5576);
nand UO_1308 (O_1308,N_6469,N_6813);
xnor UO_1309 (O_1309,N_9779,N_8476);
xnor UO_1310 (O_1310,N_6406,N_6029);
nor UO_1311 (O_1311,N_5083,N_6827);
xnor UO_1312 (O_1312,N_6914,N_8478);
and UO_1313 (O_1313,N_5204,N_5070);
xnor UO_1314 (O_1314,N_5041,N_5434);
nand UO_1315 (O_1315,N_5107,N_8485);
and UO_1316 (O_1316,N_7071,N_7796);
nor UO_1317 (O_1317,N_9210,N_6317);
nor UO_1318 (O_1318,N_5726,N_9510);
nand UO_1319 (O_1319,N_8015,N_6500);
nor UO_1320 (O_1320,N_6177,N_7069);
nand UO_1321 (O_1321,N_8594,N_7415);
and UO_1322 (O_1322,N_9205,N_6892);
or UO_1323 (O_1323,N_6497,N_8075);
and UO_1324 (O_1324,N_5794,N_6679);
or UO_1325 (O_1325,N_6147,N_9755);
xor UO_1326 (O_1326,N_9451,N_7715);
or UO_1327 (O_1327,N_7548,N_6976);
and UO_1328 (O_1328,N_8929,N_5528);
and UO_1329 (O_1329,N_6682,N_7165);
and UO_1330 (O_1330,N_5629,N_9074);
and UO_1331 (O_1331,N_5645,N_5238);
and UO_1332 (O_1332,N_5044,N_8842);
xor UO_1333 (O_1333,N_5001,N_6132);
and UO_1334 (O_1334,N_8944,N_7289);
and UO_1335 (O_1335,N_8600,N_9961);
and UO_1336 (O_1336,N_5961,N_8423);
and UO_1337 (O_1337,N_9002,N_7183);
xnor UO_1338 (O_1338,N_6797,N_8833);
xnor UO_1339 (O_1339,N_7453,N_5128);
xnor UO_1340 (O_1340,N_9817,N_8266);
nand UO_1341 (O_1341,N_7406,N_7618);
nor UO_1342 (O_1342,N_7085,N_6690);
xnor UO_1343 (O_1343,N_7874,N_8108);
nor UO_1344 (O_1344,N_8260,N_6693);
nand UO_1345 (O_1345,N_9190,N_5213);
and UO_1346 (O_1346,N_7153,N_8298);
and UO_1347 (O_1347,N_7870,N_8321);
nor UO_1348 (O_1348,N_9948,N_7776);
and UO_1349 (O_1349,N_7007,N_7127);
nand UO_1350 (O_1350,N_7898,N_7506);
xnor UO_1351 (O_1351,N_9813,N_5331);
and UO_1352 (O_1352,N_8175,N_7083);
and UO_1353 (O_1353,N_7323,N_9668);
nor UO_1354 (O_1354,N_9448,N_5137);
or UO_1355 (O_1355,N_7782,N_7729);
xnor UO_1356 (O_1356,N_7852,N_7311);
or UO_1357 (O_1357,N_8925,N_6425);
xnor UO_1358 (O_1358,N_8799,N_9746);
nand UO_1359 (O_1359,N_5835,N_9195);
nor UO_1360 (O_1360,N_7674,N_9652);
xor UO_1361 (O_1361,N_8487,N_7686);
xor UO_1362 (O_1362,N_7848,N_8975);
and UO_1363 (O_1363,N_8336,N_7322);
or UO_1364 (O_1364,N_5720,N_8696);
or UO_1365 (O_1365,N_7025,N_7885);
xnor UO_1366 (O_1366,N_9877,N_8300);
nor UO_1367 (O_1367,N_8123,N_5253);
nand UO_1368 (O_1368,N_8076,N_9474);
nand UO_1369 (O_1369,N_5570,N_7649);
and UO_1370 (O_1370,N_6843,N_7418);
nor UO_1371 (O_1371,N_5439,N_6382);
and UO_1372 (O_1372,N_6003,N_9963);
nand UO_1373 (O_1373,N_8011,N_8408);
xor UO_1374 (O_1374,N_6054,N_5502);
nor UO_1375 (O_1375,N_8543,N_9345);
xnor UO_1376 (O_1376,N_6773,N_6436);
xnor UO_1377 (O_1377,N_5690,N_8169);
nand UO_1378 (O_1378,N_8914,N_5646);
xor UO_1379 (O_1379,N_7070,N_6557);
or UO_1380 (O_1380,N_5722,N_7919);
xnor UO_1381 (O_1381,N_8919,N_5586);
nor UO_1382 (O_1382,N_6774,N_5147);
xnor UO_1383 (O_1383,N_5426,N_6830);
nand UO_1384 (O_1384,N_9256,N_5481);
or UO_1385 (O_1385,N_9102,N_6312);
or UO_1386 (O_1386,N_6929,N_7228);
xor UO_1387 (O_1387,N_9981,N_5180);
or UO_1388 (O_1388,N_5315,N_5457);
or UO_1389 (O_1389,N_8576,N_5197);
or UO_1390 (O_1390,N_6121,N_8028);
or UO_1391 (O_1391,N_8659,N_5664);
nor UO_1392 (O_1392,N_5679,N_9805);
nor UO_1393 (O_1393,N_8912,N_8051);
nand UO_1394 (O_1394,N_5977,N_7303);
nor UO_1395 (O_1395,N_8533,N_5440);
or UO_1396 (O_1396,N_6264,N_5307);
and UO_1397 (O_1397,N_8737,N_6414);
nor UO_1398 (O_1398,N_6254,N_7748);
or UO_1399 (O_1399,N_5533,N_9692);
and UO_1400 (O_1400,N_7751,N_6302);
or UO_1401 (O_1401,N_7354,N_6341);
xnor UO_1402 (O_1402,N_8869,N_6622);
and UO_1403 (O_1403,N_9255,N_7801);
nor UO_1404 (O_1404,N_9605,N_6295);
nand UO_1405 (O_1405,N_6917,N_9821);
and UO_1406 (O_1406,N_7061,N_9110);
or UO_1407 (O_1407,N_5775,N_8591);
nand UO_1408 (O_1408,N_9837,N_8334);
xor UO_1409 (O_1409,N_8824,N_6252);
nor UO_1410 (O_1410,N_8479,N_9549);
nand UO_1411 (O_1411,N_5748,N_9534);
or UO_1412 (O_1412,N_5006,N_7720);
and UO_1413 (O_1413,N_8762,N_6160);
or UO_1414 (O_1414,N_9373,N_8130);
nor UO_1415 (O_1415,N_9835,N_9901);
or UO_1416 (O_1416,N_7032,N_9403);
nand UO_1417 (O_1417,N_6285,N_8339);
nand UO_1418 (O_1418,N_8379,N_8749);
nand UO_1419 (O_1419,N_5247,N_6464);
nor UO_1420 (O_1420,N_5822,N_7583);
xnor UO_1421 (O_1421,N_7341,N_7486);
or UO_1422 (O_1422,N_5606,N_8122);
and UO_1423 (O_1423,N_6450,N_7814);
xnor UO_1424 (O_1424,N_9952,N_6809);
or UO_1425 (O_1425,N_5881,N_5077);
nand UO_1426 (O_1426,N_7004,N_9188);
nor UO_1427 (O_1427,N_5781,N_5554);
and UO_1428 (O_1428,N_5127,N_9567);
or UO_1429 (O_1429,N_9666,N_7872);
or UO_1430 (O_1430,N_5305,N_9945);
and UO_1431 (O_1431,N_9797,N_7831);
or UO_1432 (O_1432,N_7267,N_6556);
or UO_1433 (O_1433,N_9336,N_9438);
nor UO_1434 (O_1434,N_7978,N_8192);
or UO_1435 (O_1435,N_5339,N_8397);
and UO_1436 (O_1436,N_6600,N_8018);
and UO_1437 (O_1437,N_6426,N_5093);
nor UO_1438 (O_1438,N_6936,N_5651);
nand UO_1439 (O_1439,N_6900,N_9576);
nand UO_1440 (O_1440,N_5261,N_7895);
xnor UO_1441 (O_1441,N_7420,N_9550);
or UO_1442 (O_1442,N_8907,N_5052);
or UO_1443 (O_1443,N_6205,N_8288);
nand UO_1444 (O_1444,N_9301,N_7065);
nand UO_1445 (O_1445,N_6718,N_9979);
and UO_1446 (O_1446,N_8721,N_8374);
nand UO_1447 (O_1447,N_8014,N_7625);
or UO_1448 (O_1448,N_6961,N_6488);
and UO_1449 (O_1449,N_7637,N_8540);
xnor UO_1450 (O_1450,N_5303,N_6684);
nand UO_1451 (O_1451,N_8056,N_5729);
and UO_1452 (O_1452,N_7881,N_9178);
and UO_1453 (O_1453,N_9958,N_6041);
nand UO_1454 (O_1454,N_5221,N_7273);
nor UO_1455 (O_1455,N_6716,N_8222);
nor UO_1456 (O_1456,N_5810,N_6169);
nor UO_1457 (O_1457,N_5600,N_6453);
or UO_1458 (O_1458,N_5194,N_6059);
xor UO_1459 (O_1459,N_9623,N_9378);
nand UO_1460 (O_1460,N_5392,N_7507);
and UO_1461 (O_1461,N_6524,N_7628);
and UO_1462 (O_1462,N_6247,N_6262);
or UO_1463 (O_1463,N_6974,N_8161);
xnor UO_1464 (O_1464,N_8365,N_7539);
nand UO_1465 (O_1465,N_9935,N_6576);
or UO_1466 (O_1466,N_6318,N_8817);
and UO_1467 (O_1467,N_9328,N_5895);
nor UO_1468 (O_1468,N_6580,N_8514);
nor UO_1469 (O_1469,N_8796,N_9857);
nor UO_1470 (O_1470,N_7141,N_9996);
nand UO_1471 (O_1471,N_8628,N_7469);
xnor UO_1472 (O_1472,N_8189,N_8249);
nor UO_1473 (O_1473,N_7146,N_9441);
and UO_1474 (O_1474,N_8566,N_8403);
nand UO_1475 (O_1475,N_7136,N_5171);
nand UO_1476 (O_1476,N_7560,N_9645);
nor UO_1477 (O_1477,N_7089,N_8427);
nor UO_1478 (O_1478,N_9753,N_6962);
nand UO_1479 (O_1479,N_5029,N_9924);
or UO_1480 (O_1480,N_5840,N_9091);
xnor UO_1481 (O_1481,N_6388,N_6759);
or UO_1482 (O_1482,N_7636,N_7138);
or UO_1483 (O_1483,N_7970,N_6528);
nand UO_1484 (O_1484,N_9297,N_8995);
nor UO_1485 (O_1485,N_7119,N_8578);
nand UO_1486 (O_1486,N_9364,N_9504);
and UO_1487 (O_1487,N_5143,N_9088);
xor UO_1488 (O_1488,N_6920,N_7052);
xnor UO_1489 (O_1489,N_7713,N_8138);
nor UO_1490 (O_1490,N_6145,N_7496);
nand UO_1491 (O_1491,N_8285,N_9919);
and UO_1492 (O_1492,N_8898,N_5050);
or UO_1493 (O_1493,N_9587,N_6810);
and UO_1494 (O_1494,N_7460,N_9281);
nand UO_1495 (O_1495,N_6747,N_7655);
or UO_1496 (O_1496,N_5566,N_6348);
xor UO_1497 (O_1497,N_8652,N_9938);
xor UO_1498 (O_1498,N_6209,N_8574);
or UO_1499 (O_1499,N_5124,N_7053);
endmodule