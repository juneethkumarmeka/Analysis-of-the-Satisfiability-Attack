module basic_2000_20000_2500_40_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_1949,In_1547);
and U1 (N_1,In_456,In_436);
or U2 (N_2,In_550,In_1584);
nand U3 (N_3,In_236,In_527);
or U4 (N_4,In_1112,In_156);
or U5 (N_5,In_1895,In_900);
nand U6 (N_6,In_351,In_779);
and U7 (N_7,In_1155,In_1992);
xnor U8 (N_8,In_1807,In_1859);
nor U9 (N_9,In_1700,In_478);
nor U10 (N_10,In_796,In_266);
xor U11 (N_11,In_1211,In_503);
or U12 (N_12,In_404,In_1068);
xor U13 (N_13,In_98,In_954);
and U14 (N_14,In_539,In_188);
xnor U15 (N_15,In_1989,In_1986);
nand U16 (N_16,In_402,In_1438);
nor U17 (N_17,In_845,In_1014);
nand U18 (N_18,In_441,In_386);
nor U19 (N_19,In_907,In_234);
nor U20 (N_20,In_6,In_488);
nor U21 (N_21,In_1149,In_659);
nand U22 (N_22,In_1387,In_480);
and U23 (N_23,In_35,In_1133);
nand U24 (N_24,In_809,In_1210);
nor U25 (N_25,In_18,In_1001);
or U26 (N_26,In_803,In_1143);
nor U27 (N_27,In_226,In_312);
xnor U28 (N_28,In_901,In_93);
and U29 (N_29,In_1128,In_1307);
and U30 (N_30,In_1216,In_590);
and U31 (N_31,In_1994,In_1504);
or U32 (N_32,In_1317,In_356);
nand U33 (N_33,In_1689,In_915);
nand U34 (N_34,In_768,In_1559);
and U35 (N_35,In_71,In_1714);
xnor U36 (N_36,In_338,In_1728);
or U37 (N_37,In_1623,In_426);
nor U38 (N_38,In_667,In_1668);
nor U39 (N_39,In_105,In_693);
nor U40 (N_40,In_1159,In_1640);
nand U41 (N_41,In_567,In_135);
or U42 (N_42,In_538,In_1738);
xnor U43 (N_43,In_339,In_1785);
and U44 (N_44,In_1719,In_1087);
nor U45 (N_45,In_101,In_1196);
and U46 (N_46,In_1748,In_96);
or U47 (N_47,In_1290,In_52);
and U48 (N_48,In_573,In_1398);
or U49 (N_49,In_1433,In_640);
nor U50 (N_50,In_1270,In_1255);
nor U51 (N_51,In_1548,In_620);
or U52 (N_52,In_649,In_846);
and U53 (N_53,In_1957,In_701);
nor U54 (N_54,In_955,In_1578);
and U55 (N_55,In_995,In_116);
nor U56 (N_56,In_1043,In_760);
nand U57 (N_57,In_267,In_741);
nand U58 (N_58,In_139,In_1184);
or U59 (N_59,In_1840,In_1792);
nand U60 (N_60,In_1884,In_1570);
nor U61 (N_61,In_1301,In_1075);
and U62 (N_62,In_1261,In_165);
or U63 (N_63,In_1786,In_1090);
nor U64 (N_64,In_160,In_1636);
nor U65 (N_65,In_1976,In_1931);
or U66 (N_66,In_137,In_576);
or U67 (N_67,In_1698,In_1421);
or U68 (N_68,In_318,In_124);
xnor U69 (N_69,In_1222,In_189);
and U70 (N_70,In_601,In_844);
xor U71 (N_71,In_1380,In_401);
xnor U72 (N_72,In_1338,In_932);
nand U73 (N_73,In_1500,In_1172);
xor U74 (N_74,In_1049,In_560);
and U75 (N_75,In_1970,In_1188);
nand U76 (N_76,In_1522,In_286);
xnor U77 (N_77,In_1120,In_1424);
nor U78 (N_78,In_350,In_1289);
nand U79 (N_79,In_973,In_618);
xor U80 (N_80,In_63,In_792);
nand U81 (N_81,In_1315,In_1551);
nand U82 (N_82,In_1019,In_512);
xor U83 (N_83,In_1590,In_1140);
or U84 (N_84,In_1612,In_1896);
nor U85 (N_85,In_990,In_1803);
and U86 (N_86,In_542,In_981);
and U87 (N_87,In_662,In_199);
and U88 (N_88,In_1798,In_883);
and U89 (N_89,In_1830,In_1973);
and U90 (N_90,In_737,In_1069);
nand U91 (N_91,In_1660,In_1088);
nand U92 (N_92,In_1635,In_818);
nand U93 (N_93,In_825,In_893);
or U94 (N_94,In_1793,In_1524);
nand U95 (N_95,In_974,In_664);
nor U96 (N_96,In_656,In_802);
or U97 (N_97,In_1875,In_157);
xnor U98 (N_98,In_507,In_738);
nor U99 (N_99,In_1560,In_1499);
or U100 (N_100,In_562,In_604);
and U101 (N_101,In_1634,In_9);
nor U102 (N_102,In_834,In_1580);
xnor U103 (N_103,In_1384,In_869);
nand U104 (N_104,In_819,In_1263);
xor U105 (N_105,In_1930,In_43);
xor U106 (N_106,In_1705,In_721);
nand U107 (N_107,In_914,In_1228);
nand U108 (N_108,In_798,In_1562);
nor U109 (N_109,In_1519,In_1103);
or U110 (N_110,In_1028,In_36);
and U111 (N_111,In_1162,In_1180);
or U112 (N_112,In_1906,In_905);
xor U113 (N_113,In_1052,In_24);
xnor U114 (N_114,In_1557,In_887);
nand U115 (N_115,In_222,In_730);
xor U116 (N_116,In_966,In_1111);
nor U117 (N_117,In_1246,In_1170);
and U118 (N_118,In_1709,In_1688);
and U119 (N_119,In_1611,In_1343);
and U120 (N_120,In_1477,In_1395);
or U121 (N_121,In_686,In_638);
and U122 (N_122,In_599,In_1536);
and U123 (N_123,In_427,In_1409);
nand U124 (N_124,In_1825,In_377);
or U125 (N_125,In_1359,In_1000);
or U126 (N_126,In_1865,In_598);
or U127 (N_127,In_549,In_671);
and U128 (N_128,In_1532,In_676);
and U129 (N_129,In_1476,In_370);
nor U130 (N_130,In_1783,In_578);
nand U131 (N_131,In_559,In_1329);
or U132 (N_132,In_502,In_722);
nand U133 (N_133,In_215,In_922);
and U134 (N_134,In_1824,In_147);
nor U135 (N_135,In_150,In_384);
nor U136 (N_136,In_1201,In_1432);
or U137 (N_137,In_1072,In_976);
or U138 (N_138,In_1776,In_1165);
xnor U139 (N_139,In_675,In_1911);
nand U140 (N_140,In_1481,In_1682);
or U141 (N_141,In_704,In_496);
nor U142 (N_142,In_1595,In_1749);
nand U143 (N_143,In_1773,In_1979);
or U144 (N_144,In_1953,In_1061);
nor U145 (N_145,In_1036,In_1721);
nand U146 (N_146,In_252,In_1491);
nand U147 (N_147,In_1483,In_820);
nand U148 (N_148,In_308,In_710);
nand U149 (N_149,In_574,In_581);
nand U150 (N_150,In_57,In_1065);
or U151 (N_151,In_1236,In_655);
nand U152 (N_152,In_1761,In_183);
nor U153 (N_153,In_1313,In_1566);
nor U154 (N_154,In_1126,In_1005);
or U155 (N_155,In_1730,In_164);
nor U156 (N_156,In_315,In_484);
and U157 (N_157,In_1206,In_1944);
xnor U158 (N_158,In_1663,In_1404);
nand U159 (N_159,In_870,In_906);
xor U160 (N_160,In_1053,In_1495);
nor U161 (N_161,In_968,In_528);
nor U162 (N_162,In_608,In_1017);
nor U163 (N_163,In_536,In_635);
nand U164 (N_164,In_1959,In_1443);
and U165 (N_165,In_1391,In_1084);
nor U166 (N_166,In_469,In_1877);
and U167 (N_167,In_621,In_211);
nor U168 (N_168,In_669,In_394);
xnor U169 (N_169,In_761,In_442);
nand U170 (N_170,In_780,In_218);
nand U171 (N_171,In_1051,In_866);
and U172 (N_172,In_191,In_513);
nand U173 (N_173,In_1981,In_904);
or U174 (N_174,In_1975,In_1034);
nand U175 (N_175,In_145,In_1412);
or U176 (N_176,In_849,In_1811);
xnor U177 (N_177,In_1939,In_87);
xor U178 (N_178,In_534,In_46);
xnor U179 (N_179,In_735,In_1235);
nand U180 (N_180,In_1240,In_933);
nor U181 (N_181,In_657,In_1956);
and U182 (N_182,In_313,In_133);
nor U183 (N_183,In_1279,In_1815);
xor U184 (N_184,In_886,In_716);
nor U185 (N_185,In_207,In_94);
nand U186 (N_186,In_1687,In_747);
and U187 (N_187,In_1330,In_1407);
xor U188 (N_188,In_73,In_852);
nor U189 (N_189,In_674,In_962);
xnor U190 (N_190,In_518,In_917);
nor U191 (N_191,In_944,In_924);
nand U192 (N_192,In_986,In_50);
xnor U193 (N_193,In_872,In_609);
nand U194 (N_194,In_1488,In_847);
nand U195 (N_195,In_1630,In_1493);
and U196 (N_196,In_531,In_1645);
nor U197 (N_197,In_764,In_162);
or U198 (N_198,In_1633,In_719);
nand U199 (N_199,In_0,In_541);
and U200 (N_200,In_882,In_1517);
or U201 (N_201,In_324,In_1269);
xnor U202 (N_202,In_1958,In_1987);
xor U203 (N_203,In_1675,In_1239);
nand U204 (N_204,In_45,In_364);
nand U205 (N_205,In_134,In_1616);
nand U206 (N_206,In_949,In_774);
nand U207 (N_207,In_595,In_1135);
or U208 (N_208,In_317,In_1486);
nand U209 (N_209,In_611,In_1214);
nor U210 (N_210,In_321,In_1984);
or U211 (N_211,In_622,In_103);
or U212 (N_212,In_477,In_1520);
nand U213 (N_213,In_1708,In_374);
xnor U214 (N_214,In_987,In_212);
nand U215 (N_215,In_696,In_34);
and U216 (N_216,In_1641,In_1801);
xor U217 (N_217,In_1555,In_1249);
or U218 (N_218,In_1231,In_1335);
and U219 (N_219,In_1469,In_1962);
and U220 (N_220,In_397,In_107);
and U221 (N_221,In_930,In_592);
xor U222 (N_222,In_84,In_255);
and U223 (N_223,In_612,In_500);
and U224 (N_224,In_1377,In_354);
and U225 (N_225,In_89,In_1971);
and U226 (N_226,In_1265,In_1403);
xor U227 (N_227,In_514,In_1742);
nand U228 (N_228,In_1209,In_1567);
nand U229 (N_229,In_126,In_1813);
and U230 (N_230,In_1134,In_1574);
and U231 (N_231,In_1346,In_879);
nor U232 (N_232,In_1918,In_1494);
and U233 (N_233,In_789,In_691);
and U234 (N_234,In_828,In_1784);
nor U235 (N_235,In_1870,In_1601);
and U236 (N_236,In_1631,In_1339);
xnor U237 (N_237,In_1608,In_1224);
xnor U238 (N_238,In_935,In_127);
nor U239 (N_239,In_556,In_1701);
xor U240 (N_240,In_833,In_228);
xor U241 (N_241,In_448,In_1074);
nor U242 (N_242,In_443,In_245);
nor U243 (N_243,In_1765,In_749);
and U244 (N_244,In_1961,In_432);
or U245 (N_245,In_648,In_311);
and U246 (N_246,In_176,In_1321);
nand U247 (N_247,In_1629,In_947);
nand U248 (N_248,In_916,In_336);
or U249 (N_249,In_1379,In_498);
and U250 (N_250,In_1734,In_1545);
and U251 (N_251,In_1046,In_272);
xor U252 (N_252,In_1280,In_1440);
nor U253 (N_253,In_501,In_110);
and U254 (N_254,In_79,In_787);
nor U255 (N_255,In_1720,In_524);
xnor U256 (N_256,In_1581,In_1478);
and U257 (N_257,In_1579,In_654);
nand U258 (N_258,In_1285,In_358);
or U259 (N_259,In_632,In_593);
xnor U260 (N_260,In_1809,In_65);
xor U261 (N_261,In_1422,In_1527);
nand U262 (N_262,In_1370,In_1406);
nor U263 (N_263,In_85,In_299);
nor U264 (N_264,In_673,In_1552);
and U265 (N_265,In_277,In_837);
nand U266 (N_266,In_1010,In_706);
nor U267 (N_267,In_850,In_1592);
nor U268 (N_268,In_60,In_617);
nor U269 (N_269,In_977,In_864);
nand U270 (N_270,In_1295,In_1006);
xor U271 (N_271,In_964,In_613);
or U272 (N_272,In_74,In_1369);
nor U273 (N_273,In_1510,In_1456);
nand U274 (N_274,In_115,In_969);
or U275 (N_275,In_1031,In_1839);
or U276 (N_276,In_304,In_810);
or U277 (N_277,In_510,In_1460);
nor U278 (N_278,In_1376,In_1383);
or U279 (N_279,In_970,In_1841);
nor U280 (N_280,In_860,In_335);
and U281 (N_281,In_1681,In_388);
nor U282 (N_282,In_815,In_361);
xnor U283 (N_283,In_1610,In_1251);
xnor U284 (N_284,In_1648,In_1789);
nor U285 (N_285,In_1889,In_1232);
xor U286 (N_286,In_300,In_533);
nand U287 (N_287,In_714,In_1300);
nor U288 (N_288,In_51,In_457);
xnor U289 (N_289,In_1503,In_1713);
or U290 (N_290,In_1205,In_1942);
xor U291 (N_291,In_637,In_1602);
or U292 (N_292,In_1800,In_167);
or U293 (N_293,In_631,In_1587);
xnor U294 (N_294,In_425,In_807);
or U295 (N_295,In_13,In_284);
or U296 (N_296,In_1041,In_1646);
nand U297 (N_297,In_1131,In_1024);
or U298 (N_298,In_1843,In_537);
nor U299 (N_299,In_1033,In_890);
and U300 (N_300,In_522,In_1442);
xnor U301 (N_301,In_1271,In_138);
or U302 (N_302,In_1258,In_965);
and U303 (N_303,In_122,In_169);
nand U304 (N_304,In_476,In_1026);
nor U305 (N_305,In_600,In_1400);
and U306 (N_306,In_1711,In_1966);
nand U307 (N_307,In_1909,In_1819);
xor U308 (N_308,In_171,In_1350);
nand U309 (N_309,In_1462,In_1177);
nand U310 (N_310,In_455,In_1855);
and U311 (N_311,In_931,In_603);
or U312 (N_312,In_1914,In_1558);
nor U313 (N_313,In_231,In_630);
xnor U314 (N_314,In_1101,In_170);
and U315 (N_315,In_128,In_1325);
or U316 (N_316,In_1680,In_1308);
and U317 (N_317,In_1319,In_1955);
nand U318 (N_318,In_1079,In_734);
xnor U319 (N_319,In_238,In_1729);
xnor U320 (N_320,In_253,In_544);
nor U321 (N_321,In_42,In_713);
nor U322 (N_322,In_1123,In_1874);
xnor U323 (N_323,In_69,In_1326);
nand U324 (N_324,In_519,In_1297);
or U325 (N_325,In_435,In_417);
or U326 (N_326,In_261,In_1960);
xor U327 (N_327,In_1397,In_423);
xnor U328 (N_328,In_1203,In_1563);
nor U329 (N_329,In_454,In_1725);
or U330 (N_330,In_1368,In_1227);
nor U331 (N_331,In_1405,In_1402);
and U332 (N_332,In_331,In_1366);
nand U333 (N_333,In_1810,In_274);
or U334 (N_334,In_874,In_1181);
and U335 (N_335,In_395,In_95);
nor U336 (N_336,In_7,In_1764);
nor U337 (N_337,In_1732,In_132);
or U338 (N_338,In_1080,In_1879);
nand U339 (N_339,In_1735,In_619);
or U340 (N_340,In_982,In_262);
nand U341 (N_341,In_237,In_569);
nand U342 (N_342,In_830,In_1304);
and U343 (N_343,In_695,In_217);
nand U344 (N_344,In_1736,In_332);
xnor U345 (N_345,In_310,In_1791);
and U346 (N_346,In_241,In_1167);
nor U347 (N_347,In_979,In_1439);
and U348 (N_348,In_554,In_1436);
nand U349 (N_349,In_763,In_639);
or U350 (N_350,In_1081,In_1145);
xor U351 (N_351,In_1474,In_1968);
or U352 (N_352,In_1144,In_129);
or U353 (N_353,In_345,In_1684);
or U354 (N_354,In_1670,In_772);
and U355 (N_355,In_1928,In_1861);
nand U356 (N_356,In_434,In_1834);
and U357 (N_357,In_1686,In_428);
nand U358 (N_358,In_1553,In_878);
xnor U359 (N_359,In_249,In_1199);
or U360 (N_360,In_991,In_666);
or U361 (N_361,In_808,In_260);
or U362 (N_362,In_1647,In_1132);
nand U363 (N_363,In_334,In_1022);
nor U364 (N_364,In_948,In_1213);
or U365 (N_365,In_1922,In_1259);
or U366 (N_366,In_888,In_1582);
nand U367 (N_367,In_1950,In_1788);
xnor U368 (N_368,In_28,In_452);
or U369 (N_369,In_1790,In_1980);
and U370 (N_370,In_941,In_337);
or U371 (N_371,In_707,In_1322);
nand U372 (N_372,In_1336,In_918);
and U373 (N_373,In_950,In_1193);
nand U374 (N_374,In_584,In_1082);
or U375 (N_375,In_929,In_464);
and U376 (N_376,In_1885,In_757);
and U377 (N_377,In_862,In_1544);
and U378 (N_378,In_329,In_1299);
nor U379 (N_379,In_985,In_996);
xor U380 (N_380,In_1417,In_1915);
or U381 (N_381,In_543,In_1187);
and U382 (N_382,In_1607,In_572);
xnor U383 (N_383,In_92,In_1910);
and U384 (N_384,In_152,In_682);
nor U385 (N_385,In_1974,In_1217);
nand U386 (N_386,In_992,In_967);
xor U387 (N_387,In_1569,In_1782);
or U388 (N_388,In_1244,In_16);
nor U389 (N_389,In_348,In_77);
nand U390 (N_390,In_1157,In_285);
xnor U391 (N_391,In_489,In_438);
nor U392 (N_392,In_1154,In_1221);
nand U393 (N_393,In_1946,In_399);
nor U394 (N_394,In_685,In_487);
and U395 (N_395,In_634,In_227);
and U396 (N_396,In_349,In_646);
nor U397 (N_397,In_1655,In_1091);
or U398 (N_398,In_1963,In_327);
and U399 (N_399,In_1237,In_511);
nor U400 (N_400,In_1455,In_151);
or U401 (N_401,In_1769,In_699);
nor U402 (N_402,In_739,In_1018);
or U403 (N_403,In_1932,In_1964);
and U404 (N_404,In_280,In_733);
nor U405 (N_405,In_407,In_389);
or U406 (N_406,In_1160,In_1344);
xor U407 (N_407,In_39,In_999);
nand U408 (N_408,In_1489,In_292);
xor U409 (N_409,In_1820,In_446);
xor U410 (N_410,In_409,In_951);
xnor U411 (N_411,In_1386,In_1195);
nand U412 (N_412,In_1223,In_1583);
and U413 (N_413,In_22,In_1286);
or U414 (N_414,In_254,In_475);
and U415 (N_415,In_322,In_53);
nor U416 (N_416,In_1990,In_445);
nand U417 (N_417,In_1445,In_142);
and U418 (N_418,In_1042,In_347);
nor U419 (N_419,In_195,In_1515);
nand U420 (N_420,In_895,In_1250);
nand U421 (N_421,In_1866,In_927);
and U422 (N_422,In_1998,In_460);
xor U423 (N_423,In_1148,In_602);
nor U424 (N_424,In_1334,In_1363);
nor U425 (N_425,In_585,In_1355);
nor U426 (N_426,In_10,In_314);
nand U427 (N_427,In_1662,In_114);
and U428 (N_428,In_1873,In_1367);
xnor U429 (N_429,In_458,In_759);
xor U430 (N_430,In_1292,In_419);
and U431 (N_431,In_1045,In_140);
and U432 (N_432,In_1055,In_1428);
or U433 (N_433,In_470,In_1260);
and U434 (N_434,In_323,In_1303);
and U435 (N_435,In_119,In_55);
or U436 (N_436,In_978,In_1745);
xnor U437 (N_437,In_229,In_31);
nand U438 (N_438,In_783,In_307);
nand U439 (N_439,In_1624,In_1858);
and U440 (N_440,In_1845,In_216);
and U441 (N_441,In_605,In_1168);
xor U442 (N_442,In_1020,In_1067);
nor U443 (N_443,In_471,In_698);
and U444 (N_444,In_1716,In_606);
nand U445 (N_445,In_1718,In_1854);
xnor U446 (N_446,In_453,In_627);
nor U447 (N_447,In_1900,In_748);
or U448 (N_448,In_1871,In_1179);
nor U449 (N_449,In_1744,In_751);
nand U450 (N_450,In_1278,In_1107);
or U451 (N_451,In_1538,In_1356);
and U452 (N_452,In_418,In_1243);
or U453 (N_453,In_889,In_1204);
xnor U454 (N_454,In_744,In_1463);
or U455 (N_455,In_344,In_281);
nor U456 (N_456,In_1862,In_876);
or U457 (N_457,In_1781,In_1467);
or U458 (N_458,In_1257,In_1886);
nand U459 (N_459,In_1450,In_1753);
nand U460 (N_460,In_1674,In_1449);
and U461 (N_461,In_571,In_1755);
xnor U462 (N_462,In_1995,In_449);
or U463 (N_463,In_1969,In_1337);
nor U464 (N_464,In_683,In_251);
or U465 (N_465,In_858,In_58);
nand U466 (N_466,In_346,In_832);
nand U467 (N_467,In_1831,In_424);
and U468 (N_468,In_29,In_466);
and U469 (N_469,In_1272,In_1459);
nor U470 (N_470,In_643,In_805);
xnor U471 (N_471,In_1622,In_450);
and U472 (N_472,In_909,In_1652);
nand U473 (N_473,In_210,In_596);
nor U474 (N_474,In_884,In_357);
or U475 (N_475,In_433,In_1318);
or U476 (N_476,In_1508,In_867);
nor U477 (N_477,In_369,In_781);
nor U478 (N_478,In_1283,In_1929);
and U479 (N_479,In_30,In_410);
or U480 (N_480,In_1371,In_1448);
and U481 (N_481,In_1408,In_755);
or U482 (N_482,In_1340,In_1076);
nand U483 (N_483,In_175,In_728);
nor U484 (N_484,In_1281,In_902);
xor U485 (N_485,In_791,In_1632);
and U486 (N_486,In_1757,In_297);
or U487 (N_487,In_80,In_942);
xor U488 (N_488,In_1868,In_1332);
xor U489 (N_489,In_269,In_1044);
and U490 (N_490,In_835,In_1190);
nand U491 (N_491,In_1097,In_661);
nand U492 (N_492,In_1588,In_81);
nor U493 (N_493,In_1361,In_697);
or U494 (N_494,In_1039,In_381);
nand U495 (N_495,In_68,In_1642);
nand U496 (N_496,In_1653,In_1710);
and U497 (N_497,In_756,In_1565);
xor U498 (N_498,In_681,In_246);
xnor U499 (N_499,In_920,In_652);
or U500 (N_500,In_1921,In_1795);
xor U501 (N_501,In_1419,In_1715);
and U502 (N_502,In_509,In_1712);
or U503 (N_503,N_461,In_1277);
xnor U504 (N_504,In_1485,N_387);
or U505 (N_505,In_1661,In_1549);
nor U506 (N_506,N_311,In_1978);
xnor U507 (N_507,N_476,N_149);
and U508 (N_508,In_1004,N_107);
and U509 (N_509,In_37,In_1507);
and U510 (N_510,N_477,In_1169);
or U511 (N_511,In_400,In_1779);
and U512 (N_512,N_98,N_300);
nor U513 (N_513,N_41,In_1095);
and U514 (N_514,In_777,In_1345);
and U515 (N_515,N_15,N_5);
nand U516 (N_516,In_1468,In_1175);
or U517 (N_517,In_1100,N_96);
or U518 (N_518,In_213,In_1890);
or U519 (N_519,N_76,In_963);
nor U520 (N_520,N_455,In_271);
nor U521 (N_521,N_71,In_928);
nand U522 (N_522,In_1118,N_200);
and U523 (N_523,N_373,N_213);
nor U524 (N_524,In_474,In_997);
or U525 (N_525,In_1596,In_1306);
nor U526 (N_526,N_441,N_434);
or U527 (N_527,In_1901,In_1099);
or U528 (N_528,In_1309,N_372);
or U529 (N_529,N_312,N_398);
nor U530 (N_530,In_1983,In_1501);
and U531 (N_531,N_334,N_123);
or U532 (N_532,In_564,In_806);
or U533 (N_533,In_66,In_607);
nor U534 (N_534,In_960,In_1627);
or U535 (N_535,N_313,In_1530);
and U536 (N_536,In_1092,In_382);
xnor U537 (N_537,N_296,In_1775);
nor U538 (N_538,In_826,In_1759);
nor U539 (N_539,N_192,In_429);
or U540 (N_540,In_1637,N_290);
nor U541 (N_541,In_1654,In_391);
nand U542 (N_542,In_1724,N_427);
nand U543 (N_543,In_679,In_62);
and U544 (N_544,N_72,N_177);
nor U545 (N_545,In_118,N_390);
and U546 (N_546,N_407,In_670);
and U547 (N_547,In_993,N_191);
nor U548 (N_548,In_1934,In_1047);
and U549 (N_549,N_487,N_499);
or U550 (N_550,In_1750,N_308);
nor U551 (N_551,N_86,In_379);
nor U552 (N_552,N_113,N_406);
nor U553 (N_553,In_1842,N_247);
nor U554 (N_554,In_1829,In_473);
nand U555 (N_555,In_373,In_998);
and U556 (N_556,In_125,In_1427);
nor U557 (N_557,N_248,N_282);
or U558 (N_558,In_242,In_25);
or U559 (N_559,N_80,N_362);
and U560 (N_560,In_1762,In_1697);
or U561 (N_561,N_424,In_642);
or U562 (N_562,N_285,In_214);
nor U563 (N_563,In_1372,N_433);
xor U564 (N_564,N_227,N_131);
and U565 (N_565,In_295,In_1360);
nand U566 (N_566,N_397,In_1606);
and U567 (N_567,In_1385,In_937);
and U568 (N_568,In_545,In_1945);
nor U569 (N_569,N_325,In_1733);
and U570 (N_570,In_750,In_444);
nand U571 (N_571,In_2,In_153);
xnor U572 (N_572,In_1110,In_589);
xnor U573 (N_573,In_557,In_725);
nand U574 (N_574,In_790,In_1691);
nor U575 (N_575,In_1938,N_482);
or U576 (N_576,In_715,N_47);
xor U577 (N_577,In_279,In_1902);
nand U578 (N_578,In_516,In_881);
nand U579 (N_579,In_1770,In_333);
nor U580 (N_580,In_291,In_919);
or U581 (N_581,In_1105,In_1311);
xor U582 (N_582,In_306,N_489);
and U583 (N_583,N_229,N_422);
or U584 (N_584,N_148,In_897);
xor U585 (N_585,In_1248,N_10);
or U586 (N_586,N_190,In_485);
nand U587 (N_587,In_1988,In_405);
nor U588 (N_588,In_703,N_167);
nor U589 (N_589,N_180,N_297);
or U590 (N_590,In_1643,N_347);
or U591 (N_591,In_1158,In_495);
or U592 (N_592,N_498,In_582);
and U593 (N_593,In_1999,In_680);
xor U594 (N_594,In_1638,In_1651);
nand U595 (N_595,In_185,In_472);
and U596 (N_596,In_1056,N_19);
nand U597 (N_597,In_192,N_197);
nor U598 (N_598,In_1917,In_1837);
nand U599 (N_599,In_1893,N_22);
nand U600 (N_600,In_690,N_234);
nor U601 (N_601,N_179,In_1649);
nand U602 (N_602,In_1594,In_1410);
or U603 (N_603,N_233,In_1836);
or U604 (N_604,In_1600,N_114);
or U605 (N_605,In_1287,N_94);
or U606 (N_606,In_1245,N_232);
nor U607 (N_607,In_1746,In_532);
xnor U608 (N_608,In_1161,N_274);
nor U609 (N_609,N_212,In_1907);
or U610 (N_610,In_1252,In_1511);
nand U611 (N_611,In_555,In_865);
and U612 (N_612,N_216,In_1529);
nor U613 (N_613,In_4,N_186);
and U614 (N_614,N_294,In_1693);
xor U615 (N_615,In_1763,In_1274);
and U616 (N_616,In_1537,In_416);
nand U617 (N_617,In_1920,In_184);
and U618 (N_618,In_390,In_302);
and U619 (N_619,In_113,In_1991);
nor U620 (N_620,In_288,In_745);
or U621 (N_621,In_1717,In_247);
or U622 (N_622,In_1751,In_106);
xor U623 (N_623,In_1919,N_122);
and U624 (N_624,In_49,In_173);
or U625 (N_625,In_813,In_1878);
nor U626 (N_626,N_30,N_472);
nor U627 (N_627,In_823,In_1706);
xor U628 (N_628,In_1314,In_1215);
and U629 (N_629,In_980,In_575);
nand U630 (N_630,In_1756,In_1951);
or U631 (N_631,In_1207,N_160);
and U632 (N_632,N_188,N_411);
xor U633 (N_633,In_1451,In_838);
nor U634 (N_634,In_770,In_1573);
nor U635 (N_635,N_465,In_1381);
xor U636 (N_636,N_473,In_1516);
or U637 (N_637,In_1038,N_306);
and U638 (N_638,In_159,In_1437);
or U639 (N_639,In_1093,In_15);
nor U640 (N_640,N_193,In_1694);
and U641 (N_641,In_1993,In_1804);
nor U642 (N_642,N_298,In_1341);
xnor U643 (N_643,N_159,In_1426);
or U644 (N_644,N_272,In_540);
nor U645 (N_645,In_320,N_262);
xor U646 (N_646,In_1202,In_936);
nor U647 (N_647,In_1275,N_439);
xor U648 (N_648,In_3,In_1621);
xnor U649 (N_649,N_337,In_1512);
xor U650 (N_650,N_224,In_385);
nand U651 (N_651,N_42,In_988);
nand U652 (N_652,N_417,In_1166);
xnor U653 (N_653,In_1521,In_1497);
nor U654 (N_654,In_1525,In_76);
and U655 (N_655,In_717,N_56);
xnor U656 (N_656,In_403,N_51);
nor U657 (N_657,In_1833,In_708);
xor U658 (N_658,In_1740,In_1658);
xor U659 (N_659,In_483,In_482);
or U660 (N_660,In_913,In_678);
xnor U661 (N_661,N_176,In_1310);
nand U662 (N_662,In_1543,In_795);
or U663 (N_663,N_432,In_660);
and U664 (N_664,In_1294,N_369);
nand U665 (N_665,In_871,N_403);
xnor U666 (N_666,N_151,In_276);
and U667 (N_667,In_1797,In_1673);
or U668 (N_668,In_1888,In_359);
and U669 (N_669,In_1212,N_389);
or U670 (N_670,In_190,N_0);
nand U671 (N_671,N_365,In_1234);
or U672 (N_672,In_1598,In_880);
and U673 (N_673,N_118,In_1766);
nand U674 (N_674,N_437,N_310);
and U675 (N_675,N_275,N_53);
and U676 (N_676,In_1933,In_1977);
nor U677 (N_677,In_1,In_1575);
nand U678 (N_678,In_1869,In_923);
and U679 (N_679,In_1835,In_1472);
nor U680 (N_680,In_821,In_372);
xor U681 (N_681,N_23,In_1293);
and U682 (N_682,In_1117,In_505);
nand U683 (N_683,In_1822,N_414);
and U684 (N_684,N_267,In_903);
nand U685 (N_685,N_382,N_253);
or U686 (N_686,N_116,In_1924);
xnor U687 (N_687,N_84,In_863);
and U688 (N_688,N_73,N_45);
xor U689 (N_689,In_786,In_1617);
or U690 (N_690,N_235,N_359);
xnor U691 (N_691,N_48,In_1850);
nand U692 (N_692,In_565,In_1666);
or U693 (N_693,In_1071,In_462);
nor U694 (N_694,N_319,In_20);
nor U695 (N_695,In_1650,In_1899);
and U696 (N_696,In_1479,In_290);
xnor U697 (N_697,N_185,N_450);
nand U698 (N_698,In_355,In_1390);
nor U699 (N_699,In_1778,N_355);
nand U700 (N_700,In_1794,In_1130);
xnor U701 (N_701,In_896,In_1722);
and U702 (N_702,In_552,In_99);
and U703 (N_703,N_302,In_1062);
nor U704 (N_704,In_1078,In_1799);
and U705 (N_705,N_2,In_396);
or U706 (N_706,In_258,N_462);
or U707 (N_707,N_448,In_1296);
or U708 (N_708,In_88,In_367);
or U709 (N_709,In_1351,In_1023);
and U710 (N_710,In_1013,In_1241);
or U711 (N_711,N_318,N_361);
or U712 (N_712,In_1818,In_197);
nand U713 (N_713,In_1702,N_493);
nand U714 (N_714,N_173,N_103);
nand U715 (N_715,N_345,In_1083);
or U716 (N_716,In_1589,In_1142);
nand U717 (N_717,N_115,In_56);
and U718 (N_718,N_49,In_273);
or U719 (N_719,In_366,In_82);
nor U720 (N_720,In_117,N_305);
or U721 (N_721,N_95,In_563);
xor U722 (N_722,In_1050,N_65);
nand U723 (N_723,N_388,In_861);
nor U724 (N_724,In_23,In_201);
nand U725 (N_725,In_1656,N_241);
xor U726 (N_726,N_292,In_972);
nand U727 (N_727,N_136,In_268);
nand U728 (N_728,N_101,In_1064);
and U729 (N_729,In_827,In_836);
or U730 (N_730,In_1739,In_1678);
xnor U731 (N_731,N_364,N_242);
and U732 (N_732,In_1452,In_1009);
and U733 (N_733,In_148,In_393);
nand U734 (N_734,In_753,N_444);
and U735 (N_735,In_182,In_1016);
nor U736 (N_736,In_154,N_279);
and U737 (N_737,N_341,In_957);
or U738 (N_738,In_1996,N_215);
or U739 (N_739,In_1388,N_237);
nor U740 (N_740,N_425,In_769);
and U741 (N_741,In_1639,In_1707);
or U742 (N_742,N_440,In_899);
or U743 (N_743,In_1672,N_323);
nor U744 (N_744,In_1229,N_386);
or U745 (N_745,In_1473,N_78);
or U746 (N_746,In_1288,In_521);
or U747 (N_747,N_126,In_1965);
nor U748 (N_748,In_911,N_29);
or U749 (N_749,In_614,In_925);
nand U750 (N_750,In_120,In_204);
xnor U751 (N_751,In_136,In_1114);
or U752 (N_752,In_1077,N_349);
xnor U753 (N_753,In_1683,N_286);
and U754 (N_754,N_420,N_481);
xnor U755 (N_755,N_479,N_332);
nand U756 (N_756,N_60,In_206);
nand U757 (N_757,In_1185,N_491);
or U758 (N_758,In_665,In_1882);
xnor U759 (N_759,In_220,In_1528);
nand U760 (N_760,N_106,N_194);
nor U761 (N_761,In_778,In_256);
and U762 (N_762,N_436,N_281);
nand U763 (N_763,N_172,N_206);
or U764 (N_764,N_451,N_459);
xnor U765 (N_765,N_187,In_1302);
nand U766 (N_766,In_1108,N_399);
and U767 (N_767,In_301,N_82);
and U768 (N_768,In_1737,In_146);
nand U769 (N_769,N_273,In_1113);
and U770 (N_770,N_431,In_1365);
nand U771 (N_771,In_1150,In_1832);
or U772 (N_772,In_1760,In_672);
nor U773 (N_773,In_91,N_246);
nor U774 (N_774,N_463,In_1912);
nand U775 (N_775,In_1089,In_293);
and U776 (N_776,In_677,In_406);
nand U777 (N_777,N_485,N_154);
and U778 (N_778,In_1119,N_196);
and U779 (N_779,N_11,In_580);
nor U780 (N_780,In_1431,In_767);
nand U781 (N_781,In_1219,In_1848);
nor U782 (N_782,In_684,N_37);
nand U783 (N_783,In_1916,In_1826);
nor U784 (N_784,N_426,In_158);
or U785 (N_785,N_132,In_1480);
or U786 (N_786,In_375,N_327);
nand U787 (N_787,In_956,In_422);
xor U788 (N_788,In_583,N_263);
nor U789 (N_789,N_214,N_3);
nor U790 (N_790,N_475,N_340);
or U791 (N_791,In_1613,N_402);
and U792 (N_792,In_1821,N_494);
or U793 (N_793,N_360,In_1353);
nand U794 (N_794,N_16,In_1357);
nor U795 (N_795,In_412,In_921);
xnor U796 (N_796,In_1571,In_1396);
and U797 (N_797,In_1354,N_418);
or U798 (N_798,In_221,N_169);
nand U799 (N_799,In_1593,In_1805);
xnor U800 (N_800,N_374,N_478);
and U801 (N_801,N_348,In_111);
or U802 (N_802,In_305,In_1591);
and U803 (N_803,In_177,In_1506);
xor U804 (N_804,In_468,In_1425);
and U805 (N_805,N_429,N_356);
xnor U806 (N_806,In_14,In_1151);
nor U807 (N_807,In_1940,N_423);
xor U808 (N_808,In_1191,In_1771);
and U809 (N_809,N_140,N_1);
and U810 (N_810,N_63,In_1171);
or U811 (N_811,In_1374,In_1115);
xor U812 (N_812,In_633,In_934);
and U813 (N_813,In_1905,In_1471);
or U814 (N_814,In_1021,In_265);
nor U815 (N_815,N_70,In_731);
and U816 (N_816,N_64,In_688);
or U817 (N_817,In_198,In_1863);
nor U818 (N_818,In_459,N_243);
nand U819 (N_819,N_165,N_93);
nand U820 (N_820,N_385,In_499);
nand U821 (N_821,N_483,N_321);
xnor U822 (N_822,In_1189,In_736);
nor U823 (N_823,N_351,N_166);
xnor U824 (N_824,In_303,In_1894);
xnor U825 (N_825,In_90,In_1327);
xnor U826 (N_826,In_793,In_1768);
and U827 (N_827,In_1466,In_1628);
or U828 (N_828,In_1373,In_180);
nor U829 (N_829,In_1262,N_363);
nand U830 (N_830,N_486,In_1692);
xor U831 (N_831,In_1767,N_328);
or U832 (N_832,In_1011,N_404);
nand U833 (N_833,In_1743,In_54);
or U834 (N_834,In_259,In_724);
and U835 (N_835,N_170,N_120);
nor U836 (N_836,In_232,N_121);
or U837 (N_837,In_1872,N_57);
nor U838 (N_838,In_187,In_196);
xnor U839 (N_839,N_108,In_447);
or U840 (N_840,In_517,N_320);
nand U841 (N_841,In_854,N_54);
nor U842 (N_842,In_309,In_19);
or U843 (N_843,In_451,N_336);
or U844 (N_844,N_409,In_224);
nand U845 (N_845,In_910,In_1015);
and U846 (N_846,In_1948,In_17);
nor U847 (N_847,In_525,N_304);
and U848 (N_848,N_18,In_1002);
nor U849 (N_849,In_1264,In_1276);
nor U850 (N_850,In_1540,In_629);
xor U851 (N_851,N_152,In_1586);
nand U852 (N_852,In_752,In_1853);
xor U853 (N_853,In_78,In_689);
nor U854 (N_854,In_326,N_326);
xor U855 (N_855,In_566,In_1032);
nor U856 (N_856,In_1585,In_645);
xnor U857 (N_857,In_1454,N_375);
xor U858 (N_858,N_339,In_1796);
and U859 (N_859,In_41,In_1644);
and U860 (N_860,In_378,In_971);
or U861 (N_861,N_307,In_1619);
nor U862 (N_862,In_1534,In_1164);
nand U863 (N_863,In_239,N_458);
xor U864 (N_864,In_794,In_1554);
nor U865 (N_865,In_711,In_1482);
nand U866 (N_866,N_400,N_6);
and U867 (N_867,In_1389,In_1604);
nor U868 (N_868,In_1129,N_416);
nand U869 (N_869,In_1541,N_309);
nor U870 (N_870,In_1464,In_848);
xnor U871 (N_871,In_1435,In_61);
or U872 (N_872,In_841,N_357);
nor U873 (N_873,N_413,In_328);
nand U874 (N_874,In_771,In_1535);
xnor U875 (N_875,N_184,N_240);
or U876 (N_876,In_1182,In_668);
and U877 (N_877,In_47,In_822);
nand U878 (N_878,In_694,N_97);
or U879 (N_879,In_1518,In_624);
nor U880 (N_880,N_303,In_1925);
xnor U881 (N_881,In_558,In_1094);
nor U882 (N_882,In_1887,In_727);
xnor U883 (N_883,N_141,In_812);
nand U884 (N_884,In_1411,N_333);
xor U885 (N_885,In_766,N_111);
nand U886 (N_886,In_1324,In_420);
nor U887 (N_887,In_1282,In_1153);
and U888 (N_888,In_547,In_1935);
nand U889 (N_889,In_1457,In_782);
nand U890 (N_890,In_1747,In_801);
nor U891 (N_891,In_376,In_799);
nand U892 (N_892,In_1667,N_219);
nor U893 (N_893,In_1273,In_1012);
nor U894 (N_894,In_1664,In_1927);
and U895 (N_895,In_908,In_200);
xnor U896 (N_896,In_342,In_437);
or U897 (N_897,N_146,In_1985);
or U898 (N_898,In_83,In_1096);
nor U899 (N_899,In_233,In_1802);
or U900 (N_900,In_1152,In_282);
or U901 (N_901,In_1513,N_88);
or U902 (N_902,In_926,In_700);
nor U903 (N_903,N_17,In_1008);
nor U904 (N_904,N_139,In_240);
and U905 (N_905,In_989,N_182);
or U906 (N_906,N_244,N_324);
nand U907 (N_907,N_155,N_105);
and U908 (N_908,In_353,In_141);
xnor U909 (N_909,In_270,In_26);
xor U910 (N_910,N_412,N_8);
xnor U911 (N_911,In_1137,In_202);
nor U912 (N_912,In_853,N_236);
nand U913 (N_913,N_410,In_230);
nand U914 (N_914,In_121,N_394);
nor U915 (N_915,N_379,N_238);
xnor U916 (N_916,In_1186,In_12);
nor U917 (N_917,In_1291,In_1659);
xnor U918 (N_918,In_1124,N_75);
and U919 (N_919,In_1254,N_59);
or U920 (N_920,N_396,N_446);
nor U921 (N_921,N_183,In_1599);
xnor U922 (N_922,In_287,In_1060);
or U923 (N_923,In_885,In_892);
and U924 (N_924,In_1484,N_55);
or U925 (N_925,In_1007,In_1218);
xor U926 (N_926,N_250,N_153);
or U927 (N_927,N_354,N_195);
nor U928 (N_928,In_131,N_331);
and U929 (N_929,N_383,N_314);
nand U930 (N_930,In_726,In_776);
and U931 (N_931,N_284,In_508);
nand U932 (N_932,In_548,In_1857);
or U933 (N_933,N_299,N_469);
xor U934 (N_934,N_480,In_205);
nor U935 (N_935,In_278,In_1903);
nand U936 (N_936,In_636,N_145);
xor U937 (N_937,In_651,N_91);
nand U938 (N_938,In_824,N_230);
or U939 (N_939,In_1926,In_1851);
and U940 (N_940,In_492,In_898);
nand U941 (N_941,In_163,In_831);
xor U942 (N_942,In_1816,N_36);
xor U943 (N_943,N_384,In_1550);
nor U944 (N_944,In_1267,In_1141);
nand U945 (N_945,In_856,In_1420);
and U946 (N_946,In_223,N_92);
nand U947 (N_947,In_1726,In_1030);
and U948 (N_948,N_156,N_207);
nand U949 (N_949,In_1844,In_155);
nand U950 (N_950,In_961,In_811);
nor U951 (N_951,In_440,N_378);
nand U952 (N_952,In_1104,N_44);
nand U953 (N_953,N_443,In_515);
xnor U954 (N_954,N_401,In_1358);
nor U955 (N_955,N_466,In_319);
xnor U956 (N_956,In_1533,In_494);
and U957 (N_957,N_39,In_709);
or U958 (N_958,N_471,In_720);
xor U959 (N_959,In_647,In_520);
xor U960 (N_960,N_112,N_69);
and U961 (N_961,N_61,N_495);
nand U962 (N_962,In_1174,N_391);
nor U963 (N_963,N_415,In_1247);
and U964 (N_964,N_454,In_97);
and U965 (N_965,In_894,N_171);
nand U966 (N_966,N_33,In_467);
xor U967 (N_967,In_526,N_168);
nand U968 (N_968,N_317,In_1127);
xnor U969 (N_969,In_663,N_198);
and U970 (N_970,In_257,In_1603);
and U971 (N_971,In_1183,In_1677);
or U972 (N_972,In_33,N_291);
nor U973 (N_973,In_392,In_398);
nand U974 (N_974,In_411,In_11);
nand U975 (N_975,In_765,In_64);
xnor U976 (N_976,N_370,In_1465);
nand U977 (N_977,In_161,N_252);
or U978 (N_978,In_316,In_742);
or U979 (N_979,N_202,N_85);
nor U980 (N_980,In_1777,In_1898);
nand U981 (N_981,N_143,In_343);
nand U982 (N_982,In_264,In_360);
xor U983 (N_983,N_492,In_1695);
or U984 (N_984,N_158,In_1444);
xor U985 (N_985,In_1256,In_650);
nor U986 (N_986,In_1787,In_72);
or U987 (N_987,In_1305,N_162);
or U988 (N_988,In_829,In_86);
nand U989 (N_989,In_430,N_342);
and U990 (N_990,N_497,In_1058);
and U991 (N_991,In_362,In_1676);
nor U992 (N_992,N_338,In_1847);
or U993 (N_993,N_218,In_1741);
or U994 (N_994,N_266,In_1526);
and U995 (N_995,In_243,N_74);
nand U996 (N_996,In_1941,In_408);
and U997 (N_997,N_134,In_27);
or U998 (N_998,N_408,N_377);
nor U999 (N_999,N_322,In_235);
nand U1000 (N_1000,N_225,N_631);
and U1001 (N_1001,N_611,N_702);
nor U1002 (N_1002,N_102,N_778);
or U1003 (N_1003,N_926,N_707);
nor U1004 (N_1004,In_623,N_430);
xor U1005 (N_1005,N_817,In_1772);
nand U1006 (N_1006,In_178,N_563);
nor U1007 (N_1007,In_851,N_52);
or U1008 (N_1008,N_632,N_548);
or U1009 (N_1009,In_579,N_996);
or U1010 (N_1010,N_556,N_518);
and U1011 (N_1011,N_899,N_960);
nand U1012 (N_1012,N_888,In_712);
and U1013 (N_1013,In_1814,N_83);
nand U1014 (N_1014,N_813,N_344);
and U1015 (N_1015,In_40,N_34);
nand U1016 (N_1016,N_175,N_825);
xnor U1017 (N_1017,In_1679,N_613);
nor U1018 (N_1018,N_615,N_128);
xnor U1019 (N_1019,N_438,In_939);
nor U1020 (N_1020,In_225,N_330);
xor U1021 (N_1021,N_792,N_217);
nor U1022 (N_1022,In_1066,N_514);
and U1023 (N_1023,In_1881,N_142);
or U1024 (N_1024,N_898,N_808);
nand U1025 (N_1025,N_496,N_289);
nand U1026 (N_1026,N_650,N_694);
and U1027 (N_1027,In_1849,In_1947);
or U1028 (N_1028,N_917,N_671);
xnor U1029 (N_1029,In_1808,N_755);
nand U1030 (N_1030,N_852,N_280);
nor U1031 (N_1031,In_983,N_834);
and U1032 (N_1032,N_405,In_1352);
or U1033 (N_1033,N_699,N_245);
nor U1034 (N_1034,In_1542,In_1897);
or U1035 (N_1035,In_1348,N_593);
or U1036 (N_1036,N_659,N_978);
nand U1037 (N_1037,N_643,N_958);
nor U1038 (N_1038,N_784,N_468);
xnor U1039 (N_1039,N_648,In_102);
nand U1040 (N_1040,N_622,N_768);
and U1041 (N_1041,N_823,In_568);
or U1042 (N_1042,N_594,N_666);
nor U1043 (N_1043,In_168,In_1758);
xnor U1044 (N_1044,In_746,In_1242);
or U1045 (N_1045,N_603,N_638);
or U1046 (N_1046,In_1423,N_315);
nor U1047 (N_1047,In_577,In_644);
and U1048 (N_1048,N_447,N_785);
nor U1049 (N_1049,In_1208,In_1752);
or U1050 (N_1050,N_535,N_929);
nand U1051 (N_1051,In_100,N_221);
or U1052 (N_1052,N_881,In_705);
or U1053 (N_1053,N_258,N_963);
xnor U1054 (N_1054,N_585,In_1704);
and U1055 (N_1055,N_517,N_617);
or U1056 (N_1056,N_681,In_1727);
nor U1057 (N_1057,N_343,N_110);
and U1058 (N_1058,N_791,N_844);
nand U1059 (N_1059,In_946,N_809);
and U1060 (N_1060,N_565,N_581);
nand U1061 (N_1061,N_979,N_862);
nor U1062 (N_1062,In_1393,N_876);
or U1063 (N_1063,In_181,N_829);
xor U1064 (N_1064,N_679,In_1487);
and U1065 (N_1065,N_124,In_1198);
nand U1066 (N_1066,N_738,In_1394);
and U1067 (N_1067,N_68,In_814);
or U1068 (N_1068,In_1035,In_729);
xnor U1069 (N_1069,N_922,N_634);
or U1070 (N_1070,In_1531,N_606);
nand U1071 (N_1071,N_977,N_419);
or U1072 (N_1072,N_226,In_1867);
and U1073 (N_1073,N_704,N_14);
or U1074 (N_1074,N_705,In_1846);
xnor U1075 (N_1075,N_949,N_395);
nor U1076 (N_1076,N_625,N_783);
or U1077 (N_1077,N_381,In_1192);
and U1078 (N_1078,N_586,N_203);
nor U1079 (N_1079,In_953,In_1546);
nor U1080 (N_1080,N_449,In_1194);
and U1081 (N_1081,N_596,N_729);
or U1082 (N_1082,In_1523,N_376);
or U1083 (N_1083,In_1685,N_740);
nand U1084 (N_1084,N_510,In_1806);
or U1085 (N_1085,In_1098,N_77);
nand U1086 (N_1086,N_627,N_26);
nor U1087 (N_1087,In_1037,N_691);
xnor U1088 (N_1088,In_1572,N_32);
and U1089 (N_1089,N_803,In_123);
nand U1090 (N_1090,N_665,N_754);
nor U1091 (N_1091,N_997,N_647);
xnor U1092 (N_1092,N_739,In_1268);
nand U1093 (N_1093,In_1539,N_368);
nand U1094 (N_1094,N_780,N_519);
and U1095 (N_1095,In_104,N_980);
nand U1096 (N_1096,N_27,N_689);
and U1097 (N_1097,In_75,N_505);
nor U1098 (N_1098,In_529,In_788);
nor U1099 (N_1099,N_900,In_1731);
xnor U1100 (N_1100,N_553,N_981);
or U1101 (N_1101,N_133,N_753);
and U1102 (N_1102,In_352,In_1027);
xnor U1103 (N_1103,N_927,N_688);
nand U1104 (N_1104,N_993,N_661);
xor U1105 (N_1105,N_574,N_804);
or U1106 (N_1106,N_641,In_1116);
nor U1107 (N_1107,In_530,N_748);
nand U1108 (N_1108,In_1496,In_283);
or U1109 (N_1109,N_873,In_1364);
xnor U1110 (N_1110,N_961,N_835);
nand U1111 (N_1111,In_1331,N_964);
and U1112 (N_1112,N_500,In_493);
or U1113 (N_1113,N_610,In_1399);
or U1114 (N_1114,In_166,N_520);
nor U1115 (N_1115,In_740,N_592);
nand U1116 (N_1116,N_524,N_90);
nor U1117 (N_1117,In_1147,N_658);
and U1118 (N_1118,N_764,N_144);
nor U1119 (N_1119,N_807,N_826);
xnor U1120 (N_1120,N_600,N_79);
or U1121 (N_1121,In_1576,N_119);
and U1122 (N_1122,N_800,N_529);
xor U1123 (N_1123,N_453,N_211);
nand U1124 (N_1124,In_465,N_637);
nand U1125 (N_1125,N_860,In_38);
and U1126 (N_1126,In_1102,N_569);
nor U1127 (N_1127,In_1892,N_870);
or U1128 (N_1128,In_250,In_1178);
xor U1129 (N_1129,N_912,N_690);
nand U1130 (N_1130,In_1073,In_1375);
xor U1131 (N_1131,In_912,In_365);
xor U1132 (N_1132,In_1085,In_843);
or U1133 (N_1133,In_108,N_838);
and U1134 (N_1134,In_1577,N_966);
xor U1135 (N_1135,N_867,N_547);
nand U1136 (N_1136,N_598,In_431);
and U1137 (N_1137,N_255,N_786);
xor U1138 (N_1138,N_653,N_117);
and U1139 (N_1139,N_787,N_591);
xor U1140 (N_1140,N_502,N_947);
or U1141 (N_1141,N_549,In_958);
xor U1142 (N_1142,N_670,In_219);
or U1143 (N_1143,In_1312,In_1967);
and U1144 (N_1144,N_21,N_575);
or U1145 (N_1145,N_770,N_710);
xor U1146 (N_1146,In_975,N_731);
or U1147 (N_1147,In_1502,In_1864);
nand U1148 (N_1148,N_828,In_1446);
or U1149 (N_1149,N_204,N_847);
nor U1150 (N_1150,In_1561,In_1392);
or U1151 (N_1151,In_1609,In_194);
nand U1152 (N_1152,N_692,N_868);
nand U1153 (N_1153,In_506,N_257);
xnor U1154 (N_1154,N_584,N_682);
or U1155 (N_1155,N_543,In_368);
xor U1156 (N_1156,N_352,N_712);
and U1157 (N_1157,In_325,N_507);
nand U1158 (N_1158,N_544,In_59);
xor U1159 (N_1159,N_295,N_767);
or U1160 (N_1160,N_935,In_70);
and U1161 (N_1161,N_725,In_490);
or U1162 (N_1162,In_1490,N_793);
nor U1163 (N_1163,N_820,In_626);
xor U1164 (N_1164,N_999,In_415);
nor U1165 (N_1165,In_298,N_35);
and U1166 (N_1166,In_551,N_40);
or U1167 (N_1167,In_628,In_1972);
nor U1168 (N_1168,In_1342,N_910);
nand U1169 (N_1169,N_589,In_561);
xor U1170 (N_1170,N_570,N_727);
nor U1171 (N_1171,N_608,N_38);
or U1172 (N_1172,In_535,In_1139);
and U1173 (N_1173,N_649,N_685);
or U1174 (N_1174,In_1475,In_1690);
xnor U1175 (N_1175,N_660,N_189);
nor U1176 (N_1176,N_655,N_223);
or U1177 (N_1177,N_781,N_861);
or U1178 (N_1178,In_1382,In_414);
or U1179 (N_1179,N_677,N_129);
xor U1180 (N_1180,N_722,In_1121);
xnor U1181 (N_1181,In_723,In_773);
nand U1182 (N_1182,In_1620,In_263);
xor U1183 (N_1183,In_1106,N_837);
or U1184 (N_1184,N_668,N_827);
or U1185 (N_1185,In_553,In_1284);
nor U1186 (N_1186,In_1817,N_905);
nor U1187 (N_1187,N_12,N_695);
nand U1188 (N_1188,N_693,In_587);
nand U1189 (N_1189,N_164,N_442);
and U1190 (N_1190,N_872,N_893);
nor U1191 (N_1191,N_989,N_512);
or U1192 (N_1192,N_558,N_664);
or U1193 (N_1193,In_1498,N_890);
nor U1194 (N_1194,In_112,N_875);
nand U1195 (N_1195,In_1614,N_616);
nand U1196 (N_1196,N_902,In_784);
xor U1197 (N_1197,N_464,In_1048);
nor U1198 (N_1198,N_621,N_87);
or U1199 (N_1199,In_1823,N_756);
or U1200 (N_1200,In_1349,N_794);
nor U1201 (N_1201,N_777,N_525);
and U1202 (N_1202,N_938,In_1429);
xor U1203 (N_1203,N_474,N_675);
and U1204 (N_1204,N_889,In_1908);
nor U1205 (N_1205,In_943,In_1447);
or U1206 (N_1206,In_1029,In_1703);
or U1207 (N_1207,N_771,N_816);
and U1208 (N_1208,In_1828,N_560);
xnor U1209 (N_1209,N_588,In_1470);
nand U1210 (N_1210,In_1615,N_564);
nor U1211 (N_1211,N_762,N_605);
nand U1212 (N_1212,N_766,N_703);
xor U1213 (N_1213,N_533,N_604);
or U1214 (N_1214,N_283,In_32);
nand U1215 (N_1215,In_1936,In_174);
nor U1216 (N_1216,In_380,N_836);
xnor U1217 (N_1217,In_1040,In_193);
xnor U1218 (N_1218,N_580,In_1568);
and U1219 (N_1219,N_163,In_421);
or U1220 (N_1220,N_259,N_254);
nand U1221 (N_1221,In_732,In_1320);
or U1222 (N_1222,In_546,In_504);
nand U1223 (N_1223,N_944,N_20);
and U1224 (N_1224,N_392,In_1416);
or U1225 (N_1225,N_523,N_428);
xor U1226 (N_1226,N_714,N_645);
xor U1227 (N_1227,N_205,N_567);
and U1228 (N_1228,In_857,N_43);
xnor U1229 (N_1229,N_100,In_743);
or U1230 (N_1230,N_954,N_915);
nand U1231 (N_1231,N_31,N_950);
and U1232 (N_1232,In_1225,In_1220);
or U1233 (N_1233,N_965,In_1774);
nor U1234 (N_1234,N_975,N_13);
nor U1235 (N_1235,In_1138,In_653);
or U1236 (N_1236,N_268,In_855);
or U1237 (N_1237,In_1954,N_967);
and U1238 (N_1238,N_445,N_745);
and U1239 (N_1239,In_1298,N_104);
xor U1240 (N_1240,N_821,In_952);
xnor U1241 (N_1241,In_591,In_594);
and U1242 (N_1242,N_571,N_948);
and U1243 (N_1243,In_1827,N_550);
or U1244 (N_1244,N_251,N_990);
or U1245 (N_1245,N_943,N_855);
and U1246 (N_1246,In_5,N_635);
xnor U1247 (N_1247,N_46,In_186);
or U1248 (N_1248,N_630,In_21);
and U1249 (N_1249,N_857,N_335);
and U1250 (N_1250,N_654,N_576);
or U1251 (N_1251,N_726,N_928);
nor U1252 (N_1252,In_1696,N_846);
nand U1253 (N_1253,N_994,In_1173);
xor U1254 (N_1254,N_972,N_708);
and U1255 (N_1255,N_456,N_790);
or U1256 (N_1256,N_752,N_109);
xor U1257 (N_1257,N_998,N_733);
nand U1258 (N_1258,N_467,In_1063);
nand U1259 (N_1259,N_810,In_1054);
and U1260 (N_1260,N_538,N_956);
and U1261 (N_1261,N_573,In_1891);
nor U1262 (N_1262,N_680,In_1415);
nand U1263 (N_1263,N_736,In_144);
or U1264 (N_1264,In_1441,N_178);
nor U1265 (N_1265,N_460,In_1156);
nor U1266 (N_1266,N_67,N_612);
or U1267 (N_1267,N_772,N_393);
nor U1268 (N_1268,In_816,In_754);
and U1269 (N_1269,N_150,N_676);
nand U1270 (N_1270,In_1669,In_615);
or U1271 (N_1271,N_812,N_824);
nand U1272 (N_1272,In_1333,In_1226);
or U1273 (N_1273,In_938,N_923);
or U1274 (N_1274,N_125,In_1564);
and U1275 (N_1275,In_891,In_1982);
and U1276 (N_1276,N_718,N_882);
or U1277 (N_1277,N_856,N_858);
nor U1278 (N_1278,N_222,In_1253);
and U1279 (N_1279,In_1856,N_541);
nor U1280 (N_1280,N_955,N_628);
or U1281 (N_1281,N_181,In_1230);
nor U1282 (N_1282,N_537,N_278);
or U1283 (N_1283,N_536,N_228);
nor U1284 (N_1284,N_723,N_161);
and U1285 (N_1285,In_1860,N_644);
or U1286 (N_1286,N_908,In_1316);
and U1287 (N_1287,In_1780,N_983);
xnor U1288 (N_1288,N_509,In_1458);
xnor U1289 (N_1289,In_44,N_269);
xor U1290 (N_1290,N_663,N_618);
xor U1291 (N_1291,In_1070,N_851);
xnor U1292 (N_1292,N_350,In_1025);
xor U1293 (N_1293,In_1937,In_1625);
xnor U1294 (N_1294,N_747,N_757);
and U1295 (N_1295,In_940,N_871);
nor U1296 (N_1296,N_894,N_316);
or U1297 (N_1297,In_1997,N_895);
and U1298 (N_1298,N_865,N_788);
and U1299 (N_1299,N_522,N_848);
or U1300 (N_1300,In_1086,N_231);
nor U1301 (N_1301,N_911,N_732);
and U1302 (N_1302,In_588,N_276);
xor U1303 (N_1303,In_1605,N_942);
and U1304 (N_1304,N_946,In_1057);
or U1305 (N_1305,In_275,N_562);
or U1306 (N_1306,N_678,N_698);
nor U1307 (N_1307,In_1453,N_735);
xnor U1308 (N_1308,N_619,N_624);
or U1309 (N_1309,N_578,N_50);
and U1310 (N_1310,N_795,N_763);
and U1311 (N_1311,N_457,In_797);
or U1312 (N_1312,N_806,In_945);
xnor U1313 (N_1313,N_913,N_832);
xor U1314 (N_1314,N_174,N_531);
nor U1315 (N_1315,N_623,N_937);
nand U1316 (N_1316,In_1122,N_874);
and U1317 (N_1317,N_782,N_371);
nand U1318 (N_1318,N_199,In_877);
or U1319 (N_1319,N_789,N_843);
or U1320 (N_1320,N_864,N_730);
xor U1321 (N_1321,In_842,In_762);
and U1322 (N_1322,N_982,N_551);
and U1323 (N_1323,N_734,N_62);
xor U1324 (N_1324,In_586,N_945);
xor U1325 (N_1325,In_785,N_737);
nand U1326 (N_1326,N_559,N_590);
nor U1327 (N_1327,In_1876,N_89);
nor U1328 (N_1328,N_815,N_897);
and U1329 (N_1329,N_684,N_614);
nand U1330 (N_1330,N_683,N_561);
and U1331 (N_1331,N_850,N_501);
nand U1332 (N_1332,In_840,In_1505);
or U1333 (N_1333,In_616,N_540);
and U1334 (N_1334,In_67,In_570);
and U1335 (N_1335,N_742,In_994);
or U1336 (N_1336,In_687,N_854);
or U1337 (N_1337,N_779,N_716);
and U1338 (N_1338,N_885,N_511);
nand U1339 (N_1339,In_1514,N_962);
nor U1340 (N_1340,N_830,In_1626);
nand U1341 (N_1341,N_157,N_528);
xor U1342 (N_1342,In_1003,In_658);
and U1343 (N_1343,N_987,N_721);
nor U1344 (N_1344,In_859,N_887);
and U1345 (N_1345,N_58,N_220);
or U1346 (N_1346,N_796,N_892);
or U1347 (N_1347,N_353,N_7);
xor U1348 (N_1348,N_506,N_81);
xnor U1349 (N_1349,N_744,In_800);
and U1350 (N_1350,N_743,N_907);
or U1351 (N_1351,In_984,N_640);
xnor U1352 (N_1352,N_884,N_799);
and U1353 (N_1353,In_1434,N_687);
xnor U1354 (N_1354,N_920,N_859);
and U1355 (N_1355,N_329,N_358);
and U1356 (N_1356,N_9,In_839);
nor U1357 (N_1357,N_277,N_566);
and U1358 (N_1358,In_625,In_497);
or U1359 (N_1359,N_845,In_294);
or U1360 (N_1360,N_959,In_1883);
xnor U1361 (N_1361,In_1943,N_933);
or U1362 (N_1362,N_891,In_1418);
xor U1363 (N_1363,N_265,N_674);
or U1364 (N_1364,N_515,N_992);
xnor U1365 (N_1365,N_879,N_819);
or U1366 (N_1366,N_805,N_435);
nor U1367 (N_1367,N_99,N_934);
or U1368 (N_1368,N_595,N_741);
and U1369 (N_1369,N_249,In_1838);
nor U1370 (N_1370,N_957,N_750);
and U1371 (N_1371,N_470,N_652);
and U1372 (N_1372,In_1904,N_526);
or U1373 (N_1373,N_208,N_554);
or U1374 (N_1374,In_1699,In_1200);
xor U1375 (N_1375,N_287,In_1413);
or U1376 (N_1376,In_1401,N_918);
and U1377 (N_1377,N_719,N_545);
nor U1378 (N_1378,In_289,In_172);
and U1379 (N_1379,N_599,In_1414);
nor U1380 (N_1380,In_481,In_1556);
and U1381 (N_1381,N_831,N_904);
nand U1382 (N_1382,N_260,N_597);
xor U1383 (N_1383,N_642,N_903);
or U1384 (N_1384,N_818,N_909);
or U1385 (N_1385,N_749,N_713);
xnor U1386 (N_1386,In_1492,N_720);
and U1387 (N_1387,In_610,N_973);
or U1388 (N_1388,N_530,N_209);
and U1389 (N_1389,N_840,N_970);
nand U1390 (N_1390,N_346,In_718);
and U1391 (N_1391,N_759,In_775);
or U1392 (N_1392,N_696,N_4);
xor U1393 (N_1393,N_147,N_504);
nor U1394 (N_1394,In_1197,In_868);
xor U1395 (N_1395,N_775,In_1665);
and U1396 (N_1396,N_672,N_991);
xnor U1397 (N_1397,In_1812,In_48);
or U1398 (N_1398,N_751,N_421);
and U1399 (N_1399,In_461,N_896);
xor U1400 (N_1400,N_583,N_264);
nand U1401 (N_1401,In_1671,N_686);
or U1402 (N_1402,N_916,N_697);
xnor U1403 (N_1403,N_717,N_853);
or U1404 (N_1404,N_24,N_814);
nor U1405 (N_1405,In_1378,In_959);
or U1406 (N_1406,N_639,In_1125);
and U1407 (N_1407,In_179,N_931);
or U1408 (N_1408,N_880,N_802);
nand U1409 (N_1409,In_149,In_371);
xnor U1410 (N_1410,N_138,In_1923);
xor U1411 (N_1411,N_636,In_597);
nand U1412 (N_1412,N_288,N_866);
and U1413 (N_1413,N_503,N_761);
and U1414 (N_1414,N_380,N_646);
nand U1415 (N_1415,N_552,N_877);
nor U1416 (N_1416,N_261,N_629);
nor U1417 (N_1417,N_490,In_1430);
or U1418 (N_1418,N_662,N_774);
or U1419 (N_1419,N_811,N_711);
and U1420 (N_1420,N_728,N_127);
xor U1421 (N_1421,N_201,In_383);
and U1422 (N_1422,N_776,In_491);
nor U1423 (N_1423,N_28,In_244);
or U1424 (N_1424,In_1323,N_932);
or U1425 (N_1425,N_527,In_486);
or U1426 (N_1426,N_724,N_953);
nand U1427 (N_1427,In_817,N_842);
and U1428 (N_1428,N_607,In_1266);
nor U1429 (N_1429,N_626,In_1238);
or U1430 (N_1430,N_839,N_521);
and U1431 (N_1431,In_1059,In_873);
nand U1432 (N_1432,N_513,In_1913);
and U1433 (N_1433,N_301,N_941);
nand U1434 (N_1434,N_633,N_271);
nand U1435 (N_1435,N_715,In_203);
xnor U1436 (N_1436,N_976,In_479);
xor U1437 (N_1437,N_609,In_875);
nand U1438 (N_1438,In_1952,N_25);
xnor U1439 (N_1439,N_135,N_936);
nand U1440 (N_1440,In_1509,N_940);
nor U1441 (N_1441,In_130,In_1362);
nor U1442 (N_1442,N_656,N_971);
or U1443 (N_1443,In_1880,N_367);
and U1444 (N_1444,N_130,N_984);
xnor U1445 (N_1445,N_577,In_1176);
xor U1446 (N_1446,N_914,N_921);
xnor U1447 (N_1447,N_869,N_270);
nand U1448 (N_1448,N_667,N_939);
or U1449 (N_1449,N_66,N_568);
nand U1450 (N_1450,In_1618,N_906);
and U1451 (N_1451,N_366,In_363);
and U1452 (N_1452,N_701,N_539);
and U1453 (N_1453,N_969,In_804);
nand U1454 (N_1454,N_137,N_706);
nor U1455 (N_1455,N_760,In_341);
xor U1456 (N_1456,N_801,N_452);
nand U1457 (N_1457,In_1109,In_1146);
and U1458 (N_1458,In_758,In_641);
or U1459 (N_1459,In_330,In_248);
or U1460 (N_1460,N_532,In_1723);
or U1461 (N_1461,In_340,N_765);
nor U1462 (N_1462,In_702,N_951);
or U1463 (N_1463,In_1163,In_439);
xnor U1464 (N_1464,N_256,N_968);
nand U1465 (N_1465,N_924,N_985);
nand U1466 (N_1466,N_919,N_709);
nor U1467 (N_1467,In_208,In_463);
or U1468 (N_1468,In_1233,In_1657);
and U1469 (N_1469,N_657,N_952);
and U1470 (N_1470,N_601,In_1597);
xor U1471 (N_1471,N_239,N_516);
and U1472 (N_1472,In_209,N_822);
nor U1473 (N_1473,In_143,N_534);
and U1474 (N_1474,N_651,In_1328);
or U1475 (N_1475,N_883,N_587);
or U1476 (N_1476,N_758,N_797);
or U1477 (N_1477,N_988,N_210);
nor U1478 (N_1478,N_542,In_413);
nand U1479 (N_1479,N_833,N_773);
nand U1480 (N_1480,N_925,N_863);
nand U1481 (N_1481,In_1461,N_484);
xor U1482 (N_1482,In_8,N_582);
xnor U1483 (N_1483,N_700,In_1754);
nand U1484 (N_1484,N_557,N_746);
or U1485 (N_1485,N_901,In_1852);
xnor U1486 (N_1486,In_523,N_849);
nor U1487 (N_1487,In_1347,N_293);
nor U1488 (N_1488,In_109,N_995);
or U1489 (N_1489,In_692,N_508);
xnor U1490 (N_1490,N_620,In_1136);
and U1491 (N_1491,N_669,N_798);
or U1492 (N_1492,N_769,N_986);
xnor U1493 (N_1493,In_296,N_886);
and U1494 (N_1494,N_673,N_572);
and U1495 (N_1495,N_546,N_878);
and U1496 (N_1496,N_602,N_974);
or U1497 (N_1497,N_930,In_387);
nand U1498 (N_1498,N_555,N_579);
xor U1499 (N_1499,N_488,N_841);
nand U1500 (N_1500,N_1041,N_1304);
and U1501 (N_1501,N_1019,N_1440);
nand U1502 (N_1502,N_1089,N_1322);
or U1503 (N_1503,N_1005,N_1119);
nand U1504 (N_1504,N_1441,N_1141);
nor U1505 (N_1505,N_1299,N_1284);
nor U1506 (N_1506,N_1374,N_1061);
and U1507 (N_1507,N_1283,N_1271);
nand U1508 (N_1508,N_1031,N_1050);
nor U1509 (N_1509,N_1082,N_1477);
nand U1510 (N_1510,N_1191,N_1045);
or U1511 (N_1511,N_1242,N_1454);
nor U1512 (N_1512,N_1189,N_1091);
and U1513 (N_1513,N_1260,N_1408);
or U1514 (N_1514,N_1121,N_1088);
and U1515 (N_1515,N_1334,N_1330);
or U1516 (N_1516,N_1067,N_1449);
nor U1517 (N_1517,N_1007,N_1390);
xnor U1518 (N_1518,N_1318,N_1154);
xnor U1519 (N_1519,N_1377,N_1384);
xor U1520 (N_1520,N_1354,N_1149);
xnor U1521 (N_1521,N_1020,N_1338);
nor U1522 (N_1522,N_1383,N_1275);
xnor U1523 (N_1523,N_1410,N_1074);
xnor U1524 (N_1524,N_1348,N_1225);
xor U1525 (N_1525,N_1496,N_1286);
and U1526 (N_1526,N_1052,N_1212);
or U1527 (N_1527,N_1493,N_1169);
nand U1528 (N_1528,N_1195,N_1240);
nand U1529 (N_1529,N_1439,N_1073);
or U1530 (N_1530,N_1300,N_1126);
nand U1531 (N_1531,N_1401,N_1103);
or U1532 (N_1532,N_1112,N_1219);
nor U1533 (N_1533,N_1499,N_1349);
xnor U1534 (N_1534,N_1210,N_1062);
and U1535 (N_1535,N_1267,N_1072);
or U1536 (N_1536,N_1016,N_1035);
or U1537 (N_1537,N_1162,N_1261);
xnor U1538 (N_1538,N_1167,N_1340);
and U1539 (N_1539,N_1176,N_1312);
nor U1540 (N_1540,N_1385,N_1458);
nand U1541 (N_1541,N_1053,N_1131);
or U1542 (N_1542,N_1382,N_1178);
or U1543 (N_1543,N_1469,N_1209);
xor U1544 (N_1544,N_1317,N_1185);
and U1545 (N_1545,N_1277,N_1264);
xor U1546 (N_1546,N_1353,N_1307);
and U1547 (N_1547,N_1258,N_1319);
nor U1548 (N_1548,N_1190,N_1151);
xor U1549 (N_1549,N_1339,N_1101);
xnor U1550 (N_1550,N_1234,N_1237);
xor U1551 (N_1551,N_1206,N_1485);
xnor U1552 (N_1552,N_1259,N_1280);
and U1553 (N_1553,N_1389,N_1118);
xor U1554 (N_1554,N_1093,N_1415);
and U1555 (N_1555,N_1297,N_1044);
and U1556 (N_1556,N_1180,N_1294);
nand U1557 (N_1557,N_1246,N_1253);
or U1558 (N_1558,N_1243,N_1222);
xor U1559 (N_1559,N_1163,N_1314);
and U1560 (N_1560,N_1305,N_1023);
nor U1561 (N_1561,N_1282,N_1398);
or U1562 (N_1562,N_1160,N_1328);
nor U1563 (N_1563,N_1065,N_1288);
nor U1564 (N_1564,N_1100,N_1129);
and U1565 (N_1565,N_1086,N_1452);
or U1566 (N_1566,N_1059,N_1120);
xor U1567 (N_1567,N_1342,N_1373);
xnor U1568 (N_1568,N_1012,N_1343);
and U1569 (N_1569,N_1022,N_1245);
xnor U1570 (N_1570,N_1177,N_1140);
nand U1571 (N_1571,N_1227,N_1236);
nand U1572 (N_1572,N_1473,N_1098);
and U1573 (N_1573,N_1250,N_1173);
xnor U1574 (N_1574,N_1064,N_1460);
xnor U1575 (N_1575,N_1087,N_1308);
or U1576 (N_1576,N_1431,N_1158);
or U1577 (N_1577,N_1428,N_1376);
nand U1578 (N_1578,N_1347,N_1432);
and U1579 (N_1579,N_1226,N_1329);
and U1580 (N_1580,N_1276,N_1287);
nor U1581 (N_1581,N_1302,N_1278);
and U1582 (N_1582,N_1381,N_1488);
and U1583 (N_1583,N_1028,N_1213);
nand U1584 (N_1584,N_1116,N_1256);
nor U1585 (N_1585,N_1155,N_1033);
xnor U1586 (N_1586,N_1010,N_1337);
nor U1587 (N_1587,N_1198,N_1069);
and U1588 (N_1588,N_1133,N_1462);
or U1589 (N_1589,N_1139,N_1203);
or U1590 (N_1590,N_1375,N_1196);
nor U1591 (N_1591,N_1459,N_1193);
or U1592 (N_1592,N_1036,N_1427);
and U1593 (N_1593,N_1168,N_1057);
nor U1594 (N_1594,N_1128,N_1405);
nand U1595 (N_1595,N_1156,N_1388);
and U1596 (N_1596,N_1221,N_1336);
and U1597 (N_1597,N_1181,N_1251);
xnor U1598 (N_1598,N_1268,N_1455);
nand U1599 (N_1599,N_1172,N_1111);
nor U1600 (N_1600,N_1105,N_1331);
and U1601 (N_1601,N_1184,N_1451);
and U1602 (N_1602,N_1450,N_1396);
xor U1603 (N_1603,N_1363,N_1144);
nand U1604 (N_1604,N_1060,N_1255);
xnor U1605 (N_1605,N_1147,N_1403);
xor U1606 (N_1606,N_1194,N_1241);
xnor U1607 (N_1607,N_1335,N_1166);
nor U1608 (N_1608,N_1372,N_1456);
xor U1609 (N_1609,N_1368,N_1444);
nor U1610 (N_1610,N_1358,N_1137);
nand U1611 (N_1611,N_1402,N_1081);
and U1612 (N_1612,N_1084,N_1487);
nor U1613 (N_1613,N_1003,N_1179);
xor U1614 (N_1614,N_1266,N_1494);
xnor U1615 (N_1615,N_1008,N_1365);
nor U1616 (N_1616,N_1327,N_1114);
xor U1617 (N_1617,N_1110,N_1483);
or U1618 (N_1618,N_1395,N_1482);
nand U1619 (N_1619,N_1068,N_1433);
or U1620 (N_1620,N_1438,N_1475);
xor U1621 (N_1621,N_1479,N_1490);
and U1622 (N_1622,N_1182,N_1341);
nor U1623 (N_1623,N_1040,N_1159);
or U1624 (N_1624,N_1076,N_1257);
and U1625 (N_1625,N_1421,N_1400);
nor U1626 (N_1626,N_1097,N_1006);
xor U1627 (N_1627,N_1208,N_1351);
or U1628 (N_1628,N_1071,N_1362);
or U1629 (N_1629,N_1371,N_1078);
nor U1630 (N_1630,N_1369,N_1292);
xnor U1631 (N_1631,N_1229,N_1332);
nor U1632 (N_1632,N_1143,N_1430);
or U1633 (N_1633,N_1115,N_1484);
or U1634 (N_1634,N_1476,N_1090);
xnor U1635 (N_1635,N_1051,N_1435);
xor U1636 (N_1636,N_1000,N_1011);
and U1637 (N_1637,N_1047,N_1218);
and U1638 (N_1638,N_1165,N_1325);
nor U1639 (N_1639,N_1094,N_1379);
nor U1640 (N_1640,N_1175,N_1254);
nand U1641 (N_1641,N_1009,N_1345);
nor U1642 (N_1642,N_1146,N_1446);
xor U1643 (N_1643,N_1448,N_1124);
nand U1644 (N_1644,N_1027,N_1148);
nor U1645 (N_1645,N_1070,N_1085);
nand U1646 (N_1646,N_1130,N_1002);
xnor U1647 (N_1647,N_1316,N_1406);
and U1648 (N_1648,N_1486,N_1333);
nor U1649 (N_1649,N_1230,N_1192);
and U1650 (N_1650,N_1214,N_1471);
nand U1651 (N_1651,N_1021,N_1056);
nor U1652 (N_1652,N_1443,N_1004);
xor U1653 (N_1653,N_1232,N_1049);
nor U1654 (N_1654,N_1491,N_1272);
nand U1655 (N_1655,N_1216,N_1295);
or U1656 (N_1656,N_1407,N_1411);
xor U1657 (N_1657,N_1249,N_1058);
xor U1658 (N_1658,N_1024,N_1472);
nor U1659 (N_1659,N_1030,N_1387);
and U1660 (N_1660,N_1346,N_1252);
xor U1661 (N_1661,N_1066,N_1039);
nor U1662 (N_1662,N_1293,N_1157);
nand U1663 (N_1663,N_1095,N_1001);
nand U1664 (N_1664,N_1138,N_1248);
xnor U1665 (N_1665,N_1220,N_1313);
nand U1666 (N_1666,N_1127,N_1239);
or U1667 (N_1667,N_1017,N_1034);
or U1668 (N_1668,N_1352,N_1026);
or U1669 (N_1669,N_1122,N_1392);
nor U1670 (N_1670,N_1055,N_1359);
xor U1671 (N_1671,N_1291,N_1018);
and U1672 (N_1672,N_1200,N_1048);
or U1673 (N_1673,N_1397,N_1145);
xnor U1674 (N_1674,N_1037,N_1104);
nor U1675 (N_1675,N_1077,N_1478);
nand U1676 (N_1676,N_1289,N_1075);
nand U1677 (N_1677,N_1270,N_1262);
nor U1678 (N_1678,N_1422,N_1466);
or U1679 (N_1679,N_1215,N_1301);
nand U1680 (N_1680,N_1366,N_1391);
or U1681 (N_1681,N_1107,N_1153);
or U1682 (N_1682,N_1425,N_1265);
xor U1683 (N_1683,N_1386,N_1350);
nor U1684 (N_1684,N_1360,N_1187);
nand U1685 (N_1685,N_1470,N_1063);
or U1686 (N_1686,N_1233,N_1323);
nor U1687 (N_1687,N_1205,N_1436);
xnor U1688 (N_1688,N_1303,N_1412);
nand U1689 (N_1689,N_1281,N_1224);
and U1690 (N_1690,N_1054,N_1361);
nor U1691 (N_1691,N_1013,N_1269);
or U1692 (N_1692,N_1099,N_1150);
or U1693 (N_1693,N_1217,N_1461);
nor U1694 (N_1694,N_1419,N_1378);
nand U1695 (N_1695,N_1492,N_1201);
and U1696 (N_1696,N_1102,N_1474);
and U1697 (N_1697,N_1467,N_1424);
and U1698 (N_1698,N_1413,N_1279);
and U1699 (N_1699,N_1274,N_1238);
or U1700 (N_1700,N_1025,N_1247);
and U1701 (N_1701,N_1235,N_1092);
nand U1702 (N_1702,N_1465,N_1046);
and U1703 (N_1703,N_1426,N_1109);
or U1704 (N_1704,N_1014,N_1186);
nand U1705 (N_1705,N_1170,N_1480);
and U1706 (N_1706,N_1197,N_1263);
nand U1707 (N_1707,N_1481,N_1357);
and U1708 (N_1708,N_1498,N_1453);
and U1709 (N_1709,N_1188,N_1414);
or U1710 (N_1710,N_1029,N_1106);
or U1711 (N_1711,N_1142,N_1315);
and U1712 (N_1712,N_1364,N_1320);
nand U1713 (N_1713,N_1096,N_1290);
xnor U1714 (N_1714,N_1296,N_1306);
xor U1715 (N_1715,N_1298,N_1273);
and U1716 (N_1716,N_1404,N_1211);
and U1717 (N_1717,N_1202,N_1457);
and U1718 (N_1718,N_1409,N_1309);
and U1719 (N_1719,N_1416,N_1042);
xnor U1720 (N_1720,N_1032,N_1370);
nor U1721 (N_1721,N_1135,N_1420);
and U1722 (N_1722,N_1324,N_1463);
nor U1723 (N_1723,N_1489,N_1117);
xnor U1724 (N_1724,N_1495,N_1380);
nand U1725 (N_1725,N_1321,N_1174);
and U1726 (N_1726,N_1079,N_1134);
and U1727 (N_1727,N_1417,N_1123);
nand U1728 (N_1728,N_1231,N_1356);
xor U1729 (N_1729,N_1399,N_1464);
nor U1730 (N_1730,N_1164,N_1355);
and U1731 (N_1731,N_1497,N_1429);
nand U1732 (N_1732,N_1038,N_1108);
nor U1733 (N_1733,N_1199,N_1113);
or U1734 (N_1734,N_1394,N_1311);
and U1735 (N_1735,N_1125,N_1468);
xnor U1736 (N_1736,N_1204,N_1437);
or U1737 (N_1737,N_1161,N_1171);
or U1738 (N_1738,N_1447,N_1244);
and U1739 (N_1739,N_1434,N_1043);
xor U1740 (N_1740,N_1344,N_1183);
xor U1741 (N_1741,N_1310,N_1393);
nor U1742 (N_1742,N_1423,N_1228);
or U1743 (N_1743,N_1285,N_1083);
xor U1744 (N_1744,N_1207,N_1442);
and U1745 (N_1745,N_1015,N_1367);
and U1746 (N_1746,N_1445,N_1326);
xnor U1747 (N_1747,N_1223,N_1080);
or U1748 (N_1748,N_1132,N_1418);
nor U1749 (N_1749,N_1136,N_1152);
xor U1750 (N_1750,N_1499,N_1397);
and U1751 (N_1751,N_1416,N_1105);
or U1752 (N_1752,N_1281,N_1366);
and U1753 (N_1753,N_1446,N_1118);
xor U1754 (N_1754,N_1309,N_1382);
nand U1755 (N_1755,N_1280,N_1154);
and U1756 (N_1756,N_1061,N_1469);
nor U1757 (N_1757,N_1041,N_1161);
nand U1758 (N_1758,N_1065,N_1392);
nand U1759 (N_1759,N_1130,N_1447);
nand U1760 (N_1760,N_1469,N_1300);
nor U1761 (N_1761,N_1056,N_1403);
nand U1762 (N_1762,N_1155,N_1437);
nor U1763 (N_1763,N_1141,N_1056);
nand U1764 (N_1764,N_1083,N_1120);
xnor U1765 (N_1765,N_1155,N_1020);
or U1766 (N_1766,N_1466,N_1454);
or U1767 (N_1767,N_1483,N_1133);
or U1768 (N_1768,N_1443,N_1094);
nand U1769 (N_1769,N_1025,N_1334);
nand U1770 (N_1770,N_1362,N_1022);
and U1771 (N_1771,N_1473,N_1466);
nor U1772 (N_1772,N_1468,N_1415);
nor U1773 (N_1773,N_1243,N_1250);
or U1774 (N_1774,N_1342,N_1413);
xor U1775 (N_1775,N_1212,N_1254);
nor U1776 (N_1776,N_1209,N_1152);
and U1777 (N_1777,N_1467,N_1292);
or U1778 (N_1778,N_1283,N_1335);
or U1779 (N_1779,N_1246,N_1318);
and U1780 (N_1780,N_1396,N_1419);
nand U1781 (N_1781,N_1359,N_1073);
and U1782 (N_1782,N_1463,N_1013);
xor U1783 (N_1783,N_1219,N_1021);
xnor U1784 (N_1784,N_1422,N_1459);
xor U1785 (N_1785,N_1418,N_1259);
and U1786 (N_1786,N_1094,N_1046);
nand U1787 (N_1787,N_1330,N_1286);
nand U1788 (N_1788,N_1399,N_1442);
and U1789 (N_1789,N_1004,N_1054);
and U1790 (N_1790,N_1450,N_1194);
or U1791 (N_1791,N_1201,N_1309);
or U1792 (N_1792,N_1453,N_1212);
nand U1793 (N_1793,N_1317,N_1340);
nand U1794 (N_1794,N_1178,N_1113);
xor U1795 (N_1795,N_1352,N_1025);
nor U1796 (N_1796,N_1235,N_1312);
nor U1797 (N_1797,N_1258,N_1374);
xnor U1798 (N_1798,N_1440,N_1472);
nand U1799 (N_1799,N_1350,N_1318);
or U1800 (N_1800,N_1191,N_1227);
nor U1801 (N_1801,N_1328,N_1112);
or U1802 (N_1802,N_1167,N_1201);
or U1803 (N_1803,N_1247,N_1178);
nand U1804 (N_1804,N_1086,N_1422);
or U1805 (N_1805,N_1372,N_1279);
nand U1806 (N_1806,N_1465,N_1034);
nor U1807 (N_1807,N_1117,N_1306);
nand U1808 (N_1808,N_1484,N_1308);
nand U1809 (N_1809,N_1156,N_1453);
or U1810 (N_1810,N_1266,N_1480);
nor U1811 (N_1811,N_1267,N_1148);
or U1812 (N_1812,N_1377,N_1481);
or U1813 (N_1813,N_1020,N_1449);
nand U1814 (N_1814,N_1420,N_1097);
nand U1815 (N_1815,N_1249,N_1021);
nor U1816 (N_1816,N_1051,N_1333);
and U1817 (N_1817,N_1001,N_1420);
xnor U1818 (N_1818,N_1017,N_1005);
nand U1819 (N_1819,N_1010,N_1377);
nor U1820 (N_1820,N_1471,N_1450);
or U1821 (N_1821,N_1401,N_1340);
nand U1822 (N_1822,N_1400,N_1283);
or U1823 (N_1823,N_1018,N_1097);
and U1824 (N_1824,N_1422,N_1300);
nand U1825 (N_1825,N_1042,N_1351);
nor U1826 (N_1826,N_1087,N_1100);
and U1827 (N_1827,N_1308,N_1333);
or U1828 (N_1828,N_1363,N_1134);
and U1829 (N_1829,N_1147,N_1393);
nand U1830 (N_1830,N_1067,N_1485);
xnor U1831 (N_1831,N_1369,N_1278);
nand U1832 (N_1832,N_1116,N_1176);
xnor U1833 (N_1833,N_1014,N_1361);
nor U1834 (N_1834,N_1144,N_1083);
nand U1835 (N_1835,N_1239,N_1484);
xor U1836 (N_1836,N_1219,N_1124);
or U1837 (N_1837,N_1419,N_1332);
or U1838 (N_1838,N_1321,N_1102);
xnor U1839 (N_1839,N_1183,N_1227);
or U1840 (N_1840,N_1246,N_1325);
nor U1841 (N_1841,N_1297,N_1377);
and U1842 (N_1842,N_1247,N_1407);
xnor U1843 (N_1843,N_1212,N_1067);
xnor U1844 (N_1844,N_1236,N_1420);
nand U1845 (N_1845,N_1140,N_1132);
nand U1846 (N_1846,N_1104,N_1058);
or U1847 (N_1847,N_1161,N_1319);
and U1848 (N_1848,N_1445,N_1302);
and U1849 (N_1849,N_1222,N_1014);
nor U1850 (N_1850,N_1134,N_1140);
or U1851 (N_1851,N_1213,N_1338);
xnor U1852 (N_1852,N_1027,N_1068);
nand U1853 (N_1853,N_1240,N_1129);
and U1854 (N_1854,N_1071,N_1321);
xnor U1855 (N_1855,N_1393,N_1142);
and U1856 (N_1856,N_1328,N_1415);
and U1857 (N_1857,N_1411,N_1480);
and U1858 (N_1858,N_1307,N_1216);
or U1859 (N_1859,N_1430,N_1450);
or U1860 (N_1860,N_1370,N_1441);
and U1861 (N_1861,N_1219,N_1068);
xnor U1862 (N_1862,N_1444,N_1191);
xnor U1863 (N_1863,N_1374,N_1049);
nand U1864 (N_1864,N_1469,N_1033);
nor U1865 (N_1865,N_1483,N_1016);
nand U1866 (N_1866,N_1159,N_1262);
nand U1867 (N_1867,N_1232,N_1383);
or U1868 (N_1868,N_1068,N_1333);
nand U1869 (N_1869,N_1494,N_1108);
nor U1870 (N_1870,N_1215,N_1225);
nor U1871 (N_1871,N_1281,N_1054);
nand U1872 (N_1872,N_1045,N_1144);
xor U1873 (N_1873,N_1072,N_1420);
xnor U1874 (N_1874,N_1278,N_1276);
nor U1875 (N_1875,N_1304,N_1130);
xor U1876 (N_1876,N_1053,N_1178);
or U1877 (N_1877,N_1295,N_1416);
and U1878 (N_1878,N_1354,N_1126);
or U1879 (N_1879,N_1268,N_1481);
nand U1880 (N_1880,N_1274,N_1023);
xor U1881 (N_1881,N_1411,N_1209);
nand U1882 (N_1882,N_1390,N_1117);
or U1883 (N_1883,N_1236,N_1335);
and U1884 (N_1884,N_1109,N_1051);
and U1885 (N_1885,N_1165,N_1135);
and U1886 (N_1886,N_1025,N_1178);
xor U1887 (N_1887,N_1436,N_1426);
or U1888 (N_1888,N_1056,N_1492);
nor U1889 (N_1889,N_1179,N_1262);
xor U1890 (N_1890,N_1331,N_1365);
xnor U1891 (N_1891,N_1239,N_1057);
or U1892 (N_1892,N_1464,N_1113);
or U1893 (N_1893,N_1437,N_1073);
or U1894 (N_1894,N_1213,N_1379);
nand U1895 (N_1895,N_1423,N_1055);
and U1896 (N_1896,N_1261,N_1474);
nand U1897 (N_1897,N_1440,N_1001);
or U1898 (N_1898,N_1039,N_1400);
xor U1899 (N_1899,N_1428,N_1440);
or U1900 (N_1900,N_1424,N_1465);
nand U1901 (N_1901,N_1159,N_1142);
and U1902 (N_1902,N_1236,N_1389);
nand U1903 (N_1903,N_1402,N_1388);
or U1904 (N_1904,N_1373,N_1437);
nand U1905 (N_1905,N_1417,N_1020);
or U1906 (N_1906,N_1435,N_1031);
or U1907 (N_1907,N_1227,N_1117);
and U1908 (N_1908,N_1054,N_1191);
or U1909 (N_1909,N_1290,N_1315);
nand U1910 (N_1910,N_1059,N_1382);
nand U1911 (N_1911,N_1144,N_1141);
xnor U1912 (N_1912,N_1459,N_1372);
and U1913 (N_1913,N_1109,N_1147);
xor U1914 (N_1914,N_1333,N_1231);
nor U1915 (N_1915,N_1481,N_1334);
nor U1916 (N_1916,N_1344,N_1193);
xor U1917 (N_1917,N_1413,N_1300);
nand U1918 (N_1918,N_1241,N_1021);
or U1919 (N_1919,N_1451,N_1263);
nand U1920 (N_1920,N_1347,N_1158);
nand U1921 (N_1921,N_1240,N_1076);
and U1922 (N_1922,N_1233,N_1455);
nand U1923 (N_1923,N_1100,N_1468);
and U1924 (N_1924,N_1270,N_1263);
or U1925 (N_1925,N_1281,N_1295);
and U1926 (N_1926,N_1275,N_1216);
xnor U1927 (N_1927,N_1435,N_1447);
and U1928 (N_1928,N_1243,N_1020);
xnor U1929 (N_1929,N_1446,N_1046);
xor U1930 (N_1930,N_1300,N_1183);
nor U1931 (N_1931,N_1093,N_1290);
xnor U1932 (N_1932,N_1496,N_1426);
or U1933 (N_1933,N_1088,N_1354);
nand U1934 (N_1934,N_1472,N_1315);
nor U1935 (N_1935,N_1186,N_1482);
and U1936 (N_1936,N_1465,N_1464);
nor U1937 (N_1937,N_1110,N_1477);
nor U1938 (N_1938,N_1388,N_1380);
nand U1939 (N_1939,N_1129,N_1440);
or U1940 (N_1940,N_1366,N_1433);
xnor U1941 (N_1941,N_1151,N_1396);
or U1942 (N_1942,N_1069,N_1351);
xor U1943 (N_1943,N_1155,N_1401);
nand U1944 (N_1944,N_1227,N_1047);
and U1945 (N_1945,N_1183,N_1004);
and U1946 (N_1946,N_1324,N_1453);
nor U1947 (N_1947,N_1291,N_1115);
nor U1948 (N_1948,N_1011,N_1024);
nor U1949 (N_1949,N_1446,N_1301);
nand U1950 (N_1950,N_1078,N_1159);
and U1951 (N_1951,N_1186,N_1125);
nor U1952 (N_1952,N_1369,N_1014);
nand U1953 (N_1953,N_1414,N_1271);
nor U1954 (N_1954,N_1179,N_1471);
or U1955 (N_1955,N_1386,N_1018);
xor U1956 (N_1956,N_1159,N_1212);
nor U1957 (N_1957,N_1210,N_1324);
or U1958 (N_1958,N_1494,N_1203);
or U1959 (N_1959,N_1104,N_1479);
or U1960 (N_1960,N_1032,N_1379);
and U1961 (N_1961,N_1104,N_1177);
nand U1962 (N_1962,N_1085,N_1438);
nand U1963 (N_1963,N_1404,N_1179);
nand U1964 (N_1964,N_1417,N_1303);
xor U1965 (N_1965,N_1484,N_1009);
nand U1966 (N_1966,N_1189,N_1458);
nor U1967 (N_1967,N_1394,N_1454);
nand U1968 (N_1968,N_1214,N_1337);
or U1969 (N_1969,N_1317,N_1231);
and U1970 (N_1970,N_1333,N_1182);
xnor U1971 (N_1971,N_1213,N_1308);
or U1972 (N_1972,N_1043,N_1050);
xnor U1973 (N_1973,N_1234,N_1151);
nand U1974 (N_1974,N_1367,N_1369);
or U1975 (N_1975,N_1006,N_1297);
or U1976 (N_1976,N_1365,N_1156);
nor U1977 (N_1977,N_1102,N_1388);
and U1978 (N_1978,N_1332,N_1271);
and U1979 (N_1979,N_1114,N_1021);
xnor U1980 (N_1980,N_1060,N_1142);
and U1981 (N_1981,N_1031,N_1188);
or U1982 (N_1982,N_1168,N_1493);
and U1983 (N_1983,N_1225,N_1389);
or U1984 (N_1984,N_1451,N_1176);
nand U1985 (N_1985,N_1304,N_1206);
xnor U1986 (N_1986,N_1164,N_1082);
nand U1987 (N_1987,N_1010,N_1090);
and U1988 (N_1988,N_1198,N_1279);
nor U1989 (N_1989,N_1004,N_1404);
or U1990 (N_1990,N_1212,N_1102);
and U1991 (N_1991,N_1062,N_1409);
xnor U1992 (N_1992,N_1298,N_1336);
nor U1993 (N_1993,N_1397,N_1061);
nor U1994 (N_1994,N_1031,N_1166);
xor U1995 (N_1995,N_1205,N_1208);
xor U1996 (N_1996,N_1493,N_1042);
or U1997 (N_1997,N_1321,N_1293);
nand U1998 (N_1998,N_1482,N_1224);
nor U1999 (N_1999,N_1452,N_1272);
or U2000 (N_2000,N_1937,N_1525);
and U2001 (N_2001,N_1934,N_1931);
or U2002 (N_2002,N_1735,N_1771);
xnor U2003 (N_2003,N_1639,N_1627);
nand U2004 (N_2004,N_1775,N_1523);
nand U2005 (N_2005,N_1812,N_1972);
nor U2006 (N_2006,N_1580,N_1708);
and U2007 (N_2007,N_1923,N_1641);
and U2008 (N_2008,N_1727,N_1784);
nand U2009 (N_2009,N_1891,N_1811);
or U2010 (N_2010,N_1926,N_1630);
xor U2011 (N_2011,N_1834,N_1738);
nand U2012 (N_2012,N_1846,N_1974);
and U2013 (N_2013,N_1616,N_1857);
nand U2014 (N_2014,N_1597,N_1572);
xnor U2015 (N_2015,N_1642,N_1541);
nand U2016 (N_2016,N_1986,N_1569);
or U2017 (N_2017,N_1791,N_1648);
or U2018 (N_2018,N_1793,N_1553);
nand U2019 (N_2019,N_1780,N_1820);
and U2020 (N_2020,N_1538,N_1875);
xnor U2021 (N_2021,N_1958,N_1505);
nor U2022 (N_2022,N_1810,N_1513);
and U2023 (N_2023,N_1506,N_1802);
nor U2024 (N_2024,N_1685,N_1595);
and U2025 (N_2025,N_1831,N_1998);
or U2026 (N_2026,N_1890,N_1660);
or U2027 (N_2027,N_1768,N_1714);
xnor U2028 (N_2028,N_1560,N_1807);
or U2029 (N_2029,N_1544,N_1767);
xor U2030 (N_2030,N_1586,N_1773);
nand U2031 (N_2031,N_1500,N_1960);
xor U2032 (N_2032,N_1678,N_1763);
and U2033 (N_2033,N_1750,N_1501);
nand U2034 (N_2034,N_1528,N_1956);
nor U2035 (N_2035,N_1593,N_1950);
nor U2036 (N_2036,N_1900,N_1969);
nor U2037 (N_2037,N_1838,N_1698);
and U2038 (N_2038,N_1815,N_1935);
and U2039 (N_2039,N_1594,N_1976);
or U2040 (N_2040,N_1650,N_1781);
or U2041 (N_2041,N_1582,N_1795);
or U2042 (N_2042,N_1679,N_1504);
xnor U2043 (N_2043,N_1720,N_1662);
xor U2044 (N_2044,N_1743,N_1529);
and U2045 (N_2045,N_1829,N_1824);
nor U2046 (N_2046,N_1840,N_1634);
xor U2047 (N_2047,N_1654,N_1861);
and U2048 (N_2048,N_1629,N_1516);
nor U2049 (N_2049,N_1539,N_1522);
and U2050 (N_2050,N_1948,N_1806);
nand U2051 (N_2051,N_1941,N_1995);
or U2052 (N_2052,N_1883,N_1870);
and U2053 (N_2053,N_1588,N_1942);
nand U2054 (N_2054,N_1576,N_1696);
nand U2055 (N_2055,N_1723,N_1693);
nor U2056 (N_2056,N_1970,N_1703);
nor U2057 (N_2057,N_1530,N_1961);
nor U2058 (N_2058,N_1589,N_1902);
or U2059 (N_2059,N_1628,N_1725);
nor U2060 (N_2060,N_1520,N_1866);
nand U2061 (N_2061,N_1567,N_1674);
and U2062 (N_2062,N_1579,N_1962);
and U2063 (N_2063,N_1524,N_1746);
nor U2064 (N_2064,N_1638,N_1963);
nand U2065 (N_2065,N_1635,N_1876);
and U2066 (N_2066,N_1692,N_1922);
nor U2067 (N_2067,N_1519,N_1980);
xor U2068 (N_2068,N_1919,N_1514);
nor U2069 (N_2069,N_1645,N_1694);
xnor U2070 (N_2070,N_1571,N_1691);
nand U2071 (N_2071,N_1554,N_1766);
nand U2072 (N_2072,N_1655,N_1837);
or U2073 (N_2073,N_1732,N_1700);
xnor U2074 (N_2074,N_1882,N_1808);
or U2075 (N_2075,N_1885,N_1591);
nand U2076 (N_2076,N_1916,N_1917);
and U2077 (N_2077,N_1796,N_1617);
and U2078 (N_2078,N_1844,N_1804);
nand U2079 (N_2079,N_1841,N_1709);
or U2080 (N_2080,N_1610,N_1813);
nand U2081 (N_2081,N_1669,N_1847);
and U2082 (N_2082,N_1981,N_1545);
xnor U2083 (N_2083,N_1666,N_1581);
or U2084 (N_2084,N_1596,N_1792);
nor U2085 (N_2085,N_1849,N_1702);
and U2086 (N_2086,N_1893,N_1799);
nor U2087 (N_2087,N_1943,N_1656);
or U2088 (N_2088,N_1949,N_1646);
and U2089 (N_2089,N_1858,N_1982);
or U2090 (N_2090,N_1584,N_1542);
nand U2091 (N_2091,N_1764,N_1879);
and U2092 (N_2092,N_1686,N_1748);
xnor U2093 (N_2093,N_1863,N_1770);
nand U2094 (N_2094,N_1653,N_1689);
nand U2095 (N_2095,N_1557,N_1825);
and U2096 (N_2096,N_1772,N_1682);
nand U2097 (N_2097,N_1587,N_1536);
or U2098 (N_2098,N_1774,N_1563);
and U2099 (N_2099,N_1758,N_1985);
xor U2100 (N_2100,N_1631,N_1573);
and U2101 (N_2101,N_1852,N_1845);
xnor U2102 (N_2102,N_1756,N_1918);
nor U2103 (N_2103,N_1622,N_1987);
or U2104 (N_2104,N_1896,N_1869);
and U2105 (N_2105,N_1953,N_1537);
nand U2106 (N_2106,N_1611,N_1790);
and U2107 (N_2107,N_1706,N_1749);
or U2108 (N_2108,N_1512,N_1871);
nand U2109 (N_2109,N_1601,N_1996);
nor U2110 (N_2110,N_1989,N_1559);
and U2111 (N_2111,N_1786,N_1994);
xnor U2112 (N_2112,N_1983,N_1535);
nand U2113 (N_2113,N_1851,N_1533);
xnor U2114 (N_2114,N_1651,N_1930);
xor U2115 (N_2115,N_1877,N_1574);
or U2116 (N_2116,N_1868,N_1924);
xnor U2117 (N_2117,N_1510,N_1992);
nor U2118 (N_2118,N_1633,N_1966);
or U2119 (N_2119,N_1733,N_1640);
xnor U2120 (N_2120,N_1690,N_1867);
and U2121 (N_2121,N_1757,N_1915);
or U2122 (N_2122,N_1687,N_1988);
or U2123 (N_2123,N_1744,N_1908);
nand U2124 (N_2124,N_1839,N_1809);
nor U2125 (N_2125,N_1929,N_1999);
nor U2126 (N_2126,N_1540,N_1776);
or U2127 (N_2127,N_1803,N_1873);
nor U2128 (N_2128,N_1978,N_1644);
xor U2129 (N_2129,N_1859,N_1788);
and U2130 (N_2130,N_1975,N_1620);
xor U2131 (N_2131,N_1719,N_1585);
nand U2132 (N_2132,N_1740,N_1564);
nand U2133 (N_2133,N_1816,N_1798);
or U2134 (N_2134,N_1680,N_1990);
xnor U2135 (N_2135,N_1979,N_1526);
nor U2136 (N_2136,N_1787,N_1637);
nand U2137 (N_2137,N_1657,N_1711);
or U2138 (N_2138,N_1624,N_1911);
or U2139 (N_2139,N_1652,N_1664);
or U2140 (N_2140,N_1614,N_1561);
and U2141 (N_2141,N_1860,N_1936);
nand U2142 (N_2142,N_1818,N_1507);
nand U2143 (N_2143,N_1736,N_1741);
nor U2144 (N_2144,N_1671,N_1668);
nand U2145 (N_2145,N_1894,N_1701);
xnor U2146 (N_2146,N_1546,N_1887);
nor U2147 (N_2147,N_1800,N_1836);
xor U2148 (N_2148,N_1862,N_1921);
nand U2149 (N_2149,N_1991,N_1697);
or U2150 (N_2150,N_1672,N_1801);
or U2151 (N_2151,N_1794,N_1747);
nand U2152 (N_2152,N_1901,N_1707);
xnor U2153 (N_2153,N_1577,N_1613);
or U2154 (N_2154,N_1575,N_1888);
xnor U2155 (N_2155,N_1716,N_1971);
and U2156 (N_2156,N_1612,N_1884);
xor U2157 (N_2157,N_1606,N_1623);
or U2158 (N_2158,N_1517,N_1889);
nor U2159 (N_2159,N_1583,N_1667);
or U2160 (N_2160,N_1615,N_1739);
nor U2161 (N_2161,N_1765,N_1555);
xor U2162 (N_2162,N_1681,N_1608);
xor U2163 (N_2163,N_1604,N_1906);
xnor U2164 (N_2164,N_1592,N_1683);
and U2165 (N_2165,N_1762,N_1932);
nand U2166 (N_2166,N_1705,N_1928);
nor U2167 (N_2167,N_1872,N_1726);
nor U2168 (N_2168,N_1946,N_1895);
nor U2169 (N_2169,N_1552,N_1676);
nand U2170 (N_2170,N_1964,N_1724);
xnor U2171 (N_2171,N_1665,N_1600);
or U2172 (N_2172,N_1827,N_1562);
xor U2173 (N_2173,N_1731,N_1778);
xor U2174 (N_2174,N_1605,N_1625);
nand U2175 (N_2175,N_1789,N_1850);
or U2176 (N_2176,N_1548,N_1854);
nand U2177 (N_2177,N_1933,N_1712);
xnor U2178 (N_2178,N_1502,N_1511);
and U2179 (N_2179,N_1543,N_1626);
and U2180 (N_2180,N_1944,N_1920);
or U2181 (N_2181,N_1997,N_1909);
or U2182 (N_2182,N_1695,N_1618);
xor U2183 (N_2183,N_1609,N_1745);
nand U2184 (N_2184,N_1968,N_1856);
xor U2185 (N_2185,N_1503,N_1797);
or U2186 (N_2186,N_1527,N_1730);
or U2187 (N_2187,N_1826,N_1602);
nor U2188 (N_2188,N_1878,N_1673);
nor U2189 (N_2189,N_1782,N_1785);
and U2190 (N_2190,N_1832,N_1759);
and U2191 (N_2191,N_1927,N_1704);
and U2192 (N_2192,N_1910,N_1547);
or U2193 (N_2193,N_1598,N_1715);
or U2194 (N_2194,N_1590,N_1955);
xor U2195 (N_2195,N_1835,N_1892);
nand U2196 (N_2196,N_1938,N_1688);
and U2197 (N_2197,N_1842,N_1855);
nor U2198 (N_2198,N_1728,N_1833);
nand U2199 (N_2199,N_1805,N_1755);
nor U2200 (N_2200,N_1549,N_1754);
nand U2201 (N_2201,N_1945,N_1951);
or U2202 (N_2202,N_1993,N_1843);
xnor U2203 (N_2203,N_1848,N_1957);
or U2204 (N_2204,N_1675,N_1534);
or U2205 (N_2205,N_1769,N_1532);
xor U2206 (N_2206,N_1753,N_1779);
xnor U2207 (N_2207,N_1722,N_1822);
and U2208 (N_2208,N_1973,N_1551);
nand U2209 (N_2209,N_1880,N_1830);
nand U2210 (N_2210,N_1737,N_1632);
xnor U2211 (N_2211,N_1649,N_1899);
nor U2212 (N_2212,N_1905,N_1670);
nand U2213 (N_2213,N_1952,N_1508);
nor U2214 (N_2214,N_1570,N_1734);
or U2215 (N_2215,N_1751,N_1578);
nand U2216 (N_2216,N_1729,N_1518);
nand U2217 (N_2217,N_1566,N_1661);
and U2218 (N_2218,N_1742,N_1959);
or U2219 (N_2219,N_1621,N_1599);
or U2220 (N_2220,N_1954,N_1828);
and U2221 (N_2221,N_1904,N_1659);
and U2222 (N_2222,N_1984,N_1761);
and U2223 (N_2223,N_1663,N_1521);
xnor U2224 (N_2224,N_1509,N_1823);
or U2225 (N_2225,N_1814,N_1515);
nand U2226 (N_2226,N_1898,N_1881);
nor U2227 (N_2227,N_1907,N_1897);
nand U2228 (N_2228,N_1607,N_1925);
or U2229 (N_2229,N_1677,N_1947);
or U2230 (N_2230,N_1550,N_1752);
or U2231 (N_2231,N_1684,N_1977);
nand U2232 (N_2232,N_1965,N_1967);
or U2233 (N_2233,N_1718,N_1821);
xnor U2234 (N_2234,N_1819,N_1817);
nor U2235 (N_2235,N_1913,N_1556);
nand U2236 (N_2236,N_1531,N_1699);
or U2237 (N_2237,N_1783,N_1939);
or U2238 (N_2238,N_1886,N_1717);
nand U2239 (N_2239,N_1903,N_1864);
xnor U2240 (N_2240,N_1710,N_1912);
nor U2241 (N_2241,N_1777,N_1874);
and U2242 (N_2242,N_1647,N_1853);
xor U2243 (N_2243,N_1721,N_1713);
nor U2244 (N_2244,N_1914,N_1940);
and U2245 (N_2245,N_1558,N_1865);
nor U2246 (N_2246,N_1658,N_1643);
nand U2247 (N_2247,N_1568,N_1636);
nor U2248 (N_2248,N_1760,N_1565);
xor U2249 (N_2249,N_1603,N_1619);
and U2250 (N_2250,N_1582,N_1536);
nor U2251 (N_2251,N_1948,N_1981);
or U2252 (N_2252,N_1880,N_1659);
and U2253 (N_2253,N_1582,N_1865);
and U2254 (N_2254,N_1636,N_1575);
and U2255 (N_2255,N_1662,N_1733);
or U2256 (N_2256,N_1906,N_1744);
nand U2257 (N_2257,N_1820,N_1518);
or U2258 (N_2258,N_1609,N_1920);
and U2259 (N_2259,N_1877,N_1905);
nor U2260 (N_2260,N_1513,N_1721);
nand U2261 (N_2261,N_1599,N_1788);
xnor U2262 (N_2262,N_1761,N_1531);
and U2263 (N_2263,N_1875,N_1782);
or U2264 (N_2264,N_1723,N_1830);
xor U2265 (N_2265,N_1687,N_1798);
and U2266 (N_2266,N_1946,N_1599);
and U2267 (N_2267,N_1716,N_1763);
or U2268 (N_2268,N_1873,N_1580);
xor U2269 (N_2269,N_1626,N_1928);
nand U2270 (N_2270,N_1626,N_1646);
nand U2271 (N_2271,N_1828,N_1935);
or U2272 (N_2272,N_1900,N_1534);
nor U2273 (N_2273,N_1846,N_1855);
nor U2274 (N_2274,N_1514,N_1589);
and U2275 (N_2275,N_1796,N_1883);
nand U2276 (N_2276,N_1527,N_1953);
xnor U2277 (N_2277,N_1540,N_1784);
nor U2278 (N_2278,N_1530,N_1635);
nor U2279 (N_2279,N_1863,N_1561);
nor U2280 (N_2280,N_1896,N_1862);
and U2281 (N_2281,N_1872,N_1630);
nor U2282 (N_2282,N_1858,N_1573);
xnor U2283 (N_2283,N_1751,N_1911);
xnor U2284 (N_2284,N_1714,N_1502);
nand U2285 (N_2285,N_1781,N_1508);
nand U2286 (N_2286,N_1523,N_1511);
xor U2287 (N_2287,N_1552,N_1931);
and U2288 (N_2288,N_1984,N_1530);
or U2289 (N_2289,N_1861,N_1895);
or U2290 (N_2290,N_1981,N_1557);
or U2291 (N_2291,N_1900,N_1927);
nand U2292 (N_2292,N_1759,N_1500);
and U2293 (N_2293,N_1542,N_1993);
nand U2294 (N_2294,N_1675,N_1925);
nor U2295 (N_2295,N_1752,N_1712);
or U2296 (N_2296,N_1775,N_1760);
nand U2297 (N_2297,N_1842,N_1811);
nand U2298 (N_2298,N_1809,N_1507);
and U2299 (N_2299,N_1620,N_1516);
nand U2300 (N_2300,N_1706,N_1893);
and U2301 (N_2301,N_1571,N_1801);
and U2302 (N_2302,N_1650,N_1904);
nand U2303 (N_2303,N_1938,N_1873);
nor U2304 (N_2304,N_1667,N_1975);
xnor U2305 (N_2305,N_1916,N_1744);
xnor U2306 (N_2306,N_1813,N_1944);
nor U2307 (N_2307,N_1588,N_1982);
or U2308 (N_2308,N_1530,N_1919);
xor U2309 (N_2309,N_1929,N_1704);
or U2310 (N_2310,N_1623,N_1959);
or U2311 (N_2311,N_1564,N_1652);
and U2312 (N_2312,N_1924,N_1584);
and U2313 (N_2313,N_1562,N_1806);
nand U2314 (N_2314,N_1867,N_1813);
or U2315 (N_2315,N_1862,N_1573);
nor U2316 (N_2316,N_1907,N_1734);
or U2317 (N_2317,N_1619,N_1630);
and U2318 (N_2318,N_1504,N_1558);
xnor U2319 (N_2319,N_1700,N_1514);
xnor U2320 (N_2320,N_1890,N_1818);
nand U2321 (N_2321,N_1893,N_1816);
xnor U2322 (N_2322,N_1930,N_1865);
nor U2323 (N_2323,N_1538,N_1578);
nor U2324 (N_2324,N_1976,N_1541);
or U2325 (N_2325,N_1550,N_1667);
and U2326 (N_2326,N_1804,N_1690);
or U2327 (N_2327,N_1989,N_1840);
and U2328 (N_2328,N_1851,N_1655);
nand U2329 (N_2329,N_1671,N_1809);
nand U2330 (N_2330,N_1547,N_1987);
nand U2331 (N_2331,N_1541,N_1752);
nor U2332 (N_2332,N_1521,N_1794);
or U2333 (N_2333,N_1683,N_1676);
or U2334 (N_2334,N_1984,N_1723);
and U2335 (N_2335,N_1507,N_1797);
or U2336 (N_2336,N_1773,N_1844);
xor U2337 (N_2337,N_1988,N_1990);
nor U2338 (N_2338,N_1532,N_1960);
nand U2339 (N_2339,N_1510,N_1985);
and U2340 (N_2340,N_1897,N_1573);
nand U2341 (N_2341,N_1596,N_1755);
or U2342 (N_2342,N_1550,N_1779);
and U2343 (N_2343,N_1639,N_1825);
nand U2344 (N_2344,N_1748,N_1901);
nor U2345 (N_2345,N_1617,N_1865);
nand U2346 (N_2346,N_1780,N_1713);
xor U2347 (N_2347,N_1701,N_1649);
and U2348 (N_2348,N_1773,N_1741);
nand U2349 (N_2349,N_1829,N_1681);
and U2350 (N_2350,N_1546,N_1929);
xnor U2351 (N_2351,N_1761,N_1791);
nand U2352 (N_2352,N_1820,N_1706);
xor U2353 (N_2353,N_1902,N_1798);
nand U2354 (N_2354,N_1948,N_1943);
or U2355 (N_2355,N_1943,N_1698);
or U2356 (N_2356,N_1566,N_1606);
and U2357 (N_2357,N_1661,N_1537);
xnor U2358 (N_2358,N_1653,N_1800);
and U2359 (N_2359,N_1606,N_1713);
or U2360 (N_2360,N_1937,N_1674);
nor U2361 (N_2361,N_1551,N_1924);
nand U2362 (N_2362,N_1590,N_1864);
nand U2363 (N_2363,N_1699,N_1682);
nor U2364 (N_2364,N_1763,N_1739);
xor U2365 (N_2365,N_1632,N_1766);
or U2366 (N_2366,N_1838,N_1586);
nor U2367 (N_2367,N_1588,N_1706);
nor U2368 (N_2368,N_1813,N_1901);
nand U2369 (N_2369,N_1632,N_1887);
nor U2370 (N_2370,N_1801,N_1877);
xor U2371 (N_2371,N_1646,N_1530);
xnor U2372 (N_2372,N_1786,N_1853);
or U2373 (N_2373,N_1847,N_1568);
or U2374 (N_2374,N_1985,N_1928);
or U2375 (N_2375,N_1661,N_1841);
nand U2376 (N_2376,N_1881,N_1877);
xnor U2377 (N_2377,N_1683,N_1934);
xnor U2378 (N_2378,N_1940,N_1800);
and U2379 (N_2379,N_1804,N_1721);
or U2380 (N_2380,N_1991,N_1900);
nor U2381 (N_2381,N_1553,N_1575);
nor U2382 (N_2382,N_1997,N_1562);
xor U2383 (N_2383,N_1955,N_1587);
xor U2384 (N_2384,N_1654,N_1728);
or U2385 (N_2385,N_1776,N_1946);
xor U2386 (N_2386,N_1538,N_1739);
xnor U2387 (N_2387,N_1543,N_1510);
nand U2388 (N_2388,N_1928,N_1547);
xnor U2389 (N_2389,N_1719,N_1514);
or U2390 (N_2390,N_1946,N_1749);
nand U2391 (N_2391,N_1939,N_1594);
or U2392 (N_2392,N_1890,N_1655);
or U2393 (N_2393,N_1511,N_1587);
and U2394 (N_2394,N_1987,N_1613);
or U2395 (N_2395,N_1999,N_1892);
xnor U2396 (N_2396,N_1636,N_1982);
or U2397 (N_2397,N_1678,N_1764);
nand U2398 (N_2398,N_1563,N_1542);
or U2399 (N_2399,N_1845,N_1623);
nor U2400 (N_2400,N_1904,N_1778);
nand U2401 (N_2401,N_1819,N_1850);
and U2402 (N_2402,N_1979,N_1793);
and U2403 (N_2403,N_1835,N_1802);
or U2404 (N_2404,N_1893,N_1906);
or U2405 (N_2405,N_1614,N_1767);
and U2406 (N_2406,N_1660,N_1885);
nor U2407 (N_2407,N_1604,N_1796);
nor U2408 (N_2408,N_1658,N_1933);
nand U2409 (N_2409,N_1846,N_1739);
xor U2410 (N_2410,N_1792,N_1855);
nand U2411 (N_2411,N_1508,N_1687);
nand U2412 (N_2412,N_1540,N_1886);
nand U2413 (N_2413,N_1577,N_1836);
xnor U2414 (N_2414,N_1502,N_1705);
or U2415 (N_2415,N_1940,N_1874);
xnor U2416 (N_2416,N_1587,N_1895);
and U2417 (N_2417,N_1831,N_1713);
or U2418 (N_2418,N_1960,N_1524);
or U2419 (N_2419,N_1741,N_1866);
nor U2420 (N_2420,N_1669,N_1744);
or U2421 (N_2421,N_1989,N_1865);
xnor U2422 (N_2422,N_1580,N_1719);
or U2423 (N_2423,N_1805,N_1992);
and U2424 (N_2424,N_1621,N_1680);
or U2425 (N_2425,N_1792,N_1896);
xnor U2426 (N_2426,N_1505,N_1645);
nand U2427 (N_2427,N_1963,N_1799);
or U2428 (N_2428,N_1592,N_1716);
xnor U2429 (N_2429,N_1779,N_1669);
nor U2430 (N_2430,N_1620,N_1538);
nand U2431 (N_2431,N_1977,N_1891);
or U2432 (N_2432,N_1578,N_1854);
xnor U2433 (N_2433,N_1845,N_1502);
and U2434 (N_2434,N_1554,N_1741);
xor U2435 (N_2435,N_1580,N_1799);
nor U2436 (N_2436,N_1572,N_1688);
xor U2437 (N_2437,N_1757,N_1843);
xor U2438 (N_2438,N_1627,N_1918);
xnor U2439 (N_2439,N_1857,N_1625);
or U2440 (N_2440,N_1636,N_1704);
xnor U2441 (N_2441,N_1673,N_1985);
and U2442 (N_2442,N_1671,N_1619);
or U2443 (N_2443,N_1761,N_1678);
nor U2444 (N_2444,N_1847,N_1622);
nor U2445 (N_2445,N_1571,N_1612);
nand U2446 (N_2446,N_1666,N_1870);
nand U2447 (N_2447,N_1505,N_1858);
nor U2448 (N_2448,N_1895,N_1974);
and U2449 (N_2449,N_1813,N_1564);
nand U2450 (N_2450,N_1571,N_1855);
or U2451 (N_2451,N_1613,N_1673);
nor U2452 (N_2452,N_1811,N_1608);
or U2453 (N_2453,N_1933,N_1972);
or U2454 (N_2454,N_1666,N_1588);
nand U2455 (N_2455,N_1947,N_1655);
or U2456 (N_2456,N_1961,N_1661);
xnor U2457 (N_2457,N_1581,N_1897);
xor U2458 (N_2458,N_1919,N_1909);
and U2459 (N_2459,N_1747,N_1984);
and U2460 (N_2460,N_1913,N_1817);
xor U2461 (N_2461,N_1539,N_1882);
and U2462 (N_2462,N_1583,N_1632);
nand U2463 (N_2463,N_1853,N_1609);
and U2464 (N_2464,N_1809,N_1954);
or U2465 (N_2465,N_1576,N_1963);
and U2466 (N_2466,N_1549,N_1718);
xnor U2467 (N_2467,N_1767,N_1562);
and U2468 (N_2468,N_1802,N_1863);
xor U2469 (N_2469,N_1768,N_1680);
and U2470 (N_2470,N_1647,N_1919);
nand U2471 (N_2471,N_1803,N_1646);
and U2472 (N_2472,N_1749,N_1783);
nand U2473 (N_2473,N_1836,N_1970);
and U2474 (N_2474,N_1516,N_1711);
nor U2475 (N_2475,N_1565,N_1901);
nand U2476 (N_2476,N_1935,N_1690);
or U2477 (N_2477,N_1603,N_1951);
nand U2478 (N_2478,N_1701,N_1665);
nor U2479 (N_2479,N_1508,N_1741);
and U2480 (N_2480,N_1829,N_1972);
and U2481 (N_2481,N_1630,N_1711);
or U2482 (N_2482,N_1718,N_1590);
nand U2483 (N_2483,N_1754,N_1589);
nor U2484 (N_2484,N_1658,N_1613);
or U2485 (N_2485,N_1541,N_1798);
and U2486 (N_2486,N_1930,N_1948);
nor U2487 (N_2487,N_1955,N_1576);
xnor U2488 (N_2488,N_1508,N_1785);
or U2489 (N_2489,N_1787,N_1577);
nand U2490 (N_2490,N_1649,N_1973);
nor U2491 (N_2491,N_1707,N_1596);
xnor U2492 (N_2492,N_1554,N_1855);
nor U2493 (N_2493,N_1687,N_1916);
xor U2494 (N_2494,N_1530,N_1603);
nand U2495 (N_2495,N_1742,N_1901);
nand U2496 (N_2496,N_1936,N_1744);
and U2497 (N_2497,N_1678,N_1548);
nor U2498 (N_2498,N_1963,N_1768);
xnor U2499 (N_2499,N_1922,N_1512);
and U2500 (N_2500,N_2326,N_2266);
xor U2501 (N_2501,N_2030,N_2377);
or U2502 (N_2502,N_2301,N_2201);
or U2503 (N_2503,N_2325,N_2258);
nor U2504 (N_2504,N_2439,N_2262);
nand U2505 (N_2505,N_2457,N_2397);
and U2506 (N_2506,N_2376,N_2108);
nor U2507 (N_2507,N_2305,N_2444);
or U2508 (N_2508,N_2464,N_2159);
and U2509 (N_2509,N_2206,N_2210);
or U2510 (N_2510,N_2128,N_2497);
and U2511 (N_2511,N_2079,N_2016);
nor U2512 (N_2512,N_2337,N_2199);
nor U2513 (N_2513,N_2282,N_2009);
nor U2514 (N_2514,N_2392,N_2374);
and U2515 (N_2515,N_2471,N_2263);
or U2516 (N_2516,N_2091,N_2174);
and U2517 (N_2517,N_2109,N_2454);
nand U2518 (N_2518,N_2003,N_2164);
xor U2519 (N_2519,N_2406,N_2387);
xor U2520 (N_2520,N_2460,N_2084);
or U2521 (N_2521,N_2130,N_2411);
nor U2522 (N_2522,N_2299,N_2092);
xnor U2523 (N_2523,N_2083,N_2099);
xnor U2524 (N_2524,N_2235,N_2456);
and U2525 (N_2525,N_2081,N_2316);
nor U2526 (N_2526,N_2488,N_2272);
nor U2527 (N_2527,N_2175,N_2469);
xnor U2528 (N_2528,N_2320,N_2297);
nand U2529 (N_2529,N_2451,N_2322);
xnor U2530 (N_2530,N_2370,N_2340);
nor U2531 (N_2531,N_2186,N_2170);
nand U2532 (N_2532,N_2293,N_2029);
or U2533 (N_2533,N_2010,N_2119);
nor U2534 (N_2534,N_2193,N_2490);
nand U2535 (N_2535,N_2167,N_2178);
or U2536 (N_2536,N_2319,N_2085);
xor U2537 (N_2537,N_2192,N_2034);
nand U2538 (N_2538,N_2239,N_2204);
nand U2539 (N_2539,N_2446,N_2462);
nand U2540 (N_2540,N_2474,N_2379);
nor U2541 (N_2541,N_2489,N_2284);
nand U2542 (N_2542,N_2314,N_2247);
and U2543 (N_2543,N_2345,N_2477);
nor U2544 (N_2544,N_2158,N_2428);
nor U2545 (N_2545,N_2063,N_2425);
and U2546 (N_2546,N_2237,N_2101);
and U2547 (N_2547,N_2220,N_2348);
or U2548 (N_2548,N_2062,N_2071);
and U2549 (N_2549,N_2172,N_2267);
or U2550 (N_2550,N_2385,N_2410);
nand U2551 (N_2551,N_2485,N_2156);
nand U2552 (N_2552,N_2389,N_2046);
nand U2553 (N_2553,N_2194,N_2097);
and U2554 (N_2554,N_2366,N_2176);
nand U2555 (N_2555,N_2346,N_2390);
and U2556 (N_2556,N_2250,N_2145);
or U2557 (N_2557,N_2227,N_2349);
nand U2558 (N_2558,N_2042,N_2278);
xor U2559 (N_2559,N_2498,N_2365);
nor U2560 (N_2560,N_2430,N_2458);
xnor U2561 (N_2561,N_2090,N_2190);
or U2562 (N_2562,N_2187,N_2226);
or U2563 (N_2563,N_2126,N_2154);
nor U2564 (N_2564,N_2219,N_2122);
and U2565 (N_2565,N_2058,N_2106);
nor U2566 (N_2566,N_2286,N_2142);
nor U2567 (N_2567,N_2173,N_2323);
or U2568 (N_2568,N_2310,N_2399);
or U2569 (N_2569,N_2086,N_2236);
nand U2570 (N_2570,N_2149,N_2221);
or U2571 (N_2571,N_2300,N_2136);
nor U2572 (N_2572,N_2036,N_2394);
nor U2573 (N_2573,N_2461,N_2495);
and U2574 (N_2574,N_2232,N_2276);
or U2575 (N_2575,N_2309,N_2017);
or U2576 (N_2576,N_2080,N_2171);
and U2577 (N_2577,N_2327,N_2165);
or U2578 (N_2578,N_2419,N_2100);
xnor U2579 (N_2579,N_2351,N_2264);
nor U2580 (N_2580,N_2089,N_2465);
nor U2581 (N_2581,N_2146,N_2115);
nor U2582 (N_2582,N_2185,N_2166);
and U2583 (N_2583,N_2358,N_2482);
and U2584 (N_2584,N_2144,N_2212);
nor U2585 (N_2585,N_2373,N_2414);
nand U2586 (N_2586,N_2254,N_2066);
and U2587 (N_2587,N_2049,N_2306);
nand U2588 (N_2588,N_2131,N_2354);
nand U2589 (N_2589,N_2007,N_2033);
nand U2590 (N_2590,N_2476,N_2015);
or U2591 (N_2591,N_2412,N_2436);
and U2592 (N_2592,N_2160,N_2055);
nand U2593 (N_2593,N_2277,N_2271);
nor U2594 (N_2594,N_2135,N_2162);
nor U2595 (N_2595,N_2118,N_2295);
nand U2596 (N_2596,N_2179,N_2259);
or U2597 (N_2597,N_2127,N_2393);
xor U2598 (N_2598,N_2381,N_2022);
xnor U2599 (N_2599,N_2112,N_2077);
and U2600 (N_2600,N_2481,N_2231);
xor U2601 (N_2601,N_2230,N_2245);
or U2602 (N_2602,N_2361,N_2150);
nor U2603 (N_2603,N_2027,N_2255);
nand U2604 (N_2604,N_2360,N_2494);
or U2605 (N_2605,N_2432,N_2496);
or U2606 (N_2606,N_2076,N_2023);
nand U2607 (N_2607,N_2296,N_2125);
xnor U2608 (N_2608,N_2478,N_2350);
and U2609 (N_2609,N_2362,N_2054);
xor U2610 (N_2610,N_2057,N_2020);
or U2611 (N_2611,N_2026,N_2208);
xor U2612 (N_2612,N_2141,N_2233);
and U2613 (N_2613,N_2211,N_2265);
nor U2614 (N_2614,N_2429,N_2243);
or U2615 (N_2615,N_2292,N_2355);
xnor U2616 (N_2616,N_2369,N_2353);
nand U2617 (N_2617,N_2396,N_2281);
and U2618 (N_2618,N_2134,N_2329);
or U2619 (N_2619,N_2438,N_2275);
nor U2620 (N_2620,N_2363,N_2068);
nor U2621 (N_2621,N_2384,N_2442);
or U2622 (N_2622,N_2422,N_2098);
nor U2623 (N_2623,N_2060,N_2487);
or U2624 (N_2624,N_2491,N_2336);
and U2625 (N_2625,N_2044,N_2308);
nor U2626 (N_2626,N_2008,N_2217);
nand U2627 (N_2627,N_2463,N_2334);
and U2628 (N_2628,N_2163,N_2143);
xnor U2629 (N_2629,N_2234,N_2242);
nand U2630 (N_2630,N_2096,N_2005);
nor U2631 (N_2631,N_2002,N_2433);
or U2632 (N_2632,N_2352,N_2484);
and U2633 (N_2633,N_2472,N_2061);
and U2634 (N_2634,N_2056,N_2018);
nor U2635 (N_2635,N_2338,N_2213);
and U2636 (N_2636,N_2486,N_2339);
nor U2637 (N_2637,N_2011,N_2424);
xor U2638 (N_2638,N_2151,N_2229);
nand U2639 (N_2639,N_2045,N_2048);
nor U2640 (N_2640,N_2116,N_2435);
or U2641 (N_2641,N_2408,N_2447);
nor U2642 (N_2642,N_2443,N_2195);
xor U2643 (N_2643,N_2386,N_2312);
and U2644 (N_2644,N_2287,N_2274);
nand U2645 (N_2645,N_2240,N_2238);
and U2646 (N_2646,N_2357,N_2391);
xor U2647 (N_2647,N_2205,N_2270);
and U2648 (N_2648,N_2417,N_2449);
and U2649 (N_2649,N_2304,N_2401);
and U2650 (N_2650,N_2431,N_2050);
xnor U2651 (N_2651,N_2480,N_2182);
and U2652 (N_2652,N_2405,N_2180);
nand U2653 (N_2653,N_2222,N_2492);
nor U2654 (N_2654,N_2133,N_2418);
nor U2655 (N_2655,N_2289,N_2398);
xnor U2656 (N_2656,N_2021,N_2333);
and U2657 (N_2657,N_2024,N_2437);
or U2658 (N_2658,N_2001,N_2403);
and U2659 (N_2659,N_2343,N_2268);
nand U2660 (N_2660,N_2177,N_2423);
or U2661 (N_2661,N_2388,N_2452);
or U2662 (N_2662,N_2285,N_2032);
or U2663 (N_2663,N_2256,N_2040);
or U2664 (N_2664,N_2012,N_2121);
xnor U2665 (N_2665,N_2123,N_2038);
and U2666 (N_2666,N_2499,N_2420);
xnor U2667 (N_2667,N_2302,N_2409);
or U2668 (N_2668,N_2196,N_2102);
or U2669 (N_2669,N_2161,N_2359);
or U2670 (N_2670,N_2198,N_2107);
or U2671 (N_2671,N_2072,N_2459);
or U2672 (N_2672,N_2468,N_2070);
or U2673 (N_2673,N_2047,N_2067);
nand U2674 (N_2674,N_2105,N_2073);
or U2675 (N_2675,N_2152,N_2241);
and U2676 (N_2676,N_2153,N_2111);
or U2677 (N_2677,N_2248,N_2004);
nor U2678 (N_2678,N_2332,N_2280);
nand U2679 (N_2679,N_2169,N_2218);
nor U2680 (N_2680,N_2069,N_2000);
and U2681 (N_2681,N_2328,N_2139);
and U2682 (N_2682,N_2244,N_2147);
nand U2683 (N_2683,N_2039,N_2183);
nor U2684 (N_2684,N_2344,N_2028);
nor U2685 (N_2685,N_2367,N_2124);
nor U2686 (N_2686,N_2426,N_2473);
nor U2687 (N_2687,N_2246,N_2455);
and U2688 (N_2688,N_2291,N_2303);
nand U2689 (N_2689,N_2202,N_2224);
or U2690 (N_2690,N_2315,N_2261);
and U2691 (N_2691,N_2014,N_2317);
or U2692 (N_2692,N_2129,N_2324);
or U2693 (N_2693,N_2382,N_2434);
xnor U2694 (N_2694,N_2228,N_2168);
and U2695 (N_2695,N_2082,N_2307);
and U2696 (N_2696,N_2019,N_2031);
nand U2697 (N_2697,N_2025,N_2203);
xor U2698 (N_2698,N_2137,N_2253);
or U2699 (N_2699,N_2257,N_2157);
xor U2700 (N_2700,N_2294,N_2037);
or U2701 (N_2701,N_2404,N_2252);
or U2702 (N_2702,N_2311,N_2260);
or U2703 (N_2703,N_2269,N_2155);
nand U2704 (N_2704,N_2402,N_2356);
or U2705 (N_2705,N_2181,N_2075);
nand U2706 (N_2706,N_2117,N_2445);
nor U2707 (N_2707,N_2197,N_2138);
or U2708 (N_2708,N_2330,N_2104);
xnor U2709 (N_2709,N_2251,N_2103);
nor U2710 (N_2710,N_2493,N_2450);
xor U2711 (N_2711,N_2216,N_2470);
and U2712 (N_2712,N_2215,N_2120);
nor U2713 (N_2713,N_2347,N_2200);
nor U2714 (N_2714,N_2207,N_2051);
nand U2715 (N_2715,N_2132,N_2368);
and U2716 (N_2716,N_2059,N_2087);
xor U2717 (N_2717,N_2148,N_2318);
nand U2718 (N_2718,N_2114,N_2052);
nand U2719 (N_2719,N_2415,N_2467);
and U2720 (N_2720,N_2380,N_2088);
and U2721 (N_2721,N_2095,N_2013);
or U2722 (N_2722,N_2093,N_2331);
nor U2723 (N_2723,N_2283,N_2298);
or U2724 (N_2724,N_2223,N_2209);
nor U2725 (N_2725,N_2078,N_2453);
or U2726 (N_2726,N_2335,N_2053);
xor U2727 (N_2727,N_2184,N_2249);
or U2728 (N_2728,N_2479,N_2372);
xor U2729 (N_2729,N_2225,N_2341);
nor U2730 (N_2730,N_2441,N_2035);
xnor U2731 (N_2731,N_2110,N_2279);
or U2732 (N_2732,N_2065,N_2427);
xor U2733 (N_2733,N_2375,N_2395);
and U2734 (N_2734,N_2191,N_2313);
xnor U2735 (N_2735,N_2189,N_2288);
and U2736 (N_2736,N_2407,N_2364);
or U2737 (N_2737,N_2041,N_2140);
nor U2738 (N_2738,N_2006,N_2383);
or U2739 (N_2739,N_2214,N_2113);
nand U2740 (N_2740,N_2273,N_2290);
xor U2741 (N_2741,N_2371,N_2416);
nor U2742 (N_2742,N_2413,N_2064);
nor U2743 (N_2743,N_2342,N_2483);
nor U2744 (N_2744,N_2188,N_2074);
and U2745 (N_2745,N_2378,N_2448);
or U2746 (N_2746,N_2475,N_2400);
xnor U2747 (N_2747,N_2321,N_2466);
or U2748 (N_2748,N_2094,N_2421);
xnor U2749 (N_2749,N_2043,N_2440);
and U2750 (N_2750,N_2004,N_2288);
xnor U2751 (N_2751,N_2074,N_2309);
nor U2752 (N_2752,N_2118,N_2463);
nand U2753 (N_2753,N_2216,N_2344);
nand U2754 (N_2754,N_2150,N_2096);
or U2755 (N_2755,N_2011,N_2469);
and U2756 (N_2756,N_2225,N_2095);
nand U2757 (N_2757,N_2376,N_2162);
xnor U2758 (N_2758,N_2285,N_2059);
and U2759 (N_2759,N_2053,N_2142);
nor U2760 (N_2760,N_2478,N_2455);
or U2761 (N_2761,N_2250,N_2183);
nand U2762 (N_2762,N_2366,N_2407);
and U2763 (N_2763,N_2163,N_2228);
xnor U2764 (N_2764,N_2310,N_2055);
xnor U2765 (N_2765,N_2067,N_2451);
xor U2766 (N_2766,N_2235,N_2325);
or U2767 (N_2767,N_2257,N_2279);
nor U2768 (N_2768,N_2382,N_2348);
xnor U2769 (N_2769,N_2122,N_2350);
or U2770 (N_2770,N_2433,N_2209);
and U2771 (N_2771,N_2313,N_2374);
or U2772 (N_2772,N_2218,N_2088);
xor U2773 (N_2773,N_2362,N_2324);
nand U2774 (N_2774,N_2477,N_2191);
and U2775 (N_2775,N_2045,N_2329);
nor U2776 (N_2776,N_2182,N_2345);
xnor U2777 (N_2777,N_2043,N_2098);
and U2778 (N_2778,N_2212,N_2172);
or U2779 (N_2779,N_2087,N_2298);
nor U2780 (N_2780,N_2138,N_2424);
nand U2781 (N_2781,N_2038,N_2476);
nand U2782 (N_2782,N_2489,N_2403);
and U2783 (N_2783,N_2198,N_2169);
nor U2784 (N_2784,N_2164,N_2478);
nand U2785 (N_2785,N_2205,N_2197);
nand U2786 (N_2786,N_2115,N_2061);
and U2787 (N_2787,N_2440,N_2366);
and U2788 (N_2788,N_2461,N_2074);
or U2789 (N_2789,N_2150,N_2485);
xnor U2790 (N_2790,N_2490,N_2110);
xnor U2791 (N_2791,N_2063,N_2421);
or U2792 (N_2792,N_2460,N_2356);
xor U2793 (N_2793,N_2385,N_2383);
nand U2794 (N_2794,N_2190,N_2404);
and U2795 (N_2795,N_2321,N_2105);
and U2796 (N_2796,N_2150,N_2161);
and U2797 (N_2797,N_2318,N_2396);
or U2798 (N_2798,N_2124,N_2361);
or U2799 (N_2799,N_2429,N_2140);
nand U2800 (N_2800,N_2343,N_2113);
xor U2801 (N_2801,N_2145,N_2489);
nand U2802 (N_2802,N_2111,N_2131);
or U2803 (N_2803,N_2424,N_2159);
or U2804 (N_2804,N_2356,N_2383);
xor U2805 (N_2805,N_2070,N_2364);
nor U2806 (N_2806,N_2456,N_2127);
xnor U2807 (N_2807,N_2443,N_2334);
and U2808 (N_2808,N_2396,N_2477);
xor U2809 (N_2809,N_2129,N_2479);
nor U2810 (N_2810,N_2404,N_2184);
nor U2811 (N_2811,N_2270,N_2055);
nand U2812 (N_2812,N_2291,N_2330);
nor U2813 (N_2813,N_2398,N_2225);
or U2814 (N_2814,N_2489,N_2057);
and U2815 (N_2815,N_2136,N_2364);
or U2816 (N_2816,N_2328,N_2064);
nor U2817 (N_2817,N_2330,N_2440);
xor U2818 (N_2818,N_2463,N_2155);
nor U2819 (N_2819,N_2427,N_2412);
nand U2820 (N_2820,N_2459,N_2402);
nor U2821 (N_2821,N_2099,N_2102);
or U2822 (N_2822,N_2365,N_2131);
nand U2823 (N_2823,N_2325,N_2120);
or U2824 (N_2824,N_2098,N_2469);
and U2825 (N_2825,N_2324,N_2165);
nor U2826 (N_2826,N_2178,N_2216);
or U2827 (N_2827,N_2173,N_2392);
nand U2828 (N_2828,N_2401,N_2414);
xnor U2829 (N_2829,N_2229,N_2065);
or U2830 (N_2830,N_2036,N_2484);
xor U2831 (N_2831,N_2283,N_2291);
xnor U2832 (N_2832,N_2293,N_2049);
or U2833 (N_2833,N_2251,N_2025);
or U2834 (N_2834,N_2306,N_2034);
and U2835 (N_2835,N_2318,N_2049);
nand U2836 (N_2836,N_2284,N_2109);
nand U2837 (N_2837,N_2073,N_2287);
nor U2838 (N_2838,N_2310,N_2226);
nor U2839 (N_2839,N_2461,N_2220);
xor U2840 (N_2840,N_2433,N_2107);
nand U2841 (N_2841,N_2488,N_2275);
xnor U2842 (N_2842,N_2248,N_2212);
and U2843 (N_2843,N_2311,N_2065);
and U2844 (N_2844,N_2464,N_2384);
or U2845 (N_2845,N_2121,N_2172);
or U2846 (N_2846,N_2284,N_2222);
nor U2847 (N_2847,N_2371,N_2000);
nand U2848 (N_2848,N_2363,N_2478);
nor U2849 (N_2849,N_2421,N_2354);
nor U2850 (N_2850,N_2078,N_2219);
nor U2851 (N_2851,N_2199,N_2069);
or U2852 (N_2852,N_2209,N_2235);
or U2853 (N_2853,N_2479,N_2373);
xor U2854 (N_2854,N_2061,N_2323);
and U2855 (N_2855,N_2136,N_2312);
nor U2856 (N_2856,N_2287,N_2093);
or U2857 (N_2857,N_2037,N_2389);
or U2858 (N_2858,N_2365,N_2233);
and U2859 (N_2859,N_2430,N_2111);
nand U2860 (N_2860,N_2181,N_2076);
nand U2861 (N_2861,N_2269,N_2480);
nor U2862 (N_2862,N_2451,N_2324);
or U2863 (N_2863,N_2484,N_2102);
or U2864 (N_2864,N_2276,N_2085);
xor U2865 (N_2865,N_2294,N_2247);
or U2866 (N_2866,N_2308,N_2312);
or U2867 (N_2867,N_2037,N_2296);
nand U2868 (N_2868,N_2212,N_2258);
or U2869 (N_2869,N_2409,N_2390);
xor U2870 (N_2870,N_2138,N_2367);
or U2871 (N_2871,N_2206,N_2232);
or U2872 (N_2872,N_2484,N_2183);
nand U2873 (N_2873,N_2127,N_2093);
or U2874 (N_2874,N_2487,N_2386);
and U2875 (N_2875,N_2327,N_2423);
nor U2876 (N_2876,N_2272,N_2067);
nand U2877 (N_2877,N_2472,N_2423);
xor U2878 (N_2878,N_2185,N_2441);
and U2879 (N_2879,N_2146,N_2167);
xor U2880 (N_2880,N_2434,N_2163);
and U2881 (N_2881,N_2038,N_2384);
xor U2882 (N_2882,N_2389,N_2242);
and U2883 (N_2883,N_2029,N_2444);
nand U2884 (N_2884,N_2272,N_2077);
xnor U2885 (N_2885,N_2166,N_2340);
and U2886 (N_2886,N_2466,N_2086);
and U2887 (N_2887,N_2036,N_2324);
or U2888 (N_2888,N_2290,N_2302);
nor U2889 (N_2889,N_2485,N_2044);
or U2890 (N_2890,N_2217,N_2204);
nor U2891 (N_2891,N_2379,N_2478);
nand U2892 (N_2892,N_2148,N_2289);
nor U2893 (N_2893,N_2143,N_2013);
xnor U2894 (N_2894,N_2495,N_2044);
nand U2895 (N_2895,N_2424,N_2300);
nor U2896 (N_2896,N_2421,N_2489);
or U2897 (N_2897,N_2160,N_2470);
nand U2898 (N_2898,N_2246,N_2066);
nor U2899 (N_2899,N_2440,N_2206);
and U2900 (N_2900,N_2077,N_2178);
xor U2901 (N_2901,N_2230,N_2065);
nand U2902 (N_2902,N_2255,N_2014);
and U2903 (N_2903,N_2298,N_2102);
nor U2904 (N_2904,N_2270,N_2256);
and U2905 (N_2905,N_2405,N_2303);
or U2906 (N_2906,N_2156,N_2298);
nor U2907 (N_2907,N_2303,N_2382);
nor U2908 (N_2908,N_2270,N_2472);
nand U2909 (N_2909,N_2250,N_2417);
nand U2910 (N_2910,N_2199,N_2089);
xnor U2911 (N_2911,N_2445,N_2191);
and U2912 (N_2912,N_2021,N_2027);
xor U2913 (N_2913,N_2473,N_2146);
nand U2914 (N_2914,N_2033,N_2378);
xor U2915 (N_2915,N_2295,N_2375);
nor U2916 (N_2916,N_2109,N_2159);
and U2917 (N_2917,N_2027,N_2063);
or U2918 (N_2918,N_2129,N_2141);
nand U2919 (N_2919,N_2255,N_2489);
xor U2920 (N_2920,N_2247,N_2109);
and U2921 (N_2921,N_2431,N_2455);
or U2922 (N_2922,N_2327,N_2331);
nand U2923 (N_2923,N_2363,N_2288);
nand U2924 (N_2924,N_2437,N_2494);
and U2925 (N_2925,N_2474,N_2371);
nand U2926 (N_2926,N_2399,N_2272);
or U2927 (N_2927,N_2230,N_2403);
xor U2928 (N_2928,N_2059,N_2484);
nor U2929 (N_2929,N_2491,N_2341);
nand U2930 (N_2930,N_2058,N_2430);
and U2931 (N_2931,N_2233,N_2204);
nand U2932 (N_2932,N_2343,N_2397);
nand U2933 (N_2933,N_2005,N_2330);
nand U2934 (N_2934,N_2446,N_2195);
nand U2935 (N_2935,N_2325,N_2441);
xor U2936 (N_2936,N_2129,N_2196);
and U2937 (N_2937,N_2430,N_2264);
nor U2938 (N_2938,N_2210,N_2098);
xnor U2939 (N_2939,N_2431,N_2264);
and U2940 (N_2940,N_2349,N_2128);
xor U2941 (N_2941,N_2343,N_2171);
and U2942 (N_2942,N_2003,N_2109);
and U2943 (N_2943,N_2171,N_2249);
or U2944 (N_2944,N_2197,N_2437);
xor U2945 (N_2945,N_2305,N_2104);
xnor U2946 (N_2946,N_2329,N_2450);
and U2947 (N_2947,N_2034,N_2378);
or U2948 (N_2948,N_2413,N_2238);
or U2949 (N_2949,N_2259,N_2140);
xor U2950 (N_2950,N_2226,N_2327);
nor U2951 (N_2951,N_2119,N_2070);
or U2952 (N_2952,N_2337,N_2382);
nor U2953 (N_2953,N_2459,N_2345);
or U2954 (N_2954,N_2086,N_2033);
nor U2955 (N_2955,N_2117,N_2289);
or U2956 (N_2956,N_2382,N_2188);
and U2957 (N_2957,N_2301,N_2369);
nor U2958 (N_2958,N_2160,N_2073);
and U2959 (N_2959,N_2176,N_2074);
and U2960 (N_2960,N_2175,N_2439);
or U2961 (N_2961,N_2155,N_2197);
nor U2962 (N_2962,N_2123,N_2477);
nand U2963 (N_2963,N_2470,N_2293);
and U2964 (N_2964,N_2460,N_2442);
and U2965 (N_2965,N_2387,N_2135);
xnor U2966 (N_2966,N_2349,N_2372);
xor U2967 (N_2967,N_2172,N_2030);
nand U2968 (N_2968,N_2030,N_2116);
and U2969 (N_2969,N_2422,N_2262);
xor U2970 (N_2970,N_2121,N_2022);
nand U2971 (N_2971,N_2013,N_2147);
nand U2972 (N_2972,N_2044,N_2413);
xnor U2973 (N_2973,N_2094,N_2322);
nand U2974 (N_2974,N_2494,N_2424);
xor U2975 (N_2975,N_2333,N_2358);
or U2976 (N_2976,N_2084,N_2080);
xnor U2977 (N_2977,N_2379,N_2346);
xnor U2978 (N_2978,N_2478,N_2361);
nand U2979 (N_2979,N_2466,N_2251);
and U2980 (N_2980,N_2233,N_2266);
nand U2981 (N_2981,N_2468,N_2451);
or U2982 (N_2982,N_2281,N_2304);
or U2983 (N_2983,N_2148,N_2434);
or U2984 (N_2984,N_2463,N_2367);
or U2985 (N_2985,N_2044,N_2065);
nor U2986 (N_2986,N_2343,N_2484);
nand U2987 (N_2987,N_2435,N_2460);
or U2988 (N_2988,N_2412,N_2312);
nor U2989 (N_2989,N_2230,N_2049);
nand U2990 (N_2990,N_2074,N_2001);
nor U2991 (N_2991,N_2021,N_2116);
and U2992 (N_2992,N_2167,N_2436);
and U2993 (N_2993,N_2268,N_2236);
or U2994 (N_2994,N_2229,N_2437);
xnor U2995 (N_2995,N_2248,N_2002);
or U2996 (N_2996,N_2042,N_2275);
and U2997 (N_2997,N_2484,N_2294);
or U2998 (N_2998,N_2441,N_2125);
and U2999 (N_2999,N_2377,N_2345);
xnor U3000 (N_3000,N_2829,N_2542);
and U3001 (N_3001,N_2513,N_2777);
xnor U3002 (N_3002,N_2602,N_2729);
nor U3003 (N_3003,N_2768,N_2921);
and U3004 (N_3004,N_2515,N_2753);
nor U3005 (N_3005,N_2675,N_2760);
xor U3006 (N_3006,N_2755,N_2703);
or U3007 (N_3007,N_2895,N_2790);
and U3008 (N_3008,N_2841,N_2506);
and U3009 (N_3009,N_2914,N_2993);
xnor U3010 (N_3010,N_2501,N_2776);
nor U3011 (N_3011,N_2764,N_2563);
and U3012 (N_3012,N_2929,N_2759);
or U3013 (N_3013,N_2652,N_2580);
nand U3014 (N_3014,N_2543,N_2836);
nor U3015 (N_3015,N_2995,N_2920);
nand U3016 (N_3016,N_2981,N_2730);
or U3017 (N_3017,N_2679,N_2527);
nor U3018 (N_3018,N_2554,N_2819);
or U3019 (N_3019,N_2880,N_2528);
and U3020 (N_3020,N_2797,N_2644);
nor U3021 (N_3021,N_2840,N_2844);
or U3022 (N_3022,N_2851,N_2524);
nand U3023 (N_3023,N_2629,N_2509);
and U3024 (N_3024,N_2556,N_2676);
or U3025 (N_3025,N_2510,N_2953);
and U3026 (N_3026,N_2909,N_2742);
nand U3027 (N_3027,N_2706,N_2511);
and U3028 (N_3028,N_2581,N_2802);
xor U3029 (N_3029,N_2884,N_2873);
nand U3030 (N_3030,N_2565,N_2561);
or U3031 (N_3031,N_2821,N_2892);
nor U3032 (N_3032,N_2839,N_2913);
xnor U3033 (N_3033,N_2664,N_2866);
and U3034 (N_3034,N_2947,N_2812);
nand U3035 (N_3035,N_2637,N_2786);
xnor U3036 (N_3036,N_2539,N_2647);
xnor U3037 (N_3037,N_2695,N_2858);
nand U3038 (N_3038,N_2864,N_2804);
or U3039 (N_3039,N_2917,N_2994);
nand U3040 (N_3040,N_2787,N_2999);
nand U3041 (N_3041,N_2737,N_2708);
xor U3042 (N_3042,N_2714,N_2888);
or U3043 (N_3043,N_2680,N_2516);
nand U3044 (N_3044,N_2535,N_2928);
xor U3045 (N_3045,N_2793,N_2525);
nor U3046 (N_3046,N_2585,N_2719);
and U3047 (N_3047,N_2867,N_2837);
nand U3048 (N_3048,N_2523,N_2620);
and U3049 (N_3049,N_2970,N_2743);
xor U3050 (N_3050,N_2627,N_2769);
nor U3051 (N_3051,N_2887,N_2983);
or U3052 (N_3052,N_2950,N_2588);
nor U3053 (N_3053,N_2908,N_2723);
xor U3054 (N_3054,N_2607,N_2733);
and U3055 (N_3055,N_2590,N_2912);
xnor U3056 (N_3056,N_2725,N_2651);
nand U3057 (N_3057,N_2617,N_2757);
nor U3058 (N_3058,N_2848,N_2538);
nand U3059 (N_3059,N_2766,N_2572);
and U3060 (N_3060,N_2842,N_2882);
or U3061 (N_3061,N_2685,N_2978);
nand U3062 (N_3062,N_2910,N_2689);
nand U3063 (N_3063,N_2943,N_2656);
nand U3064 (N_3064,N_2870,N_2838);
and U3065 (N_3065,N_2872,N_2720);
and U3066 (N_3066,N_2849,N_2726);
nor U3067 (N_3067,N_2820,N_2852);
and U3068 (N_3068,N_2750,N_2518);
nand U3069 (N_3069,N_2717,N_2876);
or U3070 (N_3070,N_2517,N_2809);
xnor U3071 (N_3071,N_2728,N_2628);
nor U3072 (N_3072,N_2775,N_2653);
xor U3073 (N_3073,N_2878,N_2765);
or U3074 (N_3074,N_2705,N_2770);
xor U3075 (N_3075,N_2871,N_2575);
and U3076 (N_3076,N_2968,N_2808);
or U3077 (N_3077,N_2500,N_2589);
nor U3078 (N_3078,N_2532,N_2857);
and U3079 (N_3079,N_2890,N_2537);
or U3080 (N_3080,N_2571,N_2562);
xor U3081 (N_3081,N_2605,N_2697);
xor U3082 (N_3082,N_2926,N_2966);
xnor U3083 (N_3083,N_2818,N_2716);
nor U3084 (N_3084,N_2860,N_2584);
or U3085 (N_3085,N_2891,N_2748);
and U3086 (N_3086,N_2683,N_2958);
and U3087 (N_3087,N_2923,N_2698);
or U3088 (N_3088,N_2788,N_2833);
nor U3089 (N_3089,N_2813,N_2996);
nor U3090 (N_3090,N_2552,N_2547);
and U3091 (N_3091,N_2560,N_2902);
nor U3092 (N_3092,N_2930,N_2877);
xor U3093 (N_3093,N_2622,N_2810);
nor U3094 (N_3094,N_2661,N_2696);
xor U3095 (N_3095,N_2530,N_2569);
or U3096 (N_3096,N_2843,N_2774);
nand U3097 (N_3097,N_2568,N_2739);
xor U3098 (N_3098,N_2938,N_2925);
or U3099 (N_3099,N_2614,N_2933);
nor U3100 (N_3100,N_2657,N_2710);
or U3101 (N_3101,N_2756,N_2896);
nor U3102 (N_3102,N_2915,N_2905);
or U3103 (N_3103,N_2754,N_2747);
nand U3104 (N_3104,N_2597,N_2798);
or U3105 (N_3105,N_2736,N_2550);
or U3106 (N_3106,N_2971,N_2713);
nor U3107 (N_3107,N_2540,N_2972);
xor U3108 (N_3108,N_2574,N_2967);
nor U3109 (N_3109,N_2988,N_2639);
nand U3110 (N_3110,N_2856,N_2514);
nor U3111 (N_3111,N_2623,N_2566);
and U3112 (N_3112,N_2507,N_2816);
and U3113 (N_3113,N_2785,N_2658);
xnor U3114 (N_3114,N_2721,N_2941);
nand U3115 (N_3115,N_2669,N_2740);
nor U3116 (N_3116,N_2519,N_2626);
nand U3117 (N_3117,N_2801,N_2603);
or U3118 (N_3118,N_2502,N_2783);
nand U3119 (N_3119,N_2612,N_2654);
nand U3120 (N_3120,N_2645,N_2951);
nand U3121 (N_3121,N_2782,N_2591);
or U3122 (N_3122,N_2897,N_2544);
and U3123 (N_3123,N_2570,N_2663);
or U3124 (N_3124,N_2799,N_2780);
and U3125 (N_3125,N_2800,N_2508);
nand U3126 (N_3126,N_2667,N_2850);
nand U3127 (N_3127,N_2702,N_2666);
nor U3128 (N_3128,N_2636,N_2650);
or U3129 (N_3129,N_2907,N_2986);
and U3130 (N_3130,N_2583,N_2903);
or U3131 (N_3131,N_2735,N_2779);
xor U3132 (N_3132,N_2611,N_2946);
or U3133 (N_3133,N_2746,N_2642);
nand U3134 (N_3134,N_2869,N_2724);
xnor U3135 (N_3135,N_2648,N_2964);
or U3136 (N_3136,N_2660,N_2604);
and U3137 (N_3137,N_2825,N_2963);
xnor U3138 (N_3138,N_2893,N_2789);
nor U3139 (N_3139,N_2635,N_2762);
nor U3140 (N_3140,N_2715,N_2973);
or U3141 (N_3141,N_2662,N_2997);
or U3142 (N_3142,N_2707,N_2618);
nor U3143 (N_3143,N_2874,N_2936);
nor U3144 (N_3144,N_2806,N_2727);
xor U3145 (N_3145,N_2805,N_2823);
nand U3146 (N_3146,N_2945,N_2734);
and U3147 (N_3147,N_2613,N_2551);
or U3148 (N_3148,N_2534,N_2633);
or U3149 (N_3149,N_2690,N_2854);
nor U3150 (N_3150,N_2558,N_2948);
nand U3151 (N_3151,N_2773,N_2791);
or U3152 (N_3152,N_2640,N_2744);
xnor U3153 (N_3153,N_2845,N_2610);
nand U3154 (N_3154,N_2646,N_2586);
nor U3155 (N_3155,N_2548,N_2886);
nor U3156 (N_3156,N_2526,N_2831);
xor U3157 (N_3157,N_2824,N_2772);
nand U3158 (N_3158,N_2582,N_2906);
xnor U3159 (N_3159,N_2670,N_2792);
and U3160 (N_3160,N_2863,N_2911);
and U3161 (N_3161,N_2985,N_2564);
and U3162 (N_3162,N_2931,N_2632);
nand U3163 (N_3163,N_2691,N_2919);
and U3164 (N_3164,N_2531,N_2522);
xnor U3165 (N_3165,N_2894,N_2932);
nor U3166 (N_3166,N_2901,N_2916);
nand U3167 (N_3167,N_2624,N_2885);
xor U3168 (N_3168,N_2763,N_2615);
nand U3169 (N_3169,N_2989,N_2593);
xor U3170 (N_3170,N_2678,N_2944);
or U3171 (N_3171,N_2541,N_2601);
nand U3172 (N_3172,N_2796,N_2606);
xor U3173 (N_3173,N_2960,N_2751);
and U3174 (N_3174,N_2828,N_2555);
or U3175 (N_3175,N_2832,N_2987);
or U3176 (N_3176,N_2795,N_2969);
nand U3177 (N_3177,N_2965,N_2974);
nor U3178 (N_3178,N_2975,N_2794);
nor U3179 (N_3179,N_2521,N_2811);
and U3180 (N_3180,N_2503,N_2577);
nand U3181 (N_3181,N_2935,N_2899);
or U3182 (N_3182,N_2784,N_2875);
nand U3183 (N_3183,N_2692,N_2942);
or U3184 (N_3184,N_2659,N_2634);
xnor U3185 (N_3185,N_2674,N_2630);
nand U3186 (N_3186,N_2701,N_2595);
and U3187 (N_3187,N_2939,N_2956);
nor U3188 (N_3188,N_2686,N_2949);
or U3189 (N_3189,N_2738,N_2937);
or U3190 (N_3190,N_2578,N_2693);
and U3191 (N_3191,N_2957,N_2573);
nand U3192 (N_3192,N_2976,N_2761);
xor U3193 (N_3193,N_2709,N_2990);
xor U3194 (N_3194,N_2668,N_2827);
and U3195 (N_3195,N_2545,N_2694);
xor U3196 (N_3196,N_2699,N_2536);
or U3197 (N_3197,N_2520,N_2980);
nor U3198 (N_3198,N_2979,N_2922);
nor U3199 (N_3199,N_2549,N_2952);
or U3200 (N_3200,N_2631,N_2940);
xnor U3201 (N_3201,N_2673,N_2862);
xor U3202 (N_3202,N_2649,N_2961);
and U3203 (N_3203,N_2883,N_2745);
xor U3204 (N_3204,N_2781,N_2619);
nand U3205 (N_3205,N_2955,N_2977);
or U3206 (N_3206,N_2767,N_2822);
and U3207 (N_3207,N_2621,N_2830);
and U3208 (N_3208,N_2722,N_2868);
or U3209 (N_3209,N_2682,N_2641);
nand U3210 (N_3210,N_2815,N_2732);
nand U3211 (N_3211,N_2553,N_2835);
nand U3212 (N_3212,N_2533,N_2879);
nand U3213 (N_3213,N_2731,N_2803);
xor U3214 (N_3214,N_2962,N_2596);
xor U3215 (N_3215,N_2557,N_2954);
nand U3216 (N_3216,N_2771,N_2579);
or U3217 (N_3217,N_2677,N_2546);
nand U3218 (N_3218,N_2700,N_2643);
xor U3219 (N_3219,N_2665,N_2688);
nor U3220 (N_3220,N_2881,N_2817);
and U3221 (N_3221,N_2600,N_2711);
nor U3222 (N_3222,N_2598,N_2861);
xor U3223 (N_3223,N_2587,N_2991);
xnor U3224 (N_3224,N_2681,N_2684);
and U3225 (N_3225,N_2992,N_2599);
or U3226 (N_3226,N_2834,N_2687);
nand U3227 (N_3227,N_2826,N_2904);
nand U3228 (N_3228,N_2655,N_2704);
nand U3229 (N_3229,N_2559,N_2859);
or U3230 (N_3230,N_2807,N_2567);
xnor U3231 (N_3231,N_2855,N_2924);
xnor U3232 (N_3232,N_2898,N_2758);
xnor U3233 (N_3233,N_2672,N_2984);
and U3234 (N_3234,N_2616,N_2594);
and U3235 (N_3235,N_2608,N_2512);
xor U3236 (N_3236,N_2576,N_2959);
or U3237 (N_3237,N_2927,N_2625);
or U3238 (N_3238,N_2505,N_2638);
and U3239 (N_3239,N_2741,N_2718);
or U3240 (N_3240,N_2934,N_2712);
nor U3241 (N_3241,N_2778,N_2865);
or U3242 (N_3242,N_2847,N_2982);
nor U3243 (N_3243,N_2889,N_2998);
or U3244 (N_3244,N_2752,N_2592);
or U3245 (N_3245,N_2918,N_2749);
nor U3246 (N_3246,N_2853,N_2671);
or U3247 (N_3247,N_2609,N_2814);
xor U3248 (N_3248,N_2846,N_2504);
and U3249 (N_3249,N_2529,N_2900);
xor U3250 (N_3250,N_2813,N_2698);
nand U3251 (N_3251,N_2519,N_2678);
or U3252 (N_3252,N_2776,N_2600);
nand U3253 (N_3253,N_2970,N_2511);
and U3254 (N_3254,N_2660,N_2978);
and U3255 (N_3255,N_2746,N_2751);
or U3256 (N_3256,N_2762,N_2537);
nand U3257 (N_3257,N_2925,N_2837);
nor U3258 (N_3258,N_2555,N_2703);
nor U3259 (N_3259,N_2581,N_2605);
nand U3260 (N_3260,N_2641,N_2918);
and U3261 (N_3261,N_2997,N_2874);
or U3262 (N_3262,N_2812,N_2789);
nand U3263 (N_3263,N_2978,N_2567);
xor U3264 (N_3264,N_2820,N_2748);
xor U3265 (N_3265,N_2523,N_2666);
nor U3266 (N_3266,N_2600,N_2660);
nor U3267 (N_3267,N_2580,N_2773);
xor U3268 (N_3268,N_2538,N_2824);
xor U3269 (N_3269,N_2595,N_2788);
nor U3270 (N_3270,N_2506,N_2843);
xor U3271 (N_3271,N_2593,N_2909);
nor U3272 (N_3272,N_2987,N_2616);
xor U3273 (N_3273,N_2785,N_2609);
xor U3274 (N_3274,N_2505,N_2587);
nor U3275 (N_3275,N_2580,N_2691);
xor U3276 (N_3276,N_2569,N_2870);
and U3277 (N_3277,N_2999,N_2937);
nor U3278 (N_3278,N_2696,N_2966);
xor U3279 (N_3279,N_2946,N_2596);
nand U3280 (N_3280,N_2768,N_2515);
nand U3281 (N_3281,N_2541,N_2713);
nor U3282 (N_3282,N_2686,N_2754);
and U3283 (N_3283,N_2509,N_2754);
nor U3284 (N_3284,N_2794,N_2868);
or U3285 (N_3285,N_2796,N_2584);
or U3286 (N_3286,N_2722,N_2718);
nor U3287 (N_3287,N_2700,N_2616);
and U3288 (N_3288,N_2699,N_2582);
nor U3289 (N_3289,N_2896,N_2542);
nand U3290 (N_3290,N_2858,N_2952);
or U3291 (N_3291,N_2581,N_2810);
xnor U3292 (N_3292,N_2943,N_2605);
and U3293 (N_3293,N_2577,N_2823);
xnor U3294 (N_3294,N_2726,N_2581);
xor U3295 (N_3295,N_2871,N_2750);
or U3296 (N_3296,N_2753,N_2651);
or U3297 (N_3297,N_2951,N_2787);
or U3298 (N_3298,N_2868,N_2813);
nor U3299 (N_3299,N_2952,N_2955);
nand U3300 (N_3300,N_2931,N_2525);
nand U3301 (N_3301,N_2528,N_2932);
and U3302 (N_3302,N_2997,N_2835);
and U3303 (N_3303,N_2718,N_2554);
nor U3304 (N_3304,N_2622,N_2916);
nor U3305 (N_3305,N_2995,N_2516);
and U3306 (N_3306,N_2675,N_2888);
and U3307 (N_3307,N_2785,N_2955);
nand U3308 (N_3308,N_2793,N_2518);
nor U3309 (N_3309,N_2601,N_2681);
or U3310 (N_3310,N_2555,N_2790);
nand U3311 (N_3311,N_2929,N_2917);
xor U3312 (N_3312,N_2664,N_2793);
xor U3313 (N_3313,N_2891,N_2622);
nor U3314 (N_3314,N_2715,N_2952);
or U3315 (N_3315,N_2889,N_2986);
xor U3316 (N_3316,N_2974,N_2510);
and U3317 (N_3317,N_2527,N_2520);
nor U3318 (N_3318,N_2772,N_2922);
or U3319 (N_3319,N_2864,N_2935);
or U3320 (N_3320,N_2530,N_2760);
nand U3321 (N_3321,N_2721,N_2881);
nor U3322 (N_3322,N_2668,N_2763);
nor U3323 (N_3323,N_2673,N_2993);
or U3324 (N_3324,N_2866,N_2718);
nor U3325 (N_3325,N_2668,N_2515);
nor U3326 (N_3326,N_2699,N_2709);
nand U3327 (N_3327,N_2504,N_2650);
nand U3328 (N_3328,N_2637,N_2521);
or U3329 (N_3329,N_2864,N_2896);
and U3330 (N_3330,N_2801,N_2535);
nor U3331 (N_3331,N_2888,N_2587);
nand U3332 (N_3332,N_2653,N_2907);
nor U3333 (N_3333,N_2685,N_2748);
nor U3334 (N_3334,N_2651,N_2837);
or U3335 (N_3335,N_2871,N_2973);
nand U3336 (N_3336,N_2965,N_2712);
or U3337 (N_3337,N_2842,N_2827);
and U3338 (N_3338,N_2511,N_2948);
or U3339 (N_3339,N_2786,N_2917);
or U3340 (N_3340,N_2520,N_2748);
nand U3341 (N_3341,N_2508,N_2604);
nand U3342 (N_3342,N_2531,N_2650);
and U3343 (N_3343,N_2936,N_2816);
or U3344 (N_3344,N_2919,N_2915);
xor U3345 (N_3345,N_2561,N_2798);
or U3346 (N_3346,N_2914,N_2879);
nor U3347 (N_3347,N_2600,N_2808);
nand U3348 (N_3348,N_2672,N_2640);
or U3349 (N_3349,N_2691,N_2546);
or U3350 (N_3350,N_2676,N_2937);
or U3351 (N_3351,N_2863,N_2754);
nand U3352 (N_3352,N_2692,N_2523);
nor U3353 (N_3353,N_2858,N_2891);
xor U3354 (N_3354,N_2923,N_2846);
and U3355 (N_3355,N_2689,N_2810);
nor U3356 (N_3356,N_2514,N_2669);
nor U3357 (N_3357,N_2943,N_2922);
nor U3358 (N_3358,N_2998,N_2677);
or U3359 (N_3359,N_2706,N_2582);
xor U3360 (N_3360,N_2576,N_2561);
xnor U3361 (N_3361,N_2510,N_2542);
nand U3362 (N_3362,N_2974,N_2828);
and U3363 (N_3363,N_2742,N_2948);
nand U3364 (N_3364,N_2665,N_2827);
nand U3365 (N_3365,N_2723,N_2758);
nand U3366 (N_3366,N_2595,N_2808);
and U3367 (N_3367,N_2722,N_2737);
nand U3368 (N_3368,N_2683,N_2874);
nor U3369 (N_3369,N_2951,N_2543);
or U3370 (N_3370,N_2585,N_2705);
or U3371 (N_3371,N_2612,N_2927);
nand U3372 (N_3372,N_2563,N_2703);
nand U3373 (N_3373,N_2681,N_2607);
nor U3374 (N_3374,N_2924,N_2522);
and U3375 (N_3375,N_2694,N_2730);
and U3376 (N_3376,N_2882,N_2854);
xor U3377 (N_3377,N_2693,N_2709);
and U3378 (N_3378,N_2940,N_2914);
nand U3379 (N_3379,N_2655,N_2700);
and U3380 (N_3380,N_2978,N_2779);
nand U3381 (N_3381,N_2541,N_2968);
xor U3382 (N_3382,N_2723,N_2559);
nor U3383 (N_3383,N_2595,N_2778);
nand U3384 (N_3384,N_2542,N_2697);
nand U3385 (N_3385,N_2693,N_2577);
or U3386 (N_3386,N_2668,N_2728);
nand U3387 (N_3387,N_2860,N_2605);
or U3388 (N_3388,N_2900,N_2787);
and U3389 (N_3389,N_2892,N_2693);
or U3390 (N_3390,N_2605,N_2982);
and U3391 (N_3391,N_2956,N_2587);
nor U3392 (N_3392,N_2706,N_2559);
nand U3393 (N_3393,N_2622,N_2856);
nand U3394 (N_3394,N_2701,N_2864);
nand U3395 (N_3395,N_2810,N_2786);
nor U3396 (N_3396,N_2752,N_2593);
and U3397 (N_3397,N_2812,N_2711);
and U3398 (N_3398,N_2574,N_2805);
nand U3399 (N_3399,N_2885,N_2700);
xor U3400 (N_3400,N_2584,N_2659);
nand U3401 (N_3401,N_2558,N_2813);
and U3402 (N_3402,N_2647,N_2735);
and U3403 (N_3403,N_2543,N_2554);
and U3404 (N_3404,N_2939,N_2569);
or U3405 (N_3405,N_2619,N_2868);
or U3406 (N_3406,N_2993,N_2632);
nand U3407 (N_3407,N_2761,N_2843);
or U3408 (N_3408,N_2564,N_2855);
or U3409 (N_3409,N_2970,N_2883);
xnor U3410 (N_3410,N_2604,N_2909);
or U3411 (N_3411,N_2982,N_2698);
or U3412 (N_3412,N_2644,N_2569);
nor U3413 (N_3413,N_2527,N_2608);
nor U3414 (N_3414,N_2818,N_2636);
xor U3415 (N_3415,N_2992,N_2634);
xor U3416 (N_3416,N_2557,N_2990);
nand U3417 (N_3417,N_2931,N_2605);
nor U3418 (N_3418,N_2823,N_2760);
and U3419 (N_3419,N_2862,N_2924);
or U3420 (N_3420,N_2982,N_2676);
nor U3421 (N_3421,N_2774,N_2944);
xor U3422 (N_3422,N_2571,N_2642);
xor U3423 (N_3423,N_2662,N_2984);
and U3424 (N_3424,N_2948,N_2777);
nand U3425 (N_3425,N_2834,N_2658);
or U3426 (N_3426,N_2884,N_2653);
nor U3427 (N_3427,N_2881,N_2888);
nand U3428 (N_3428,N_2665,N_2634);
nor U3429 (N_3429,N_2602,N_2654);
or U3430 (N_3430,N_2891,N_2740);
and U3431 (N_3431,N_2690,N_2663);
nor U3432 (N_3432,N_2877,N_2619);
nand U3433 (N_3433,N_2504,N_2714);
xor U3434 (N_3434,N_2865,N_2523);
nand U3435 (N_3435,N_2836,N_2808);
or U3436 (N_3436,N_2502,N_2988);
or U3437 (N_3437,N_2652,N_2600);
nor U3438 (N_3438,N_2985,N_2535);
or U3439 (N_3439,N_2664,N_2538);
and U3440 (N_3440,N_2826,N_2647);
or U3441 (N_3441,N_2807,N_2861);
nor U3442 (N_3442,N_2994,N_2769);
nor U3443 (N_3443,N_2568,N_2666);
or U3444 (N_3444,N_2910,N_2671);
nand U3445 (N_3445,N_2627,N_2588);
nor U3446 (N_3446,N_2950,N_2594);
nor U3447 (N_3447,N_2835,N_2596);
and U3448 (N_3448,N_2889,N_2645);
nor U3449 (N_3449,N_2670,N_2651);
and U3450 (N_3450,N_2607,N_2972);
nand U3451 (N_3451,N_2874,N_2761);
and U3452 (N_3452,N_2817,N_2949);
and U3453 (N_3453,N_2996,N_2857);
nor U3454 (N_3454,N_2848,N_2508);
xnor U3455 (N_3455,N_2566,N_2596);
or U3456 (N_3456,N_2546,N_2986);
nor U3457 (N_3457,N_2844,N_2588);
nand U3458 (N_3458,N_2968,N_2690);
nor U3459 (N_3459,N_2829,N_2603);
or U3460 (N_3460,N_2667,N_2735);
xnor U3461 (N_3461,N_2767,N_2998);
nand U3462 (N_3462,N_2562,N_2779);
or U3463 (N_3463,N_2853,N_2966);
nor U3464 (N_3464,N_2532,N_2888);
and U3465 (N_3465,N_2785,N_2564);
nand U3466 (N_3466,N_2743,N_2966);
and U3467 (N_3467,N_2661,N_2862);
nand U3468 (N_3468,N_2948,N_2539);
or U3469 (N_3469,N_2627,N_2863);
nand U3470 (N_3470,N_2732,N_2819);
xnor U3471 (N_3471,N_2847,N_2792);
nor U3472 (N_3472,N_2510,N_2788);
or U3473 (N_3473,N_2825,N_2925);
xor U3474 (N_3474,N_2723,N_2754);
nor U3475 (N_3475,N_2623,N_2680);
or U3476 (N_3476,N_2627,N_2842);
and U3477 (N_3477,N_2554,N_2972);
or U3478 (N_3478,N_2869,N_2777);
or U3479 (N_3479,N_2909,N_2847);
xor U3480 (N_3480,N_2659,N_2600);
and U3481 (N_3481,N_2813,N_2646);
and U3482 (N_3482,N_2867,N_2999);
or U3483 (N_3483,N_2781,N_2542);
nor U3484 (N_3484,N_2794,N_2749);
xor U3485 (N_3485,N_2601,N_2546);
or U3486 (N_3486,N_2884,N_2795);
or U3487 (N_3487,N_2768,N_2964);
nand U3488 (N_3488,N_2664,N_2910);
xnor U3489 (N_3489,N_2710,N_2777);
nand U3490 (N_3490,N_2942,N_2789);
xnor U3491 (N_3491,N_2675,N_2872);
nor U3492 (N_3492,N_2560,N_2599);
xnor U3493 (N_3493,N_2766,N_2982);
nand U3494 (N_3494,N_2750,N_2663);
xnor U3495 (N_3495,N_2625,N_2887);
nor U3496 (N_3496,N_2557,N_2946);
or U3497 (N_3497,N_2738,N_2510);
or U3498 (N_3498,N_2708,N_2672);
and U3499 (N_3499,N_2908,N_2649);
nand U3500 (N_3500,N_3128,N_3069);
nor U3501 (N_3501,N_3327,N_3169);
xnor U3502 (N_3502,N_3223,N_3314);
and U3503 (N_3503,N_3288,N_3489);
nor U3504 (N_3504,N_3221,N_3397);
nor U3505 (N_3505,N_3260,N_3036);
xnor U3506 (N_3506,N_3256,N_3152);
and U3507 (N_3507,N_3182,N_3303);
xor U3508 (N_3508,N_3264,N_3282);
and U3509 (N_3509,N_3173,N_3296);
nor U3510 (N_3510,N_3337,N_3029);
nor U3511 (N_3511,N_3410,N_3392);
nor U3512 (N_3512,N_3156,N_3484);
xnor U3513 (N_3513,N_3449,N_3079);
nor U3514 (N_3514,N_3185,N_3209);
and U3515 (N_3515,N_3460,N_3091);
nand U3516 (N_3516,N_3318,N_3432);
nand U3517 (N_3517,N_3174,N_3271);
nor U3518 (N_3518,N_3006,N_3428);
xor U3519 (N_3519,N_3019,N_3162);
nor U3520 (N_3520,N_3080,N_3194);
or U3521 (N_3521,N_3159,N_3382);
nor U3522 (N_3522,N_3160,N_3086);
and U3523 (N_3523,N_3468,N_3081);
or U3524 (N_3524,N_3283,N_3301);
and U3525 (N_3525,N_3110,N_3493);
and U3526 (N_3526,N_3299,N_3139);
nand U3527 (N_3527,N_3055,N_3202);
xor U3528 (N_3528,N_3144,N_3300);
nand U3529 (N_3529,N_3437,N_3100);
or U3530 (N_3530,N_3125,N_3157);
xor U3531 (N_3531,N_3431,N_3050);
or U3532 (N_3532,N_3088,N_3023);
nor U3533 (N_3533,N_3181,N_3092);
or U3534 (N_3534,N_3304,N_3328);
and U3535 (N_3535,N_3307,N_3113);
xor U3536 (N_3536,N_3012,N_3374);
nand U3537 (N_3537,N_3268,N_3298);
and U3538 (N_3538,N_3481,N_3045);
xor U3539 (N_3539,N_3232,N_3393);
or U3540 (N_3540,N_3040,N_3197);
xor U3541 (N_3541,N_3261,N_3380);
nand U3542 (N_3542,N_3241,N_3370);
nor U3543 (N_3543,N_3007,N_3022);
xor U3544 (N_3544,N_3373,N_3207);
and U3545 (N_3545,N_3341,N_3123);
nand U3546 (N_3546,N_3378,N_3132);
xnor U3547 (N_3547,N_3364,N_3124);
nand U3548 (N_3548,N_3490,N_3353);
nor U3549 (N_3549,N_3339,N_3039);
and U3550 (N_3550,N_3429,N_3073);
or U3551 (N_3551,N_3131,N_3010);
nand U3552 (N_3552,N_3320,N_3452);
nor U3553 (N_3553,N_3014,N_3458);
and U3554 (N_3554,N_3383,N_3058);
nand U3555 (N_3555,N_3367,N_3455);
nor U3556 (N_3556,N_3406,N_3401);
or U3557 (N_3557,N_3195,N_3136);
or U3558 (N_3558,N_3211,N_3099);
and U3559 (N_3559,N_3016,N_3361);
xnor U3560 (N_3560,N_3206,N_3056);
or U3561 (N_3561,N_3239,N_3352);
nor U3562 (N_3562,N_3179,N_3222);
and U3563 (N_3563,N_3254,N_3097);
nor U3564 (N_3564,N_3135,N_3008);
nand U3565 (N_3565,N_3400,N_3026);
nand U3566 (N_3566,N_3395,N_3281);
xor U3567 (N_3567,N_3321,N_3279);
xnor U3568 (N_3568,N_3426,N_3037);
and U3569 (N_3569,N_3018,N_3051);
xor U3570 (N_3570,N_3285,N_3054);
xnor U3571 (N_3571,N_3255,N_3001);
xor U3572 (N_3572,N_3457,N_3329);
nor U3573 (N_3573,N_3478,N_3453);
or U3574 (N_3574,N_3280,N_3137);
nor U3575 (N_3575,N_3423,N_3147);
and U3576 (N_3576,N_3448,N_3251);
and U3577 (N_3577,N_3002,N_3275);
nor U3578 (N_3578,N_3473,N_3388);
and U3579 (N_3579,N_3362,N_3356);
or U3580 (N_3580,N_3163,N_3068);
and U3581 (N_3581,N_3143,N_3053);
nand U3582 (N_3582,N_3138,N_3461);
or U3583 (N_3583,N_3035,N_3451);
or U3584 (N_3584,N_3496,N_3189);
or U3585 (N_3585,N_3020,N_3114);
nor U3586 (N_3586,N_3176,N_3440);
xnor U3587 (N_3587,N_3064,N_3272);
and U3588 (N_3588,N_3379,N_3442);
xnor U3589 (N_3589,N_3456,N_3387);
and U3590 (N_3590,N_3177,N_3161);
nor U3591 (N_3591,N_3192,N_3308);
and U3592 (N_3592,N_3474,N_3150);
and U3593 (N_3593,N_3077,N_3433);
nand U3594 (N_3594,N_3273,N_3404);
nor U3595 (N_3595,N_3096,N_3447);
or U3596 (N_3596,N_3263,N_3444);
or U3597 (N_3597,N_3258,N_3421);
nor U3598 (N_3598,N_3061,N_3483);
and U3599 (N_3599,N_3122,N_3398);
or U3600 (N_3600,N_3291,N_3316);
nand U3601 (N_3601,N_3032,N_3234);
nand U3602 (N_3602,N_3441,N_3278);
and U3603 (N_3603,N_3266,N_3435);
xor U3604 (N_3604,N_3305,N_3498);
or U3605 (N_3605,N_3365,N_3193);
nor U3606 (N_3606,N_3188,N_3306);
and U3607 (N_3607,N_3359,N_3215);
or U3608 (N_3608,N_3477,N_3067);
and U3609 (N_3609,N_3116,N_3425);
xor U3610 (N_3610,N_3357,N_3237);
and U3611 (N_3611,N_3171,N_3236);
or U3612 (N_3612,N_3322,N_3292);
and U3613 (N_3613,N_3411,N_3219);
or U3614 (N_3614,N_3063,N_3089);
nor U3615 (N_3615,N_3191,N_3470);
nor U3616 (N_3616,N_3253,N_3052);
nand U3617 (N_3617,N_3294,N_3065);
and U3618 (N_3618,N_3075,N_3025);
xnor U3619 (N_3619,N_3027,N_3409);
and U3620 (N_3620,N_3034,N_3118);
and U3621 (N_3621,N_3497,N_3252);
or U3622 (N_3622,N_3438,N_3366);
xor U3623 (N_3623,N_3491,N_3000);
nand U3624 (N_3624,N_3231,N_3480);
nand U3625 (N_3625,N_3347,N_3041);
xnor U3626 (N_3626,N_3047,N_3270);
nor U3627 (N_3627,N_3030,N_3333);
xnor U3628 (N_3628,N_3106,N_3021);
nor U3629 (N_3629,N_3345,N_3396);
or U3630 (N_3630,N_3024,N_3003);
or U3631 (N_3631,N_3229,N_3276);
nor U3632 (N_3632,N_3350,N_3004);
nand U3633 (N_3633,N_3059,N_3213);
nand U3634 (N_3634,N_3293,N_3355);
and U3635 (N_3635,N_3098,N_3459);
or U3636 (N_3636,N_3205,N_3319);
nand U3637 (N_3637,N_3057,N_3071);
nor U3638 (N_3638,N_3228,N_3471);
and U3639 (N_3639,N_3046,N_3145);
nand U3640 (N_3640,N_3129,N_3220);
and U3641 (N_3641,N_3094,N_3297);
nor U3642 (N_3642,N_3133,N_3416);
nand U3643 (N_3643,N_3492,N_3208);
nand U3644 (N_3644,N_3153,N_3408);
nand U3645 (N_3645,N_3107,N_3302);
nand U3646 (N_3646,N_3178,N_3149);
nor U3647 (N_3647,N_3127,N_3414);
or U3648 (N_3648,N_3164,N_3289);
or U3649 (N_3649,N_3464,N_3074);
or U3650 (N_3650,N_3115,N_3070);
nor U3651 (N_3651,N_3499,N_3117);
and U3652 (N_3652,N_3184,N_3267);
nand U3653 (N_3653,N_3033,N_3265);
xor U3654 (N_3654,N_3072,N_3101);
xnor U3655 (N_3655,N_3436,N_3485);
nor U3656 (N_3656,N_3463,N_3028);
nand U3657 (N_3657,N_3286,N_3227);
and U3658 (N_3658,N_3167,N_3204);
nand U3659 (N_3659,N_3405,N_3242);
nand U3660 (N_3660,N_3082,N_3472);
or U3661 (N_3661,N_3317,N_3412);
xor U3662 (N_3662,N_3257,N_3439);
or U3663 (N_3663,N_3338,N_3476);
nor U3664 (N_3664,N_3119,N_3391);
nor U3665 (N_3665,N_3358,N_3332);
nor U3666 (N_3666,N_3418,N_3262);
nor U3667 (N_3667,N_3134,N_3172);
nand U3668 (N_3668,N_3375,N_3402);
or U3669 (N_3669,N_3465,N_3415);
or U3670 (N_3670,N_3372,N_3462);
nand U3671 (N_3671,N_3313,N_3335);
xor U3672 (N_3672,N_3377,N_3331);
nor U3673 (N_3673,N_3390,N_3446);
nand U3674 (N_3674,N_3422,N_3290);
xnor U3675 (N_3675,N_3469,N_3102);
and U3676 (N_3676,N_3200,N_3407);
xor U3677 (N_3677,N_3454,N_3495);
and U3678 (N_3678,N_3371,N_3486);
xor U3679 (N_3679,N_3269,N_3225);
nor U3680 (N_3680,N_3015,N_3198);
or U3681 (N_3681,N_3005,N_3140);
nand U3682 (N_3682,N_3203,N_3038);
and U3683 (N_3683,N_3354,N_3247);
and U3684 (N_3684,N_3363,N_3466);
xnor U3685 (N_3685,N_3434,N_3103);
and U3686 (N_3686,N_3450,N_3336);
or U3687 (N_3687,N_3168,N_3233);
and U3688 (N_3688,N_3130,N_3017);
and U3689 (N_3689,N_3243,N_3111);
or U3690 (N_3690,N_3180,N_3230);
nor U3691 (N_3691,N_3467,N_3403);
or U3692 (N_3692,N_3166,N_3245);
xor U3693 (N_3693,N_3310,N_3226);
nor U3694 (N_3694,N_3494,N_3043);
xnor U3695 (N_3695,N_3482,N_3344);
or U3696 (N_3696,N_3044,N_3093);
and U3697 (N_3697,N_3218,N_3413);
nor U3698 (N_3698,N_3108,N_3346);
xor U3699 (N_3699,N_3384,N_3274);
xnor U3700 (N_3700,N_3284,N_3295);
or U3701 (N_3701,N_3155,N_3210);
nor U3702 (N_3702,N_3196,N_3095);
and U3703 (N_3703,N_3201,N_3151);
nand U3704 (N_3704,N_3084,N_3424);
nand U3705 (N_3705,N_3175,N_3386);
or U3706 (N_3706,N_3190,N_3249);
or U3707 (N_3707,N_3121,N_3090);
nor U3708 (N_3708,N_3430,N_3287);
or U3709 (N_3709,N_3488,N_3158);
xnor U3710 (N_3710,N_3238,N_3312);
and U3711 (N_3711,N_3348,N_3146);
or U3712 (N_3712,N_3487,N_3154);
nor U3713 (N_3713,N_3076,N_3479);
nand U3714 (N_3714,N_3148,N_3186);
xor U3715 (N_3715,N_3011,N_3031);
and U3716 (N_3716,N_3325,N_3351);
or U3717 (N_3717,N_3246,N_3248);
nor U3718 (N_3718,N_3235,N_3126);
nor U3719 (N_3719,N_3214,N_3066);
nor U3720 (N_3720,N_3427,N_3087);
xor U3721 (N_3721,N_3109,N_3078);
or U3722 (N_3722,N_3323,N_3112);
nand U3723 (N_3723,N_3217,N_3083);
nor U3724 (N_3724,N_3187,N_3105);
nor U3725 (N_3725,N_3376,N_3340);
xor U3726 (N_3726,N_3049,N_3334);
and U3727 (N_3727,N_3385,N_3165);
nor U3728 (N_3728,N_3342,N_3060);
xnor U3729 (N_3729,N_3216,N_3224);
or U3730 (N_3730,N_3311,N_3240);
and U3731 (N_3731,N_3062,N_3399);
nor U3732 (N_3732,N_3259,N_3183);
nand U3733 (N_3733,N_3042,N_3212);
or U3734 (N_3734,N_3475,N_3085);
nand U3735 (N_3735,N_3369,N_3445);
and U3736 (N_3736,N_3048,N_3104);
nand U3737 (N_3737,N_3309,N_3417);
nor U3738 (N_3738,N_3170,N_3326);
xor U3739 (N_3739,N_3009,N_3343);
nor U3740 (N_3740,N_3315,N_3420);
or U3741 (N_3741,N_3244,N_3443);
nor U3742 (N_3742,N_3141,N_3330);
or U3743 (N_3743,N_3349,N_3324);
nor U3744 (N_3744,N_3368,N_3389);
or U3745 (N_3745,N_3120,N_3394);
nor U3746 (N_3746,N_3381,N_3277);
and U3747 (N_3747,N_3013,N_3142);
nand U3748 (N_3748,N_3250,N_3419);
nand U3749 (N_3749,N_3199,N_3360);
xnor U3750 (N_3750,N_3364,N_3302);
nand U3751 (N_3751,N_3337,N_3330);
nand U3752 (N_3752,N_3284,N_3246);
and U3753 (N_3753,N_3229,N_3323);
nor U3754 (N_3754,N_3011,N_3050);
xor U3755 (N_3755,N_3100,N_3390);
and U3756 (N_3756,N_3323,N_3018);
nand U3757 (N_3757,N_3290,N_3002);
nor U3758 (N_3758,N_3033,N_3196);
and U3759 (N_3759,N_3426,N_3407);
nand U3760 (N_3760,N_3323,N_3086);
nor U3761 (N_3761,N_3441,N_3150);
and U3762 (N_3762,N_3210,N_3467);
or U3763 (N_3763,N_3185,N_3289);
nor U3764 (N_3764,N_3264,N_3329);
or U3765 (N_3765,N_3314,N_3336);
xor U3766 (N_3766,N_3357,N_3128);
or U3767 (N_3767,N_3286,N_3061);
and U3768 (N_3768,N_3308,N_3477);
xnor U3769 (N_3769,N_3400,N_3153);
and U3770 (N_3770,N_3295,N_3338);
and U3771 (N_3771,N_3133,N_3358);
and U3772 (N_3772,N_3306,N_3173);
or U3773 (N_3773,N_3260,N_3085);
or U3774 (N_3774,N_3187,N_3488);
nand U3775 (N_3775,N_3239,N_3055);
nand U3776 (N_3776,N_3261,N_3195);
and U3777 (N_3777,N_3464,N_3270);
and U3778 (N_3778,N_3313,N_3444);
xor U3779 (N_3779,N_3070,N_3036);
nor U3780 (N_3780,N_3314,N_3164);
xor U3781 (N_3781,N_3223,N_3229);
nand U3782 (N_3782,N_3457,N_3165);
or U3783 (N_3783,N_3108,N_3400);
xor U3784 (N_3784,N_3253,N_3051);
or U3785 (N_3785,N_3482,N_3341);
nand U3786 (N_3786,N_3166,N_3318);
or U3787 (N_3787,N_3377,N_3314);
nor U3788 (N_3788,N_3484,N_3056);
or U3789 (N_3789,N_3450,N_3056);
nand U3790 (N_3790,N_3270,N_3474);
nand U3791 (N_3791,N_3492,N_3011);
nor U3792 (N_3792,N_3041,N_3139);
nor U3793 (N_3793,N_3100,N_3487);
xor U3794 (N_3794,N_3471,N_3248);
and U3795 (N_3795,N_3270,N_3428);
and U3796 (N_3796,N_3392,N_3403);
xnor U3797 (N_3797,N_3044,N_3404);
xnor U3798 (N_3798,N_3353,N_3217);
xor U3799 (N_3799,N_3178,N_3461);
or U3800 (N_3800,N_3310,N_3258);
xnor U3801 (N_3801,N_3047,N_3220);
xor U3802 (N_3802,N_3073,N_3489);
and U3803 (N_3803,N_3077,N_3253);
nor U3804 (N_3804,N_3389,N_3125);
or U3805 (N_3805,N_3365,N_3102);
nand U3806 (N_3806,N_3175,N_3373);
nand U3807 (N_3807,N_3235,N_3318);
or U3808 (N_3808,N_3421,N_3133);
or U3809 (N_3809,N_3088,N_3086);
nor U3810 (N_3810,N_3368,N_3371);
xnor U3811 (N_3811,N_3019,N_3214);
xor U3812 (N_3812,N_3323,N_3266);
and U3813 (N_3813,N_3404,N_3200);
nand U3814 (N_3814,N_3177,N_3050);
xnor U3815 (N_3815,N_3175,N_3274);
and U3816 (N_3816,N_3172,N_3145);
nand U3817 (N_3817,N_3383,N_3030);
or U3818 (N_3818,N_3259,N_3012);
or U3819 (N_3819,N_3084,N_3011);
and U3820 (N_3820,N_3087,N_3052);
nor U3821 (N_3821,N_3410,N_3464);
xor U3822 (N_3822,N_3294,N_3429);
or U3823 (N_3823,N_3391,N_3312);
and U3824 (N_3824,N_3346,N_3275);
or U3825 (N_3825,N_3401,N_3099);
nand U3826 (N_3826,N_3413,N_3205);
xnor U3827 (N_3827,N_3340,N_3261);
and U3828 (N_3828,N_3465,N_3136);
or U3829 (N_3829,N_3303,N_3348);
nand U3830 (N_3830,N_3344,N_3090);
nand U3831 (N_3831,N_3107,N_3321);
nand U3832 (N_3832,N_3229,N_3356);
xnor U3833 (N_3833,N_3213,N_3436);
or U3834 (N_3834,N_3232,N_3469);
or U3835 (N_3835,N_3120,N_3300);
nor U3836 (N_3836,N_3160,N_3078);
nor U3837 (N_3837,N_3055,N_3021);
xnor U3838 (N_3838,N_3360,N_3212);
and U3839 (N_3839,N_3241,N_3069);
nand U3840 (N_3840,N_3200,N_3248);
nor U3841 (N_3841,N_3069,N_3346);
xnor U3842 (N_3842,N_3031,N_3306);
nor U3843 (N_3843,N_3088,N_3064);
xor U3844 (N_3844,N_3082,N_3390);
nor U3845 (N_3845,N_3439,N_3248);
nand U3846 (N_3846,N_3136,N_3249);
and U3847 (N_3847,N_3045,N_3348);
nor U3848 (N_3848,N_3088,N_3267);
and U3849 (N_3849,N_3209,N_3154);
and U3850 (N_3850,N_3359,N_3256);
or U3851 (N_3851,N_3101,N_3326);
xor U3852 (N_3852,N_3442,N_3155);
or U3853 (N_3853,N_3101,N_3208);
xnor U3854 (N_3854,N_3428,N_3416);
and U3855 (N_3855,N_3249,N_3139);
or U3856 (N_3856,N_3107,N_3080);
or U3857 (N_3857,N_3243,N_3385);
nand U3858 (N_3858,N_3384,N_3006);
or U3859 (N_3859,N_3154,N_3024);
nor U3860 (N_3860,N_3402,N_3073);
and U3861 (N_3861,N_3050,N_3015);
nand U3862 (N_3862,N_3352,N_3070);
and U3863 (N_3863,N_3145,N_3444);
nor U3864 (N_3864,N_3333,N_3410);
nand U3865 (N_3865,N_3117,N_3414);
or U3866 (N_3866,N_3276,N_3327);
nand U3867 (N_3867,N_3156,N_3312);
nand U3868 (N_3868,N_3273,N_3127);
xor U3869 (N_3869,N_3431,N_3315);
nand U3870 (N_3870,N_3434,N_3195);
nand U3871 (N_3871,N_3260,N_3197);
and U3872 (N_3872,N_3363,N_3272);
nand U3873 (N_3873,N_3405,N_3108);
nand U3874 (N_3874,N_3010,N_3479);
and U3875 (N_3875,N_3221,N_3121);
nand U3876 (N_3876,N_3344,N_3048);
nand U3877 (N_3877,N_3258,N_3264);
and U3878 (N_3878,N_3461,N_3002);
and U3879 (N_3879,N_3427,N_3481);
and U3880 (N_3880,N_3116,N_3292);
nor U3881 (N_3881,N_3094,N_3174);
nand U3882 (N_3882,N_3165,N_3243);
xor U3883 (N_3883,N_3479,N_3077);
and U3884 (N_3884,N_3178,N_3284);
nand U3885 (N_3885,N_3318,N_3273);
xor U3886 (N_3886,N_3121,N_3261);
nand U3887 (N_3887,N_3424,N_3126);
nor U3888 (N_3888,N_3485,N_3272);
and U3889 (N_3889,N_3394,N_3323);
nor U3890 (N_3890,N_3321,N_3471);
and U3891 (N_3891,N_3239,N_3006);
nand U3892 (N_3892,N_3244,N_3232);
and U3893 (N_3893,N_3184,N_3043);
and U3894 (N_3894,N_3059,N_3010);
nor U3895 (N_3895,N_3169,N_3336);
xnor U3896 (N_3896,N_3367,N_3161);
nand U3897 (N_3897,N_3113,N_3050);
and U3898 (N_3898,N_3499,N_3336);
or U3899 (N_3899,N_3339,N_3236);
nor U3900 (N_3900,N_3499,N_3233);
nand U3901 (N_3901,N_3405,N_3058);
or U3902 (N_3902,N_3123,N_3202);
nand U3903 (N_3903,N_3139,N_3496);
nand U3904 (N_3904,N_3439,N_3075);
nand U3905 (N_3905,N_3472,N_3449);
and U3906 (N_3906,N_3010,N_3195);
nand U3907 (N_3907,N_3469,N_3476);
nand U3908 (N_3908,N_3342,N_3025);
and U3909 (N_3909,N_3218,N_3314);
and U3910 (N_3910,N_3206,N_3227);
or U3911 (N_3911,N_3384,N_3292);
nand U3912 (N_3912,N_3013,N_3377);
xnor U3913 (N_3913,N_3420,N_3163);
xor U3914 (N_3914,N_3154,N_3176);
or U3915 (N_3915,N_3171,N_3198);
and U3916 (N_3916,N_3366,N_3224);
nand U3917 (N_3917,N_3330,N_3278);
nand U3918 (N_3918,N_3381,N_3294);
xnor U3919 (N_3919,N_3180,N_3123);
or U3920 (N_3920,N_3186,N_3307);
nor U3921 (N_3921,N_3233,N_3492);
nor U3922 (N_3922,N_3246,N_3444);
xor U3923 (N_3923,N_3363,N_3220);
or U3924 (N_3924,N_3255,N_3263);
xnor U3925 (N_3925,N_3117,N_3140);
xnor U3926 (N_3926,N_3388,N_3237);
xor U3927 (N_3927,N_3483,N_3490);
nand U3928 (N_3928,N_3300,N_3389);
xnor U3929 (N_3929,N_3080,N_3444);
xnor U3930 (N_3930,N_3399,N_3413);
or U3931 (N_3931,N_3052,N_3035);
and U3932 (N_3932,N_3237,N_3380);
or U3933 (N_3933,N_3112,N_3405);
and U3934 (N_3934,N_3031,N_3049);
nor U3935 (N_3935,N_3229,N_3445);
nand U3936 (N_3936,N_3352,N_3080);
nor U3937 (N_3937,N_3421,N_3047);
nor U3938 (N_3938,N_3468,N_3110);
or U3939 (N_3939,N_3384,N_3141);
nand U3940 (N_3940,N_3372,N_3023);
xnor U3941 (N_3941,N_3016,N_3007);
or U3942 (N_3942,N_3117,N_3325);
or U3943 (N_3943,N_3191,N_3478);
nand U3944 (N_3944,N_3499,N_3382);
xnor U3945 (N_3945,N_3078,N_3008);
and U3946 (N_3946,N_3446,N_3144);
xor U3947 (N_3947,N_3499,N_3320);
or U3948 (N_3948,N_3265,N_3235);
nand U3949 (N_3949,N_3145,N_3169);
and U3950 (N_3950,N_3143,N_3082);
or U3951 (N_3951,N_3028,N_3298);
and U3952 (N_3952,N_3119,N_3172);
or U3953 (N_3953,N_3074,N_3191);
nor U3954 (N_3954,N_3334,N_3283);
or U3955 (N_3955,N_3416,N_3267);
and U3956 (N_3956,N_3176,N_3088);
xor U3957 (N_3957,N_3353,N_3165);
xor U3958 (N_3958,N_3089,N_3362);
nor U3959 (N_3959,N_3045,N_3450);
nand U3960 (N_3960,N_3417,N_3117);
or U3961 (N_3961,N_3144,N_3487);
xnor U3962 (N_3962,N_3420,N_3129);
or U3963 (N_3963,N_3343,N_3205);
and U3964 (N_3964,N_3368,N_3330);
nor U3965 (N_3965,N_3054,N_3243);
or U3966 (N_3966,N_3304,N_3092);
nand U3967 (N_3967,N_3164,N_3130);
and U3968 (N_3968,N_3277,N_3315);
nor U3969 (N_3969,N_3288,N_3442);
nand U3970 (N_3970,N_3160,N_3011);
and U3971 (N_3971,N_3442,N_3293);
nand U3972 (N_3972,N_3039,N_3242);
and U3973 (N_3973,N_3226,N_3384);
xor U3974 (N_3974,N_3116,N_3366);
or U3975 (N_3975,N_3074,N_3272);
nor U3976 (N_3976,N_3409,N_3127);
or U3977 (N_3977,N_3136,N_3448);
and U3978 (N_3978,N_3372,N_3376);
and U3979 (N_3979,N_3090,N_3146);
and U3980 (N_3980,N_3231,N_3308);
xor U3981 (N_3981,N_3055,N_3073);
nand U3982 (N_3982,N_3240,N_3107);
xor U3983 (N_3983,N_3487,N_3394);
xnor U3984 (N_3984,N_3408,N_3025);
nor U3985 (N_3985,N_3369,N_3166);
xnor U3986 (N_3986,N_3122,N_3138);
or U3987 (N_3987,N_3169,N_3107);
xnor U3988 (N_3988,N_3465,N_3247);
xor U3989 (N_3989,N_3206,N_3172);
nand U3990 (N_3990,N_3488,N_3264);
or U3991 (N_3991,N_3106,N_3469);
nand U3992 (N_3992,N_3166,N_3014);
or U3993 (N_3993,N_3470,N_3004);
or U3994 (N_3994,N_3396,N_3287);
nand U3995 (N_3995,N_3220,N_3415);
and U3996 (N_3996,N_3096,N_3188);
nor U3997 (N_3997,N_3064,N_3469);
nand U3998 (N_3998,N_3388,N_3231);
and U3999 (N_3999,N_3200,N_3362);
nand U4000 (N_4000,N_3522,N_3925);
xor U4001 (N_4001,N_3658,N_3962);
and U4002 (N_4002,N_3995,N_3849);
and U4003 (N_4003,N_3991,N_3570);
or U4004 (N_4004,N_3538,N_3690);
or U4005 (N_4005,N_3847,N_3916);
xor U4006 (N_4006,N_3556,N_3567);
nand U4007 (N_4007,N_3561,N_3784);
or U4008 (N_4008,N_3766,N_3646);
and U4009 (N_4009,N_3754,N_3516);
and U4010 (N_4010,N_3968,N_3949);
and U4011 (N_4011,N_3665,N_3612);
nand U4012 (N_4012,N_3909,N_3714);
nand U4013 (N_4013,N_3560,N_3929);
or U4014 (N_4014,N_3677,N_3871);
xnor U4015 (N_4015,N_3844,N_3793);
and U4016 (N_4016,N_3700,N_3912);
nand U4017 (N_4017,N_3777,N_3720);
nand U4018 (N_4018,N_3530,N_3748);
nand U4019 (N_4019,N_3926,N_3892);
xnor U4020 (N_4020,N_3838,N_3649);
nand U4021 (N_4021,N_3662,N_3708);
xnor U4022 (N_4022,N_3947,N_3903);
nand U4023 (N_4023,N_3952,N_3577);
xnor U4024 (N_4024,N_3756,N_3502);
or U4025 (N_4025,N_3951,N_3999);
xor U4026 (N_4026,N_3632,N_3536);
or U4027 (N_4027,N_3590,N_3686);
or U4028 (N_4028,N_3548,N_3666);
nand U4029 (N_4029,N_3563,N_3940);
and U4030 (N_4030,N_3997,N_3965);
nand U4031 (N_4031,N_3939,N_3505);
nor U4032 (N_4032,N_3687,N_3703);
xnor U4033 (N_4033,N_3851,N_3723);
nand U4034 (N_4034,N_3931,N_3582);
nor U4035 (N_4035,N_3622,N_3834);
nand U4036 (N_4036,N_3616,N_3858);
nand U4037 (N_4037,N_3565,N_3865);
or U4038 (N_4038,N_3963,N_3906);
or U4039 (N_4039,N_3883,N_3924);
or U4040 (N_4040,N_3990,N_3675);
nand U4041 (N_4041,N_3866,N_3895);
and U4042 (N_4042,N_3500,N_3759);
nand U4043 (N_4043,N_3648,N_3518);
nor U4044 (N_4044,N_3730,N_3989);
nand U4045 (N_4045,N_3633,N_3890);
or U4046 (N_4046,N_3814,N_3606);
nor U4047 (N_4047,N_3569,N_3812);
nand U4048 (N_4048,N_3868,N_3881);
and U4049 (N_4049,N_3957,N_3694);
nor U4050 (N_4050,N_3550,N_3899);
nand U4051 (N_4051,N_3765,N_3992);
nor U4052 (N_4052,N_3613,N_3840);
xnor U4053 (N_4053,N_3525,N_3634);
nor U4054 (N_4054,N_3880,N_3535);
nand U4055 (N_4055,N_3531,N_3933);
nand U4056 (N_4056,N_3555,N_3807);
xnor U4057 (N_4057,N_3791,N_3600);
or U4058 (N_4058,N_3914,N_3678);
xnor U4059 (N_4059,N_3994,N_3578);
xnor U4060 (N_4060,N_3543,N_3679);
and U4061 (N_4061,N_3620,N_3710);
nand U4062 (N_4062,N_3534,N_3636);
nor U4063 (N_4063,N_3693,N_3943);
xor U4064 (N_4064,N_3734,N_3819);
nand U4065 (N_4065,N_3755,N_3950);
xnor U4066 (N_4066,N_3749,N_3904);
nor U4067 (N_4067,N_3668,N_3961);
nand U4068 (N_4068,N_3571,N_3659);
or U4069 (N_4069,N_3798,N_3732);
xnor U4070 (N_4070,N_3850,N_3683);
and U4071 (N_4071,N_3719,N_3935);
nand U4072 (N_4072,N_3862,N_3878);
nor U4073 (N_4073,N_3542,N_3780);
xor U4074 (N_4074,N_3757,N_3581);
or U4075 (N_4075,N_3855,N_3729);
nand U4076 (N_4076,N_3592,N_3964);
xnor U4077 (N_4077,N_3815,N_3827);
and U4078 (N_4078,N_3831,N_3523);
nor U4079 (N_4079,N_3911,N_3680);
and U4080 (N_4080,N_3512,N_3857);
nor U4081 (N_4081,N_3510,N_3617);
xor U4082 (N_4082,N_3846,N_3872);
or U4083 (N_4083,N_3586,N_3809);
xor U4084 (N_4084,N_3603,N_3789);
or U4085 (N_4085,N_3795,N_3764);
nand U4086 (N_4086,N_3650,N_3702);
or U4087 (N_4087,N_3837,N_3737);
nand U4088 (N_4088,N_3938,N_3721);
nand U4089 (N_4089,N_3547,N_3768);
nor U4090 (N_4090,N_3651,N_3958);
nor U4091 (N_4091,N_3882,N_3697);
xor U4092 (N_4092,N_3704,N_3937);
nor U4093 (N_4093,N_3978,N_3724);
nand U4094 (N_4094,N_3954,N_3656);
xor U4095 (N_4095,N_3948,N_3967);
nor U4096 (N_4096,N_3551,N_3705);
nor U4097 (N_4097,N_3922,N_3830);
nor U4098 (N_4098,N_3836,N_3741);
nor U4099 (N_4099,N_3716,N_3736);
and U4100 (N_4100,N_3514,N_3879);
xor U4101 (N_4101,N_3923,N_3982);
and U4102 (N_4102,N_3977,N_3682);
nand U4103 (N_4103,N_3905,N_3744);
nand U4104 (N_4104,N_3860,N_3552);
and U4105 (N_4105,N_3685,N_3944);
xnor U4106 (N_4106,N_3739,N_3828);
nor U4107 (N_4107,N_3568,N_3527);
nor U4108 (N_4108,N_3804,N_3504);
xor U4109 (N_4109,N_3747,N_3753);
xor U4110 (N_4110,N_3718,N_3971);
nand U4111 (N_4111,N_3618,N_3652);
nor U4112 (N_4112,N_3645,N_3605);
nor U4113 (N_4113,N_3631,N_3790);
and U4114 (N_4114,N_3526,N_3657);
nor U4115 (N_4115,N_3821,N_3886);
or U4116 (N_4116,N_3654,N_3508);
or U4117 (N_4117,N_3558,N_3667);
nand U4118 (N_4118,N_3774,N_3996);
xor U4119 (N_4119,N_3772,N_3663);
nand U4120 (N_4120,N_3509,N_3698);
nor U4121 (N_4121,N_3779,N_3712);
or U4122 (N_4122,N_3801,N_3873);
or U4123 (N_4123,N_3524,N_3727);
nor U4124 (N_4124,N_3853,N_3671);
or U4125 (N_4125,N_3826,N_3845);
and U4126 (N_4126,N_3520,N_3579);
and U4127 (N_4127,N_3921,N_3988);
xnor U4128 (N_4128,N_3945,N_3588);
or U4129 (N_4129,N_3630,N_3559);
xnor U4130 (N_4130,N_3792,N_3614);
nand U4131 (N_4131,N_3597,N_3981);
xnor U4132 (N_4132,N_3876,N_3896);
nand U4133 (N_4133,N_3684,N_3993);
xor U4134 (N_4134,N_3595,N_3781);
or U4135 (N_4135,N_3507,N_3628);
nor U4136 (N_4136,N_3908,N_3515);
and U4137 (N_4137,N_3701,N_3717);
xnor U4138 (N_4138,N_3713,N_3893);
nor U4139 (N_4139,N_3998,N_3856);
nor U4140 (N_4140,N_3841,N_3824);
or U4141 (N_4141,N_3915,N_3692);
xor U4142 (N_4142,N_3927,N_3803);
nand U4143 (N_4143,N_3611,N_3574);
xor U4144 (N_4144,N_3517,N_3762);
or U4145 (N_4145,N_3820,N_3788);
and U4146 (N_4146,N_3805,N_3740);
and U4147 (N_4147,N_3533,N_3709);
nand U4148 (N_4148,N_3771,N_3623);
nand U4149 (N_4149,N_3553,N_3775);
nor U4150 (N_4150,N_3624,N_3959);
xnor U4151 (N_4151,N_3859,N_3575);
nand U4152 (N_4152,N_3738,N_3707);
xor U4153 (N_4153,N_3573,N_3681);
xor U4154 (N_4154,N_3842,N_3576);
nor U4155 (N_4155,N_3975,N_3731);
nand U4156 (N_4156,N_3888,N_3673);
and U4157 (N_4157,N_3742,N_3875);
xor U4158 (N_4158,N_3802,N_3797);
and U4159 (N_4159,N_3691,N_3786);
or U4160 (N_4160,N_3832,N_3810);
xnor U4161 (N_4161,N_3825,N_3867);
nand U4162 (N_4162,N_3580,N_3806);
nand U4163 (N_4163,N_3621,N_3885);
nand U4164 (N_4164,N_3767,N_3848);
or U4165 (N_4165,N_3672,N_3593);
xor U4166 (N_4166,N_3557,N_3918);
xor U4167 (N_4167,N_3609,N_3979);
and U4168 (N_4168,N_3726,N_3778);
xnor U4169 (N_4169,N_3639,N_3589);
or U4170 (N_4170,N_3884,N_3974);
or U4171 (N_4171,N_3970,N_3562);
nand U4172 (N_4172,N_3539,N_3808);
nand U4173 (N_4173,N_3554,N_3537);
or U4174 (N_4174,N_3907,N_3604);
and U4175 (N_4175,N_3919,N_3644);
nor U4176 (N_4176,N_3769,N_3549);
nor U4177 (N_4177,N_3898,N_3902);
nand U4178 (N_4178,N_3887,N_3607);
nand U4179 (N_4179,N_3642,N_3894);
nor U4180 (N_4180,N_3913,N_3513);
and U4181 (N_4181,N_3799,N_3540);
nor U4182 (N_4182,N_3936,N_3584);
and U4183 (N_4183,N_3751,N_3591);
nor U4184 (N_4184,N_3521,N_3980);
nand U4185 (N_4185,N_3752,N_3889);
or U4186 (N_4186,N_3598,N_3863);
nor U4187 (N_4187,N_3966,N_3643);
nor U4188 (N_4188,N_3528,N_3969);
nand U4189 (N_4189,N_3897,N_3901);
or U4190 (N_4190,N_3546,N_3758);
xnor U4191 (N_4191,N_3688,N_3506);
and U4192 (N_4192,N_3647,N_3874);
xor U4193 (N_4193,N_3869,N_3545);
xnor U4194 (N_4194,N_3699,N_3635);
nand U4195 (N_4195,N_3532,N_3900);
nand U4196 (N_4196,N_3760,N_3669);
and U4197 (N_4197,N_3861,N_3956);
or U4198 (N_4198,N_3987,N_3572);
nor U4199 (N_4199,N_3641,N_3930);
nor U4200 (N_4200,N_3785,N_3519);
nand U4201 (N_4201,N_3664,N_3796);
nand U4202 (N_4202,N_3782,N_3776);
nor U4203 (N_4203,N_3615,N_3529);
xnor U4204 (N_4204,N_3670,N_3816);
nor U4205 (N_4205,N_3829,N_3715);
xor U4206 (N_4206,N_3722,N_3676);
or U4207 (N_4207,N_3864,N_3750);
and U4208 (N_4208,N_3627,N_3783);
xnor U4209 (N_4209,N_3610,N_3544);
nand U4210 (N_4210,N_3696,N_3583);
or U4211 (N_4211,N_3852,N_3833);
xnor U4212 (N_4212,N_3728,N_3835);
nand U4213 (N_4213,N_3955,N_3800);
and U4214 (N_4214,N_3920,N_3746);
nand U4215 (N_4215,N_3501,N_3934);
or U4216 (N_4216,N_3960,N_3566);
xnor U4217 (N_4217,N_3745,N_3695);
xnor U4218 (N_4218,N_3711,N_3910);
or U4219 (N_4219,N_3811,N_3985);
xnor U4220 (N_4220,N_3794,N_3770);
or U4221 (N_4221,N_3823,N_3870);
nor U4222 (N_4222,N_3735,N_3655);
xnor U4223 (N_4223,N_3773,N_3511);
nor U4224 (N_4224,N_3733,N_3976);
xor U4225 (N_4225,N_3585,N_3629);
nor U4226 (N_4226,N_3594,N_3596);
and U4227 (N_4227,N_3608,N_3601);
nand U4228 (N_4228,N_3660,N_3653);
and U4229 (N_4229,N_3986,N_3689);
nor U4230 (N_4230,N_3928,N_3972);
or U4231 (N_4231,N_3599,N_3674);
or U4232 (N_4232,N_3725,N_3640);
nor U4233 (N_4233,N_3932,N_3743);
nand U4234 (N_4234,N_3941,N_3787);
nand U4235 (N_4235,N_3619,N_3839);
or U4236 (N_4236,N_3761,N_3953);
and U4237 (N_4237,N_3877,N_3843);
nor U4238 (N_4238,N_3942,N_3817);
nor U4239 (N_4239,N_3503,N_3661);
xor U4240 (N_4240,N_3637,N_3626);
nor U4241 (N_4241,N_3602,N_3625);
and U4242 (N_4242,N_3822,N_3983);
and U4243 (N_4243,N_3564,N_3984);
or U4244 (N_4244,N_3854,N_3818);
and U4245 (N_4245,N_3973,N_3917);
nand U4246 (N_4246,N_3541,N_3813);
and U4247 (N_4247,N_3706,N_3763);
nor U4248 (N_4248,N_3638,N_3891);
nor U4249 (N_4249,N_3587,N_3946);
nor U4250 (N_4250,N_3744,N_3635);
and U4251 (N_4251,N_3653,N_3646);
xor U4252 (N_4252,N_3899,N_3788);
xnor U4253 (N_4253,N_3867,N_3667);
nand U4254 (N_4254,N_3788,N_3735);
or U4255 (N_4255,N_3750,N_3968);
nand U4256 (N_4256,N_3745,N_3889);
and U4257 (N_4257,N_3828,N_3721);
xor U4258 (N_4258,N_3676,N_3980);
or U4259 (N_4259,N_3530,N_3616);
nor U4260 (N_4260,N_3727,N_3676);
and U4261 (N_4261,N_3971,N_3901);
nor U4262 (N_4262,N_3631,N_3731);
and U4263 (N_4263,N_3825,N_3868);
nor U4264 (N_4264,N_3956,N_3942);
xor U4265 (N_4265,N_3679,N_3514);
nor U4266 (N_4266,N_3813,N_3680);
and U4267 (N_4267,N_3905,N_3523);
nor U4268 (N_4268,N_3647,N_3753);
nand U4269 (N_4269,N_3658,N_3818);
and U4270 (N_4270,N_3982,N_3526);
or U4271 (N_4271,N_3677,N_3845);
xor U4272 (N_4272,N_3950,N_3824);
or U4273 (N_4273,N_3573,N_3801);
nor U4274 (N_4274,N_3580,N_3630);
and U4275 (N_4275,N_3952,N_3967);
nand U4276 (N_4276,N_3737,N_3666);
or U4277 (N_4277,N_3507,N_3928);
xnor U4278 (N_4278,N_3615,N_3967);
or U4279 (N_4279,N_3506,N_3759);
xor U4280 (N_4280,N_3596,N_3909);
nand U4281 (N_4281,N_3976,N_3902);
nand U4282 (N_4282,N_3992,N_3820);
and U4283 (N_4283,N_3964,N_3555);
and U4284 (N_4284,N_3915,N_3913);
or U4285 (N_4285,N_3635,N_3664);
and U4286 (N_4286,N_3997,N_3658);
nand U4287 (N_4287,N_3567,N_3603);
and U4288 (N_4288,N_3733,N_3883);
nor U4289 (N_4289,N_3697,N_3929);
or U4290 (N_4290,N_3702,N_3658);
and U4291 (N_4291,N_3506,N_3777);
and U4292 (N_4292,N_3847,N_3792);
and U4293 (N_4293,N_3753,N_3738);
xnor U4294 (N_4294,N_3992,N_3630);
and U4295 (N_4295,N_3945,N_3956);
nor U4296 (N_4296,N_3644,N_3555);
or U4297 (N_4297,N_3719,N_3956);
nand U4298 (N_4298,N_3909,N_3600);
nor U4299 (N_4299,N_3922,N_3969);
and U4300 (N_4300,N_3678,N_3806);
nor U4301 (N_4301,N_3670,N_3572);
or U4302 (N_4302,N_3873,N_3532);
nand U4303 (N_4303,N_3642,N_3760);
nor U4304 (N_4304,N_3588,N_3929);
nor U4305 (N_4305,N_3878,N_3789);
xnor U4306 (N_4306,N_3528,N_3637);
nor U4307 (N_4307,N_3908,N_3959);
nor U4308 (N_4308,N_3531,N_3722);
and U4309 (N_4309,N_3569,N_3785);
or U4310 (N_4310,N_3570,N_3562);
or U4311 (N_4311,N_3683,N_3694);
nand U4312 (N_4312,N_3725,N_3798);
nor U4313 (N_4313,N_3834,N_3836);
or U4314 (N_4314,N_3960,N_3984);
nand U4315 (N_4315,N_3874,N_3737);
xor U4316 (N_4316,N_3547,N_3801);
and U4317 (N_4317,N_3526,N_3993);
and U4318 (N_4318,N_3779,N_3752);
and U4319 (N_4319,N_3619,N_3798);
xor U4320 (N_4320,N_3782,N_3820);
and U4321 (N_4321,N_3617,N_3802);
xnor U4322 (N_4322,N_3573,N_3887);
or U4323 (N_4323,N_3938,N_3764);
or U4324 (N_4324,N_3810,N_3818);
nand U4325 (N_4325,N_3730,N_3971);
or U4326 (N_4326,N_3945,N_3680);
nand U4327 (N_4327,N_3889,N_3877);
or U4328 (N_4328,N_3648,N_3680);
xor U4329 (N_4329,N_3745,N_3709);
xnor U4330 (N_4330,N_3820,N_3967);
or U4331 (N_4331,N_3796,N_3722);
nand U4332 (N_4332,N_3513,N_3895);
nor U4333 (N_4333,N_3666,N_3812);
xnor U4334 (N_4334,N_3673,N_3738);
xor U4335 (N_4335,N_3746,N_3651);
nor U4336 (N_4336,N_3822,N_3785);
nand U4337 (N_4337,N_3668,N_3562);
nor U4338 (N_4338,N_3958,N_3681);
and U4339 (N_4339,N_3911,N_3946);
nand U4340 (N_4340,N_3587,N_3562);
xnor U4341 (N_4341,N_3609,N_3965);
or U4342 (N_4342,N_3718,N_3988);
xnor U4343 (N_4343,N_3934,N_3622);
xor U4344 (N_4344,N_3574,N_3513);
xnor U4345 (N_4345,N_3813,N_3796);
xor U4346 (N_4346,N_3842,N_3561);
and U4347 (N_4347,N_3971,N_3815);
xnor U4348 (N_4348,N_3789,N_3902);
and U4349 (N_4349,N_3969,N_3587);
nand U4350 (N_4350,N_3878,N_3621);
or U4351 (N_4351,N_3575,N_3662);
xor U4352 (N_4352,N_3582,N_3916);
nor U4353 (N_4353,N_3782,N_3783);
xnor U4354 (N_4354,N_3671,N_3528);
xor U4355 (N_4355,N_3889,N_3973);
xnor U4356 (N_4356,N_3947,N_3989);
and U4357 (N_4357,N_3614,N_3882);
or U4358 (N_4358,N_3729,N_3670);
or U4359 (N_4359,N_3716,N_3842);
and U4360 (N_4360,N_3844,N_3796);
xnor U4361 (N_4361,N_3835,N_3742);
nor U4362 (N_4362,N_3613,N_3582);
and U4363 (N_4363,N_3801,N_3797);
or U4364 (N_4364,N_3706,N_3773);
or U4365 (N_4365,N_3854,N_3806);
or U4366 (N_4366,N_3744,N_3807);
nand U4367 (N_4367,N_3572,N_3621);
nor U4368 (N_4368,N_3571,N_3725);
nand U4369 (N_4369,N_3887,N_3948);
and U4370 (N_4370,N_3936,N_3788);
and U4371 (N_4371,N_3902,N_3740);
and U4372 (N_4372,N_3535,N_3761);
nor U4373 (N_4373,N_3669,N_3926);
nand U4374 (N_4374,N_3809,N_3543);
nand U4375 (N_4375,N_3994,N_3687);
xor U4376 (N_4376,N_3888,N_3621);
nand U4377 (N_4377,N_3589,N_3893);
nor U4378 (N_4378,N_3517,N_3976);
nor U4379 (N_4379,N_3795,N_3533);
nand U4380 (N_4380,N_3699,N_3874);
nor U4381 (N_4381,N_3850,N_3822);
nand U4382 (N_4382,N_3842,N_3661);
nor U4383 (N_4383,N_3665,N_3945);
and U4384 (N_4384,N_3888,N_3716);
and U4385 (N_4385,N_3997,N_3857);
or U4386 (N_4386,N_3863,N_3959);
nand U4387 (N_4387,N_3501,N_3577);
nand U4388 (N_4388,N_3591,N_3635);
nor U4389 (N_4389,N_3772,N_3658);
nor U4390 (N_4390,N_3786,N_3957);
xor U4391 (N_4391,N_3735,N_3505);
and U4392 (N_4392,N_3722,N_3951);
or U4393 (N_4393,N_3588,N_3835);
nand U4394 (N_4394,N_3776,N_3773);
nor U4395 (N_4395,N_3959,N_3979);
nand U4396 (N_4396,N_3922,N_3828);
xor U4397 (N_4397,N_3575,N_3753);
nor U4398 (N_4398,N_3879,N_3771);
or U4399 (N_4399,N_3927,N_3520);
and U4400 (N_4400,N_3915,N_3856);
xnor U4401 (N_4401,N_3918,N_3990);
or U4402 (N_4402,N_3615,N_3943);
nor U4403 (N_4403,N_3508,N_3684);
nand U4404 (N_4404,N_3714,N_3934);
xor U4405 (N_4405,N_3744,N_3607);
nor U4406 (N_4406,N_3530,N_3648);
and U4407 (N_4407,N_3860,N_3642);
or U4408 (N_4408,N_3826,N_3670);
nand U4409 (N_4409,N_3926,N_3594);
xnor U4410 (N_4410,N_3932,N_3908);
nor U4411 (N_4411,N_3555,N_3929);
nand U4412 (N_4412,N_3995,N_3984);
or U4413 (N_4413,N_3961,N_3764);
xor U4414 (N_4414,N_3867,N_3703);
nor U4415 (N_4415,N_3664,N_3579);
xor U4416 (N_4416,N_3538,N_3550);
and U4417 (N_4417,N_3953,N_3890);
and U4418 (N_4418,N_3682,N_3620);
nand U4419 (N_4419,N_3783,N_3685);
nand U4420 (N_4420,N_3636,N_3873);
nor U4421 (N_4421,N_3870,N_3961);
and U4422 (N_4422,N_3515,N_3567);
nor U4423 (N_4423,N_3868,N_3798);
and U4424 (N_4424,N_3918,N_3769);
xnor U4425 (N_4425,N_3955,N_3845);
xor U4426 (N_4426,N_3813,N_3985);
nor U4427 (N_4427,N_3924,N_3815);
nand U4428 (N_4428,N_3753,N_3542);
or U4429 (N_4429,N_3746,N_3672);
and U4430 (N_4430,N_3793,N_3887);
nand U4431 (N_4431,N_3797,N_3844);
xor U4432 (N_4432,N_3758,N_3613);
and U4433 (N_4433,N_3912,N_3768);
nand U4434 (N_4434,N_3718,N_3559);
xnor U4435 (N_4435,N_3636,N_3518);
and U4436 (N_4436,N_3842,N_3933);
nand U4437 (N_4437,N_3701,N_3938);
xnor U4438 (N_4438,N_3661,N_3793);
nor U4439 (N_4439,N_3753,N_3993);
nor U4440 (N_4440,N_3661,N_3829);
or U4441 (N_4441,N_3816,N_3865);
or U4442 (N_4442,N_3793,N_3517);
or U4443 (N_4443,N_3507,N_3538);
and U4444 (N_4444,N_3658,N_3825);
nand U4445 (N_4445,N_3922,N_3758);
xnor U4446 (N_4446,N_3501,N_3527);
xnor U4447 (N_4447,N_3610,N_3896);
nor U4448 (N_4448,N_3589,N_3800);
nor U4449 (N_4449,N_3941,N_3986);
xnor U4450 (N_4450,N_3603,N_3706);
or U4451 (N_4451,N_3676,N_3545);
nor U4452 (N_4452,N_3647,N_3571);
nand U4453 (N_4453,N_3570,N_3505);
or U4454 (N_4454,N_3758,N_3948);
or U4455 (N_4455,N_3609,N_3703);
nor U4456 (N_4456,N_3707,N_3925);
nor U4457 (N_4457,N_3673,N_3955);
nand U4458 (N_4458,N_3559,N_3709);
or U4459 (N_4459,N_3644,N_3540);
or U4460 (N_4460,N_3670,N_3515);
nand U4461 (N_4461,N_3562,N_3574);
nor U4462 (N_4462,N_3755,N_3927);
nand U4463 (N_4463,N_3647,N_3990);
nor U4464 (N_4464,N_3836,N_3728);
nor U4465 (N_4465,N_3999,N_3747);
and U4466 (N_4466,N_3736,N_3906);
and U4467 (N_4467,N_3541,N_3700);
and U4468 (N_4468,N_3781,N_3753);
or U4469 (N_4469,N_3927,N_3834);
nand U4470 (N_4470,N_3947,N_3742);
nand U4471 (N_4471,N_3582,N_3787);
nor U4472 (N_4472,N_3909,N_3650);
nand U4473 (N_4473,N_3867,N_3700);
and U4474 (N_4474,N_3944,N_3910);
xnor U4475 (N_4475,N_3675,N_3981);
xor U4476 (N_4476,N_3901,N_3898);
and U4477 (N_4477,N_3670,N_3678);
and U4478 (N_4478,N_3968,N_3583);
nor U4479 (N_4479,N_3907,N_3613);
xnor U4480 (N_4480,N_3919,N_3993);
or U4481 (N_4481,N_3507,N_3589);
nor U4482 (N_4482,N_3608,N_3609);
or U4483 (N_4483,N_3947,N_3806);
nor U4484 (N_4484,N_3760,N_3974);
and U4485 (N_4485,N_3853,N_3775);
nor U4486 (N_4486,N_3757,N_3707);
and U4487 (N_4487,N_3832,N_3886);
or U4488 (N_4488,N_3882,N_3954);
nor U4489 (N_4489,N_3739,N_3514);
xnor U4490 (N_4490,N_3629,N_3920);
or U4491 (N_4491,N_3595,N_3848);
or U4492 (N_4492,N_3646,N_3703);
and U4493 (N_4493,N_3788,N_3894);
nor U4494 (N_4494,N_3636,N_3676);
xnor U4495 (N_4495,N_3848,N_3613);
and U4496 (N_4496,N_3646,N_3635);
or U4497 (N_4497,N_3668,N_3969);
nor U4498 (N_4498,N_3872,N_3858);
nor U4499 (N_4499,N_3644,N_3709);
nand U4500 (N_4500,N_4108,N_4081);
nand U4501 (N_4501,N_4302,N_4490);
nor U4502 (N_4502,N_4013,N_4179);
and U4503 (N_4503,N_4232,N_4330);
nand U4504 (N_4504,N_4198,N_4489);
and U4505 (N_4505,N_4225,N_4461);
and U4506 (N_4506,N_4216,N_4364);
nor U4507 (N_4507,N_4460,N_4438);
nor U4508 (N_4508,N_4261,N_4235);
and U4509 (N_4509,N_4095,N_4060);
nand U4510 (N_4510,N_4498,N_4337);
nand U4511 (N_4511,N_4488,N_4007);
nand U4512 (N_4512,N_4247,N_4286);
nor U4513 (N_4513,N_4105,N_4205);
or U4514 (N_4514,N_4413,N_4213);
nor U4515 (N_4515,N_4383,N_4174);
nand U4516 (N_4516,N_4113,N_4030);
and U4517 (N_4517,N_4285,N_4079);
nor U4518 (N_4518,N_4431,N_4069);
xor U4519 (N_4519,N_4208,N_4097);
and U4520 (N_4520,N_4355,N_4047);
xor U4521 (N_4521,N_4037,N_4196);
nand U4522 (N_4522,N_4085,N_4019);
xor U4523 (N_4523,N_4416,N_4146);
and U4524 (N_4524,N_4478,N_4022);
nand U4525 (N_4525,N_4031,N_4207);
nor U4526 (N_4526,N_4137,N_4011);
and U4527 (N_4527,N_4428,N_4058);
nand U4528 (N_4528,N_4424,N_4126);
and U4529 (N_4529,N_4064,N_4088);
nand U4530 (N_4530,N_4094,N_4118);
or U4531 (N_4531,N_4408,N_4270);
nand U4532 (N_4532,N_4300,N_4417);
or U4533 (N_4533,N_4138,N_4115);
and U4534 (N_4534,N_4362,N_4437);
or U4535 (N_4535,N_4410,N_4005);
or U4536 (N_4536,N_4200,N_4131);
or U4537 (N_4537,N_4043,N_4173);
xnor U4538 (N_4538,N_4432,N_4176);
xnor U4539 (N_4539,N_4405,N_4068);
nand U4540 (N_4540,N_4393,N_4376);
nand U4541 (N_4541,N_4091,N_4481);
nand U4542 (N_4542,N_4296,N_4497);
nor U4543 (N_4543,N_4499,N_4434);
or U4544 (N_4544,N_4483,N_4074);
xnor U4545 (N_4545,N_4239,N_4293);
and U4546 (N_4546,N_4443,N_4275);
xor U4547 (N_4547,N_4280,N_4243);
or U4548 (N_4548,N_4265,N_4283);
nor U4549 (N_4549,N_4002,N_4096);
nand U4550 (N_4550,N_4229,N_4429);
xnor U4551 (N_4551,N_4345,N_4394);
xor U4552 (N_4552,N_4082,N_4375);
nor U4553 (N_4553,N_4199,N_4034);
nor U4554 (N_4554,N_4366,N_4320);
nand U4555 (N_4555,N_4441,N_4141);
nor U4556 (N_4556,N_4258,N_4365);
nor U4557 (N_4557,N_4358,N_4197);
nor U4558 (N_4558,N_4324,N_4440);
or U4559 (N_4559,N_4476,N_4127);
nand U4560 (N_4560,N_4363,N_4316);
xor U4561 (N_4561,N_4192,N_4400);
or U4562 (N_4562,N_4103,N_4252);
or U4563 (N_4563,N_4214,N_4122);
or U4564 (N_4564,N_4102,N_4160);
nor U4565 (N_4565,N_4397,N_4426);
and U4566 (N_4566,N_4249,N_4189);
or U4567 (N_4567,N_4224,N_4299);
nor U4568 (N_4568,N_4396,N_4350);
and U4569 (N_4569,N_4399,N_4412);
xnor U4570 (N_4570,N_4238,N_4303);
nand U4571 (N_4571,N_4178,N_4301);
or U4572 (N_4572,N_4430,N_4486);
nand U4573 (N_4573,N_4382,N_4215);
or U4574 (N_4574,N_4304,N_4023);
and U4575 (N_4575,N_4052,N_4371);
and U4576 (N_4576,N_4143,N_4253);
and U4577 (N_4577,N_4260,N_4279);
nor U4578 (N_4578,N_4020,N_4256);
xnor U4579 (N_4579,N_4480,N_4357);
nand U4580 (N_4580,N_4310,N_4177);
nor U4581 (N_4581,N_4202,N_4346);
or U4582 (N_4582,N_4090,N_4361);
or U4583 (N_4583,N_4334,N_4028);
xnor U4584 (N_4584,N_4152,N_4435);
nand U4585 (N_4585,N_4464,N_4135);
and U4586 (N_4586,N_4193,N_4297);
nor U4587 (N_4587,N_4233,N_4185);
or U4588 (N_4588,N_4419,N_4191);
nand U4589 (N_4589,N_4356,N_4231);
nand U4590 (N_4590,N_4289,N_4351);
xor U4591 (N_4591,N_4084,N_4341);
xor U4592 (N_4592,N_4133,N_4264);
or U4593 (N_4593,N_4164,N_4445);
nand U4594 (N_4594,N_4159,N_4099);
nor U4595 (N_4595,N_4277,N_4487);
or U4596 (N_4596,N_4271,N_4388);
xor U4597 (N_4597,N_4495,N_4251);
xor U4598 (N_4598,N_4325,N_4244);
nand U4599 (N_4599,N_4479,N_4121);
nor U4600 (N_4600,N_4147,N_4041);
nor U4601 (N_4601,N_4015,N_4267);
nor U4602 (N_4602,N_4234,N_4162);
or U4603 (N_4603,N_4403,N_4306);
or U4604 (N_4604,N_4190,N_4378);
xor U4605 (N_4605,N_4001,N_4077);
nand U4606 (N_4606,N_4117,N_4292);
nand U4607 (N_4607,N_4312,N_4448);
nor U4608 (N_4608,N_4046,N_4009);
nor U4609 (N_4609,N_4457,N_4245);
and U4610 (N_4610,N_4427,N_4183);
xnor U4611 (N_4611,N_4053,N_4367);
and U4612 (N_4612,N_4067,N_4452);
and U4613 (N_4613,N_4421,N_4212);
nor U4614 (N_4614,N_4402,N_4153);
xnor U4615 (N_4615,N_4175,N_4093);
xor U4616 (N_4616,N_4398,N_4401);
and U4617 (N_4617,N_4107,N_4321);
and U4618 (N_4618,N_4033,N_4278);
xor U4619 (N_4619,N_4282,N_4418);
or U4620 (N_4620,N_4469,N_4161);
nor U4621 (N_4621,N_4230,N_4119);
or U4622 (N_4622,N_4142,N_4101);
nor U4623 (N_4623,N_4467,N_4057);
or U4624 (N_4624,N_4054,N_4468);
nor U4625 (N_4625,N_4112,N_4257);
xnor U4626 (N_4626,N_4343,N_4169);
or U4627 (N_4627,N_4317,N_4444);
or U4628 (N_4628,N_4227,N_4336);
and U4629 (N_4629,N_4311,N_4262);
and U4630 (N_4630,N_4106,N_4027);
xnor U4631 (N_4631,N_4433,N_4342);
and U4632 (N_4632,N_4063,N_4080);
or U4633 (N_4633,N_4319,N_4474);
or U4634 (N_4634,N_4423,N_4014);
or U4635 (N_4635,N_4032,N_4184);
nand U4636 (N_4636,N_4470,N_4222);
xor U4637 (N_4637,N_4129,N_4315);
nand U4638 (N_4638,N_4166,N_4255);
nor U4639 (N_4639,N_4092,N_4048);
xor U4640 (N_4640,N_4484,N_4287);
xor U4641 (N_4641,N_4349,N_4450);
or U4642 (N_4642,N_4026,N_4273);
xor U4643 (N_4643,N_4422,N_4295);
or U4644 (N_4644,N_4132,N_4110);
xor U4645 (N_4645,N_4347,N_4078);
nand U4646 (N_4646,N_4409,N_4328);
nand U4647 (N_4647,N_4195,N_4155);
nand U4648 (N_4648,N_4272,N_4274);
or U4649 (N_4649,N_4242,N_4259);
xnor U4650 (N_4650,N_4477,N_4309);
xor U4651 (N_4651,N_4045,N_4021);
xor U4652 (N_4652,N_4220,N_4368);
and U4653 (N_4653,N_4018,N_4136);
xor U4654 (N_4654,N_4145,N_4459);
nor U4655 (N_4655,N_4024,N_4050);
and U4656 (N_4656,N_4236,N_4056);
nand U4657 (N_4657,N_4223,N_4254);
or U4658 (N_4658,N_4010,N_4348);
nor U4659 (N_4659,N_4333,N_4327);
and U4660 (N_4660,N_4447,N_4065);
or U4661 (N_4661,N_4210,N_4128);
or U4662 (N_4662,N_4298,N_4455);
xnor U4663 (N_4663,N_4114,N_4016);
nor U4664 (N_4664,N_4111,N_4322);
or U4665 (N_4665,N_4269,N_4439);
nor U4666 (N_4666,N_4218,N_4458);
or U4667 (N_4667,N_4151,N_4389);
nor U4668 (N_4668,N_4241,N_4221);
or U4669 (N_4669,N_4237,N_4449);
xor U4670 (N_4670,N_4462,N_4339);
or U4671 (N_4671,N_4039,N_4062);
and U4672 (N_4672,N_4250,N_4149);
nor U4673 (N_4673,N_4124,N_4381);
xnor U4674 (N_4674,N_4130,N_4150);
nor U4675 (N_4675,N_4073,N_4456);
xnor U4676 (N_4676,N_4000,N_4465);
nor U4677 (N_4677,N_4171,N_4109);
and U4678 (N_4678,N_4219,N_4120);
xnor U4679 (N_4679,N_4370,N_4475);
nor U4680 (N_4680,N_4036,N_4288);
or U4681 (N_4681,N_4003,N_4305);
and U4682 (N_4682,N_4411,N_4385);
xor U4683 (N_4683,N_4029,N_4211);
xnor U4684 (N_4684,N_4331,N_4042);
and U4685 (N_4685,N_4466,N_4025);
nand U4686 (N_4686,N_4040,N_4471);
xor U4687 (N_4687,N_4201,N_4404);
nand U4688 (N_4688,N_4374,N_4387);
nand U4689 (N_4689,N_4463,N_4061);
and U4690 (N_4690,N_4104,N_4359);
nand U4691 (N_4691,N_4318,N_4436);
xor U4692 (N_4692,N_4246,N_4494);
and U4693 (N_4693,N_4167,N_4390);
and U4694 (N_4694,N_4072,N_4194);
and U4695 (N_4695,N_4116,N_4071);
or U4696 (N_4696,N_4144,N_4360);
nand U4697 (N_4697,N_4098,N_4075);
or U4698 (N_4698,N_4485,N_4181);
nand U4699 (N_4699,N_4323,N_4313);
nor U4700 (N_4700,N_4188,N_4373);
nor U4701 (N_4701,N_4496,N_4377);
nor U4702 (N_4702,N_4384,N_4157);
and U4703 (N_4703,N_4154,N_4386);
xor U4704 (N_4704,N_4380,N_4482);
xor U4705 (N_4705,N_4172,N_4035);
nand U4706 (N_4706,N_4148,N_4392);
xor U4707 (N_4707,N_4017,N_4406);
or U4708 (N_4708,N_4086,N_4228);
and U4709 (N_4709,N_4492,N_4281);
xor U4710 (N_4710,N_4168,N_4240);
and U4711 (N_4711,N_4263,N_4472);
nor U4712 (N_4712,N_4070,N_4170);
nand U4713 (N_4713,N_4055,N_4049);
or U4714 (N_4714,N_4206,N_4451);
nand U4715 (N_4715,N_4326,N_4180);
xnor U4716 (N_4716,N_4446,N_4407);
xor U4717 (N_4717,N_4187,N_4209);
and U4718 (N_4718,N_4051,N_4415);
nand U4719 (N_4719,N_4268,N_4493);
and U4720 (N_4720,N_4308,N_4248);
nor U4721 (N_4721,N_4352,N_4414);
nand U4722 (N_4722,N_4044,N_4083);
nand U4723 (N_4723,N_4266,N_4395);
nor U4724 (N_4724,N_4332,N_4038);
and U4725 (N_4725,N_4089,N_4291);
and U4726 (N_4726,N_4491,N_4217);
or U4727 (N_4727,N_4156,N_4134);
xnor U4728 (N_4728,N_4165,N_4123);
or U4729 (N_4729,N_4307,N_4425);
or U4730 (N_4730,N_4008,N_4454);
and U4731 (N_4731,N_4158,N_4182);
nor U4732 (N_4732,N_4329,N_4276);
or U4733 (N_4733,N_4353,N_4294);
xnor U4734 (N_4734,N_4006,N_4284);
or U4735 (N_4735,N_4453,N_4369);
xor U4736 (N_4736,N_4335,N_4163);
and U4737 (N_4737,N_4473,N_4354);
or U4738 (N_4738,N_4139,N_4076);
xor U4739 (N_4739,N_4420,N_4066);
and U4740 (N_4740,N_4100,N_4203);
xnor U4741 (N_4741,N_4391,N_4340);
nand U4742 (N_4742,N_4087,N_4442);
nor U4743 (N_4743,N_4004,N_4290);
nand U4744 (N_4744,N_4338,N_4012);
or U4745 (N_4745,N_4372,N_4125);
or U4746 (N_4746,N_4059,N_4140);
nor U4747 (N_4747,N_4186,N_4226);
nand U4748 (N_4748,N_4314,N_4204);
nand U4749 (N_4749,N_4379,N_4344);
nand U4750 (N_4750,N_4085,N_4284);
or U4751 (N_4751,N_4057,N_4377);
xnor U4752 (N_4752,N_4058,N_4293);
nor U4753 (N_4753,N_4400,N_4415);
xnor U4754 (N_4754,N_4499,N_4081);
and U4755 (N_4755,N_4151,N_4452);
or U4756 (N_4756,N_4249,N_4379);
or U4757 (N_4757,N_4401,N_4335);
nand U4758 (N_4758,N_4110,N_4170);
or U4759 (N_4759,N_4334,N_4391);
and U4760 (N_4760,N_4277,N_4281);
nand U4761 (N_4761,N_4138,N_4129);
nor U4762 (N_4762,N_4456,N_4375);
and U4763 (N_4763,N_4154,N_4176);
nor U4764 (N_4764,N_4278,N_4213);
and U4765 (N_4765,N_4374,N_4234);
nand U4766 (N_4766,N_4243,N_4189);
or U4767 (N_4767,N_4445,N_4409);
nand U4768 (N_4768,N_4461,N_4490);
or U4769 (N_4769,N_4303,N_4015);
nor U4770 (N_4770,N_4088,N_4058);
and U4771 (N_4771,N_4346,N_4294);
xor U4772 (N_4772,N_4364,N_4420);
nor U4773 (N_4773,N_4474,N_4011);
nand U4774 (N_4774,N_4047,N_4368);
or U4775 (N_4775,N_4050,N_4068);
xor U4776 (N_4776,N_4316,N_4300);
nor U4777 (N_4777,N_4260,N_4061);
or U4778 (N_4778,N_4380,N_4468);
nand U4779 (N_4779,N_4460,N_4256);
nand U4780 (N_4780,N_4386,N_4091);
nor U4781 (N_4781,N_4157,N_4088);
or U4782 (N_4782,N_4006,N_4019);
nor U4783 (N_4783,N_4289,N_4184);
and U4784 (N_4784,N_4027,N_4428);
xnor U4785 (N_4785,N_4401,N_4071);
xnor U4786 (N_4786,N_4123,N_4402);
xor U4787 (N_4787,N_4347,N_4007);
xor U4788 (N_4788,N_4259,N_4225);
xnor U4789 (N_4789,N_4470,N_4447);
xnor U4790 (N_4790,N_4269,N_4422);
nor U4791 (N_4791,N_4361,N_4196);
and U4792 (N_4792,N_4155,N_4391);
and U4793 (N_4793,N_4042,N_4271);
nor U4794 (N_4794,N_4473,N_4453);
or U4795 (N_4795,N_4328,N_4119);
nand U4796 (N_4796,N_4184,N_4118);
or U4797 (N_4797,N_4097,N_4015);
xor U4798 (N_4798,N_4078,N_4425);
and U4799 (N_4799,N_4227,N_4394);
nand U4800 (N_4800,N_4064,N_4149);
nand U4801 (N_4801,N_4229,N_4038);
nand U4802 (N_4802,N_4234,N_4186);
or U4803 (N_4803,N_4479,N_4246);
nor U4804 (N_4804,N_4380,N_4083);
or U4805 (N_4805,N_4306,N_4013);
xnor U4806 (N_4806,N_4295,N_4019);
or U4807 (N_4807,N_4219,N_4195);
and U4808 (N_4808,N_4349,N_4306);
and U4809 (N_4809,N_4264,N_4386);
or U4810 (N_4810,N_4437,N_4374);
nand U4811 (N_4811,N_4371,N_4349);
nand U4812 (N_4812,N_4368,N_4064);
nand U4813 (N_4813,N_4356,N_4191);
xor U4814 (N_4814,N_4137,N_4230);
nor U4815 (N_4815,N_4398,N_4305);
xnor U4816 (N_4816,N_4055,N_4499);
or U4817 (N_4817,N_4374,N_4109);
xor U4818 (N_4818,N_4112,N_4118);
xnor U4819 (N_4819,N_4271,N_4380);
nand U4820 (N_4820,N_4074,N_4449);
and U4821 (N_4821,N_4182,N_4029);
nand U4822 (N_4822,N_4128,N_4197);
and U4823 (N_4823,N_4446,N_4495);
xor U4824 (N_4824,N_4332,N_4122);
xor U4825 (N_4825,N_4193,N_4027);
and U4826 (N_4826,N_4222,N_4199);
nand U4827 (N_4827,N_4213,N_4406);
and U4828 (N_4828,N_4356,N_4319);
or U4829 (N_4829,N_4217,N_4131);
xor U4830 (N_4830,N_4115,N_4175);
xnor U4831 (N_4831,N_4450,N_4130);
nor U4832 (N_4832,N_4233,N_4326);
nor U4833 (N_4833,N_4469,N_4453);
or U4834 (N_4834,N_4286,N_4149);
nand U4835 (N_4835,N_4081,N_4264);
xnor U4836 (N_4836,N_4287,N_4470);
and U4837 (N_4837,N_4057,N_4073);
or U4838 (N_4838,N_4411,N_4302);
and U4839 (N_4839,N_4076,N_4407);
xor U4840 (N_4840,N_4157,N_4232);
or U4841 (N_4841,N_4313,N_4106);
or U4842 (N_4842,N_4203,N_4175);
nand U4843 (N_4843,N_4311,N_4463);
or U4844 (N_4844,N_4476,N_4364);
nand U4845 (N_4845,N_4189,N_4410);
nor U4846 (N_4846,N_4110,N_4159);
or U4847 (N_4847,N_4121,N_4134);
or U4848 (N_4848,N_4240,N_4103);
nor U4849 (N_4849,N_4125,N_4149);
or U4850 (N_4850,N_4312,N_4218);
xnor U4851 (N_4851,N_4029,N_4400);
or U4852 (N_4852,N_4098,N_4466);
nor U4853 (N_4853,N_4234,N_4214);
xnor U4854 (N_4854,N_4050,N_4265);
and U4855 (N_4855,N_4041,N_4466);
xor U4856 (N_4856,N_4487,N_4240);
nor U4857 (N_4857,N_4249,N_4460);
or U4858 (N_4858,N_4271,N_4167);
xnor U4859 (N_4859,N_4392,N_4364);
nor U4860 (N_4860,N_4022,N_4446);
and U4861 (N_4861,N_4260,N_4418);
xor U4862 (N_4862,N_4299,N_4334);
nor U4863 (N_4863,N_4266,N_4050);
nor U4864 (N_4864,N_4049,N_4310);
nand U4865 (N_4865,N_4482,N_4105);
xnor U4866 (N_4866,N_4056,N_4065);
nand U4867 (N_4867,N_4231,N_4209);
nand U4868 (N_4868,N_4494,N_4191);
and U4869 (N_4869,N_4128,N_4227);
nand U4870 (N_4870,N_4375,N_4353);
or U4871 (N_4871,N_4221,N_4402);
or U4872 (N_4872,N_4329,N_4416);
xnor U4873 (N_4873,N_4359,N_4453);
xor U4874 (N_4874,N_4459,N_4110);
xor U4875 (N_4875,N_4290,N_4074);
or U4876 (N_4876,N_4124,N_4463);
nor U4877 (N_4877,N_4065,N_4336);
or U4878 (N_4878,N_4236,N_4174);
nor U4879 (N_4879,N_4191,N_4440);
nor U4880 (N_4880,N_4087,N_4227);
nor U4881 (N_4881,N_4386,N_4380);
or U4882 (N_4882,N_4469,N_4230);
nand U4883 (N_4883,N_4149,N_4264);
nand U4884 (N_4884,N_4055,N_4011);
and U4885 (N_4885,N_4237,N_4430);
and U4886 (N_4886,N_4434,N_4245);
nand U4887 (N_4887,N_4414,N_4072);
nand U4888 (N_4888,N_4116,N_4121);
nor U4889 (N_4889,N_4217,N_4213);
nand U4890 (N_4890,N_4100,N_4306);
or U4891 (N_4891,N_4243,N_4402);
nand U4892 (N_4892,N_4394,N_4082);
or U4893 (N_4893,N_4476,N_4133);
nand U4894 (N_4894,N_4164,N_4385);
nor U4895 (N_4895,N_4457,N_4376);
xor U4896 (N_4896,N_4209,N_4470);
nand U4897 (N_4897,N_4157,N_4255);
nor U4898 (N_4898,N_4454,N_4105);
and U4899 (N_4899,N_4402,N_4356);
xor U4900 (N_4900,N_4174,N_4283);
or U4901 (N_4901,N_4177,N_4012);
or U4902 (N_4902,N_4121,N_4448);
or U4903 (N_4903,N_4405,N_4193);
nor U4904 (N_4904,N_4363,N_4042);
or U4905 (N_4905,N_4495,N_4059);
and U4906 (N_4906,N_4292,N_4375);
xnor U4907 (N_4907,N_4033,N_4047);
and U4908 (N_4908,N_4495,N_4126);
nor U4909 (N_4909,N_4005,N_4456);
and U4910 (N_4910,N_4195,N_4442);
nor U4911 (N_4911,N_4131,N_4462);
and U4912 (N_4912,N_4370,N_4429);
nand U4913 (N_4913,N_4367,N_4113);
xnor U4914 (N_4914,N_4087,N_4237);
xor U4915 (N_4915,N_4312,N_4066);
and U4916 (N_4916,N_4323,N_4258);
nand U4917 (N_4917,N_4337,N_4014);
nand U4918 (N_4918,N_4200,N_4079);
nand U4919 (N_4919,N_4492,N_4201);
or U4920 (N_4920,N_4347,N_4140);
xor U4921 (N_4921,N_4046,N_4375);
and U4922 (N_4922,N_4216,N_4078);
nand U4923 (N_4923,N_4465,N_4374);
or U4924 (N_4924,N_4311,N_4219);
and U4925 (N_4925,N_4337,N_4490);
nor U4926 (N_4926,N_4457,N_4178);
and U4927 (N_4927,N_4360,N_4283);
or U4928 (N_4928,N_4075,N_4343);
nand U4929 (N_4929,N_4179,N_4286);
or U4930 (N_4930,N_4288,N_4081);
xnor U4931 (N_4931,N_4169,N_4295);
and U4932 (N_4932,N_4293,N_4254);
nor U4933 (N_4933,N_4021,N_4203);
xor U4934 (N_4934,N_4451,N_4462);
nor U4935 (N_4935,N_4125,N_4246);
nand U4936 (N_4936,N_4027,N_4011);
and U4937 (N_4937,N_4008,N_4441);
nor U4938 (N_4938,N_4193,N_4285);
or U4939 (N_4939,N_4309,N_4342);
nand U4940 (N_4940,N_4418,N_4087);
nor U4941 (N_4941,N_4481,N_4378);
xnor U4942 (N_4942,N_4286,N_4352);
xnor U4943 (N_4943,N_4084,N_4398);
or U4944 (N_4944,N_4455,N_4012);
or U4945 (N_4945,N_4496,N_4024);
or U4946 (N_4946,N_4450,N_4470);
xnor U4947 (N_4947,N_4299,N_4292);
and U4948 (N_4948,N_4120,N_4254);
nor U4949 (N_4949,N_4366,N_4400);
and U4950 (N_4950,N_4317,N_4341);
nor U4951 (N_4951,N_4355,N_4342);
and U4952 (N_4952,N_4109,N_4371);
xor U4953 (N_4953,N_4024,N_4272);
nor U4954 (N_4954,N_4189,N_4074);
or U4955 (N_4955,N_4485,N_4093);
nor U4956 (N_4956,N_4112,N_4233);
nor U4957 (N_4957,N_4178,N_4413);
nor U4958 (N_4958,N_4434,N_4382);
nand U4959 (N_4959,N_4407,N_4036);
nor U4960 (N_4960,N_4405,N_4243);
or U4961 (N_4961,N_4200,N_4165);
xor U4962 (N_4962,N_4391,N_4307);
xor U4963 (N_4963,N_4102,N_4238);
nor U4964 (N_4964,N_4306,N_4266);
xnor U4965 (N_4965,N_4172,N_4085);
nand U4966 (N_4966,N_4244,N_4136);
nor U4967 (N_4967,N_4040,N_4461);
nor U4968 (N_4968,N_4344,N_4223);
nand U4969 (N_4969,N_4001,N_4410);
xor U4970 (N_4970,N_4265,N_4070);
nor U4971 (N_4971,N_4069,N_4024);
xnor U4972 (N_4972,N_4224,N_4033);
nand U4973 (N_4973,N_4080,N_4400);
and U4974 (N_4974,N_4281,N_4280);
xnor U4975 (N_4975,N_4124,N_4087);
xnor U4976 (N_4976,N_4135,N_4432);
xnor U4977 (N_4977,N_4321,N_4046);
xnor U4978 (N_4978,N_4431,N_4422);
xor U4979 (N_4979,N_4430,N_4474);
nor U4980 (N_4980,N_4191,N_4046);
nand U4981 (N_4981,N_4415,N_4049);
nor U4982 (N_4982,N_4419,N_4178);
nor U4983 (N_4983,N_4042,N_4255);
xnor U4984 (N_4984,N_4011,N_4300);
xnor U4985 (N_4985,N_4072,N_4339);
nand U4986 (N_4986,N_4403,N_4383);
nor U4987 (N_4987,N_4097,N_4480);
nor U4988 (N_4988,N_4463,N_4138);
xnor U4989 (N_4989,N_4447,N_4011);
or U4990 (N_4990,N_4023,N_4250);
or U4991 (N_4991,N_4321,N_4058);
nand U4992 (N_4992,N_4026,N_4048);
nor U4993 (N_4993,N_4418,N_4284);
or U4994 (N_4994,N_4194,N_4394);
and U4995 (N_4995,N_4484,N_4191);
and U4996 (N_4996,N_4142,N_4377);
nor U4997 (N_4997,N_4086,N_4461);
nand U4998 (N_4998,N_4403,N_4099);
nand U4999 (N_4999,N_4070,N_4420);
and U5000 (N_5000,N_4685,N_4523);
or U5001 (N_5001,N_4540,N_4802);
and U5002 (N_5002,N_4681,N_4987);
nor U5003 (N_5003,N_4677,N_4580);
xor U5004 (N_5004,N_4882,N_4786);
nand U5005 (N_5005,N_4625,N_4683);
nor U5006 (N_5006,N_4745,N_4964);
nor U5007 (N_5007,N_4817,N_4945);
xor U5008 (N_5008,N_4597,N_4521);
and U5009 (N_5009,N_4844,N_4503);
or U5010 (N_5010,N_4759,N_4660);
or U5011 (N_5011,N_4637,N_4848);
xor U5012 (N_5012,N_4651,N_4618);
nor U5013 (N_5013,N_4881,N_4722);
or U5014 (N_5014,N_4859,N_4500);
nand U5015 (N_5015,N_4914,N_4729);
or U5016 (N_5016,N_4734,N_4510);
nand U5017 (N_5017,N_4645,N_4505);
and U5018 (N_5018,N_4575,N_4943);
and U5019 (N_5019,N_4546,N_4872);
and U5020 (N_5020,N_4902,N_4849);
xor U5021 (N_5021,N_4838,N_4811);
or U5022 (N_5022,N_4871,N_4696);
nand U5023 (N_5023,N_4702,N_4958);
nor U5024 (N_5024,N_4531,N_4530);
nor U5025 (N_5025,N_4732,N_4843);
nor U5026 (N_5026,N_4669,N_4918);
or U5027 (N_5027,N_4993,N_4930);
and U5028 (N_5028,N_4558,N_4852);
nor U5029 (N_5029,N_4887,N_4717);
and U5030 (N_5030,N_4690,N_4524);
xor U5031 (N_5031,N_4527,N_4782);
or U5032 (N_5032,N_4954,N_4536);
nand U5033 (N_5033,N_4623,N_4674);
nand U5034 (N_5034,N_4513,N_4680);
and U5035 (N_5035,N_4877,N_4707);
xnor U5036 (N_5036,N_4790,N_4659);
and U5037 (N_5037,N_4648,N_4661);
and U5038 (N_5038,N_4746,N_4551);
or U5039 (N_5039,N_4856,N_4547);
or U5040 (N_5040,N_4762,N_4989);
nand U5041 (N_5041,N_4619,N_4827);
nor U5042 (N_5042,N_4553,N_4678);
xnor U5043 (N_5043,N_4665,N_4839);
nor U5044 (N_5044,N_4658,N_4529);
xor U5045 (N_5045,N_4628,N_4990);
and U5046 (N_5046,N_4956,N_4721);
nand U5047 (N_5047,N_4919,N_4915);
xnor U5048 (N_5048,N_4591,N_4911);
and U5049 (N_5049,N_4953,N_4772);
or U5050 (N_5050,N_4894,N_4761);
xnor U5051 (N_5051,N_4544,N_4641);
xor U5052 (N_5052,N_4832,N_4886);
xor U5053 (N_5053,N_4944,N_4765);
nand U5054 (N_5054,N_4905,N_4506);
nor U5055 (N_5055,N_4507,N_4569);
and U5056 (N_5056,N_4635,N_4560);
xor U5057 (N_5057,N_4955,N_4692);
nor U5058 (N_5058,N_4596,N_4592);
and U5059 (N_5059,N_4809,N_4846);
xor U5060 (N_5060,N_4785,N_4508);
nor U5061 (N_5061,N_4663,N_4925);
and U5062 (N_5062,N_4627,N_4691);
nand U5063 (N_5063,N_4920,N_4934);
xnor U5064 (N_5064,N_4720,N_4939);
and U5065 (N_5065,N_4907,N_4766);
nand U5066 (N_5066,N_4948,N_4899);
and U5067 (N_5067,N_4537,N_4741);
nor U5068 (N_5068,N_4601,N_4781);
nor U5069 (N_5069,N_4855,N_4686);
or U5070 (N_5070,N_4795,N_4897);
or U5071 (N_5071,N_4815,N_4788);
and U5072 (N_5072,N_4584,N_4821);
nand U5073 (N_5073,N_4857,N_4824);
and U5074 (N_5074,N_4794,N_4805);
xnor U5075 (N_5075,N_4965,N_4552);
nand U5076 (N_5076,N_4727,N_4836);
or U5077 (N_5077,N_4937,N_4676);
xor U5078 (N_5078,N_4576,N_4869);
nor U5079 (N_5079,N_4906,N_4622);
nand U5080 (N_5080,N_4556,N_4992);
nor U5081 (N_5081,N_4779,N_4978);
xor U5082 (N_5082,N_4554,N_4797);
nand U5083 (N_5083,N_4563,N_4543);
nor U5084 (N_5084,N_4688,N_4742);
nand U5085 (N_5085,N_4895,N_4968);
and U5086 (N_5086,N_4800,N_4985);
or U5087 (N_5087,N_4578,N_4929);
xnor U5088 (N_5088,N_4583,N_4861);
and U5089 (N_5089,N_4644,N_4594);
nand U5090 (N_5090,N_4555,N_4670);
and U5091 (N_5091,N_4582,N_4853);
nand U5092 (N_5092,N_4643,N_4892);
nand U5093 (N_5093,N_4921,N_4932);
xor U5094 (N_5094,N_4514,N_4726);
or U5095 (N_5095,N_4896,N_4997);
nand U5096 (N_5096,N_4988,N_4977);
nand U5097 (N_5097,N_4776,N_4614);
or U5098 (N_5098,N_4890,N_4962);
xor U5099 (N_5099,N_4737,N_4705);
xor U5100 (N_5100,N_4784,N_4878);
or U5101 (N_5101,N_4769,N_4512);
nor U5102 (N_5102,N_4708,N_4980);
nand U5103 (N_5103,N_4862,N_4571);
or U5104 (N_5104,N_4868,N_4501);
and U5105 (N_5105,N_4866,N_4655);
nor U5106 (N_5106,N_4947,N_4996);
nand U5107 (N_5107,N_4664,N_4972);
and U5108 (N_5108,N_4751,N_4840);
or U5109 (N_5109,N_4940,N_4983);
xor U5110 (N_5110,N_4652,N_4998);
nand U5111 (N_5111,N_4904,N_4753);
xor U5112 (N_5112,N_4653,N_4697);
nand U5113 (N_5113,N_4917,N_4668);
xnor U5114 (N_5114,N_4783,N_4796);
nor U5115 (N_5115,N_4662,N_4960);
and U5116 (N_5116,N_4710,N_4842);
or U5117 (N_5117,N_4608,N_4851);
nor U5118 (N_5118,N_4957,N_4778);
nor U5119 (N_5119,N_4740,N_4654);
or U5120 (N_5120,N_4775,N_4963);
and U5121 (N_5121,N_4565,N_4928);
or U5122 (N_5122,N_4585,N_4548);
nand U5123 (N_5123,N_4950,N_4870);
and U5124 (N_5124,N_4981,N_4528);
and U5125 (N_5125,N_4716,N_4936);
xnor U5126 (N_5126,N_4994,N_4703);
or U5127 (N_5127,N_4874,N_4718);
and U5128 (N_5128,N_4952,N_4864);
or U5129 (N_5129,N_4519,N_4946);
xnor U5130 (N_5130,N_4709,N_4656);
nand U5131 (N_5131,N_4819,N_4533);
nand U5132 (N_5132,N_4646,N_4908);
nor U5133 (N_5133,N_4793,N_4901);
xor U5134 (N_5134,N_4822,N_4995);
xor U5135 (N_5135,N_4700,N_4538);
nand U5136 (N_5136,N_4876,N_4679);
xnor U5137 (N_5137,N_4941,N_4572);
nand U5138 (N_5138,N_4704,N_4739);
nand U5139 (N_5139,N_4682,N_4912);
nor U5140 (N_5140,N_4756,N_4639);
and U5141 (N_5141,N_4748,N_4595);
and U5142 (N_5142,N_4550,N_4603);
xnor U5143 (N_5143,N_4823,N_4975);
or U5144 (N_5144,N_4750,N_4615);
and U5145 (N_5145,N_4693,N_4673);
nor U5146 (N_5146,N_4933,N_4638);
and U5147 (N_5147,N_4774,N_4699);
xnor U5148 (N_5148,N_4816,N_4879);
xor U5149 (N_5149,N_4589,N_4806);
and U5150 (N_5150,N_4828,N_4631);
nand U5151 (N_5151,N_4675,N_4787);
nand U5152 (N_5152,N_4731,N_4599);
and U5153 (N_5153,N_4612,N_4620);
xor U5154 (N_5154,N_4557,N_4789);
nor U5155 (N_5155,N_4684,N_4758);
or U5156 (N_5156,N_4586,N_4567);
xor U5157 (N_5157,N_4974,N_4516);
nand U5158 (N_5158,N_4517,N_4967);
and U5159 (N_5159,N_4632,N_4723);
xnor U5160 (N_5160,N_4671,N_4949);
or U5161 (N_5161,N_4649,N_4860);
xor U5162 (N_5162,N_4728,N_4780);
nand U5163 (N_5163,N_4970,N_4971);
nand U5164 (N_5164,N_4520,N_4698);
nor U5165 (N_5165,N_4573,N_4830);
nor U5166 (N_5166,N_4885,N_4574);
or U5167 (N_5167,N_4518,N_4961);
nor U5168 (N_5168,N_4873,N_4744);
and U5169 (N_5169,N_4719,N_4770);
and U5170 (N_5170,N_4509,N_4714);
xnor U5171 (N_5171,N_4672,N_4791);
or U5172 (N_5172,N_4916,N_4969);
xor U5173 (N_5173,N_4511,N_4733);
or U5174 (N_5174,N_4755,N_4642);
xnor U5175 (N_5175,N_4834,N_4807);
or U5176 (N_5176,N_4711,N_4942);
or U5177 (N_5177,N_4845,N_4559);
and U5178 (N_5178,N_4837,N_4566);
nor U5179 (N_5179,N_4535,N_4754);
xnor U5180 (N_5180,N_4991,N_4689);
or U5181 (N_5181,N_4883,N_4577);
nand U5182 (N_5182,N_4854,N_4522);
or U5183 (N_5183,N_4799,N_4606);
or U5184 (N_5184,N_4621,N_4813);
nand U5185 (N_5185,N_4598,N_4561);
or U5186 (N_5186,N_4609,N_4630);
nor U5187 (N_5187,N_4835,N_4898);
nand U5188 (N_5188,N_4926,N_4979);
nor U5189 (N_5189,N_4951,N_4626);
nor U5190 (N_5190,N_4624,N_4613);
nor U5191 (N_5191,N_4777,N_4743);
nor U5192 (N_5192,N_4579,N_4590);
or U5193 (N_5193,N_4923,N_4810);
and U5194 (N_5194,N_4984,N_4829);
nor U5195 (N_5195,N_4549,N_4867);
or U5196 (N_5196,N_4713,N_4850);
and U5197 (N_5197,N_4910,N_4747);
nor U5198 (N_5198,N_4541,N_4938);
or U5199 (N_5199,N_4833,N_4636);
nand U5200 (N_5200,N_4735,N_4650);
or U5201 (N_5201,N_4924,N_4935);
and U5202 (N_5202,N_4738,N_4736);
or U5203 (N_5203,N_4647,N_4752);
nor U5204 (N_5204,N_4602,N_4767);
and U5205 (N_5205,N_4768,N_4927);
xnor U5206 (N_5206,N_4863,N_4808);
nor U5207 (N_5207,N_4875,N_4760);
nand U5208 (N_5208,N_4986,N_4525);
xnor U5209 (N_5209,N_4633,N_4812);
nor U5210 (N_5210,N_4730,N_4889);
nand U5211 (N_5211,N_4982,N_4600);
xnor U5212 (N_5212,N_4634,N_4803);
and U5213 (N_5213,N_4611,N_4706);
and U5214 (N_5214,N_4818,N_4909);
xnor U5215 (N_5215,N_4605,N_4564);
nor U5216 (N_5216,N_4562,N_4900);
xor U5217 (N_5217,N_4891,N_4826);
nand U5218 (N_5218,N_4712,N_4763);
xor U5219 (N_5219,N_4804,N_4913);
nor U5220 (N_5220,N_4667,N_4771);
nor U5221 (N_5221,N_4880,N_4757);
and U5222 (N_5222,N_4847,N_4568);
nor U5223 (N_5223,N_4903,N_4931);
nand U5224 (N_5224,N_4884,N_4966);
nand U5225 (N_5225,N_4616,N_4715);
nor U5226 (N_5226,N_4545,N_4841);
and U5227 (N_5227,N_4526,N_4687);
and U5228 (N_5228,N_4504,N_4502);
nand U5229 (N_5229,N_4640,N_4515);
nand U5230 (N_5230,N_4725,N_4666);
or U5231 (N_5231,N_4724,N_4749);
or U5232 (N_5232,N_4922,N_4593);
nor U5233 (N_5233,N_4657,N_4581);
or U5234 (N_5234,N_4865,N_4542);
and U5235 (N_5235,N_4695,N_4825);
or U5236 (N_5236,N_4893,N_4999);
and U5237 (N_5237,N_4801,N_4858);
xnor U5238 (N_5238,N_4604,N_4973);
or U5239 (N_5239,N_4798,N_4792);
xnor U5240 (N_5240,N_4831,N_4814);
nand U5241 (N_5241,N_4764,N_4570);
xnor U5242 (N_5242,N_4959,N_4694);
nand U5243 (N_5243,N_4701,N_4610);
nor U5244 (N_5244,N_4629,N_4888);
xnor U5245 (N_5245,N_4820,N_4588);
nor U5246 (N_5246,N_4539,N_4617);
xor U5247 (N_5247,N_4534,N_4532);
nor U5248 (N_5248,N_4607,N_4773);
xnor U5249 (N_5249,N_4976,N_4587);
and U5250 (N_5250,N_4946,N_4875);
or U5251 (N_5251,N_4567,N_4509);
nand U5252 (N_5252,N_4741,N_4573);
and U5253 (N_5253,N_4959,N_4508);
xor U5254 (N_5254,N_4543,N_4950);
and U5255 (N_5255,N_4912,N_4600);
xor U5256 (N_5256,N_4858,N_4585);
and U5257 (N_5257,N_4742,N_4556);
nor U5258 (N_5258,N_4811,N_4948);
xor U5259 (N_5259,N_4794,N_4834);
and U5260 (N_5260,N_4904,N_4744);
nand U5261 (N_5261,N_4798,N_4720);
nand U5262 (N_5262,N_4893,N_4798);
nand U5263 (N_5263,N_4906,N_4594);
xnor U5264 (N_5264,N_4567,N_4639);
nand U5265 (N_5265,N_4537,N_4513);
nor U5266 (N_5266,N_4765,N_4848);
or U5267 (N_5267,N_4979,N_4964);
and U5268 (N_5268,N_4873,N_4651);
nor U5269 (N_5269,N_4790,N_4847);
or U5270 (N_5270,N_4958,N_4980);
xor U5271 (N_5271,N_4555,N_4704);
or U5272 (N_5272,N_4846,N_4756);
and U5273 (N_5273,N_4533,N_4530);
nand U5274 (N_5274,N_4983,N_4719);
or U5275 (N_5275,N_4708,N_4919);
and U5276 (N_5276,N_4772,N_4985);
or U5277 (N_5277,N_4501,N_4819);
nor U5278 (N_5278,N_4993,N_4885);
nor U5279 (N_5279,N_4770,N_4812);
xnor U5280 (N_5280,N_4874,N_4553);
nand U5281 (N_5281,N_4764,N_4726);
xor U5282 (N_5282,N_4619,N_4925);
or U5283 (N_5283,N_4865,N_4710);
or U5284 (N_5284,N_4646,N_4753);
xor U5285 (N_5285,N_4796,N_4622);
xnor U5286 (N_5286,N_4717,N_4697);
xnor U5287 (N_5287,N_4734,N_4978);
and U5288 (N_5288,N_4661,N_4564);
nand U5289 (N_5289,N_4711,N_4753);
nand U5290 (N_5290,N_4656,N_4845);
or U5291 (N_5291,N_4505,N_4633);
xnor U5292 (N_5292,N_4580,N_4500);
nor U5293 (N_5293,N_4765,N_4760);
xor U5294 (N_5294,N_4816,N_4844);
nand U5295 (N_5295,N_4695,N_4711);
or U5296 (N_5296,N_4567,N_4797);
nand U5297 (N_5297,N_4624,N_4645);
nor U5298 (N_5298,N_4866,N_4989);
and U5299 (N_5299,N_4860,N_4747);
nand U5300 (N_5300,N_4736,N_4776);
or U5301 (N_5301,N_4590,N_4843);
nand U5302 (N_5302,N_4909,N_4838);
nand U5303 (N_5303,N_4915,N_4967);
and U5304 (N_5304,N_4957,N_4729);
or U5305 (N_5305,N_4539,N_4606);
and U5306 (N_5306,N_4573,N_4686);
xor U5307 (N_5307,N_4981,N_4944);
nor U5308 (N_5308,N_4907,N_4950);
nand U5309 (N_5309,N_4736,N_4667);
or U5310 (N_5310,N_4746,N_4868);
or U5311 (N_5311,N_4965,N_4885);
or U5312 (N_5312,N_4942,N_4521);
or U5313 (N_5313,N_4786,N_4778);
xnor U5314 (N_5314,N_4983,N_4753);
or U5315 (N_5315,N_4929,N_4567);
or U5316 (N_5316,N_4825,N_4676);
nand U5317 (N_5317,N_4792,N_4854);
and U5318 (N_5318,N_4956,N_4533);
or U5319 (N_5319,N_4619,N_4741);
or U5320 (N_5320,N_4594,N_4987);
nand U5321 (N_5321,N_4951,N_4912);
xnor U5322 (N_5322,N_4909,N_4597);
xnor U5323 (N_5323,N_4523,N_4969);
nand U5324 (N_5324,N_4541,N_4665);
and U5325 (N_5325,N_4642,N_4563);
nand U5326 (N_5326,N_4773,N_4867);
xnor U5327 (N_5327,N_4654,N_4584);
nor U5328 (N_5328,N_4919,N_4501);
nor U5329 (N_5329,N_4929,N_4855);
nor U5330 (N_5330,N_4520,N_4784);
and U5331 (N_5331,N_4617,N_4560);
xor U5332 (N_5332,N_4632,N_4824);
nand U5333 (N_5333,N_4605,N_4872);
xor U5334 (N_5334,N_4871,N_4523);
nor U5335 (N_5335,N_4577,N_4752);
nand U5336 (N_5336,N_4728,N_4882);
nand U5337 (N_5337,N_4851,N_4780);
or U5338 (N_5338,N_4858,N_4909);
nand U5339 (N_5339,N_4758,N_4734);
and U5340 (N_5340,N_4933,N_4968);
or U5341 (N_5341,N_4931,N_4507);
or U5342 (N_5342,N_4865,N_4789);
nand U5343 (N_5343,N_4869,N_4735);
or U5344 (N_5344,N_4713,N_4782);
and U5345 (N_5345,N_4679,N_4574);
nor U5346 (N_5346,N_4547,N_4792);
nand U5347 (N_5347,N_4502,N_4511);
xnor U5348 (N_5348,N_4826,N_4525);
or U5349 (N_5349,N_4609,N_4524);
and U5350 (N_5350,N_4862,N_4902);
xnor U5351 (N_5351,N_4654,N_4559);
xnor U5352 (N_5352,N_4649,N_4710);
xor U5353 (N_5353,N_4593,N_4508);
nand U5354 (N_5354,N_4980,N_4766);
xor U5355 (N_5355,N_4526,N_4714);
or U5356 (N_5356,N_4724,N_4551);
or U5357 (N_5357,N_4873,N_4925);
xor U5358 (N_5358,N_4684,N_4960);
nor U5359 (N_5359,N_4726,N_4684);
nand U5360 (N_5360,N_4597,N_4971);
and U5361 (N_5361,N_4858,N_4505);
nor U5362 (N_5362,N_4642,N_4886);
nor U5363 (N_5363,N_4685,N_4606);
and U5364 (N_5364,N_4853,N_4940);
and U5365 (N_5365,N_4735,N_4720);
or U5366 (N_5366,N_4771,N_4778);
xor U5367 (N_5367,N_4622,N_4992);
nand U5368 (N_5368,N_4848,N_4586);
or U5369 (N_5369,N_4809,N_4968);
xnor U5370 (N_5370,N_4983,N_4945);
nor U5371 (N_5371,N_4625,N_4669);
nand U5372 (N_5372,N_4937,N_4739);
nor U5373 (N_5373,N_4511,N_4517);
or U5374 (N_5374,N_4680,N_4659);
nor U5375 (N_5375,N_4810,N_4756);
nor U5376 (N_5376,N_4780,N_4942);
or U5377 (N_5377,N_4680,N_4988);
nand U5378 (N_5378,N_4555,N_4690);
or U5379 (N_5379,N_4808,N_4541);
and U5380 (N_5380,N_4872,N_4890);
nand U5381 (N_5381,N_4907,N_4565);
nor U5382 (N_5382,N_4849,N_4695);
nor U5383 (N_5383,N_4506,N_4701);
xnor U5384 (N_5384,N_4523,N_4609);
and U5385 (N_5385,N_4706,N_4964);
or U5386 (N_5386,N_4799,N_4877);
xor U5387 (N_5387,N_4895,N_4919);
or U5388 (N_5388,N_4572,N_4552);
and U5389 (N_5389,N_4690,N_4936);
xnor U5390 (N_5390,N_4673,N_4818);
or U5391 (N_5391,N_4713,N_4894);
and U5392 (N_5392,N_4879,N_4587);
xor U5393 (N_5393,N_4856,N_4731);
nor U5394 (N_5394,N_4895,N_4743);
or U5395 (N_5395,N_4979,N_4787);
and U5396 (N_5396,N_4536,N_4999);
nand U5397 (N_5397,N_4846,N_4632);
nand U5398 (N_5398,N_4630,N_4759);
nor U5399 (N_5399,N_4967,N_4765);
or U5400 (N_5400,N_4957,N_4934);
and U5401 (N_5401,N_4539,N_4784);
nor U5402 (N_5402,N_4828,N_4528);
xor U5403 (N_5403,N_4805,N_4812);
or U5404 (N_5404,N_4846,N_4858);
nor U5405 (N_5405,N_4596,N_4938);
or U5406 (N_5406,N_4906,N_4572);
nand U5407 (N_5407,N_4970,N_4593);
and U5408 (N_5408,N_4810,N_4598);
xnor U5409 (N_5409,N_4640,N_4875);
or U5410 (N_5410,N_4996,N_4690);
and U5411 (N_5411,N_4802,N_4613);
nor U5412 (N_5412,N_4866,N_4776);
nor U5413 (N_5413,N_4501,N_4797);
nor U5414 (N_5414,N_4656,N_4674);
nor U5415 (N_5415,N_4802,N_4655);
xnor U5416 (N_5416,N_4577,N_4882);
nand U5417 (N_5417,N_4739,N_4850);
nand U5418 (N_5418,N_4663,N_4980);
or U5419 (N_5419,N_4592,N_4669);
or U5420 (N_5420,N_4866,N_4974);
nor U5421 (N_5421,N_4747,N_4667);
nand U5422 (N_5422,N_4944,N_4889);
or U5423 (N_5423,N_4529,N_4855);
or U5424 (N_5424,N_4938,N_4922);
xor U5425 (N_5425,N_4846,N_4891);
nor U5426 (N_5426,N_4735,N_4871);
and U5427 (N_5427,N_4745,N_4937);
or U5428 (N_5428,N_4750,N_4923);
and U5429 (N_5429,N_4558,N_4782);
nand U5430 (N_5430,N_4755,N_4547);
nor U5431 (N_5431,N_4567,N_4916);
and U5432 (N_5432,N_4840,N_4726);
nand U5433 (N_5433,N_4778,N_4683);
xnor U5434 (N_5434,N_4886,N_4723);
xnor U5435 (N_5435,N_4650,N_4749);
or U5436 (N_5436,N_4989,N_4701);
nor U5437 (N_5437,N_4812,N_4840);
and U5438 (N_5438,N_4811,N_4665);
nor U5439 (N_5439,N_4957,N_4642);
nand U5440 (N_5440,N_4921,N_4819);
or U5441 (N_5441,N_4936,N_4599);
nand U5442 (N_5442,N_4644,N_4971);
nor U5443 (N_5443,N_4854,N_4684);
or U5444 (N_5444,N_4596,N_4500);
or U5445 (N_5445,N_4501,N_4684);
nor U5446 (N_5446,N_4935,N_4822);
nand U5447 (N_5447,N_4801,N_4819);
nor U5448 (N_5448,N_4563,N_4722);
or U5449 (N_5449,N_4551,N_4844);
xnor U5450 (N_5450,N_4767,N_4799);
and U5451 (N_5451,N_4951,N_4701);
or U5452 (N_5452,N_4853,N_4768);
or U5453 (N_5453,N_4532,N_4827);
xor U5454 (N_5454,N_4710,N_4518);
xnor U5455 (N_5455,N_4813,N_4935);
nand U5456 (N_5456,N_4991,N_4830);
and U5457 (N_5457,N_4726,N_4984);
xor U5458 (N_5458,N_4722,N_4509);
xnor U5459 (N_5459,N_4863,N_4676);
nor U5460 (N_5460,N_4674,N_4842);
nand U5461 (N_5461,N_4672,N_4563);
xor U5462 (N_5462,N_4976,N_4833);
nand U5463 (N_5463,N_4995,N_4931);
nor U5464 (N_5464,N_4893,N_4823);
nor U5465 (N_5465,N_4595,N_4570);
nor U5466 (N_5466,N_4511,N_4984);
xnor U5467 (N_5467,N_4984,N_4988);
nor U5468 (N_5468,N_4584,N_4756);
nand U5469 (N_5469,N_4688,N_4804);
and U5470 (N_5470,N_4542,N_4552);
nor U5471 (N_5471,N_4805,N_4775);
nor U5472 (N_5472,N_4619,N_4892);
nand U5473 (N_5473,N_4906,N_4609);
and U5474 (N_5474,N_4658,N_4731);
nor U5475 (N_5475,N_4625,N_4526);
or U5476 (N_5476,N_4517,N_4727);
xor U5477 (N_5477,N_4985,N_4687);
or U5478 (N_5478,N_4774,N_4783);
and U5479 (N_5479,N_4886,N_4976);
xnor U5480 (N_5480,N_4529,N_4837);
xnor U5481 (N_5481,N_4598,N_4545);
xor U5482 (N_5482,N_4599,N_4699);
nor U5483 (N_5483,N_4633,N_4960);
and U5484 (N_5484,N_4871,N_4657);
or U5485 (N_5485,N_4539,N_4533);
nor U5486 (N_5486,N_4607,N_4504);
nor U5487 (N_5487,N_4764,N_4814);
nand U5488 (N_5488,N_4636,N_4720);
or U5489 (N_5489,N_4541,N_4979);
xnor U5490 (N_5490,N_4917,N_4661);
nand U5491 (N_5491,N_4639,N_4538);
and U5492 (N_5492,N_4942,N_4551);
and U5493 (N_5493,N_4672,N_4544);
xnor U5494 (N_5494,N_4621,N_4964);
xor U5495 (N_5495,N_4506,N_4543);
xnor U5496 (N_5496,N_4970,N_4920);
xor U5497 (N_5497,N_4940,N_4567);
nand U5498 (N_5498,N_4615,N_4980);
and U5499 (N_5499,N_4578,N_4774);
and U5500 (N_5500,N_5059,N_5206);
xnor U5501 (N_5501,N_5265,N_5451);
nand U5502 (N_5502,N_5383,N_5327);
and U5503 (N_5503,N_5027,N_5332);
and U5504 (N_5504,N_5227,N_5184);
nand U5505 (N_5505,N_5358,N_5065);
and U5506 (N_5506,N_5448,N_5072);
or U5507 (N_5507,N_5437,N_5414);
xnor U5508 (N_5508,N_5234,N_5142);
or U5509 (N_5509,N_5028,N_5443);
and U5510 (N_5510,N_5097,N_5317);
xor U5511 (N_5511,N_5345,N_5338);
and U5512 (N_5512,N_5203,N_5402);
and U5513 (N_5513,N_5287,N_5409);
or U5514 (N_5514,N_5458,N_5201);
nor U5515 (N_5515,N_5377,N_5374);
xnor U5516 (N_5516,N_5488,N_5013);
nor U5517 (N_5517,N_5223,N_5092);
nand U5518 (N_5518,N_5104,N_5336);
xor U5519 (N_5519,N_5271,N_5038);
nor U5520 (N_5520,N_5387,N_5043);
xor U5521 (N_5521,N_5479,N_5406);
nor U5522 (N_5522,N_5325,N_5042);
nand U5523 (N_5523,N_5121,N_5424);
nor U5524 (N_5524,N_5172,N_5357);
or U5525 (N_5525,N_5470,N_5426);
or U5526 (N_5526,N_5034,N_5207);
and U5527 (N_5527,N_5257,N_5318);
or U5528 (N_5528,N_5083,N_5047);
and U5529 (N_5529,N_5438,N_5453);
and U5530 (N_5530,N_5032,N_5017);
and U5531 (N_5531,N_5471,N_5212);
nand U5532 (N_5532,N_5395,N_5081);
nor U5533 (N_5533,N_5288,N_5280);
nand U5534 (N_5534,N_5302,N_5045);
nand U5535 (N_5535,N_5214,N_5118);
or U5536 (N_5536,N_5159,N_5362);
nor U5537 (N_5537,N_5303,N_5480);
or U5538 (N_5538,N_5127,N_5421);
xor U5539 (N_5539,N_5306,N_5391);
nor U5540 (N_5540,N_5343,N_5132);
nand U5541 (N_5541,N_5068,N_5329);
xor U5542 (N_5542,N_5205,N_5024);
nor U5543 (N_5543,N_5090,N_5269);
xor U5544 (N_5544,N_5260,N_5449);
or U5545 (N_5545,N_5293,N_5139);
nor U5546 (N_5546,N_5394,N_5009);
nor U5547 (N_5547,N_5157,N_5103);
or U5548 (N_5548,N_5093,N_5069);
nand U5549 (N_5549,N_5131,N_5133);
xnor U5550 (N_5550,N_5330,N_5080);
nand U5551 (N_5551,N_5433,N_5169);
or U5552 (N_5552,N_5167,N_5368);
or U5553 (N_5553,N_5099,N_5228);
xor U5554 (N_5554,N_5372,N_5145);
xnor U5555 (N_5555,N_5369,N_5089);
nand U5556 (N_5556,N_5404,N_5188);
xor U5557 (N_5557,N_5185,N_5460);
or U5558 (N_5558,N_5180,N_5040);
nor U5559 (N_5559,N_5225,N_5373);
and U5560 (N_5560,N_5352,N_5146);
xnor U5561 (N_5561,N_5376,N_5183);
nand U5562 (N_5562,N_5209,N_5199);
xnor U5563 (N_5563,N_5001,N_5454);
nand U5564 (N_5564,N_5447,N_5495);
and U5565 (N_5565,N_5224,N_5016);
nor U5566 (N_5566,N_5179,N_5254);
nand U5567 (N_5567,N_5420,N_5096);
nor U5568 (N_5568,N_5305,N_5276);
xnor U5569 (N_5569,N_5173,N_5241);
and U5570 (N_5570,N_5235,N_5450);
or U5571 (N_5571,N_5348,N_5039);
xor U5572 (N_5572,N_5164,N_5396);
or U5573 (N_5573,N_5412,N_5346);
xnor U5574 (N_5574,N_5363,N_5176);
xnor U5575 (N_5575,N_5249,N_5114);
or U5576 (N_5576,N_5434,N_5095);
xnor U5577 (N_5577,N_5217,N_5291);
nor U5578 (N_5578,N_5490,N_5098);
and U5579 (N_5579,N_5378,N_5286);
or U5580 (N_5580,N_5138,N_5380);
nor U5581 (N_5581,N_5469,N_5101);
nand U5582 (N_5582,N_5189,N_5117);
xor U5583 (N_5583,N_5175,N_5314);
nor U5584 (N_5584,N_5401,N_5353);
xnor U5585 (N_5585,N_5337,N_5066);
xnor U5586 (N_5586,N_5370,N_5410);
nor U5587 (N_5587,N_5151,N_5422);
xor U5588 (N_5588,N_5128,N_5025);
xnor U5589 (N_5589,N_5278,N_5459);
nor U5590 (N_5590,N_5486,N_5143);
nand U5591 (N_5591,N_5191,N_5324);
nand U5592 (N_5592,N_5168,N_5386);
xor U5593 (N_5593,N_5148,N_5197);
and U5594 (N_5594,N_5137,N_5171);
nor U5595 (N_5595,N_5279,N_5295);
or U5596 (N_5596,N_5481,N_5186);
or U5597 (N_5597,N_5216,N_5166);
xnor U5598 (N_5598,N_5416,N_5379);
xor U5599 (N_5599,N_5285,N_5273);
and U5600 (N_5600,N_5311,N_5196);
or U5601 (N_5601,N_5026,N_5482);
or U5602 (N_5602,N_5054,N_5489);
nand U5603 (N_5603,N_5382,N_5181);
and U5604 (N_5604,N_5468,N_5229);
and U5605 (N_5605,N_5445,N_5392);
xor U5606 (N_5606,N_5002,N_5244);
or U5607 (N_5607,N_5063,N_5282);
xnor U5608 (N_5608,N_5226,N_5425);
and U5609 (N_5609,N_5156,N_5112);
or U5610 (N_5610,N_5456,N_5094);
nor U5611 (N_5611,N_5497,N_5182);
and U5612 (N_5612,N_5149,N_5023);
and U5613 (N_5613,N_5312,N_5067);
and U5614 (N_5614,N_5411,N_5010);
xor U5615 (N_5615,N_5477,N_5494);
or U5616 (N_5616,N_5105,N_5339);
and U5617 (N_5617,N_5084,N_5270);
and U5618 (N_5618,N_5218,N_5030);
nand U5619 (N_5619,N_5439,N_5060);
and U5620 (N_5620,N_5272,N_5004);
or U5621 (N_5621,N_5408,N_5474);
or U5622 (N_5622,N_5154,N_5008);
nor U5623 (N_5623,N_5077,N_5140);
and U5624 (N_5624,N_5236,N_5195);
or U5625 (N_5625,N_5122,N_5141);
nand U5626 (N_5626,N_5048,N_5087);
xnor U5627 (N_5627,N_5299,N_5487);
nand U5628 (N_5628,N_5334,N_5021);
or U5629 (N_5629,N_5163,N_5165);
and U5630 (N_5630,N_5162,N_5484);
nand U5631 (N_5631,N_5463,N_5022);
nand U5632 (N_5632,N_5116,N_5220);
xor U5633 (N_5633,N_5309,N_5070);
nand U5634 (N_5634,N_5284,N_5135);
nor U5635 (N_5635,N_5233,N_5499);
nor U5636 (N_5636,N_5294,N_5031);
xor U5637 (N_5637,N_5473,N_5413);
xnor U5638 (N_5638,N_5058,N_5230);
or U5639 (N_5639,N_5301,N_5277);
nor U5640 (N_5640,N_5290,N_5385);
xnor U5641 (N_5641,N_5014,N_5431);
or U5642 (N_5642,N_5085,N_5261);
nand U5643 (N_5643,N_5323,N_5100);
or U5644 (N_5644,N_5292,N_5297);
xor U5645 (N_5645,N_5019,N_5457);
nand U5646 (N_5646,N_5354,N_5056);
nand U5647 (N_5647,N_5129,N_5152);
xor U5648 (N_5648,N_5442,N_5136);
nor U5649 (N_5649,N_5111,N_5036);
xnor U5650 (N_5650,N_5005,N_5304);
nor U5651 (N_5651,N_5177,N_5259);
and U5652 (N_5652,N_5478,N_5222);
xor U5653 (N_5653,N_5446,N_5011);
nand U5654 (N_5654,N_5472,N_5384);
nor U5655 (N_5655,N_5365,N_5423);
and U5656 (N_5656,N_5342,N_5455);
nand U5657 (N_5657,N_5018,N_5240);
xor U5658 (N_5658,N_5307,N_5155);
xnor U5659 (N_5659,N_5247,N_5263);
nand U5660 (N_5660,N_5211,N_5476);
nand U5661 (N_5661,N_5262,N_5115);
or U5662 (N_5662,N_5326,N_5267);
nor U5663 (N_5663,N_5427,N_5300);
nor U5664 (N_5664,N_5246,N_5064);
nor U5665 (N_5665,N_5239,N_5316);
nand U5666 (N_5666,N_5091,N_5341);
nand U5667 (N_5667,N_5248,N_5335);
nand U5668 (N_5668,N_5250,N_5086);
nor U5669 (N_5669,N_5243,N_5253);
xnor U5670 (N_5670,N_5071,N_5035);
nand U5671 (N_5671,N_5367,N_5428);
nand U5672 (N_5672,N_5258,N_5242);
or U5673 (N_5673,N_5255,N_5088);
and U5674 (N_5674,N_5440,N_5296);
or U5675 (N_5675,N_5340,N_5388);
nand U5676 (N_5676,N_5381,N_5475);
nand U5677 (N_5677,N_5134,N_5298);
xnor U5678 (N_5678,N_5000,N_5390);
and U5679 (N_5679,N_5397,N_5347);
and U5680 (N_5680,N_5020,N_5275);
nand U5681 (N_5681,N_5078,N_5232);
xor U5682 (N_5682,N_5074,N_5107);
xnor U5683 (N_5683,N_5398,N_5359);
nor U5684 (N_5684,N_5144,N_5328);
nand U5685 (N_5685,N_5485,N_5436);
and U5686 (N_5686,N_5007,N_5208);
xnor U5687 (N_5687,N_5405,N_5464);
nand U5688 (N_5688,N_5268,N_5015);
xor U5689 (N_5689,N_5124,N_5462);
xor U5690 (N_5690,N_5308,N_5213);
nand U5691 (N_5691,N_5106,N_5153);
nor U5692 (N_5692,N_5187,N_5113);
nor U5693 (N_5693,N_5498,N_5194);
xor U5694 (N_5694,N_5356,N_5200);
xor U5695 (N_5695,N_5281,N_5310);
xnor U5696 (N_5696,N_5125,N_5037);
nor U5697 (N_5697,N_5349,N_5256);
nor U5698 (N_5698,N_5466,N_5493);
nand U5699 (N_5699,N_5350,N_5237);
nor U5700 (N_5700,N_5351,N_5215);
nand U5701 (N_5701,N_5366,N_5178);
nand U5702 (N_5702,N_5496,N_5289);
xnor U5703 (N_5703,N_5245,N_5052);
xnor U5704 (N_5704,N_5079,N_5119);
and U5705 (N_5705,N_5319,N_5483);
nor U5706 (N_5706,N_5238,N_5198);
and U5707 (N_5707,N_5221,N_5161);
and U5708 (N_5708,N_5012,N_5429);
and U5709 (N_5709,N_5333,N_5399);
and U5710 (N_5710,N_5061,N_5375);
nand U5711 (N_5711,N_5344,N_5331);
xnor U5712 (N_5712,N_5174,N_5057);
xor U5713 (N_5713,N_5283,N_5400);
or U5714 (N_5714,N_5355,N_5150);
and U5715 (N_5715,N_5322,N_5418);
or U5716 (N_5716,N_5192,N_5044);
and U5717 (N_5717,N_5491,N_5062);
xnor U5718 (N_5718,N_5371,N_5110);
and U5719 (N_5719,N_5160,N_5252);
nand U5720 (N_5720,N_5321,N_5492);
and U5721 (N_5721,N_5202,N_5219);
nor U5722 (N_5722,N_5441,N_5315);
and U5723 (N_5723,N_5006,N_5075);
and U5724 (N_5724,N_5082,N_5403);
nand U5725 (N_5725,N_5461,N_5467);
nor U5726 (N_5726,N_5076,N_5320);
xnor U5727 (N_5727,N_5130,N_5251);
and U5728 (N_5728,N_5266,N_5055);
and U5729 (N_5729,N_5465,N_5430);
or U5730 (N_5730,N_5193,N_5053);
xor U5731 (N_5731,N_5102,N_5147);
and U5732 (N_5732,N_5041,N_5073);
or U5733 (N_5733,N_5190,N_5108);
xor U5734 (N_5734,N_5360,N_5029);
xnor U5735 (N_5735,N_5444,N_5126);
xnor U5736 (N_5736,N_5231,N_5170);
nand U5737 (N_5737,N_5003,N_5046);
xnor U5738 (N_5738,N_5432,N_5452);
and U5739 (N_5739,N_5049,N_5264);
nand U5740 (N_5740,N_5435,N_5393);
nor U5741 (N_5741,N_5313,N_5210);
xnor U5742 (N_5742,N_5120,N_5050);
nor U5743 (N_5743,N_5417,N_5361);
xor U5744 (N_5744,N_5123,N_5407);
or U5745 (N_5745,N_5109,N_5158);
or U5746 (N_5746,N_5274,N_5419);
or U5747 (N_5747,N_5033,N_5389);
or U5748 (N_5748,N_5364,N_5415);
or U5749 (N_5749,N_5204,N_5051);
nand U5750 (N_5750,N_5468,N_5212);
nor U5751 (N_5751,N_5358,N_5441);
nand U5752 (N_5752,N_5361,N_5083);
nor U5753 (N_5753,N_5189,N_5367);
and U5754 (N_5754,N_5259,N_5060);
or U5755 (N_5755,N_5410,N_5002);
nor U5756 (N_5756,N_5195,N_5425);
or U5757 (N_5757,N_5080,N_5054);
nor U5758 (N_5758,N_5129,N_5270);
nor U5759 (N_5759,N_5193,N_5065);
nor U5760 (N_5760,N_5047,N_5436);
nor U5761 (N_5761,N_5346,N_5252);
and U5762 (N_5762,N_5102,N_5182);
or U5763 (N_5763,N_5166,N_5278);
and U5764 (N_5764,N_5333,N_5177);
nand U5765 (N_5765,N_5325,N_5285);
nor U5766 (N_5766,N_5102,N_5473);
or U5767 (N_5767,N_5488,N_5426);
nand U5768 (N_5768,N_5394,N_5385);
nand U5769 (N_5769,N_5477,N_5303);
or U5770 (N_5770,N_5376,N_5219);
or U5771 (N_5771,N_5349,N_5258);
nand U5772 (N_5772,N_5053,N_5451);
or U5773 (N_5773,N_5116,N_5493);
xor U5774 (N_5774,N_5397,N_5432);
nand U5775 (N_5775,N_5043,N_5211);
or U5776 (N_5776,N_5214,N_5149);
or U5777 (N_5777,N_5204,N_5293);
nor U5778 (N_5778,N_5270,N_5291);
nor U5779 (N_5779,N_5206,N_5346);
or U5780 (N_5780,N_5147,N_5414);
nand U5781 (N_5781,N_5448,N_5276);
nand U5782 (N_5782,N_5141,N_5478);
nand U5783 (N_5783,N_5247,N_5310);
nand U5784 (N_5784,N_5380,N_5007);
and U5785 (N_5785,N_5087,N_5137);
nand U5786 (N_5786,N_5076,N_5412);
and U5787 (N_5787,N_5181,N_5486);
and U5788 (N_5788,N_5117,N_5273);
nand U5789 (N_5789,N_5223,N_5247);
xor U5790 (N_5790,N_5186,N_5202);
xnor U5791 (N_5791,N_5048,N_5403);
xor U5792 (N_5792,N_5495,N_5257);
and U5793 (N_5793,N_5305,N_5085);
and U5794 (N_5794,N_5401,N_5066);
or U5795 (N_5795,N_5374,N_5456);
and U5796 (N_5796,N_5486,N_5275);
or U5797 (N_5797,N_5158,N_5191);
nand U5798 (N_5798,N_5321,N_5155);
and U5799 (N_5799,N_5365,N_5276);
nor U5800 (N_5800,N_5206,N_5162);
xnor U5801 (N_5801,N_5190,N_5279);
and U5802 (N_5802,N_5251,N_5133);
or U5803 (N_5803,N_5467,N_5004);
or U5804 (N_5804,N_5317,N_5499);
and U5805 (N_5805,N_5481,N_5436);
or U5806 (N_5806,N_5068,N_5491);
nand U5807 (N_5807,N_5236,N_5064);
xor U5808 (N_5808,N_5267,N_5149);
xor U5809 (N_5809,N_5250,N_5478);
nand U5810 (N_5810,N_5310,N_5254);
nand U5811 (N_5811,N_5471,N_5136);
nand U5812 (N_5812,N_5347,N_5316);
nor U5813 (N_5813,N_5019,N_5465);
nor U5814 (N_5814,N_5315,N_5458);
or U5815 (N_5815,N_5355,N_5346);
nor U5816 (N_5816,N_5448,N_5252);
or U5817 (N_5817,N_5345,N_5302);
and U5818 (N_5818,N_5214,N_5318);
nor U5819 (N_5819,N_5346,N_5301);
and U5820 (N_5820,N_5160,N_5477);
or U5821 (N_5821,N_5070,N_5079);
xor U5822 (N_5822,N_5152,N_5450);
and U5823 (N_5823,N_5014,N_5339);
xor U5824 (N_5824,N_5169,N_5235);
or U5825 (N_5825,N_5389,N_5069);
or U5826 (N_5826,N_5457,N_5469);
nand U5827 (N_5827,N_5478,N_5055);
and U5828 (N_5828,N_5365,N_5146);
nand U5829 (N_5829,N_5378,N_5323);
nor U5830 (N_5830,N_5464,N_5239);
or U5831 (N_5831,N_5255,N_5490);
nor U5832 (N_5832,N_5277,N_5124);
nor U5833 (N_5833,N_5306,N_5318);
nand U5834 (N_5834,N_5248,N_5035);
nand U5835 (N_5835,N_5124,N_5030);
or U5836 (N_5836,N_5064,N_5022);
nand U5837 (N_5837,N_5160,N_5014);
and U5838 (N_5838,N_5440,N_5142);
nand U5839 (N_5839,N_5158,N_5232);
nand U5840 (N_5840,N_5047,N_5048);
nor U5841 (N_5841,N_5378,N_5424);
nor U5842 (N_5842,N_5069,N_5204);
nor U5843 (N_5843,N_5283,N_5059);
nor U5844 (N_5844,N_5192,N_5339);
nand U5845 (N_5845,N_5489,N_5081);
nand U5846 (N_5846,N_5063,N_5248);
nor U5847 (N_5847,N_5416,N_5220);
xor U5848 (N_5848,N_5095,N_5324);
or U5849 (N_5849,N_5029,N_5165);
nor U5850 (N_5850,N_5214,N_5444);
nor U5851 (N_5851,N_5180,N_5468);
xnor U5852 (N_5852,N_5396,N_5108);
and U5853 (N_5853,N_5037,N_5159);
nand U5854 (N_5854,N_5366,N_5189);
or U5855 (N_5855,N_5100,N_5005);
and U5856 (N_5856,N_5329,N_5484);
or U5857 (N_5857,N_5093,N_5274);
or U5858 (N_5858,N_5252,N_5229);
nand U5859 (N_5859,N_5486,N_5256);
xor U5860 (N_5860,N_5493,N_5328);
nor U5861 (N_5861,N_5099,N_5113);
and U5862 (N_5862,N_5497,N_5390);
or U5863 (N_5863,N_5091,N_5358);
xnor U5864 (N_5864,N_5403,N_5068);
or U5865 (N_5865,N_5248,N_5455);
or U5866 (N_5866,N_5046,N_5026);
or U5867 (N_5867,N_5185,N_5056);
xor U5868 (N_5868,N_5116,N_5395);
xor U5869 (N_5869,N_5157,N_5116);
nor U5870 (N_5870,N_5147,N_5439);
or U5871 (N_5871,N_5396,N_5057);
xnor U5872 (N_5872,N_5094,N_5220);
nor U5873 (N_5873,N_5153,N_5096);
nand U5874 (N_5874,N_5371,N_5059);
xnor U5875 (N_5875,N_5492,N_5326);
and U5876 (N_5876,N_5256,N_5023);
nor U5877 (N_5877,N_5465,N_5084);
or U5878 (N_5878,N_5390,N_5429);
nand U5879 (N_5879,N_5372,N_5261);
nand U5880 (N_5880,N_5285,N_5319);
xor U5881 (N_5881,N_5290,N_5024);
nand U5882 (N_5882,N_5395,N_5067);
nor U5883 (N_5883,N_5245,N_5400);
nand U5884 (N_5884,N_5397,N_5278);
xor U5885 (N_5885,N_5261,N_5242);
and U5886 (N_5886,N_5271,N_5420);
and U5887 (N_5887,N_5298,N_5105);
nand U5888 (N_5888,N_5072,N_5423);
and U5889 (N_5889,N_5265,N_5013);
nand U5890 (N_5890,N_5204,N_5326);
nor U5891 (N_5891,N_5292,N_5381);
nor U5892 (N_5892,N_5216,N_5347);
and U5893 (N_5893,N_5170,N_5341);
xnor U5894 (N_5894,N_5028,N_5280);
xnor U5895 (N_5895,N_5297,N_5003);
nor U5896 (N_5896,N_5337,N_5467);
and U5897 (N_5897,N_5305,N_5233);
and U5898 (N_5898,N_5096,N_5068);
and U5899 (N_5899,N_5341,N_5291);
and U5900 (N_5900,N_5383,N_5334);
nor U5901 (N_5901,N_5009,N_5358);
or U5902 (N_5902,N_5318,N_5042);
nand U5903 (N_5903,N_5175,N_5495);
nand U5904 (N_5904,N_5058,N_5195);
nor U5905 (N_5905,N_5324,N_5138);
xnor U5906 (N_5906,N_5273,N_5421);
nor U5907 (N_5907,N_5459,N_5297);
and U5908 (N_5908,N_5465,N_5257);
nor U5909 (N_5909,N_5108,N_5238);
nand U5910 (N_5910,N_5359,N_5297);
and U5911 (N_5911,N_5285,N_5022);
nor U5912 (N_5912,N_5468,N_5463);
or U5913 (N_5913,N_5389,N_5084);
nand U5914 (N_5914,N_5171,N_5204);
and U5915 (N_5915,N_5045,N_5245);
and U5916 (N_5916,N_5141,N_5260);
xnor U5917 (N_5917,N_5477,N_5294);
nand U5918 (N_5918,N_5250,N_5333);
xor U5919 (N_5919,N_5380,N_5122);
or U5920 (N_5920,N_5327,N_5330);
xor U5921 (N_5921,N_5435,N_5156);
nand U5922 (N_5922,N_5337,N_5196);
xor U5923 (N_5923,N_5275,N_5225);
nand U5924 (N_5924,N_5447,N_5468);
xor U5925 (N_5925,N_5073,N_5052);
and U5926 (N_5926,N_5030,N_5085);
or U5927 (N_5927,N_5452,N_5122);
xor U5928 (N_5928,N_5254,N_5141);
nand U5929 (N_5929,N_5441,N_5335);
nor U5930 (N_5930,N_5375,N_5163);
nand U5931 (N_5931,N_5191,N_5463);
xor U5932 (N_5932,N_5351,N_5257);
or U5933 (N_5933,N_5160,N_5010);
nand U5934 (N_5934,N_5196,N_5320);
or U5935 (N_5935,N_5142,N_5496);
and U5936 (N_5936,N_5025,N_5443);
and U5937 (N_5937,N_5268,N_5136);
xor U5938 (N_5938,N_5397,N_5473);
nor U5939 (N_5939,N_5073,N_5196);
xor U5940 (N_5940,N_5395,N_5001);
nor U5941 (N_5941,N_5460,N_5382);
nand U5942 (N_5942,N_5445,N_5473);
and U5943 (N_5943,N_5024,N_5054);
xor U5944 (N_5944,N_5490,N_5010);
nand U5945 (N_5945,N_5454,N_5292);
xor U5946 (N_5946,N_5309,N_5495);
nor U5947 (N_5947,N_5074,N_5041);
nand U5948 (N_5948,N_5120,N_5398);
or U5949 (N_5949,N_5459,N_5225);
nor U5950 (N_5950,N_5116,N_5124);
xor U5951 (N_5951,N_5348,N_5383);
xnor U5952 (N_5952,N_5162,N_5050);
xor U5953 (N_5953,N_5385,N_5444);
nor U5954 (N_5954,N_5122,N_5212);
xor U5955 (N_5955,N_5337,N_5312);
and U5956 (N_5956,N_5462,N_5388);
and U5957 (N_5957,N_5301,N_5201);
and U5958 (N_5958,N_5103,N_5416);
nor U5959 (N_5959,N_5075,N_5303);
xor U5960 (N_5960,N_5110,N_5314);
and U5961 (N_5961,N_5170,N_5392);
or U5962 (N_5962,N_5110,N_5320);
or U5963 (N_5963,N_5099,N_5097);
or U5964 (N_5964,N_5233,N_5104);
nand U5965 (N_5965,N_5308,N_5177);
xnor U5966 (N_5966,N_5287,N_5088);
xor U5967 (N_5967,N_5366,N_5351);
nor U5968 (N_5968,N_5449,N_5337);
or U5969 (N_5969,N_5207,N_5384);
or U5970 (N_5970,N_5403,N_5465);
nor U5971 (N_5971,N_5468,N_5093);
nor U5972 (N_5972,N_5378,N_5161);
and U5973 (N_5973,N_5382,N_5435);
xor U5974 (N_5974,N_5114,N_5338);
nand U5975 (N_5975,N_5312,N_5202);
nand U5976 (N_5976,N_5373,N_5241);
nor U5977 (N_5977,N_5312,N_5361);
and U5978 (N_5978,N_5318,N_5457);
nand U5979 (N_5979,N_5365,N_5056);
nand U5980 (N_5980,N_5411,N_5175);
xor U5981 (N_5981,N_5183,N_5238);
or U5982 (N_5982,N_5218,N_5288);
nor U5983 (N_5983,N_5207,N_5458);
nor U5984 (N_5984,N_5143,N_5208);
or U5985 (N_5985,N_5349,N_5219);
nand U5986 (N_5986,N_5156,N_5153);
or U5987 (N_5987,N_5090,N_5106);
or U5988 (N_5988,N_5264,N_5335);
and U5989 (N_5989,N_5494,N_5394);
nand U5990 (N_5990,N_5437,N_5355);
nand U5991 (N_5991,N_5125,N_5179);
and U5992 (N_5992,N_5074,N_5424);
nand U5993 (N_5993,N_5139,N_5085);
xor U5994 (N_5994,N_5323,N_5366);
nor U5995 (N_5995,N_5161,N_5285);
xnor U5996 (N_5996,N_5362,N_5041);
xnor U5997 (N_5997,N_5228,N_5072);
and U5998 (N_5998,N_5155,N_5344);
nand U5999 (N_5999,N_5339,N_5393);
and U6000 (N_6000,N_5533,N_5656);
nor U6001 (N_6001,N_5974,N_5815);
nand U6002 (N_6002,N_5769,N_5582);
nor U6003 (N_6003,N_5876,N_5632);
nor U6004 (N_6004,N_5862,N_5960);
xnor U6005 (N_6005,N_5861,N_5562);
nand U6006 (N_6006,N_5528,N_5848);
xnor U6007 (N_6007,N_5684,N_5685);
and U6008 (N_6008,N_5933,N_5972);
or U6009 (N_6009,N_5732,N_5995);
nand U6010 (N_6010,N_5761,N_5673);
xnor U6011 (N_6011,N_5926,N_5942);
and U6012 (N_6012,N_5838,N_5696);
or U6013 (N_6013,N_5931,N_5625);
nor U6014 (N_6014,N_5921,N_5952);
nand U6015 (N_6015,N_5789,N_5904);
nor U6016 (N_6016,N_5882,N_5885);
nand U6017 (N_6017,N_5634,N_5527);
xor U6018 (N_6018,N_5713,N_5664);
nand U6019 (N_6019,N_5585,N_5944);
nand U6020 (N_6020,N_5653,N_5660);
xor U6021 (N_6021,N_5801,N_5538);
nor U6022 (N_6022,N_5677,N_5821);
nor U6023 (N_6023,N_5524,N_5907);
nand U6024 (N_6024,N_5503,N_5934);
nand U6025 (N_6025,N_5791,N_5602);
nor U6026 (N_6026,N_5768,N_5786);
or U6027 (N_6027,N_5520,N_5557);
nand U6028 (N_6028,N_5780,N_5607);
nor U6029 (N_6029,N_5820,N_5980);
nor U6030 (N_6030,N_5908,N_5554);
xnor U6031 (N_6031,N_5877,N_5746);
nor U6032 (N_6032,N_5999,N_5819);
nor U6033 (N_6033,N_5920,N_5806);
and U6034 (N_6034,N_5630,N_5911);
and U6035 (N_6035,N_5730,N_5612);
nor U6036 (N_6036,N_5729,N_5679);
nor U6037 (N_6037,N_5967,N_5597);
and U6038 (N_6038,N_5758,N_5866);
or U6039 (N_6039,N_5859,N_5515);
and U6040 (N_6040,N_5704,N_5894);
and U6041 (N_6041,N_5833,N_5683);
or U6042 (N_6042,N_5940,N_5832);
xnor U6043 (N_6043,N_5519,N_5643);
xor U6044 (N_6044,N_5521,N_5808);
and U6045 (N_6045,N_5903,N_5924);
and U6046 (N_6046,N_5662,N_5760);
or U6047 (N_6047,N_5539,N_5626);
or U6048 (N_6048,N_5666,N_5797);
or U6049 (N_6049,N_5724,N_5970);
xor U6050 (N_6050,N_5818,N_5592);
xnor U6051 (N_6051,N_5959,N_5541);
and U6052 (N_6052,N_5707,N_5689);
and U6053 (N_6053,N_5743,N_5896);
nor U6054 (N_6054,N_5558,N_5699);
and U6055 (N_6055,N_5556,N_5657);
or U6056 (N_6056,N_5932,N_5793);
or U6057 (N_6057,N_5963,N_5681);
and U6058 (N_6058,N_5802,N_5694);
and U6059 (N_6059,N_5796,N_5545);
nand U6060 (N_6060,N_5914,N_5693);
nand U6061 (N_6061,N_5839,N_5869);
nand U6062 (N_6062,N_5569,N_5883);
or U6063 (N_6063,N_5635,N_5517);
or U6064 (N_6064,N_5608,N_5993);
and U6065 (N_6065,N_5956,N_5864);
nand U6066 (N_6066,N_5845,N_5502);
nor U6067 (N_6067,N_5831,N_5510);
or U6068 (N_6068,N_5709,N_5698);
xor U6069 (N_6069,N_5898,N_5955);
and U6070 (N_6070,N_5733,N_5575);
nor U6071 (N_6071,N_5826,N_5957);
nand U6072 (N_6072,N_5773,N_5890);
or U6073 (N_6073,N_5688,N_5697);
or U6074 (N_6074,N_5771,N_5714);
nand U6075 (N_6075,N_5954,N_5621);
or U6076 (N_6076,N_5588,N_5830);
and U6077 (N_6077,N_5923,N_5583);
and U6078 (N_6078,N_5649,N_5794);
nor U6079 (N_6079,N_5619,N_5889);
and U6080 (N_6080,N_5540,N_5675);
nor U6081 (N_6081,N_5984,N_5770);
xor U6082 (N_6082,N_5580,N_5912);
and U6083 (N_6083,N_5508,N_5599);
or U6084 (N_6084,N_5928,N_5576);
and U6085 (N_6085,N_5814,N_5505);
or U6086 (N_6086,N_5750,N_5631);
or U6087 (N_6087,N_5740,N_5899);
and U6088 (N_6088,N_5561,N_5902);
or U6089 (N_6089,N_5706,N_5950);
nor U6090 (N_6090,N_5840,N_5629);
nor U6091 (N_6091,N_5586,N_5572);
nand U6092 (N_6092,N_5712,N_5616);
nand U6093 (N_6093,N_5705,N_5738);
nor U6094 (N_6094,N_5927,N_5905);
or U6095 (N_6095,N_5553,N_5687);
nand U6096 (N_6096,N_5717,N_5555);
or U6097 (N_6097,N_5915,N_5971);
nand U6098 (N_6098,N_5951,N_5596);
and U6099 (N_6099,N_5594,N_5731);
nand U6100 (N_6100,N_5860,N_5560);
nor U6101 (N_6101,N_5804,N_5529);
or U6102 (N_6102,N_5721,N_5506);
and U6103 (N_6103,N_5711,N_5728);
xnor U6104 (N_6104,N_5982,N_5975);
or U6105 (N_6105,N_5670,N_5996);
or U6106 (N_6106,N_5638,N_5754);
xnor U6107 (N_6107,N_5736,N_5930);
and U6108 (N_6108,N_5851,N_5537);
or U6109 (N_6109,N_5719,N_5739);
xor U6110 (N_6110,N_5535,N_5800);
and U6111 (N_6111,N_5976,N_5642);
nor U6112 (N_6112,N_5946,N_5567);
xor U6113 (N_6113,N_5941,N_5737);
xnor U6114 (N_6114,N_5991,N_5901);
xor U6115 (N_6115,N_5986,N_5628);
nor U6116 (N_6116,N_5548,N_5753);
xor U6117 (N_6117,N_5803,N_5525);
or U6118 (N_6118,N_5606,N_5741);
and U6119 (N_6119,N_5601,N_5522);
nor U6120 (N_6120,N_5526,N_5849);
xnor U6121 (N_6121,N_5501,N_5661);
nand U6122 (N_6122,N_5584,N_5891);
nand U6123 (N_6123,N_5735,N_5600);
nor U6124 (N_6124,N_5672,N_5658);
or U6125 (N_6125,N_5825,N_5591);
nor U6126 (N_6126,N_5563,N_5674);
nor U6127 (N_6127,N_5775,N_5659);
xor U6128 (N_6128,N_5722,N_5847);
nor U6129 (N_6129,N_5922,N_5604);
nor U6130 (N_6130,N_5756,N_5841);
nor U6131 (N_6131,N_5858,N_5647);
and U6132 (N_6132,N_5766,N_5570);
or U6133 (N_6133,N_5726,N_5764);
and U6134 (N_6134,N_5663,N_5835);
nor U6135 (N_6135,N_5690,N_5985);
or U6136 (N_6136,N_5551,N_5822);
xnor U6137 (N_6137,N_5917,N_5874);
and U6138 (N_6138,N_5611,N_5948);
nand U6139 (N_6139,N_5834,N_5617);
xnor U6140 (N_6140,N_5813,N_5645);
nand U6141 (N_6141,N_5752,N_5992);
or U6142 (N_6142,N_5990,N_5929);
nor U6143 (N_6143,N_5938,N_5574);
or U6144 (N_6144,N_5745,N_5700);
nor U6145 (N_6145,N_5846,N_5962);
or U6146 (N_6146,N_5667,N_5623);
and U6147 (N_6147,N_5777,N_5895);
xor U6148 (N_6148,N_5781,N_5610);
and U6149 (N_6149,N_5725,N_5913);
nor U6150 (N_6150,N_5983,N_5590);
nand U6151 (N_6151,N_5865,N_5511);
xor U6152 (N_6152,N_5857,N_5509);
xor U6153 (N_6153,N_5897,N_5816);
or U6154 (N_6154,N_5961,N_5772);
or U6155 (N_6155,N_5978,N_5828);
nor U6156 (N_6156,N_5886,N_5748);
nor U6157 (N_6157,N_5641,N_5549);
nor U6158 (N_6158,N_5947,N_5867);
xnor U6159 (N_6159,N_5755,N_5784);
nand U6160 (N_6160,N_5836,N_5843);
nand U6161 (N_6161,N_5581,N_5720);
or U6162 (N_6162,N_5817,N_5723);
xnor U6163 (N_6163,N_5514,N_5906);
or U6164 (N_6164,N_5881,N_5795);
nand U6165 (N_6165,N_5778,N_5531);
xnor U6166 (N_6166,N_5964,N_5682);
or U6167 (N_6167,N_5516,N_5523);
nor U6168 (N_6168,N_5937,N_5759);
and U6169 (N_6169,N_5747,N_5863);
nor U6170 (N_6170,N_5751,N_5650);
xnor U6171 (N_6171,N_5648,N_5577);
nor U6172 (N_6172,N_5762,N_5757);
or U6173 (N_6173,N_5850,N_5564);
and U6174 (N_6174,N_5716,N_5613);
nor U6175 (N_6175,N_5744,N_5870);
nor U6176 (N_6176,N_5918,N_5695);
nor U6177 (N_6177,N_5609,N_5703);
xnor U6178 (N_6178,N_5550,N_5598);
xor U6179 (N_6179,N_5678,N_5779);
and U6180 (N_6180,N_5568,N_5546);
and U6181 (N_6181,N_5998,N_5639);
nand U6182 (N_6182,N_5844,N_5742);
nor U6183 (N_6183,N_5878,N_5969);
nand U6184 (N_6184,N_5792,N_5783);
xnor U6185 (N_6185,N_5812,N_5652);
or U6186 (N_6186,N_5798,N_5676);
or U6187 (N_6187,N_5566,N_5871);
or U6188 (N_6188,N_5710,N_5827);
or U6189 (N_6189,N_5979,N_5749);
or U6190 (N_6190,N_5855,N_5782);
nand U6191 (N_6191,N_5935,N_5587);
nand U6192 (N_6192,N_5785,N_5953);
xor U6193 (N_6193,N_5893,N_5776);
or U6194 (N_6194,N_5949,N_5680);
nand U6195 (N_6195,N_5790,N_5977);
or U6196 (N_6196,N_5853,N_5842);
nand U6197 (N_6197,N_5603,N_5987);
nand U6198 (N_6198,N_5981,N_5943);
or U6199 (N_6199,N_5936,N_5966);
nor U6200 (N_6200,N_5856,N_5542);
nand U6201 (N_6201,N_5973,N_5512);
nor U6202 (N_6202,N_5945,N_5559);
xor U6203 (N_6203,N_5655,N_5787);
nor U6204 (N_6204,N_5875,N_5734);
nor U6205 (N_6205,N_5854,N_5686);
and U6206 (N_6206,N_5810,N_5605);
or U6207 (N_6207,N_5988,N_5788);
nor U6208 (N_6208,N_5805,N_5637);
xor U6209 (N_6209,N_5532,N_5765);
nor U6210 (N_6210,N_5873,N_5708);
or U6211 (N_6211,N_5852,N_5888);
nand U6212 (N_6212,N_5671,N_5571);
xor U6213 (N_6213,N_5919,N_5900);
nand U6214 (N_6214,N_5593,N_5892);
or U6215 (N_6215,N_5884,N_5958);
xnor U6216 (N_6216,N_5692,N_5518);
or U6217 (N_6217,N_5887,N_5573);
and U6218 (N_6218,N_5763,N_5552);
and U6219 (N_6219,N_5702,N_5651);
nand U6220 (N_6220,N_5644,N_5640);
nor U6221 (N_6221,N_5799,N_5534);
nor U6222 (N_6222,N_5727,N_5579);
xnor U6223 (N_6223,N_5824,N_5595);
nand U6224 (N_6224,N_5691,N_5622);
or U6225 (N_6225,N_5615,N_5880);
or U6226 (N_6226,N_5767,N_5774);
and U6227 (N_6227,N_5636,N_5618);
and U6228 (N_6228,N_5939,N_5868);
nand U6229 (N_6229,N_5589,N_5654);
nor U6230 (N_6230,N_5823,N_5624);
xor U6231 (N_6231,N_5669,N_5997);
nand U6232 (N_6232,N_5718,N_5909);
and U6233 (N_6233,N_5627,N_5701);
or U6234 (N_6234,N_5837,N_5665);
xor U6235 (N_6235,N_5994,N_5620);
nor U6236 (N_6236,N_5530,N_5910);
nor U6237 (N_6237,N_5925,N_5543);
or U6238 (N_6238,N_5507,N_5989);
and U6239 (N_6239,N_5829,N_5504);
and U6240 (N_6240,N_5544,N_5916);
and U6241 (N_6241,N_5811,N_5872);
nor U6242 (N_6242,N_5500,N_5807);
and U6243 (N_6243,N_5715,N_5513);
nand U6244 (N_6244,N_5668,N_5879);
or U6245 (N_6245,N_5968,N_5809);
xnor U6246 (N_6246,N_5565,N_5536);
or U6247 (N_6247,N_5578,N_5614);
or U6248 (N_6248,N_5646,N_5633);
xor U6249 (N_6249,N_5965,N_5547);
and U6250 (N_6250,N_5747,N_5506);
and U6251 (N_6251,N_5631,N_5673);
and U6252 (N_6252,N_5904,N_5635);
or U6253 (N_6253,N_5500,N_5707);
and U6254 (N_6254,N_5593,N_5902);
xor U6255 (N_6255,N_5895,N_5826);
nand U6256 (N_6256,N_5533,N_5679);
or U6257 (N_6257,N_5741,N_5988);
and U6258 (N_6258,N_5672,N_5931);
nand U6259 (N_6259,N_5947,N_5665);
xor U6260 (N_6260,N_5807,N_5561);
nor U6261 (N_6261,N_5866,N_5844);
and U6262 (N_6262,N_5508,N_5946);
or U6263 (N_6263,N_5532,N_5828);
and U6264 (N_6264,N_5509,N_5710);
nand U6265 (N_6265,N_5515,N_5880);
nor U6266 (N_6266,N_5835,N_5823);
nor U6267 (N_6267,N_5706,N_5850);
xnor U6268 (N_6268,N_5985,N_5830);
xnor U6269 (N_6269,N_5884,N_5955);
xor U6270 (N_6270,N_5585,N_5718);
xor U6271 (N_6271,N_5544,N_5723);
or U6272 (N_6272,N_5500,N_5598);
nor U6273 (N_6273,N_5977,N_5990);
xnor U6274 (N_6274,N_5988,N_5664);
xor U6275 (N_6275,N_5899,N_5795);
xor U6276 (N_6276,N_5947,N_5732);
xor U6277 (N_6277,N_5618,N_5896);
or U6278 (N_6278,N_5553,N_5823);
nor U6279 (N_6279,N_5795,N_5999);
nand U6280 (N_6280,N_5557,N_5672);
nand U6281 (N_6281,N_5604,N_5729);
xor U6282 (N_6282,N_5701,N_5863);
nor U6283 (N_6283,N_5554,N_5696);
nand U6284 (N_6284,N_5738,N_5782);
or U6285 (N_6285,N_5663,N_5627);
nor U6286 (N_6286,N_5982,N_5506);
nor U6287 (N_6287,N_5788,N_5823);
and U6288 (N_6288,N_5807,N_5925);
nand U6289 (N_6289,N_5920,N_5988);
nand U6290 (N_6290,N_5832,N_5521);
and U6291 (N_6291,N_5860,N_5935);
and U6292 (N_6292,N_5591,N_5751);
or U6293 (N_6293,N_5723,N_5610);
nor U6294 (N_6294,N_5634,N_5501);
and U6295 (N_6295,N_5935,N_5572);
and U6296 (N_6296,N_5852,N_5904);
or U6297 (N_6297,N_5640,N_5605);
and U6298 (N_6298,N_5811,N_5784);
and U6299 (N_6299,N_5504,N_5963);
nor U6300 (N_6300,N_5717,N_5904);
or U6301 (N_6301,N_5949,N_5662);
or U6302 (N_6302,N_5727,N_5546);
nor U6303 (N_6303,N_5515,N_5757);
nor U6304 (N_6304,N_5920,N_5565);
nand U6305 (N_6305,N_5838,N_5615);
xnor U6306 (N_6306,N_5580,N_5668);
or U6307 (N_6307,N_5844,N_5916);
nand U6308 (N_6308,N_5976,N_5791);
nor U6309 (N_6309,N_5635,N_5925);
nand U6310 (N_6310,N_5792,N_5868);
nand U6311 (N_6311,N_5539,N_5536);
xor U6312 (N_6312,N_5962,N_5820);
nand U6313 (N_6313,N_5538,N_5513);
and U6314 (N_6314,N_5665,N_5869);
nand U6315 (N_6315,N_5729,N_5991);
nor U6316 (N_6316,N_5940,N_5828);
and U6317 (N_6317,N_5965,N_5673);
or U6318 (N_6318,N_5857,N_5641);
nand U6319 (N_6319,N_5674,N_5967);
or U6320 (N_6320,N_5793,N_5603);
or U6321 (N_6321,N_5821,N_5622);
and U6322 (N_6322,N_5520,N_5920);
nand U6323 (N_6323,N_5966,N_5948);
nand U6324 (N_6324,N_5760,N_5769);
nor U6325 (N_6325,N_5770,N_5564);
xnor U6326 (N_6326,N_5705,N_5922);
or U6327 (N_6327,N_5812,N_5996);
xor U6328 (N_6328,N_5882,N_5677);
xnor U6329 (N_6329,N_5891,N_5887);
or U6330 (N_6330,N_5818,N_5652);
or U6331 (N_6331,N_5874,N_5611);
or U6332 (N_6332,N_5986,N_5721);
or U6333 (N_6333,N_5715,N_5548);
and U6334 (N_6334,N_5625,N_5671);
nand U6335 (N_6335,N_5766,N_5605);
nand U6336 (N_6336,N_5574,N_5504);
or U6337 (N_6337,N_5690,N_5755);
xnor U6338 (N_6338,N_5546,N_5786);
xor U6339 (N_6339,N_5702,N_5772);
and U6340 (N_6340,N_5698,N_5818);
or U6341 (N_6341,N_5629,N_5881);
nor U6342 (N_6342,N_5579,N_5800);
xor U6343 (N_6343,N_5852,N_5868);
nor U6344 (N_6344,N_5597,N_5530);
nor U6345 (N_6345,N_5685,N_5995);
xnor U6346 (N_6346,N_5613,N_5586);
nor U6347 (N_6347,N_5613,N_5868);
xnor U6348 (N_6348,N_5776,N_5884);
and U6349 (N_6349,N_5684,N_5566);
or U6350 (N_6350,N_5673,N_5749);
or U6351 (N_6351,N_5719,N_5895);
or U6352 (N_6352,N_5715,N_5752);
nand U6353 (N_6353,N_5795,N_5504);
and U6354 (N_6354,N_5874,N_5550);
xor U6355 (N_6355,N_5587,N_5709);
nor U6356 (N_6356,N_5732,N_5939);
nor U6357 (N_6357,N_5887,N_5514);
xnor U6358 (N_6358,N_5579,N_5620);
nor U6359 (N_6359,N_5558,N_5529);
and U6360 (N_6360,N_5806,N_5771);
nor U6361 (N_6361,N_5654,N_5745);
nand U6362 (N_6362,N_5720,N_5696);
and U6363 (N_6363,N_5986,N_5517);
and U6364 (N_6364,N_5514,N_5742);
or U6365 (N_6365,N_5645,N_5808);
or U6366 (N_6366,N_5986,N_5723);
or U6367 (N_6367,N_5798,N_5657);
nor U6368 (N_6368,N_5767,N_5789);
nand U6369 (N_6369,N_5531,N_5686);
or U6370 (N_6370,N_5824,N_5729);
nor U6371 (N_6371,N_5969,N_5716);
nand U6372 (N_6372,N_5844,N_5562);
and U6373 (N_6373,N_5980,N_5895);
nand U6374 (N_6374,N_5756,N_5911);
nor U6375 (N_6375,N_5518,N_5793);
and U6376 (N_6376,N_5859,N_5898);
nor U6377 (N_6377,N_5932,N_5608);
nand U6378 (N_6378,N_5533,N_5516);
or U6379 (N_6379,N_5505,N_5751);
xnor U6380 (N_6380,N_5528,N_5786);
and U6381 (N_6381,N_5689,N_5985);
xnor U6382 (N_6382,N_5637,N_5680);
and U6383 (N_6383,N_5805,N_5674);
nand U6384 (N_6384,N_5729,N_5701);
nand U6385 (N_6385,N_5982,N_5754);
xnor U6386 (N_6386,N_5514,N_5950);
xnor U6387 (N_6387,N_5686,N_5602);
nand U6388 (N_6388,N_5751,N_5560);
xnor U6389 (N_6389,N_5755,N_5857);
nor U6390 (N_6390,N_5971,N_5595);
nand U6391 (N_6391,N_5778,N_5931);
xnor U6392 (N_6392,N_5632,N_5842);
nand U6393 (N_6393,N_5699,N_5747);
nand U6394 (N_6394,N_5855,N_5792);
xnor U6395 (N_6395,N_5679,N_5884);
and U6396 (N_6396,N_5681,N_5538);
xnor U6397 (N_6397,N_5761,N_5781);
nand U6398 (N_6398,N_5926,N_5980);
and U6399 (N_6399,N_5767,N_5917);
nor U6400 (N_6400,N_5783,N_5555);
xnor U6401 (N_6401,N_5716,N_5592);
and U6402 (N_6402,N_5866,N_5679);
or U6403 (N_6403,N_5718,N_5829);
or U6404 (N_6404,N_5519,N_5554);
or U6405 (N_6405,N_5680,N_5615);
and U6406 (N_6406,N_5836,N_5688);
or U6407 (N_6407,N_5589,N_5769);
xnor U6408 (N_6408,N_5543,N_5650);
nand U6409 (N_6409,N_5735,N_5840);
xor U6410 (N_6410,N_5910,N_5695);
nor U6411 (N_6411,N_5896,N_5878);
or U6412 (N_6412,N_5733,N_5623);
or U6413 (N_6413,N_5849,N_5903);
and U6414 (N_6414,N_5765,N_5660);
nand U6415 (N_6415,N_5748,N_5929);
and U6416 (N_6416,N_5559,N_5717);
and U6417 (N_6417,N_5513,N_5537);
or U6418 (N_6418,N_5844,N_5529);
nor U6419 (N_6419,N_5794,N_5777);
nor U6420 (N_6420,N_5513,N_5919);
xnor U6421 (N_6421,N_5641,N_5720);
and U6422 (N_6422,N_5923,N_5821);
nor U6423 (N_6423,N_5662,N_5763);
xor U6424 (N_6424,N_5859,N_5966);
nand U6425 (N_6425,N_5723,N_5506);
or U6426 (N_6426,N_5663,N_5960);
or U6427 (N_6427,N_5529,N_5711);
and U6428 (N_6428,N_5911,N_5974);
nand U6429 (N_6429,N_5530,N_5738);
and U6430 (N_6430,N_5774,N_5988);
and U6431 (N_6431,N_5891,N_5824);
xnor U6432 (N_6432,N_5985,N_5922);
nor U6433 (N_6433,N_5557,N_5841);
xor U6434 (N_6434,N_5906,N_5945);
or U6435 (N_6435,N_5802,N_5604);
xnor U6436 (N_6436,N_5540,N_5691);
and U6437 (N_6437,N_5975,N_5640);
xor U6438 (N_6438,N_5884,N_5946);
and U6439 (N_6439,N_5550,N_5820);
nand U6440 (N_6440,N_5982,N_5550);
xnor U6441 (N_6441,N_5870,N_5507);
or U6442 (N_6442,N_5549,N_5855);
nor U6443 (N_6443,N_5881,N_5583);
nor U6444 (N_6444,N_5525,N_5604);
nor U6445 (N_6445,N_5805,N_5817);
xor U6446 (N_6446,N_5910,N_5692);
or U6447 (N_6447,N_5578,N_5682);
or U6448 (N_6448,N_5900,N_5993);
and U6449 (N_6449,N_5863,N_5930);
or U6450 (N_6450,N_5909,N_5700);
and U6451 (N_6451,N_5516,N_5755);
or U6452 (N_6452,N_5974,N_5669);
or U6453 (N_6453,N_5542,N_5930);
nor U6454 (N_6454,N_5929,N_5871);
xor U6455 (N_6455,N_5997,N_5698);
and U6456 (N_6456,N_5685,N_5956);
or U6457 (N_6457,N_5593,N_5715);
xnor U6458 (N_6458,N_5573,N_5803);
nand U6459 (N_6459,N_5780,N_5760);
xnor U6460 (N_6460,N_5560,N_5909);
xor U6461 (N_6461,N_5788,N_5949);
nor U6462 (N_6462,N_5611,N_5820);
nor U6463 (N_6463,N_5823,N_5724);
nand U6464 (N_6464,N_5696,N_5927);
and U6465 (N_6465,N_5847,N_5588);
or U6466 (N_6466,N_5798,N_5708);
xnor U6467 (N_6467,N_5733,N_5917);
nor U6468 (N_6468,N_5629,N_5940);
nand U6469 (N_6469,N_5946,N_5682);
nand U6470 (N_6470,N_5866,N_5968);
and U6471 (N_6471,N_5720,N_5871);
nor U6472 (N_6472,N_5919,N_5681);
or U6473 (N_6473,N_5855,N_5774);
nor U6474 (N_6474,N_5841,N_5750);
xnor U6475 (N_6475,N_5901,N_5705);
xnor U6476 (N_6476,N_5552,N_5575);
nand U6477 (N_6477,N_5718,N_5695);
or U6478 (N_6478,N_5662,N_5796);
xnor U6479 (N_6479,N_5830,N_5556);
and U6480 (N_6480,N_5789,N_5943);
xnor U6481 (N_6481,N_5636,N_5792);
xnor U6482 (N_6482,N_5955,N_5901);
nor U6483 (N_6483,N_5815,N_5899);
and U6484 (N_6484,N_5618,N_5619);
and U6485 (N_6485,N_5923,N_5834);
nor U6486 (N_6486,N_5681,N_5518);
or U6487 (N_6487,N_5928,N_5943);
or U6488 (N_6488,N_5632,N_5784);
or U6489 (N_6489,N_5686,N_5890);
xor U6490 (N_6490,N_5803,N_5774);
or U6491 (N_6491,N_5808,N_5905);
or U6492 (N_6492,N_5849,N_5770);
and U6493 (N_6493,N_5583,N_5666);
and U6494 (N_6494,N_5773,N_5785);
and U6495 (N_6495,N_5938,N_5597);
xnor U6496 (N_6496,N_5707,N_5539);
nor U6497 (N_6497,N_5770,N_5632);
xnor U6498 (N_6498,N_5939,N_5689);
nand U6499 (N_6499,N_5974,N_5582);
or U6500 (N_6500,N_6462,N_6351);
and U6501 (N_6501,N_6398,N_6267);
or U6502 (N_6502,N_6404,N_6205);
nor U6503 (N_6503,N_6246,N_6052);
nand U6504 (N_6504,N_6341,N_6131);
and U6505 (N_6505,N_6279,N_6356);
nor U6506 (N_6506,N_6295,N_6028);
xor U6507 (N_6507,N_6250,N_6484);
nand U6508 (N_6508,N_6416,N_6474);
or U6509 (N_6509,N_6387,N_6082);
or U6510 (N_6510,N_6411,N_6059);
xor U6511 (N_6511,N_6227,N_6033);
nand U6512 (N_6512,N_6147,N_6034);
nor U6513 (N_6513,N_6044,N_6296);
and U6514 (N_6514,N_6190,N_6446);
xor U6515 (N_6515,N_6208,N_6090);
nand U6516 (N_6516,N_6083,N_6156);
and U6517 (N_6517,N_6013,N_6247);
nor U6518 (N_6518,N_6268,N_6198);
nand U6519 (N_6519,N_6266,N_6107);
and U6520 (N_6520,N_6130,N_6135);
or U6521 (N_6521,N_6277,N_6382);
nand U6522 (N_6522,N_6001,N_6333);
and U6523 (N_6523,N_6461,N_6392);
or U6524 (N_6524,N_6389,N_6449);
and U6525 (N_6525,N_6138,N_6240);
nor U6526 (N_6526,N_6016,N_6496);
xnor U6527 (N_6527,N_6290,N_6085);
or U6528 (N_6528,N_6451,N_6039);
xnor U6529 (N_6529,N_6467,N_6414);
and U6530 (N_6530,N_6081,N_6282);
xor U6531 (N_6531,N_6364,N_6415);
or U6532 (N_6532,N_6353,N_6079);
and U6533 (N_6533,N_6084,N_6217);
nor U6534 (N_6534,N_6045,N_6197);
and U6535 (N_6535,N_6062,N_6212);
nor U6536 (N_6536,N_6106,N_6287);
nand U6537 (N_6537,N_6284,N_6271);
or U6538 (N_6538,N_6168,N_6298);
or U6539 (N_6539,N_6313,N_6174);
nor U6540 (N_6540,N_6248,N_6146);
and U6541 (N_6541,N_6409,N_6068);
or U6542 (N_6542,N_6256,N_6063);
nand U6543 (N_6543,N_6098,N_6096);
nand U6544 (N_6544,N_6380,N_6302);
xor U6545 (N_6545,N_6216,N_6148);
nor U6546 (N_6546,N_6127,N_6143);
xor U6547 (N_6547,N_6358,N_6487);
nand U6548 (N_6548,N_6196,N_6021);
nand U6549 (N_6549,N_6308,N_6064);
or U6550 (N_6550,N_6038,N_6325);
nand U6551 (N_6551,N_6157,N_6188);
xnor U6552 (N_6552,N_6065,N_6365);
xnor U6553 (N_6553,N_6465,N_6225);
xor U6554 (N_6554,N_6383,N_6219);
nand U6555 (N_6555,N_6192,N_6043);
or U6556 (N_6556,N_6057,N_6281);
nor U6557 (N_6557,N_6195,N_6306);
nor U6558 (N_6558,N_6099,N_6032);
xnor U6559 (N_6559,N_6428,N_6122);
or U6560 (N_6560,N_6361,N_6498);
or U6561 (N_6561,N_6150,N_6490);
nor U6562 (N_6562,N_6373,N_6105);
xnor U6563 (N_6563,N_6421,N_6483);
nand U6564 (N_6564,N_6340,N_6441);
nand U6565 (N_6565,N_6152,N_6088);
nor U6566 (N_6566,N_6024,N_6432);
or U6567 (N_6567,N_6104,N_6259);
or U6568 (N_6568,N_6211,N_6257);
or U6569 (N_6569,N_6445,N_6407);
nand U6570 (N_6570,N_6425,N_6172);
xnor U6571 (N_6571,N_6352,N_6234);
nor U6572 (N_6572,N_6301,N_6347);
and U6573 (N_6573,N_6471,N_6426);
xor U6574 (N_6574,N_6453,N_6381);
nand U6575 (N_6575,N_6184,N_6324);
or U6576 (N_6576,N_6419,N_6374);
nor U6577 (N_6577,N_6137,N_6086);
and U6578 (N_6578,N_6242,N_6417);
xor U6579 (N_6579,N_6393,N_6454);
and U6580 (N_6580,N_6254,N_6288);
or U6581 (N_6581,N_6022,N_6476);
nand U6582 (N_6582,N_6331,N_6166);
and U6583 (N_6583,N_6236,N_6493);
xor U6584 (N_6584,N_6424,N_6376);
xor U6585 (N_6585,N_6220,N_6486);
xor U6586 (N_6586,N_6073,N_6226);
nor U6587 (N_6587,N_6488,N_6164);
xnor U6588 (N_6588,N_6204,N_6093);
nor U6589 (N_6589,N_6434,N_6109);
or U6590 (N_6590,N_6307,N_6078);
nand U6591 (N_6591,N_6468,N_6323);
xor U6592 (N_6592,N_6187,N_6355);
or U6593 (N_6593,N_6263,N_6115);
or U6594 (N_6594,N_6452,N_6158);
xor U6595 (N_6595,N_6470,N_6144);
nor U6596 (N_6596,N_6249,N_6186);
and U6597 (N_6597,N_6151,N_6004);
xor U6598 (N_6598,N_6489,N_6299);
xor U6599 (N_6599,N_6218,N_6485);
nand U6600 (N_6600,N_6280,N_6019);
xnor U6601 (N_6601,N_6473,N_6260);
or U6602 (N_6602,N_6423,N_6049);
xnor U6603 (N_6603,N_6179,N_6456);
nor U6604 (N_6604,N_6114,N_6349);
and U6605 (N_6605,N_6206,N_6436);
nand U6606 (N_6606,N_6342,N_6007);
nand U6607 (N_6607,N_6481,N_6371);
nor U6608 (N_6608,N_6275,N_6181);
nor U6609 (N_6609,N_6286,N_6011);
and U6610 (N_6610,N_6031,N_6309);
and U6611 (N_6611,N_6350,N_6053);
xnor U6612 (N_6612,N_6326,N_6047);
xor U6613 (N_6613,N_6119,N_6455);
nor U6614 (N_6614,N_6403,N_6274);
and U6615 (N_6615,N_6343,N_6029);
and U6616 (N_6616,N_6182,N_6113);
or U6617 (N_6617,N_6189,N_6291);
and U6618 (N_6618,N_6080,N_6317);
nand U6619 (N_6619,N_6050,N_6066);
or U6620 (N_6620,N_6023,N_6163);
nor U6621 (N_6621,N_6366,N_6067);
and U6622 (N_6622,N_6191,N_6231);
nor U6623 (N_6623,N_6310,N_6435);
nand U6624 (N_6624,N_6167,N_6477);
xnor U6625 (N_6625,N_6431,N_6162);
nor U6626 (N_6626,N_6338,N_6040);
or U6627 (N_6627,N_6345,N_6141);
nand U6628 (N_6628,N_6292,N_6395);
xor U6629 (N_6629,N_6475,N_6178);
and U6630 (N_6630,N_6076,N_6170);
nand U6631 (N_6631,N_6367,N_6129);
and U6632 (N_6632,N_6095,N_6273);
or U6633 (N_6633,N_6289,N_6092);
xor U6634 (N_6634,N_6229,N_6177);
nand U6635 (N_6635,N_6153,N_6041);
nand U6636 (N_6636,N_6140,N_6030);
nand U6637 (N_6637,N_6450,N_6069);
or U6638 (N_6638,N_6311,N_6399);
and U6639 (N_6639,N_6003,N_6457);
nor U6640 (N_6640,N_6386,N_6091);
nand U6641 (N_6641,N_6094,N_6264);
or U6642 (N_6642,N_6017,N_6169);
or U6643 (N_6643,N_6401,N_6125);
xnor U6644 (N_6644,N_6000,N_6370);
xor U6645 (N_6645,N_6334,N_6132);
or U6646 (N_6646,N_6482,N_6075);
or U6647 (N_6647,N_6133,N_6176);
nor U6648 (N_6648,N_6448,N_6012);
or U6649 (N_6649,N_6036,N_6402);
nor U6650 (N_6650,N_6100,N_6117);
and U6651 (N_6651,N_6270,N_6077);
nor U6652 (N_6652,N_6276,N_6293);
or U6653 (N_6653,N_6244,N_6269);
nor U6654 (N_6654,N_6232,N_6479);
nand U6655 (N_6655,N_6165,N_6430);
and U6656 (N_6656,N_6362,N_6026);
nor U6657 (N_6657,N_6251,N_6139);
nand U6658 (N_6658,N_6018,N_6228);
or U6659 (N_6659,N_6201,N_6327);
nand U6660 (N_6660,N_6438,N_6002);
nand U6661 (N_6661,N_6285,N_6253);
and U6662 (N_6662,N_6121,N_6110);
nand U6663 (N_6663,N_6390,N_6058);
or U6664 (N_6664,N_6222,N_6009);
xnor U6665 (N_6665,N_6388,N_6329);
nor U6666 (N_6666,N_6061,N_6173);
nor U6667 (N_6667,N_6339,N_6429);
and U6668 (N_6668,N_6112,N_6346);
or U6669 (N_6669,N_6006,N_6161);
xnor U6670 (N_6670,N_6027,N_6305);
and U6671 (N_6671,N_6149,N_6159);
xnor U6672 (N_6672,N_6480,N_6335);
nand U6673 (N_6673,N_6116,N_6303);
nor U6674 (N_6674,N_6214,N_6258);
and U6675 (N_6675,N_6202,N_6363);
and U6676 (N_6676,N_6294,N_6048);
nor U6677 (N_6677,N_6348,N_6444);
xor U6678 (N_6678,N_6321,N_6055);
or U6679 (N_6679,N_6304,N_6492);
and U6680 (N_6680,N_6262,N_6375);
and U6681 (N_6681,N_6283,N_6315);
nor U6682 (N_6682,N_6224,N_6418);
xor U6683 (N_6683,N_6359,N_6037);
nor U6684 (N_6684,N_6297,N_6108);
or U6685 (N_6685,N_6193,N_6255);
nor U6686 (N_6686,N_6175,N_6272);
nor U6687 (N_6687,N_6210,N_6491);
xnor U6688 (N_6688,N_6396,N_6200);
nor U6689 (N_6689,N_6447,N_6203);
xor U6690 (N_6690,N_6463,N_6070);
xor U6691 (N_6691,N_6494,N_6397);
nand U6692 (N_6692,N_6378,N_6042);
nor U6693 (N_6693,N_6221,N_6103);
nor U6694 (N_6694,N_6372,N_6469);
and U6695 (N_6695,N_6472,N_6408);
and U6696 (N_6696,N_6405,N_6239);
and U6697 (N_6697,N_6120,N_6459);
xnor U6698 (N_6698,N_6422,N_6025);
nand U6699 (N_6699,N_6391,N_6213);
nand U6700 (N_6700,N_6142,N_6406);
nand U6701 (N_6701,N_6035,N_6278);
nand U6702 (N_6702,N_6233,N_6209);
and U6703 (N_6703,N_6154,N_6183);
nand U6704 (N_6704,N_6433,N_6199);
nand U6705 (N_6705,N_6466,N_6368);
and U6706 (N_6706,N_6437,N_6439);
or U6707 (N_6707,N_6443,N_6413);
or U6708 (N_6708,N_6336,N_6235);
nor U6709 (N_6709,N_6360,N_6410);
nand U6710 (N_6710,N_6440,N_6160);
nand U6711 (N_6711,N_6322,N_6060);
and U6712 (N_6712,N_6412,N_6332);
and U6713 (N_6713,N_6015,N_6230);
nor U6714 (N_6714,N_6427,N_6111);
nor U6715 (N_6715,N_6010,N_6499);
nor U6716 (N_6716,N_6330,N_6237);
or U6717 (N_6717,N_6155,N_6128);
nor U6718 (N_6718,N_6379,N_6369);
or U6719 (N_6719,N_6126,N_6243);
or U6720 (N_6720,N_6420,N_6344);
and U6721 (N_6721,N_6136,N_6008);
xor U6722 (N_6722,N_6497,N_6354);
and U6723 (N_6723,N_6337,N_6185);
nand U6724 (N_6724,N_6072,N_6241);
xor U6725 (N_6725,N_6377,N_6056);
and U6726 (N_6726,N_6238,N_6495);
nand U6727 (N_6727,N_6458,N_6215);
and U6728 (N_6728,N_6384,N_6261);
nand U6729 (N_6729,N_6020,N_6314);
and U6730 (N_6730,N_6087,N_6385);
nor U6731 (N_6731,N_6312,N_6318);
nand U6732 (N_6732,N_6097,N_6265);
or U6733 (N_6733,N_6394,N_6171);
xor U6734 (N_6734,N_6118,N_6319);
xnor U6735 (N_6735,N_6328,N_6180);
nor U6736 (N_6736,N_6194,N_6320);
or U6737 (N_6737,N_6014,N_6046);
or U6738 (N_6738,N_6207,N_6460);
nor U6739 (N_6739,N_6005,N_6223);
xnor U6740 (N_6740,N_6300,N_6123);
nor U6741 (N_6741,N_6074,N_6357);
xor U6742 (N_6742,N_6478,N_6102);
xor U6743 (N_6743,N_6071,N_6400);
xor U6744 (N_6744,N_6145,N_6316);
or U6745 (N_6745,N_6134,N_6054);
and U6746 (N_6746,N_6101,N_6051);
or U6747 (N_6747,N_6252,N_6464);
nor U6748 (N_6748,N_6245,N_6124);
xnor U6749 (N_6749,N_6442,N_6089);
and U6750 (N_6750,N_6467,N_6492);
nor U6751 (N_6751,N_6482,N_6379);
nand U6752 (N_6752,N_6019,N_6028);
or U6753 (N_6753,N_6051,N_6169);
nor U6754 (N_6754,N_6499,N_6346);
xor U6755 (N_6755,N_6011,N_6203);
nor U6756 (N_6756,N_6224,N_6153);
or U6757 (N_6757,N_6163,N_6168);
nor U6758 (N_6758,N_6484,N_6210);
nor U6759 (N_6759,N_6142,N_6171);
nor U6760 (N_6760,N_6051,N_6279);
xnor U6761 (N_6761,N_6488,N_6207);
and U6762 (N_6762,N_6459,N_6350);
xnor U6763 (N_6763,N_6199,N_6499);
and U6764 (N_6764,N_6363,N_6133);
or U6765 (N_6765,N_6102,N_6354);
or U6766 (N_6766,N_6320,N_6356);
xnor U6767 (N_6767,N_6344,N_6068);
or U6768 (N_6768,N_6425,N_6326);
xor U6769 (N_6769,N_6143,N_6133);
nand U6770 (N_6770,N_6456,N_6310);
nand U6771 (N_6771,N_6093,N_6313);
nand U6772 (N_6772,N_6058,N_6150);
and U6773 (N_6773,N_6480,N_6384);
nand U6774 (N_6774,N_6470,N_6026);
and U6775 (N_6775,N_6022,N_6141);
nor U6776 (N_6776,N_6392,N_6293);
xor U6777 (N_6777,N_6154,N_6246);
nor U6778 (N_6778,N_6205,N_6224);
nand U6779 (N_6779,N_6357,N_6058);
xnor U6780 (N_6780,N_6106,N_6110);
nor U6781 (N_6781,N_6354,N_6088);
nand U6782 (N_6782,N_6186,N_6051);
and U6783 (N_6783,N_6138,N_6356);
nand U6784 (N_6784,N_6277,N_6276);
nand U6785 (N_6785,N_6001,N_6386);
xor U6786 (N_6786,N_6291,N_6078);
nor U6787 (N_6787,N_6489,N_6311);
and U6788 (N_6788,N_6471,N_6445);
xor U6789 (N_6789,N_6354,N_6122);
and U6790 (N_6790,N_6008,N_6360);
and U6791 (N_6791,N_6108,N_6371);
or U6792 (N_6792,N_6084,N_6403);
nor U6793 (N_6793,N_6180,N_6269);
and U6794 (N_6794,N_6340,N_6390);
or U6795 (N_6795,N_6176,N_6460);
nand U6796 (N_6796,N_6319,N_6015);
and U6797 (N_6797,N_6078,N_6026);
nand U6798 (N_6798,N_6089,N_6031);
xor U6799 (N_6799,N_6227,N_6056);
and U6800 (N_6800,N_6083,N_6373);
xor U6801 (N_6801,N_6047,N_6445);
nor U6802 (N_6802,N_6410,N_6274);
nand U6803 (N_6803,N_6276,N_6184);
or U6804 (N_6804,N_6327,N_6479);
xnor U6805 (N_6805,N_6389,N_6347);
xnor U6806 (N_6806,N_6173,N_6214);
and U6807 (N_6807,N_6035,N_6157);
nor U6808 (N_6808,N_6387,N_6088);
xnor U6809 (N_6809,N_6011,N_6484);
and U6810 (N_6810,N_6337,N_6455);
and U6811 (N_6811,N_6449,N_6109);
nor U6812 (N_6812,N_6115,N_6299);
nor U6813 (N_6813,N_6243,N_6305);
nor U6814 (N_6814,N_6429,N_6017);
xnor U6815 (N_6815,N_6128,N_6274);
or U6816 (N_6816,N_6037,N_6449);
and U6817 (N_6817,N_6396,N_6320);
nand U6818 (N_6818,N_6413,N_6288);
nor U6819 (N_6819,N_6071,N_6346);
xor U6820 (N_6820,N_6172,N_6340);
xor U6821 (N_6821,N_6228,N_6448);
and U6822 (N_6822,N_6041,N_6005);
nor U6823 (N_6823,N_6068,N_6185);
nor U6824 (N_6824,N_6457,N_6337);
nand U6825 (N_6825,N_6108,N_6274);
or U6826 (N_6826,N_6104,N_6364);
nand U6827 (N_6827,N_6192,N_6131);
or U6828 (N_6828,N_6310,N_6306);
xnor U6829 (N_6829,N_6308,N_6485);
or U6830 (N_6830,N_6201,N_6232);
and U6831 (N_6831,N_6426,N_6351);
or U6832 (N_6832,N_6457,N_6069);
nand U6833 (N_6833,N_6447,N_6163);
nor U6834 (N_6834,N_6149,N_6021);
and U6835 (N_6835,N_6224,N_6201);
nor U6836 (N_6836,N_6222,N_6347);
nand U6837 (N_6837,N_6015,N_6376);
or U6838 (N_6838,N_6294,N_6034);
and U6839 (N_6839,N_6046,N_6035);
and U6840 (N_6840,N_6021,N_6163);
xnor U6841 (N_6841,N_6259,N_6049);
or U6842 (N_6842,N_6188,N_6104);
nor U6843 (N_6843,N_6281,N_6285);
or U6844 (N_6844,N_6149,N_6101);
nand U6845 (N_6845,N_6283,N_6001);
xnor U6846 (N_6846,N_6182,N_6150);
nor U6847 (N_6847,N_6365,N_6226);
or U6848 (N_6848,N_6191,N_6103);
xor U6849 (N_6849,N_6228,N_6411);
nor U6850 (N_6850,N_6063,N_6002);
nand U6851 (N_6851,N_6084,N_6369);
or U6852 (N_6852,N_6416,N_6188);
nand U6853 (N_6853,N_6379,N_6357);
nor U6854 (N_6854,N_6477,N_6390);
nor U6855 (N_6855,N_6491,N_6149);
nand U6856 (N_6856,N_6380,N_6421);
and U6857 (N_6857,N_6296,N_6242);
and U6858 (N_6858,N_6113,N_6306);
and U6859 (N_6859,N_6330,N_6177);
or U6860 (N_6860,N_6345,N_6464);
and U6861 (N_6861,N_6242,N_6243);
xor U6862 (N_6862,N_6413,N_6437);
xnor U6863 (N_6863,N_6366,N_6436);
nand U6864 (N_6864,N_6424,N_6056);
nor U6865 (N_6865,N_6483,N_6188);
and U6866 (N_6866,N_6312,N_6410);
or U6867 (N_6867,N_6358,N_6281);
nand U6868 (N_6868,N_6319,N_6398);
xor U6869 (N_6869,N_6362,N_6377);
or U6870 (N_6870,N_6256,N_6008);
nand U6871 (N_6871,N_6359,N_6405);
nand U6872 (N_6872,N_6425,N_6448);
or U6873 (N_6873,N_6193,N_6171);
nor U6874 (N_6874,N_6206,N_6366);
and U6875 (N_6875,N_6404,N_6491);
xnor U6876 (N_6876,N_6308,N_6046);
or U6877 (N_6877,N_6068,N_6247);
xor U6878 (N_6878,N_6203,N_6130);
nand U6879 (N_6879,N_6468,N_6145);
nand U6880 (N_6880,N_6392,N_6228);
and U6881 (N_6881,N_6306,N_6218);
and U6882 (N_6882,N_6328,N_6193);
or U6883 (N_6883,N_6499,N_6384);
xor U6884 (N_6884,N_6146,N_6203);
nand U6885 (N_6885,N_6490,N_6454);
nor U6886 (N_6886,N_6049,N_6112);
nand U6887 (N_6887,N_6257,N_6131);
or U6888 (N_6888,N_6160,N_6067);
nand U6889 (N_6889,N_6305,N_6092);
or U6890 (N_6890,N_6045,N_6490);
and U6891 (N_6891,N_6033,N_6167);
xnor U6892 (N_6892,N_6249,N_6288);
nand U6893 (N_6893,N_6034,N_6229);
xor U6894 (N_6894,N_6453,N_6380);
or U6895 (N_6895,N_6366,N_6154);
nand U6896 (N_6896,N_6370,N_6460);
nor U6897 (N_6897,N_6277,N_6156);
and U6898 (N_6898,N_6101,N_6408);
xnor U6899 (N_6899,N_6043,N_6002);
nor U6900 (N_6900,N_6422,N_6188);
nand U6901 (N_6901,N_6140,N_6258);
nand U6902 (N_6902,N_6428,N_6192);
nor U6903 (N_6903,N_6132,N_6262);
or U6904 (N_6904,N_6273,N_6363);
and U6905 (N_6905,N_6062,N_6348);
and U6906 (N_6906,N_6321,N_6272);
nor U6907 (N_6907,N_6147,N_6008);
nand U6908 (N_6908,N_6017,N_6189);
and U6909 (N_6909,N_6036,N_6419);
and U6910 (N_6910,N_6072,N_6208);
or U6911 (N_6911,N_6494,N_6280);
nand U6912 (N_6912,N_6474,N_6386);
or U6913 (N_6913,N_6215,N_6116);
nand U6914 (N_6914,N_6182,N_6340);
xor U6915 (N_6915,N_6449,N_6221);
xor U6916 (N_6916,N_6389,N_6043);
nand U6917 (N_6917,N_6068,N_6434);
and U6918 (N_6918,N_6480,N_6126);
nand U6919 (N_6919,N_6339,N_6351);
and U6920 (N_6920,N_6264,N_6432);
or U6921 (N_6921,N_6282,N_6442);
and U6922 (N_6922,N_6205,N_6251);
or U6923 (N_6923,N_6073,N_6198);
and U6924 (N_6924,N_6363,N_6498);
nand U6925 (N_6925,N_6120,N_6289);
nand U6926 (N_6926,N_6299,N_6331);
and U6927 (N_6927,N_6396,N_6434);
nor U6928 (N_6928,N_6445,N_6367);
nor U6929 (N_6929,N_6423,N_6055);
nor U6930 (N_6930,N_6216,N_6417);
nand U6931 (N_6931,N_6226,N_6148);
nor U6932 (N_6932,N_6377,N_6038);
or U6933 (N_6933,N_6107,N_6410);
nand U6934 (N_6934,N_6383,N_6067);
and U6935 (N_6935,N_6347,N_6299);
xnor U6936 (N_6936,N_6307,N_6350);
nor U6937 (N_6937,N_6307,N_6449);
nor U6938 (N_6938,N_6237,N_6053);
nor U6939 (N_6939,N_6083,N_6205);
nor U6940 (N_6940,N_6392,N_6407);
and U6941 (N_6941,N_6453,N_6418);
or U6942 (N_6942,N_6003,N_6382);
nor U6943 (N_6943,N_6358,N_6158);
and U6944 (N_6944,N_6078,N_6212);
and U6945 (N_6945,N_6187,N_6292);
nand U6946 (N_6946,N_6286,N_6066);
nor U6947 (N_6947,N_6429,N_6221);
and U6948 (N_6948,N_6175,N_6408);
xor U6949 (N_6949,N_6134,N_6461);
and U6950 (N_6950,N_6329,N_6392);
or U6951 (N_6951,N_6219,N_6192);
nor U6952 (N_6952,N_6415,N_6287);
nand U6953 (N_6953,N_6478,N_6057);
nor U6954 (N_6954,N_6425,N_6294);
xnor U6955 (N_6955,N_6399,N_6374);
nand U6956 (N_6956,N_6070,N_6370);
and U6957 (N_6957,N_6190,N_6257);
nand U6958 (N_6958,N_6220,N_6218);
and U6959 (N_6959,N_6090,N_6247);
and U6960 (N_6960,N_6181,N_6140);
and U6961 (N_6961,N_6218,N_6152);
and U6962 (N_6962,N_6222,N_6130);
nand U6963 (N_6963,N_6071,N_6227);
xnor U6964 (N_6964,N_6261,N_6117);
nand U6965 (N_6965,N_6366,N_6170);
nor U6966 (N_6966,N_6166,N_6104);
nor U6967 (N_6967,N_6236,N_6391);
xnor U6968 (N_6968,N_6330,N_6328);
nor U6969 (N_6969,N_6066,N_6387);
and U6970 (N_6970,N_6243,N_6116);
nor U6971 (N_6971,N_6087,N_6056);
and U6972 (N_6972,N_6476,N_6030);
nor U6973 (N_6973,N_6401,N_6331);
or U6974 (N_6974,N_6384,N_6344);
or U6975 (N_6975,N_6068,N_6472);
nand U6976 (N_6976,N_6147,N_6491);
and U6977 (N_6977,N_6381,N_6286);
and U6978 (N_6978,N_6092,N_6450);
or U6979 (N_6979,N_6374,N_6417);
or U6980 (N_6980,N_6113,N_6021);
and U6981 (N_6981,N_6038,N_6167);
nor U6982 (N_6982,N_6040,N_6415);
nor U6983 (N_6983,N_6155,N_6318);
nor U6984 (N_6984,N_6056,N_6216);
nand U6985 (N_6985,N_6332,N_6113);
nor U6986 (N_6986,N_6470,N_6136);
and U6987 (N_6987,N_6053,N_6343);
xnor U6988 (N_6988,N_6279,N_6317);
nand U6989 (N_6989,N_6117,N_6200);
or U6990 (N_6990,N_6140,N_6108);
xnor U6991 (N_6991,N_6420,N_6436);
nor U6992 (N_6992,N_6086,N_6095);
nand U6993 (N_6993,N_6218,N_6040);
xor U6994 (N_6994,N_6445,N_6038);
nand U6995 (N_6995,N_6331,N_6473);
or U6996 (N_6996,N_6304,N_6331);
or U6997 (N_6997,N_6358,N_6284);
nor U6998 (N_6998,N_6038,N_6495);
or U6999 (N_6999,N_6465,N_6398);
xnor U7000 (N_7000,N_6679,N_6515);
nor U7001 (N_7001,N_6902,N_6773);
and U7002 (N_7002,N_6960,N_6741);
nand U7003 (N_7003,N_6596,N_6635);
xor U7004 (N_7004,N_6796,N_6705);
and U7005 (N_7005,N_6771,N_6573);
or U7006 (N_7006,N_6787,N_6988);
nor U7007 (N_7007,N_6670,N_6912);
nand U7008 (N_7008,N_6744,N_6614);
xor U7009 (N_7009,N_6520,N_6671);
nand U7010 (N_7010,N_6860,N_6973);
or U7011 (N_7011,N_6729,N_6948);
xnor U7012 (N_7012,N_6502,N_6828);
and U7013 (N_7013,N_6687,N_6721);
xor U7014 (N_7014,N_6666,N_6688);
nor U7015 (N_7015,N_6602,N_6969);
nor U7016 (N_7016,N_6563,N_6930);
or U7017 (N_7017,N_6881,N_6662);
and U7018 (N_7018,N_6816,N_6581);
nor U7019 (N_7019,N_6768,N_6663);
nor U7020 (N_7020,N_6636,N_6511);
or U7021 (N_7021,N_6939,N_6975);
and U7022 (N_7022,N_6879,N_6629);
or U7023 (N_7023,N_6922,N_6704);
and U7024 (N_7024,N_6594,N_6691);
nand U7025 (N_7025,N_6780,N_6616);
and U7026 (N_7026,N_6605,N_6595);
nand U7027 (N_7027,N_6880,N_6833);
nand U7028 (N_7028,N_6901,N_6858);
xnor U7029 (N_7029,N_6947,N_6755);
nor U7030 (N_7030,N_6999,N_6588);
or U7031 (N_7031,N_6774,N_6634);
nand U7032 (N_7032,N_6737,N_6720);
or U7033 (N_7033,N_6590,N_6844);
or U7034 (N_7034,N_6577,N_6536);
and U7035 (N_7035,N_6644,N_6785);
nor U7036 (N_7036,N_6713,N_6758);
nand U7037 (N_7037,N_6503,N_6598);
nor U7038 (N_7038,N_6946,N_6829);
and U7039 (N_7039,N_6501,N_6897);
and U7040 (N_7040,N_6990,N_6541);
nor U7041 (N_7041,N_6877,N_6994);
xor U7042 (N_7042,N_6798,N_6586);
or U7043 (N_7043,N_6809,N_6891);
and U7044 (N_7044,N_6748,N_6898);
xnor U7045 (N_7045,N_6706,N_6587);
nand U7046 (N_7046,N_6625,N_6921);
or U7047 (N_7047,N_6507,N_6963);
or U7048 (N_7048,N_6509,N_6795);
and U7049 (N_7049,N_6826,N_6915);
nand U7050 (N_7050,N_6832,N_6653);
and U7051 (N_7051,N_6801,N_6820);
or U7052 (N_7052,N_6791,N_6840);
nand U7053 (N_7053,N_6628,N_6556);
xor U7054 (N_7054,N_6583,N_6531);
and U7055 (N_7055,N_6980,N_6945);
nand U7056 (N_7056,N_6893,N_6845);
xnor U7057 (N_7057,N_6732,N_6923);
nor U7058 (N_7058,N_6876,N_6557);
and U7059 (N_7059,N_6643,N_6637);
nor U7060 (N_7060,N_6778,N_6950);
or U7061 (N_7061,N_6872,N_6895);
or U7062 (N_7062,N_6976,N_6807);
or U7063 (N_7063,N_6730,N_6609);
nor U7064 (N_7064,N_6918,N_6709);
xor U7065 (N_7065,N_6576,N_6538);
or U7066 (N_7066,N_6514,N_6522);
nand U7067 (N_7067,N_6917,N_6797);
and U7068 (N_7068,N_6674,N_6851);
nor U7069 (N_7069,N_6633,N_6677);
nor U7070 (N_7070,N_6943,N_6769);
nand U7071 (N_7071,N_6838,N_6567);
nor U7072 (N_7072,N_6937,N_6841);
nor U7073 (N_7073,N_6718,N_6523);
nor U7074 (N_7074,N_6570,N_6689);
or U7075 (N_7075,N_6660,N_6743);
or U7076 (N_7076,N_6823,N_6938);
and U7077 (N_7077,N_6537,N_6953);
and U7078 (N_7078,N_6804,N_6642);
nor U7079 (N_7079,N_6699,N_6597);
nor U7080 (N_7080,N_6665,N_6986);
nor U7081 (N_7081,N_6885,N_6626);
xnor U7082 (N_7082,N_6714,N_6600);
or U7083 (N_7083,N_6672,N_6961);
nor U7084 (N_7084,N_6776,N_6919);
nand U7085 (N_7085,N_6683,N_6924);
or U7086 (N_7086,N_6746,N_6690);
and U7087 (N_7087,N_6813,N_6708);
nand U7088 (N_7088,N_6914,N_6545);
and U7089 (N_7089,N_6886,N_6608);
or U7090 (N_7090,N_6955,N_6967);
and U7091 (N_7091,N_6562,N_6604);
nand U7092 (N_7092,N_6640,N_6516);
and U7093 (N_7093,N_6652,N_6848);
xor U7094 (N_7094,N_6763,N_6727);
or U7095 (N_7095,N_6676,N_6977);
nand U7096 (N_7096,N_6752,N_6834);
or U7097 (N_7097,N_6623,N_6649);
nand U7098 (N_7098,N_6906,N_6781);
or U7099 (N_7099,N_6942,N_6651);
and U7100 (N_7100,N_6717,N_6592);
or U7101 (N_7101,N_6874,N_6822);
and U7102 (N_7102,N_6610,N_6681);
nand U7103 (N_7103,N_6611,N_6749);
xnor U7104 (N_7104,N_6504,N_6772);
and U7105 (N_7105,N_6814,N_6508);
xor U7106 (N_7106,N_6530,N_6971);
nand U7107 (N_7107,N_6770,N_6534);
nor U7108 (N_7108,N_6951,N_6742);
xnor U7109 (N_7109,N_6571,N_6540);
xor U7110 (N_7110,N_6551,N_6944);
xnor U7111 (N_7111,N_6964,N_6928);
nor U7112 (N_7112,N_6892,N_6997);
and U7113 (N_7113,N_6751,N_6655);
nand U7114 (N_7114,N_6675,N_6542);
or U7115 (N_7115,N_6959,N_6533);
xnor U7116 (N_7116,N_6871,N_6680);
and U7117 (N_7117,N_6788,N_6631);
nor U7118 (N_7118,N_6574,N_6527);
xor U7119 (N_7119,N_6936,N_6510);
nor U7120 (N_7120,N_6726,N_6849);
and U7121 (N_7121,N_6618,N_6517);
nor U7122 (N_7122,N_6529,N_6673);
nand U7123 (N_7123,N_6933,N_6831);
nand U7124 (N_7124,N_6852,N_6544);
nor U7125 (N_7125,N_6935,N_6965);
xnor U7126 (N_7126,N_6888,N_6966);
nand U7127 (N_7127,N_6722,N_6613);
nand U7128 (N_7128,N_6981,N_6684);
xor U7129 (N_7129,N_6782,N_6993);
or U7130 (N_7130,N_6932,N_6750);
nor U7131 (N_7131,N_6646,N_6696);
nand U7132 (N_7132,N_6558,N_6546);
and U7133 (N_7133,N_6926,N_6512);
and U7134 (N_7134,N_6745,N_6856);
nor U7135 (N_7135,N_6850,N_6870);
nand U7136 (N_7136,N_6925,N_6524);
or U7137 (N_7137,N_6621,N_6548);
xor U7138 (N_7138,N_6836,N_6547);
nand U7139 (N_7139,N_6799,N_6747);
nor U7140 (N_7140,N_6612,N_6995);
or U7141 (N_7141,N_6916,N_6606);
xnor U7142 (N_7142,N_6593,N_6783);
and U7143 (N_7143,N_6575,N_6572);
nand U7144 (N_7144,N_6827,N_6728);
xnor U7145 (N_7145,N_6695,N_6911);
nand U7146 (N_7146,N_6599,N_6528);
nor U7147 (N_7147,N_6878,N_6985);
and U7148 (N_7148,N_6927,N_6910);
nor U7149 (N_7149,N_6957,N_6884);
nand U7150 (N_7150,N_6535,N_6979);
or U7151 (N_7151,N_6686,N_6630);
xnor U7152 (N_7152,N_6875,N_6835);
xnor U7153 (N_7153,N_6920,N_6735);
and U7154 (N_7154,N_6553,N_6661);
xor U7155 (N_7155,N_6913,N_6733);
or U7156 (N_7156,N_6724,N_6810);
nand U7157 (N_7157,N_6700,N_6865);
xor U7158 (N_7158,N_6775,N_6707);
xor U7159 (N_7159,N_6759,N_6580);
nand U7160 (N_7160,N_6561,N_6521);
nor U7161 (N_7161,N_6989,N_6817);
xnor U7162 (N_7162,N_6615,N_6941);
nand U7163 (N_7163,N_6786,N_6903);
nor U7164 (N_7164,N_6837,N_6641);
and U7165 (N_7165,N_6624,N_6802);
xnor U7166 (N_7166,N_6703,N_6894);
nor U7167 (N_7167,N_6949,N_6899);
or U7168 (N_7168,N_6552,N_6821);
or U7169 (N_7169,N_6698,N_6754);
nand U7170 (N_7170,N_6736,N_6519);
nand U7171 (N_7171,N_6762,N_6929);
nor U7172 (N_7172,N_6702,N_6991);
or U7173 (N_7173,N_6582,N_6761);
or U7174 (N_7174,N_6591,N_6719);
and U7175 (N_7175,N_6697,N_6907);
or U7176 (N_7176,N_6792,N_6734);
nor U7177 (N_7177,N_6806,N_6617);
and U7178 (N_7178,N_6603,N_6882);
xor U7179 (N_7179,N_6819,N_6970);
xor U7180 (N_7180,N_6863,N_6701);
nor U7181 (N_7181,N_6659,N_6998);
and U7182 (N_7182,N_6668,N_6711);
or U7183 (N_7183,N_6765,N_6805);
nand U7184 (N_7184,N_6525,N_6532);
or U7185 (N_7185,N_6958,N_6650);
nand U7186 (N_7186,N_6984,N_6694);
nor U7187 (N_7187,N_6667,N_6723);
nand U7188 (N_7188,N_6585,N_6956);
nand U7189 (N_7189,N_6757,N_6794);
or U7190 (N_7190,N_6864,N_6908);
xnor U7191 (N_7191,N_6555,N_6506);
xor U7192 (N_7192,N_6518,N_6873);
or U7193 (N_7193,N_6554,N_6738);
xor U7194 (N_7194,N_6808,N_6900);
nand U7195 (N_7195,N_6658,N_6766);
nor U7196 (N_7196,N_6622,N_6992);
and U7197 (N_7197,N_6607,N_6818);
or U7198 (N_7198,N_6500,N_6861);
xnor U7199 (N_7199,N_6559,N_6867);
xor U7200 (N_7200,N_6620,N_6934);
xor U7201 (N_7201,N_6824,N_6657);
nor U7202 (N_7202,N_6756,N_6815);
and U7203 (N_7203,N_6568,N_6682);
and U7204 (N_7204,N_6692,N_6855);
and U7205 (N_7205,N_6853,N_6846);
nand U7206 (N_7206,N_6789,N_6560);
xor U7207 (N_7207,N_6645,N_6793);
or U7208 (N_7208,N_6656,N_6862);
nand U7209 (N_7209,N_6859,N_6725);
nand U7210 (N_7210,N_6678,N_6803);
and U7211 (N_7211,N_6790,N_6647);
nand U7212 (N_7212,N_6664,N_6952);
or U7213 (N_7213,N_6962,N_6526);
xnor U7214 (N_7214,N_6578,N_6983);
xnor U7215 (N_7215,N_6830,N_6539);
nor U7216 (N_7216,N_6764,N_6693);
nor U7217 (N_7217,N_6905,N_6619);
and U7218 (N_7218,N_6648,N_6669);
nand U7219 (N_7219,N_6839,N_6584);
and U7220 (N_7220,N_6825,N_6543);
or U7221 (N_7221,N_6731,N_6800);
xnor U7222 (N_7222,N_6996,N_6566);
xnor U7223 (N_7223,N_6889,N_6654);
nor U7224 (N_7224,N_6904,N_6896);
nor U7225 (N_7225,N_6638,N_6710);
or U7226 (N_7226,N_6847,N_6866);
nand U7227 (N_7227,N_6854,N_6974);
nand U7228 (N_7228,N_6940,N_6890);
or U7229 (N_7229,N_6968,N_6887);
nand U7230 (N_7230,N_6601,N_6812);
nand U7231 (N_7231,N_6740,N_6779);
and U7232 (N_7232,N_6857,N_6627);
nand U7233 (N_7233,N_6513,N_6978);
xnor U7234 (N_7234,N_6883,N_6550);
xnor U7235 (N_7235,N_6753,N_6767);
nor U7236 (N_7236,N_6564,N_6987);
xnor U7237 (N_7237,N_6972,N_6843);
or U7238 (N_7238,N_6868,N_6589);
xor U7239 (N_7239,N_6632,N_6982);
xnor U7240 (N_7240,N_6842,N_6565);
and U7241 (N_7241,N_6811,N_6760);
nor U7242 (N_7242,N_6739,N_6685);
and U7243 (N_7243,N_6715,N_6549);
or U7244 (N_7244,N_6716,N_6569);
or U7245 (N_7245,N_6712,N_6639);
and U7246 (N_7246,N_6784,N_6954);
and U7247 (N_7247,N_6869,N_6505);
xnor U7248 (N_7248,N_6909,N_6777);
nand U7249 (N_7249,N_6931,N_6579);
xnor U7250 (N_7250,N_6675,N_6551);
nor U7251 (N_7251,N_6933,N_6776);
nor U7252 (N_7252,N_6731,N_6842);
nand U7253 (N_7253,N_6580,N_6602);
or U7254 (N_7254,N_6717,N_6778);
nor U7255 (N_7255,N_6852,N_6905);
xor U7256 (N_7256,N_6734,N_6927);
nor U7257 (N_7257,N_6570,N_6519);
nand U7258 (N_7258,N_6841,N_6899);
xnor U7259 (N_7259,N_6781,N_6780);
nor U7260 (N_7260,N_6927,N_6685);
or U7261 (N_7261,N_6733,N_6668);
nand U7262 (N_7262,N_6717,N_6609);
xor U7263 (N_7263,N_6634,N_6884);
xor U7264 (N_7264,N_6686,N_6861);
xor U7265 (N_7265,N_6562,N_6590);
and U7266 (N_7266,N_6613,N_6646);
nand U7267 (N_7267,N_6500,N_6815);
nand U7268 (N_7268,N_6739,N_6920);
or U7269 (N_7269,N_6527,N_6909);
and U7270 (N_7270,N_6619,N_6742);
and U7271 (N_7271,N_6563,N_6722);
nor U7272 (N_7272,N_6774,N_6757);
nor U7273 (N_7273,N_6786,N_6956);
and U7274 (N_7274,N_6891,N_6572);
xnor U7275 (N_7275,N_6681,N_6851);
or U7276 (N_7276,N_6726,N_6672);
xor U7277 (N_7277,N_6549,N_6621);
nand U7278 (N_7278,N_6693,N_6683);
xor U7279 (N_7279,N_6863,N_6616);
nor U7280 (N_7280,N_6507,N_6846);
nand U7281 (N_7281,N_6631,N_6907);
xor U7282 (N_7282,N_6942,N_6809);
and U7283 (N_7283,N_6848,N_6680);
xnor U7284 (N_7284,N_6844,N_6856);
nor U7285 (N_7285,N_6996,N_6887);
xor U7286 (N_7286,N_6753,N_6778);
and U7287 (N_7287,N_6505,N_6969);
xor U7288 (N_7288,N_6733,N_6666);
nor U7289 (N_7289,N_6539,N_6613);
xnor U7290 (N_7290,N_6794,N_6668);
nor U7291 (N_7291,N_6866,N_6856);
or U7292 (N_7292,N_6937,N_6821);
nand U7293 (N_7293,N_6569,N_6941);
nand U7294 (N_7294,N_6970,N_6759);
or U7295 (N_7295,N_6862,N_6884);
or U7296 (N_7296,N_6547,N_6763);
nand U7297 (N_7297,N_6626,N_6631);
xor U7298 (N_7298,N_6642,N_6800);
nor U7299 (N_7299,N_6812,N_6663);
xnor U7300 (N_7300,N_6968,N_6899);
or U7301 (N_7301,N_6759,N_6528);
nand U7302 (N_7302,N_6995,N_6515);
or U7303 (N_7303,N_6773,N_6825);
nor U7304 (N_7304,N_6792,N_6757);
nor U7305 (N_7305,N_6546,N_6500);
nand U7306 (N_7306,N_6812,N_6721);
and U7307 (N_7307,N_6888,N_6622);
or U7308 (N_7308,N_6551,N_6669);
nor U7309 (N_7309,N_6567,N_6842);
xnor U7310 (N_7310,N_6906,N_6624);
or U7311 (N_7311,N_6932,N_6981);
and U7312 (N_7312,N_6513,N_6645);
nor U7313 (N_7313,N_6773,N_6842);
nand U7314 (N_7314,N_6737,N_6685);
and U7315 (N_7315,N_6685,N_6645);
xnor U7316 (N_7316,N_6887,N_6732);
nor U7317 (N_7317,N_6905,N_6715);
nand U7318 (N_7318,N_6858,N_6553);
nand U7319 (N_7319,N_6659,N_6797);
and U7320 (N_7320,N_6519,N_6562);
xnor U7321 (N_7321,N_6806,N_6653);
nand U7322 (N_7322,N_6563,N_6749);
xor U7323 (N_7323,N_6978,N_6636);
nand U7324 (N_7324,N_6535,N_6884);
xnor U7325 (N_7325,N_6839,N_6988);
nand U7326 (N_7326,N_6848,N_6737);
and U7327 (N_7327,N_6505,N_6788);
or U7328 (N_7328,N_6848,N_6937);
or U7329 (N_7329,N_6613,N_6623);
nand U7330 (N_7330,N_6552,N_6625);
nand U7331 (N_7331,N_6966,N_6760);
or U7332 (N_7332,N_6875,N_6707);
nand U7333 (N_7333,N_6626,N_6519);
nor U7334 (N_7334,N_6725,N_6587);
nor U7335 (N_7335,N_6754,N_6997);
and U7336 (N_7336,N_6647,N_6770);
nand U7337 (N_7337,N_6829,N_6766);
nor U7338 (N_7338,N_6582,N_6816);
xnor U7339 (N_7339,N_6901,N_6831);
nor U7340 (N_7340,N_6575,N_6895);
or U7341 (N_7341,N_6805,N_6801);
nand U7342 (N_7342,N_6668,N_6819);
and U7343 (N_7343,N_6934,N_6947);
or U7344 (N_7344,N_6738,N_6823);
nor U7345 (N_7345,N_6890,N_6993);
xor U7346 (N_7346,N_6849,N_6876);
or U7347 (N_7347,N_6734,N_6650);
and U7348 (N_7348,N_6798,N_6926);
xnor U7349 (N_7349,N_6755,N_6698);
nand U7350 (N_7350,N_6818,N_6522);
and U7351 (N_7351,N_6698,N_6769);
or U7352 (N_7352,N_6688,N_6864);
nand U7353 (N_7353,N_6593,N_6894);
and U7354 (N_7354,N_6873,N_6596);
or U7355 (N_7355,N_6811,N_6520);
xor U7356 (N_7356,N_6876,N_6642);
xor U7357 (N_7357,N_6758,N_6903);
xnor U7358 (N_7358,N_6577,N_6539);
nor U7359 (N_7359,N_6930,N_6972);
nor U7360 (N_7360,N_6973,N_6736);
nor U7361 (N_7361,N_6868,N_6824);
xor U7362 (N_7362,N_6616,N_6760);
or U7363 (N_7363,N_6660,N_6811);
xnor U7364 (N_7364,N_6961,N_6820);
xnor U7365 (N_7365,N_6857,N_6865);
xnor U7366 (N_7366,N_6973,N_6547);
xnor U7367 (N_7367,N_6674,N_6962);
nand U7368 (N_7368,N_6542,N_6898);
and U7369 (N_7369,N_6619,N_6769);
or U7370 (N_7370,N_6990,N_6859);
or U7371 (N_7371,N_6673,N_6774);
and U7372 (N_7372,N_6801,N_6534);
or U7373 (N_7373,N_6601,N_6619);
nand U7374 (N_7374,N_6875,N_6682);
and U7375 (N_7375,N_6922,N_6592);
nor U7376 (N_7376,N_6668,N_6692);
nor U7377 (N_7377,N_6995,N_6677);
or U7378 (N_7378,N_6868,N_6736);
xnor U7379 (N_7379,N_6567,N_6624);
or U7380 (N_7380,N_6803,N_6515);
xor U7381 (N_7381,N_6769,N_6692);
and U7382 (N_7382,N_6747,N_6574);
nand U7383 (N_7383,N_6777,N_6648);
or U7384 (N_7384,N_6764,N_6578);
xnor U7385 (N_7385,N_6917,N_6729);
and U7386 (N_7386,N_6936,N_6547);
or U7387 (N_7387,N_6856,N_6952);
nor U7388 (N_7388,N_6506,N_6976);
xnor U7389 (N_7389,N_6735,N_6669);
xor U7390 (N_7390,N_6787,N_6807);
xnor U7391 (N_7391,N_6821,N_6607);
or U7392 (N_7392,N_6640,N_6810);
nand U7393 (N_7393,N_6652,N_6880);
nor U7394 (N_7394,N_6555,N_6531);
or U7395 (N_7395,N_6808,N_6778);
or U7396 (N_7396,N_6827,N_6594);
and U7397 (N_7397,N_6773,N_6512);
nand U7398 (N_7398,N_6752,N_6527);
nor U7399 (N_7399,N_6940,N_6621);
xnor U7400 (N_7400,N_6894,N_6505);
and U7401 (N_7401,N_6550,N_6871);
nor U7402 (N_7402,N_6801,N_6861);
nand U7403 (N_7403,N_6595,N_6780);
nand U7404 (N_7404,N_6795,N_6674);
xnor U7405 (N_7405,N_6807,N_6815);
nand U7406 (N_7406,N_6771,N_6954);
nand U7407 (N_7407,N_6796,N_6730);
and U7408 (N_7408,N_6604,N_6912);
or U7409 (N_7409,N_6766,N_6668);
nand U7410 (N_7410,N_6880,N_6510);
xor U7411 (N_7411,N_6893,N_6715);
and U7412 (N_7412,N_6933,N_6940);
or U7413 (N_7413,N_6652,N_6655);
xor U7414 (N_7414,N_6927,N_6999);
nand U7415 (N_7415,N_6870,N_6940);
nor U7416 (N_7416,N_6743,N_6960);
nand U7417 (N_7417,N_6845,N_6732);
and U7418 (N_7418,N_6697,N_6723);
and U7419 (N_7419,N_6599,N_6652);
or U7420 (N_7420,N_6693,N_6933);
and U7421 (N_7421,N_6756,N_6856);
xnor U7422 (N_7422,N_6502,N_6767);
nor U7423 (N_7423,N_6846,N_6573);
nor U7424 (N_7424,N_6929,N_6535);
nor U7425 (N_7425,N_6526,N_6869);
nand U7426 (N_7426,N_6798,N_6820);
nor U7427 (N_7427,N_6604,N_6635);
or U7428 (N_7428,N_6925,N_6526);
xnor U7429 (N_7429,N_6779,N_6743);
nor U7430 (N_7430,N_6659,N_6862);
and U7431 (N_7431,N_6870,N_6650);
or U7432 (N_7432,N_6685,N_6883);
nand U7433 (N_7433,N_6986,N_6564);
and U7434 (N_7434,N_6685,N_6592);
nand U7435 (N_7435,N_6678,N_6587);
and U7436 (N_7436,N_6903,N_6930);
xor U7437 (N_7437,N_6840,N_6703);
xor U7438 (N_7438,N_6725,N_6701);
and U7439 (N_7439,N_6806,N_6557);
nor U7440 (N_7440,N_6773,N_6520);
xor U7441 (N_7441,N_6731,N_6942);
or U7442 (N_7442,N_6512,N_6757);
nor U7443 (N_7443,N_6903,N_6747);
or U7444 (N_7444,N_6592,N_6947);
xor U7445 (N_7445,N_6986,N_6949);
and U7446 (N_7446,N_6955,N_6929);
xnor U7447 (N_7447,N_6859,N_6549);
or U7448 (N_7448,N_6641,N_6899);
nand U7449 (N_7449,N_6953,N_6911);
xnor U7450 (N_7450,N_6802,N_6984);
xor U7451 (N_7451,N_6865,N_6856);
nand U7452 (N_7452,N_6860,N_6545);
nand U7453 (N_7453,N_6916,N_6580);
nand U7454 (N_7454,N_6907,N_6824);
or U7455 (N_7455,N_6907,N_6834);
or U7456 (N_7456,N_6974,N_6587);
and U7457 (N_7457,N_6903,N_6909);
and U7458 (N_7458,N_6843,N_6798);
or U7459 (N_7459,N_6791,N_6751);
and U7460 (N_7460,N_6597,N_6792);
nand U7461 (N_7461,N_6834,N_6823);
nor U7462 (N_7462,N_6992,N_6798);
and U7463 (N_7463,N_6596,N_6989);
or U7464 (N_7464,N_6881,N_6852);
nor U7465 (N_7465,N_6782,N_6613);
or U7466 (N_7466,N_6621,N_6530);
and U7467 (N_7467,N_6536,N_6880);
xnor U7468 (N_7468,N_6809,N_6774);
xor U7469 (N_7469,N_6694,N_6746);
nor U7470 (N_7470,N_6969,N_6835);
and U7471 (N_7471,N_6507,N_6728);
nand U7472 (N_7472,N_6545,N_6850);
or U7473 (N_7473,N_6599,N_6899);
or U7474 (N_7474,N_6694,N_6753);
nand U7475 (N_7475,N_6623,N_6547);
xor U7476 (N_7476,N_6566,N_6821);
nor U7477 (N_7477,N_6876,N_6823);
nand U7478 (N_7478,N_6612,N_6656);
nand U7479 (N_7479,N_6607,N_6580);
nand U7480 (N_7480,N_6891,N_6663);
nor U7481 (N_7481,N_6606,N_6821);
and U7482 (N_7482,N_6646,N_6764);
nand U7483 (N_7483,N_6933,N_6775);
or U7484 (N_7484,N_6827,N_6658);
nor U7485 (N_7485,N_6597,N_6752);
and U7486 (N_7486,N_6709,N_6616);
and U7487 (N_7487,N_6976,N_6783);
nand U7488 (N_7488,N_6975,N_6965);
or U7489 (N_7489,N_6875,N_6583);
nor U7490 (N_7490,N_6943,N_6807);
nand U7491 (N_7491,N_6514,N_6554);
nor U7492 (N_7492,N_6895,N_6736);
nor U7493 (N_7493,N_6947,N_6778);
nand U7494 (N_7494,N_6622,N_6634);
nor U7495 (N_7495,N_6619,N_6705);
xor U7496 (N_7496,N_6974,N_6718);
nand U7497 (N_7497,N_6883,N_6659);
xnor U7498 (N_7498,N_6943,N_6919);
or U7499 (N_7499,N_6533,N_6716);
nor U7500 (N_7500,N_7381,N_7222);
nor U7501 (N_7501,N_7483,N_7051);
nor U7502 (N_7502,N_7333,N_7340);
or U7503 (N_7503,N_7418,N_7213);
and U7504 (N_7504,N_7071,N_7034);
nand U7505 (N_7505,N_7374,N_7150);
nor U7506 (N_7506,N_7154,N_7290);
xor U7507 (N_7507,N_7323,N_7411);
or U7508 (N_7508,N_7301,N_7014);
xnor U7509 (N_7509,N_7389,N_7028);
and U7510 (N_7510,N_7322,N_7457);
nor U7511 (N_7511,N_7405,N_7084);
or U7512 (N_7512,N_7268,N_7189);
and U7513 (N_7513,N_7440,N_7258);
xnor U7514 (N_7514,N_7414,N_7027);
or U7515 (N_7515,N_7209,N_7036);
or U7516 (N_7516,N_7047,N_7168);
nor U7517 (N_7517,N_7196,N_7248);
xor U7518 (N_7518,N_7021,N_7250);
nand U7519 (N_7519,N_7033,N_7151);
and U7520 (N_7520,N_7139,N_7193);
nand U7521 (N_7521,N_7052,N_7184);
nand U7522 (N_7522,N_7498,N_7486);
xor U7523 (N_7523,N_7353,N_7026);
and U7524 (N_7524,N_7306,N_7360);
nand U7525 (N_7525,N_7382,N_7073);
nand U7526 (N_7526,N_7309,N_7284);
and U7527 (N_7527,N_7126,N_7271);
nor U7528 (N_7528,N_7491,N_7128);
or U7529 (N_7529,N_7287,N_7335);
xnor U7530 (N_7530,N_7467,N_7439);
nand U7531 (N_7531,N_7468,N_7143);
and U7532 (N_7532,N_7015,N_7485);
or U7533 (N_7533,N_7078,N_7183);
or U7534 (N_7534,N_7140,N_7198);
nor U7535 (N_7535,N_7424,N_7282);
and U7536 (N_7536,N_7180,N_7165);
or U7537 (N_7537,N_7104,N_7499);
nand U7538 (N_7538,N_7283,N_7155);
nor U7539 (N_7539,N_7002,N_7080);
and U7540 (N_7540,N_7096,N_7495);
or U7541 (N_7541,N_7355,N_7390);
nor U7542 (N_7542,N_7362,N_7227);
or U7543 (N_7543,N_7305,N_7315);
nor U7544 (N_7544,N_7492,N_7138);
and U7545 (N_7545,N_7378,N_7347);
or U7546 (N_7546,N_7386,N_7477);
nand U7547 (N_7547,N_7384,N_7293);
xnor U7548 (N_7548,N_7324,N_7197);
nor U7549 (N_7549,N_7089,N_7387);
and U7550 (N_7550,N_7408,N_7229);
and U7551 (N_7551,N_7063,N_7233);
and U7552 (N_7552,N_7112,N_7211);
or U7553 (N_7553,N_7449,N_7370);
xor U7554 (N_7554,N_7242,N_7101);
or U7555 (N_7555,N_7441,N_7275);
and U7556 (N_7556,N_7019,N_7235);
xnor U7557 (N_7557,N_7373,N_7044);
nor U7558 (N_7558,N_7496,N_7473);
and U7559 (N_7559,N_7296,N_7456);
nor U7560 (N_7560,N_7075,N_7447);
and U7561 (N_7561,N_7228,N_7177);
and U7562 (N_7562,N_7380,N_7115);
nor U7563 (N_7563,N_7095,N_7407);
and U7564 (N_7564,N_7169,N_7016);
or U7565 (N_7565,N_7404,N_7218);
and U7566 (N_7566,N_7035,N_7281);
nor U7567 (N_7567,N_7246,N_7247);
and U7568 (N_7568,N_7182,N_7334);
nand U7569 (N_7569,N_7300,N_7023);
and U7570 (N_7570,N_7307,N_7413);
nor U7571 (N_7571,N_7412,N_7176);
xor U7572 (N_7572,N_7121,N_7348);
nor U7573 (N_7573,N_7158,N_7167);
nand U7574 (N_7574,N_7292,N_7453);
nand U7575 (N_7575,N_7402,N_7039);
or U7576 (N_7576,N_7337,N_7267);
nand U7577 (N_7577,N_7363,N_7256);
or U7578 (N_7578,N_7427,N_7444);
or U7579 (N_7579,N_7472,N_7102);
nor U7580 (N_7580,N_7396,N_7043);
or U7581 (N_7581,N_7142,N_7436);
or U7582 (N_7582,N_7025,N_7480);
nor U7583 (N_7583,N_7001,N_7437);
xor U7584 (N_7584,N_7186,N_7288);
and U7585 (N_7585,N_7215,N_7354);
nor U7586 (N_7586,N_7216,N_7254);
xnor U7587 (N_7587,N_7105,N_7391);
nor U7588 (N_7588,N_7448,N_7316);
xor U7589 (N_7589,N_7311,N_7107);
xnor U7590 (N_7590,N_7310,N_7379);
or U7591 (N_7591,N_7129,N_7147);
nor U7592 (N_7592,N_7372,N_7365);
xnor U7593 (N_7593,N_7127,N_7217);
and U7594 (N_7594,N_7286,N_7137);
nor U7595 (N_7595,N_7383,N_7329);
nand U7596 (N_7596,N_7463,N_7234);
or U7597 (N_7597,N_7156,N_7125);
nor U7598 (N_7598,N_7471,N_7304);
xor U7599 (N_7599,N_7231,N_7050);
or U7600 (N_7600,N_7345,N_7343);
xor U7601 (N_7601,N_7000,N_7313);
and U7602 (N_7602,N_7433,N_7490);
xor U7603 (N_7603,N_7079,N_7270);
xor U7604 (N_7604,N_7067,N_7109);
nand U7605 (N_7605,N_7048,N_7484);
nand U7606 (N_7606,N_7103,N_7114);
and U7607 (N_7607,N_7190,N_7007);
or U7608 (N_7608,N_7116,N_7435);
and U7609 (N_7609,N_7420,N_7022);
nor U7610 (N_7610,N_7342,N_7395);
nand U7611 (N_7611,N_7032,N_7081);
nand U7612 (N_7612,N_7289,N_7450);
nand U7613 (N_7613,N_7132,N_7274);
nor U7614 (N_7614,N_7312,N_7061);
nor U7615 (N_7615,N_7244,N_7291);
nand U7616 (N_7616,N_7219,N_7438);
nor U7617 (N_7617,N_7086,N_7172);
and U7618 (N_7618,N_7469,N_7461);
and U7619 (N_7619,N_7053,N_7245);
nor U7620 (N_7620,N_7331,N_7187);
nor U7621 (N_7621,N_7458,N_7403);
nand U7622 (N_7622,N_7314,N_7120);
and U7623 (N_7623,N_7249,N_7356);
and U7624 (N_7624,N_7462,N_7194);
or U7625 (N_7625,N_7210,N_7263);
and U7626 (N_7626,N_7111,N_7181);
and U7627 (N_7627,N_7170,N_7171);
xor U7628 (N_7628,N_7240,N_7452);
xnor U7629 (N_7629,N_7141,N_7098);
nand U7630 (N_7630,N_7200,N_7376);
nor U7631 (N_7631,N_7358,N_7269);
nor U7632 (N_7632,N_7351,N_7066);
nor U7633 (N_7633,N_7265,N_7350);
xor U7634 (N_7634,N_7020,N_7011);
nand U7635 (N_7635,N_7493,N_7024);
and U7636 (N_7636,N_7070,N_7173);
or U7637 (N_7637,N_7037,N_7366);
xnor U7638 (N_7638,N_7157,N_7057);
nand U7639 (N_7639,N_7401,N_7317);
xor U7640 (N_7640,N_7359,N_7392);
or U7641 (N_7641,N_7415,N_7208);
nand U7642 (N_7642,N_7232,N_7454);
or U7643 (N_7643,N_7065,N_7397);
nor U7644 (N_7644,N_7308,N_7091);
or U7645 (N_7645,N_7161,N_7042);
nor U7646 (N_7646,N_7199,N_7262);
nor U7647 (N_7647,N_7475,N_7224);
nand U7648 (N_7648,N_7017,N_7319);
nand U7649 (N_7649,N_7226,N_7205);
xor U7650 (N_7650,N_7394,N_7174);
nor U7651 (N_7651,N_7178,N_7489);
and U7652 (N_7652,N_7442,N_7009);
or U7653 (N_7653,N_7201,N_7195);
nand U7654 (N_7654,N_7152,N_7478);
xor U7655 (N_7655,N_7136,N_7093);
or U7656 (N_7656,N_7188,N_7432);
nand U7657 (N_7657,N_7464,N_7297);
and U7658 (N_7658,N_7388,N_7191);
and U7659 (N_7659,N_7299,N_7393);
xor U7660 (N_7660,N_7214,N_7398);
or U7661 (N_7661,N_7431,N_7465);
and U7662 (N_7662,N_7417,N_7207);
nor U7663 (N_7663,N_7175,N_7321);
nor U7664 (N_7664,N_7423,N_7164);
nor U7665 (N_7665,N_7399,N_7460);
nor U7666 (N_7666,N_7459,N_7122);
nand U7667 (N_7667,N_7251,N_7425);
and U7668 (N_7668,N_7266,N_7145);
or U7669 (N_7669,N_7082,N_7325);
nor U7670 (N_7670,N_7364,N_7083);
xnor U7671 (N_7671,N_7385,N_7361);
and U7672 (N_7672,N_7367,N_7487);
and U7673 (N_7673,N_7466,N_7099);
nor U7674 (N_7674,N_7088,N_7338);
nand U7675 (N_7675,N_7159,N_7006);
nor U7676 (N_7676,N_7476,N_7430);
and U7677 (N_7677,N_7488,N_7253);
xnor U7678 (N_7678,N_7400,N_7276);
nand U7679 (N_7679,N_7261,N_7069);
nand U7680 (N_7680,N_7236,N_7339);
nand U7681 (N_7681,N_7445,N_7106);
xnor U7682 (N_7682,N_7119,N_7326);
nand U7683 (N_7683,N_7349,N_7260);
xor U7684 (N_7684,N_7076,N_7055);
or U7685 (N_7685,N_7077,N_7153);
or U7686 (N_7686,N_7072,N_7192);
nand U7687 (N_7687,N_7446,N_7357);
or U7688 (N_7688,N_7241,N_7225);
nand U7689 (N_7689,N_7264,N_7278);
xnor U7690 (N_7690,N_7133,N_7030);
and U7691 (N_7691,N_7202,N_7285);
and U7692 (N_7692,N_7074,N_7004);
and U7693 (N_7693,N_7204,N_7045);
or U7694 (N_7694,N_7332,N_7238);
and U7695 (N_7695,N_7494,N_7113);
or U7696 (N_7696,N_7419,N_7010);
nor U7697 (N_7697,N_7406,N_7421);
and U7698 (N_7698,N_7163,N_7124);
xnor U7699 (N_7699,N_7206,N_7482);
and U7700 (N_7700,N_7108,N_7148);
xor U7701 (N_7701,N_7303,N_7123);
or U7702 (N_7702,N_7018,N_7371);
nor U7703 (N_7703,N_7135,N_7062);
nor U7704 (N_7704,N_7474,N_7346);
or U7705 (N_7705,N_7259,N_7318);
xor U7706 (N_7706,N_7220,N_7330);
and U7707 (N_7707,N_7272,N_7443);
nor U7708 (N_7708,N_7279,N_7295);
nor U7709 (N_7709,N_7239,N_7049);
or U7710 (N_7710,N_7162,N_7377);
xnor U7711 (N_7711,N_7230,N_7410);
and U7712 (N_7712,N_7144,N_7255);
nand U7713 (N_7713,N_7455,N_7094);
nor U7714 (N_7714,N_7090,N_7185);
nor U7715 (N_7715,N_7005,N_7257);
nor U7716 (N_7716,N_7059,N_7179);
xnor U7717 (N_7717,N_7092,N_7294);
nand U7718 (N_7718,N_7003,N_7273);
or U7719 (N_7719,N_7479,N_7375);
or U7720 (N_7720,N_7131,N_7428);
nand U7721 (N_7721,N_7277,N_7146);
xor U7722 (N_7722,N_7046,N_7416);
or U7723 (N_7723,N_7203,N_7166);
nor U7724 (N_7724,N_7012,N_7031);
xnor U7725 (N_7725,N_7341,N_7298);
and U7726 (N_7726,N_7100,N_7118);
and U7727 (N_7727,N_7481,N_7344);
and U7728 (N_7728,N_7008,N_7429);
and U7729 (N_7729,N_7060,N_7368);
nor U7730 (N_7730,N_7223,N_7160);
nand U7731 (N_7731,N_7110,N_7280);
xnor U7732 (N_7732,N_7369,N_7054);
xor U7733 (N_7733,N_7117,N_7038);
nand U7734 (N_7734,N_7352,N_7064);
nor U7735 (N_7735,N_7058,N_7097);
or U7736 (N_7736,N_7327,N_7336);
xnor U7737 (N_7737,N_7130,N_7013);
and U7738 (N_7738,N_7422,N_7212);
nand U7739 (N_7739,N_7085,N_7434);
and U7740 (N_7740,N_7320,N_7409);
or U7741 (N_7741,N_7497,N_7237);
nand U7742 (N_7742,N_7056,N_7252);
nor U7743 (N_7743,N_7041,N_7328);
and U7744 (N_7744,N_7149,N_7243);
nand U7745 (N_7745,N_7029,N_7068);
xor U7746 (N_7746,N_7302,N_7087);
and U7747 (N_7747,N_7451,N_7426);
nand U7748 (N_7748,N_7221,N_7470);
and U7749 (N_7749,N_7134,N_7040);
nand U7750 (N_7750,N_7441,N_7203);
and U7751 (N_7751,N_7060,N_7252);
nor U7752 (N_7752,N_7011,N_7420);
nor U7753 (N_7753,N_7345,N_7463);
nand U7754 (N_7754,N_7268,N_7491);
nand U7755 (N_7755,N_7100,N_7409);
and U7756 (N_7756,N_7082,N_7346);
xor U7757 (N_7757,N_7070,N_7065);
nand U7758 (N_7758,N_7065,N_7499);
xnor U7759 (N_7759,N_7051,N_7107);
nor U7760 (N_7760,N_7013,N_7480);
and U7761 (N_7761,N_7139,N_7467);
nor U7762 (N_7762,N_7339,N_7094);
nand U7763 (N_7763,N_7101,N_7356);
xnor U7764 (N_7764,N_7207,N_7175);
nor U7765 (N_7765,N_7135,N_7205);
and U7766 (N_7766,N_7182,N_7039);
nand U7767 (N_7767,N_7104,N_7252);
and U7768 (N_7768,N_7305,N_7042);
or U7769 (N_7769,N_7082,N_7269);
and U7770 (N_7770,N_7321,N_7482);
and U7771 (N_7771,N_7263,N_7011);
nand U7772 (N_7772,N_7167,N_7444);
and U7773 (N_7773,N_7495,N_7174);
nor U7774 (N_7774,N_7009,N_7346);
or U7775 (N_7775,N_7146,N_7188);
and U7776 (N_7776,N_7075,N_7182);
nand U7777 (N_7777,N_7340,N_7148);
and U7778 (N_7778,N_7413,N_7198);
xor U7779 (N_7779,N_7414,N_7391);
xor U7780 (N_7780,N_7214,N_7423);
nor U7781 (N_7781,N_7111,N_7476);
nand U7782 (N_7782,N_7152,N_7497);
nand U7783 (N_7783,N_7288,N_7191);
or U7784 (N_7784,N_7045,N_7447);
or U7785 (N_7785,N_7173,N_7476);
and U7786 (N_7786,N_7005,N_7318);
xor U7787 (N_7787,N_7202,N_7160);
nand U7788 (N_7788,N_7354,N_7116);
xor U7789 (N_7789,N_7037,N_7348);
nand U7790 (N_7790,N_7436,N_7206);
nand U7791 (N_7791,N_7010,N_7109);
xor U7792 (N_7792,N_7085,N_7062);
or U7793 (N_7793,N_7259,N_7251);
nand U7794 (N_7794,N_7420,N_7366);
and U7795 (N_7795,N_7121,N_7211);
nand U7796 (N_7796,N_7173,N_7290);
nand U7797 (N_7797,N_7153,N_7057);
or U7798 (N_7798,N_7093,N_7198);
nand U7799 (N_7799,N_7007,N_7418);
nand U7800 (N_7800,N_7064,N_7039);
and U7801 (N_7801,N_7449,N_7302);
xnor U7802 (N_7802,N_7406,N_7261);
nand U7803 (N_7803,N_7246,N_7029);
and U7804 (N_7804,N_7406,N_7467);
nand U7805 (N_7805,N_7439,N_7291);
nand U7806 (N_7806,N_7390,N_7048);
nor U7807 (N_7807,N_7176,N_7226);
xnor U7808 (N_7808,N_7029,N_7181);
nand U7809 (N_7809,N_7217,N_7229);
and U7810 (N_7810,N_7003,N_7474);
xor U7811 (N_7811,N_7426,N_7472);
xor U7812 (N_7812,N_7230,N_7141);
and U7813 (N_7813,N_7231,N_7225);
xor U7814 (N_7814,N_7286,N_7087);
xnor U7815 (N_7815,N_7077,N_7312);
nor U7816 (N_7816,N_7297,N_7153);
xor U7817 (N_7817,N_7120,N_7432);
and U7818 (N_7818,N_7014,N_7152);
nand U7819 (N_7819,N_7112,N_7354);
nor U7820 (N_7820,N_7148,N_7421);
xor U7821 (N_7821,N_7029,N_7474);
nor U7822 (N_7822,N_7478,N_7349);
xor U7823 (N_7823,N_7060,N_7233);
or U7824 (N_7824,N_7277,N_7140);
xor U7825 (N_7825,N_7481,N_7244);
nor U7826 (N_7826,N_7246,N_7373);
nand U7827 (N_7827,N_7451,N_7242);
nand U7828 (N_7828,N_7245,N_7015);
and U7829 (N_7829,N_7252,N_7319);
nand U7830 (N_7830,N_7380,N_7184);
nand U7831 (N_7831,N_7429,N_7102);
xor U7832 (N_7832,N_7068,N_7439);
and U7833 (N_7833,N_7448,N_7272);
xor U7834 (N_7834,N_7384,N_7460);
or U7835 (N_7835,N_7159,N_7249);
nand U7836 (N_7836,N_7037,N_7164);
or U7837 (N_7837,N_7166,N_7489);
nand U7838 (N_7838,N_7002,N_7495);
and U7839 (N_7839,N_7059,N_7307);
nand U7840 (N_7840,N_7091,N_7059);
nor U7841 (N_7841,N_7355,N_7342);
and U7842 (N_7842,N_7378,N_7206);
nand U7843 (N_7843,N_7129,N_7463);
or U7844 (N_7844,N_7385,N_7271);
nand U7845 (N_7845,N_7456,N_7472);
or U7846 (N_7846,N_7462,N_7215);
nor U7847 (N_7847,N_7016,N_7483);
or U7848 (N_7848,N_7057,N_7011);
nand U7849 (N_7849,N_7144,N_7097);
nor U7850 (N_7850,N_7136,N_7110);
or U7851 (N_7851,N_7300,N_7063);
nand U7852 (N_7852,N_7094,N_7258);
xor U7853 (N_7853,N_7097,N_7402);
and U7854 (N_7854,N_7026,N_7429);
nand U7855 (N_7855,N_7344,N_7254);
nand U7856 (N_7856,N_7205,N_7359);
or U7857 (N_7857,N_7356,N_7054);
nand U7858 (N_7858,N_7313,N_7446);
or U7859 (N_7859,N_7084,N_7288);
or U7860 (N_7860,N_7405,N_7471);
or U7861 (N_7861,N_7144,N_7125);
and U7862 (N_7862,N_7050,N_7435);
xor U7863 (N_7863,N_7134,N_7084);
or U7864 (N_7864,N_7369,N_7483);
and U7865 (N_7865,N_7254,N_7180);
xor U7866 (N_7866,N_7104,N_7498);
xnor U7867 (N_7867,N_7182,N_7434);
or U7868 (N_7868,N_7062,N_7302);
nor U7869 (N_7869,N_7050,N_7342);
nand U7870 (N_7870,N_7256,N_7328);
nor U7871 (N_7871,N_7141,N_7275);
nor U7872 (N_7872,N_7349,N_7012);
or U7873 (N_7873,N_7076,N_7408);
and U7874 (N_7874,N_7333,N_7085);
nor U7875 (N_7875,N_7475,N_7044);
nor U7876 (N_7876,N_7313,N_7424);
nor U7877 (N_7877,N_7080,N_7168);
xnor U7878 (N_7878,N_7435,N_7156);
and U7879 (N_7879,N_7444,N_7250);
nand U7880 (N_7880,N_7102,N_7410);
or U7881 (N_7881,N_7396,N_7398);
nand U7882 (N_7882,N_7118,N_7455);
nand U7883 (N_7883,N_7418,N_7299);
xnor U7884 (N_7884,N_7136,N_7085);
nand U7885 (N_7885,N_7268,N_7047);
nor U7886 (N_7886,N_7394,N_7356);
and U7887 (N_7887,N_7281,N_7268);
xor U7888 (N_7888,N_7446,N_7259);
xnor U7889 (N_7889,N_7279,N_7147);
or U7890 (N_7890,N_7085,N_7234);
nand U7891 (N_7891,N_7009,N_7369);
xor U7892 (N_7892,N_7302,N_7340);
nor U7893 (N_7893,N_7189,N_7192);
nand U7894 (N_7894,N_7098,N_7481);
nand U7895 (N_7895,N_7199,N_7316);
nor U7896 (N_7896,N_7336,N_7163);
or U7897 (N_7897,N_7117,N_7149);
or U7898 (N_7898,N_7001,N_7195);
and U7899 (N_7899,N_7283,N_7018);
nand U7900 (N_7900,N_7426,N_7217);
xnor U7901 (N_7901,N_7466,N_7473);
nor U7902 (N_7902,N_7225,N_7499);
nor U7903 (N_7903,N_7444,N_7395);
and U7904 (N_7904,N_7329,N_7295);
or U7905 (N_7905,N_7001,N_7123);
nor U7906 (N_7906,N_7393,N_7159);
or U7907 (N_7907,N_7162,N_7491);
xor U7908 (N_7908,N_7077,N_7065);
or U7909 (N_7909,N_7461,N_7156);
nand U7910 (N_7910,N_7173,N_7061);
or U7911 (N_7911,N_7412,N_7258);
or U7912 (N_7912,N_7294,N_7486);
nand U7913 (N_7913,N_7220,N_7083);
xor U7914 (N_7914,N_7208,N_7196);
or U7915 (N_7915,N_7003,N_7062);
and U7916 (N_7916,N_7454,N_7158);
nor U7917 (N_7917,N_7014,N_7164);
nor U7918 (N_7918,N_7117,N_7100);
xor U7919 (N_7919,N_7060,N_7407);
xor U7920 (N_7920,N_7357,N_7136);
and U7921 (N_7921,N_7274,N_7065);
nor U7922 (N_7922,N_7113,N_7049);
or U7923 (N_7923,N_7495,N_7078);
or U7924 (N_7924,N_7239,N_7300);
nand U7925 (N_7925,N_7332,N_7180);
xnor U7926 (N_7926,N_7238,N_7103);
or U7927 (N_7927,N_7458,N_7116);
and U7928 (N_7928,N_7361,N_7232);
xor U7929 (N_7929,N_7253,N_7109);
and U7930 (N_7930,N_7120,N_7387);
and U7931 (N_7931,N_7341,N_7228);
nand U7932 (N_7932,N_7484,N_7237);
nor U7933 (N_7933,N_7072,N_7228);
nor U7934 (N_7934,N_7333,N_7130);
or U7935 (N_7935,N_7343,N_7008);
and U7936 (N_7936,N_7418,N_7231);
nand U7937 (N_7937,N_7133,N_7427);
xnor U7938 (N_7938,N_7445,N_7457);
or U7939 (N_7939,N_7311,N_7498);
or U7940 (N_7940,N_7481,N_7101);
nand U7941 (N_7941,N_7249,N_7290);
nor U7942 (N_7942,N_7384,N_7137);
nand U7943 (N_7943,N_7397,N_7362);
xor U7944 (N_7944,N_7066,N_7386);
xnor U7945 (N_7945,N_7309,N_7182);
nand U7946 (N_7946,N_7333,N_7386);
and U7947 (N_7947,N_7000,N_7197);
nor U7948 (N_7948,N_7419,N_7389);
and U7949 (N_7949,N_7085,N_7330);
nand U7950 (N_7950,N_7174,N_7428);
and U7951 (N_7951,N_7388,N_7219);
xor U7952 (N_7952,N_7223,N_7193);
nor U7953 (N_7953,N_7497,N_7095);
and U7954 (N_7954,N_7435,N_7213);
and U7955 (N_7955,N_7358,N_7215);
nand U7956 (N_7956,N_7110,N_7413);
nand U7957 (N_7957,N_7202,N_7427);
xor U7958 (N_7958,N_7420,N_7460);
and U7959 (N_7959,N_7249,N_7444);
nor U7960 (N_7960,N_7273,N_7397);
xnor U7961 (N_7961,N_7205,N_7343);
or U7962 (N_7962,N_7231,N_7316);
nor U7963 (N_7963,N_7259,N_7205);
nor U7964 (N_7964,N_7423,N_7343);
or U7965 (N_7965,N_7387,N_7447);
or U7966 (N_7966,N_7391,N_7025);
xnor U7967 (N_7967,N_7157,N_7434);
nor U7968 (N_7968,N_7333,N_7151);
or U7969 (N_7969,N_7086,N_7497);
or U7970 (N_7970,N_7356,N_7387);
nand U7971 (N_7971,N_7164,N_7258);
nor U7972 (N_7972,N_7287,N_7470);
xor U7973 (N_7973,N_7483,N_7443);
or U7974 (N_7974,N_7261,N_7235);
nor U7975 (N_7975,N_7448,N_7110);
and U7976 (N_7976,N_7273,N_7461);
nor U7977 (N_7977,N_7037,N_7235);
xor U7978 (N_7978,N_7374,N_7303);
nand U7979 (N_7979,N_7446,N_7460);
xnor U7980 (N_7980,N_7025,N_7016);
nor U7981 (N_7981,N_7374,N_7432);
nand U7982 (N_7982,N_7213,N_7451);
and U7983 (N_7983,N_7335,N_7005);
nor U7984 (N_7984,N_7152,N_7151);
xnor U7985 (N_7985,N_7048,N_7074);
or U7986 (N_7986,N_7161,N_7052);
and U7987 (N_7987,N_7089,N_7449);
or U7988 (N_7988,N_7290,N_7086);
or U7989 (N_7989,N_7123,N_7418);
xnor U7990 (N_7990,N_7110,N_7493);
and U7991 (N_7991,N_7159,N_7149);
nor U7992 (N_7992,N_7364,N_7283);
and U7993 (N_7993,N_7080,N_7228);
nand U7994 (N_7994,N_7270,N_7025);
xnor U7995 (N_7995,N_7323,N_7217);
xnor U7996 (N_7996,N_7192,N_7473);
and U7997 (N_7997,N_7232,N_7241);
xnor U7998 (N_7998,N_7209,N_7444);
or U7999 (N_7999,N_7453,N_7321);
nand U8000 (N_8000,N_7870,N_7864);
or U8001 (N_8001,N_7680,N_7625);
or U8002 (N_8002,N_7552,N_7783);
or U8003 (N_8003,N_7745,N_7645);
nand U8004 (N_8004,N_7767,N_7940);
or U8005 (N_8005,N_7577,N_7535);
nor U8006 (N_8006,N_7628,N_7950);
and U8007 (N_8007,N_7749,N_7525);
nand U8008 (N_8008,N_7939,N_7534);
nand U8009 (N_8009,N_7918,N_7548);
or U8010 (N_8010,N_7545,N_7520);
nand U8011 (N_8011,N_7995,N_7543);
nand U8012 (N_8012,N_7523,N_7937);
and U8013 (N_8013,N_7629,N_7536);
nand U8014 (N_8014,N_7764,N_7926);
nor U8015 (N_8015,N_7696,N_7959);
nor U8016 (N_8016,N_7921,N_7707);
or U8017 (N_8017,N_7916,N_7507);
nor U8018 (N_8018,N_7579,N_7729);
xnor U8019 (N_8019,N_7681,N_7989);
and U8020 (N_8020,N_7831,N_7857);
or U8021 (N_8021,N_7955,N_7717);
or U8022 (N_8022,N_7566,N_7692);
or U8023 (N_8023,N_7938,N_7758);
or U8024 (N_8024,N_7683,N_7691);
and U8025 (N_8025,N_7952,N_7732);
nand U8026 (N_8026,N_7929,N_7632);
or U8027 (N_8027,N_7798,N_7542);
or U8028 (N_8028,N_7866,N_7801);
xnor U8029 (N_8029,N_7725,N_7816);
nand U8030 (N_8030,N_7787,N_7568);
nand U8031 (N_8031,N_7872,N_7634);
nor U8032 (N_8032,N_7742,N_7901);
nor U8033 (N_8033,N_7968,N_7792);
nand U8034 (N_8034,N_7606,N_7698);
and U8035 (N_8035,N_7987,N_7641);
nand U8036 (N_8036,N_7694,N_7677);
nor U8037 (N_8037,N_7956,N_7890);
nor U8038 (N_8038,N_7540,N_7687);
and U8039 (N_8039,N_7867,N_7927);
nand U8040 (N_8040,N_7999,N_7903);
nand U8041 (N_8041,N_7560,N_7796);
xor U8042 (N_8042,N_7815,N_7851);
nand U8043 (N_8043,N_7727,N_7817);
xnor U8044 (N_8044,N_7704,N_7856);
xor U8045 (N_8045,N_7557,N_7572);
nand U8046 (N_8046,N_7573,N_7909);
nor U8047 (N_8047,N_7919,N_7752);
xnor U8048 (N_8048,N_7514,N_7904);
or U8049 (N_8049,N_7547,N_7669);
or U8050 (N_8050,N_7527,N_7617);
and U8051 (N_8051,N_7762,N_7781);
or U8052 (N_8052,N_7737,N_7602);
and U8053 (N_8053,N_7873,N_7772);
xor U8054 (N_8054,N_7795,N_7728);
xor U8055 (N_8055,N_7612,N_7679);
or U8056 (N_8056,N_7848,N_7825);
or U8057 (N_8057,N_7649,N_7978);
nand U8058 (N_8058,N_7779,N_7963);
nor U8059 (N_8059,N_7503,N_7891);
nor U8060 (N_8060,N_7914,N_7674);
or U8061 (N_8061,N_7554,N_7622);
or U8062 (N_8062,N_7569,N_7824);
and U8063 (N_8063,N_7899,N_7946);
and U8064 (N_8064,N_7847,N_7807);
nor U8065 (N_8065,N_7650,N_7934);
or U8066 (N_8066,N_7733,N_7794);
nor U8067 (N_8067,N_7721,N_7593);
and U8068 (N_8068,N_7962,N_7667);
and U8069 (N_8069,N_7763,N_7510);
or U8070 (N_8070,N_7853,N_7591);
or U8071 (N_8071,N_7666,N_7609);
and U8072 (N_8072,N_7556,N_7965);
nor U8073 (N_8073,N_7971,N_7601);
nor U8074 (N_8074,N_7912,N_7574);
nand U8075 (N_8075,N_7553,N_7583);
nand U8076 (N_8076,N_7673,N_7699);
or U8077 (N_8077,N_7973,N_7607);
or U8078 (N_8078,N_7874,N_7835);
or U8079 (N_8079,N_7690,N_7842);
or U8080 (N_8080,N_7880,N_7878);
nand U8081 (N_8081,N_7898,N_7636);
nor U8082 (N_8082,N_7539,N_7608);
or U8083 (N_8083,N_7822,N_7706);
xnor U8084 (N_8084,N_7935,N_7575);
nor U8085 (N_8085,N_7998,N_7715);
xor U8086 (N_8086,N_7659,N_7757);
and U8087 (N_8087,N_7741,N_7718);
or U8088 (N_8088,N_7664,N_7885);
xor U8089 (N_8089,N_7521,N_7723);
nor U8090 (N_8090,N_7977,N_7562);
nor U8091 (N_8091,N_7571,N_7653);
nand U8092 (N_8092,N_7695,N_7614);
and U8093 (N_8093,N_7689,N_7746);
nor U8094 (N_8094,N_7906,N_7887);
or U8095 (N_8095,N_7697,N_7708);
xnor U8096 (N_8096,N_7850,N_7892);
and U8097 (N_8097,N_7982,N_7981);
nand U8098 (N_8098,N_7902,N_7626);
nand U8099 (N_8099,N_7654,N_7502);
and U8100 (N_8100,N_7592,N_7883);
nor U8101 (N_8101,N_7972,N_7668);
or U8102 (N_8102,N_7671,N_7778);
and U8103 (N_8103,N_7701,N_7945);
and U8104 (N_8104,N_7685,N_7893);
xor U8105 (N_8105,N_7970,N_7549);
xnor U8106 (N_8106,N_7537,N_7907);
nor U8107 (N_8107,N_7643,N_7505);
or U8108 (N_8108,N_7693,N_7845);
xnor U8109 (N_8109,N_7802,N_7623);
or U8110 (N_8110,N_7805,N_7777);
and U8111 (N_8111,N_7513,N_7944);
and U8112 (N_8112,N_7610,N_7586);
xor U8113 (N_8113,N_7604,N_7790);
and U8114 (N_8114,N_7541,N_7900);
nor U8115 (N_8115,N_7877,N_7594);
nor U8116 (N_8116,N_7911,N_7598);
xnor U8117 (N_8117,N_7682,N_7797);
and U8118 (N_8118,N_7735,N_7960);
or U8119 (N_8119,N_7600,N_7886);
or U8120 (N_8120,N_7841,N_7849);
xnor U8121 (N_8121,N_7544,N_7776);
or U8122 (N_8122,N_7923,N_7633);
and U8123 (N_8123,N_7941,N_7879);
nand U8124 (N_8124,N_7821,N_7518);
and U8125 (N_8125,N_7766,N_7843);
nand U8126 (N_8126,N_7538,N_7894);
or U8127 (N_8127,N_7932,N_7871);
and U8128 (N_8128,N_7730,N_7876);
nor U8129 (N_8129,N_7588,N_7551);
and U8130 (N_8130,N_7834,N_7522);
or U8131 (N_8131,N_7905,N_7512);
or U8132 (N_8132,N_7760,N_7975);
nand U8133 (N_8133,N_7589,N_7996);
and U8134 (N_8134,N_7550,N_7726);
and U8135 (N_8135,N_7770,N_7581);
nor U8136 (N_8136,N_7785,N_7823);
nand U8137 (N_8137,N_7517,N_7615);
or U8138 (N_8138,N_7930,N_7931);
nand U8139 (N_8139,N_7859,N_7703);
or U8140 (N_8140,N_7670,N_7678);
xor U8141 (N_8141,N_7528,N_7736);
and U8142 (N_8142,N_7846,N_7624);
or U8143 (N_8143,N_7854,N_7928);
nor U8144 (N_8144,N_7951,N_7774);
and U8145 (N_8145,N_7747,N_7943);
or U8146 (N_8146,N_7976,N_7958);
or U8147 (N_8147,N_7675,N_7631);
nor U8148 (N_8148,N_7936,N_7660);
nor U8149 (N_8149,N_7786,N_7563);
nor U8150 (N_8150,N_7565,N_7910);
or U8151 (N_8151,N_7642,N_7710);
xnor U8152 (N_8152,N_7861,N_7947);
or U8153 (N_8153,N_7637,N_7827);
xor U8154 (N_8154,N_7705,N_7804);
nand U8155 (N_8155,N_7780,N_7888);
and U8156 (N_8156,N_7775,N_7855);
xnor U8157 (N_8157,N_7869,N_7724);
nand U8158 (N_8158,N_7754,N_7915);
and U8159 (N_8159,N_7639,N_7702);
or U8160 (N_8160,N_7875,N_7722);
and U8161 (N_8161,N_7686,N_7896);
or U8162 (N_8162,N_7509,N_7922);
and U8163 (N_8163,N_7578,N_7753);
nor U8164 (N_8164,N_7812,N_7748);
nand U8165 (N_8165,N_7948,N_7840);
xor U8166 (N_8166,N_7655,N_7720);
xnor U8167 (N_8167,N_7858,N_7828);
or U8168 (N_8168,N_7515,N_7969);
nand U8169 (N_8169,N_7913,N_7844);
nor U8170 (N_8170,N_7992,N_7627);
and U8171 (N_8171,N_7576,N_7833);
or U8172 (N_8172,N_7529,N_7961);
or U8173 (N_8173,N_7743,N_7744);
nand U8174 (N_8174,N_7789,N_7665);
and U8175 (N_8175,N_7558,N_7567);
or U8176 (N_8176,N_7852,N_7897);
xor U8177 (N_8177,N_7676,N_7799);
xor U8178 (N_8178,N_7587,N_7908);
or U8179 (N_8179,N_7803,N_7773);
nand U8180 (N_8180,N_7983,N_7646);
nor U8181 (N_8181,N_7719,N_7635);
or U8182 (N_8182,N_7994,N_7769);
xnor U8183 (N_8183,N_7832,N_7647);
nand U8184 (N_8184,N_7818,N_7644);
or U8185 (N_8185,N_7533,N_7986);
nand U8186 (N_8186,N_7964,N_7920);
nor U8187 (N_8187,N_7613,N_7688);
nand U8188 (N_8188,N_7838,N_7806);
nand U8189 (N_8189,N_7656,N_7788);
and U8190 (N_8190,N_7648,N_7530);
xor U8191 (N_8191,N_7739,N_7811);
xor U8192 (N_8192,N_7813,N_7755);
nand U8193 (N_8193,N_7657,N_7651);
and U8194 (N_8194,N_7917,N_7555);
or U8195 (N_8195,N_7889,N_7712);
and U8196 (N_8196,N_7991,N_7546);
xor U8197 (N_8197,N_7953,N_7784);
xnor U8198 (N_8198,N_7988,N_7782);
and U8199 (N_8199,N_7862,N_7768);
or U8200 (N_8200,N_7611,N_7532);
nor U8201 (N_8201,N_7662,N_7761);
and U8202 (N_8202,N_7597,N_7700);
nand U8203 (N_8203,N_7511,N_7564);
xnor U8204 (N_8204,N_7500,N_7711);
xor U8205 (N_8205,N_7621,N_7508);
nor U8206 (N_8206,N_7814,N_7584);
and U8207 (N_8207,N_7925,N_7882);
nand U8208 (N_8208,N_7504,N_7618);
nor U8209 (N_8209,N_7709,N_7516);
nand U8210 (N_8210,N_7808,N_7590);
xor U8211 (N_8211,N_7949,N_7638);
nand U8212 (N_8212,N_7865,N_7884);
nor U8213 (N_8213,N_7501,N_7716);
or U8214 (N_8214,N_7984,N_7661);
nor U8215 (N_8215,N_7979,N_7596);
xnor U8216 (N_8216,N_7658,N_7559);
and U8217 (N_8217,N_7759,N_7595);
or U8218 (N_8218,N_7997,N_7526);
or U8219 (N_8219,N_7966,N_7837);
and U8220 (N_8220,N_7531,N_7895);
and U8221 (N_8221,N_7830,N_7771);
nor U8222 (N_8222,N_7570,N_7993);
xnor U8223 (N_8223,N_7868,N_7751);
xnor U8224 (N_8224,N_7630,N_7738);
and U8225 (N_8225,N_7616,N_7985);
nand U8226 (N_8226,N_7603,N_7605);
nor U8227 (N_8227,N_7974,N_7640);
and U8228 (N_8228,N_7734,N_7839);
or U8229 (N_8229,N_7524,N_7582);
or U8230 (N_8230,N_7980,N_7765);
xnor U8231 (N_8231,N_7967,N_7933);
and U8232 (N_8232,N_7672,N_7826);
nand U8233 (N_8233,N_7829,N_7810);
and U8234 (N_8234,N_7561,N_7506);
nor U8235 (N_8235,N_7819,N_7519);
and U8236 (N_8236,N_7990,N_7836);
or U8237 (N_8237,N_7820,N_7740);
or U8238 (N_8238,N_7800,N_7580);
or U8239 (N_8239,N_7756,N_7957);
and U8240 (N_8240,N_7731,N_7599);
nor U8241 (N_8241,N_7750,N_7954);
nand U8242 (N_8242,N_7863,N_7942);
and U8243 (N_8243,N_7585,N_7881);
nor U8244 (N_8244,N_7793,N_7714);
xnor U8245 (N_8245,N_7619,N_7713);
xnor U8246 (N_8246,N_7663,N_7652);
and U8247 (N_8247,N_7809,N_7924);
nor U8248 (N_8248,N_7860,N_7620);
and U8249 (N_8249,N_7684,N_7791);
nand U8250 (N_8250,N_7879,N_7719);
and U8251 (N_8251,N_7628,N_7698);
or U8252 (N_8252,N_7511,N_7939);
xnor U8253 (N_8253,N_7958,N_7906);
nand U8254 (N_8254,N_7985,N_7569);
and U8255 (N_8255,N_7675,N_7853);
nor U8256 (N_8256,N_7577,N_7712);
nor U8257 (N_8257,N_7668,N_7804);
or U8258 (N_8258,N_7752,N_7881);
and U8259 (N_8259,N_7882,N_7514);
xor U8260 (N_8260,N_7545,N_7728);
and U8261 (N_8261,N_7567,N_7638);
and U8262 (N_8262,N_7609,N_7500);
xor U8263 (N_8263,N_7809,N_7797);
or U8264 (N_8264,N_7727,N_7978);
xor U8265 (N_8265,N_7685,N_7552);
xor U8266 (N_8266,N_7776,N_7597);
xor U8267 (N_8267,N_7514,N_7705);
or U8268 (N_8268,N_7972,N_7738);
and U8269 (N_8269,N_7996,N_7653);
and U8270 (N_8270,N_7997,N_7849);
xnor U8271 (N_8271,N_7572,N_7648);
and U8272 (N_8272,N_7741,N_7751);
nand U8273 (N_8273,N_7952,N_7659);
xor U8274 (N_8274,N_7961,N_7875);
nand U8275 (N_8275,N_7767,N_7747);
or U8276 (N_8276,N_7861,N_7957);
nand U8277 (N_8277,N_7542,N_7568);
and U8278 (N_8278,N_7824,N_7815);
xor U8279 (N_8279,N_7742,N_7798);
nand U8280 (N_8280,N_7780,N_7841);
nor U8281 (N_8281,N_7767,N_7980);
or U8282 (N_8282,N_7943,N_7679);
and U8283 (N_8283,N_7976,N_7511);
or U8284 (N_8284,N_7874,N_7882);
xor U8285 (N_8285,N_7687,N_7965);
nand U8286 (N_8286,N_7661,N_7727);
nand U8287 (N_8287,N_7614,N_7913);
nand U8288 (N_8288,N_7618,N_7726);
nor U8289 (N_8289,N_7812,N_7668);
or U8290 (N_8290,N_7672,N_7695);
nor U8291 (N_8291,N_7565,N_7988);
nand U8292 (N_8292,N_7611,N_7725);
nor U8293 (N_8293,N_7822,N_7811);
nand U8294 (N_8294,N_7564,N_7570);
xnor U8295 (N_8295,N_7563,N_7734);
and U8296 (N_8296,N_7788,N_7974);
xnor U8297 (N_8297,N_7517,N_7608);
xor U8298 (N_8298,N_7738,N_7577);
nand U8299 (N_8299,N_7942,N_7887);
xor U8300 (N_8300,N_7929,N_7577);
xnor U8301 (N_8301,N_7624,N_7673);
nand U8302 (N_8302,N_7522,N_7766);
xnor U8303 (N_8303,N_7657,N_7762);
xor U8304 (N_8304,N_7562,N_7612);
nand U8305 (N_8305,N_7744,N_7662);
and U8306 (N_8306,N_7724,N_7668);
and U8307 (N_8307,N_7688,N_7546);
nand U8308 (N_8308,N_7713,N_7727);
nand U8309 (N_8309,N_7847,N_7534);
xnor U8310 (N_8310,N_7718,N_7639);
nand U8311 (N_8311,N_7696,N_7885);
xor U8312 (N_8312,N_7858,N_7958);
nand U8313 (N_8313,N_7988,N_7948);
or U8314 (N_8314,N_7808,N_7882);
nand U8315 (N_8315,N_7515,N_7938);
and U8316 (N_8316,N_7850,N_7942);
xnor U8317 (N_8317,N_7906,N_7731);
and U8318 (N_8318,N_7894,N_7909);
and U8319 (N_8319,N_7508,N_7516);
nand U8320 (N_8320,N_7962,N_7919);
nor U8321 (N_8321,N_7549,N_7814);
nand U8322 (N_8322,N_7500,N_7700);
nand U8323 (N_8323,N_7910,N_7957);
nor U8324 (N_8324,N_7524,N_7790);
and U8325 (N_8325,N_7513,N_7701);
and U8326 (N_8326,N_7928,N_7746);
nor U8327 (N_8327,N_7777,N_7722);
and U8328 (N_8328,N_7902,N_7717);
and U8329 (N_8329,N_7530,N_7501);
xor U8330 (N_8330,N_7539,N_7520);
or U8331 (N_8331,N_7814,N_7905);
or U8332 (N_8332,N_7624,N_7681);
or U8333 (N_8333,N_7791,N_7969);
or U8334 (N_8334,N_7638,N_7741);
and U8335 (N_8335,N_7993,N_7501);
nor U8336 (N_8336,N_7978,N_7698);
nand U8337 (N_8337,N_7803,N_7704);
xor U8338 (N_8338,N_7881,N_7900);
and U8339 (N_8339,N_7879,N_7578);
xor U8340 (N_8340,N_7972,N_7599);
nor U8341 (N_8341,N_7917,N_7718);
and U8342 (N_8342,N_7982,N_7956);
nand U8343 (N_8343,N_7808,N_7539);
or U8344 (N_8344,N_7544,N_7921);
nor U8345 (N_8345,N_7736,N_7604);
nand U8346 (N_8346,N_7510,N_7779);
nand U8347 (N_8347,N_7802,N_7599);
or U8348 (N_8348,N_7788,N_7557);
or U8349 (N_8349,N_7684,N_7800);
xnor U8350 (N_8350,N_7796,N_7916);
or U8351 (N_8351,N_7675,N_7839);
nor U8352 (N_8352,N_7564,N_7783);
and U8353 (N_8353,N_7991,N_7736);
nand U8354 (N_8354,N_7729,N_7897);
and U8355 (N_8355,N_7751,N_7853);
or U8356 (N_8356,N_7578,N_7943);
nand U8357 (N_8357,N_7524,N_7600);
xnor U8358 (N_8358,N_7840,N_7721);
nand U8359 (N_8359,N_7787,N_7565);
xnor U8360 (N_8360,N_7626,N_7961);
or U8361 (N_8361,N_7825,N_7833);
nand U8362 (N_8362,N_7990,N_7903);
or U8363 (N_8363,N_7705,N_7722);
nor U8364 (N_8364,N_7602,N_7698);
xor U8365 (N_8365,N_7538,N_7645);
nand U8366 (N_8366,N_7699,N_7623);
xor U8367 (N_8367,N_7975,N_7795);
and U8368 (N_8368,N_7836,N_7780);
nand U8369 (N_8369,N_7747,N_7888);
or U8370 (N_8370,N_7918,N_7927);
or U8371 (N_8371,N_7700,N_7987);
nand U8372 (N_8372,N_7722,N_7932);
nand U8373 (N_8373,N_7936,N_7576);
or U8374 (N_8374,N_7704,N_7962);
nand U8375 (N_8375,N_7897,N_7782);
or U8376 (N_8376,N_7773,N_7706);
or U8377 (N_8377,N_7972,N_7602);
nand U8378 (N_8378,N_7671,N_7669);
nor U8379 (N_8379,N_7810,N_7761);
and U8380 (N_8380,N_7516,N_7529);
xor U8381 (N_8381,N_7561,N_7743);
nand U8382 (N_8382,N_7772,N_7842);
and U8383 (N_8383,N_7981,N_7877);
xnor U8384 (N_8384,N_7970,N_7563);
nor U8385 (N_8385,N_7516,N_7938);
nor U8386 (N_8386,N_7615,N_7879);
xnor U8387 (N_8387,N_7989,N_7838);
and U8388 (N_8388,N_7684,N_7517);
nand U8389 (N_8389,N_7587,N_7828);
xnor U8390 (N_8390,N_7519,N_7670);
nor U8391 (N_8391,N_7610,N_7773);
xnor U8392 (N_8392,N_7898,N_7952);
nand U8393 (N_8393,N_7576,N_7642);
and U8394 (N_8394,N_7511,N_7774);
or U8395 (N_8395,N_7817,N_7818);
and U8396 (N_8396,N_7680,N_7838);
and U8397 (N_8397,N_7713,N_7956);
and U8398 (N_8398,N_7802,N_7944);
and U8399 (N_8399,N_7974,N_7910);
nor U8400 (N_8400,N_7937,N_7537);
or U8401 (N_8401,N_7660,N_7962);
nor U8402 (N_8402,N_7595,N_7896);
nor U8403 (N_8403,N_7782,N_7955);
nor U8404 (N_8404,N_7616,N_7604);
or U8405 (N_8405,N_7705,N_7783);
and U8406 (N_8406,N_7670,N_7788);
xnor U8407 (N_8407,N_7944,N_7568);
and U8408 (N_8408,N_7567,N_7752);
xor U8409 (N_8409,N_7867,N_7748);
nand U8410 (N_8410,N_7969,N_7675);
and U8411 (N_8411,N_7801,N_7582);
nand U8412 (N_8412,N_7932,N_7850);
or U8413 (N_8413,N_7798,N_7856);
or U8414 (N_8414,N_7551,N_7510);
nand U8415 (N_8415,N_7724,N_7903);
and U8416 (N_8416,N_7734,N_7785);
nand U8417 (N_8417,N_7507,N_7854);
xor U8418 (N_8418,N_7565,N_7563);
nor U8419 (N_8419,N_7787,N_7701);
and U8420 (N_8420,N_7506,N_7895);
nand U8421 (N_8421,N_7768,N_7724);
xor U8422 (N_8422,N_7982,N_7965);
nor U8423 (N_8423,N_7817,N_7576);
nor U8424 (N_8424,N_7658,N_7705);
nand U8425 (N_8425,N_7559,N_7887);
nor U8426 (N_8426,N_7522,N_7559);
nand U8427 (N_8427,N_7951,N_7730);
xor U8428 (N_8428,N_7762,N_7814);
nor U8429 (N_8429,N_7886,N_7815);
nand U8430 (N_8430,N_7777,N_7677);
and U8431 (N_8431,N_7683,N_7710);
and U8432 (N_8432,N_7693,N_7679);
nor U8433 (N_8433,N_7681,N_7751);
nor U8434 (N_8434,N_7921,N_7537);
and U8435 (N_8435,N_7647,N_7718);
and U8436 (N_8436,N_7517,N_7704);
nand U8437 (N_8437,N_7936,N_7793);
xnor U8438 (N_8438,N_7687,N_7684);
nor U8439 (N_8439,N_7975,N_7669);
or U8440 (N_8440,N_7688,N_7616);
and U8441 (N_8441,N_7881,N_7643);
or U8442 (N_8442,N_7986,N_7588);
nand U8443 (N_8443,N_7626,N_7656);
nand U8444 (N_8444,N_7526,N_7728);
and U8445 (N_8445,N_7652,N_7549);
nor U8446 (N_8446,N_7770,N_7648);
nand U8447 (N_8447,N_7531,N_7938);
xnor U8448 (N_8448,N_7661,N_7681);
and U8449 (N_8449,N_7901,N_7976);
or U8450 (N_8450,N_7573,N_7858);
and U8451 (N_8451,N_7523,N_7514);
nor U8452 (N_8452,N_7697,N_7519);
nor U8453 (N_8453,N_7688,N_7662);
nand U8454 (N_8454,N_7922,N_7657);
nand U8455 (N_8455,N_7939,N_7954);
nor U8456 (N_8456,N_7792,N_7688);
nand U8457 (N_8457,N_7955,N_7884);
xor U8458 (N_8458,N_7667,N_7975);
nor U8459 (N_8459,N_7559,N_7562);
nand U8460 (N_8460,N_7854,N_7632);
nor U8461 (N_8461,N_7937,N_7936);
nor U8462 (N_8462,N_7586,N_7712);
xnor U8463 (N_8463,N_7723,N_7978);
nor U8464 (N_8464,N_7941,N_7784);
and U8465 (N_8465,N_7807,N_7915);
nand U8466 (N_8466,N_7870,N_7989);
or U8467 (N_8467,N_7670,N_7879);
nor U8468 (N_8468,N_7750,N_7828);
nor U8469 (N_8469,N_7893,N_7573);
nand U8470 (N_8470,N_7960,N_7550);
xnor U8471 (N_8471,N_7970,N_7727);
and U8472 (N_8472,N_7956,N_7826);
and U8473 (N_8473,N_7570,N_7653);
nand U8474 (N_8474,N_7814,N_7697);
nand U8475 (N_8475,N_7731,N_7811);
or U8476 (N_8476,N_7876,N_7613);
or U8477 (N_8477,N_7719,N_7918);
xnor U8478 (N_8478,N_7926,N_7674);
nand U8479 (N_8479,N_7821,N_7951);
and U8480 (N_8480,N_7891,N_7802);
nand U8481 (N_8481,N_7815,N_7603);
xor U8482 (N_8482,N_7696,N_7907);
xnor U8483 (N_8483,N_7811,N_7523);
or U8484 (N_8484,N_7521,N_7677);
or U8485 (N_8485,N_7934,N_7676);
nand U8486 (N_8486,N_7962,N_7906);
xnor U8487 (N_8487,N_7679,N_7783);
and U8488 (N_8488,N_7562,N_7702);
or U8489 (N_8489,N_7874,N_7732);
and U8490 (N_8490,N_7788,N_7612);
nor U8491 (N_8491,N_7735,N_7824);
nand U8492 (N_8492,N_7583,N_7890);
and U8493 (N_8493,N_7695,N_7753);
nor U8494 (N_8494,N_7987,N_7609);
nor U8495 (N_8495,N_7693,N_7831);
nand U8496 (N_8496,N_7687,N_7966);
xnor U8497 (N_8497,N_7919,N_7809);
nand U8498 (N_8498,N_7671,N_7813);
nand U8499 (N_8499,N_7757,N_7598);
and U8500 (N_8500,N_8274,N_8442);
and U8501 (N_8501,N_8022,N_8306);
and U8502 (N_8502,N_8480,N_8178);
or U8503 (N_8503,N_8266,N_8261);
or U8504 (N_8504,N_8408,N_8337);
and U8505 (N_8505,N_8237,N_8453);
nor U8506 (N_8506,N_8210,N_8315);
nor U8507 (N_8507,N_8486,N_8054);
and U8508 (N_8508,N_8186,N_8242);
or U8509 (N_8509,N_8025,N_8427);
or U8510 (N_8510,N_8253,N_8272);
or U8511 (N_8511,N_8461,N_8437);
nand U8512 (N_8512,N_8343,N_8355);
xor U8513 (N_8513,N_8299,N_8038);
xnor U8514 (N_8514,N_8198,N_8405);
or U8515 (N_8515,N_8234,N_8216);
nor U8516 (N_8516,N_8397,N_8466);
nand U8517 (N_8517,N_8016,N_8230);
or U8518 (N_8518,N_8106,N_8262);
nand U8519 (N_8519,N_8363,N_8339);
or U8520 (N_8520,N_8460,N_8148);
nand U8521 (N_8521,N_8328,N_8130);
nor U8522 (N_8522,N_8100,N_8428);
nand U8523 (N_8523,N_8477,N_8332);
or U8524 (N_8524,N_8029,N_8206);
xnor U8525 (N_8525,N_8043,N_8215);
and U8526 (N_8526,N_8050,N_8135);
xor U8527 (N_8527,N_8137,N_8103);
or U8528 (N_8528,N_8340,N_8244);
nand U8529 (N_8529,N_8387,N_8342);
xnor U8530 (N_8530,N_8011,N_8170);
and U8531 (N_8531,N_8443,N_8245);
and U8532 (N_8532,N_8000,N_8147);
xor U8533 (N_8533,N_8324,N_8371);
nand U8534 (N_8534,N_8260,N_8149);
or U8535 (N_8535,N_8412,N_8194);
or U8536 (N_8536,N_8113,N_8400);
nor U8537 (N_8537,N_8150,N_8346);
or U8538 (N_8538,N_8456,N_8138);
or U8539 (N_8539,N_8421,N_8468);
xnor U8540 (N_8540,N_8192,N_8263);
and U8541 (N_8541,N_8154,N_8096);
nand U8542 (N_8542,N_8065,N_8241);
nor U8543 (N_8543,N_8479,N_8284);
and U8544 (N_8544,N_8356,N_8490);
or U8545 (N_8545,N_8099,N_8478);
or U8546 (N_8546,N_8398,N_8257);
or U8547 (N_8547,N_8067,N_8182);
nand U8548 (N_8548,N_8063,N_8472);
or U8549 (N_8549,N_8354,N_8329);
xor U8550 (N_8550,N_8086,N_8401);
nor U8551 (N_8551,N_8309,N_8047);
nor U8552 (N_8552,N_8098,N_8108);
xnor U8553 (N_8553,N_8014,N_8243);
xnor U8554 (N_8554,N_8037,N_8080);
xnor U8555 (N_8555,N_8450,N_8350);
or U8556 (N_8556,N_8191,N_8247);
nand U8557 (N_8557,N_8302,N_8021);
or U8558 (N_8558,N_8205,N_8173);
nand U8559 (N_8559,N_8376,N_8226);
xnor U8560 (N_8560,N_8140,N_8289);
or U8561 (N_8561,N_8345,N_8270);
xnor U8562 (N_8562,N_8035,N_8297);
nand U8563 (N_8563,N_8141,N_8423);
nor U8564 (N_8564,N_8483,N_8118);
xnor U8565 (N_8565,N_8134,N_8197);
xnor U8566 (N_8566,N_8463,N_8120);
nand U8567 (N_8567,N_8171,N_8122);
nor U8568 (N_8568,N_8325,N_8109);
and U8569 (N_8569,N_8300,N_8018);
nor U8570 (N_8570,N_8026,N_8174);
and U8571 (N_8571,N_8322,N_8385);
nand U8572 (N_8572,N_8061,N_8105);
or U8573 (N_8573,N_8048,N_8180);
or U8574 (N_8574,N_8347,N_8365);
xor U8575 (N_8575,N_8494,N_8030);
and U8576 (N_8576,N_8402,N_8326);
nor U8577 (N_8577,N_8458,N_8276);
nand U8578 (N_8578,N_8088,N_8277);
nand U8579 (N_8579,N_8114,N_8367);
and U8580 (N_8580,N_8286,N_8042);
and U8581 (N_8581,N_8331,N_8469);
xor U8582 (N_8582,N_8471,N_8406);
and U8583 (N_8583,N_8143,N_8188);
xor U8584 (N_8584,N_8227,N_8092);
xnor U8585 (N_8585,N_8200,N_8012);
nor U8586 (N_8586,N_8217,N_8003);
nor U8587 (N_8587,N_8064,N_8203);
nand U8588 (N_8588,N_8199,N_8316);
or U8589 (N_8589,N_8124,N_8159);
and U8590 (N_8590,N_8489,N_8288);
and U8591 (N_8591,N_8475,N_8333);
nand U8592 (N_8592,N_8110,N_8267);
nor U8593 (N_8593,N_8444,N_8256);
nor U8594 (N_8594,N_8314,N_8418);
or U8595 (N_8595,N_8294,N_8057);
nor U8596 (N_8596,N_8298,N_8032);
or U8597 (N_8597,N_8485,N_8183);
nand U8598 (N_8598,N_8128,N_8295);
or U8599 (N_8599,N_8313,N_8019);
nor U8600 (N_8600,N_8465,N_8164);
or U8601 (N_8601,N_8358,N_8059);
xor U8602 (N_8602,N_8291,N_8323);
xnor U8603 (N_8603,N_8386,N_8179);
and U8604 (N_8604,N_8033,N_8410);
or U8605 (N_8605,N_8318,N_8344);
nor U8606 (N_8606,N_8498,N_8368);
nor U8607 (N_8607,N_8083,N_8349);
nand U8608 (N_8608,N_8133,N_8013);
or U8609 (N_8609,N_8434,N_8395);
nor U8610 (N_8610,N_8090,N_8155);
or U8611 (N_8611,N_8378,N_8087);
and U8612 (N_8612,N_8319,N_8055);
xor U8613 (N_8613,N_8268,N_8404);
or U8614 (N_8614,N_8010,N_8379);
and U8615 (N_8615,N_8167,N_8484);
or U8616 (N_8616,N_8422,N_8462);
xnor U8617 (N_8617,N_8269,N_8290);
nor U8618 (N_8618,N_8305,N_8015);
and U8619 (N_8619,N_8177,N_8089);
nand U8620 (N_8620,N_8467,N_8036);
or U8621 (N_8621,N_8211,N_8181);
xor U8622 (N_8622,N_8123,N_8381);
and U8623 (N_8623,N_8496,N_8020);
and U8624 (N_8624,N_8034,N_8076);
or U8625 (N_8625,N_8238,N_8207);
or U8626 (N_8626,N_8101,N_8375);
nor U8627 (N_8627,N_8360,N_8078);
nand U8628 (N_8628,N_8071,N_8066);
and U8629 (N_8629,N_8499,N_8094);
nand U8630 (N_8630,N_8366,N_8429);
and U8631 (N_8631,N_8310,N_8228);
nor U8632 (N_8632,N_8474,N_8415);
or U8633 (N_8633,N_8362,N_8144);
and U8634 (N_8634,N_8495,N_8449);
nand U8635 (N_8635,N_8165,N_8233);
nor U8636 (N_8636,N_8455,N_8005);
nor U8637 (N_8637,N_8341,N_8185);
or U8638 (N_8638,N_8491,N_8334);
nand U8639 (N_8639,N_8424,N_8258);
xor U8640 (N_8640,N_8209,N_8327);
nor U8641 (N_8641,N_8024,N_8431);
nand U8642 (N_8642,N_8028,N_8414);
nand U8643 (N_8643,N_8218,N_8396);
nand U8644 (N_8644,N_8436,N_8044);
nor U8645 (N_8645,N_8419,N_8007);
xor U8646 (N_8646,N_8482,N_8470);
nor U8647 (N_8647,N_8152,N_8204);
nand U8648 (N_8648,N_8119,N_8493);
nand U8649 (N_8649,N_8049,N_8190);
xnor U8650 (N_8650,N_8040,N_8432);
nand U8651 (N_8651,N_8158,N_8002);
or U8652 (N_8652,N_8189,N_8220);
nand U8653 (N_8653,N_8487,N_8214);
and U8654 (N_8654,N_8196,N_8184);
nor U8655 (N_8655,N_8279,N_8353);
xor U8656 (N_8656,N_8338,N_8031);
xor U8657 (N_8657,N_8212,N_8085);
or U8658 (N_8658,N_8407,N_8392);
nor U8659 (N_8659,N_8389,N_8166);
nand U8660 (N_8660,N_8438,N_8053);
xnor U8661 (N_8661,N_8320,N_8255);
xor U8662 (N_8662,N_8041,N_8104);
or U8663 (N_8663,N_8153,N_8452);
and U8664 (N_8664,N_8492,N_8045);
or U8665 (N_8665,N_8239,N_8307);
or U8666 (N_8666,N_8107,N_8001);
xnor U8667 (N_8667,N_8006,N_8052);
nand U8668 (N_8668,N_8240,N_8102);
or U8669 (N_8669,N_8273,N_8370);
xor U8670 (N_8670,N_8481,N_8303);
xor U8671 (N_8671,N_8382,N_8287);
xnor U8672 (N_8672,N_8208,N_8433);
and U8673 (N_8673,N_8121,N_8317);
and U8674 (N_8674,N_8169,N_8446);
xnor U8675 (N_8675,N_8265,N_8027);
nor U8676 (N_8676,N_8136,N_8369);
or U8677 (N_8677,N_8292,N_8112);
xnor U8678 (N_8678,N_8070,N_8077);
and U8679 (N_8679,N_8377,N_8426);
nor U8680 (N_8680,N_8116,N_8201);
or U8681 (N_8681,N_8157,N_8093);
xnor U8682 (N_8682,N_8380,N_8447);
nand U8683 (N_8683,N_8372,N_8359);
xor U8684 (N_8684,N_8457,N_8008);
nand U8685 (N_8685,N_8004,N_8068);
nand U8686 (N_8686,N_8497,N_8079);
nand U8687 (N_8687,N_8278,N_8417);
and U8688 (N_8688,N_8283,N_8357);
nand U8689 (N_8689,N_8441,N_8361);
nand U8690 (N_8690,N_8330,N_8308);
nand U8691 (N_8691,N_8213,N_8095);
xor U8692 (N_8692,N_8430,N_8249);
nor U8693 (N_8693,N_8202,N_8399);
nand U8694 (N_8694,N_8409,N_8388);
and U8695 (N_8695,N_8231,N_8160);
and U8696 (N_8696,N_8236,N_8251);
nor U8697 (N_8697,N_8225,N_8445);
nor U8698 (N_8698,N_8187,N_8373);
xor U8699 (N_8699,N_8451,N_8411);
and U8700 (N_8700,N_8056,N_8440);
and U8701 (N_8701,N_8296,N_8311);
nor U8702 (N_8702,N_8097,N_8248);
or U8703 (N_8703,N_8132,N_8082);
nor U8704 (N_8704,N_8280,N_8454);
nor U8705 (N_8705,N_8293,N_8221);
and U8706 (N_8706,N_8115,N_8403);
xor U8707 (N_8707,N_8139,N_8439);
or U8708 (N_8708,N_8252,N_8156);
and U8709 (N_8709,N_8058,N_8074);
nor U8710 (N_8710,N_8282,N_8129);
nand U8711 (N_8711,N_8352,N_8229);
and U8712 (N_8712,N_8390,N_8459);
xor U8713 (N_8713,N_8464,N_8195);
and U8714 (N_8714,N_8172,N_8264);
nand U8715 (N_8715,N_8473,N_8073);
or U8716 (N_8716,N_8384,N_8348);
nor U8717 (N_8717,N_8163,N_8259);
xnor U8718 (N_8718,N_8254,N_8304);
nor U8719 (N_8719,N_8336,N_8072);
xnor U8720 (N_8720,N_8413,N_8127);
nor U8721 (N_8721,N_8364,N_8222);
xnor U8722 (N_8722,N_8084,N_8393);
or U8723 (N_8723,N_8075,N_8235);
and U8724 (N_8724,N_8023,N_8351);
or U8725 (N_8725,N_8476,N_8246);
or U8726 (N_8726,N_8168,N_8321);
xnor U8727 (N_8727,N_8250,N_8176);
or U8728 (N_8728,N_8062,N_8117);
and U8729 (N_8729,N_8111,N_8142);
and U8730 (N_8730,N_8146,N_8193);
nand U8731 (N_8731,N_8312,N_8069);
nand U8732 (N_8732,N_8060,N_8435);
or U8733 (N_8733,N_8394,N_8383);
nor U8734 (N_8734,N_8162,N_8285);
xor U8735 (N_8735,N_8271,N_8281);
xor U8736 (N_8736,N_8224,N_8046);
nand U8737 (N_8737,N_8017,N_8151);
and U8738 (N_8738,N_8091,N_8391);
nand U8739 (N_8739,N_8161,N_8275);
or U8740 (N_8740,N_8420,N_8009);
nor U8741 (N_8741,N_8488,N_8126);
or U8742 (N_8742,N_8232,N_8374);
and U8743 (N_8743,N_8051,N_8131);
or U8744 (N_8744,N_8145,N_8081);
or U8745 (N_8745,N_8301,N_8448);
or U8746 (N_8746,N_8175,N_8335);
and U8747 (N_8747,N_8125,N_8425);
nand U8748 (N_8748,N_8219,N_8416);
or U8749 (N_8749,N_8223,N_8039);
xor U8750 (N_8750,N_8120,N_8059);
nand U8751 (N_8751,N_8109,N_8234);
nand U8752 (N_8752,N_8129,N_8009);
and U8753 (N_8753,N_8463,N_8118);
and U8754 (N_8754,N_8229,N_8297);
and U8755 (N_8755,N_8054,N_8139);
nor U8756 (N_8756,N_8137,N_8398);
or U8757 (N_8757,N_8153,N_8031);
or U8758 (N_8758,N_8077,N_8281);
or U8759 (N_8759,N_8127,N_8498);
xnor U8760 (N_8760,N_8363,N_8163);
or U8761 (N_8761,N_8067,N_8276);
nand U8762 (N_8762,N_8086,N_8372);
or U8763 (N_8763,N_8477,N_8329);
nand U8764 (N_8764,N_8039,N_8401);
or U8765 (N_8765,N_8248,N_8011);
nand U8766 (N_8766,N_8021,N_8316);
xnor U8767 (N_8767,N_8064,N_8126);
or U8768 (N_8768,N_8065,N_8459);
and U8769 (N_8769,N_8244,N_8243);
nor U8770 (N_8770,N_8365,N_8123);
nor U8771 (N_8771,N_8419,N_8147);
and U8772 (N_8772,N_8185,N_8453);
nand U8773 (N_8773,N_8087,N_8460);
xor U8774 (N_8774,N_8404,N_8452);
nand U8775 (N_8775,N_8348,N_8195);
and U8776 (N_8776,N_8087,N_8357);
nand U8777 (N_8777,N_8394,N_8136);
nor U8778 (N_8778,N_8013,N_8418);
or U8779 (N_8779,N_8430,N_8002);
or U8780 (N_8780,N_8133,N_8402);
and U8781 (N_8781,N_8498,N_8113);
or U8782 (N_8782,N_8388,N_8266);
or U8783 (N_8783,N_8203,N_8011);
and U8784 (N_8784,N_8428,N_8319);
or U8785 (N_8785,N_8119,N_8357);
and U8786 (N_8786,N_8097,N_8333);
xnor U8787 (N_8787,N_8233,N_8368);
nand U8788 (N_8788,N_8062,N_8318);
or U8789 (N_8789,N_8495,N_8288);
xnor U8790 (N_8790,N_8201,N_8300);
nor U8791 (N_8791,N_8450,N_8041);
nand U8792 (N_8792,N_8291,N_8450);
and U8793 (N_8793,N_8345,N_8171);
and U8794 (N_8794,N_8405,N_8215);
and U8795 (N_8795,N_8499,N_8072);
and U8796 (N_8796,N_8166,N_8046);
or U8797 (N_8797,N_8150,N_8326);
nor U8798 (N_8798,N_8217,N_8095);
nor U8799 (N_8799,N_8265,N_8254);
nand U8800 (N_8800,N_8355,N_8426);
nand U8801 (N_8801,N_8289,N_8342);
and U8802 (N_8802,N_8146,N_8006);
nand U8803 (N_8803,N_8236,N_8376);
nor U8804 (N_8804,N_8006,N_8083);
or U8805 (N_8805,N_8384,N_8071);
and U8806 (N_8806,N_8046,N_8180);
nor U8807 (N_8807,N_8272,N_8046);
xnor U8808 (N_8808,N_8252,N_8053);
nand U8809 (N_8809,N_8407,N_8070);
xor U8810 (N_8810,N_8412,N_8470);
xor U8811 (N_8811,N_8468,N_8446);
and U8812 (N_8812,N_8236,N_8279);
and U8813 (N_8813,N_8142,N_8268);
nor U8814 (N_8814,N_8345,N_8356);
xnor U8815 (N_8815,N_8058,N_8206);
or U8816 (N_8816,N_8144,N_8294);
nand U8817 (N_8817,N_8390,N_8204);
nor U8818 (N_8818,N_8168,N_8212);
nand U8819 (N_8819,N_8080,N_8314);
and U8820 (N_8820,N_8123,N_8310);
nand U8821 (N_8821,N_8076,N_8094);
nor U8822 (N_8822,N_8260,N_8280);
or U8823 (N_8823,N_8016,N_8372);
nor U8824 (N_8824,N_8364,N_8233);
nor U8825 (N_8825,N_8108,N_8229);
and U8826 (N_8826,N_8054,N_8329);
xor U8827 (N_8827,N_8001,N_8190);
xor U8828 (N_8828,N_8054,N_8290);
and U8829 (N_8829,N_8433,N_8147);
nand U8830 (N_8830,N_8029,N_8173);
nand U8831 (N_8831,N_8349,N_8411);
and U8832 (N_8832,N_8203,N_8247);
or U8833 (N_8833,N_8373,N_8458);
nor U8834 (N_8834,N_8178,N_8186);
and U8835 (N_8835,N_8304,N_8107);
xnor U8836 (N_8836,N_8318,N_8416);
nor U8837 (N_8837,N_8200,N_8081);
or U8838 (N_8838,N_8454,N_8162);
xnor U8839 (N_8839,N_8252,N_8181);
or U8840 (N_8840,N_8197,N_8303);
xnor U8841 (N_8841,N_8299,N_8412);
and U8842 (N_8842,N_8310,N_8115);
nand U8843 (N_8843,N_8467,N_8289);
nand U8844 (N_8844,N_8112,N_8366);
or U8845 (N_8845,N_8354,N_8216);
xor U8846 (N_8846,N_8413,N_8316);
or U8847 (N_8847,N_8475,N_8478);
nand U8848 (N_8848,N_8334,N_8323);
and U8849 (N_8849,N_8102,N_8185);
nor U8850 (N_8850,N_8307,N_8160);
xnor U8851 (N_8851,N_8178,N_8417);
nor U8852 (N_8852,N_8337,N_8331);
and U8853 (N_8853,N_8450,N_8347);
xnor U8854 (N_8854,N_8344,N_8406);
nand U8855 (N_8855,N_8269,N_8135);
or U8856 (N_8856,N_8195,N_8271);
nand U8857 (N_8857,N_8093,N_8406);
and U8858 (N_8858,N_8328,N_8416);
and U8859 (N_8859,N_8185,N_8181);
nor U8860 (N_8860,N_8137,N_8187);
nand U8861 (N_8861,N_8366,N_8420);
nand U8862 (N_8862,N_8265,N_8381);
or U8863 (N_8863,N_8226,N_8125);
or U8864 (N_8864,N_8168,N_8387);
nand U8865 (N_8865,N_8274,N_8386);
or U8866 (N_8866,N_8462,N_8416);
and U8867 (N_8867,N_8366,N_8367);
xnor U8868 (N_8868,N_8294,N_8473);
xor U8869 (N_8869,N_8292,N_8298);
nand U8870 (N_8870,N_8378,N_8367);
nor U8871 (N_8871,N_8209,N_8098);
nor U8872 (N_8872,N_8432,N_8352);
xnor U8873 (N_8873,N_8371,N_8173);
xor U8874 (N_8874,N_8184,N_8091);
xnor U8875 (N_8875,N_8177,N_8453);
and U8876 (N_8876,N_8483,N_8438);
or U8877 (N_8877,N_8039,N_8372);
or U8878 (N_8878,N_8330,N_8461);
nor U8879 (N_8879,N_8347,N_8494);
or U8880 (N_8880,N_8253,N_8401);
xor U8881 (N_8881,N_8127,N_8401);
nor U8882 (N_8882,N_8032,N_8299);
xnor U8883 (N_8883,N_8131,N_8331);
nor U8884 (N_8884,N_8369,N_8335);
nand U8885 (N_8885,N_8049,N_8394);
nand U8886 (N_8886,N_8473,N_8059);
and U8887 (N_8887,N_8289,N_8311);
and U8888 (N_8888,N_8091,N_8432);
nand U8889 (N_8889,N_8311,N_8028);
xnor U8890 (N_8890,N_8444,N_8468);
and U8891 (N_8891,N_8097,N_8271);
nor U8892 (N_8892,N_8411,N_8003);
nand U8893 (N_8893,N_8304,N_8456);
nand U8894 (N_8894,N_8216,N_8459);
xnor U8895 (N_8895,N_8221,N_8402);
nand U8896 (N_8896,N_8298,N_8042);
nor U8897 (N_8897,N_8213,N_8170);
xor U8898 (N_8898,N_8295,N_8154);
xor U8899 (N_8899,N_8312,N_8235);
nor U8900 (N_8900,N_8489,N_8333);
nand U8901 (N_8901,N_8370,N_8323);
or U8902 (N_8902,N_8039,N_8105);
nor U8903 (N_8903,N_8415,N_8069);
or U8904 (N_8904,N_8131,N_8408);
xnor U8905 (N_8905,N_8231,N_8470);
nand U8906 (N_8906,N_8207,N_8435);
and U8907 (N_8907,N_8315,N_8411);
nand U8908 (N_8908,N_8117,N_8386);
nand U8909 (N_8909,N_8123,N_8200);
or U8910 (N_8910,N_8103,N_8214);
and U8911 (N_8911,N_8283,N_8247);
or U8912 (N_8912,N_8313,N_8209);
nand U8913 (N_8913,N_8296,N_8261);
nand U8914 (N_8914,N_8345,N_8387);
xnor U8915 (N_8915,N_8359,N_8085);
nand U8916 (N_8916,N_8300,N_8009);
nor U8917 (N_8917,N_8462,N_8423);
and U8918 (N_8918,N_8093,N_8325);
and U8919 (N_8919,N_8359,N_8280);
or U8920 (N_8920,N_8438,N_8269);
or U8921 (N_8921,N_8056,N_8157);
xor U8922 (N_8922,N_8197,N_8364);
nand U8923 (N_8923,N_8085,N_8262);
xnor U8924 (N_8924,N_8062,N_8143);
xor U8925 (N_8925,N_8110,N_8392);
nand U8926 (N_8926,N_8453,N_8373);
nand U8927 (N_8927,N_8248,N_8423);
or U8928 (N_8928,N_8408,N_8220);
or U8929 (N_8929,N_8007,N_8377);
xor U8930 (N_8930,N_8119,N_8085);
nor U8931 (N_8931,N_8017,N_8363);
xnor U8932 (N_8932,N_8316,N_8353);
nor U8933 (N_8933,N_8300,N_8238);
nor U8934 (N_8934,N_8244,N_8224);
nand U8935 (N_8935,N_8289,N_8119);
or U8936 (N_8936,N_8467,N_8336);
nor U8937 (N_8937,N_8253,N_8297);
xor U8938 (N_8938,N_8339,N_8240);
nor U8939 (N_8939,N_8348,N_8176);
xnor U8940 (N_8940,N_8315,N_8431);
or U8941 (N_8941,N_8331,N_8309);
and U8942 (N_8942,N_8299,N_8357);
and U8943 (N_8943,N_8159,N_8092);
nor U8944 (N_8944,N_8290,N_8369);
or U8945 (N_8945,N_8018,N_8159);
nor U8946 (N_8946,N_8453,N_8046);
and U8947 (N_8947,N_8030,N_8454);
nand U8948 (N_8948,N_8043,N_8271);
nand U8949 (N_8949,N_8402,N_8132);
nor U8950 (N_8950,N_8017,N_8387);
and U8951 (N_8951,N_8115,N_8096);
xnor U8952 (N_8952,N_8398,N_8102);
nor U8953 (N_8953,N_8280,N_8147);
nand U8954 (N_8954,N_8049,N_8029);
and U8955 (N_8955,N_8467,N_8026);
or U8956 (N_8956,N_8295,N_8301);
nor U8957 (N_8957,N_8383,N_8022);
nor U8958 (N_8958,N_8178,N_8366);
or U8959 (N_8959,N_8378,N_8470);
nor U8960 (N_8960,N_8443,N_8475);
or U8961 (N_8961,N_8293,N_8135);
xor U8962 (N_8962,N_8204,N_8178);
xor U8963 (N_8963,N_8339,N_8027);
nand U8964 (N_8964,N_8276,N_8151);
xor U8965 (N_8965,N_8496,N_8439);
nand U8966 (N_8966,N_8264,N_8001);
nor U8967 (N_8967,N_8411,N_8374);
nor U8968 (N_8968,N_8351,N_8079);
or U8969 (N_8969,N_8034,N_8250);
or U8970 (N_8970,N_8065,N_8496);
and U8971 (N_8971,N_8057,N_8034);
xor U8972 (N_8972,N_8333,N_8065);
nor U8973 (N_8973,N_8200,N_8205);
or U8974 (N_8974,N_8116,N_8242);
xor U8975 (N_8975,N_8269,N_8277);
xnor U8976 (N_8976,N_8154,N_8241);
nor U8977 (N_8977,N_8047,N_8208);
nand U8978 (N_8978,N_8208,N_8307);
xnor U8979 (N_8979,N_8083,N_8413);
xor U8980 (N_8980,N_8056,N_8038);
or U8981 (N_8981,N_8032,N_8389);
and U8982 (N_8982,N_8009,N_8379);
or U8983 (N_8983,N_8459,N_8152);
and U8984 (N_8984,N_8368,N_8206);
or U8985 (N_8985,N_8167,N_8187);
and U8986 (N_8986,N_8069,N_8201);
or U8987 (N_8987,N_8397,N_8355);
nor U8988 (N_8988,N_8155,N_8304);
or U8989 (N_8989,N_8453,N_8347);
and U8990 (N_8990,N_8318,N_8341);
nand U8991 (N_8991,N_8245,N_8346);
xor U8992 (N_8992,N_8050,N_8229);
and U8993 (N_8993,N_8223,N_8033);
or U8994 (N_8994,N_8214,N_8087);
or U8995 (N_8995,N_8270,N_8115);
and U8996 (N_8996,N_8326,N_8219);
xnor U8997 (N_8997,N_8105,N_8187);
nor U8998 (N_8998,N_8058,N_8338);
xnor U8999 (N_8999,N_8498,N_8323);
xor U9000 (N_9000,N_8860,N_8721);
and U9001 (N_9001,N_8900,N_8965);
and U9002 (N_9002,N_8799,N_8573);
or U9003 (N_9003,N_8856,N_8703);
xor U9004 (N_9004,N_8607,N_8908);
nand U9005 (N_9005,N_8613,N_8976);
xnor U9006 (N_9006,N_8905,N_8540);
xnor U9007 (N_9007,N_8830,N_8763);
nand U9008 (N_9008,N_8864,N_8862);
and U9009 (N_9009,N_8876,N_8816);
nor U9010 (N_9010,N_8624,N_8601);
xnor U9011 (N_9011,N_8632,N_8514);
nor U9012 (N_9012,N_8815,N_8519);
xor U9013 (N_9013,N_8853,N_8887);
xnor U9014 (N_9014,N_8738,N_8604);
nand U9015 (N_9015,N_8814,N_8709);
xor U9016 (N_9016,N_8777,N_8733);
nor U9017 (N_9017,N_8962,N_8953);
nor U9018 (N_9018,N_8509,N_8500);
or U9019 (N_9019,N_8930,N_8707);
xnor U9020 (N_9020,N_8701,N_8880);
or U9021 (N_9021,N_8669,N_8939);
or U9022 (N_9022,N_8575,N_8787);
nand U9023 (N_9023,N_8751,N_8995);
nor U9024 (N_9024,N_8524,N_8626);
or U9025 (N_9025,N_8505,N_8739);
and U9026 (N_9026,N_8837,N_8821);
and U9027 (N_9027,N_8757,N_8768);
or U9028 (N_9028,N_8541,N_8857);
and U9029 (N_9029,N_8903,N_8952);
nor U9030 (N_9030,N_8960,N_8620);
and U9031 (N_9031,N_8841,N_8502);
or U9032 (N_9032,N_8752,N_8531);
nand U9033 (N_9033,N_8718,N_8817);
or U9034 (N_9034,N_8973,N_8801);
nor U9035 (N_9035,N_8746,N_8537);
nand U9036 (N_9036,N_8772,N_8981);
and U9037 (N_9037,N_8923,N_8726);
xor U9038 (N_9038,N_8614,N_8569);
and U9039 (N_9039,N_8641,N_8854);
xor U9040 (N_9040,N_8650,N_8566);
xor U9041 (N_9041,N_8651,N_8679);
xnor U9042 (N_9042,N_8518,N_8783);
xor U9043 (N_9043,N_8542,N_8647);
and U9044 (N_9044,N_8728,N_8873);
xnor U9045 (N_9045,N_8562,N_8686);
nor U9046 (N_9046,N_8661,N_8936);
xor U9047 (N_9047,N_8740,N_8512);
xor U9048 (N_9048,N_8587,N_8576);
nand U9049 (N_9049,N_8670,N_8565);
nand U9050 (N_9050,N_8530,N_8889);
and U9051 (N_9051,N_8517,N_8684);
xor U9052 (N_9052,N_8767,N_8780);
nor U9053 (N_9053,N_8700,N_8765);
and U9054 (N_9054,N_8781,N_8720);
and U9055 (N_9055,N_8805,N_8828);
nand U9056 (N_9056,N_8547,N_8695);
xor U9057 (N_9057,N_8997,N_8957);
nor U9058 (N_9058,N_8527,N_8634);
nor U9059 (N_9059,N_8636,N_8774);
xor U9060 (N_9060,N_8773,N_8642);
nor U9061 (N_9061,N_8983,N_8653);
nor U9062 (N_9062,N_8605,N_8513);
and U9063 (N_9063,N_8741,N_8769);
xnor U9064 (N_9064,N_8825,N_8748);
and U9065 (N_9065,N_8858,N_8951);
nor U9066 (N_9066,N_8802,N_8894);
or U9067 (N_9067,N_8663,N_8849);
and U9068 (N_9068,N_8550,N_8994);
nand U9069 (N_9069,N_8646,N_8680);
nand U9070 (N_9070,N_8657,N_8682);
or U9071 (N_9071,N_8567,N_8975);
nor U9072 (N_9072,N_8929,N_8598);
xor U9073 (N_9073,N_8941,N_8836);
nand U9074 (N_9074,N_8938,N_8654);
nor U9075 (N_9075,N_8879,N_8611);
nand U9076 (N_9076,N_8789,N_8696);
nor U9077 (N_9077,N_8883,N_8870);
nand U9078 (N_9078,N_8974,N_8667);
nand U9079 (N_9079,N_8592,N_8711);
nand U9080 (N_9080,N_8539,N_8599);
nand U9081 (N_9081,N_8621,N_8627);
xnor U9082 (N_9082,N_8762,N_8984);
nor U9083 (N_9083,N_8600,N_8612);
and U9084 (N_9084,N_8675,N_8998);
nor U9085 (N_9085,N_8618,N_8940);
nand U9086 (N_9086,N_8737,N_8759);
xor U9087 (N_9087,N_8919,N_8788);
or U9088 (N_9088,N_8779,N_8943);
nand U9089 (N_9089,N_8723,N_8866);
or U9090 (N_9090,N_8840,N_8590);
xor U9091 (N_9091,N_8988,N_8552);
nand U9092 (N_9092,N_8888,N_8526);
nor U9093 (N_9093,N_8949,N_8616);
xnor U9094 (N_9094,N_8784,N_8557);
nor U9095 (N_9095,N_8520,N_8843);
and U9096 (N_9096,N_8735,N_8833);
and U9097 (N_9097,N_8672,N_8794);
nor U9098 (N_9098,N_8898,N_8503);
and U9099 (N_9099,N_8555,N_8570);
xnor U9100 (N_9100,N_8778,N_8515);
and U9101 (N_9101,N_8832,N_8609);
xor U9102 (N_9102,N_8764,N_8822);
nand U9103 (N_9103,N_8591,N_8804);
xnor U9104 (N_9104,N_8619,N_8807);
xnor U9105 (N_9105,N_8851,N_8553);
or U9106 (N_9106,N_8610,N_8544);
or U9107 (N_9107,N_8648,N_8705);
xor U9108 (N_9108,N_8945,N_8715);
nor U9109 (N_9109,N_8831,N_8872);
xor U9110 (N_9110,N_8572,N_8508);
and U9111 (N_9111,N_8538,N_8596);
or U9112 (N_9112,N_8734,N_8956);
or U9113 (N_9113,N_8745,N_8895);
xor U9114 (N_9114,N_8980,N_8834);
and U9115 (N_9115,N_8885,N_8676);
and U9116 (N_9116,N_8645,N_8693);
and U9117 (N_9117,N_8971,N_8913);
or U9118 (N_9118,N_8820,N_8637);
nor U9119 (N_9119,N_8685,N_8969);
nand U9120 (N_9120,N_8691,N_8776);
nand U9121 (N_9121,N_8589,N_8692);
and U9122 (N_9122,N_8623,N_8747);
xor U9123 (N_9123,N_8568,N_8838);
xor U9124 (N_9124,N_8749,N_8925);
nand U9125 (N_9125,N_8800,N_8533);
and U9126 (N_9126,N_8934,N_8933);
nand U9127 (N_9127,N_8717,N_8617);
nor U9128 (N_9128,N_8795,N_8699);
nor U9129 (N_9129,N_8855,N_8668);
and U9130 (N_9130,N_8683,N_8716);
xor U9131 (N_9131,N_8558,N_8595);
nand U9132 (N_9132,N_8847,N_8593);
xnor U9133 (N_9133,N_8602,N_8797);
nor U9134 (N_9134,N_8608,N_8775);
or U9135 (N_9135,N_8631,N_8659);
nand U9136 (N_9136,N_8506,N_8761);
and U9137 (N_9137,N_8875,N_8755);
xor U9138 (N_9138,N_8708,N_8750);
and U9139 (N_9139,N_8697,N_8852);
xnor U9140 (N_9140,N_8766,N_8916);
or U9141 (N_9141,N_8990,N_8977);
and U9142 (N_9142,N_8991,N_8992);
and U9143 (N_9143,N_8574,N_8829);
and U9144 (N_9144,N_8730,N_8986);
xnor U9145 (N_9145,N_8525,N_8877);
nand U9146 (N_9146,N_8850,N_8603);
nand U9147 (N_9147,N_8656,N_8736);
nand U9148 (N_9148,N_8897,N_8742);
or U9149 (N_9149,N_8551,N_8674);
and U9150 (N_9150,N_8694,N_8996);
or U9151 (N_9151,N_8665,N_8982);
or U9152 (N_9152,N_8978,N_8606);
and U9153 (N_9153,N_8811,N_8989);
nand U9154 (N_9154,N_8944,N_8630);
and U9155 (N_9155,N_8867,N_8993);
nand U9156 (N_9156,N_8655,N_8892);
xor U9157 (N_9157,N_8678,N_8891);
xnor U9158 (N_9158,N_8688,N_8523);
nor U9159 (N_9159,N_8810,N_8724);
nor U9160 (N_9160,N_8536,N_8844);
and U9161 (N_9161,N_8871,N_8644);
nand U9162 (N_9162,N_8863,N_8842);
or U9163 (N_9163,N_8690,N_8658);
or U9164 (N_9164,N_8921,N_8543);
or U9165 (N_9165,N_8588,N_8535);
nor U9166 (N_9166,N_8987,N_8947);
or U9167 (N_9167,N_8687,N_8958);
nand U9168 (N_9168,N_8886,N_8760);
and U9169 (N_9169,N_8564,N_8578);
nor U9170 (N_9170,N_8970,N_8639);
and U9171 (N_9171,N_8652,N_8791);
nor U9172 (N_9172,N_8560,N_8706);
nand U9173 (N_9173,N_8926,N_8985);
xor U9174 (N_9174,N_8964,N_8848);
nand U9175 (N_9175,N_8556,N_8909);
and U9176 (N_9176,N_8979,N_8999);
xnor U9177 (N_9177,N_8809,N_8677);
xor U9178 (N_9178,N_8731,N_8704);
xor U9179 (N_9179,N_8580,N_8702);
nand U9180 (N_9180,N_8950,N_8722);
and U9181 (N_9181,N_8671,N_8826);
or U9182 (N_9182,N_8754,N_8615);
and U9183 (N_9183,N_8827,N_8968);
xnor U9184 (N_9184,N_8664,N_8920);
nand U9185 (N_9185,N_8744,N_8666);
xnor U9186 (N_9186,N_8845,N_8579);
and U9187 (N_9187,N_8638,N_8522);
nand U9188 (N_9188,N_8963,N_8549);
and U9189 (N_9189,N_8689,N_8725);
and U9190 (N_9190,N_8922,N_8545);
nand U9191 (N_9191,N_8582,N_8790);
xor U9192 (N_9192,N_8823,N_8594);
xnor U9193 (N_9193,N_8961,N_8899);
xor U9194 (N_9194,N_8782,N_8714);
nand U9195 (N_9195,N_8554,N_8559);
nand U9196 (N_9196,N_8698,N_8884);
nand U9197 (N_9197,N_8597,N_8803);
nand U9198 (N_9198,N_8808,N_8946);
and U9199 (N_9199,N_8902,N_8532);
or U9200 (N_9200,N_8918,N_8625);
nand U9201 (N_9201,N_8901,N_8510);
or U9202 (N_9202,N_8758,N_8924);
xnor U9203 (N_9203,N_8910,N_8622);
or U9204 (N_9204,N_8511,N_8874);
xor U9205 (N_9205,N_8629,N_8548);
and U9206 (N_9206,N_8584,N_8907);
nor U9207 (N_9207,N_8640,N_8914);
xor U9208 (N_9208,N_8585,N_8660);
xor U9209 (N_9209,N_8896,N_8959);
nand U9210 (N_9210,N_8915,N_8534);
nand U9211 (N_9211,N_8906,N_8927);
xor U9212 (N_9212,N_8528,N_8729);
nor U9213 (N_9213,N_8516,N_8793);
xnor U9214 (N_9214,N_8966,N_8846);
or U9215 (N_9215,N_8812,N_8882);
or U9216 (N_9216,N_8948,N_8917);
or U9217 (N_9217,N_8861,N_8628);
nor U9218 (N_9218,N_8865,N_8643);
and U9219 (N_9219,N_8571,N_8911);
nand U9220 (N_9220,N_8662,N_8868);
and U9221 (N_9221,N_8635,N_8546);
or U9222 (N_9222,N_8818,N_8869);
nor U9223 (N_9223,N_8521,N_8792);
nor U9224 (N_9224,N_8785,N_8786);
xor U9225 (N_9225,N_8942,N_8932);
or U9226 (N_9226,N_8935,N_8713);
nand U9227 (N_9227,N_8904,N_8753);
xnor U9228 (N_9228,N_8756,N_8881);
nand U9229 (N_9229,N_8743,N_8732);
xnor U9230 (N_9230,N_8681,N_8586);
nor U9231 (N_9231,N_8824,N_8563);
and U9232 (N_9232,N_8937,N_8727);
xnor U9233 (N_9233,N_8955,N_8710);
and U9234 (N_9234,N_8806,N_8581);
xnor U9235 (N_9235,N_8859,N_8931);
nor U9236 (N_9236,N_8912,N_8673);
or U9237 (N_9237,N_8813,N_8504);
nand U9238 (N_9238,N_8529,N_8501);
and U9239 (N_9239,N_8633,N_8583);
or U9240 (N_9240,N_8719,N_8796);
nand U9241 (N_9241,N_8798,N_8878);
nand U9242 (N_9242,N_8771,N_8577);
and U9243 (N_9243,N_8972,N_8890);
xnor U9244 (N_9244,N_8819,N_8649);
or U9245 (N_9245,N_8712,N_8561);
xnor U9246 (N_9246,N_8893,N_8954);
xnor U9247 (N_9247,N_8928,N_8770);
xnor U9248 (N_9248,N_8507,N_8835);
nand U9249 (N_9249,N_8967,N_8839);
and U9250 (N_9250,N_8948,N_8786);
nand U9251 (N_9251,N_8784,N_8733);
and U9252 (N_9252,N_8811,N_8814);
nor U9253 (N_9253,N_8768,N_8639);
or U9254 (N_9254,N_8781,N_8899);
nand U9255 (N_9255,N_8727,N_8571);
xnor U9256 (N_9256,N_8918,N_8761);
nand U9257 (N_9257,N_8502,N_8939);
or U9258 (N_9258,N_8635,N_8913);
or U9259 (N_9259,N_8825,N_8563);
nand U9260 (N_9260,N_8582,N_8868);
and U9261 (N_9261,N_8776,N_8503);
and U9262 (N_9262,N_8947,N_8893);
xor U9263 (N_9263,N_8710,N_8630);
xor U9264 (N_9264,N_8564,N_8681);
and U9265 (N_9265,N_8954,N_8607);
or U9266 (N_9266,N_8664,N_8598);
or U9267 (N_9267,N_8973,N_8761);
nor U9268 (N_9268,N_8565,N_8924);
nand U9269 (N_9269,N_8810,N_8588);
nor U9270 (N_9270,N_8683,N_8807);
nor U9271 (N_9271,N_8949,N_8635);
nor U9272 (N_9272,N_8655,N_8707);
xnor U9273 (N_9273,N_8936,N_8762);
and U9274 (N_9274,N_8881,N_8966);
or U9275 (N_9275,N_8607,N_8969);
or U9276 (N_9276,N_8833,N_8795);
and U9277 (N_9277,N_8796,N_8569);
and U9278 (N_9278,N_8996,N_8541);
nand U9279 (N_9279,N_8751,N_8845);
nand U9280 (N_9280,N_8620,N_8539);
nand U9281 (N_9281,N_8651,N_8670);
xor U9282 (N_9282,N_8917,N_8765);
and U9283 (N_9283,N_8635,N_8958);
xnor U9284 (N_9284,N_8975,N_8972);
nand U9285 (N_9285,N_8757,N_8840);
xnor U9286 (N_9286,N_8515,N_8790);
nand U9287 (N_9287,N_8522,N_8775);
and U9288 (N_9288,N_8779,N_8829);
xnor U9289 (N_9289,N_8656,N_8647);
xnor U9290 (N_9290,N_8656,N_8563);
or U9291 (N_9291,N_8975,N_8933);
nand U9292 (N_9292,N_8927,N_8615);
and U9293 (N_9293,N_8817,N_8569);
nand U9294 (N_9294,N_8831,N_8747);
or U9295 (N_9295,N_8870,N_8731);
nor U9296 (N_9296,N_8671,N_8591);
and U9297 (N_9297,N_8940,N_8906);
and U9298 (N_9298,N_8855,N_8894);
nor U9299 (N_9299,N_8921,N_8957);
xnor U9300 (N_9300,N_8963,N_8790);
and U9301 (N_9301,N_8777,N_8862);
and U9302 (N_9302,N_8883,N_8963);
and U9303 (N_9303,N_8606,N_8663);
nor U9304 (N_9304,N_8850,N_8890);
or U9305 (N_9305,N_8784,N_8519);
nor U9306 (N_9306,N_8817,N_8794);
or U9307 (N_9307,N_8841,N_8571);
and U9308 (N_9308,N_8891,N_8818);
xnor U9309 (N_9309,N_8783,N_8762);
or U9310 (N_9310,N_8803,N_8827);
and U9311 (N_9311,N_8717,N_8995);
nor U9312 (N_9312,N_8950,N_8995);
nor U9313 (N_9313,N_8609,N_8988);
nor U9314 (N_9314,N_8813,N_8952);
or U9315 (N_9315,N_8630,N_8589);
nor U9316 (N_9316,N_8555,N_8681);
or U9317 (N_9317,N_8983,N_8984);
and U9318 (N_9318,N_8655,N_8516);
nor U9319 (N_9319,N_8575,N_8747);
nand U9320 (N_9320,N_8651,N_8821);
nor U9321 (N_9321,N_8681,N_8615);
and U9322 (N_9322,N_8563,N_8807);
or U9323 (N_9323,N_8855,N_8879);
or U9324 (N_9324,N_8880,N_8856);
nand U9325 (N_9325,N_8846,N_8738);
nand U9326 (N_9326,N_8999,N_8909);
or U9327 (N_9327,N_8715,N_8890);
or U9328 (N_9328,N_8508,N_8606);
nor U9329 (N_9329,N_8913,N_8664);
and U9330 (N_9330,N_8989,N_8618);
xnor U9331 (N_9331,N_8698,N_8625);
xnor U9332 (N_9332,N_8707,N_8532);
xor U9333 (N_9333,N_8980,N_8869);
nand U9334 (N_9334,N_8632,N_8858);
and U9335 (N_9335,N_8949,N_8803);
or U9336 (N_9336,N_8884,N_8739);
and U9337 (N_9337,N_8988,N_8531);
nor U9338 (N_9338,N_8802,N_8917);
nand U9339 (N_9339,N_8877,N_8747);
or U9340 (N_9340,N_8868,N_8791);
xor U9341 (N_9341,N_8892,N_8710);
nor U9342 (N_9342,N_8949,N_8668);
nand U9343 (N_9343,N_8886,N_8515);
or U9344 (N_9344,N_8514,N_8566);
nand U9345 (N_9345,N_8544,N_8904);
nand U9346 (N_9346,N_8817,N_8676);
xnor U9347 (N_9347,N_8962,N_8731);
xnor U9348 (N_9348,N_8735,N_8563);
nor U9349 (N_9349,N_8933,N_8514);
nor U9350 (N_9350,N_8975,N_8834);
xnor U9351 (N_9351,N_8675,N_8933);
and U9352 (N_9352,N_8655,N_8955);
and U9353 (N_9353,N_8804,N_8780);
xor U9354 (N_9354,N_8588,N_8943);
or U9355 (N_9355,N_8915,N_8537);
xnor U9356 (N_9356,N_8939,N_8653);
and U9357 (N_9357,N_8697,N_8747);
nor U9358 (N_9358,N_8558,N_8913);
xnor U9359 (N_9359,N_8678,N_8663);
or U9360 (N_9360,N_8946,N_8763);
xor U9361 (N_9361,N_8793,N_8521);
and U9362 (N_9362,N_8608,N_8742);
xor U9363 (N_9363,N_8881,N_8784);
and U9364 (N_9364,N_8526,N_8814);
nand U9365 (N_9365,N_8820,N_8947);
nand U9366 (N_9366,N_8788,N_8861);
and U9367 (N_9367,N_8523,N_8631);
xnor U9368 (N_9368,N_8846,N_8606);
or U9369 (N_9369,N_8596,N_8513);
or U9370 (N_9370,N_8796,N_8654);
nand U9371 (N_9371,N_8754,N_8749);
nor U9372 (N_9372,N_8601,N_8820);
nor U9373 (N_9373,N_8671,N_8906);
xor U9374 (N_9374,N_8910,N_8517);
and U9375 (N_9375,N_8960,N_8704);
and U9376 (N_9376,N_8552,N_8951);
and U9377 (N_9377,N_8838,N_8805);
and U9378 (N_9378,N_8703,N_8584);
xor U9379 (N_9379,N_8904,N_8932);
xnor U9380 (N_9380,N_8789,N_8798);
nand U9381 (N_9381,N_8761,N_8999);
or U9382 (N_9382,N_8907,N_8952);
xor U9383 (N_9383,N_8594,N_8724);
nand U9384 (N_9384,N_8525,N_8752);
or U9385 (N_9385,N_8768,N_8676);
xnor U9386 (N_9386,N_8892,N_8998);
nor U9387 (N_9387,N_8680,N_8773);
nor U9388 (N_9388,N_8839,N_8598);
nor U9389 (N_9389,N_8955,N_8532);
or U9390 (N_9390,N_8878,N_8875);
and U9391 (N_9391,N_8864,N_8850);
nor U9392 (N_9392,N_8818,N_8706);
nor U9393 (N_9393,N_8912,N_8582);
xor U9394 (N_9394,N_8719,N_8662);
or U9395 (N_9395,N_8586,N_8851);
xor U9396 (N_9396,N_8599,N_8622);
nand U9397 (N_9397,N_8900,N_8630);
nand U9398 (N_9398,N_8674,N_8639);
nand U9399 (N_9399,N_8648,N_8938);
xnor U9400 (N_9400,N_8829,N_8971);
nand U9401 (N_9401,N_8672,N_8834);
or U9402 (N_9402,N_8504,N_8729);
nor U9403 (N_9403,N_8877,N_8928);
nand U9404 (N_9404,N_8863,N_8548);
and U9405 (N_9405,N_8677,N_8837);
and U9406 (N_9406,N_8712,N_8641);
and U9407 (N_9407,N_8685,N_8688);
or U9408 (N_9408,N_8674,N_8515);
nand U9409 (N_9409,N_8910,N_8690);
nor U9410 (N_9410,N_8809,N_8591);
nor U9411 (N_9411,N_8651,N_8515);
nand U9412 (N_9412,N_8501,N_8852);
nor U9413 (N_9413,N_8770,N_8811);
and U9414 (N_9414,N_8826,N_8760);
or U9415 (N_9415,N_8598,N_8943);
xnor U9416 (N_9416,N_8537,N_8800);
xor U9417 (N_9417,N_8825,N_8610);
and U9418 (N_9418,N_8895,N_8776);
and U9419 (N_9419,N_8761,N_8849);
or U9420 (N_9420,N_8786,N_8797);
nand U9421 (N_9421,N_8749,N_8676);
and U9422 (N_9422,N_8915,N_8685);
xor U9423 (N_9423,N_8897,N_8978);
and U9424 (N_9424,N_8866,N_8520);
and U9425 (N_9425,N_8731,N_8588);
or U9426 (N_9426,N_8939,N_8817);
or U9427 (N_9427,N_8553,N_8587);
or U9428 (N_9428,N_8914,N_8810);
nand U9429 (N_9429,N_8551,N_8582);
nand U9430 (N_9430,N_8593,N_8568);
or U9431 (N_9431,N_8718,N_8516);
xor U9432 (N_9432,N_8977,N_8967);
nor U9433 (N_9433,N_8848,N_8669);
or U9434 (N_9434,N_8861,N_8958);
nand U9435 (N_9435,N_8841,N_8998);
nor U9436 (N_9436,N_8918,N_8757);
and U9437 (N_9437,N_8692,N_8507);
and U9438 (N_9438,N_8887,N_8843);
or U9439 (N_9439,N_8931,N_8892);
nand U9440 (N_9440,N_8592,N_8973);
or U9441 (N_9441,N_8767,N_8517);
or U9442 (N_9442,N_8726,N_8859);
xor U9443 (N_9443,N_8920,N_8631);
xnor U9444 (N_9444,N_8659,N_8853);
nand U9445 (N_9445,N_8572,N_8846);
xor U9446 (N_9446,N_8992,N_8722);
nand U9447 (N_9447,N_8593,N_8741);
nand U9448 (N_9448,N_8591,N_8865);
nand U9449 (N_9449,N_8947,N_8589);
xnor U9450 (N_9450,N_8602,N_8550);
nor U9451 (N_9451,N_8926,N_8971);
or U9452 (N_9452,N_8764,N_8556);
and U9453 (N_9453,N_8581,N_8615);
and U9454 (N_9454,N_8561,N_8507);
or U9455 (N_9455,N_8681,N_8659);
or U9456 (N_9456,N_8788,N_8778);
and U9457 (N_9457,N_8664,N_8503);
nor U9458 (N_9458,N_8598,N_8722);
and U9459 (N_9459,N_8577,N_8705);
or U9460 (N_9460,N_8883,N_8874);
and U9461 (N_9461,N_8749,N_8736);
xor U9462 (N_9462,N_8651,N_8537);
nor U9463 (N_9463,N_8808,N_8611);
and U9464 (N_9464,N_8901,N_8637);
nand U9465 (N_9465,N_8815,N_8792);
xor U9466 (N_9466,N_8755,N_8995);
xor U9467 (N_9467,N_8675,N_8532);
nand U9468 (N_9468,N_8957,N_8999);
xnor U9469 (N_9469,N_8668,N_8718);
xnor U9470 (N_9470,N_8630,N_8919);
and U9471 (N_9471,N_8559,N_8771);
xnor U9472 (N_9472,N_8980,N_8833);
nor U9473 (N_9473,N_8669,N_8777);
and U9474 (N_9474,N_8629,N_8669);
nor U9475 (N_9475,N_8764,N_8754);
xor U9476 (N_9476,N_8960,N_8861);
nand U9477 (N_9477,N_8678,N_8928);
and U9478 (N_9478,N_8658,N_8992);
xnor U9479 (N_9479,N_8974,N_8914);
or U9480 (N_9480,N_8678,N_8672);
xor U9481 (N_9481,N_8818,N_8899);
nor U9482 (N_9482,N_8560,N_8566);
xnor U9483 (N_9483,N_8580,N_8944);
or U9484 (N_9484,N_8611,N_8680);
nor U9485 (N_9485,N_8508,N_8741);
and U9486 (N_9486,N_8717,N_8619);
and U9487 (N_9487,N_8943,N_8762);
xor U9488 (N_9488,N_8507,N_8628);
xnor U9489 (N_9489,N_8508,N_8694);
nand U9490 (N_9490,N_8599,N_8699);
and U9491 (N_9491,N_8964,N_8973);
xnor U9492 (N_9492,N_8731,N_8692);
and U9493 (N_9493,N_8566,N_8616);
xnor U9494 (N_9494,N_8856,N_8622);
and U9495 (N_9495,N_8829,N_8973);
nand U9496 (N_9496,N_8767,N_8543);
nand U9497 (N_9497,N_8998,N_8802);
nor U9498 (N_9498,N_8887,N_8836);
and U9499 (N_9499,N_8603,N_8562);
nand U9500 (N_9500,N_9482,N_9448);
xnor U9501 (N_9501,N_9041,N_9086);
or U9502 (N_9502,N_9020,N_9431);
xor U9503 (N_9503,N_9375,N_9472);
xor U9504 (N_9504,N_9009,N_9222);
or U9505 (N_9505,N_9475,N_9489);
nor U9506 (N_9506,N_9125,N_9220);
and U9507 (N_9507,N_9329,N_9164);
nor U9508 (N_9508,N_9387,N_9171);
and U9509 (N_9509,N_9066,N_9207);
nor U9510 (N_9510,N_9002,N_9240);
nor U9511 (N_9511,N_9301,N_9403);
and U9512 (N_9512,N_9254,N_9025);
nand U9513 (N_9513,N_9186,N_9257);
nor U9514 (N_9514,N_9130,N_9269);
xnor U9515 (N_9515,N_9335,N_9298);
nor U9516 (N_9516,N_9366,N_9132);
nor U9517 (N_9517,N_9296,N_9261);
and U9518 (N_9518,N_9076,N_9116);
nor U9519 (N_9519,N_9377,N_9305);
xnor U9520 (N_9520,N_9189,N_9121);
nor U9521 (N_9521,N_9445,N_9050);
xor U9522 (N_9522,N_9049,N_9229);
or U9523 (N_9523,N_9061,N_9182);
or U9524 (N_9524,N_9043,N_9058);
xor U9525 (N_9525,N_9036,N_9427);
or U9526 (N_9526,N_9200,N_9410);
or U9527 (N_9527,N_9462,N_9409);
xnor U9528 (N_9528,N_9317,N_9196);
xnor U9529 (N_9529,N_9215,N_9102);
nor U9530 (N_9530,N_9468,N_9374);
or U9531 (N_9531,N_9415,N_9339);
or U9532 (N_9532,N_9178,N_9242);
or U9533 (N_9533,N_9423,N_9424);
xnor U9534 (N_9534,N_9350,N_9248);
nor U9535 (N_9535,N_9413,N_9358);
nor U9536 (N_9536,N_9490,N_9247);
nand U9537 (N_9537,N_9223,N_9465);
nor U9538 (N_9538,N_9162,N_9143);
nor U9539 (N_9539,N_9059,N_9080);
or U9540 (N_9540,N_9429,N_9372);
nand U9541 (N_9541,N_9297,N_9003);
and U9542 (N_9542,N_9417,N_9053);
nand U9543 (N_9543,N_9253,N_9068);
nor U9544 (N_9544,N_9149,N_9163);
xor U9545 (N_9545,N_9219,N_9213);
or U9546 (N_9546,N_9395,N_9360);
nor U9547 (N_9547,N_9195,N_9477);
xor U9548 (N_9548,N_9359,N_9141);
xnor U9549 (N_9549,N_9302,N_9032);
xnor U9550 (N_9550,N_9176,N_9106);
xnor U9551 (N_9551,N_9451,N_9113);
and U9552 (N_9552,N_9264,N_9390);
nor U9553 (N_9553,N_9293,N_9040);
and U9554 (N_9554,N_9190,N_9150);
xnor U9555 (N_9555,N_9383,N_9496);
nand U9556 (N_9556,N_9478,N_9031);
nor U9557 (N_9557,N_9396,N_9225);
nor U9558 (N_9558,N_9291,N_9203);
nand U9559 (N_9559,N_9382,N_9405);
and U9560 (N_9560,N_9425,N_9000);
nand U9561 (N_9561,N_9193,N_9142);
and U9562 (N_9562,N_9385,N_9259);
nand U9563 (N_9563,N_9100,N_9498);
nor U9564 (N_9564,N_9288,N_9202);
and U9565 (N_9565,N_9124,N_9140);
and U9566 (N_9566,N_9093,N_9177);
nand U9567 (N_9567,N_9233,N_9211);
xor U9568 (N_9568,N_9401,N_9243);
nand U9569 (N_9569,N_9273,N_9354);
and U9570 (N_9570,N_9459,N_9318);
and U9571 (N_9571,N_9241,N_9098);
nor U9572 (N_9572,N_9493,N_9333);
and U9573 (N_9573,N_9416,N_9208);
nor U9574 (N_9574,N_9268,N_9173);
and U9575 (N_9575,N_9275,N_9316);
xor U9576 (N_9576,N_9037,N_9338);
and U9577 (N_9577,N_9436,N_9327);
nor U9578 (N_9578,N_9393,N_9309);
or U9579 (N_9579,N_9353,N_9276);
xor U9580 (N_9580,N_9146,N_9007);
or U9581 (N_9581,N_9485,N_9209);
or U9582 (N_9582,N_9251,N_9394);
xor U9583 (N_9583,N_9089,N_9038);
nor U9584 (N_9584,N_9079,N_9055);
or U9585 (N_9585,N_9008,N_9384);
xor U9586 (N_9586,N_9446,N_9073);
nor U9587 (N_9587,N_9016,N_9322);
and U9588 (N_9588,N_9012,N_9308);
or U9589 (N_9589,N_9197,N_9105);
nand U9590 (N_9590,N_9342,N_9029);
or U9591 (N_9591,N_9289,N_9330);
or U9592 (N_9592,N_9062,N_9454);
and U9593 (N_9593,N_9152,N_9054);
nand U9594 (N_9594,N_9277,N_9048);
or U9595 (N_9595,N_9167,N_9274);
nand U9596 (N_9596,N_9314,N_9456);
and U9597 (N_9597,N_9255,N_9123);
nand U9598 (N_9598,N_9292,N_9306);
and U9599 (N_9599,N_9450,N_9075);
nand U9600 (N_9600,N_9487,N_9001);
xnor U9601 (N_9601,N_9328,N_9379);
nor U9602 (N_9602,N_9045,N_9434);
nor U9603 (N_9603,N_9381,N_9131);
and U9604 (N_9604,N_9422,N_9249);
xnor U9605 (N_9605,N_9426,N_9161);
xnor U9606 (N_9606,N_9380,N_9299);
nand U9607 (N_9607,N_9082,N_9227);
xor U9608 (N_9608,N_9090,N_9217);
nor U9609 (N_9609,N_9440,N_9072);
nor U9610 (N_9610,N_9170,N_9226);
or U9611 (N_9611,N_9421,N_9185);
nand U9612 (N_9612,N_9109,N_9165);
or U9613 (N_9613,N_9461,N_9244);
xnor U9614 (N_9614,N_9119,N_9087);
nor U9615 (N_9615,N_9096,N_9432);
nand U9616 (N_9616,N_9480,N_9024);
xnor U9617 (N_9617,N_9371,N_9057);
nand U9618 (N_9618,N_9237,N_9260);
nor U9619 (N_9619,N_9285,N_9144);
and U9620 (N_9620,N_9046,N_9136);
xor U9621 (N_9621,N_9444,N_9204);
nor U9622 (N_9622,N_9357,N_9246);
nand U9623 (N_9623,N_9026,N_9348);
and U9624 (N_9624,N_9460,N_9010);
nor U9625 (N_9625,N_9402,N_9078);
nor U9626 (N_9626,N_9351,N_9341);
nand U9627 (N_9627,N_9452,N_9439);
nand U9628 (N_9628,N_9312,N_9155);
and U9629 (N_9629,N_9224,N_9334);
and U9630 (N_9630,N_9303,N_9013);
or U9631 (N_9631,N_9370,N_9457);
nor U9632 (N_9632,N_9412,N_9278);
nand U9633 (N_9633,N_9464,N_9221);
xnor U9634 (N_9634,N_9187,N_9287);
or U9635 (N_9635,N_9214,N_9127);
or U9636 (N_9636,N_9343,N_9271);
and U9637 (N_9637,N_9332,N_9212);
or U9638 (N_9638,N_9210,N_9077);
and U9639 (N_9639,N_9158,N_9216);
nor U9640 (N_9640,N_9014,N_9151);
and U9641 (N_9641,N_9272,N_9104);
and U9642 (N_9642,N_9138,N_9258);
nor U9643 (N_9643,N_9199,N_9320);
or U9644 (N_9644,N_9304,N_9326);
nor U9645 (N_9645,N_9435,N_9463);
xnor U9646 (N_9646,N_9018,N_9284);
xnor U9647 (N_9647,N_9070,N_9122);
xnor U9648 (N_9648,N_9028,N_9107);
xnor U9649 (N_9649,N_9315,N_9331);
and U9650 (N_9650,N_9033,N_9336);
or U9651 (N_9651,N_9184,N_9117);
or U9652 (N_9652,N_9408,N_9071);
nor U9653 (N_9653,N_9133,N_9458);
xnor U9654 (N_9654,N_9019,N_9263);
xnor U9655 (N_9655,N_9443,N_9154);
and U9656 (N_9656,N_9129,N_9235);
and U9657 (N_9657,N_9349,N_9039);
xnor U9658 (N_9658,N_9438,N_9356);
xor U9659 (N_9659,N_9455,N_9491);
xor U9660 (N_9660,N_9245,N_9433);
nand U9661 (N_9661,N_9499,N_9407);
xnor U9662 (N_9662,N_9386,N_9364);
nand U9663 (N_9663,N_9476,N_9497);
nor U9664 (N_9664,N_9188,N_9112);
or U9665 (N_9665,N_9192,N_9313);
nor U9666 (N_9666,N_9231,N_9365);
xor U9667 (N_9667,N_9323,N_9174);
nor U9668 (N_9668,N_9198,N_9428);
xnor U9669 (N_9669,N_9294,N_9483);
and U9670 (N_9670,N_9183,N_9191);
nor U9671 (N_9671,N_9005,N_9091);
or U9672 (N_9672,N_9419,N_9266);
nand U9673 (N_9673,N_9056,N_9236);
nor U9674 (N_9674,N_9234,N_9051);
nand U9675 (N_9675,N_9420,N_9111);
xor U9676 (N_9676,N_9034,N_9118);
xnor U9677 (N_9677,N_9368,N_9324);
nor U9678 (N_9678,N_9027,N_9256);
nand U9679 (N_9679,N_9230,N_9344);
and U9680 (N_9680,N_9239,N_9437);
nor U9681 (N_9681,N_9282,N_9280);
and U9682 (N_9682,N_9169,N_9414);
nand U9683 (N_9683,N_9267,N_9494);
xor U9684 (N_9684,N_9181,N_9145);
nand U9685 (N_9685,N_9290,N_9265);
or U9686 (N_9686,N_9442,N_9120);
or U9687 (N_9687,N_9388,N_9147);
and U9688 (N_9688,N_9362,N_9373);
nor U9689 (N_9689,N_9252,N_9250);
xor U9690 (N_9690,N_9114,N_9023);
and U9691 (N_9691,N_9069,N_9378);
nor U9692 (N_9692,N_9126,N_9495);
xnor U9693 (N_9693,N_9406,N_9347);
nand U9694 (N_9694,N_9017,N_9411);
nor U9695 (N_9695,N_9398,N_9063);
or U9696 (N_9696,N_9135,N_9307);
xnor U9697 (N_9697,N_9300,N_9065);
nand U9698 (N_9698,N_9172,N_9389);
nor U9699 (N_9699,N_9047,N_9418);
nand U9700 (N_9700,N_9035,N_9492);
nand U9701 (N_9701,N_9201,N_9270);
and U9702 (N_9702,N_9281,N_9168);
and U9703 (N_9703,N_9015,N_9484);
or U9704 (N_9704,N_9473,N_9139);
xnor U9705 (N_9705,N_9488,N_9470);
or U9706 (N_9706,N_9115,N_9092);
or U9707 (N_9707,N_9232,N_9004);
nand U9708 (N_9708,N_9180,N_9337);
or U9709 (N_9709,N_9134,N_9262);
and U9710 (N_9710,N_9449,N_9083);
nand U9711 (N_9711,N_9352,N_9030);
xor U9712 (N_9712,N_9159,N_9006);
and U9713 (N_9713,N_9279,N_9042);
nor U9714 (N_9714,N_9361,N_9404);
or U9715 (N_9715,N_9011,N_9311);
nor U9716 (N_9716,N_9325,N_9022);
and U9717 (N_9717,N_9108,N_9453);
and U9718 (N_9718,N_9156,N_9179);
and U9719 (N_9719,N_9218,N_9286);
nor U9720 (N_9720,N_9346,N_9153);
nand U9721 (N_9721,N_9392,N_9085);
xnor U9722 (N_9722,N_9376,N_9467);
and U9723 (N_9723,N_9094,N_9084);
nor U9724 (N_9724,N_9391,N_9148);
xnor U9725 (N_9725,N_9295,N_9474);
and U9726 (N_9726,N_9469,N_9157);
nand U9727 (N_9727,N_9369,N_9099);
xnor U9728 (N_9728,N_9319,N_9160);
and U9729 (N_9729,N_9430,N_9097);
nor U9730 (N_9730,N_9081,N_9166);
and U9731 (N_9731,N_9064,N_9044);
nand U9732 (N_9732,N_9074,N_9238);
and U9733 (N_9733,N_9021,N_9400);
xor U9734 (N_9734,N_9088,N_9194);
or U9735 (N_9735,N_9397,N_9052);
nand U9736 (N_9736,N_9103,N_9283);
xor U9737 (N_9737,N_9175,N_9355);
nand U9738 (N_9738,N_9310,N_9060);
nand U9739 (N_9739,N_9466,N_9340);
nand U9740 (N_9740,N_9441,N_9321);
or U9741 (N_9741,N_9205,N_9481);
or U9742 (N_9742,N_9101,N_9110);
or U9743 (N_9743,N_9363,N_9399);
xor U9744 (N_9744,N_9128,N_9137);
or U9745 (N_9745,N_9447,N_9367);
nor U9746 (N_9746,N_9228,N_9067);
nor U9747 (N_9747,N_9479,N_9345);
and U9748 (N_9748,N_9095,N_9486);
nor U9749 (N_9749,N_9471,N_9206);
nor U9750 (N_9750,N_9441,N_9260);
or U9751 (N_9751,N_9126,N_9427);
xnor U9752 (N_9752,N_9059,N_9053);
nand U9753 (N_9753,N_9082,N_9496);
nor U9754 (N_9754,N_9249,N_9247);
nand U9755 (N_9755,N_9494,N_9271);
nand U9756 (N_9756,N_9162,N_9396);
nand U9757 (N_9757,N_9319,N_9042);
nor U9758 (N_9758,N_9232,N_9451);
nand U9759 (N_9759,N_9153,N_9368);
xor U9760 (N_9760,N_9314,N_9373);
nor U9761 (N_9761,N_9225,N_9416);
xnor U9762 (N_9762,N_9485,N_9330);
and U9763 (N_9763,N_9064,N_9184);
or U9764 (N_9764,N_9306,N_9396);
and U9765 (N_9765,N_9094,N_9482);
or U9766 (N_9766,N_9397,N_9138);
or U9767 (N_9767,N_9087,N_9014);
nand U9768 (N_9768,N_9267,N_9415);
nand U9769 (N_9769,N_9443,N_9188);
nor U9770 (N_9770,N_9381,N_9449);
or U9771 (N_9771,N_9263,N_9316);
nand U9772 (N_9772,N_9287,N_9466);
and U9773 (N_9773,N_9319,N_9079);
nor U9774 (N_9774,N_9484,N_9116);
nand U9775 (N_9775,N_9279,N_9159);
nor U9776 (N_9776,N_9347,N_9004);
or U9777 (N_9777,N_9372,N_9352);
nand U9778 (N_9778,N_9366,N_9339);
nand U9779 (N_9779,N_9008,N_9451);
nand U9780 (N_9780,N_9307,N_9427);
or U9781 (N_9781,N_9242,N_9133);
nor U9782 (N_9782,N_9058,N_9492);
and U9783 (N_9783,N_9025,N_9343);
and U9784 (N_9784,N_9207,N_9366);
nor U9785 (N_9785,N_9353,N_9292);
nand U9786 (N_9786,N_9141,N_9480);
and U9787 (N_9787,N_9134,N_9092);
xor U9788 (N_9788,N_9497,N_9368);
nor U9789 (N_9789,N_9349,N_9122);
nand U9790 (N_9790,N_9497,N_9448);
nor U9791 (N_9791,N_9477,N_9361);
or U9792 (N_9792,N_9137,N_9202);
xnor U9793 (N_9793,N_9007,N_9302);
nor U9794 (N_9794,N_9110,N_9419);
or U9795 (N_9795,N_9363,N_9206);
nor U9796 (N_9796,N_9169,N_9129);
nor U9797 (N_9797,N_9319,N_9313);
nand U9798 (N_9798,N_9418,N_9021);
xor U9799 (N_9799,N_9411,N_9053);
xor U9800 (N_9800,N_9156,N_9137);
nor U9801 (N_9801,N_9385,N_9161);
or U9802 (N_9802,N_9264,N_9196);
nor U9803 (N_9803,N_9186,N_9373);
or U9804 (N_9804,N_9231,N_9267);
nand U9805 (N_9805,N_9386,N_9422);
and U9806 (N_9806,N_9316,N_9494);
nor U9807 (N_9807,N_9237,N_9347);
nor U9808 (N_9808,N_9042,N_9373);
xnor U9809 (N_9809,N_9217,N_9143);
nor U9810 (N_9810,N_9408,N_9079);
and U9811 (N_9811,N_9054,N_9307);
nand U9812 (N_9812,N_9268,N_9483);
xor U9813 (N_9813,N_9361,N_9138);
or U9814 (N_9814,N_9168,N_9061);
and U9815 (N_9815,N_9407,N_9065);
nand U9816 (N_9816,N_9462,N_9411);
nor U9817 (N_9817,N_9226,N_9442);
xnor U9818 (N_9818,N_9495,N_9401);
or U9819 (N_9819,N_9030,N_9405);
nand U9820 (N_9820,N_9357,N_9329);
xnor U9821 (N_9821,N_9054,N_9381);
xnor U9822 (N_9822,N_9462,N_9092);
nor U9823 (N_9823,N_9298,N_9282);
nand U9824 (N_9824,N_9066,N_9399);
nor U9825 (N_9825,N_9001,N_9279);
and U9826 (N_9826,N_9347,N_9041);
nor U9827 (N_9827,N_9053,N_9124);
and U9828 (N_9828,N_9223,N_9076);
nor U9829 (N_9829,N_9135,N_9143);
nor U9830 (N_9830,N_9145,N_9162);
or U9831 (N_9831,N_9029,N_9374);
nor U9832 (N_9832,N_9364,N_9036);
nand U9833 (N_9833,N_9492,N_9041);
and U9834 (N_9834,N_9168,N_9073);
nor U9835 (N_9835,N_9352,N_9115);
and U9836 (N_9836,N_9381,N_9407);
and U9837 (N_9837,N_9422,N_9276);
xor U9838 (N_9838,N_9499,N_9019);
xnor U9839 (N_9839,N_9033,N_9498);
xor U9840 (N_9840,N_9000,N_9077);
xnor U9841 (N_9841,N_9370,N_9458);
and U9842 (N_9842,N_9024,N_9072);
and U9843 (N_9843,N_9134,N_9036);
or U9844 (N_9844,N_9320,N_9256);
and U9845 (N_9845,N_9382,N_9406);
nor U9846 (N_9846,N_9186,N_9015);
and U9847 (N_9847,N_9154,N_9271);
xor U9848 (N_9848,N_9455,N_9304);
nand U9849 (N_9849,N_9387,N_9009);
and U9850 (N_9850,N_9189,N_9158);
and U9851 (N_9851,N_9181,N_9292);
and U9852 (N_9852,N_9222,N_9469);
or U9853 (N_9853,N_9298,N_9211);
xnor U9854 (N_9854,N_9062,N_9030);
and U9855 (N_9855,N_9083,N_9262);
and U9856 (N_9856,N_9492,N_9417);
or U9857 (N_9857,N_9003,N_9059);
xnor U9858 (N_9858,N_9282,N_9236);
or U9859 (N_9859,N_9173,N_9224);
nand U9860 (N_9860,N_9284,N_9259);
nand U9861 (N_9861,N_9354,N_9142);
nand U9862 (N_9862,N_9378,N_9321);
and U9863 (N_9863,N_9068,N_9126);
nor U9864 (N_9864,N_9303,N_9494);
or U9865 (N_9865,N_9023,N_9088);
nor U9866 (N_9866,N_9352,N_9368);
nor U9867 (N_9867,N_9276,N_9078);
or U9868 (N_9868,N_9064,N_9247);
or U9869 (N_9869,N_9173,N_9280);
or U9870 (N_9870,N_9449,N_9405);
nand U9871 (N_9871,N_9116,N_9347);
or U9872 (N_9872,N_9436,N_9246);
nand U9873 (N_9873,N_9127,N_9386);
xor U9874 (N_9874,N_9032,N_9114);
xnor U9875 (N_9875,N_9358,N_9028);
nor U9876 (N_9876,N_9132,N_9432);
xor U9877 (N_9877,N_9131,N_9134);
and U9878 (N_9878,N_9447,N_9269);
or U9879 (N_9879,N_9299,N_9025);
xor U9880 (N_9880,N_9238,N_9007);
nand U9881 (N_9881,N_9032,N_9409);
nand U9882 (N_9882,N_9328,N_9363);
and U9883 (N_9883,N_9277,N_9253);
xnor U9884 (N_9884,N_9251,N_9010);
nand U9885 (N_9885,N_9426,N_9194);
or U9886 (N_9886,N_9235,N_9451);
nand U9887 (N_9887,N_9272,N_9048);
or U9888 (N_9888,N_9225,N_9178);
and U9889 (N_9889,N_9363,N_9026);
or U9890 (N_9890,N_9285,N_9333);
nand U9891 (N_9891,N_9096,N_9471);
nor U9892 (N_9892,N_9339,N_9496);
and U9893 (N_9893,N_9206,N_9238);
or U9894 (N_9894,N_9406,N_9445);
nor U9895 (N_9895,N_9115,N_9228);
and U9896 (N_9896,N_9242,N_9120);
and U9897 (N_9897,N_9290,N_9072);
or U9898 (N_9898,N_9263,N_9021);
or U9899 (N_9899,N_9174,N_9458);
nand U9900 (N_9900,N_9428,N_9258);
and U9901 (N_9901,N_9382,N_9422);
xor U9902 (N_9902,N_9453,N_9432);
nand U9903 (N_9903,N_9323,N_9018);
xnor U9904 (N_9904,N_9200,N_9206);
and U9905 (N_9905,N_9440,N_9100);
xor U9906 (N_9906,N_9404,N_9173);
or U9907 (N_9907,N_9053,N_9462);
nor U9908 (N_9908,N_9083,N_9194);
nand U9909 (N_9909,N_9061,N_9002);
or U9910 (N_9910,N_9147,N_9306);
nor U9911 (N_9911,N_9271,N_9088);
nor U9912 (N_9912,N_9484,N_9495);
xor U9913 (N_9913,N_9095,N_9074);
and U9914 (N_9914,N_9047,N_9454);
and U9915 (N_9915,N_9343,N_9258);
or U9916 (N_9916,N_9492,N_9172);
nor U9917 (N_9917,N_9405,N_9185);
nand U9918 (N_9918,N_9278,N_9443);
xnor U9919 (N_9919,N_9300,N_9428);
xor U9920 (N_9920,N_9448,N_9209);
and U9921 (N_9921,N_9346,N_9215);
xnor U9922 (N_9922,N_9275,N_9354);
or U9923 (N_9923,N_9086,N_9019);
and U9924 (N_9924,N_9344,N_9172);
nand U9925 (N_9925,N_9030,N_9069);
nand U9926 (N_9926,N_9013,N_9346);
and U9927 (N_9927,N_9369,N_9395);
xnor U9928 (N_9928,N_9309,N_9453);
nand U9929 (N_9929,N_9243,N_9071);
nor U9930 (N_9930,N_9137,N_9037);
nor U9931 (N_9931,N_9345,N_9068);
nand U9932 (N_9932,N_9174,N_9467);
or U9933 (N_9933,N_9066,N_9406);
and U9934 (N_9934,N_9174,N_9151);
and U9935 (N_9935,N_9118,N_9002);
or U9936 (N_9936,N_9051,N_9386);
and U9937 (N_9937,N_9409,N_9378);
and U9938 (N_9938,N_9494,N_9300);
nor U9939 (N_9939,N_9082,N_9294);
or U9940 (N_9940,N_9155,N_9109);
or U9941 (N_9941,N_9342,N_9287);
or U9942 (N_9942,N_9313,N_9383);
xor U9943 (N_9943,N_9124,N_9222);
and U9944 (N_9944,N_9280,N_9210);
or U9945 (N_9945,N_9252,N_9001);
nor U9946 (N_9946,N_9071,N_9049);
nand U9947 (N_9947,N_9499,N_9328);
nand U9948 (N_9948,N_9160,N_9100);
or U9949 (N_9949,N_9248,N_9045);
or U9950 (N_9950,N_9328,N_9449);
and U9951 (N_9951,N_9463,N_9076);
and U9952 (N_9952,N_9456,N_9336);
nand U9953 (N_9953,N_9084,N_9431);
xnor U9954 (N_9954,N_9340,N_9465);
xnor U9955 (N_9955,N_9066,N_9485);
nor U9956 (N_9956,N_9203,N_9086);
or U9957 (N_9957,N_9295,N_9044);
or U9958 (N_9958,N_9410,N_9237);
nand U9959 (N_9959,N_9361,N_9473);
nor U9960 (N_9960,N_9065,N_9144);
and U9961 (N_9961,N_9043,N_9349);
nand U9962 (N_9962,N_9061,N_9284);
or U9963 (N_9963,N_9028,N_9324);
nor U9964 (N_9964,N_9238,N_9172);
or U9965 (N_9965,N_9035,N_9087);
nand U9966 (N_9966,N_9167,N_9233);
and U9967 (N_9967,N_9243,N_9208);
nand U9968 (N_9968,N_9483,N_9259);
and U9969 (N_9969,N_9076,N_9207);
nand U9970 (N_9970,N_9309,N_9238);
and U9971 (N_9971,N_9067,N_9150);
nor U9972 (N_9972,N_9344,N_9167);
xor U9973 (N_9973,N_9302,N_9257);
or U9974 (N_9974,N_9430,N_9383);
xnor U9975 (N_9975,N_9292,N_9003);
or U9976 (N_9976,N_9068,N_9201);
and U9977 (N_9977,N_9385,N_9477);
xor U9978 (N_9978,N_9031,N_9075);
xor U9979 (N_9979,N_9246,N_9329);
nand U9980 (N_9980,N_9362,N_9229);
nor U9981 (N_9981,N_9132,N_9373);
nand U9982 (N_9982,N_9419,N_9115);
nor U9983 (N_9983,N_9084,N_9482);
or U9984 (N_9984,N_9375,N_9249);
and U9985 (N_9985,N_9454,N_9241);
nand U9986 (N_9986,N_9337,N_9191);
or U9987 (N_9987,N_9432,N_9391);
or U9988 (N_9988,N_9332,N_9084);
nand U9989 (N_9989,N_9158,N_9114);
or U9990 (N_9990,N_9259,N_9188);
or U9991 (N_9991,N_9127,N_9302);
and U9992 (N_9992,N_9266,N_9320);
or U9993 (N_9993,N_9167,N_9104);
nand U9994 (N_9994,N_9207,N_9319);
nand U9995 (N_9995,N_9299,N_9454);
and U9996 (N_9996,N_9161,N_9271);
nand U9997 (N_9997,N_9046,N_9269);
xnor U9998 (N_9998,N_9413,N_9259);
nor U9999 (N_9999,N_9303,N_9176);
xor U10000 (N_10000,N_9814,N_9789);
and U10001 (N_10001,N_9762,N_9958);
or U10002 (N_10002,N_9643,N_9927);
nor U10003 (N_10003,N_9959,N_9585);
xor U10004 (N_10004,N_9882,N_9987);
and U10005 (N_10005,N_9887,N_9595);
nand U10006 (N_10006,N_9972,N_9936);
xnor U10007 (N_10007,N_9978,N_9630);
nor U10008 (N_10008,N_9700,N_9589);
and U10009 (N_10009,N_9827,N_9939);
xor U10010 (N_10010,N_9629,N_9813);
nand U10011 (N_10011,N_9581,N_9672);
and U10012 (N_10012,N_9916,N_9898);
nor U10013 (N_10013,N_9949,N_9593);
and U10014 (N_10014,N_9596,N_9893);
xor U10015 (N_10015,N_9655,N_9508);
nand U10016 (N_10016,N_9962,N_9802);
xor U10017 (N_10017,N_9851,N_9966);
or U10018 (N_10018,N_9710,N_9714);
xnor U10019 (N_10019,N_9905,N_9664);
nand U10020 (N_10020,N_9872,N_9708);
and U10021 (N_10021,N_9942,N_9976);
nor U10022 (N_10022,N_9839,N_9723);
nor U10023 (N_10023,N_9575,N_9863);
xor U10024 (N_10024,N_9734,N_9638);
nand U10025 (N_10025,N_9536,N_9716);
or U10026 (N_10026,N_9844,N_9721);
nor U10027 (N_10027,N_9766,N_9564);
xor U10028 (N_10028,N_9828,N_9569);
and U10029 (N_10029,N_9786,N_9590);
or U10030 (N_10030,N_9707,N_9731);
and U10031 (N_10031,N_9907,N_9545);
nand U10032 (N_10032,N_9746,N_9877);
nor U10033 (N_10033,N_9832,N_9873);
or U10034 (N_10034,N_9718,N_9588);
nand U10035 (N_10035,N_9522,N_9791);
xnor U10036 (N_10036,N_9689,N_9621);
xnor U10037 (N_10037,N_9546,N_9777);
nor U10038 (N_10038,N_9678,N_9523);
and U10039 (N_10039,N_9729,N_9561);
nor U10040 (N_10040,N_9835,N_9822);
or U10041 (N_10041,N_9687,N_9517);
nor U10042 (N_10042,N_9598,N_9850);
nand U10043 (N_10043,N_9560,N_9651);
nand U10044 (N_10044,N_9684,N_9500);
or U10045 (N_10045,N_9566,N_9625);
xnor U10046 (N_10046,N_9904,N_9914);
xnor U10047 (N_10047,N_9864,N_9792);
and U10048 (N_10048,N_9856,N_9520);
xnor U10049 (N_10049,N_9954,N_9506);
nand U10050 (N_10050,N_9549,N_9940);
nand U10051 (N_10051,N_9645,N_9610);
or U10052 (N_10052,N_9849,N_9909);
xnor U10053 (N_10053,N_9741,N_9885);
nor U10054 (N_10054,N_9799,N_9556);
xor U10055 (N_10055,N_9930,N_9986);
xnor U10056 (N_10056,N_9899,N_9830);
xnor U10057 (N_10057,N_9964,N_9913);
or U10058 (N_10058,N_9519,N_9858);
or U10059 (N_10059,N_9997,N_9558);
xnor U10060 (N_10060,N_9815,N_9703);
xnor U10061 (N_10061,N_9695,N_9511);
or U10062 (N_10062,N_9646,N_9884);
xor U10063 (N_10063,N_9715,N_9807);
xnor U10064 (N_10064,N_9670,N_9539);
or U10065 (N_10065,N_9749,N_9597);
or U10066 (N_10066,N_9552,N_9870);
and U10067 (N_10067,N_9614,N_9915);
or U10068 (N_10068,N_9578,N_9767);
xnor U10069 (N_10069,N_9607,N_9618);
nor U10070 (N_10070,N_9823,N_9737);
nand U10071 (N_10071,N_9859,N_9572);
and U10072 (N_10072,N_9640,N_9768);
and U10073 (N_10073,N_9763,N_9674);
nor U10074 (N_10074,N_9793,N_9754);
xor U10075 (N_10075,N_9676,N_9975);
and U10076 (N_10076,N_9981,N_9960);
or U10077 (N_10077,N_9953,N_9881);
and U10078 (N_10078,N_9696,N_9609);
nand U10079 (N_10079,N_9837,N_9748);
xnor U10080 (N_10080,N_9803,N_9977);
and U10081 (N_10081,N_9626,N_9557);
and U10082 (N_10082,N_9667,N_9925);
or U10083 (N_10083,N_9753,N_9888);
nor U10084 (N_10084,N_9613,N_9804);
xor U10085 (N_10085,N_9761,N_9886);
or U10086 (N_10086,N_9796,N_9562);
nand U10087 (N_10087,N_9509,N_9834);
or U10088 (N_10088,N_9603,N_9711);
or U10089 (N_10089,N_9658,N_9847);
nor U10090 (N_10090,N_9820,N_9554);
xnor U10091 (N_10091,N_9620,N_9635);
or U10092 (N_10092,N_9512,N_9961);
or U10093 (N_10093,N_9633,N_9984);
xor U10094 (N_10094,N_9669,N_9829);
xnor U10095 (N_10095,N_9713,N_9782);
nor U10096 (N_10096,N_9533,N_9866);
xor U10097 (N_10097,N_9883,N_9892);
xor U10098 (N_10098,N_9704,N_9662);
or U10099 (N_10099,N_9547,N_9769);
or U10100 (N_10100,N_9524,N_9602);
or U10101 (N_10101,N_9908,N_9518);
or U10102 (N_10102,N_9636,N_9526);
or U10103 (N_10103,N_9974,N_9994);
nand U10104 (N_10104,N_9648,N_9957);
or U10105 (N_10105,N_9706,N_9649);
xor U10106 (N_10106,N_9641,N_9502);
nand U10107 (N_10107,N_9995,N_9501);
and U10108 (N_10108,N_9642,N_9673);
xnor U10109 (N_10109,N_9969,N_9542);
or U10110 (N_10110,N_9559,N_9826);
and U10111 (N_10111,N_9819,N_9751);
nand U10112 (N_10112,N_9611,N_9776);
and U10113 (N_10113,N_9697,N_9513);
or U10114 (N_10114,N_9982,N_9805);
nand U10115 (N_10115,N_9660,N_9910);
nand U10116 (N_10116,N_9929,N_9817);
or U10117 (N_10117,N_9816,N_9586);
xor U10118 (N_10118,N_9623,N_9604);
and U10119 (N_10119,N_9875,N_9699);
and U10120 (N_10120,N_9926,N_9808);
xnor U10121 (N_10121,N_9980,N_9783);
or U10122 (N_10122,N_9568,N_9920);
nand U10123 (N_10123,N_9690,N_9738);
and U10124 (N_10124,N_9727,N_9685);
nor U10125 (N_10125,N_9967,N_9529);
and U10126 (N_10126,N_9686,N_9553);
xor U10127 (N_10127,N_9652,N_9668);
or U10128 (N_10128,N_9531,N_9582);
and U10129 (N_10129,N_9608,N_9730);
nand U10130 (N_10130,N_9945,N_9989);
or U10131 (N_10131,N_9831,N_9999);
or U10132 (N_10132,N_9965,N_9579);
and U10133 (N_10133,N_9891,N_9911);
nor U10134 (N_10134,N_9983,N_9797);
nor U10135 (N_10135,N_9944,N_9938);
nor U10136 (N_10136,N_9902,N_9567);
nor U10137 (N_10137,N_9505,N_9950);
or U10138 (N_10138,N_9871,N_9855);
or U10139 (N_10139,N_9532,N_9912);
or U10140 (N_10140,N_9860,N_9724);
nor U10141 (N_10141,N_9992,N_9903);
nand U10142 (N_10142,N_9933,N_9548);
or U10143 (N_10143,N_9628,N_9919);
or U10144 (N_10144,N_9906,N_9683);
xnor U10145 (N_10145,N_9555,N_9865);
nand U10146 (N_10146,N_9812,N_9771);
nand U10147 (N_10147,N_9922,N_9979);
nand U10148 (N_10148,N_9778,N_9504);
and U10149 (N_10149,N_9712,N_9619);
and U10150 (N_10150,N_9795,N_9833);
xor U10151 (N_10151,N_9759,N_9848);
nor U10152 (N_10152,N_9874,N_9921);
nand U10153 (N_10153,N_9756,N_9631);
xor U10154 (N_10154,N_9634,N_9681);
xnor U10155 (N_10155,N_9719,N_9698);
nand U10156 (N_10156,N_9565,N_9838);
or U10157 (N_10157,N_9601,N_9750);
nand U10158 (N_10158,N_9988,N_9900);
or U10159 (N_10159,N_9705,N_9514);
nor U10160 (N_10160,N_9679,N_9653);
and U10161 (N_10161,N_9993,N_9781);
nand U10162 (N_10162,N_9709,N_9809);
or U10163 (N_10163,N_9854,N_9811);
or U10164 (N_10164,N_9970,N_9541);
and U10165 (N_10165,N_9946,N_9800);
xnor U10166 (N_10166,N_9740,N_9991);
or U10167 (N_10167,N_9821,N_9600);
xnor U10168 (N_10168,N_9507,N_9963);
nand U10169 (N_10169,N_9790,N_9901);
or U10170 (N_10170,N_9896,N_9757);
or U10171 (N_10171,N_9580,N_9521);
and U10172 (N_10172,N_9592,N_9842);
or U10173 (N_10173,N_9510,N_9932);
or U10174 (N_10174,N_9726,N_9682);
nor U10175 (N_10175,N_9952,N_9617);
nor U10176 (N_10176,N_9694,N_9841);
nor U10177 (N_10177,N_9576,N_9570);
or U10178 (N_10178,N_9563,N_9606);
nor U10179 (N_10179,N_9971,N_9722);
nor U10180 (N_10180,N_9535,N_9943);
nand U10181 (N_10181,N_9890,N_9889);
nand U10182 (N_10182,N_9528,N_9632);
nor U10183 (N_10183,N_9540,N_9515);
xor U10184 (N_10184,N_9654,N_9675);
nor U10185 (N_10185,N_9772,N_9941);
and U10186 (N_10186,N_9587,N_9937);
xor U10187 (N_10187,N_9503,N_9878);
nand U10188 (N_10188,N_9798,N_9577);
nor U10189 (N_10189,N_9573,N_9801);
nand U10190 (N_10190,N_9880,N_9951);
and U10191 (N_10191,N_9845,N_9584);
xnor U10192 (N_10192,N_9665,N_9998);
xor U10193 (N_10193,N_9717,N_9876);
nand U10194 (N_10194,N_9680,N_9612);
xnor U10195 (N_10195,N_9825,N_9773);
nand U10196 (N_10196,N_9760,N_9846);
and U10197 (N_10197,N_9571,N_9948);
or U10198 (N_10198,N_9688,N_9968);
xnor U10199 (N_10199,N_9840,N_9671);
or U10200 (N_10200,N_9692,N_9583);
nand U10201 (N_10201,N_9810,N_9770);
or U10202 (N_10202,N_9534,N_9639);
nor U10203 (N_10203,N_9666,N_9544);
nor U10204 (N_10204,N_9551,N_9947);
nor U10205 (N_10205,N_9918,N_9764);
nor U10206 (N_10206,N_9934,N_9543);
or U10207 (N_10207,N_9897,N_9720);
xor U10208 (N_10208,N_9869,N_9599);
xor U10209 (N_10209,N_9867,N_9996);
or U10210 (N_10210,N_9853,N_9659);
and U10211 (N_10211,N_9765,N_9806);
nand U10212 (N_10212,N_9787,N_9591);
nor U10213 (N_10213,N_9924,N_9574);
nand U10214 (N_10214,N_9743,N_9616);
and U10215 (N_10215,N_9538,N_9693);
and U10216 (N_10216,N_9733,N_9794);
or U10217 (N_10217,N_9985,N_9917);
xor U10218 (N_10218,N_9656,N_9928);
or U10219 (N_10219,N_9857,N_9879);
nor U10220 (N_10220,N_9702,N_9661);
xor U10221 (N_10221,N_9663,N_9728);
and U10222 (N_10222,N_9862,N_9605);
and U10223 (N_10223,N_9627,N_9736);
xor U10224 (N_10224,N_9657,N_9650);
or U10225 (N_10225,N_9824,N_9752);
xnor U10226 (N_10226,N_9550,N_9742);
and U10227 (N_10227,N_9990,N_9691);
and U10228 (N_10228,N_9747,N_9931);
xnor U10229 (N_10229,N_9774,N_9868);
nor U10230 (N_10230,N_9852,N_9755);
and U10231 (N_10231,N_9677,N_9894);
nor U10232 (N_10232,N_9923,N_9537);
or U10233 (N_10233,N_9732,N_9594);
nor U10234 (N_10234,N_9784,N_9836);
nor U10235 (N_10235,N_9956,N_9780);
nor U10236 (N_10236,N_9739,N_9779);
xnor U10237 (N_10237,N_9725,N_9955);
nand U10238 (N_10238,N_9530,N_9843);
nand U10239 (N_10239,N_9615,N_9745);
or U10240 (N_10240,N_9624,N_9701);
nand U10241 (N_10241,N_9758,N_9644);
nand U10242 (N_10242,N_9818,N_9647);
nor U10243 (N_10243,N_9735,N_9516);
xnor U10244 (N_10244,N_9525,N_9775);
xor U10245 (N_10245,N_9637,N_9895);
or U10246 (N_10246,N_9744,N_9622);
nor U10247 (N_10247,N_9973,N_9788);
nand U10248 (N_10248,N_9785,N_9527);
or U10249 (N_10249,N_9935,N_9861);
nand U10250 (N_10250,N_9741,N_9991);
nand U10251 (N_10251,N_9540,N_9555);
nand U10252 (N_10252,N_9973,N_9989);
nand U10253 (N_10253,N_9602,N_9749);
nor U10254 (N_10254,N_9878,N_9970);
and U10255 (N_10255,N_9685,N_9983);
and U10256 (N_10256,N_9770,N_9713);
nand U10257 (N_10257,N_9829,N_9891);
and U10258 (N_10258,N_9757,N_9783);
nor U10259 (N_10259,N_9630,N_9971);
and U10260 (N_10260,N_9751,N_9871);
nor U10261 (N_10261,N_9851,N_9855);
or U10262 (N_10262,N_9978,N_9857);
nor U10263 (N_10263,N_9996,N_9906);
or U10264 (N_10264,N_9834,N_9936);
and U10265 (N_10265,N_9623,N_9737);
nand U10266 (N_10266,N_9988,N_9979);
xnor U10267 (N_10267,N_9704,N_9567);
nor U10268 (N_10268,N_9726,N_9844);
and U10269 (N_10269,N_9781,N_9904);
xnor U10270 (N_10270,N_9946,N_9546);
and U10271 (N_10271,N_9946,N_9972);
or U10272 (N_10272,N_9858,N_9784);
xnor U10273 (N_10273,N_9887,N_9738);
nor U10274 (N_10274,N_9714,N_9816);
nand U10275 (N_10275,N_9651,N_9801);
xnor U10276 (N_10276,N_9697,N_9787);
nor U10277 (N_10277,N_9638,N_9699);
and U10278 (N_10278,N_9606,N_9921);
nor U10279 (N_10279,N_9513,N_9562);
nand U10280 (N_10280,N_9872,N_9621);
and U10281 (N_10281,N_9571,N_9591);
xnor U10282 (N_10282,N_9526,N_9746);
nor U10283 (N_10283,N_9936,N_9963);
nand U10284 (N_10284,N_9777,N_9940);
nand U10285 (N_10285,N_9765,N_9695);
or U10286 (N_10286,N_9567,N_9682);
or U10287 (N_10287,N_9985,N_9600);
or U10288 (N_10288,N_9542,N_9729);
or U10289 (N_10289,N_9858,N_9926);
xnor U10290 (N_10290,N_9923,N_9590);
and U10291 (N_10291,N_9576,N_9580);
nand U10292 (N_10292,N_9863,N_9547);
nor U10293 (N_10293,N_9623,N_9725);
and U10294 (N_10294,N_9801,N_9716);
and U10295 (N_10295,N_9754,N_9685);
and U10296 (N_10296,N_9840,N_9960);
or U10297 (N_10297,N_9771,N_9510);
nand U10298 (N_10298,N_9629,N_9845);
xnor U10299 (N_10299,N_9742,N_9861);
nor U10300 (N_10300,N_9860,N_9891);
nor U10301 (N_10301,N_9981,N_9762);
nand U10302 (N_10302,N_9545,N_9827);
nor U10303 (N_10303,N_9541,N_9921);
nor U10304 (N_10304,N_9963,N_9957);
xor U10305 (N_10305,N_9653,N_9749);
or U10306 (N_10306,N_9732,N_9599);
or U10307 (N_10307,N_9580,N_9849);
and U10308 (N_10308,N_9998,N_9666);
nand U10309 (N_10309,N_9651,N_9671);
nand U10310 (N_10310,N_9664,N_9833);
xor U10311 (N_10311,N_9995,N_9538);
xnor U10312 (N_10312,N_9900,N_9857);
xor U10313 (N_10313,N_9683,N_9596);
or U10314 (N_10314,N_9807,N_9674);
nor U10315 (N_10315,N_9643,N_9926);
xor U10316 (N_10316,N_9670,N_9642);
or U10317 (N_10317,N_9836,N_9580);
nor U10318 (N_10318,N_9569,N_9566);
or U10319 (N_10319,N_9854,N_9559);
nand U10320 (N_10320,N_9914,N_9997);
or U10321 (N_10321,N_9982,N_9948);
or U10322 (N_10322,N_9867,N_9799);
or U10323 (N_10323,N_9697,N_9722);
or U10324 (N_10324,N_9715,N_9826);
and U10325 (N_10325,N_9994,N_9647);
nand U10326 (N_10326,N_9635,N_9751);
or U10327 (N_10327,N_9979,N_9602);
xnor U10328 (N_10328,N_9922,N_9765);
nand U10329 (N_10329,N_9834,N_9553);
and U10330 (N_10330,N_9590,N_9567);
xnor U10331 (N_10331,N_9933,N_9630);
and U10332 (N_10332,N_9590,N_9652);
or U10333 (N_10333,N_9789,N_9925);
nor U10334 (N_10334,N_9558,N_9515);
nand U10335 (N_10335,N_9634,N_9582);
nand U10336 (N_10336,N_9877,N_9955);
nor U10337 (N_10337,N_9785,N_9973);
or U10338 (N_10338,N_9962,N_9572);
or U10339 (N_10339,N_9866,N_9706);
nand U10340 (N_10340,N_9652,N_9536);
nand U10341 (N_10341,N_9971,N_9718);
or U10342 (N_10342,N_9952,N_9766);
or U10343 (N_10343,N_9795,N_9859);
nand U10344 (N_10344,N_9595,N_9650);
nand U10345 (N_10345,N_9901,N_9615);
xor U10346 (N_10346,N_9503,N_9930);
and U10347 (N_10347,N_9792,N_9906);
and U10348 (N_10348,N_9916,N_9808);
or U10349 (N_10349,N_9995,N_9973);
nand U10350 (N_10350,N_9900,N_9791);
nand U10351 (N_10351,N_9766,N_9508);
and U10352 (N_10352,N_9607,N_9521);
nor U10353 (N_10353,N_9789,N_9680);
or U10354 (N_10354,N_9998,N_9632);
nor U10355 (N_10355,N_9929,N_9755);
and U10356 (N_10356,N_9739,N_9718);
or U10357 (N_10357,N_9859,N_9732);
and U10358 (N_10358,N_9930,N_9586);
nor U10359 (N_10359,N_9835,N_9616);
nand U10360 (N_10360,N_9886,N_9752);
nand U10361 (N_10361,N_9948,N_9860);
nor U10362 (N_10362,N_9531,N_9794);
or U10363 (N_10363,N_9537,N_9574);
xnor U10364 (N_10364,N_9635,N_9892);
nor U10365 (N_10365,N_9884,N_9597);
and U10366 (N_10366,N_9655,N_9645);
xor U10367 (N_10367,N_9840,N_9810);
and U10368 (N_10368,N_9761,N_9901);
or U10369 (N_10369,N_9978,N_9688);
nand U10370 (N_10370,N_9776,N_9644);
nand U10371 (N_10371,N_9816,N_9631);
nand U10372 (N_10372,N_9700,N_9896);
and U10373 (N_10373,N_9920,N_9889);
and U10374 (N_10374,N_9745,N_9949);
nand U10375 (N_10375,N_9749,N_9768);
or U10376 (N_10376,N_9843,N_9754);
nor U10377 (N_10377,N_9521,N_9643);
and U10378 (N_10378,N_9563,N_9863);
or U10379 (N_10379,N_9691,N_9768);
xor U10380 (N_10380,N_9536,N_9516);
and U10381 (N_10381,N_9951,N_9585);
and U10382 (N_10382,N_9772,N_9698);
nor U10383 (N_10383,N_9831,N_9757);
nand U10384 (N_10384,N_9778,N_9951);
and U10385 (N_10385,N_9951,N_9714);
or U10386 (N_10386,N_9805,N_9577);
and U10387 (N_10387,N_9529,N_9897);
or U10388 (N_10388,N_9633,N_9919);
nor U10389 (N_10389,N_9836,N_9883);
xor U10390 (N_10390,N_9692,N_9994);
and U10391 (N_10391,N_9789,N_9775);
or U10392 (N_10392,N_9750,N_9652);
xnor U10393 (N_10393,N_9988,N_9660);
xor U10394 (N_10394,N_9922,N_9956);
nor U10395 (N_10395,N_9688,N_9903);
xor U10396 (N_10396,N_9595,N_9592);
xnor U10397 (N_10397,N_9722,N_9621);
nor U10398 (N_10398,N_9708,N_9978);
xor U10399 (N_10399,N_9535,N_9841);
nand U10400 (N_10400,N_9990,N_9804);
xnor U10401 (N_10401,N_9726,N_9894);
and U10402 (N_10402,N_9713,N_9832);
xor U10403 (N_10403,N_9903,N_9984);
nand U10404 (N_10404,N_9986,N_9940);
nor U10405 (N_10405,N_9838,N_9928);
xor U10406 (N_10406,N_9547,N_9527);
or U10407 (N_10407,N_9848,N_9640);
or U10408 (N_10408,N_9717,N_9568);
xor U10409 (N_10409,N_9536,N_9971);
and U10410 (N_10410,N_9720,N_9667);
nor U10411 (N_10411,N_9901,N_9839);
nand U10412 (N_10412,N_9963,N_9921);
or U10413 (N_10413,N_9812,N_9558);
nand U10414 (N_10414,N_9733,N_9789);
nor U10415 (N_10415,N_9866,N_9861);
nor U10416 (N_10416,N_9957,N_9774);
xnor U10417 (N_10417,N_9882,N_9694);
and U10418 (N_10418,N_9704,N_9929);
and U10419 (N_10419,N_9730,N_9959);
nand U10420 (N_10420,N_9873,N_9765);
or U10421 (N_10421,N_9893,N_9659);
and U10422 (N_10422,N_9621,N_9940);
and U10423 (N_10423,N_9533,N_9540);
and U10424 (N_10424,N_9907,N_9945);
xnor U10425 (N_10425,N_9839,N_9846);
and U10426 (N_10426,N_9726,N_9924);
nor U10427 (N_10427,N_9967,N_9773);
and U10428 (N_10428,N_9867,N_9904);
xnor U10429 (N_10429,N_9533,N_9810);
nor U10430 (N_10430,N_9802,N_9523);
nand U10431 (N_10431,N_9965,N_9525);
or U10432 (N_10432,N_9995,N_9700);
xnor U10433 (N_10433,N_9689,N_9788);
nand U10434 (N_10434,N_9694,N_9759);
xnor U10435 (N_10435,N_9841,N_9633);
and U10436 (N_10436,N_9739,N_9622);
nor U10437 (N_10437,N_9614,N_9575);
and U10438 (N_10438,N_9887,N_9901);
and U10439 (N_10439,N_9554,N_9518);
and U10440 (N_10440,N_9735,N_9525);
xor U10441 (N_10441,N_9917,N_9554);
nand U10442 (N_10442,N_9995,N_9686);
xnor U10443 (N_10443,N_9941,N_9602);
nor U10444 (N_10444,N_9812,N_9508);
nand U10445 (N_10445,N_9595,N_9893);
or U10446 (N_10446,N_9907,N_9755);
and U10447 (N_10447,N_9822,N_9839);
xnor U10448 (N_10448,N_9972,N_9806);
xor U10449 (N_10449,N_9547,N_9737);
or U10450 (N_10450,N_9540,N_9874);
nand U10451 (N_10451,N_9697,N_9639);
xnor U10452 (N_10452,N_9901,N_9512);
xor U10453 (N_10453,N_9645,N_9852);
and U10454 (N_10454,N_9895,N_9584);
or U10455 (N_10455,N_9699,N_9886);
xnor U10456 (N_10456,N_9520,N_9660);
nand U10457 (N_10457,N_9513,N_9639);
xor U10458 (N_10458,N_9783,N_9551);
xor U10459 (N_10459,N_9847,N_9662);
xnor U10460 (N_10460,N_9949,N_9727);
nor U10461 (N_10461,N_9690,N_9976);
nand U10462 (N_10462,N_9540,N_9822);
nor U10463 (N_10463,N_9925,N_9666);
or U10464 (N_10464,N_9565,N_9568);
xnor U10465 (N_10465,N_9791,N_9830);
nor U10466 (N_10466,N_9592,N_9699);
or U10467 (N_10467,N_9769,N_9546);
xnor U10468 (N_10468,N_9751,N_9703);
nor U10469 (N_10469,N_9629,N_9530);
nand U10470 (N_10470,N_9751,N_9860);
and U10471 (N_10471,N_9860,N_9768);
xnor U10472 (N_10472,N_9783,N_9941);
and U10473 (N_10473,N_9608,N_9751);
nand U10474 (N_10474,N_9501,N_9712);
nand U10475 (N_10475,N_9953,N_9579);
or U10476 (N_10476,N_9700,N_9526);
nand U10477 (N_10477,N_9567,N_9842);
and U10478 (N_10478,N_9777,N_9724);
nand U10479 (N_10479,N_9915,N_9621);
and U10480 (N_10480,N_9551,N_9507);
and U10481 (N_10481,N_9736,N_9692);
nand U10482 (N_10482,N_9980,N_9978);
xnor U10483 (N_10483,N_9876,N_9950);
or U10484 (N_10484,N_9833,N_9672);
and U10485 (N_10485,N_9825,N_9503);
nor U10486 (N_10486,N_9635,N_9873);
xor U10487 (N_10487,N_9629,N_9992);
xor U10488 (N_10488,N_9564,N_9986);
and U10489 (N_10489,N_9740,N_9771);
nor U10490 (N_10490,N_9570,N_9639);
nor U10491 (N_10491,N_9942,N_9888);
nor U10492 (N_10492,N_9848,N_9905);
and U10493 (N_10493,N_9960,N_9835);
xnor U10494 (N_10494,N_9594,N_9776);
xnor U10495 (N_10495,N_9708,N_9681);
or U10496 (N_10496,N_9574,N_9949);
nor U10497 (N_10497,N_9978,N_9930);
or U10498 (N_10498,N_9730,N_9860);
nand U10499 (N_10499,N_9627,N_9721);
and U10500 (N_10500,N_10371,N_10335);
nand U10501 (N_10501,N_10245,N_10295);
nand U10502 (N_10502,N_10006,N_10142);
nor U10503 (N_10503,N_10201,N_10067);
and U10504 (N_10504,N_10186,N_10499);
xor U10505 (N_10505,N_10431,N_10430);
or U10506 (N_10506,N_10450,N_10210);
or U10507 (N_10507,N_10372,N_10265);
nor U10508 (N_10508,N_10158,N_10133);
and U10509 (N_10509,N_10338,N_10438);
nand U10510 (N_10510,N_10051,N_10012);
xor U10511 (N_10511,N_10028,N_10079);
and U10512 (N_10512,N_10283,N_10428);
nor U10513 (N_10513,N_10345,N_10364);
or U10514 (N_10514,N_10030,N_10073);
nor U10515 (N_10515,N_10203,N_10426);
nand U10516 (N_10516,N_10026,N_10437);
xor U10517 (N_10517,N_10064,N_10116);
nor U10518 (N_10518,N_10417,N_10191);
and U10519 (N_10519,N_10358,N_10395);
xor U10520 (N_10520,N_10149,N_10435);
xor U10521 (N_10521,N_10241,N_10134);
or U10522 (N_10522,N_10069,N_10071);
and U10523 (N_10523,N_10453,N_10488);
or U10524 (N_10524,N_10369,N_10261);
or U10525 (N_10525,N_10192,N_10167);
and U10526 (N_10526,N_10316,N_10083);
xnor U10527 (N_10527,N_10093,N_10443);
or U10528 (N_10528,N_10301,N_10224);
or U10529 (N_10529,N_10419,N_10234);
nor U10530 (N_10530,N_10282,N_10185);
nor U10531 (N_10531,N_10470,N_10042);
nand U10532 (N_10532,N_10127,N_10351);
xnor U10533 (N_10533,N_10378,N_10180);
and U10534 (N_10534,N_10065,N_10289);
xnor U10535 (N_10535,N_10412,N_10441);
xor U10536 (N_10536,N_10390,N_10409);
and U10537 (N_10537,N_10498,N_10009);
or U10538 (N_10538,N_10125,N_10355);
nor U10539 (N_10539,N_10477,N_10005);
nand U10540 (N_10540,N_10015,N_10476);
or U10541 (N_10541,N_10198,N_10161);
or U10542 (N_10542,N_10175,N_10264);
and U10543 (N_10543,N_10494,N_10197);
and U10544 (N_10544,N_10391,N_10056);
or U10545 (N_10545,N_10460,N_10243);
xor U10546 (N_10546,N_10341,N_10023);
xnor U10547 (N_10547,N_10250,N_10456);
nor U10548 (N_10548,N_10052,N_10278);
nand U10549 (N_10549,N_10220,N_10445);
and U10550 (N_10550,N_10034,N_10074);
or U10551 (N_10551,N_10209,N_10386);
xnor U10552 (N_10552,N_10043,N_10267);
nor U10553 (N_10553,N_10266,N_10483);
or U10554 (N_10554,N_10287,N_10454);
or U10555 (N_10555,N_10270,N_10200);
and U10556 (N_10556,N_10085,N_10002);
nor U10557 (N_10557,N_10379,N_10318);
or U10558 (N_10558,N_10172,N_10084);
nor U10559 (N_10559,N_10121,N_10407);
and U10560 (N_10560,N_10225,N_10478);
nand U10561 (N_10561,N_10076,N_10060);
and U10562 (N_10562,N_10216,N_10370);
and U10563 (N_10563,N_10362,N_10349);
xnor U10564 (N_10564,N_10434,N_10162);
nand U10565 (N_10565,N_10296,N_10157);
and U10566 (N_10566,N_10096,N_10363);
or U10567 (N_10567,N_10276,N_10202);
nand U10568 (N_10568,N_10174,N_10353);
and U10569 (N_10569,N_10336,N_10377);
or U10570 (N_10570,N_10360,N_10022);
or U10571 (N_10571,N_10080,N_10277);
or U10572 (N_10572,N_10179,N_10217);
xnor U10573 (N_10573,N_10306,N_10122);
nor U10574 (N_10574,N_10422,N_10410);
nand U10575 (N_10575,N_10135,N_10465);
and U10576 (N_10576,N_10115,N_10150);
or U10577 (N_10577,N_10100,N_10144);
nand U10578 (N_10578,N_10236,N_10053);
nand U10579 (N_10579,N_10413,N_10485);
nand U10580 (N_10580,N_10469,N_10467);
xnor U10581 (N_10581,N_10048,N_10258);
xnor U10582 (N_10582,N_10061,N_10229);
xnor U10583 (N_10583,N_10111,N_10082);
xor U10584 (N_10584,N_10094,N_10109);
or U10585 (N_10585,N_10331,N_10442);
nor U10586 (N_10586,N_10151,N_10171);
or U10587 (N_10587,N_10021,N_10031);
xnor U10588 (N_10588,N_10325,N_10046);
nor U10589 (N_10589,N_10447,N_10350);
or U10590 (N_10590,N_10457,N_10000);
and U10591 (N_10591,N_10237,N_10376);
nor U10592 (N_10592,N_10466,N_10184);
nor U10593 (N_10593,N_10455,N_10105);
nor U10594 (N_10594,N_10248,N_10346);
or U10595 (N_10595,N_10177,N_10327);
and U10596 (N_10596,N_10029,N_10472);
xnor U10597 (N_10597,N_10078,N_10130);
nand U10598 (N_10598,N_10156,N_10496);
xnor U10599 (N_10599,N_10054,N_10396);
or U10600 (N_10600,N_10070,N_10168);
and U10601 (N_10601,N_10380,N_10219);
and U10602 (N_10602,N_10152,N_10155);
xor U10603 (N_10603,N_10050,N_10285);
xnor U10604 (N_10604,N_10032,N_10420);
or U10605 (N_10605,N_10092,N_10057);
nand U10606 (N_10606,N_10354,N_10401);
or U10607 (N_10607,N_10439,N_10309);
xnor U10608 (N_10608,N_10193,N_10091);
nor U10609 (N_10609,N_10400,N_10367);
nand U10610 (N_10610,N_10406,N_10062);
nor U10611 (N_10611,N_10044,N_10313);
and U10612 (N_10612,N_10408,N_10337);
or U10613 (N_10613,N_10486,N_10464);
xor U10614 (N_10614,N_10249,N_10039);
and U10615 (N_10615,N_10275,N_10113);
nand U10616 (N_10616,N_10387,N_10329);
nand U10617 (N_10617,N_10189,N_10007);
and U10618 (N_10618,N_10238,N_10099);
nor U10619 (N_10619,N_10104,N_10246);
nand U10620 (N_10620,N_10356,N_10231);
or U10621 (N_10621,N_10024,N_10001);
or U10622 (N_10622,N_10359,N_10211);
nand U10623 (N_10623,N_10132,N_10473);
and U10624 (N_10624,N_10374,N_10147);
and U10625 (N_10625,N_10286,N_10047);
nor U10626 (N_10626,N_10214,N_10291);
and U10627 (N_10627,N_10187,N_10199);
nor U10628 (N_10628,N_10223,N_10148);
nand U10629 (N_10629,N_10041,N_10206);
nor U10630 (N_10630,N_10143,N_10178);
xnor U10631 (N_10631,N_10230,N_10452);
and U10632 (N_10632,N_10288,N_10448);
and U10633 (N_10633,N_10242,N_10305);
or U10634 (N_10634,N_10108,N_10205);
nand U10635 (N_10635,N_10375,N_10268);
xnor U10636 (N_10636,N_10361,N_10011);
or U10637 (N_10637,N_10495,N_10257);
nand U10638 (N_10638,N_10321,N_10089);
nor U10639 (N_10639,N_10424,N_10118);
nand U10640 (N_10640,N_10339,N_10036);
nand U10641 (N_10641,N_10415,N_10497);
or U10642 (N_10642,N_10344,N_10433);
or U10643 (N_10643,N_10310,N_10263);
xnor U10644 (N_10644,N_10117,N_10418);
nand U10645 (N_10645,N_10357,N_10019);
nor U10646 (N_10646,N_10397,N_10239);
xnor U10647 (N_10647,N_10013,N_10394);
and U10648 (N_10648,N_10416,N_10334);
or U10649 (N_10649,N_10482,N_10342);
nand U10650 (N_10650,N_10131,N_10468);
or U10651 (N_10651,N_10228,N_10163);
xor U10652 (N_10652,N_10256,N_10181);
and U10653 (N_10653,N_10382,N_10146);
xnor U10654 (N_10654,N_10110,N_10173);
and U10655 (N_10655,N_10008,N_10385);
or U10656 (N_10656,N_10055,N_10490);
and U10657 (N_10657,N_10294,N_10253);
nor U10658 (N_10658,N_10269,N_10399);
and U10659 (N_10659,N_10004,N_10095);
nand U10660 (N_10660,N_10381,N_10204);
nor U10661 (N_10661,N_10451,N_10479);
nand U10662 (N_10662,N_10170,N_10293);
and U10663 (N_10663,N_10087,N_10302);
and U10664 (N_10664,N_10059,N_10440);
or U10665 (N_10665,N_10492,N_10058);
xnor U10666 (N_10666,N_10014,N_10402);
nor U10667 (N_10667,N_10398,N_10368);
xor U10668 (N_10668,N_10255,N_10297);
xor U10669 (N_10669,N_10075,N_10190);
or U10670 (N_10670,N_10033,N_10328);
and U10671 (N_10671,N_10040,N_10112);
or U10672 (N_10672,N_10195,N_10025);
nor U10673 (N_10673,N_10352,N_10481);
nand U10674 (N_10674,N_10326,N_10348);
nor U10675 (N_10675,N_10347,N_10252);
and U10676 (N_10676,N_10102,N_10388);
or U10677 (N_10677,N_10366,N_10303);
xor U10678 (N_10678,N_10323,N_10487);
nor U10679 (N_10679,N_10273,N_10218);
and U10680 (N_10680,N_10254,N_10188);
and U10681 (N_10681,N_10081,N_10298);
or U10682 (N_10682,N_10279,N_10153);
nor U10683 (N_10683,N_10165,N_10103);
nor U10684 (N_10684,N_10429,N_10123);
nor U10685 (N_10685,N_10090,N_10383);
or U10686 (N_10686,N_10129,N_10307);
or U10687 (N_10687,N_10137,N_10097);
xnor U10688 (N_10688,N_10314,N_10140);
or U10689 (N_10689,N_10027,N_10427);
or U10690 (N_10690,N_10471,N_10232);
and U10691 (N_10691,N_10221,N_10333);
or U10692 (N_10692,N_10101,N_10458);
or U10693 (N_10693,N_10425,N_10141);
and U10694 (N_10694,N_10207,N_10304);
or U10695 (N_10695,N_10045,N_10183);
xor U10696 (N_10696,N_10444,N_10423);
nand U10697 (N_10697,N_10139,N_10077);
xnor U10698 (N_10698,N_10322,N_10330);
and U10699 (N_10699,N_10324,N_10365);
xnor U10700 (N_10700,N_10068,N_10475);
nand U10701 (N_10701,N_10421,N_10284);
xnor U10702 (N_10702,N_10405,N_10119);
nor U10703 (N_10703,N_10393,N_10160);
and U10704 (N_10704,N_10213,N_10145);
xor U10705 (N_10705,N_10020,N_10138);
nand U10706 (N_10706,N_10340,N_10164);
xnor U10707 (N_10707,N_10280,N_10315);
or U10708 (N_10708,N_10066,N_10154);
xnor U10709 (N_10709,N_10226,N_10262);
and U10710 (N_10710,N_10251,N_10194);
xor U10711 (N_10711,N_10403,N_10126);
xnor U10712 (N_10712,N_10461,N_10493);
and U10713 (N_10713,N_10235,N_10392);
and U10714 (N_10714,N_10247,N_10389);
nor U10715 (N_10715,N_10271,N_10244);
nor U10716 (N_10716,N_10332,N_10107);
or U10717 (N_10717,N_10016,N_10136);
nor U10718 (N_10718,N_10292,N_10449);
and U10719 (N_10719,N_10233,N_10159);
and U10720 (N_10720,N_10018,N_10035);
nor U10721 (N_10721,N_10459,N_10088);
nand U10722 (N_10722,N_10484,N_10373);
xor U10723 (N_10723,N_10196,N_10300);
nor U10724 (N_10724,N_10259,N_10227);
nor U10725 (N_10725,N_10072,N_10462);
nor U10726 (N_10726,N_10208,N_10446);
xnor U10727 (N_10727,N_10114,N_10176);
xor U10728 (N_10728,N_10272,N_10240);
nand U10729 (N_10729,N_10463,N_10049);
nor U10730 (N_10730,N_10308,N_10166);
and U10731 (N_10731,N_10124,N_10299);
and U10732 (N_10732,N_10003,N_10290);
nand U10733 (N_10733,N_10384,N_10274);
and U10734 (N_10734,N_10281,N_10086);
nor U10735 (N_10735,N_10320,N_10063);
or U10736 (N_10736,N_10480,N_10432);
or U10737 (N_10737,N_10489,N_10474);
or U10738 (N_10738,N_10317,N_10017);
xnor U10739 (N_10739,N_10010,N_10260);
nor U10740 (N_10740,N_10212,N_10106);
nand U10741 (N_10741,N_10120,N_10343);
and U10742 (N_10742,N_10128,N_10169);
xor U10743 (N_10743,N_10319,N_10311);
xor U10744 (N_10744,N_10037,N_10411);
and U10745 (N_10745,N_10215,N_10436);
xnor U10746 (N_10746,N_10491,N_10404);
nand U10747 (N_10747,N_10098,N_10414);
nand U10748 (N_10748,N_10312,N_10038);
or U10749 (N_10749,N_10182,N_10222);
xnor U10750 (N_10750,N_10073,N_10439);
or U10751 (N_10751,N_10244,N_10461);
xor U10752 (N_10752,N_10336,N_10313);
nand U10753 (N_10753,N_10401,N_10443);
nand U10754 (N_10754,N_10350,N_10096);
xor U10755 (N_10755,N_10173,N_10373);
nand U10756 (N_10756,N_10400,N_10283);
or U10757 (N_10757,N_10108,N_10483);
and U10758 (N_10758,N_10212,N_10427);
nor U10759 (N_10759,N_10089,N_10322);
or U10760 (N_10760,N_10143,N_10033);
xor U10761 (N_10761,N_10448,N_10156);
xor U10762 (N_10762,N_10191,N_10030);
or U10763 (N_10763,N_10122,N_10440);
nor U10764 (N_10764,N_10079,N_10440);
nand U10765 (N_10765,N_10291,N_10481);
xor U10766 (N_10766,N_10234,N_10393);
nand U10767 (N_10767,N_10197,N_10474);
xnor U10768 (N_10768,N_10009,N_10079);
nand U10769 (N_10769,N_10194,N_10071);
and U10770 (N_10770,N_10246,N_10072);
nor U10771 (N_10771,N_10152,N_10334);
nor U10772 (N_10772,N_10309,N_10117);
xnor U10773 (N_10773,N_10131,N_10028);
nor U10774 (N_10774,N_10356,N_10246);
nand U10775 (N_10775,N_10338,N_10157);
nand U10776 (N_10776,N_10246,N_10070);
xor U10777 (N_10777,N_10297,N_10090);
nor U10778 (N_10778,N_10460,N_10462);
xor U10779 (N_10779,N_10236,N_10267);
xnor U10780 (N_10780,N_10125,N_10476);
and U10781 (N_10781,N_10258,N_10406);
nand U10782 (N_10782,N_10067,N_10332);
nor U10783 (N_10783,N_10019,N_10340);
nor U10784 (N_10784,N_10344,N_10273);
nor U10785 (N_10785,N_10176,N_10102);
nand U10786 (N_10786,N_10183,N_10390);
or U10787 (N_10787,N_10395,N_10332);
and U10788 (N_10788,N_10421,N_10093);
or U10789 (N_10789,N_10447,N_10204);
nor U10790 (N_10790,N_10401,N_10130);
and U10791 (N_10791,N_10496,N_10492);
and U10792 (N_10792,N_10106,N_10319);
nand U10793 (N_10793,N_10168,N_10248);
nand U10794 (N_10794,N_10258,N_10316);
or U10795 (N_10795,N_10206,N_10453);
nand U10796 (N_10796,N_10378,N_10117);
nor U10797 (N_10797,N_10277,N_10005);
xnor U10798 (N_10798,N_10037,N_10045);
nand U10799 (N_10799,N_10441,N_10293);
xor U10800 (N_10800,N_10184,N_10083);
or U10801 (N_10801,N_10194,N_10012);
or U10802 (N_10802,N_10257,N_10068);
or U10803 (N_10803,N_10106,N_10139);
nor U10804 (N_10804,N_10398,N_10401);
or U10805 (N_10805,N_10392,N_10287);
nor U10806 (N_10806,N_10464,N_10123);
nand U10807 (N_10807,N_10018,N_10229);
or U10808 (N_10808,N_10109,N_10431);
nand U10809 (N_10809,N_10131,N_10390);
xor U10810 (N_10810,N_10046,N_10085);
nand U10811 (N_10811,N_10462,N_10433);
xnor U10812 (N_10812,N_10270,N_10297);
xnor U10813 (N_10813,N_10443,N_10067);
or U10814 (N_10814,N_10154,N_10030);
nor U10815 (N_10815,N_10159,N_10065);
nand U10816 (N_10816,N_10483,N_10128);
xnor U10817 (N_10817,N_10287,N_10497);
and U10818 (N_10818,N_10208,N_10365);
nand U10819 (N_10819,N_10279,N_10090);
nand U10820 (N_10820,N_10449,N_10163);
nand U10821 (N_10821,N_10367,N_10369);
and U10822 (N_10822,N_10207,N_10488);
xnor U10823 (N_10823,N_10260,N_10088);
nand U10824 (N_10824,N_10149,N_10196);
and U10825 (N_10825,N_10076,N_10329);
and U10826 (N_10826,N_10444,N_10078);
or U10827 (N_10827,N_10355,N_10415);
or U10828 (N_10828,N_10376,N_10329);
xor U10829 (N_10829,N_10294,N_10197);
or U10830 (N_10830,N_10236,N_10383);
xnor U10831 (N_10831,N_10437,N_10057);
or U10832 (N_10832,N_10402,N_10095);
or U10833 (N_10833,N_10042,N_10278);
or U10834 (N_10834,N_10031,N_10380);
xor U10835 (N_10835,N_10055,N_10179);
nand U10836 (N_10836,N_10068,N_10225);
or U10837 (N_10837,N_10300,N_10128);
nor U10838 (N_10838,N_10470,N_10025);
nor U10839 (N_10839,N_10011,N_10126);
nor U10840 (N_10840,N_10464,N_10473);
and U10841 (N_10841,N_10276,N_10489);
nand U10842 (N_10842,N_10270,N_10363);
or U10843 (N_10843,N_10022,N_10207);
and U10844 (N_10844,N_10182,N_10401);
xnor U10845 (N_10845,N_10102,N_10188);
or U10846 (N_10846,N_10448,N_10415);
or U10847 (N_10847,N_10405,N_10096);
or U10848 (N_10848,N_10175,N_10393);
nor U10849 (N_10849,N_10492,N_10296);
nor U10850 (N_10850,N_10455,N_10442);
or U10851 (N_10851,N_10083,N_10467);
xor U10852 (N_10852,N_10088,N_10342);
xor U10853 (N_10853,N_10210,N_10106);
xnor U10854 (N_10854,N_10043,N_10019);
and U10855 (N_10855,N_10485,N_10162);
and U10856 (N_10856,N_10360,N_10209);
nand U10857 (N_10857,N_10221,N_10380);
nor U10858 (N_10858,N_10452,N_10402);
xnor U10859 (N_10859,N_10248,N_10005);
or U10860 (N_10860,N_10118,N_10308);
nor U10861 (N_10861,N_10225,N_10117);
nor U10862 (N_10862,N_10310,N_10456);
and U10863 (N_10863,N_10454,N_10330);
and U10864 (N_10864,N_10201,N_10163);
nor U10865 (N_10865,N_10012,N_10019);
or U10866 (N_10866,N_10199,N_10246);
and U10867 (N_10867,N_10321,N_10412);
nand U10868 (N_10868,N_10366,N_10258);
xor U10869 (N_10869,N_10288,N_10261);
nand U10870 (N_10870,N_10115,N_10151);
nand U10871 (N_10871,N_10493,N_10393);
nand U10872 (N_10872,N_10458,N_10494);
nor U10873 (N_10873,N_10349,N_10368);
xnor U10874 (N_10874,N_10130,N_10259);
nor U10875 (N_10875,N_10430,N_10366);
xor U10876 (N_10876,N_10284,N_10376);
or U10877 (N_10877,N_10435,N_10364);
nor U10878 (N_10878,N_10286,N_10014);
or U10879 (N_10879,N_10351,N_10188);
xor U10880 (N_10880,N_10161,N_10099);
or U10881 (N_10881,N_10416,N_10452);
nand U10882 (N_10882,N_10326,N_10347);
and U10883 (N_10883,N_10409,N_10448);
and U10884 (N_10884,N_10168,N_10091);
and U10885 (N_10885,N_10367,N_10370);
nand U10886 (N_10886,N_10351,N_10363);
and U10887 (N_10887,N_10179,N_10224);
or U10888 (N_10888,N_10041,N_10166);
nor U10889 (N_10889,N_10062,N_10218);
nor U10890 (N_10890,N_10094,N_10122);
or U10891 (N_10891,N_10317,N_10241);
or U10892 (N_10892,N_10459,N_10241);
or U10893 (N_10893,N_10321,N_10315);
nand U10894 (N_10894,N_10083,N_10078);
or U10895 (N_10895,N_10164,N_10467);
xor U10896 (N_10896,N_10158,N_10003);
or U10897 (N_10897,N_10430,N_10497);
or U10898 (N_10898,N_10045,N_10380);
and U10899 (N_10899,N_10370,N_10365);
and U10900 (N_10900,N_10384,N_10423);
nor U10901 (N_10901,N_10159,N_10034);
xnor U10902 (N_10902,N_10338,N_10238);
nand U10903 (N_10903,N_10032,N_10418);
and U10904 (N_10904,N_10151,N_10235);
nand U10905 (N_10905,N_10489,N_10464);
or U10906 (N_10906,N_10158,N_10295);
or U10907 (N_10907,N_10316,N_10211);
or U10908 (N_10908,N_10395,N_10388);
xor U10909 (N_10909,N_10271,N_10289);
nor U10910 (N_10910,N_10248,N_10151);
and U10911 (N_10911,N_10431,N_10195);
or U10912 (N_10912,N_10112,N_10041);
xor U10913 (N_10913,N_10287,N_10171);
nor U10914 (N_10914,N_10463,N_10222);
nor U10915 (N_10915,N_10155,N_10440);
nand U10916 (N_10916,N_10458,N_10440);
xor U10917 (N_10917,N_10409,N_10433);
or U10918 (N_10918,N_10329,N_10321);
xor U10919 (N_10919,N_10255,N_10366);
and U10920 (N_10920,N_10158,N_10449);
and U10921 (N_10921,N_10473,N_10161);
xnor U10922 (N_10922,N_10384,N_10157);
xnor U10923 (N_10923,N_10261,N_10344);
nand U10924 (N_10924,N_10057,N_10064);
xnor U10925 (N_10925,N_10270,N_10295);
and U10926 (N_10926,N_10473,N_10216);
or U10927 (N_10927,N_10136,N_10121);
nand U10928 (N_10928,N_10294,N_10018);
xnor U10929 (N_10929,N_10451,N_10099);
xnor U10930 (N_10930,N_10160,N_10240);
nor U10931 (N_10931,N_10444,N_10362);
nand U10932 (N_10932,N_10222,N_10487);
xor U10933 (N_10933,N_10280,N_10240);
and U10934 (N_10934,N_10067,N_10255);
xnor U10935 (N_10935,N_10221,N_10070);
or U10936 (N_10936,N_10156,N_10336);
xnor U10937 (N_10937,N_10375,N_10395);
nand U10938 (N_10938,N_10295,N_10496);
xnor U10939 (N_10939,N_10494,N_10191);
nand U10940 (N_10940,N_10204,N_10234);
and U10941 (N_10941,N_10005,N_10489);
and U10942 (N_10942,N_10116,N_10348);
or U10943 (N_10943,N_10458,N_10000);
xnor U10944 (N_10944,N_10367,N_10309);
or U10945 (N_10945,N_10066,N_10100);
nor U10946 (N_10946,N_10430,N_10488);
and U10947 (N_10947,N_10288,N_10433);
nand U10948 (N_10948,N_10198,N_10478);
or U10949 (N_10949,N_10200,N_10429);
nor U10950 (N_10950,N_10341,N_10396);
or U10951 (N_10951,N_10151,N_10212);
or U10952 (N_10952,N_10149,N_10256);
nor U10953 (N_10953,N_10368,N_10300);
and U10954 (N_10954,N_10183,N_10472);
nand U10955 (N_10955,N_10068,N_10098);
nor U10956 (N_10956,N_10367,N_10139);
nand U10957 (N_10957,N_10357,N_10186);
and U10958 (N_10958,N_10271,N_10389);
nor U10959 (N_10959,N_10071,N_10055);
nor U10960 (N_10960,N_10381,N_10358);
nand U10961 (N_10961,N_10063,N_10412);
xnor U10962 (N_10962,N_10118,N_10301);
and U10963 (N_10963,N_10254,N_10343);
nor U10964 (N_10964,N_10012,N_10246);
nor U10965 (N_10965,N_10087,N_10462);
xor U10966 (N_10966,N_10345,N_10331);
xnor U10967 (N_10967,N_10368,N_10125);
or U10968 (N_10968,N_10123,N_10062);
nor U10969 (N_10969,N_10317,N_10134);
nor U10970 (N_10970,N_10348,N_10022);
nor U10971 (N_10971,N_10124,N_10094);
nor U10972 (N_10972,N_10253,N_10072);
or U10973 (N_10973,N_10177,N_10382);
xor U10974 (N_10974,N_10484,N_10080);
xnor U10975 (N_10975,N_10405,N_10033);
nor U10976 (N_10976,N_10394,N_10154);
xnor U10977 (N_10977,N_10431,N_10416);
or U10978 (N_10978,N_10179,N_10047);
or U10979 (N_10979,N_10374,N_10492);
nor U10980 (N_10980,N_10304,N_10049);
or U10981 (N_10981,N_10149,N_10344);
and U10982 (N_10982,N_10447,N_10095);
and U10983 (N_10983,N_10166,N_10342);
and U10984 (N_10984,N_10035,N_10225);
xor U10985 (N_10985,N_10344,N_10439);
nand U10986 (N_10986,N_10032,N_10067);
nand U10987 (N_10987,N_10287,N_10272);
nor U10988 (N_10988,N_10182,N_10405);
xnor U10989 (N_10989,N_10222,N_10113);
and U10990 (N_10990,N_10345,N_10154);
nand U10991 (N_10991,N_10020,N_10005);
and U10992 (N_10992,N_10201,N_10216);
or U10993 (N_10993,N_10163,N_10082);
xor U10994 (N_10994,N_10386,N_10210);
nor U10995 (N_10995,N_10454,N_10044);
nor U10996 (N_10996,N_10021,N_10257);
and U10997 (N_10997,N_10210,N_10434);
or U10998 (N_10998,N_10223,N_10438);
and U10999 (N_10999,N_10208,N_10294);
xnor U11000 (N_11000,N_10680,N_10940);
nor U11001 (N_11001,N_10743,N_10722);
nor U11002 (N_11002,N_10922,N_10591);
nand U11003 (N_11003,N_10965,N_10769);
or U11004 (N_11004,N_10634,N_10828);
nand U11005 (N_11005,N_10737,N_10970);
nand U11006 (N_11006,N_10806,N_10555);
and U11007 (N_11007,N_10839,N_10520);
and U11008 (N_11008,N_10625,N_10945);
and U11009 (N_11009,N_10862,N_10985);
nand U11010 (N_11010,N_10919,N_10647);
or U11011 (N_11011,N_10502,N_10579);
nand U11012 (N_11012,N_10646,N_10780);
or U11013 (N_11013,N_10913,N_10611);
nand U11014 (N_11014,N_10799,N_10650);
or U11015 (N_11015,N_10954,N_10800);
nor U11016 (N_11016,N_10939,N_10918);
and U11017 (N_11017,N_10716,N_10968);
xor U11018 (N_11018,N_10717,N_10869);
and U11019 (N_11019,N_10648,N_10884);
or U11020 (N_11020,N_10896,N_10760);
nand U11021 (N_11021,N_10691,N_10866);
xnor U11022 (N_11022,N_10908,N_10997);
nand U11023 (N_11023,N_10781,N_10524);
and U11024 (N_11024,N_10629,N_10802);
nand U11025 (N_11025,N_10912,N_10926);
xor U11026 (N_11026,N_10563,N_10885);
and U11027 (N_11027,N_10715,N_10888);
nor U11028 (N_11028,N_10552,N_10775);
nand U11029 (N_11029,N_10515,N_10533);
nand U11030 (N_11030,N_10557,N_10822);
and U11031 (N_11031,N_10607,N_10641);
or U11032 (N_11032,N_10543,N_10957);
xnor U11033 (N_11033,N_10794,N_10617);
xor U11034 (N_11034,N_10952,N_10848);
or U11035 (N_11035,N_10695,N_10897);
and U11036 (N_11036,N_10675,N_10793);
or U11037 (N_11037,N_10705,N_10724);
xnor U11038 (N_11038,N_10678,N_10924);
nand U11039 (N_11039,N_10521,N_10854);
nand U11040 (N_11040,N_10774,N_10701);
xor U11041 (N_11041,N_10762,N_10654);
nor U11042 (N_11042,N_10993,N_10895);
nand U11043 (N_11043,N_10714,N_10796);
xnor U11044 (N_11044,N_10636,N_10829);
or U11045 (N_11045,N_10811,N_10728);
and U11046 (N_11046,N_10766,N_10645);
nand U11047 (N_11047,N_10910,N_10596);
or U11048 (N_11048,N_10668,N_10528);
or U11049 (N_11049,N_10711,N_10682);
nor U11050 (N_11050,N_10814,N_10783);
nand U11051 (N_11051,N_10981,N_10638);
xor U11052 (N_11052,N_10972,N_10577);
xnor U11053 (N_11053,N_10601,N_10523);
nor U11054 (N_11054,N_10891,N_10764);
or U11055 (N_11055,N_10843,N_10999);
nor U11056 (N_11056,N_10619,N_10580);
and U11057 (N_11057,N_10827,N_10748);
nor U11058 (N_11058,N_10730,N_10639);
and U11059 (N_11059,N_10697,N_10545);
and U11060 (N_11060,N_10944,N_10739);
and U11061 (N_11061,N_10670,N_10816);
nand U11062 (N_11062,N_10627,N_10672);
or U11063 (N_11063,N_10784,N_10534);
and U11064 (N_11064,N_10558,N_10763);
nor U11065 (N_11065,N_10902,N_10674);
nand U11066 (N_11066,N_10978,N_10798);
nor U11067 (N_11067,N_10614,N_10556);
xnor U11068 (N_11068,N_10637,N_10538);
xor U11069 (N_11069,N_10589,N_10905);
nor U11070 (N_11070,N_10621,N_10788);
or U11071 (N_11071,N_10504,N_10583);
nand U11072 (N_11072,N_10566,N_10805);
and U11073 (N_11073,N_10966,N_10842);
or U11074 (N_11074,N_10947,N_10809);
xor U11075 (N_11075,N_10786,N_10911);
nand U11076 (N_11076,N_10610,N_10688);
nor U11077 (N_11077,N_10958,N_10626);
nand U11078 (N_11078,N_10928,N_10936);
xor U11079 (N_11079,N_10850,N_10801);
nand U11080 (N_11080,N_10880,N_10946);
and U11081 (N_11081,N_10852,N_10853);
or U11082 (N_11082,N_10628,N_10770);
and U11083 (N_11083,N_10804,N_10949);
nand U11084 (N_11084,N_10667,N_10747);
or U11085 (N_11085,N_10980,N_10676);
xor U11086 (N_11086,N_10643,N_10756);
or U11087 (N_11087,N_10588,N_10740);
xnor U11088 (N_11088,N_10785,N_10567);
nand U11089 (N_11089,N_10983,N_10530);
xnor U11090 (N_11090,N_10883,N_10511);
nor U11091 (N_11091,N_10642,N_10597);
nor U11092 (N_11092,N_10584,N_10787);
nor U11093 (N_11093,N_10903,N_10974);
nand U11094 (N_11094,N_10844,N_10677);
nand U11095 (N_11095,N_10967,N_10706);
nand U11096 (N_11096,N_10909,N_10878);
xor U11097 (N_11097,N_10821,N_10734);
and U11098 (N_11098,N_10603,N_10573);
nand U11099 (N_11099,N_10778,N_10693);
nor U11100 (N_11100,N_10679,N_10516);
nor U11101 (N_11101,N_10602,N_10624);
nand U11102 (N_11102,N_10548,N_10605);
nand U11103 (N_11103,N_10824,N_10574);
or U11104 (N_11104,N_10535,N_10586);
nor U11105 (N_11105,N_10700,N_10790);
or U11106 (N_11106,N_10731,N_10810);
xor U11107 (N_11107,N_10640,N_10836);
nand U11108 (N_11108,N_10592,N_10518);
nand U11109 (N_11109,N_10750,N_10789);
nand U11110 (N_11110,N_10633,N_10820);
xor U11111 (N_11111,N_10735,N_10559);
and U11112 (N_11112,N_10941,N_10501);
nor U11113 (N_11113,N_10873,N_10698);
xnor U11114 (N_11114,N_10808,N_10560);
or U11115 (N_11115,N_10608,N_10898);
nand U11116 (N_11116,N_10948,N_10998);
or U11117 (N_11117,N_10917,N_10719);
xor U11118 (N_11118,N_10582,N_10525);
or U11119 (N_11119,N_10595,N_10660);
nand U11120 (N_11120,N_10522,N_10777);
or U11121 (N_11121,N_10835,N_10819);
and U11122 (N_11122,N_10925,N_10510);
and U11123 (N_11123,N_10553,N_10606);
or U11124 (N_11124,N_10581,N_10609);
or U11125 (N_11125,N_10632,N_10791);
nand U11126 (N_11126,N_10539,N_10702);
nand U11127 (N_11127,N_10565,N_10755);
and U11128 (N_11128,N_10673,N_10823);
nor U11129 (N_11129,N_10870,N_10877);
xnor U11130 (N_11130,N_10933,N_10865);
or U11131 (N_11131,N_10613,N_10507);
and U11132 (N_11132,N_10761,N_10527);
nand U11133 (N_11133,N_10838,N_10532);
and U11134 (N_11134,N_10568,N_10593);
nor U11135 (N_11135,N_10860,N_10961);
and U11136 (N_11136,N_10564,N_10859);
xor U11137 (N_11137,N_10686,N_10951);
xnor U11138 (N_11138,N_10807,N_10635);
nand U11139 (N_11139,N_10841,N_10846);
nor U11140 (N_11140,N_10694,N_10631);
xnor U11141 (N_11141,N_10547,N_10696);
or U11142 (N_11142,N_10749,N_10585);
or U11143 (N_11143,N_10973,N_10955);
and U11144 (N_11144,N_10754,N_10669);
xnor U11145 (N_11145,N_10540,N_10868);
and U11146 (N_11146,N_10704,N_10962);
and U11147 (N_11147,N_10817,N_10757);
xor U11148 (N_11148,N_10689,N_10847);
xnor U11149 (N_11149,N_10834,N_10923);
xor U11150 (N_11150,N_10622,N_10832);
nor U11151 (N_11151,N_10773,N_10707);
and U11152 (N_11152,N_10906,N_10746);
xor U11153 (N_11153,N_10992,N_10879);
nand U11154 (N_11154,N_10792,N_10779);
or U11155 (N_11155,N_10681,N_10994);
nand U11156 (N_11156,N_10623,N_10931);
or U11157 (N_11157,N_10513,N_10765);
nor U11158 (N_11158,N_10536,N_10576);
and U11159 (N_11159,N_10709,N_10875);
xnor U11160 (N_11160,N_10971,N_10509);
nor U11161 (N_11161,N_10699,N_10901);
xnor U11162 (N_11162,N_10744,N_10512);
and U11163 (N_11163,N_10758,N_10826);
xor U11164 (N_11164,N_10503,N_10943);
nor U11165 (N_11165,N_10963,N_10658);
nand U11166 (N_11166,N_10508,N_10753);
nand U11167 (N_11167,N_10721,N_10861);
or U11168 (N_11168,N_10935,N_10818);
nand U11169 (N_11169,N_10649,N_10894);
xnor U11170 (N_11170,N_10987,N_10550);
nand U11171 (N_11171,N_10575,N_10953);
or U11172 (N_11172,N_10703,N_10690);
nor U11173 (N_11173,N_10803,N_10887);
xnor U11174 (N_11174,N_10876,N_10657);
nand U11175 (N_11175,N_10616,N_10920);
nor U11176 (N_11176,N_10687,N_10651);
nand U11177 (N_11177,N_10561,N_10914);
or U11178 (N_11178,N_10982,N_10984);
or U11179 (N_11179,N_10713,N_10988);
or U11180 (N_11180,N_10745,N_10544);
xnor U11181 (N_11181,N_10546,N_10929);
xnor U11182 (N_11182,N_10727,N_10882);
nand U11183 (N_11183,N_10812,N_10767);
xor U11184 (N_11184,N_10587,N_10813);
nor U11185 (N_11185,N_10932,N_10529);
nor U11186 (N_11186,N_10976,N_10500);
and U11187 (N_11187,N_10514,N_10708);
xnor U11188 (N_11188,N_10710,N_10692);
nand U11189 (N_11189,N_10921,N_10930);
and U11190 (N_11190,N_10618,N_10526);
nor U11191 (N_11191,N_10519,N_10892);
xnor U11192 (N_11192,N_10505,N_10975);
and U11193 (N_11193,N_10732,N_10837);
or U11194 (N_11194,N_10915,N_10831);
and U11195 (N_11195,N_10950,N_10537);
or U11196 (N_11196,N_10795,N_10578);
xnor U11197 (N_11197,N_10942,N_10927);
and U11198 (N_11198,N_10990,N_10825);
nand U11199 (N_11199,N_10517,N_10900);
or U11200 (N_11200,N_10867,N_10864);
nor U11201 (N_11201,N_10684,N_10979);
xor U11202 (N_11202,N_10886,N_10845);
nand U11203 (N_11203,N_10772,N_10652);
nor U11204 (N_11204,N_10833,N_10849);
and U11205 (N_11205,N_10815,N_10663);
nand U11206 (N_11206,N_10771,N_10549);
and U11207 (N_11207,N_10656,N_10934);
and U11208 (N_11208,N_10893,N_10570);
nand U11209 (N_11209,N_10742,N_10995);
or U11210 (N_11210,N_10594,N_10531);
and U11211 (N_11211,N_10683,N_10991);
xor U11212 (N_11212,N_10551,N_10986);
xor U11213 (N_11213,N_10907,N_10506);
nor U11214 (N_11214,N_10554,N_10653);
and U11215 (N_11215,N_10956,N_10662);
and U11216 (N_11216,N_10712,N_10644);
xnor U11217 (N_11217,N_10664,N_10797);
and U11218 (N_11218,N_10615,N_10959);
xnor U11219 (N_11219,N_10733,N_10964);
nand U11220 (N_11220,N_10720,N_10590);
or U11221 (N_11221,N_10759,N_10723);
or U11222 (N_11222,N_10612,N_10671);
xor U11223 (N_11223,N_10729,N_10572);
nor U11224 (N_11224,N_10856,N_10840);
nor U11225 (N_11225,N_10741,N_10960);
xor U11226 (N_11226,N_10881,N_10989);
and U11227 (N_11227,N_10916,N_10890);
or U11228 (N_11228,N_10855,N_10969);
nor U11229 (N_11229,N_10782,N_10666);
xor U11230 (N_11230,N_10541,N_10752);
or U11231 (N_11231,N_10661,N_10904);
nand U11232 (N_11232,N_10599,N_10751);
or U11233 (N_11233,N_10996,N_10604);
or U11234 (N_11234,N_10598,N_10665);
xnor U11235 (N_11235,N_10889,N_10871);
nand U11236 (N_11236,N_10830,N_10571);
nor U11237 (N_11237,N_10736,N_10685);
xnor U11238 (N_11238,N_10938,N_10562);
xnor U11239 (N_11239,N_10768,N_10738);
xor U11240 (N_11240,N_10600,N_10569);
and U11241 (N_11241,N_10726,N_10874);
nor U11242 (N_11242,N_10851,N_10630);
nand U11243 (N_11243,N_10857,N_10542);
or U11244 (N_11244,N_10858,N_10776);
or U11245 (N_11245,N_10655,N_10872);
or U11246 (N_11246,N_10937,N_10725);
nand U11247 (N_11247,N_10899,N_10977);
nand U11248 (N_11248,N_10659,N_10620);
nand U11249 (N_11249,N_10718,N_10863);
nor U11250 (N_11250,N_10935,N_10888);
nor U11251 (N_11251,N_10885,N_10747);
or U11252 (N_11252,N_10673,N_10666);
and U11253 (N_11253,N_10864,N_10730);
nor U11254 (N_11254,N_10582,N_10597);
xnor U11255 (N_11255,N_10817,N_10639);
or U11256 (N_11256,N_10826,N_10589);
and U11257 (N_11257,N_10576,N_10785);
and U11258 (N_11258,N_10598,N_10937);
nand U11259 (N_11259,N_10911,N_10806);
nand U11260 (N_11260,N_10578,N_10813);
xnor U11261 (N_11261,N_10533,N_10687);
nand U11262 (N_11262,N_10964,N_10987);
xor U11263 (N_11263,N_10958,N_10640);
nor U11264 (N_11264,N_10726,N_10971);
nor U11265 (N_11265,N_10688,N_10563);
and U11266 (N_11266,N_10504,N_10961);
or U11267 (N_11267,N_10900,N_10652);
nand U11268 (N_11268,N_10827,N_10595);
nand U11269 (N_11269,N_10717,N_10880);
or U11270 (N_11270,N_10604,N_10520);
nand U11271 (N_11271,N_10791,N_10594);
and U11272 (N_11272,N_10989,N_10587);
xnor U11273 (N_11273,N_10568,N_10721);
xor U11274 (N_11274,N_10781,N_10858);
nand U11275 (N_11275,N_10756,N_10689);
nor U11276 (N_11276,N_10620,N_10576);
and U11277 (N_11277,N_10719,N_10641);
nand U11278 (N_11278,N_10774,N_10987);
or U11279 (N_11279,N_10624,N_10652);
nor U11280 (N_11280,N_10733,N_10514);
and U11281 (N_11281,N_10809,N_10763);
and U11282 (N_11282,N_10636,N_10767);
and U11283 (N_11283,N_10965,N_10668);
xor U11284 (N_11284,N_10992,N_10642);
nor U11285 (N_11285,N_10567,N_10806);
xor U11286 (N_11286,N_10632,N_10947);
xor U11287 (N_11287,N_10658,N_10541);
and U11288 (N_11288,N_10889,N_10716);
nand U11289 (N_11289,N_10816,N_10922);
and U11290 (N_11290,N_10826,N_10892);
or U11291 (N_11291,N_10744,N_10815);
xor U11292 (N_11292,N_10847,N_10988);
nor U11293 (N_11293,N_10721,N_10793);
or U11294 (N_11294,N_10631,N_10897);
nor U11295 (N_11295,N_10785,N_10857);
and U11296 (N_11296,N_10667,N_10962);
or U11297 (N_11297,N_10522,N_10505);
nor U11298 (N_11298,N_10741,N_10546);
nor U11299 (N_11299,N_10880,N_10667);
nand U11300 (N_11300,N_10763,N_10697);
nor U11301 (N_11301,N_10713,N_10566);
xor U11302 (N_11302,N_10818,N_10536);
and U11303 (N_11303,N_10790,N_10512);
and U11304 (N_11304,N_10700,N_10831);
or U11305 (N_11305,N_10608,N_10858);
nor U11306 (N_11306,N_10918,N_10796);
nor U11307 (N_11307,N_10842,N_10988);
or U11308 (N_11308,N_10530,N_10768);
nand U11309 (N_11309,N_10681,N_10602);
or U11310 (N_11310,N_10744,N_10842);
or U11311 (N_11311,N_10629,N_10964);
nor U11312 (N_11312,N_10915,N_10896);
or U11313 (N_11313,N_10604,N_10778);
xor U11314 (N_11314,N_10593,N_10583);
or U11315 (N_11315,N_10779,N_10627);
nor U11316 (N_11316,N_10655,N_10563);
or U11317 (N_11317,N_10908,N_10911);
or U11318 (N_11318,N_10952,N_10950);
and U11319 (N_11319,N_10964,N_10544);
xor U11320 (N_11320,N_10787,N_10885);
nor U11321 (N_11321,N_10630,N_10560);
or U11322 (N_11322,N_10911,N_10776);
nor U11323 (N_11323,N_10771,N_10989);
and U11324 (N_11324,N_10624,N_10846);
nor U11325 (N_11325,N_10656,N_10930);
nor U11326 (N_11326,N_10631,N_10548);
xor U11327 (N_11327,N_10595,N_10518);
nor U11328 (N_11328,N_10685,N_10851);
or U11329 (N_11329,N_10774,N_10692);
xor U11330 (N_11330,N_10718,N_10699);
and U11331 (N_11331,N_10614,N_10534);
nand U11332 (N_11332,N_10861,N_10811);
nor U11333 (N_11333,N_10683,N_10865);
xnor U11334 (N_11334,N_10973,N_10902);
nor U11335 (N_11335,N_10947,N_10987);
nor U11336 (N_11336,N_10500,N_10875);
and U11337 (N_11337,N_10741,N_10711);
nor U11338 (N_11338,N_10713,N_10743);
nand U11339 (N_11339,N_10945,N_10947);
and U11340 (N_11340,N_10966,N_10684);
nand U11341 (N_11341,N_10853,N_10581);
xnor U11342 (N_11342,N_10784,N_10916);
or U11343 (N_11343,N_10922,N_10657);
nand U11344 (N_11344,N_10551,N_10959);
xor U11345 (N_11345,N_10685,N_10689);
xnor U11346 (N_11346,N_10937,N_10881);
nand U11347 (N_11347,N_10736,N_10624);
or U11348 (N_11348,N_10826,N_10582);
xor U11349 (N_11349,N_10559,N_10954);
xnor U11350 (N_11350,N_10684,N_10984);
nand U11351 (N_11351,N_10795,N_10910);
nand U11352 (N_11352,N_10678,N_10518);
nor U11353 (N_11353,N_10556,N_10780);
nor U11354 (N_11354,N_10819,N_10753);
xor U11355 (N_11355,N_10578,N_10518);
nor U11356 (N_11356,N_10816,N_10903);
nand U11357 (N_11357,N_10772,N_10936);
nor U11358 (N_11358,N_10811,N_10505);
or U11359 (N_11359,N_10597,N_10706);
xnor U11360 (N_11360,N_10973,N_10992);
xnor U11361 (N_11361,N_10529,N_10747);
and U11362 (N_11362,N_10979,N_10649);
or U11363 (N_11363,N_10943,N_10933);
or U11364 (N_11364,N_10633,N_10848);
xor U11365 (N_11365,N_10518,N_10876);
and U11366 (N_11366,N_10869,N_10753);
nand U11367 (N_11367,N_10780,N_10636);
or U11368 (N_11368,N_10986,N_10565);
and U11369 (N_11369,N_10767,N_10574);
xnor U11370 (N_11370,N_10679,N_10606);
xor U11371 (N_11371,N_10815,N_10918);
nand U11372 (N_11372,N_10684,N_10522);
nor U11373 (N_11373,N_10940,N_10581);
and U11374 (N_11374,N_10672,N_10990);
xor U11375 (N_11375,N_10765,N_10997);
nand U11376 (N_11376,N_10678,N_10625);
nor U11377 (N_11377,N_10597,N_10501);
nor U11378 (N_11378,N_10833,N_10827);
xor U11379 (N_11379,N_10683,N_10896);
nor U11380 (N_11380,N_10788,N_10714);
nand U11381 (N_11381,N_10590,N_10609);
or U11382 (N_11382,N_10684,N_10880);
nor U11383 (N_11383,N_10969,N_10808);
or U11384 (N_11384,N_10853,N_10948);
xor U11385 (N_11385,N_10988,N_10699);
or U11386 (N_11386,N_10521,N_10549);
nor U11387 (N_11387,N_10970,N_10574);
xor U11388 (N_11388,N_10718,N_10894);
or U11389 (N_11389,N_10539,N_10787);
nor U11390 (N_11390,N_10844,N_10773);
nand U11391 (N_11391,N_10852,N_10960);
nand U11392 (N_11392,N_10728,N_10659);
or U11393 (N_11393,N_10670,N_10698);
nand U11394 (N_11394,N_10673,N_10645);
nand U11395 (N_11395,N_10852,N_10826);
nand U11396 (N_11396,N_10559,N_10543);
nand U11397 (N_11397,N_10659,N_10910);
nor U11398 (N_11398,N_10519,N_10705);
xnor U11399 (N_11399,N_10578,N_10668);
nor U11400 (N_11400,N_10628,N_10555);
xnor U11401 (N_11401,N_10942,N_10722);
nand U11402 (N_11402,N_10705,N_10872);
and U11403 (N_11403,N_10751,N_10674);
xnor U11404 (N_11404,N_10818,N_10839);
xnor U11405 (N_11405,N_10842,N_10637);
nand U11406 (N_11406,N_10908,N_10701);
nor U11407 (N_11407,N_10626,N_10743);
nand U11408 (N_11408,N_10975,N_10608);
and U11409 (N_11409,N_10648,N_10547);
nor U11410 (N_11410,N_10617,N_10832);
nor U11411 (N_11411,N_10887,N_10824);
nor U11412 (N_11412,N_10524,N_10742);
and U11413 (N_11413,N_10833,N_10991);
and U11414 (N_11414,N_10870,N_10654);
nor U11415 (N_11415,N_10870,N_10687);
nor U11416 (N_11416,N_10799,N_10608);
nor U11417 (N_11417,N_10737,N_10713);
nor U11418 (N_11418,N_10929,N_10549);
nand U11419 (N_11419,N_10652,N_10969);
or U11420 (N_11420,N_10730,N_10913);
or U11421 (N_11421,N_10966,N_10900);
nand U11422 (N_11422,N_10865,N_10807);
xnor U11423 (N_11423,N_10983,N_10744);
xor U11424 (N_11424,N_10683,N_10698);
and U11425 (N_11425,N_10592,N_10775);
nand U11426 (N_11426,N_10597,N_10958);
xor U11427 (N_11427,N_10737,N_10586);
and U11428 (N_11428,N_10648,N_10812);
nand U11429 (N_11429,N_10813,N_10685);
nand U11430 (N_11430,N_10638,N_10822);
nor U11431 (N_11431,N_10653,N_10559);
or U11432 (N_11432,N_10588,N_10933);
xnor U11433 (N_11433,N_10922,N_10757);
or U11434 (N_11434,N_10714,N_10844);
or U11435 (N_11435,N_10619,N_10575);
and U11436 (N_11436,N_10912,N_10776);
xor U11437 (N_11437,N_10810,N_10924);
or U11438 (N_11438,N_10740,N_10522);
xnor U11439 (N_11439,N_10507,N_10599);
nor U11440 (N_11440,N_10662,N_10588);
nand U11441 (N_11441,N_10626,N_10658);
or U11442 (N_11442,N_10585,N_10997);
nor U11443 (N_11443,N_10731,N_10637);
or U11444 (N_11444,N_10858,N_10508);
nand U11445 (N_11445,N_10827,N_10580);
nand U11446 (N_11446,N_10747,N_10918);
xor U11447 (N_11447,N_10504,N_10587);
xor U11448 (N_11448,N_10593,N_10934);
nor U11449 (N_11449,N_10889,N_10527);
xor U11450 (N_11450,N_10791,N_10524);
nand U11451 (N_11451,N_10839,N_10722);
xor U11452 (N_11452,N_10699,N_10871);
xor U11453 (N_11453,N_10647,N_10736);
nand U11454 (N_11454,N_10689,N_10647);
or U11455 (N_11455,N_10691,N_10987);
or U11456 (N_11456,N_10538,N_10994);
nor U11457 (N_11457,N_10813,N_10912);
xor U11458 (N_11458,N_10804,N_10676);
nand U11459 (N_11459,N_10737,N_10740);
and U11460 (N_11460,N_10529,N_10788);
nand U11461 (N_11461,N_10952,N_10565);
or U11462 (N_11462,N_10815,N_10501);
or U11463 (N_11463,N_10562,N_10679);
nand U11464 (N_11464,N_10904,N_10927);
and U11465 (N_11465,N_10996,N_10508);
nand U11466 (N_11466,N_10775,N_10869);
nand U11467 (N_11467,N_10563,N_10799);
nand U11468 (N_11468,N_10547,N_10637);
nor U11469 (N_11469,N_10653,N_10970);
and U11470 (N_11470,N_10505,N_10752);
and U11471 (N_11471,N_10874,N_10989);
and U11472 (N_11472,N_10963,N_10808);
nor U11473 (N_11473,N_10521,N_10697);
or U11474 (N_11474,N_10642,N_10701);
xnor U11475 (N_11475,N_10977,N_10904);
or U11476 (N_11476,N_10686,N_10721);
xnor U11477 (N_11477,N_10766,N_10613);
and U11478 (N_11478,N_10906,N_10526);
nand U11479 (N_11479,N_10656,N_10623);
or U11480 (N_11480,N_10546,N_10796);
or U11481 (N_11481,N_10726,N_10705);
nand U11482 (N_11482,N_10868,N_10605);
nand U11483 (N_11483,N_10851,N_10855);
nor U11484 (N_11484,N_10653,N_10879);
nand U11485 (N_11485,N_10640,N_10651);
nor U11486 (N_11486,N_10892,N_10966);
nand U11487 (N_11487,N_10607,N_10814);
and U11488 (N_11488,N_10993,N_10561);
or U11489 (N_11489,N_10553,N_10958);
or U11490 (N_11490,N_10692,N_10596);
nand U11491 (N_11491,N_10539,N_10541);
or U11492 (N_11492,N_10554,N_10733);
and U11493 (N_11493,N_10515,N_10604);
and U11494 (N_11494,N_10507,N_10582);
nand U11495 (N_11495,N_10966,N_10979);
xor U11496 (N_11496,N_10811,N_10910);
and U11497 (N_11497,N_10750,N_10716);
nor U11498 (N_11498,N_10715,N_10582);
nor U11499 (N_11499,N_10728,N_10550);
and U11500 (N_11500,N_11363,N_11171);
nand U11501 (N_11501,N_11205,N_11396);
or U11502 (N_11502,N_11028,N_11178);
xor U11503 (N_11503,N_11223,N_11295);
nand U11504 (N_11504,N_11119,N_11072);
nor U11505 (N_11505,N_11381,N_11388);
and U11506 (N_11506,N_11261,N_11096);
nor U11507 (N_11507,N_11282,N_11300);
or U11508 (N_11508,N_11471,N_11418);
or U11509 (N_11509,N_11422,N_11234);
and U11510 (N_11510,N_11122,N_11177);
xor U11511 (N_11511,N_11137,N_11366);
xnor U11512 (N_11512,N_11196,N_11309);
nand U11513 (N_11513,N_11324,N_11395);
nand U11514 (N_11514,N_11085,N_11157);
nor U11515 (N_11515,N_11461,N_11315);
nor U11516 (N_11516,N_11424,N_11148);
nand U11517 (N_11517,N_11293,N_11145);
xor U11518 (N_11518,N_11308,N_11139);
and U11519 (N_11519,N_11417,N_11018);
or U11520 (N_11520,N_11345,N_11033);
nor U11521 (N_11521,N_11252,N_11380);
and U11522 (N_11522,N_11231,N_11022);
or U11523 (N_11523,N_11064,N_11184);
nor U11524 (N_11524,N_11495,N_11128);
or U11525 (N_11525,N_11399,N_11191);
and U11526 (N_11526,N_11368,N_11106);
and U11527 (N_11527,N_11089,N_11450);
xnor U11528 (N_11528,N_11311,N_11305);
or U11529 (N_11529,N_11485,N_11135);
and U11530 (N_11530,N_11406,N_11431);
and U11531 (N_11531,N_11480,N_11220);
and U11532 (N_11532,N_11218,N_11056);
and U11533 (N_11533,N_11365,N_11006);
nand U11534 (N_11534,N_11465,N_11049);
xor U11535 (N_11535,N_11172,N_11004);
or U11536 (N_11536,N_11116,N_11207);
or U11537 (N_11537,N_11012,N_11247);
and U11538 (N_11538,N_11038,N_11105);
nand U11539 (N_11539,N_11151,N_11017);
or U11540 (N_11540,N_11425,N_11025);
nand U11541 (N_11541,N_11158,N_11244);
xor U11542 (N_11542,N_11419,N_11156);
nand U11543 (N_11543,N_11270,N_11228);
xnor U11544 (N_11544,N_11246,N_11109);
and U11545 (N_11545,N_11074,N_11059);
or U11546 (N_11546,N_11445,N_11164);
xor U11547 (N_11547,N_11052,N_11199);
and U11548 (N_11548,N_11313,N_11120);
nor U11549 (N_11549,N_11267,N_11041);
xnor U11550 (N_11550,N_11389,N_11131);
xnor U11551 (N_11551,N_11376,N_11273);
nand U11552 (N_11552,N_11217,N_11159);
or U11553 (N_11553,N_11352,N_11414);
xor U11554 (N_11554,N_11342,N_11170);
xnor U11555 (N_11555,N_11484,N_11115);
nor U11556 (N_11556,N_11254,N_11104);
nor U11557 (N_11557,N_11467,N_11113);
and U11558 (N_11558,N_11434,N_11200);
or U11559 (N_11559,N_11063,N_11264);
nand U11560 (N_11560,N_11277,N_11492);
and U11561 (N_11561,N_11369,N_11031);
and U11562 (N_11562,N_11221,N_11143);
nor U11563 (N_11563,N_11427,N_11413);
nand U11564 (N_11564,N_11092,N_11097);
nand U11565 (N_11565,N_11192,N_11426);
and U11566 (N_11566,N_11167,N_11242);
nand U11567 (N_11567,N_11343,N_11250);
and U11568 (N_11568,N_11408,N_11141);
and U11569 (N_11569,N_11144,N_11232);
or U11570 (N_11570,N_11090,N_11000);
nor U11571 (N_11571,N_11405,N_11146);
and U11572 (N_11572,N_11103,N_11360);
nand U11573 (N_11573,N_11204,N_11451);
and U11574 (N_11574,N_11454,N_11398);
or U11575 (N_11575,N_11463,N_11392);
nor U11576 (N_11576,N_11081,N_11362);
nor U11577 (N_11577,N_11374,N_11401);
xor U11578 (N_11578,N_11462,N_11168);
or U11579 (N_11579,N_11475,N_11420);
and U11580 (N_11580,N_11314,N_11444);
or U11581 (N_11581,N_11384,N_11078);
nand U11582 (N_11582,N_11227,N_11416);
xor U11583 (N_11583,N_11403,N_11130);
nor U11584 (N_11584,N_11225,N_11108);
nand U11585 (N_11585,N_11377,N_11447);
nand U11586 (N_11586,N_11235,N_11349);
or U11587 (N_11587,N_11299,N_11236);
nor U11588 (N_11588,N_11323,N_11442);
nor U11589 (N_11589,N_11358,N_11367);
nor U11590 (N_11590,N_11364,N_11446);
or U11591 (N_11591,N_11339,N_11430);
and U11592 (N_11592,N_11248,N_11002);
xor U11593 (N_11593,N_11259,N_11029);
nand U11594 (N_11594,N_11329,N_11036);
and U11595 (N_11595,N_11240,N_11320);
xor U11596 (N_11596,N_11265,N_11479);
nand U11597 (N_11597,N_11188,N_11400);
nor U11598 (N_11598,N_11147,N_11271);
or U11599 (N_11599,N_11082,N_11073);
nand U11600 (N_11600,N_11040,N_11001);
nand U11601 (N_11601,N_11125,N_11212);
xor U11602 (N_11602,N_11013,N_11140);
or U11603 (N_11603,N_11245,N_11088);
nor U11604 (N_11604,N_11015,N_11032);
and U11605 (N_11605,N_11307,N_11045);
and U11606 (N_11606,N_11276,N_11288);
and U11607 (N_11607,N_11468,N_11303);
nor U11608 (N_11608,N_11067,N_11497);
or U11609 (N_11609,N_11460,N_11043);
and U11610 (N_11610,N_11016,N_11490);
and U11611 (N_11611,N_11214,N_11292);
and U11612 (N_11612,N_11152,N_11154);
nor U11613 (N_11613,N_11283,N_11357);
xor U11614 (N_11614,N_11111,N_11331);
and U11615 (N_11615,N_11176,N_11397);
nand U11616 (N_11616,N_11173,N_11393);
nand U11617 (N_11617,N_11211,N_11213);
nor U11618 (N_11618,N_11257,N_11410);
xnor U11619 (N_11619,N_11457,N_11449);
xor U11620 (N_11620,N_11057,N_11421);
or U11621 (N_11621,N_11226,N_11356);
and U11622 (N_11622,N_11075,N_11117);
and U11623 (N_11623,N_11336,N_11243);
xor U11624 (N_11624,N_11224,N_11179);
nand U11625 (N_11625,N_11298,N_11284);
and U11626 (N_11626,N_11455,N_11316);
xnor U11627 (N_11627,N_11302,N_11438);
xnor U11628 (N_11628,N_11326,N_11373);
or U11629 (N_11629,N_11080,N_11429);
nor U11630 (N_11630,N_11290,N_11165);
nor U11631 (N_11631,N_11216,N_11286);
or U11632 (N_11632,N_11253,N_11306);
nor U11633 (N_11633,N_11155,N_11023);
or U11634 (N_11634,N_11037,N_11047);
nor U11635 (N_11635,N_11448,N_11150);
nand U11636 (N_11636,N_11436,N_11142);
nand U11637 (N_11637,N_11340,N_11107);
nand U11638 (N_11638,N_11301,N_11136);
nand U11639 (N_11639,N_11132,N_11206);
nor U11640 (N_11640,N_11354,N_11258);
nand U11641 (N_11641,N_11070,N_11432);
and U11642 (N_11642,N_11034,N_11193);
nand U11643 (N_11643,N_11325,N_11428);
xnor U11644 (N_11644,N_11269,N_11496);
nor U11645 (N_11645,N_11415,N_11337);
and U11646 (N_11646,N_11319,N_11189);
nand U11647 (N_11647,N_11441,N_11433);
nand U11648 (N_11648,N_11359,N_11394);
and U11649 (N_11649,N_11333,N_11387);
or U11650 (N_11650,N_11201,N_11190);
or U11651 (N_11651,N_11322,N_11472);
and U11652 (N_11652,N_11129,N_11327);
nand U11653 (N_11653,N_11478,N_11383);
and U11654 (N_11654,N_11249,N_11330);
or U11655 (N_11655,N_11317,N_11348);
and U11656 (N_11656,N_11035,N_11486);
xor U11657 (N_11657,N_11048,N_11102);
nor U11658 (N_11658,N_11278,N_11187);
nor U11659 (N_11659,N_11355,N_11008);
xnor U11660 (N_11660,N_11233,N_11153);
or U11661 (N_11661,N_11161,N_11412);
nor U11662 (N_11662,N_11186,N_11251);
or U11663 (N_11663,N_11378,N_11222);
nand U11664 (N_11664,N_11274,N_11112);
nand U11665 (N_11665,N_11077,N_11493);
nor U11666 (N_11666,N_11208,N_11499);
xor U11667 (N_11667,N_11439,N_11042);
nand U11668 (N_11668,N_11114,N_11239);
or U11669 (N_11669,N_11456,N_11459);
nand U11670 (N_11670,N_11066,N_11050);
nand U11671 (N_11671,N_11098,N_11382);
xor U11672 (N_11672,N_11481,N_11407);
xor U11673 (N_11673,N_11255,N_11310);
or U11674 (N_11674,N_11346,N_11044);
xor U11675 (N_11675,N_11005,N_11100);
nor U11676 (N_11676,N_11219,N_11391);
and U11677 (N_11677,N_11489,N_11021);
or U11678 (N_11678,N_11361,N_11379);
nand U11679 (N_11679,N_11210,N_11385);
xor U11680 (N_11680,N_11014,N_11160);
or U11681 (N_11681,N_11279,N_11068);
nor U11682 (N_11682,N_11477,N_11263);
or U11683 (N_11683,N_11071,N_11198);
nor U11684 (N_11684,N_11007,N_11084);
nand U11685 (N_11685,N_11076,N_11474);
nand U11686 (N_11686,N_11209,N_11423);
nor U11687 (N_11687,N_11024,N_11297);
xnor U11688 (N_11688,N_11093,N_11027);
nand U11689 (N_11689,N_11470,N_11351);
nand U11690 (N_11690,N_11046,N_11335);
or U11691 (N_11691,N_11183,N_11280);
nand U11692 (N_11692,N_11149,N_11488);
nor U11693 (N_11693,N_11118,N_11291);
xor U11694 (N_11694,N_11404,N_11241);
xor U11695 (N_11695,N_11175,N_11272);
xnor U11696 (N_11696,N_11466,N_11289);
nand U11697 (N_11697,N_11197,N_11055);
and U11698 (N_11698,N_11498,N_11126);
xor U11699 (N_11699,N_11230,N_11294);
nand U11700 (N_11700,N_11091,N_11370);
xnor U11701 (N_11701,N_11386,N_11039);
nor U11702 (N_11702,N_11347,N_11138);
nor U11703 (N_11703,N_11304,N_11341);
or U11704 (N_11704,N_11409,N_11473);
and U11705 (N_11705,N_11372,N_11215);
nor U11706 (N_11706,N_11202,N_11133);
nor U11707 (N_11707,N_11411,N_11287);
and U11708 (N_11708,N_11203,N_11443);
xnor U11709 (N_11709,N_11487,N_11229);
and U11710 (N_11710,N_11328,N_11285);
nand U11711 (N_11711,N_11318,N_11051);
and U11712 (N_11712,N_11321,N_11010);
nand U11713 (N_11713,N_11087,N_11182);
and U11714 (N_11714,N_11069,N_11237);
nor U11715 (N_11715,N_11127,N_11312);
or U11716 (N_11716,N_11053,N_11194);
or U11717 (N_11717,N_11371,N_11083);
and U11718 (N_11718,N_11494,N_11121);
xor U11719 (N_11719,N_11344,N_11060);
xnor U11720 (N_11720,N_11061,N_11062);
and U11721 (N_11721,N_11110,N_11101);
and U11722 (N_11722,N_11482,N_11453);
or U11723 (N_11723,N_11054,N_11375);
and U11724 (N_11724,N_11185,N_11390);
nand U11725 (N_11725,N_11019,N_11094);
or U11726 (N_11726,N_11268,N_11020);
nor U11727 (N_11727,N_11123,N_11058);
nand U11728 (N_11728,N_11266,N_11332);
nand U11729 (N_11729,N_11260,N_11011);
or U11730 (N_11730,N_11079,N_11464);
or U11731 (N_11731,N_11065,N_11458);
or U11732 (N_11732,N_11195,N_11469);
xor U11733 (N_11733,N_11174,N_11262);
or U11734 (N_11734,N_11350,N_11437);
and U11735 (N_11735,N_11003,N_11491);
and U11736 (N_11736,N_11181,N_11281);
or U11737 (N_11737,N_11275,N_11440);
nand U11738 (N_11738,N_11353,N_11086);
xnor U11739 (N_11739,N_11169,N_11338);
xnor U11740 (N_11740,N_11026,N_11009);
and U11741 (N_11741,N_11238,N_11402);
nor U11742 (N_11742,N_11296,N_11452);
nand U11743 (N_11743,N_11099,N_11256);
and U11744 (N_11744,N_11124,N_11030);
and U11745 (N_11745,N_11095,N_11163);
and U11746 (N_11746,N_11180,N_11166);
xnor U11747 (N_11747,N_11334,N_11134);
and U11748 (N_11748,N_11162,N_11435);
xnor U11749 (N_11749,N_11483,N_11476);
or U11750 (N_11750,N_11177,N_11499);
xnor U11751 (N_11751,N_11444,N_11084);
and U11752 (N_11752,N_11135,N_11363);
nor U11753 (N_11753,N_11146,N_11443);
xor U11754 (N_11754,N_11017,N_11131);
and U11755 (N_11755,N_11001,N_11008);
nand U11756 (N_11756,N_11304,N_11396);
and U11757 (N_11757,N_11081,N_11203);
and U11758 (N_11758,N_11414,N_11475);
nor U11759 (N_11759,N_11390,N_11303);
nand U11760 (N_11760,N_11366,N_11155);
nand U11761 (N_11761,N_11042,N_11098);
and U11762 (N_11762,N_11183,N_11190);
nand U11763 (N_11763,N_11303,N_11146);
nand U11764 (N_11764,N_11446,N_11296);
nand U11765 (N_11765,N_11214,N_11359);
nand U11766 (N_11766,N_11487,N_11242);
nand U11767 (N_11767,N_11406,N_11243);
nand U11768 (N_11768,N_11440,N_11008);
nor U11769 (N_11769,N_11241,N_11188);
nand U11770 (N_11770,N_11043,N_11041);
and U11771 (N_11771,N_11099,N_11426);
and U11772 (N_11772,N_11042,N_11212);
or U11773 (N_11773,N_11396,N_11203);
or U11774 (N_11774,N_11299,N_11371);
or U11775 (N_11775,N_11100,N_11086);
xnor U11776 (N_11776,N_11355,N_11497);
nor U11777 (N_11777,N_11492,N_11337);
nand U11778 (N_11778,N_11320,N_11073);
and U11779 (N_11779,N_11479,N_11455);
xnor U11780 (N_11780,N_11065,N_11039);
nand U11781 (N_11781,N_11100,N_11414);
or U11782 (N_11782,N_11091,N_11006);
xor U11783 (N_11783,N_11136,N_11125);
xnor U11784 (N_11784,N_11053,N_11240);
xor U11785 (N_11785,N_11046,N_11433);
xor U11786 (N_11786,N_11065,N_11429);
and U11787 (N_11787,N_11339,N_11379);
nor U11788 (N_11788,N_11251,N_11448);
nor U11789 (N_11789,N_11452,N_11392);
nand U11790 (N_11790,N_11476,N_11040);
nand U11791 (N_11791,N_11383,N_11101);
xor U11792 (N_11792,N_11348,N_11340);
nand U11793 (N_11793,N_11335,N_11339);
nand U11794 (N_11794,N_11316,N_11422);
xor U11795 (N_11795,N_11413,N_11342);
and U11796 (N_11796,N_11245,N_11288);
and U11797 (N_11797,N_11095,N_11431);
and U11798 (N_11798,N_11454,N_11053);
xnor U11799 (N_11799,N_11088,N_11365);
nand U11800 (N_11800,N_11408,N_11152);
nand U11801 (N_11801,N_11266,N_11191);
and U11802 (N_11802,N_11144,N_11117);
nand U11803 (N_11803,N_11418,N_11239);
or U11804 (N_11804,N_11421,N_11290);
and U11805 (N_11805,N_11151,N_11111);
and U11806 (N_11806,N_11001,N_11028);
and U11807 (N_11807,N_11352,N_11283);
xnor U11808 (N_11808,N_11486,N_11259);
nor U11809 (N_11809,N_11207,N_11255);
nand U11810 (N_11810,N_11401,N_11068);
xor U11811 (N_11811,N_11376,N_11415);
nor U11812 (N_11812,N_11339,N_11094);
xnor U11813 (N_11813,N_11150,N_11019);
and U11814 (N_11814,N_11212,N_11426);
nand U11815 (N_11815,N_11364,N_11325);
or U11816 (N_11816,N_11379,N_11061);
xor U11817 (N_11817,N_11056,N_11136);
nand U11818 (N_11818,N_11076,N_11346);
or U11819 (N_11819,N_11025,N_11347);
nor U11820 (N_11820,N_11405,N_11379);
xor U11821 (N_11821,N_11047,N_11049);
nor U11822 (N_11822,N_11132,N_11337);
or U11823 (N_11823,N_11170,N_11196);
nand U11824 (N_11824,N_11358,N_11322);
xnor U11825 (N_11825,N_11319,N_11473);
and U11826 (N_11826,N_11404,N_11420);
or U11827 (N_11827,N_11028,N_11258);
nand U11828 (N_11828,N_11384,N_11214);
and U11829 (N_11829,N_11130,N_11306);
and U11830 (N_11830,N_11215,N_11148);
xor U11831 (N_11831,N_11185,N_11208);
nand U11832 (N_11832,N_11195,N_11040);
and U11833 (N_11833,N_11499,N_11286);
or U11834 (N_11834,N_11124,N_11240);
and U11835 (N_11835,N_11494,N_11488);
or U11836 (N_11836,N_11008,N_11187);
or U11837 (N_11837,N_11121,N_11288);
and U11838 (N_11838,N_11038,N_11324);
nor U11839 (N_11839,N_11307,N_11243);
or U11840 (N_11840,N_11075,N_11104);
or U11841 (N_11841,N_11240,N_11147);
xor U11842 (N_11842,N_11137,N_11002);
nor U11843 (N_11843,N_11286,N_11489);
and U11844 (N_11844,N_11424,N_11468);
nand U11845 (N_11845,N_11065,N_11194);
or U11846 (N_11846,N_11495,N_11459);
nor U11847 (N_11847,N_11007,N_11102);
nand U11848 (N_11848,N_11335,N_11322);
or U11849 (N_11849,N_11086,N_11451);
xor U11850 (N_11850,N_11483,N_11098);
nand U11851 (N_11851,N_11224,N_11482);
and U11852 (N_11852,N_11308,N_11258);
and U11853 (N_11853,N_11120,N_11208);
or U11854 (N_11854,N_11393,N_11386);
nor U11855 (N_11855,N_11127,N_11247);
and U11856 (N_11856,N_11087,N_11229);
nand U11857 (N_11857,N_11383,N_11289);
xnor U11858 (N_11858,N_11029,N_11206);
xor U11859 (N_11859,N_11295,N_11061);
nand U11860 (N_11860,N_11486,N_11013);
nand U11861 (N_11861,N_11033,N_11041);
and U11862 (N_11862,N_11246,N_11080);
or U11863 (N_11863,N_11215,N_11485);
nor U11864 (N_11864,N_11009,N_11394);
nand U11865 (N_11865,N_11359,N_11468);
and U11866 (N_11866,N_11187,N_11255);
nand U11867 (N_11867,N_11008,N_11234);
or U11868 (N_11868,N_11368,N_11419);
and U11869 (N_11869,N_11047,N_11116);
and U11870 (N_11870,N_11352,N_11134);
or U11871 (N_11871,N_11029,N_11472);
xnor U11872 (N_11872,N_11238,N_11454);
and U11873 (N_11873,N_11315,N_11467);
nand U11874 (N_11874,N_11173,N_11489);
xor U11875 (N_11875,N_11486,N_11322);
or U11876 (N_11876,N_11080,N_11134);
nor U11877 (N_11877,N_11055,N_11050);
and U11878 (N_11878,N_11286,N_11111);
xor U11879 (N_11879,N_11107,N_11272);
nor U11880 (N_11880,N_11235,N_11337);
and U11881 (N_11881,N_11468,N_11094);
xnor U11882 (N_11882,N_11444,N_11289);
and U11883 (N_11883,N_11387,N_11069);
and U11884 (N_11884,N_11281,N_11068);
xnor U11885 (N_11885,N_11150,N_11112);
nor U11886 (N_11886,N_11197,N_11132);
xor U11887 (N_11887,N_11448,N_11345);
and U11888 (N_11888,N_11082,N_11394);
or U11889 (N_11889,N_11238,N_11160);
or U11890 (N_11890,N_11014,N_11161);
xnor U11891 (N_11891,N_11009,N_11074);
or U11892 (N_11892,N_11321,N_11292);
and U11893 (N_11893,N_11295,N_11200);
nor U11894 (N_11894,N_11040,N_11178);
and U11895 (N_11895,N_11135,N_11145);
or U11896 (N_11896,N_11353,N_11317);
nor U11897 (N_11897,N_11117,N_11158);
xnor U11898 (N_11898,N_11295,N_11403);
or U11899 (N_11899,N_11158,N_11070);
nand U11900 (N_11900,N_11496,N_11182);
xor U11901 (N_11901,N_11353,N_11242);
or U11902 (N_11902,N_11410,N_11194);
and U11903 (N_11903,N_11447,N_11002);
nand U11904 (N_11904,N_11380,N_11459);
and U11905 (N_11905,N_11040,N_11274);
nor U11906 (N_11906,N_11280,N_11259);
and U11907 (N_11907,N_11341,N_11388);
xnor U11908 (N_11908,N_11457,N_11426);
nand U11909 (N_11909,N_11097,N_11440);
and U11910 (N_11910,N_11334,N_11348);
or U11911 (N_11911,N_11280,N_11385);
xor U11912 (N_11912,N_11463,N_11205);
xnor U11913 (N_11913,N_11048,N_11064);
nor U11914 (N_11914,N_11357,N_11107);
xnor U11915 (N_11915,N_11297,N_11250);
nand U11916 (N_11916,N_11170,N_11291);
and U11917 (N_11917,N_11002,N_11168);
and U11918 (N_11918,N_11280,N_11129);
or U11919 (N_11919,N_11297,N_11131);
nand U11920 (N_11920,N_11174,N_11454);
nand U11921 (N_11921,N_11372,N_11159);
nand U11922 (N_11922,N_11446,N_11438);
and U11923 (N_11923,N_11404,N_11308);
or U11924 (N_11924,N_11205,N_11459);
or U11925 (N_11925,N_11160,N_11226);
or U11926 (N_11926,N_11424,N_11278);
nor U11927 (N_11927,N_11114,N_11443);
nor U11928 (N_11928,N_11104,N_11261);
xor U11929 (N_11929,N_11321,N_11324);
nor U11930 (N_11930,N_11169,N_11029);
nand U11931 (N_11931,N_11003,N_11467);
and U11932 (N_11932,N_11040,N_11170);
xor U11933 (N_11933,N_11257,N_11277);
nor U11934 (N_11934,N_11299,N_11105);
nor U11935 (N_11935,N_11324,N_11423);
and U11936 (N_11936,N_11350,N_11308);
xnor U11937 (N_11937,N_11033,N_11321);
nand U11938 (N_11938,N_11435,N_11140);
nand U11939 (N_11939,N_11376,N_11304);
nand U11940 (N_11940,N_11023,N_11434);
nand U11941 (N_11941,N_11037,N_11074);
xnor U11942 (N_11942,N_11164,N_11336);
nor U11943 (N_11943,N_11423,N_11020);
xor U11944 (N_11944,N_11240,N_11036);
and U11945 (N_11945,N_11460,N_11171);
nand U11946 (N_11946,N_11174,N_11275);
xor U11947 (N_11947,N_11188,N_11442);
xor U11948 (N_11948,N_11245,N_11273);
and U11949 (N_11949,N_11326,N_11011);
or U11950 (N_11950,N_11209,N_11400);
nor U11951 (N_11951,N_11031,N_11164);
nand U11952 (N_11952,N_11124,N_11051);
and U11953 (N_11953,N_11160,N_11211);
xnor U11954 (N_11954,N_11414,N_11306);
nand U11955 (N_11955,N_11181,N_11174);
xnor U11956 (N_11956,N_11257,N_11328);
nand U11957 (N_11957,N_11471,N_11334);
nand U11958 (N_11958,N_11039,N_11024);
or U11959 (N_11959,N_11424,N_11044);
nand U11960 (N_11960,N_11228,N_11320);
or U11961 (N_11961,N_11033,N_11346);
nor U11962 (N_11962,N_11206,N_11332);
and U11963 (N_11963,N_11464,N_11275);
and U11964 (N_11964,N_11087,N_11444);
nand U11965 (N_11965,N_11301,N_11235);
nand U11966 (N_11966,N_11324,N_11017);
or U11967 (N_11967,N_11291,N_11375);
xnor U11968 (N_11968,N_11405,N_11394);
nand U11969 (N_11969,N_11069,N_11207);
nor U11970 (N_11970,N_11252,N_11190);
xor U11971 (N_11971,N_11080,N_11142);
nor U11972 (N_11972,N_11424,N_11341);
xnor U11973 (N_11973,N_11283,N_11050);
xnor U11974 (N_11974,N_11207,N_11065);
and U11975 (N_11975,N_11471,N_11369);
xnor U11976 (N_11976,N_11061,N_11113);
or U11977 (N_11977,N_11467,N_11355);
nor U11978 (N_11978,N_11095,N_11221);
xnor U11979 (N_11979,N_11302,N_11232);
xor U11980 (N_11980,N_11001,N_11379);
or U11981 (N_11981,N_11226,N_11244);
xor U11982 (N_11982,N_11012,N_11169);
nor U11983 (N_11983,N_11071,N_11251);
and U11984 (N_11984,N_11138,N_11276);
or U11985 (N_11985,N_11194,N_11076);
nand U11986 (N_11986,N_11063,N_11164);
and U11987 (N_11987,N_11348,N_11292);
xor U11988 (N_11988,N_11417,N_11481);
nand U11989 (N_11989,N_11236,N_11326);
and U11990 (N_11990,N_11229,N_11163);
or U11991 (N_11991,N_11359,N_11356);
xor U11992 (N_11992,N_11232,N_11086);
xnor U11993 (N_11993,N_11282,N_11433);
nor U11994 (N_11994,N_11487,N_11199);
or U11995 (N_11995,N_11332,N_11383);
nand U11996 (N_11996,N_11011,N_11350);
and U11997 (N_11997,N_11100,N_11167);
and U11998 (N_11998,N_11036,N_11100);
nor U11999 (N_11999,N_11201,N_11477);
or U12000 (N_12000,N_11571,N_11969);
xor U12001 (N_12001,N_11646,N_11778);
nand U12002 (N_12002,N_11694,N_11934);
xor U12003 (N_12003,N_11864,N_11554);
or U12004 (N_12004,N_11516,N_11693);
and U12005 (N_12005,N_11574,N_11504);
or U12006 (N_12006,N_11797,N_11783);
or U12007 (N_12007,N_11922,N_11687);
and U12008 (N_12008,N_11983,N_11753);
nor U12009 (N_12009,N_11745,N_11545);
or U12010 (N_12010,N_11506,N_11820);
nor U12011 (N_12011,N_11813,N_11639);
nand U12012 (N_12012,N_11682,N_11530);
nand U12013 (N_12013,N_11696,N_11844);
xor U12014 (N_12014,N_11752,N_11588);
nand U12015 (N_12015,N_11823,N_11601);
or U12016 (N_12016,N_11621,N_11970);
xnor U12017 (N_12017,N_11622,N_11718);
or U12018 (N_12018,N_11917,N_11677);
nand U12019 (N_12019,N_11547,N_11563);
nand U12020 (N_12020,N_11559,N_11916);
nor U12021 (N_12021,N_11848,N_11873);
nand U12022 (N_12022,N_11929,N_11827);
nor U12023 (N_12023,N_11643,N_11534);
and U12024 (N_12024,N_11635,N_11722);
xnor U12025 (N_12025,N_11605,N_11985);
or U12026 (N_12026,N_11749,N_11736);
xor U12027 (N_12027,N_11793,N_11960);
or U12028 (N_12028,N_11772,N_11738);
nand U12029 (N_12029,N_11587,N_11914);
or U12030 (N_12030,N_11689,N_11940);
xor U12031 (N_12031,N_11552,N_11840);
or U12032 (N_12032,N_11791,N_11822);
and U12033 (N_12033,N_11730,N_11876);
xnor U12034 (N_12034,N_11544,N_11968);
nor U12035 (N_12035,N_11867,N_11603);
and U12036 (N_12036,N_11926,N_11888);
nand U12037 (N_12037,N_11734,N_11654);
xnor U12038 (N_12038,N_11548,N_11656);
xor U12039 (N_12039,N_11862,N_11649);
and U12040 (N_12040,N_11727,N_11598);
xnor U12041 (N_12041,N_11992,N_11626);
nand U12042 (N_12042,N_11664,N_11683);
nor U12043 (N_12043,N_11991,N_11859);
nand U12044 (N_12044,N_11742,N_11703);
and U12045 (N_12045,N_11769,N_11925);
and U12046 (N_12046,N_11755,N_11996);
nor U12047 (N_12047,N_11704,N_11511);
xor U12048 (N_12048,N_11861,N_11606);
and U12049 (N_12049,N_11828,N_11717);
xor U12050 (N_12050,N_11507,N_11855);
nor U12051 (N_12051,N_11789,N_11614);
xnor U12052 (N_12052,N_11853,N_11540);
or U12053 (N_12053,N_11774,N_11972);
or U12054 (N_12054,N_11818,N_11674);
nand U12055 (N_12055,N_11645,N_11673);
xnor U12056 (N_12056,N_11777,N_11883);
nor U12057 (N_12057,N_11653,N_11805);
or U12058 (N_12058,N_11640,N_11806);
xnor U12059 (N_12059,N_11838,N_11663);
nand U12060 (N_12060,N_11543,N_11661);
xor U12061 (N_12061,N_11939,N_11585);
xnor U12062 (N_12062,N_11651,N_11556);
and U12063 (N_12063,N_11503,N_11933);
nand U12064 (N_12064,N_11909,N_11878);
nand U12065 (N_12065,N_11636,N_11565);
and U12066 (N_12066,N_11505,N_11986);
and U12067 (N_12067,N_11566,N_11685);
or U12068 (N_12068,N_11510,N_11905);
xnor U12069 (N_12069,N_11668,N_11652);
xor U12070 (N_12070,N_11549,N_11580);
nand U12071 (N_12071,N_11583,N_11773);
xnor U12072 (N_12072,N_11965,N_11837);
and U12073 (N_12073,N_11557,N_11567);
nand U12074 (N_12074,N_11650,N_11799);
xnor U12075 (N_12075,N_11959,N_11949);
nand U12076 (N_12076,N_11898,N_11679);
xor U12077 (N_12077,N_11915,N_11942);
nand U12078 (N_12078,N_11520,N_11512);
nor U12079 (N_12079,N_11521,N_11884);
or U12080 (N_12080,N_11719,N_11961);
nand U12081 (N_12081,N_11962,N_11629);
nand U12082 (N_12082,N_11633,N_11887);
nand U12083 (N_12083,N_11569,N_11821);
or U12084 (N_12084,N_11760,N_11950);
or U12085 (N_12085,N_11714,N_11576);
nand U12086 (N_12086,N_11988,N_11570);
nor U12087 (N_12087,N_11817,N_11667);
nand U12088 (N_12088,N_11509,N_11819);
or U12089 (N_12089,N_11660,N_11766);
or U12090 (N_12090,N_11886,N_11780);
nor U12091 (N_12091,N_11947,N_11715);
or U12092 (N_12092,N_11784,N_11658);
xnor U12093 (N_12093,N_11675,N_11941);
nor U12094 (N_12094,N_11584,N_11684);
nor U12095 (N_12095,N_11918,N_11857);
xor U12096 (N_12096,N_11904,N_11731);
xor U12097 (N_12097,N_11871,N_11608);
nand U12098 (N_12098,N_11907,N_11836);
and U12099 (N_12099,N_11938,N_11692);
or U12100 (N_12100,N_11798,N_11865);
nand U12101 (N_12101,N_11558,N_11691);
xnor U12102 (N_12102,N_11958,N_11826);
or U12103 (N_12103,N_11973,N_11852);
nand U12104 (N_12104,N_11741,N_11787);
nor U12105 (N_12105,N_11816,N_11721);
nand U12106 (N_12106,N_11593,N_11690);
and U12107 (N_12107,N_11885,N_11600);
nand U12108 (N_12108,N_11644,N_11733);
xor U12109 (N_12109,N_11845,N_11634);
nand U12110 (N_12110,N_11908,N_11720);
nor U12111 (N_12111,N_11551,N_11627);
nor U12112 (N_12112,N_11604,N_11708);
or U12113 (N_12113,N_11850,N_11523);
nor U12114 (N_12114,N_11573,N_11586);
and U12115 (N_12115,N_11517,N_11589);
xnor U12116 (N_12116,N_11982,N_11804);
xor U12117 (N_12117,N_11882,N_11538);
nand U12118 (N_12118,N_11642,N_11762);
or U12119 (N_12119,N_11758,N_11901);
or U12120 (N_12120,N_11872,N_11712);
or U12121 (N_12121,N_11531,N_11782);
nor U12122 (N_12122,N_11607,N_11880);
xnor U12123 (N_12123,N_11539,N_11709);
xnor U12124 (N_12124,N_11529,N_11553);
and U12125 (N_12125,N_11666,N_11617);
or U12126 (N_12126,N_11632,N_11810);
or U12127 (N_12127,N_11648,N_11894);
xor U12128 (N_12128,N_11681,N_11781);
xnor U12129 (N_12129,N_11701,N_11832);
xor U12130 (N_12130,N_11670,N_11954);
xor U12131 (N_12131,N_11564,N_11971);
nand U12132 (N_12132,N_11863,N_11856);
or U12133 (N_12133,N_11906,N_11581);
and U12134 (N_12134,N_11868,N_11532);
or U12135 (N_12135,N_11750,N_11526);
nand U12136 (N_12136,N_11870,N_11809);
xnor U12137 (N_12137,N_11928,N_11989);
xnor U12138 (N_12138,N_11792,N_11881);
nand U12139 (N_12139,N_11524,N_11814);
or U12140 (N_12140,N_11542,N_11946);
nand U12141 (N_12141,N_11628,N_11980);
nor U12142 (N_12142,N_11609,N_11582);
xnor U12143 (N_12143,N_11611,N_11678);
xnor U12144 (N_12144,N_11525,N_11711);
and U12145 (N_12145,N_11994,N_11533);
or U12146 (N_12146,N_11619,N_11936);
and U12147 (N_12147,N_11546,N_11599);
nand U12148 (N_12148,N_11877,N_11514);
nor U12149 (N_12149,N_11515,N_11974);
nor U12150 (N_12150,N_11702,N_11808);
nor U12151 (N_12151,N_11975,N_11647);
nand U12152 (N_12152,N_11561,N_11981);
or U12153 (N_12153,N_11943,N_11843);
nor U12154 (N_12154,N_11706,N_11625);
xnor U12155 (N_12155,N_11802,N_11834);
nor U12156 (N_12156,N_11923,N_11790);
and U12157 (N_12157,N_11594,N_11978);
and U12158 (N_12158,N_11623,N_11775);
and U12159 (N_12159,N_11671,N_11785);
xor U12160 (N_12160,N_11676,N_11912);
and U12161 (N_12161,N_11964,N_11620);
and U12162 (N_12162,N_11765,N_11699);
xor U12163 (N_12163,N_11725,N_11737);
or U12164 (N_12164,N_11896,N_11579);
xnor U12165 (N_12165,N_11550,N_11747);
xnor U12166 (N_12166,N_11776,N_11815);
xnor U12167 (N_12167,N_11637,N_11860);
nand U12168 (N_12168,N_11842,N_11931);
nor U12169 (N_12169,N_11957,N_11500);
nor U12170 (N_12170,N_11732,N_11921);
xnor U12171 (N_12171,N_11841,N_11953);
nand U12172 (N_12172,N_11779,N_11590);
xnor U12173 (N_12173,N_11924,N_11761);
nand U12174 (N_12174,N_11578,N_11707);
nor U12175 (N_12175,N_11695,N_11669);
and U12176 (N_12176,N_11680,N_11688);
nor U12177 (N_12177,N_11613,N_11910);
or U12178 (N_12178,N_11955,N_11657);
nor U12179 (N_12179,N_11794,N_11739);
nor U12180 (N_12180,N_11522,N_11875);
or U12181 (N_12181,N_11890,N_11811);
and U12182 (N_12182,N_11560,N_11786);
and U12183 (N_12183,N_11829,N_11911);
xor U12184 (N_12184,N_11927,N_11698);
nor U12185 (N_12185,N_11631,N_11892);
and U12186 (N_12186,N_11993,N_11858);
nor U12187 (N_12187,N_11997,N_11930);
nor U12188 (N_12188,N_11746,N_11513);
nand U12189 (N_12189,N_11595,N_11630);
nor U12190 (N_12190,N_11665,N_11612);
or U12191 (N_12191,N_11879,N_11977);
nand U12192 (N_12192,N_11501,N_11768);
xnor U12193 (N_12193,N_11895,N_11979);
nand U12194 (N_12194,N_11803,N_11728);
nor U12195 (N_12195,N_11541,N_11527);
nor U12196 (N_12196,N_11830,N_11723);
or U12197 (N_12197,N_11995,N_11920);
nor U12198 (N_12198,N_11869,N_11724);
and U12199 (N_12199,N_11999,N_11903);
nand U12200 (N_12200,N_11700,N_11710);
and U12201 (N_12201,N_11502,N_11800);
and U12202 (N_12202,N_11759,N_11748);
or U12203 (N_12203,N_11568,N_11919);
nand U12204 (N_12204,N_11937,N_11935);
or U12205 (N_12205,N_11771,N_11899);
nor U12206 (N_12206,N_11610,N_11824);
and U12207 (N_12207,N_11807,N_11705);
nand U12208 (N_12208,N_11638,N_11596);
xor U12209 (N_12209,N_11913,N_11851);
and U12210 (N_12210,N_11849,N_11662);
xor U12211 (N_12211,N_11796,N_11659);
nor U12212 (N_12212,N_11754,N_11744);
xor U12213 (N_12213,N_11839,N_11562);
and U12214 (N_12214,N_11767,N_11555);
nand U12215 (N_12215,N_11575,N_11833);
or U12216 (N_12216,N_11990,N_11945);
and U12217 (N_12217,N_11729,N_11655);
nand U12218 (N_12218,N_11866,N_11891);
and U12219 (N_12219,N_11956,N_11615);
and U12220 (N_12220,N_11966,N_11812);
nand U12221 (N_12221,N_11900,N_11618);
nor U12222 (N_12222,N_11984,N_11508);
or U12223 (N_12223,N_11976,N_11519);
or U12224 (N_12224,N_11825,N_11951);
xnor U12225 (N_12225,N_11770,N_11902);
or U12226 (N_12226,N_11616,N_11686);
nor U12227 (N_12227,N_11624,N_11726);
nand U12228 (N_12228,N_11577,N_11967);
or U12229 (N_12229,N_11897,N_11735);
or U12230 (N_12230,N_11846,N_11998);
nand U12231 (N_12231,N_11963,N_11536);
nand U12232 (N_12232,N_11874,N_11889);
and U12233 (N_12233,N_11572,N_11952);
or U12234 (N_12234,N_11831,N_11763);
xnor U12235 (N_12235,N_11835,N_11893);
and U12236 (N_12236,N_11740,N_11757);
or U12237 (N_12237,N_11716,N_11944);
and U12238 (N_12238,N_11591,N_11795);
nand U12239 (N_12239,N_11528,N_11537);
nand U12240 (N_12240,N_11592,N_11713);
nor U12241 (N_12241,N_11847,N_11672);
and U12242 (N_12242,N_11987,N_11697);
xnor U12243 (N_12243,N_11751,N_11535);
nand U12244 (N_12244,N_11756,N_11948);
nand U12245 (N_12245,N_11801,N_11854);
and U12246 (N_12246,N_11602,N_11932);
nor U12247 (N_12247,N_11788,N_11743);
xor U12248 (N_12248,N_11764,N_11597);
nor U12249 (N_12249,N_11641,N_11518);
and U12250 (N_12250,N_11927,N_11649);
or U12251 (N_12251,N_11810,N_11930);
xor U12252 (N_12252,N_11838,N_11941);
or U12253 (N_12253,N_11757,N_11863);
and U12254 (N_12254,N_11844,N_11702);
nor U12255 (N_12255,N_11694,N_11561);
nor U12256 (N_12256,N_11762,N_11702);
and U12257 (N_12257,N_11585,N_11668);
and U12258 (N_12258,N_11582,N_11804);
xnor U12259 (N_12259,N_11692,N_11693);
or U12260 (N_12260,N_11688,N_11660);
or U12261 (N_12261,N_11680,N_11651);
or U12262 (N_12262,N_11632,N_11802);
or U12263 (N_12263,N_11557,N_11506);
nor U12264 (N_12264,N_11895,N_11789);
nand U12265 (N_12265,N_11715,N_11812);
or U12266 (N_12266,N_11549,N_11551);
xor U12267 (N_12267,N_11809,N_11733);
nand U12268 (N_12268,N_11554,N_11996);
and U12269 (N_12269,N_11547,N_11999);
or U12270 (N_12270,N_11987,N_11727);
xor U12271 (N_12271,N_11844,N_11593);
nand U12272 (N_12272,N_11924,N_11926);
xnor U12273 (N_12273,N_11981,N_11919);
xor U12274 (N_12274,N_11797,N_11528);
or U12275 (N_12275,N_11689,N_11883);
nor U12276 (N_12276,N_11824,N_11829);
and U12277 (N_12277,N_11948,N_11917);
or U12278 (N_12278,N_11923,N_11602);
nand U12279 (N_12279,N_11764,N_11838);
xor U12280 (N_12280,N_11511,N_11881);
nor U12281 (N_12281,N_11795,N_11663);
nand U12282 (N_12282,N_11670,N_11976);
nor U12283 (N_12283,N_11922,N_11860);
nor U12284 (N_12284,N_11794,N_11911);
xnor U12285 (N_12285,N_11735,N_11880);
and U12286 (N_12286,N_11999,N_11779);
nand U12287 (N_12287,N_11888,N_11673);
or U12288 (N_12288,N_11720,N_11749);
or U12289 (N_12289,N_11921,N_11787);
nor U12290 (N_12290,N_11546,N_11820);
nand U12291 (N_12291,N_11561,N_11879);
or U12292 (N_12292,N_11703,N_11914);
and U12293 (N_12293,N_11514,N_11783);
nor U12294 (N_12294,N_11539,N_11717);
xor U12295 (N_12295,N_11621,N_11792);
xor U12296 (N_12296,N_11740,N_11889);
or U12297 (N_12297,N_11871,N_11509);
nand U12298 (N_12298,N_11538,N_11780);
or U12299 (N_12299,N_11533,N_11882);
xor U12300 (N_12300,N_11587,N_11590);
nor U12301 (N_12301,N_11908,N_11729);
nand U12302 (N_12302,N_11552,N_11918);
or U12303 (N_12303,N_11543,N_11584);
nand U12304 (N_12304,N_11960,N_11503);
nor U12305 (N_12305,N_11865,N_11931);
nor U12306 (N_12306,N_11620,N_11977);
and U12307 (N_12307,N_11531,N_11673);
nor U12308 (N_12308,N_11845,N_11640);
nor U12309 (N_12309,N_11683,N_11938);
and U12310 (N_12310,N_11755,N_11539);
xnor U12311 (N_12311,N_11555,N_11596);
nand U12312 (N_12312,N_11805,N_11580);
nor U12313 (N_12313,N_11892,N_11973);
or U12314 (N_12314,N_11656,N_11653);
xor U12315 (N_12315,N_11825,N_11711);
or U12316 (N_12316,N_11708,N_11987);
nor U12317 (N_12317,N_11547,N_11695);
nor U12318 (N_12318,N_11710,N_11687);
nor U12319 (N_12319,N_11846,N_11806);
nor U12320 (N_12320,N_11988,N_11997);
and U12321 (N_12321,N_11981,N_11542);
and U12322 (N_12322,N_11821,N_11958);
or U12323 (N_12323,N_11600,N_11728);
nor U12324 (N_12324,N_11530,N_11527);
nand U12325 (N_12325,N_11568,N_11968);
or U12326 (N_12326,N_11719,N_11565);
and U12327 (N_12327,N_11863,N_11675);
nand U12328 (N_12328,N_11944,N_11595);
nor U12329 (N_12329,N_11545,N_11797);
and U12330 (N_12330,N_11997,N_11690);
nor U12331 (N_12331,N_11971,N_11905);
xor U12332 (N_12332,N_11541,N_11958);
nand U12333 (N_12333,N_11520,N_11763);
and U12334 (N_12334,N_11727,N_11758);
nand U12335 (N_12335,N_11903,N_11947);
xnor U12336 (N_12336,N_11591,N_11762);
and U12337 (N_12337,N_11587,N_11574);
or U12338 (N_12338,N_11824,N_11651);
nand U12339 (N_12339,N_11850,N_11599);
nor U12340 (N_12340,N_11506,N_11834);
or U12341 (N_12341,N_11973,N_11761);
xor U12342 (N_12342,N_11635,N_11815);
xnor U12343 (N_12343,N_11805,N_11629);
or U12344 (N_12344,N_11865,N_11567);
or U12345 (N_12345,N_11849,N_11581);
or U12346 (N_12346,N_11650,N_11774);
nand U12347 (N_12347,N_11686,N_11768);
and U12348 (N_12348,N_11901,N_11966);
xor U12349 (N_12349,N_11936,N_11747);
or U12350 (N_12350,N_11778,N_11838);
and U12351 (N_12351,N_11647,N_11645);
or U12352 (N_12352,N_11906,N_11707);
xor U12353 (N_12353,N_11948,N_11728);
nor U12354 (N_12354,N_11845,N_11627);
nor U12355 (N_12355,N_11893,N_11530);
xor U12356 (N_12356,N_11998,N_11502);
and U12357 (N_12357,N_11879,N_11928);
nand U12358 (N_12358,N_11652,N_11874);
nor U12359 (N_12359,N_11756,N_11518);
nor U12360 (N_12360,N_11943,N_11903);
or U12361 (N_12361,N_11768,N_11994);
or U12362 (N_12362,N_11717,N_11518);
or U12363 (N_12363,N_11600,N_11884);
xor U12364 (N_12364,N_11970,N_11840);
nand U12365 (N_12365,N_11774,N_11946);
and U12366 (N_12366,N_11898,N_11505);
xnor U12367 (N_12367,N_11822,N_11607);
nand U12368 (N_12368,N_11840,N_11889);
nand U12369 (N_12369,N_11995,N_11765);
xnor U12370 (N_12370,N_11756,N_11574);
xnor U12371 (N_12371,N_11817,N_11855);
or U12372 (N_12372,N_11981,N_11579);
nor U12373 (N_12373,N_11714,N_11925);
and U12374 (N_12374,N_11901,N_11509);
xor U12375 (N_12375,N_11818,N_11979);
or U12376 (N_12376,N_11952,N_11803);
or U12377 (N_12377,N_11749,N_11958);
nand U12378 (N_12378,N_11964,N_11743);
nand U12379 (N_12379,N_11934,N_11872);
or U12380 (N_12380,N_11760,N_11530);
and U12381 (N_12381,N_11879,N_11912);
and U12382 (N_12382,N_11917,N_11639);
and U12383 (N_12383,N_11568,N_11925);
nand U12384 (N_12384,N_11711,N_11888);
nand U12385 (N_12385,N_11807,N_11816);
nor U12386 (N_12386,N_11771,N_11897);
xor U12387 (N_12387,N_11873,N_11727);
nor U12388 (N_12388,N_11510,N_11875);
nand U12389 (N_12389,N_11694,N_11729);
and U12390 (N_12390,N_11622,N_11729);
nand U12391 (N_12391,N_11555,N_11795);
nand U12392 (N_12392,N_11785,N_11842);
nand U12393 (N_12393,N_11915,N_11551);
nand U12394 (N_12394,N_11654,N_11920);
or U12395 (N_12395,N_11719,N_11523);
and U12396 (N_12396,N_11540,N_11872);
xnor U12397 (N_12397,N_11909,N_11625);
and U12398 (N_12398,N_11810,N_11985);
nor U12399 (N_12399,N_11974,N_11558);
nor U12400 (N_12400,N_11925,N_11908);
nor U12401 (N_12401,N_11689,N_11846);
nor U12402 (N_12402,N_11864,N_11827);
and U12403 (N_12403,N_11999,N_11933);
or U12404 (N_12404,N_11625,N_11985);
nor U12405 (N_12405,N_11866,N_11741);
and U12406 (N_12406,N_11525,N_11754);
nand U12407 (N_12407,N_11662,N_11827);
nand U12408 (N_12408,N_11936,N_11559);
nand U12409 (N_12409,N_11554,N_11940);
nand U12410 (N_12410,N_11907,N_11775);
xor U12411 (N_12411,N_11523,N_11565);
or U12412 (N_12412,N_11633,N_11770);
nand U12413 (N_12413,N_11609,N_11734);
nor U12414 (N_12414,N_11796,N_11692);
nor U12415 (N_12415,N_11808,N_11615);
or U12416 (N_12416,N_11925,N_11822);
or U12417 (N_12417,N_11738,N_11905);
nor U12418 (N_12418,N_11952,N_11535);
nor U12419 (N_12419,N_11802,N_11975);
and U12420 (N_12420,N_11521,N_11661);
nand U12421 (N_12421,N_11817,N_11740);
xor U12422 (N_12422,N_11729,N_11747);
nor U12423 (N_12423,N_11580,N_11958);
and U12424 (N_12424,N_11518,N_11976);
nand U12425 (N_12425,N_11670,N_11694);
nor U12426 (N_12426,N_11643,N_11531);
and U12427 (N_12427,N_11875,N_11769);
and U12428 (N_12428,N_11935,N_11759);
or U12429 (N_12429,N_11523,N_11515);
or U12430 (N_12430,N_11858,N_11629);
or U12431 (N_12431,N_11543,N_11551);
xnor U12432 (N_12432,N_11827,N_11745);
xor U12433 (N_12433,N_11957,N_11557);
xor U12434 (N_12434,N_11905,N_11874);
or U12435 (N_12435,N_11705,N_11898);
nor U12436 (N_12436,N_11709,N_11774);
and U12437 (N_12437,N_11607,N_11845);
nor U12438 (N_12438,N_11802,N_11813);
and U12439 (N_12439,N_11874,N_11912);
and U12440 (N_12440,N_11772,N_11640);
nand U12441 (N_12441,N_11503,N_11576);
and U12442 (N_12442,N_11577,N_11927);
xnor U12443 (N_12443,N_11748,N_11549);
and U12444 (N_12444,N_11729,N_11708);
nor U12445 (N_12445,N_11616,N_11768);
and U12446 (N_12446,N_11714,N_11952);
or U12447 (N_12447,N_11828,N_11736);
and U12448 (N_12448,N_11765,N_11608);
and U12449 (N_12449,N_11751,N_11580);
xnor U12450 (N_12450,N_11503,N_11778);
or U12451 (N_12451,N_11886,N_11850);
and U12452 (N_12452,N_11732,N_11813);
xnor U12453 (N_12453,N_11897,N_11780);
xnor U12454 (N_12454,N_11855,N_11796);
xnor U12455 (N_12455,N_11519,N_11932);
nor U12456 (N_12456,N_11513,N_11807);
and U12457 (N_12457,N_11612,N_11849);
and U12458 (N_12458,N_11535,N_11636);
or U12459 (N_12459,N_11904,N_11512);
xnor U12460 (N_12460,N_11965,N_11813);
and U12461 (N_12461,N_11933,N_11654);
and U12462 (N_12462,N_11555,N_11788);
xnor U12463 (N_12463,N_11940,N_11505);
nand U12464 (N_12464,N_11773,N_11890);
or U12465 (N_12465,N_11605,N_11555);
and U12466 (N_12466,N_11716,N_11605);
nand U12467 (N_12467,N_11778,N_11756);
or U12468 (N_12468,N_11646,N_11619);
nor U12469 (N_12469,N_11952,N_11799);
xnor U12470 (N_12470,N_11680,N_11515);
xor U12471 (N_12471,N_11979,N_11906);
or U12472 (N_12472,N_11899,N_11994);
nand U12473 (N_12473,N_11848,N_11583);
and U12474 (N_12474,N_11836,N_11689);
and U12475 (N_12475,N_11721,N_11725);
and U12476 (N_12476,N_11986,N_11887);
or U12477 (N_12477,N_11624,N_11909);
nor U12478 (N_12478,N_11875,N_11593);
nand U12479 (N_12479,N_11601,N_11946);
and U12480 (N_12480,N_11690,N_11794);
or U12481 (N_12481,N_11581,N_11612);
xor U12482 (N_12482,N_11754,N_11861);
and U12483 (N_12483,N_11830,N_11737);
xor U12484 (N_12484,N_11953,N_11757);
nand U12485 (N_12485,N_11998,N_11696);
nor U12486 (N_12486,N_11715,N_11579);
or U12487 (N_12487,N_11520,N_11783);
or U12488 (N_12488,N_11506,N_11979);
nand U12489 (N_12489,N_11600,N_11694);
xnor U12490 (N_12490,N_11757,N_11931);
and U12491 (N_12491,N_11653,N_11553);
nor U12492 (N_12492,N_11687,N_11948);
and U12493 (N_12493,N_11543,N_11937);
nor U12494 (N_12494,N_11523,N_11617);
or U12495 (N_12495,N_11895,N_11823);
and U12496 (N_12496,N_11902,N_11998);
nand U12497 (N_12497,N_11632,N_11676);
nor U12498 (N_12498,N_11668,N_11654);
xnor U12499 (N_12499,N_11534,N_11807);
or U12500 (N_12500,N_12128,N_12405);
nor U12501 (N_12501,N_12332,N_12219);
nor U12502 (N_12502,N_12233,N_12062);
xnor U12503 (N_12503,N_12172,N_12455);
nand U12504 (N_12504,N_12127,N_12230);
nor U12505 (N_12505,N_12161,N_12149);
and U12506 (N_12506,N_12374,N_12220);
or U12507 (N_12507,N_12224,N_12483);
nor U12508 (N_12508,N_12415,N_12361);
xor U12509 (N_12509,N_12074,N_12002);
nand U12510 (N_12510,N_12153,N_12169);
nand U12511 (N_12511,N_12090,N_12493);
nor U12512 (N_12512,N_12260,N_12179);
xor U12513 (N_12513,N_12398,N_12178);
or U12514 (N_12514,N_12254,N_12404);
nand U12515 (N_12515,N_12466,N_12211);
and U12516 (N_12516,N_12018,N_12320);
nor U12517 (N_12517,N_12005,N_12333);
nor U12518 (N_12518,N_12006,N_12200);
nand U12519 (N_12519,N_12203,N_12016);
nor U12520 (N_12520,N_12151,N_12086);
and U12521 (N_12521,N_12221,N_12067);
nand U12522 (N_12522,N_12388,N_12034);
and U12523 (N_12523,N_12304,N_12119);
xnor U12524 (N_12524,N_12488,N_12070);
and U12525 (N_12525,N_12107,N_12206);
nand U12526 (N_12526,N_12307,N_12375);
and U12527 (N_12527,N_12245,N_12446);
and U12528 (N_12528,N_12343,N_12464);
and U12529 (N_12529,N_12058,N_12420);
or U12530 (N_12530,N_12401,N_12222);
nor U12531 (N_12531,N_12399,N_12436);
nand U12532 (N_12532,N_12449,N_12369);
and U12533 (N_12533,N_12474,N_12184);
xnor U12534 (N_12534,N_12066,N_12093);
xnor U12535 (N_12535,N_12476,N_12035);
nand U12536 (N_12536,N_12424,N_12323);
nor U12537 (N_12537,N_12114,N_12285);
nand U12538 (N_12538,N_12370,N_12262);
nand U12539 (N_12539,N_12444,N_12064);
xor U12540 (N_12540,N_12024,N_12213);
xor U12541 (N_12541,N_12232,N_12299);
nor U12542 (N_12542,N_12118,N_12156);
xor U12543 (N_12543,N_12252,N_12037);
xnor U12544 (N_12544,N_12341,N_12095);
nand U12545 (N_12545,N_12409,N_12318);
or U12546 (N_12546,N_12004,N_12044);
or U12547 (N_12547,N_12251,N_12204);
nor U12548 (N_12548,N_12432,N_12365);
or U12549 (N_12549,N_12463,N_12092);
nor U12550 (N_12550,N_12228,N_12435);
or U12551 (N_12551,N_12180,N_12396);
nor U12552 (N_12552,N_12352,N_12126);
or U12553 (N_12553,N_12083,N_12194);
or U12554 (N_12554,N_12467,N_12407);
nor U12555 (N_12555,N_12380,N_12280);
nor U12556 (N_12556,N_12071,N_12327);
nand U12557 (N_12557,N_12088,N_12000);
or U12558 (N_12558,N_12344,N_12244);
nand U12559 (N_12559,N_12185,N_12082);
nand U12560 (N_12560,N_12163,N_12102);
nand U12561 (N_12561,N_12052,N_12363);
nor U12562 (N_12562,N_12054,N_12196);
nor U12563 (N_12563,N_12250,N_12417);
or U12564 (N_12564,N_12395,N_12322);
and U12565 (N_12565,N_12281,N_12135);
nand U12566 (N_12566,N_12342,N_12356);
and U12567 (N_12567,N_12300,N_12340);
or U12568 (N_12568,N_12081,N_12084);
nand U12569 (N_12569,N_12142,N_12421);
xnor U12570 (N_12570,N_12215,N_12094);
nand U12571 (N_12571,N_12195,N_12419);
xor U12572 (N_12572,N_12129,N_12314);
nor U12573 (N_12573,N_12468,N_12392);
or U12574 (N_12574,N_12096,N_12237);
nand U12575 (N_12575,N_12471,N_12461);
nor U12576 (N_12576,N_12031,N_12288);
nand U12577 (N_12577,N_12047,N_12039);
nor U12578 (N_12578,N_12345,N_12303);
nor U12579 (N_12579,N_12384,N_12267);
xor U12580 (N_12580,N_12315,N_12110);
nand U12581 (N_12581,N_12248,N_12073);
and U12582 (N_12582,N_12470,N_12347);
nor U12583 (N_12583,N_12182,N_12326);
xnor U12584 (N_12584,N_12486,N_12152);
and U12585 (N_12585,N_12227,N_12485);
nor U12586 (N_12586,N_12150,N_12275);
and U12587 (N_12587,N_12255,N_12160);
xor U12588 (N_12588,N_12351,N_12124);
or U12589 (N_12589,N_12489,N_12240);
nor U12590 (N_12590,N_12492,N_12494);
and U12591 (N_12591,N_12116,N_12413);
or U12592 (N_12592,N_12353,N_12430);
nor U12593 (N_12593,N_12176,N_12140);
or U12594 (N_12594,N_12181,N_12308);
nor U12595 (N_12595,N_12208,N_12137);
or U12596 (N_12596,N_12033,N_12246);
or U12597 (N_12597,N_12372,N_12239);
and U12598 (N_12598,N_12197,N_12162);
nand U12599 (N_12599,N_12480,N_12367);
nand U12600 (N_12600,N_12258,N_12259);
or U12601 (N_12601,N_12223,N_12427);
nand U12602 (N_12602,N_12063,N_12324);
nor U12603 (N_12603,N_12115,N_12433);
or U12604 (N_12604,N_12053,N_12168);
nor U12605 (N_12605,N_12329,N_12029);
or U12606 (N_12606,N_12045,N_12236);
nor U12607 (N_12607,N_12061,N_12048);
or U12608 (N_12608,N_12101,N_12377);
nor U12609 (N_12609,N_12431,N_12484);
or U12610 (N_12610,N_12191,N_12122);
xnor U12611 (N_12611,N_12041,N_12282);
or U12612 (N_12612,N_12337,N_12386);
and U12613 (N_12613,N_12012,N_12289);
nor U12614 (N_12614,N_12112,N_12458);
or U12615 (N_12615,N_12261,N_12364);
xor U12616 (N_12616,N_12306,N_12186);
nand U12617 (N_12617,N_12271,N_12036);
or U12618 (N_12618,N_12428,N_12187);
and U12619 (N_12619,N_12060,N_12298);
nor U12620 (N_12620,N_12445,N_12270);
or U12621 (N_12621,N_12042,N_12411);
nand U12622 (N_12622,N_12212,N_12279);
and U12623 (N_12623,N_12422,N_12105);
and U12624 (N_12624,N_12193,N_12123);
and U12625 (N_12625,N_12269,N_12015);
or U12626 (N_12626,N_12309,N_12389);
nor U12627 (N_12627,N_12418,N_12454);
nand U12628 (N_12628,N_12216,N_12429);
nor U12629 (N_12629,N_12338,N_12209);
and U12630 (N_12630,N_12192,N_12391);
or U12631 (N_12631,N_12297,N_12134);
and U12632 (N_12632,N_12362,N_12014);
or U12633 (N_12633,N_12008,N_12201);
and U12634 (N_12634,N_12055,N_12473);
xnor U12635 (N_12635,N_12078,N_12190);
or U12636 (N_12636,N_12174,N_12453);
or U12637 (N_12637,N_12423,N_12284);
xor U12638 (N_12638,N_12143,N_12098);
xnor U12639 (N_12639,N_12167,N_12416);
and U12640 (N_12640,N_12079,N_12497);
and U12641 (N_12641,N_12155,N_12225);
xor U12642 (N_12642,N_12108,N_12013);
xnor U12643 (N_12643,N_12019,N_12460);
and U12644 (N_12644,N_12076,N_12264);
xnor U12645 (N_12645,N_12166,N_12482);
xnor U12646 (N_12646,N_12130,N_12243);
nor U12647 (N_12647,N_12434,N_12104);
nand U12648 (N_12648,N_12080,N_12120);
nor U12649 (N_12649,N_12443,N_12056);
xnor U12650 (N_12650,N_12003,N_12028);
nor U12651 (N_12651,N_12366,N_12390);
xnor U12652 (N_12652,N_12478,N_12009);
xor U12653 (N_12653,N_12157,N_12205);
and U12654 (N_12654,N_12348,N_12441);
and U12655 (N_12655,N_12292,N_12358);
nand U12656 (N_12656,N_12334,N_12360);
nor U12657 (N_12657,N_12136,N_12310);
xor U12658 (N_12658,N_12450,N_12376);
nor U12659 (N_12659,N_12164,N_12350);
xor U12660 (N_12660,N_12010,N_12030);
and U12661 (N_12661,N_12026,N_12368);
xor U12662 (N_12662,N_12226,N_12100);
xnor U12663 (N_12663,N_12043,N_12290);
xor U12664 (N_12664,N_12472,N_12456);
nand U12665 (N_12665,N_12465,N_12025);
xnor U12666 (N_12666,N_12188,N_12017);
nor U12667 (N_12667,N_12498,N_12448);
nor U12668 (N_12668,N_12402,N_12229);
or U12669 (N_12669,N_12381,N_12286);
and U12670 (N_12670,N_12406,N_12218);
or U12671 (N_12671,N_12394,N_12316);
and U12672 (N_12672,N_12051,N_12354);
nand U12673 (N_12673,N_12346,N_12040);
xor U12674 (N_12674,N_12274,N_12177);
xor U12675 (N_12675,N_12335,N_12385);
xnor U12676 (N_12676,N_12378,N_12089);
nand U12677 (N_12677,N_12302,N_12214);
and U12678 (N_12678,N_12159,N_12027);
xnor U12679 (N_12679,N_12171,N_12442);
nand U12680 (N_12680,N_12106,N_12393);
or U12681 (N_12681,N_12247,N_12154);
or U12682 (N_12682,N_12312,N_12451);
nand U12683 (N_12683,N_12400,N_12139);
nor U12684 (N_12684,N_12241,N_12481);
and U12685 (N_12685,N_12103,N_12234);
xnor U12686 (N_12686,N_12069,N_12132);
and U12687 (N_12687,N_12414,N_12452);
xnor U12688 (N_12688,N_12145,N_12294);
xor U12689 (N_12689,N_12131,N_12479);
or U12690 (N_12690,N_12469,N_12278);
nand U12691 (N_12691,N_12263,N_12057);
nor U12692 (N_12692,N_12059,N_12272);
or U12693 (N_12693,N_12266,N_12147);
and U12694 (N_12694,N_12256,N_12148);
xnor U12695 (N_12695,N_12277,N_12170);
nand U12696 (N_12696,N_12437,N_12085);
nand U12697 (N_12697,N_12109,N_12426);
or U12698 (N_12698,N_12291,N_12499);
nor U12699 (N_12699,N_12295,N_12235);
or U12700 (N_12700,N_12001,N_12487);
xnor U12701 (N_12701,N_12242,N_12077);
or U12702 (N_12702,N_12382,N_12412);
nand U12703 (N_12703,N_12273,N_12495);
xnor U12704 (N_12704,N_12183,N_12189);
nand U12705 (N_12705,N_12317,N_12410);
nand U12706 (N_12706,N_12068,N_12099);
and U12707 (N_12707,N_12355,N_12023);
nand U12708 (N_12708,N_12117,N_12268);
nor U12709 (N_12709,N_12091,N_12440);
or U12710 (N_12710,N_12328,N_12146);
nand U12711 (N_12711,N_12438,N_12447);
and U12712 (N_12712,N_12325,N_12425);
nand U12713 (N_12713,N_12202,N_12339);
or U12714 (N_12714,N_12283,N_12199);
and U12715 (N_12715,N_12125,N_12198);
xnor U12716 (N_12716,N_12383,N_12373);
xor U12717 (N_12717,N_12020,N_12097);
or U12718 (N_12718,N_12477,N_12231);
nor U12719 (N_12719,N_12021,N_12439);
nand U12720 (N_12720,N_12462,N_12011);
or U12721 (N_12721,N_12144,N_12371);
and U12722 (N_12722,N_12457,N_12330);
and U12723 (N_12723,N_12038,N_12113);
and U12724 (N_12724,N_12049,N_12359);
xnor U12725 (N_12725,N_12257,N_12065);
or U12726 (N_12726,N_12301,N_12305);
nand U12727 (N_12727,N_12490,N_12287);
or U12728 (N_12728,N_12387,N_12072);
xnor U12729 (N_12729,N_12087,N_12321);
xor U12730 (N_12730,N_12217,N_12397);
nor U12731 (N_12731,N_12475,N_12357);
or U12732 (N_12732,N_12046,N_12138);
and U12733 (N_12733,N_12459,N_12379);
xnor U12734 (N_12734,N_12408,N_12050);
nand U12735 (N_12735,N_12238,N_12311);
or U12736 (N_12736,N_12293,N_12265);
nand U12737 (N_12737,N_12403,N_12032);
nand U12738 (N_12738,N_12133,N_12158);
and U12739 (N_12739,N_12331,N_12007);
and U12740 (N_12740,N_12141,N_12336);
and U12741 (N_12741,N_12349,N_12496);
nor U12742 (N_12742,N_12319,N_12165);
nand U12743 (N_12743,N_12022,N_12210);
nor U12744 (N_12744,N_12249,N_12276);
nor U12745 (N_12745,N_12173,N_12253);
and U12746 (N_12746,N_12491,N_12175);
or U12747 (N_12747,N_12313,N_12296);
nor U12748 (N_12748,N_12121,N_12207);
xnor U12749 (N_12749,N_12111,N_12075);
xor U12750 (N_12750,N_12482,N_12226);
nor U12751 (N_12751,N_12431,N_12417);
nand U12752 (N_12752,N_12118,N_12137);
xor U12753 (N_12753,N_12286,N_12484);
and U12754 (N_12754,N_12045,N_12210);
and U12755 (N_12755,N_12255,N_12459);
nor U12756 (N_12756,N_12065,N_12013);
or U12757 (N_12757,N_12476,N_12496);
xor U12758 (N_12758,N_12420,N_12343);
xnor U12759 (N_12759,N_12080,N_12433);
or U12760 (N_12760,N_12367,N_12469);
or U12761 (N_12761,N_12491,N_12450);
and U12762 (N_12762,N_12462,N_12307);
nand U12763 (N_12763,N_12449,N_12403);
nand U12764 (N_12764,N_12004,N_12173);
or U12765 (N_12765,N_12274,N_12357);
or U12766 (N_12766,N_12187,N_12026);
xnor U12767 (N_12767,N_12087,N_12253);
or U12768 (N_12768,N_12182,N_12335);
nor U12769 (N_12769,N_12055,N_12416);
and U12770 (N_12770,N_12219,N_12403);
nand U12771 (N_12771,N_12094,N_12365);
and U12772 (N_12772,N_12118,N_12299);
and U12773 (N_12773,N_12121,N_12111);
nor U12774 (N_12774,N_12078,N_12304);
xnor U12775 (N_12775,N_12174,N_12019);
xor U12776 (N_12776,N_12124,N_12435);
nand U12777 (N_12777,N_12370,N_12299);
xnor U12778 (N_12778,N_12103,N_12222);
nor U12779 (N_12779,N_12444,N_12324);
and U12780 (N_12780,N_12028,N_12126);
or U12781 (N_12781,N_12155,N_12290);
nand U12782 (N_12782,N_12160,N_12446);
nor U12783 (N_12783,N_12351,N_12167);
xnor U12784 (N_12784,N_12182,N_12145);
or U12785 (N_12785,N_12099,N_12047);
nor U12786 (N_12786,N_12482,N_12302);
nor U12787 (N_12787,N_12199,N_12147);
and U12788 (N_12788,N_12011,N_12082);
nor U12789 (N_12789,N_12178,N_12148);
and U12790 (N_12790,N_12403,N_12092);
or U12791 (N_12791,N_12412,N_12061);
nor U12792 (N_12792,N_12138,N_12129);
and U12793 (N_12793,N_12377,N_12016);
nor U12794 (N_12794,N_12237,N_12344);
and U12795 (N_12795,N_12196,N_12298);
and U12796 (N_12796,N_12012,N_12035);
nor U12797 (N_12797,N_12396,N_12142);
xor U12798 (N_12798,N_12362,N_12307);
nor U12799 (N_12799,N_12111,N_12020);
or U12800 (N_12800,N_12042,N_12301);
nand U12801 (N_12801,N_12241,N_12014);
or U12802 (N_12802,N_12302,N_12466);
xnor U12803 (N_12803,N_12204,N_12132);
nand U12804 (N_12804,N_12355,N_12159);
xnor U12805 (N_12805,N_12021,N_12285);
nor U12806 (N_12806,N_12164,N_12361);
and U12807 (N_12807,N_12000,N_12148);
or U12808 (N_12808,N_12474,N_12138);
nand U12809 (N_12809,N_12373,N_12275);
and U12810 (N_12810,N_12493,N_12435);
and U12811 (N_12811,N_12247,N_12400);
nor U12812 (N_12812,N_12263,N_12139);
xor U12813 (N_12813,N_12408,N_12414);
xor U12814 (N_12814,N_12431,N_12429);
nand U12815 (N_12815,N_12407,N_12390);
and U12816 (N_12816,N_12415,N_12386);
or U12817 (N_12817,N_12326,N_12409);
xor U12818 (N_12818,N_12028,N_12320);
or U12819 (N_12819,N_12362,N_12137);
or U12820 (N_12820,N_12464,N_12059);
nand U12821 (N_12821,N_12427,N_12241);
xnor U12822 (N_12822,N_12001,N_12286);
xor U12823 (N_12823,N_12307,N_12459);
nor U12824 (N_12824,N_12013,N_12428);
or U12825 (N_12825,N_12487,N_12041);
and U12826 (N_12826,N_12346,N_12297);
xor U12827 (N_12827,N_12140,N_12274);
or U12828 (N_12828,N_12205,N_12464);
nand U12829 (N_12829,N_12036,N_12491);
xnor U12830 (N_12830,N_12468,N_12498);
and U12831 (N_12831,N_12242,N_12216);
or U12832 (N_12832,N_12111,N_12257);
nor U12833 (N_12833,N_12278,N_12131);
xor U12834 (N_12834,N_12484,N_12281);
nor U12835 (N_12835,N_12003,N_12431);
nand U12836 (N_12836,N_12418,N_12063);
or U12837 (N_12837,N_12040,N_12267);
nand U12838 (N_12838,N_12370,N_12177);
or U12839 (N_12839,N_12452,N_12157);
or U12840 (N_12840,N_12220,N_12148);
and U12841 (N_12841,N_12385,N_12343);
nand U12842 (N_12842,N_12362,N_12005);
nor U12843 (N_12843,N_12010,N_12125);
nand U12844 (N_12844,N_12460,N_12445);
and U12845 (N_12845,N_12038,N_12175);
xor U12846 (N_12846,N_12333,N_12169);
nand U12847 (N_12847,N_12412,N_12110);
or U12848 (N_12848,N_12157,N_12334);
and U12849 (N_12849,N_12316,N_12434);
nor U12850 (N_12850,N_12073,N_12063);
nand U12851 (N_12851,N_12050,N_12401);
nand U12852 (N_12852,N_12222,N_12142);
nand U12853 (N_12853,N_12198,N_12118);
xor U12854 (N_12854,N_12186,N_12259);
nor U12855 (N_12855,N_12008,N_12246);
and U12856 (N_12856,N_12073,N_12395);
or U12857 (N_12857,N_12097,N_12370);
nand U12858 (N_12858,N_12489,N_12170);
xnor U12859 (N_12859,N_12275,N_12187);
or U12860 (N_12860,N_12274,N_12355);
xnor U12861 (N_12861,N_12040,N_12246);
nor U12862 (N_12862,N_12365,N_12193);
nor U12863 (N_12863,N_12159,N_12171);
nor U12864 (N_12864,N_12340,N_12316);
xnor U12865 (N_12865,N_12277,N_12434);
nor U12866 (N_12866,N_12427,N_12025);
and U12867 (N_12867,N_12148,N_12325);
nand U12868 (N_12868,N_12490,N_12355);
and U12869 (N_12869,N_12298,N_12339);
xnor U12870 (N_12870,N_12147,N_12094);
nand U12871 (N_12871,N_12254,N_12092);
xnor U12872 (N_12872,N_12025,N_12279);
nor U12873 (N_12873,N_12443,N_12155);
nand U12874 (N_12874,N_12344,N_12401);
nand U12875 (N_12875,N_12016,N_12447);
nor U12876 (N_12876,N_12049,N_12477);
and U12877 (N_12877,N_12155,N_12002);
nor U12878 (N_12878,N_12108,N_12430);
xor U12879 (N_12879,N_12219,N_12089);
xnor U12880 (N_12880,N_12341,N_12059);
nand U12881 (N_12881,N_12035,N_12424);
or U12882 (N_12882,N_12415,N_12185);
or U12883 (N_12883,N_12064,N_12066);
xor U12884 (N_12884,N_12045,N_12162);
and U12885 (N_12885,N_12304,N_12406);
or U12886 (N_12886,N_12077,N_12280);
nand U12887 (N_12887,N_12037,N_12192);
and U12888 (N_12888,N_12443,N_12285);
nor U12889 (N_12889,N_12158,N_12024);
xnor U12890 (N_12890,N_12245,N_12448);
nand U12891 (N_12891,N_12066,N_12036);
xnor U12892 (N_12892,N_12345,N_12432);
nor U12893 (N_12893,N_12096,N_12228);
nor U12894 (N_12894,N_12300,N_12467);
or U12895 (N_12895,N_12064,N_12495);
nand U12896 (N_12896,N_12004,N_12228);
nor U12897 (N_12897,N_12275,N_12213);
nand U12898 (N_12898,N_12178,N_12412);
or U12899 (N_12899,N_12367,N_12035);
xor U12900 (N_12900,N_12279,N_12149);
xor U12901 (N_12901,N_12201,N_12130);
or U12902 (N_12902,N_12058,N_12330);
or U12903 (N_12903,N_12241,N_12336);
or U12904 (N_12904,N_12310,N_12289);
and U12905 (N_12905,N_12423,N_12358);
nor U12906 (N_12906,N_12193,N_12279);
or U12907 (N_12907,N_12324,N_12266);
nor U12908 (N_12908,N_12280,N_12045);
and U12909 (N_12909,N_12331,N_12167);
or U12910 (N_12910,N_12375,N_12271);
and U12911 (N_12911,N_12406,N_12214);
nand U12912 (N_12912,N_12353,N_12408);
nand U12913 (N_12913,N_12180,N_12458);
nand U12914 (N_12914,N_12454,N_12228);
nand U12915 (N_12915,N_12192,N_12489);
and U12916 (N_12916,N_12128,N_12382);
nand U12917 (N_12917,N_12037,N_12181);
and U12918 (N_12918,N_12345,N_12046);
nor U12919 (N_12919,N_12259,N_12419);
xnor U12920 (N_12920,N_12300,N_12491);
xor U12921 (N_12921,N_12082,N_12123);
xor U12922 (N_12922,N_12201,N_12000);
nor U12923 (N_12923,N_12311,N_12129);
nor U12924 (N_12924,N_12441,N_12017);
nor U12925 (N_12925,N_12434,N_12328);
xnor U12926 (N_12926,N_12242,N_12241);
or U12927 (N_12927,N_12191,N_12008);
and U12928 (N_12928,N_12184,N_12230);
xor U12929 (N_12929,N_12048,N_12374);
and U12930 (N_12930,N_12487,N_12470);
nor U12931 (N_12931,N_12340,N_12442);
xnor U12932 (N_12932,N_12334,N_12064);
xor U12933 (N_12933,N_12124,N_12234);
or U12934 (N_12934,N_12131,N_12321);
xor U12935 (N_12935,N_12046,N_12398);
nor U12936 (N_12936,N_12019,N_12242);
nor U12937 (N_12937,N_12149,N_12176);
nand U12938 (N_12938,N_12133,N_12015);
or U12939 (N_12939,N_12390,N_12100);
nand U12940 (N_12940,N_12106,N_12160);
or U12941 (N_12941,N_12269,N_12295);
and U12942 (N_12942,N_12429,N_12138);
or U12943 (N_12943,N_12423,N_12166);
and U12944 (N_12944,N_12204,N_12413);
and U12945 (N_12945,N_12490,N_12282);
and U12946 (N_12946,N_12412,N_12109);
and U12947 (N_12947,N_12419,N_12055);
and U12948 (N_12948,N_12185,N_12403);
and U12949 (N_12949,N_12317,N_12427);
nand U12950 (N_12950,N_12468,N_12423);
xnor U12951 (N_12951,N_12448,N_12011);
nand U12952 (N_12952,N_12376,N_12211);
xnor U12953 (N_12953,N_12461,N_12356);
or U12954 (N_12954,N_12263,N_12075);
and U12955 (N_12955,N_12344,N_12351);
nor U12956 (N_12956,N_12277,N_12299);
nor U12957 (N_12957,N_12155,N_12223);
and U12958 (N_12958,N_12414,N_12014);
or U12959 (N_12959,N_12063,N_12046);
nor U12960 (N_12960,N_12476,N_12355);
nor U12961 (N_12961,N_12368,N_12075);
nor U12962 (N_12962,N_12158,N_12029);
xor U12963 (N_12963,N_12203,N_12008);
and U12964 (N_12964,N_12478,N_12002);
nor U12965 (N_12965,N_12287,N_12283);
xor U12966 (N_12966,N_12273,N_12384);
nand U12967 (N_12967,N_12439,N_12301);
nor U12968 (N_12968,N_12383,N_12143);
xor U12969 (N_12969,N_12143,N_12497);
or U12970 (N_12970,N_12065,N_12056);
nand U12971 (N_12971,N_12479,N_12197);
nand U12972 (N_12972,N_12213,N_12007);
and U12973 (N_12973,N_12145,N_12220);
or U12974 (N_12974,N_12281,N_12305);
nand U12975 (N_12975,N_12265,N_12140);
or U12976 (N_12976,N_12326,N_12046);
and U12977 (N_12977,N_12166,N_12038);
and U12978 (N_12978,N_12473,N_12004);
or U12979 (N_12979,N_12325,N_12097);
and U12980 (N_12980,N_12497,N_12444);
xnor U12981 (N_12981,N_12079,N_12146);
or U12982 (N_12982,N_12463,N_12218);
nand U12983 (N_12983,N_12034,N_12070);
xnor U12984 (N_12984,N_12312,N_12094);
or U12985 (N_12985,N_12073,N_12354);
and U12986 (N_12986,N_12499,N_12255);
xnor U12987 (N_12987,N_12022,N_12298);
xor U12988 (N_12988,N_12300,N_12119);
and U12989 (N_12989,N_12476,N_12366);
nand U12990 (N_12990,N_12384,N_12323);
or U12991 (N_12991,N_12368,N_12017);
and U12992 (N_12992,N_12458,N_12408);
nand U12993 (N_12993,N_12190,N_12328);
nor U12994 (N_12994,N_12103,N_12371);
and U12995 (N_12995,N_12232,N_12039);
xor U12996 (N_12996,N_12270,N_12215);
nand U12997 (N_12997,N_12014,N_12267);
xnor U12998 (N_12998,N_12183,N_12291);
and U12999 (N_12999,N_12368,N_12448);
nor U13000 (N_13000,N_12637,N_12983);
or U13001 (N_13001,N_12635,N_12749);
nor U13002 (N_13002,N_12837,N_12632);
and U13003 (N_13003,N_12543,N_12850);
xor U13004 (N_13004,N_12709,N_12722);
xor U13005 (N_13005,N_12502,N_12613);
and U13006 (N_13006,N_12644,N_12582);
or U13007 (N_13007,N_12575,N_12534);
xor U13008 (N_13008,N_12861,N_12563);
nand U13009 (N_13009,N_12938,N_12648);
nor U13010 (N_13010,N_12597,N_12995);
xor U13011 (N_13011,N_12514,N_12858);
nor U13012 (N_13012,N_12803,N_12794);
xnor U13013 (N_13013,N_12706,N_12616);
nand U13014 (N_13014,N_12974,N_12897);
nor U13015 (N_13015,N_12958,N_12509);
and U13016 (N_13016,N_12647,N_12584);
nor U13017 (N_13017,N_12999,N_12568);
nor U13018 (N_13018,N_12501,N_12868);
nand U13019 (N_13019,N_12962,N_12838);
nor U13020 (N_13020,N_12788,N_12927);
nand U13021 (N_13021,N_12924,N_12660);
and U13022 (N_13022,N_12881,N_12907);
or U13023 (N_13023,N_12691,N_12940);
and U13024 (N_13024,N_12775,N_12664);
nand U13025 (N_13025,N_12966,N_12835);
nor U13026 (N_13026,N_12614,N_12930);
or U13027 (N_13027,N_12679,N_12681);
xnor U13028 (N_13028,N_12885,N_12760);
nor U13029 (N_13029,N_12612,N_12580);
nor U13030 (N_13030,N_12828,N_12781);
or U13031 (N_13031,N_12730,N_12887);
nand U13032 (N_13032,N_12948,N_12620);
nor U13033 (N_13033,N_12586,N_12809);
xor U13034 (N_13034,N_12685,N_12845);
or U13035 (N_13035,N_12830,N_12530);
nor U13036 (N_13036,N_12834,N_12800);
nor U13037 (N_13037,N_12742,N_12891);
and U13038 (N_13038,N_12822,N_12776);
xnor U13039 (N_13039,N_12998,N_12553);
or U13040 (N_13040,N_12625,N_12546);
nor U13041 (N_13041,N_12994,N_12646);
or U13042 (N_13042,N_12947,N_12980);
nand U13043 (N_13043,N_12990,N_12954);
nor U13044 (N_13044,N_12871,N_12951);
and U13045 (N_13045,N_12622,N_12753);
xnor U13046 (N_13046,N_12957,N_12880);
or U13047 (N_13047,N_12883,N_12799);
or U13048 (N_13048,N_12665,N_12555);
xnor U13049 (N_13049,N_12655,N_12945);
nand U13050 (N_13050,N_12738,N_12988);
nor U13051 (N_13051,N_12922,N_12900);
xnor U13052 (N_13052,N_12903,N_12688);
nand U13053 (N_13053,N_12524,N_12905);
or U13054 (N_13054,N_12937,N_12624);
and U13055 (N_13055,N_12987,N_12517);
or U13056 (N_13056,N_12968,N_12511);
nand U13057 (N_13057,N_12535,N_12591);
xor U13058 (N_13058,N_12574,N_12592);
and U13059 (N_13059,N_12588,N_12904);
and U13060 (N_13060,N_12906,N_12703);
xnor U13061 (N_13061,N_12997,N_12793);
and U13062 (N_13062,N_12728,N_12545);
nor U13063 (N_13063,N_12559,N_12532);
xor U13064 (N_13064,N_12806,N_12716);
xor U13065 (N_13065,N_12542,N_12908);
nor U13066 (N_13066,N_12508,N_12626);
nand U13067 (N_13067,N_12836,N_12857);
or U13068 (N_13068,N_12662,N_12638);
nand U13069 (N_13069,N_12692,N_12767);
and U13070 (N_13070,N_12770,N_12578);
xor U13071 (N_13071,N_12715,N_12931);
nand U13072 (N_13072,N_12864,N_12663);
xnor U13073 (N_13073,N_12736,N_12566);
nand U13074 (N_13074,N_12923,N_12533);
xnor U13075 (N_13075,N_12570,N_12627);
or U13076 (N_13076,N_12824,N_12640);
or U13077 (N_13077,N_12743,N_12755);
nand U13078 (N_13078,N_12562,N_12785);
nor U13079 (N_13079,N_12636,N_12986);
or U13080 (N_13080,N_12724,N_12848);
and U13081 (N_13081,N_12979,N_12551);
nor U13082 (N_13082,N_12550,N_12634);
xnor U13083 (N_13083,N_12929,N_12946);
nand U13084 (N_13084,N_12720,N_12593);
or U13085 (N_13085,N_12961,N_12820);
and U13086 (N_13086,N_12859,N_12500);
nor U13087 (N_13087,N_12590,N_12518);
and U13088 (N_13088,N_12710,N_12842);
nand U13089 (N_13089,N_12888,N_12818);
xor U13090 (N_13090,N_12713,N_12911);
or U13091 (N_13091,N_12917,N_12963);
and U13092 (N_13092,N_12519,N_12970);
nor U13093 (N_13093,N_12723,N_12512);
or U13094 (N_13094,N_12798,N_12942);
nand U13095 (N_13095,N_12727,N_12873);
and U13096 (N_13096,N_12556,N_12919);
or U13097 (N_13097,N_12839,N_12629);
nand U13098 (N_13098,N_12933,N_12801);
nand U13099 (N_13099,N_12650,N_12916);
xor U13100 (N_13100,N_12813,N_12950);
or U13101 (N_13101,N_12771,N_12693);
nand U13102 (N_13102,N_12805,N_12510);
and U13103 (N_13103,N_12571,N_12814);
or U13104 (N_13104,N_12827,N_12811);
xor U13105 (N_13105,N_12847,N_12649);
xnor U13106 (N_13106,N_12695,N_12522);
or U13107 (N_13107,N_12833,N_12768);
nor U13108 (N_13108,N_12505,N_12955);
nand U13109 (N_13109,N_12964,N_12849);
or U13110 (N_13110,N_12589,N_12527);
nor U13111 (N_13111,N_12577,N_12969);
or U13112 (N_13112,N_12934,N_12658);
and U13113 (N_13113,N_12603,N_12712);
nor U13114 (N_13114,N_12796,N_12773);
and U13115 (N_13115,N_12876,N_12554);
xnor U13116 (N_13116,N_12744,N_12783);
and U13117 (N_13117,N_12686,N_12884);
or U13118 (N_13118,N_12764,N_12564);
xor U13119 (N_13119,N_12867,N_12735);
and U13120 (N_13120,N_12774,N_12921);
and U13121 (N_13121,N_12993,N_12886);
nor U13122 (N_13122,N_12701,N_12872);
nand U13123 (N_13123,N_12879,N_12698);
and U13124 (N_13124,N_12526,N_12666);
xnor U13125 (N_13125,N_12856,N_12531);
nand U13126 (N_13126,N_12549,N_12734);
or U13127 (N_13127,N_12521,N_12717);
xnor U13128 (N_13128,N_12504,N_12795);
nand U13129 (N_13129,N_12972,N_12976);
xnor U13130 (N_13130,N_12731,N_12894);
nand U13131 (N_13131,N_12996,N_12746);
xor U13132 (N_13132,N_12901,N_12875);
xor U13133 (N_13133,N_12780,N_12892);
nor U13134 (N_13134,N_12747,N_12729);
xor U13135 (N_13135,N_12608,N_12628);
or U13136 (N_13136,N_12538,N_12611);
nor U13137 (N_13137,N_12936,N_12765);
and U13138 (N_13138,N_12910,N_12802);
and U13139 (N_13139,N_12769,N_12960);
nand U13140 (N_13140,N_12756,N_12704);
or U13141 (N_13141,N_12617,N_12725);
nand U13142 (N_13142,N_12677,N_12699);
or U13143 (N_13143,N_12877,N_12825);
nand U13144 (N_13144,N_12569,N_12610);
nor U13145 (N_13145,N_12890,N_12654);
nor U13146 (N_13146,N_12804,N_12866);
and U13147 (N_13147,N_12544,N_12581);
and U13148 (N_13148,N_12815,N_12705);
nand U13149 (N_13149,N_12823,N_12855);
xnor U13150 (N_13150,N_12935,N_12895);
and U13151 (N_13151,N_12596,N_12992);
nor U13152 (N_13152,N_12507,N_12784);
nor U13153 (N_13153,N_12618,N_12808);
nor U13154 (N_13154,N_12941,N_12939);
xnor U13155 (N_13155,N_12882,N_12560);
or U13156 (N_13156,N_12754,N_12841);
nor U13157 (N_13157,N_12851,N_12675);
nor U13158 (N_13158,N_12684,N_12630);
xor U13159 (N_13159,N_12680,N_12503);
nand U13160 (N_13160,N_12982,N_12557);
xnor U13161 (N_13161,N_12971,N_12641);
nor U13162 (N_13162,N_12778,N_12846);
nor U13163 (N_13163,N_12757,N_12810);
and U13164 (N_13164,N_12707,N_12565);
xor U13165 (N_13165,N_12766,N_12683);
nor U13166 (N_13166,N_12697,N_12653);
xnor U13167 (N_13167,N_12516,N_12925);
and U13168 (N_13168,N_12748,N_12573);
and U13169 (N_13169,N_12840,N_12567);
xnor U13170 (N_13170,N_12759,N_12789);
xnor U13171 (N_13171,N_12732,N_12600);
nand U13172 (N_13172,N_12893,N_12633);
or U13173 (N_13173,N_12978,N_12678);
nor U13174 (N_13174,N_12690,N_12711);
nor U13175 (N_13175,N_12540,N_12984);
and U13176 (N_13176,N_12700,N_12657);
and U13177 (N_13177,N_12965,N_12829);
or U13178 (N_13178,N_12520,N_12528);
nor U13179 (N_13179,N_12726,N_12751);
and U13180 (N_13180,N_12874,N_12843);
nand U13181 (N_13181,N_12761,N_12860);
and U13182 (N_13182,N_12708,N_12576);
and U13183 (N_13183,N_12670,N_12898);
and U13184 (N_13184,N_12676,N_12525);
or U13185 (N_13185,N_12689,N_12621);
and U13186 (N_13186,N_12797,N_12831);
nand U13187 (N_13187,N_12631,N_12741);
nand U13188 (N_13188,N_12782,N_12718);
or U13189 (N_13189,N_12949,N_12547);
nor U13190 (N_13190,N_12682,N_12607);
and U13191 (N_13191,N_12602,N_12956);
or U13192 (N_13192,N_12619,N_12787);
nand U13193 (N_13193,N_12853,N_12541);
nand U13194 (N_13194,N_12672,N_12777);
nor U13195 (N_13195,N_12740,N_12539);
xnor U13196 (N_13196,N_12523,N_12975);
xor U13197 (N_13197,N_12943,N_12721);
xnor U13198 (N_13198,N_12561,N_12737);
xnor U13199 (N_13199,N_12587,N_12659);
nor U13200 (N_13200,N_12989,N_12865);
and U13201 (N_13201,N_12953,N_12595);
nor U13202 (N_13202,N_12609,N_12967);
nand U13203 (N_13203,N_12791,N_12714);
nor U13204 (N_13204,N_12786,N_12601);
or U13205 (N_13205,N_12615,N_12854);
or U13206 (N_13206,N_12852,N_12758);
xnor U13207 (N_13207,N_12750,N_12763);
or U13208 (N_13208,N_12645,N_12790);
nor U13209 (N_13209,N_12739,N_12819);
and U13210 (N_13210,N_12896,N_12920);
nand U13211 (N_13211,N_12599,N_12889);
xor U13212 (N_13212,N_12733,N_12832);
or U13213 (N_13213,N_12844,N_12918);
and U13214 (N_13214,N_12605,N_12673);
xor U13215 (N_13215,N_12642,N_12932);
and U13216 (N_13216,N_12623,N_12694);
nor U13217 (N_13217,N_12552,N_12668);
nand U13218 (N_13218,N_12674,N_12899);
nor U13219 (N_13219,N_12652,N_12579);
or U13220 (N_13220,N_12779,N_12558);
nand U13221 (N_13221,N_12669,N_12821);
nor U13222 (N_13222,N_12914,N_12909);
nor U13223 (N_13223,N_12515,N_12651);
nor U13224 (N_13224,N_12985,N_12548);
and U13225 (N_13225,N_12973,N_12583);
or U13226 (N_13226,N_12671,N_12817);
nand U13227 (N_13227,N_12537,N_12977);
or U13228 (N_13228,N_12656,N_12869);
xor U13229 (N_13229,N_12863,N_12902);
xor U13230 (N_13230,N_12912,N_12661);
xor U13231 (N_13231,N_12991,N_12959);
nand U13232 (N_13232,N_12792,N_12585);
nor U13233 (N_13233,N_12594,N_12696);
or U13234 (N_13234,N_12513,N_12719);
or U13235 (N_13235,N_12816,N_12667);
nand U13236 (N_13236,N_12915,N_12807);
xor U13237 (N_13237,N_12598,N_12643);
and U13238 (N_13238,N_12944,N_12529);
nand U13239 (N_13239,N_12862,N_12952);
xnor U13240 (N_13240,N_12913,N_12606);
or U13241 (N_13241,N_12926,N_12702);
and U13242 (N_13242,N_12812,N_12928);
nor U13243 (N_13243,N_12687,N_12506);
nor U13244 (N_13244,N_12762,N_12870);
nand U13245 (N_13245,N_12639,N_12826);
or U13246 (N_13246,N_12745,N_12981);
or U13247 (N_13247,N_12572,N_12604);
or U13248 (N_13248,N_12752,N_12772);
xor U13249 (N_13249,N_12878,N_12536);
or U13250 (N_13250,N_12680,N_12554);
nand U13251 (N_13251,N_12568,N_12719);
or U13252 (N_13252,N_12660,N_12716);
or U13253 (N_13253,N_12688,N_12758);
or U13254 (N_13254,N_12699,N_12981);
or U13255 (N_13255,N_12782,N_12970);
xnor U13256 (N_13256,N_12726,N_12667);
or U13257 (N_13257,N_12701,N_12926);
xor U13258 (N_13258,N_12628,N_12801);
nor U13259 (N_13259,N_12910,N_12696);
and U13260 (N_13260,N_12818,N_12802);
nand U13261 (N_13261,N_12521,N_12619);
or U13262 (N_13262,N_12860,N_12942);
xor U13263 (N_13263,N_12656,N_12653);
nor U13264 (N_13264,N_12557,N_12805);
nand U13265 (N_13265,N_12696,N_12852);
or U13266 (N_13266,N_12744,N_12638);
or U13267 (N_13267,N_12675,N_12618);
nor U13268 (N_13268,N_12790,N_12566);
and U13269 (N_13269,N_12842,N_12767);
nor U13270 (N_13270,N_12586,N_12532);
xnor U13271 (N_13271,N_12635,N_12849);
nor U13272 (N_13272,N_12825,N_12706);
xor U13273 (N_13273,N_12578,N_12819);
and U13274 (N_13274,N_12651,N_12672);
xnor U13275 (N_13275,N_12568,N_12901);
or U13276 (N_13276,N_12891,N_12584);
nand U13277 (N_13277,N_12539,N_12701);
nor U13278 (N_13278,N_12715,N_12548);
or U13279 (N_13279,N_12832,N_12841);
nand U13280 (N_13280,N_12993,N_12940);
nand U13281 (N_13281,N_12980,N_12555);
or U13282 (N_13282,N_12636,N_12964);
nor U13283 (N_13283,N_12618,N_12854);
xnor U13284 (N_13284,N_12664,N_12693);
nor U13285 (N_13285,N_12644,N_12686);
xnor U13286 (N_13286,N_12532,N_12968);
or U13287 (N_13287,N_12524,N_12532);
nand U13288 (N_13288,N_12818,N_12997);
nand U13289 (N_13289,N_12565,N_12737);
and U13290 (N_13290,N_12825,N_12544);
nor U13291 (N_13291,N_12543,N_12559);
nand U13292 (N_13292,N_12895,N_12886);
nand U13293 (N_13293,N_12875,N_12836);
nand U13294 (N_13294,N_12743,N_12668);
nor U13295 (N_13295,N_12883,N_12990);
nor U13296 (N_13296,N_12800,N_12956);
and U13297 (N_13297,N_12845,N_12744);
or U13298 (N_13298,N_12551,N_12825);
nand U13299 (N_13299,N_12701,N_12793);
xnor U13300 (N_13300,N_12710,N_12841);
xnor U13301 (N_13301,N_12719,N_12949);
nand U13302 (N_13302,N_12591,N_12981);
and U13303 (N_13303,N_12552,N_12777);
nor U13304 (N_13304,N_12771,N_12659);
and U13305 (N_13305,N_12656,N_12787);
and U13306 (N_13306,N_12924,N_12880);
or U13307 (N_13307,N_12974,N_12661);
xor U13308 (N_13308,N_12688,N_12713);
and U13309 (N_13309,N_12961,N_12683);
nand U13310 (N_13310,N_12665,N_12925);
nor U13311 (N_13311,N_12914,N_12916);
nor U13312 (N_13312,N_12596,N_12647);
nand U13313 (N_13313,N_12546,N_12861);
xor U13314 (N_13314,N_12886,N_12805);
xor U13315 (N_13315,N_12899,N_12767);
nand U13316 (N_13316,N_12774,N_12758);
xor U13317 (N_13317,N_12910,N_12996);
nand U13318 (N_13318,N_12513,N_12691);
xor U13319 (N_13319,N_12903,N_12837);
nand U13320 (N_13320,N_12956,N_12967);
nor U13321 (N_13321,N_12583,N_12833);
and U13322 (N_13322,N_12585,N_12944);
xor U13323 (N_13323,N_12960,N_12955);
and U13324 (N_13324,N_12519,N_12554);
nand U13325 (N_13325,N_12858,N_12831);
nor U13326 (N_13326,N_12967,N_12785);
xnor U13327 (N_13327,N_12566,N_12906);
and U13328 (N_13328,N_12969,N_12976);
nor U13329 (N_13329,N_12877,N_12907);
xor U13330 (N_13330,N_12746,N_12954);
nand U13331 (N_13331,N_12576,N_12600);
or U13332 (N_13332,N_12611,N_12786);
and U13333 (N_13333,N_12612,N_12673);
xor U13334 (N_13334,N_12624,N_12960);
xnor U13335 (N_13335,N_12985,N_12907);
or U13336 (N_13336,N_12588,N_12800);
xor U13337 (N_13337,N_12871,N_12657);
nor U13338 (N_13338,N_12667,N_12875);
and U13339 (N_13339,N_12651,N_12735);
xnor U13340 (N_13340,N_12913,N_12898);
nor U13341 (N_13341,N_12984,N_12882);
and U13342 (N_13342,N_12692,N_12714);
xnor U13343 (N_13343,N_12889,N_12948);
and U13344 (N_13344,N_12791,N_12525);
xor U13345 (N_13345,N_12730,N_12565);
nand U13346 (N_13346,N_12849,N_12605);
xnor U13347 (N_13347,N_12713,N_12630);
nand U13348 (N_13348,N_12664,N_12707);
nor U13349 (N_13349,N_12584,N_12947);
or U13350 (N_13350,N_12500,N_12952);
or U13351 (N_13351,N_12956,N_12904);
nand U13352 (N_13352,N_12800,N_12754);
xnor U13353 (N_13353,N_12664,N_12767);
nand U13354 (N_13354,N_12531,N_12697);
nand U13355 (N_13355,N_12606,N_12803);
xnor U13356 (N_13356,N_12815,N_12909);
nand U13357 (N_13357,N_12593,N_12536);
nor U13358 (N_13358,N_12878,N_12992);
and U13359 (N_13359,N_12987,N_12827);
xnor U13360 (N_13360,N_12952,N_12602);
nor U13361 (N_13361,N_12960,N_12683);
nand U13362 (N_13362,N_12764,N_12761);
or U13363 (N_13363,N_12750,N_12996);
and U13364 (N_13364,N_12951,N_12595);
xor U13365 (N_13365,N_12882,N_12692);
xnor U13366 (N_13366,N_12615,N_12909);
xnor U13367 (N_13367,N_12961,N_12794);
or U13368 (N_13368,N_12791,N_12828);
nand U13369 (N_13369,N_12876,N_12782);
nor U13370 (N_13370,N_12639,N_12796);
nor U13371 (N_13371,N_12648,N_12972);
xnor U13372 (N_13372,N_12534,N_12966);
nand U13373 (N_13373,N_12758,N_12991);
xor U13374 (N_13374,N_12572,N_12988);
or U13375 (N_13375,N_12964,N_12950);
nand U13376 (N_13376,N_12773,N_12506);
and U13377 (N_13377,N_12867,N_12780);
xor U13378 (N_13378,N_12922,N_12817);
xnor U13379 (N_13379,N_12531,N_12947);
and U13380 (N_13380,N_12640,N_12797);
nor U13381 (N_13381,N_12985,N_12954);
and U13382 (N_13382,N_12822,N_12693);
nor U13383 (N_13383,N_12551,N_12529);
and U13384 (N_13384,N_12540,N_12699);
nor U13385 (N_13385,N_12538,N_12912);
nand U13386 (N_13386,N_12859,N_12826);
nor U13387 (N_13387,N_12912,N_12871);
nand U13388 (N_13388,N_12702,N_12601);
or U13389 (N_13389,N_12683,N_12966);
xor U13390 (N_13390,N_12887,N_12581);
xnor U13391 (N_13391,N_12876,N_12873);
or U13392 (N_13392,N_12982,N_12553);
nand U13393 (N_13393,N_12975,N_12814);
and U13394 (N_13394,N_12834,N_12924);
nand U13395 (N_13395,N_12835,N_12904);
or U13396 (N_13396,N_12678,N_12554);
or U13397 (N_13397,N_12625,N_12759);
nand U13398 (N_13398,N_12533,N_12811);
or U13399 (N_13399,N_12541,N_12513);
or U13400 (N_13400,N_12900,N_12946);
or U13401 (N_13401,N_12590,N_12764);
or U13402 (N_13402,N_12765,N_12930);
xor U13403 (N_13403,N_12844,N_12817);
and U13404 (N_13404,N_12776,N_12751);
or U13405 (N_13405,N_12876,N_12845);
or U13406 (N_13406,N_12892,N_12647);
nand U13407 (N_13407,N_12534,N_12631);
nor U13408 (N_13408,N_12838,N_12667);
nand U13409 (N_13409,N_12798,N_12692);
or U13410 (N_13410,N_12814,N_12647);
nand U13411 (N_13411,N_12775,N_12796);
nor U13412 (N_13412,N_12625,N_12739);
nor U13413 (N_13413,N_12894,N_12555);
xnor U13414 (N_13414,N_12815,N_12965);
xnor U13415 (N_13415,N_12584,N_12588);
or U13416 (N_13416,N_12507,N_12645);
nand U13417 (N_13417,N_12539,N_12858);
and U13418 (N_13418,N_12667,N_12610);
xnor U13419 (N_13419,N_12514,N_12754);
nor U13420 (N_13420,N_12540,N_12723);
nand U13421 (N_13421,N_12966,N_12580);
and U13422 (N_13422,N_12982,N_12583);
and U13423 (N_13423,N_12910,N_12810);
or U13424 (N_13424,N_12802,N_12838);
xor U13425 (N_13425,N_12814,N_12804);
and U13426 (N_13426,N_12675,N_12782);
or U13427 (N_13427,N_12766,N_12676);
and U13428 (N_13428,N_12690,N_12955);
nor U13429 (N_13429,N_12634,N_12793);
nand U13430 (N_13430,N_12598,N_12641);
xnor U13431 (N_13431,N_12519,N_12528);
nor U13432 (N_13432,N_12529,N_12856);
xnor U13433 (N_13433,N_12838,N_12509);
or U13434 (N_13434,N_12934,N_12929);
and U13435 (N_13435,N_12892,N_12763);
nor U13436 (N_13436,N_12753,N_12702);
or U13437 (N_13437,N_12662,N_12550);
nand U13438 (N_13438,N_12702,N_12783);
nor U13439 (N_13439,N_12994,N_12650);
nand U13440 (N_13440,N_12742,N_12698);
nor U13441 (N_13441,N_12685,N_12788);
and U13442 (N_13442,N_12988,N_12928);
or U13443 (N_13443,N_12599,N_12715);
nand U13444 (N_13444,N_12560,N_12921);
nand U13445 (N_13445,N_12671,N_12871);
xnor U13446 (N_13446,N_12637,N_12556);
or U13447 (N_13447,N_12701,N_12608);
or U13448 (N_13448,N_12843,N_12691);
or U13449 (N_13449,N_12950,N_12730);
and U13450 (N_13450,N_12646,N_12821);
or U13451 (N_13451,N_12913,N_12691);
xor U13452 (N_13452,N_12531,N_12781);
xor U13453 (N_13453,N_12554,N_12849);
and U13454 (N_13454,N_12993,N_12805);
xor U13455 (N_13455,N_12835,N_12833);
nand U13456 (N_13456,N_12841,N_12765);
or U13457 (N_13457,N_12877,N_12995);
xor U13458 (N_13458,N_12665,N_12577);
or U13459 (N_13459,N_12573,N_12642);
or U13460 (N_13460,N_12508,N_12827);
nor U13461 (N_13461,N_12901,N_12757);
nand U13462 (N_13462,N_12791,N_12767);
nor U13463 (N_13463,N_12668,N_12661);
and U13464 (N_13464,N_12689,N_12832);
xnor U13465 (N_13465,N_12898,N_12999);
and U13466 (N_13466,N_12919,N_12941);
nor U13467 (N_13467,N_12814,N_12883);
or U13468 (N_13468,N_12954,N_12775);
nor U13469 (N_13469,N_12912,N_12614);
and U13470 (N_13470,N_12705,N_12747);
and U13471 (N_13471,N_12856,N_12813);
and U13472 (N_13472,N_12591,N_12617);
xor U13473 (N_13473,N_12711,N_12858);
xnor U13474 (N_13474,N_12545,N_12786);
nand U13475 (N_13475,N_12606,N_12726);
or U13476 (N_13476,N_12908,N_12994);
and U13477 (N_13477,N_12674,N_12838);
and U13478 (N_13478,N_12614,N_12779);
xnor U13479 (N_13479,N_12649,N_12565);
and U13480 (N_13480,N_12811,N_12820);
and U13481 (N_13481,N_12994,N_12806);
nand U13482 (N_13482,N_12988,N_12599);
or U13483 (N_13483,N_12627,N_12985);
or U13484 (N_13484,N_12955,N_12883);
nor U13485 (N_13485,N_12771,N_12601);
and U13486 (N_13486,N_12513,N_12688);
nor U13487 (N_13487,N_12924,N_12955);
and U13488 (N_13488,N_12678,N_12526);
nor U13489 (N_13489,N_12531,N_12937);
nor U13490 (N_13490,N_12643,N_12691);
nand U13491 (N_13491,N_12688,N_12783);
nor U13492 (N_13492,N_12762,N_12879);
xor U13493 (N_13493,N_12591,N_12794);
nor U13494 (N_13494,N_12997,N_12940);
or U13495 (N_13495,N_12763,N_12826);
and U13496 (N_13496,N_12681,N_12950);
nand U13497 (N_13497,N_12794,N_12786);
nand U13498 (N_13498,N_12582,N_12838);
and U13499 (N_13499,N_12742,N_12633);
or U13500 (N_13500,N_13204,N_13160);
nor U13501 (N_13501,N_13411,N_13255);
or U13502 (N_13502,N_13226,N_13124);
nor U13503 (N_13503,N_13444,N_13278);
or U13504 (N_13504,N_13198,N_13326);
nor U13505 (N_13505,N_13053,N_13484);
and U13506 (N_13506,N_13289,N_13424);
xnor U13507 (N_13507,N_13400,N_13183);
or U13508 (N_13508,N_13246,N_13005);
nor U13509 (N_13509,N_13401,N_13364);
xor U13510 (N_13510,N_13426,N_13138);
xnor U13511 (N_13511,N_13331,N_13024);
nand U13512 (N_13512,N_13154,N_13354);
nand U13513 (N_13513,N_13136,N_13311);
and U13514 (N_13514,N_13271,N_13279);
and U13515 (N_13515,N_13052,N_13387);
or U13516 (N_13516,N_13223,N_13001);
nand U13517 (N_13517,N_13039,N_13429);
nand U13518 (N_13518,N_13458,N_13245);
or U13519 (N_13519,N_13383,N_13064);
and U13520 (N_13520,N_13152,N_13362);
xnor U13521 (N_13521,N_13067,N_13352);
nor U13522 (N_13522,N_13098,N_13149);
xnor U13523 (N_13523,N_13155,N_13211);
xnor U13524 (N_13524,N_13475,N_13378);
nor U13525 (N_13525,N_13442,N_13283);
nor U13526 (N_13526,N_13402,N_13302);
or U13527 (N_13527,N_13242,N_13269);
or U13528 (N_13528,N_13170,N_13186);
xnor U13529 (N_13529,N_13294,N_13292);
nor U13530 (N_13530,N_13035,N_13079);
and U13531 (N_13531,N_13057,N_13435);
or U13532 (N_13532,N_13405,N_13389);
nor U13533 (N_13533,N_13494,N_13384);
nor U13534 (N_13534,N_13277,N_13129);
xnor U13535 (N_13535,N_13158,N_13325);
nor U13536 (N_13536,N_13000,N_13410);
or U13537 (N_13537,N_13290,N_13011);
nor U13538 (N_13538,N_13036,N_13119);
nor U13539 (N_13539,N_13252,N_13372);
nand U13540 (N_13540,N_13111,N_13376);
nor U13541 (N_13541,N_13371,N_13247);
or U13542 (N_13542,N_13355,N_13254);
nor U13543 (N_13543,N_13237,N_13340);
or U13544 (N_13544,N_13034,N_13218);
xnor U13545 (N_13545,N_13100,N_13133);
nor U13546 (N_13546,N_13356,N_13055);
xor U13547 (N_13547,N_13492,N_13162);
nand U13548 (N_13548,N_13105,N_13134);
nor U13549 (N_13549,N_13425,N_13438);
nor U13550 (N_13550,N_13126,N_13346);
and U13551 (N_13551,N_13249,N_13320);
and U13552 (N_13552,N_13224,N_13443);
nand U13553 (N_13553,N_13392,N_13151);
nor U13554 (N_13554,N_13409,N_13153);
and U13555 (N_13555,N_13256,N_13343);
nor U13556 (N_13556,N_13301,N_13214);
nand U13557 (N_13557,N_13122,N_13359);
or U13558 (N_13558,N_13447,N_13228);
nand U13559 (N_13559,N_13436,N_13069);
or U13560 (N_13560,N_13396,N_13422);
nand U13561 (N_13561,N_13399,N_13025);
xor U13562 (N_13562,N_13212,N_13167);
nor U13563 (N_13563,N_13490,N_13293);
and U13564 (N_13564,N_13415,N_13201);
or U13565 (N_13565,N_13106,N_13262);
xor U13566 (N_13566,N_13266,N_13303);
nor U13567 (N_13567,N_13465,N_13179);
nand U13568 (N_13568,N_13070,N_13207);
xnor U13569 (N_13569,N_13274,N_13470);
and U13570 (N_13570,N_13107,N_13093);
xor U13571 (N_13571,N_13434,N_13299);
nand U13572 (N_13572,N_13339,N_13193);
nor U13573 (N_13573,N_13091,N_13413);
or U13574 (N_13574,N_13412,N_13141);
and U13575 (N_13575,N_13419,N_13157);
nand U13576 (N_13576,N_13042,N_13403);
xnor U13577 (N_13577,N_13408,N_13188);
nand U13578 (N_13578,N_13463,N_13008);
xnor U13579 (N_13579,N_13081,N_13472);
nand U13580 (N_13580,N_13088,N_13427);
nor U13581 (N_13581,N_13022,N_13075);
nand U13582 (N_13582,N_13385,N_13431);
nor U13583 (N_13583,N_13197,N_13227);
nor U13584 (N_13584,N_13307,N_13488);
nor U13585 (N_13585,N_13464,N_13496);
xor U13586 (N_13586,N_13441,N_13027);
nand U13587 (N_13587,N_13112,N_13280);
xor U13588 (N_13588,N_13043,N_13267);
and U13589 (N_13589,N_13456,N_13369);
nand U13590 (N_13590,N_13483,N_13082);
nor U13591 (N_13591,N_13108,N_13049);
nand U13592 (N_13592,N_13144,N_13391);
xnor U13593 (N_13593,N_13377,N_13131);
and U13594 (N_13594,N_13213,N_13086);
nand U13595 (N_13595,N_13234,N_13322);
nand U13596 (N_13596,N_13020,N_13048);
and U13597 (N_13597,N_13169,N_13499);
nor U13598 (N_13598,N_13261,N_13316);
or U13599 (N_13599,N_13338,N_13397);
and U13600 (N_13600,N_13139,N_13386);
nand U13601 (N_13601,N_13121,N_13099);
or U13602 (N_13602,N_13459,N_13478);
nand U13603 (N_13603,N_13404,N_13103);
xor U13604 (N_13604,N_13077,N_13466);
and U13605 (N_13605,N_13469,N_13394);
nand U13606 (N_13606,N_13231,N_13063);
nand U13607 (N_13607,N_13321,N_13215);
nand U13608 (N_13608,N_13379,N_13018);
nor U13609 (N_13609,N_13440,N_13040);
nor U13610 (N_13610,N_13332,N_13461);
nand U13611 (N_13611,N_13272,N_13172);
nor U13612 (N_13612,N_13113,N_13491);
and U13613 (N_13613,N_13178,N_13327);
nor U13614 (N_13614,N_13002,N_13334);
nand U13615 (N_13615,N_13467,N_13328);
or U13616 (N_13616,N_13350,N_13295);
nand U13617 (N_13617,N_13284,N_13176);
or U13618 (N_13618,N_13497,N_13480);
nor U13619 (N_13619,N_13166,N_13263);
xnor U13620 (N_13620,N_13357,N_13208);
or U13621 (N_13621,N_13360,N_13014);
or U13622 (N_13622,N_13473,N_13140);
nor U13623 (N_13623,N_13406,N_13095);
or U13624 (N_13624,N_13446,N_13184);
and U13625 (N_13625,N_13233,N_13033);
or U13626 (N_13626,N_13324,N_13353);
and U13627 (N_13627,N_13418,N_13071);
nor U13628 (N_13628,N_13310,N_13417);
nor U13629 (N_13629,N_13109,N_13021);
or U13630 (N_13630,N_13090,N_13205);
nand U13631 (N_13631,N_13457,N_13333);
nand U13632 (N_13632,N_13433,N_13248);
xor U13633 (N_13633,N_13031,N_13056);
nand U13634 (N_13634,N_13460,N_13217);
xnor U13635 (N_13635,N_13335,N_13045);
xnor U13636 (N_13636,N_13341,N_13060);
and U13637 (N_13637,N_13381,N_13150);
or U13638 (N_13638,N_13250,N_13072);
nand U13639 (N_13639,N_13029,N_13462);
xnor U13640 (N_13640,N_13146,N_13388);
xnor U13641 (N_13641,N_13319,N_13368);
or U13642 (N_13642,N_13486,N_13199);
nand U13643 (N_13643,N_13323,N_13062);
nor U13644 (N_13644,N_13448,N_13165);
xnor U13645 (N_13645,N_13287,N_13312);
nor U13646 (N_13646,N_13159,N_13414);
nor U13647 (N_13647,N_13454,N_13143);
nor U13648 (N_13648,N_13078,N_13087);
and U13649 (N_13649,N_13317,N_13315);
or U13650 (N_13650,N_13192,N_13210);
xor U13651 (N_13651,N_13244,N_13161);
xnor U13652 (N_13652,N_13330,N_13276);
xor U13653 (N_13653,N_13230,N_13085);
nor U13654 (N_13654,N_13127,N_13206);
xor U13655 (N_13655,N_13373,N_13265);
nor U13656 (N_13656,N_13345,N_13061);
or U13657 (N_13657,N_13222,N_13285);
nor U13658 (N_13658,N_13185,N_13375);
nand U13659 (N_13659,N_13164,N_13498);
nor U13660 (N_13660,N_13175,N_13296);
and U13661 (N_13661,N_13259,N_13065);
or U13662 (N_13662,N_13382,N_13037);
nand U13663 (N_13663,N_13370,N_13398);
and U13664 (N_13664,N_13125,N_13195);
nand U13665 (N_13665,N_13174,N_13239);
or U13666 (N_13666,N_13041,N_13474);
or U13667 (N_13667,N_13297,N_13110);
nand U13668 (N_13668,N_13051,N_13300);
xor U13669 (N_13669,N_13380,N_13349);
nor U13670 (N_13670,N_13337,N_13291);
xnor U13671 (N_13671,N_13135,N_13187);
or U13672 (N_13672,N_13275,N_13481);
and U13673 (N_13673,N_13445,N_13468);
nor U13674 (N_13674,N_13240,N_13485);
nor U13675 (N_13675,N_13342,N_13200);
nand U13676 (N_13676,N_13102,N_13050);
nand U13677 (N_13677,N_13257,N_13089);
and U13678 (N_13678,N_13073,N_13471);
and U13679 (N_13679,N_13015,N_13238);
and U13680 (N_13680,N_13083,N_13028);
nand U13681 (N_13681,N_13298,N_13305);
xnor U13682 (N_13682,N_13117,N_13004);
nand U13683 (N_13683,N_13329,N_13009);
nand U13684 (N_13684,N_13288,N_13148);
nand U13685 (N_13685,N_13006,N_13455);
and U13686 (N_13686,N_13177,N_13452);
xor U13687 (N_13687,N_13147,N_13236);
or U13688 (N_13688,N_13016,N_13286);
nand U13689 (N_13689,N_13066,N_13428);
nor U13690 (N_13690,N_13281,N_13420);
or U13691 (N_13691,N_13010,N_13495);
xnor U13692 (N_13692,N_13358,N_13104);
xor U13693 (N_13693,N_13390,N_13476);
nand U13694 (N_13694,N_13351,N_13074);
xor U13695 (N_13695,N_13437,N_13229);
nand U13696 (N_13696,N_13023,N_13258);
xnor U13697 (N_13697,N_13130,N_13235);
or U13698 (N_13698,N_13080,N_13407);
nor U13699 (N_13699,N_13260,N_13173);
nand U13700 (N_13700,N_13116,N_13309);
nor U13701 (N_13701,N_13493,N_13479);
nor U13702 (N_13702,N_13251,N_13190);
xnor U13703 (N_13703,N_13209,N_13374);
or U13704 (N_13704,N_13363,N_13221);
xnor U13705 (N_13705,N_13038,N_13365);
or U13706 (N_13706,N_13423,N_13304);
or U13707 (N_13707,N_13241,N_13189);
xnor U13708 (N_13708,N_13076,N_13450);
nor U13709 (N_13709,N_13449,N_13168);
or U13710 (N_13710,N_13046,N_13007);
and U13711 (N_13711,N_13084,N_13344);
xor U13712 (N_13712,N_13253,N_13115);
and U13713 (N_13713,N_13306,N_13453);
nand U13714 (N_13714,N_13273,N_13094);
and U13715 (N_13715,N_13120,N_13264);
and U13716 (N_13716,N_13058,N_13044);
and U13717 (N_13717,N_13318,N_13012);
or U13718 (N_13718,N_13219,N_13118);
or U13719 (N_13719,N_13092,N_13156);
or U13720 (N_13720,N_13132,N_13439);
xor U13721 (N_13721,N_13482,N_13416);
nand U13722 (N_13722,N_13477,N_13003);
nor U13723 (N_13723,N_13019,N_13243);
and U13724 (N_13724,N_13196,N_13270);
nand U13725 (N_13725,N_13313,N_13203);
xnor U13726 (N_13726,N_13220,N_13393);
nand U13727 (N_13727,N_13101,N_13421);
or U13728 (N_13728,N_13308,N_13145);
nand U13729 (N_13729,N_13128,N_13097);
nand U13730 (N_13730,N_13026,N_13171);
nand U13731 (N_13731,N_13432,N_13347);
nand U13732 (N_13732,N_13142,N_13366);
nor U13733 (N_13733,N_13030,N_13367);
xnor U13734 (N_13734,N_13032,N_13282);
or U13735 (N_13735,N_13194,N_13202);
nand U13736 (N_13736,N_13180,N_13430);
and U13737 (N_13737,N_13013,N_13054);
nand U13738 (N_13738,N_13163,N_13114);
or U13739 (N_13739,N_13348,N_13268);
xor U13740 (N_13740,N_13182,N_13068);
or U13741 (N_13741,N_13059,N_13181);
xor U13742 (N_13742,N_13216,N_13395);
and U13743 (N_13743,N_13047,N_13336);
xnor U13744 (N_13744,N_13017,N_13191);
and U13745 (N_13745,N_13487,N_13314);
nand U13746 (N_13746,N_13123,N_13096);
xor U13747 (N_13747,N_13225,N_13137);
xnor U13748 (N_13748,N_13361,N_13451);
nor U13749 (N_13749,N_13489,N_13232);
and U13750 (N_13750,N_13301,N_13130);
and U13751 (N_13751,N_13248,N_13396);
or U13752 (N_13752,N_13159,N_13245);
nand U13753 (N_13753,N_13473,N_13411);
nor U13754 (N_13754,N_13166,N_13347);
nor U13755 (N_13755,N_13369,N_13054);
xnor U13756 (N_13756,N_13484,N_13049);
xnor U13757 (N_13757,N_13210,N_13209);
and U13758 (N_13758,N_13421,N_13043);
xnor U13759 (N_13759,N_13455,N_13342);
nand U13760 (N_13760,N_13238,N_13264);
nor U13761 (N_13761,N_13027,N_13159);
xor U13762 (N_13762,N_13403,N_13136);
xnor U13763 (N_13763,N_13165,N_13411);
nand U13764 (N_13764,N_13421,N_13390);
xor U13765 (N_13765,N_13299,N_13445);
or U13766 (N_13766,N_13303,N_13158);
xor U13767 (N_13767,N_13357,N_13447);
nor U13768 (N_13768,N_13290,N_13065);
nand U13769 (N_13769,N_13422,N_13052);
xnor U13770 (N_13770,N_13401,N_13306);
and U13771 (N_13771,N_13280,N_13091);
nor U13772 (N_13772,N_13462,N_13128);
or U13773 (N_13773,N_13484,N_13163);
nor U13774 (N_13774,N_13163,N_13357);
xnor U13775 (N_13775,N_13163,N_13383);
xor U13776 (N_13776,N_13263,N_13077);
nand U13777 (N_13777,N_13411,N_13003);
nor U13778 (N_13778,N_13080,N_13010);
and U13779 (N_13779,N_13284,N_13410);
nand U13780 (N_13780,N_13405,N_13339);
and U13781 (N_13781,N_13305,N_13409);
xnor U13782 (N_13782,N_13290,N_13028);
nor U13783 (N_13783,N_13266,N_13006);
nand U13784 (N_13784,N_13424,N_13113);
xnor U13785 (N_13785,N_13236,N_13398);
nand U13786 (N_13786,N_13175,N_13325);
and U13787 (N_13787,N_13360,N_13079);
nor U13788 (N_13788,N_13385,N_13042);
or U13789 (N_13789,N_13068,N_13028);
or U13790 (N_13790,N_13082,N_13187);
nor U13791 (N_13791,N_13354,N_13494);
xnor U13792 (N_13792,N_13315,N_13349);
nand U13793 (N_13793,N_13156,N_13206);
xor U13794 (N_13794,N_13128,N_13182);
and U13795 (N_13795,N_13274,N_13040);
nand U13796 (N_13796,N_13451,N_13229);
and U13797 (N_13797,N_13309,N_13105);
nor U13798 (N_13798,N_13473,N_13118);
nand U13799 (N_13799,N_13195,N_13026);
nand U13800 (N_13800,N_13005,N_13081);
nand U13801 (N_13801,N_13127,N_13003);
or U13802 (N_13802,N_13404,N_13475);
and U13803 (N_13803,N_13393,N_13165);
nand U13804 (N_13804,N_13170,N_13178);
nand U13805 (N_13805,N_13481,N_13398);
and U13806 (N_13806,N_13319,N_13104);
or U13807 (N_13807,N_13039,N_13414);
nor U13808 (N_13808,N_13390,N_13284);
nand U13809 (N_13809,N_13477,N_13468);
nand U13810 (N_13810,N_13248,N_13497);
and U13811 (N_13811,N_13127,N_13122);
and U13812 (N_13812,N_13203,N_13493);
or U13813 (N_13813,N_13149,N_13272);
xor U13814 (N_13814,N_13060,N_13203);
or U13815 (N_13815,N_13215,N_13104);
nand U13816 (N_13816,N_13069,N_13219);
xnor U13817 (N_13817,N_13471,N_13293);
xor U13818 (N_13818,N_13394,N_13384);
nand U13819 (N_13819,N_13450,N_13400);
xnor U13820 (N_13820,N_13085,N_13389);
and U13821 (N_13821,N_13155,N_13149);
nor U13822 (N_13822,N_13247,N_13478);
or U13823 (N_13823,N_13403,N_13008);
nor U13824 (N_13824,N_13032,N_13395);
nand U13825 (N_13825,N_13017,N_13055);
or U13826 (N_13826,N_13107,N_13018);
and U13827 (N_13827,N_13220,N_13323);
or U13828 (N_13828,N_13403,N_13106);
nor U13829 (N_13829,N_13474,N_13195);
nor U13830 (N_13830,N_13330,N_13454);
xnor U13831 (N_13831,N_13145,N_13269);
nand U13832 (N_13832,N_13185,N_13105);
or U13833 (N_13833,N_13355,N_13442);
and U13834 (N_13834,N_13295,N_13229);
nor U13835 (N_13835,N_13037,N_13028);
nand U13836 (N_13836,N_13071,N_13206);
nor U13837 (N_13837,N_13487,N_13055);
or U13838 (N_13838,N_13044,N_13056);
nor U13839 (N_13839,N_13321,N_13045);
and U13840 (N_13840,N_13266,N_13434);
nor U13841 (N_13841,N_13461,N_13413);
nor U13842 (N_13842,N_13465,N_13126);
or U13843 (N_13843,N_13405,N_13007);
nor U13844 (N_13844,N_13291,N_13466);
nand U13845 (N_13845,N_13352,N_13092);
or U13846 (N_13846,N_13107,N_13039);
or U13847 (N_13847,N_13022,N_13004);
or U13848 (N_13848,N_13495,N_13377);
and U13849 (N_13849,N_13149,N_13403);
nor U13850 (N_13850,N_13373,N_13273);
nand U13851 (N_13851,N_13027,N_13352);
or U13852 (N_13852,N_13399,N_13135);
xnor U13853 (N_13853,N_13384,N_13029);
nor U13854 (N_13854,N_13175,N_13499);
nor U13855 (N_13855,N_13103,N_13193);
nand U13856 (N_13856,N_13209,N_13078);
nor U13857 (N_13857,N_13052,N_13386);
and U13858 (N_13858,N_13006,N_13139);
nor U13859 (N_13859,N_13119,N_13228);
nand U13860 (N_13860,N_13207,N_13076);
nor U13861 (N_13861,N_13398,N_13102);
nor U13862 (N_13862,N_13295,N_13274);
xnor U13863 (N_13863,N_13465,N_13323);
and U13864 (N_13864,N_13119,N_13165);
and U13865 (N_13865,N_13277,N_13463);
xnor U13866 (N_13866,N_13313,N_13043);
nor U13867 (N_13867,N_13202,N_13097);
nor U13868 (N_13868,N_13126,N_13317);
or U13869 (N_13869,N_13110,N_13404);
and U13870 (N_13870,N_13170,N_13474);
and U13871 (N_13871,N_13212,N_13344);
xor U13872 (N_13872,N_13368,N_13419);
and U13873 (N_13873,N_13265,N_13089);
xor U13874 (N_13874,N_13270,N_13314);
nand U13875 (N_13875,N_13375,N_13031);
nand U13876 (N_13876,N_13485,N_13057);
xor U13877 (N_13877,N_13451,N_13334);
nor U13878 (N_13878,N_13478,N_13260);
and U13879 (N_13879,N_13388,N_13108);
and U13880 (N_13880,N_13189,N_13462);
nor U13881 (N_13881,N_13458,N_13255);
and U13882 (N_13882,N_13384,N_13445);
and U13883 (N_13883,N_13146,N_13362);
nor U13884 (N_13884,N_13446,N_13080);
or U13885 (N_13885,N_13279,N_13289);
xor U13886 (N_13886,N_13423,N_13290);
nor U13887 (N_13887,N_13101,N_13145);
or U13888 (N_13888,N_13274,N_13276);
nand U13889 (N_13889,N_13435,N_13095);
and U13890 (N_13890,N_13437,N_13119);
or U13891 (N_13891,N_13068,N_13047);
nor U13892 (N_13892,N_13268,N_13003);
or U13893 (N_13893,N_13328,N_13464);
nand U13894 (N_13894,N_13028,N_13259);
nor U13895 (N_13895,N_13259,N_13390);
or U13896 (N_13896,N_13074,N_13111);
or U13897 (N_13897,N_13152,N_13342);
nand U13898 (N_13898,N_13375,N_13405);
or U13899 (N_13899,N_13369,N_13106);
xor U13900 (N_13900,N_13247,N_13128);
nand U13901 (N_13901,N_13237,N_13481);
nor U13902 (N_13902,N_13416,N_13262);
xor U13903 (N_13903,N_13372,N_13480);
and U13904 (N_13904,N_13105,N_13117);
xor U13905 (N_13905,N_13205,N_13497);
and U13906 (N_13906,N_13054,N_13360);
xnor U13907 (N_13907,N_13348,N_13301);
nand U13908 (N_13908,N_13235,N_13465);
or U13909 (N_13909,N_13412,N_13321);
xnor U13910 (N_13910,N_13450,N_13439);
nor U13911 (N_13911,N_13492,N_13064);
xor U13912 (N_13912,N_13109,N_13206);
nand U13913 (N_13913,N_13206,N_13128);
nand U13914 (N_13914,N_13106,N_13376);
and U13915 (N_13915,N_13284,N_13159);
or U13916 (N_13916,N_13466,N_13118);
xor U13917 (N_13917,N_13003,N_13181);
nand U13918 (N_13918,N_13304,N_13405);
and U13919 (N_13919,N_13021,N_13173);
xor U13920 (N_13920,N_13325,N_13454);
xor U13921 (N_13921,N_13426,N_13302);
nor U13922 (N_13922,N_13079,N_13325);
nand U13923 (N_13923,N_13046,N_13364);
or U13924 (N_13924,N_13049,N_13497);
nor U13925 (N_13925,N_13417,N_13223);
nand U13926 (N_13926,N_13450,N_13443);
xor U13927 (N_13927,N_13410,N_13170);
nand U13928 (N_13928,N_13038,N_13260);
nor U13929 (N_13929,N_13064,N_13052);
and U13930 (N_13930,N_13055,N_13193);
and U13931 (N_13931,N_13427,N_13197);
nor U13932 (N_13932,N_13470,N_13204);
xnor U13933 (N_13933,N_13019,N_13460);
nor U13934 (N_13934,N_13008,N_13110);
and U13935 (N_13935,N_13330,N_13352);
nand U13936 (N_13936,N_13236,N_13187);
xnor U13937 (N_13937,N_13011,N_13159);
or U13938 (N_13938,N_13032,N_13499);
nor U13939 (N_13939,N_13150,N_13047);
xor U13940 (N_13940,N_13240,N_13121);
and U13941 (N_13941,N_13046,N_13035);
or U13942 (N_13942,N_13356,N_13319);
nand U13943 (N_13943,N_13474,N_13409);
nor U13944 (N_13944,N_13421,N_13307);
or U13945 (N_13945,N_13068,N_13364);
and U13946 (N_13946,N_13108,N_13217);
xor U13947 (N_13947,N_13207,N_13159);
nand U13948 (N_13948,N_13483,N_13221);
nand U13949 (N_13949,N_13095,N_13139);
nor U13950 (N_13950,N_13109,N_13210);
nand U13951 (N_13951,N_13156,N_13412);
nand U13952 (N_13952,N_13369,N_13278);
and U13953 (N_13953,N_13030,N_13497);
nor U13954 (N_13954,N_13170,N_13369);
or U13955 (N_13955,N_13199,N_13192);
and U13956 (N_13956,N_13215,N_13006);
and U13957 (N_13957,N_13233,N_13026);
xnor U13958 (N_13958,N_13365,N_13251);
or U13959 (N_13959,N_13248,N_13394);
and U13960 (N_13960,N_13281,N_13271);
and U13961 (N_13961,N_13336,N_13142);
nor U13962 (N_13962,N_13351,N_13464);
or U13963 (N_13963,N_13383,N_13272);
and U13964 (N_13964,N_13209,N_13202);
nand U13965 (N_13965,N_13360,N_13332);
nand U13966 (N_13966,N_13410,N_13344);
nand U13967 (N_13967,N_13043,N_13094);
nand U13968 (N_13968,N_13057,N_13208);
nor U13969 (N_13969,N_13033,N_13087);
xnor U13970 (N_13970,N_13304,N_13302);
nor U13971 (N_13971,N_13331,N_13334);
nor U13972 (N_13972,N_13320,N_13099);
and U13973 (N_13973,N_13249,N_13219);
nand U13974 (N_13974,N_13118,N_13313);
and U13975 (N_13975,N_13154,N_13227);
nor U13976 (N_13976,N_13234,N_13443);
nand U13977 (N_13977,N_13242,N_13143);
nor U13978 (N_13978,N_13470,N_13466);
nand U13979 (N_13979,N_13454,N_13455);
nand U13980 (N_13980,N_13391,N_13186);
nor U13981 (N_13981,N_13321,N_13094);
xnor U13982 (N_13982,N_13238,N_13379);
nor U13983 (N_13983,N_13131,N_13420);
or U13984 (N_13984,N_13299,N_13458);
nor U13985 (N_13985,N_13270,N_13408);
xor U13986 (N_13986,N_13161,N_13150);
and U13987 (N_13987,N_13475,N_13074);
nor U13988 (N_13988,N_13181,N_13079);
xnor U13989 (N_13989,N_13351,N_13148);
nand U13990 (N_13990,N_13345,N_13383);
nand U13991 (N_13991,N_13010,N_13217);
nor U13992 (N_13992,N_13072,N_13454);
and U13993 (N_13993,N_13311,N_13046);
and U13994 (N_13994,N_13219,N_13002);
nand U13995 (N_13995,N_13266,N_13180);
nor U13996 (N_13996,N_13257,N_13455);
xor U13997 (N_13997,N_13442,N_13153);
and U13998 (N_13998,N_13488,N_13460);
nor U13999 (N_13999,N_13334,N_13273);
nor U14000 (N_14000,N_13698,N_13640);
and U14001 (N_14001,N_13511,N_13803);
xnor U14002 (N_14002,N_13593,N_13658);
nor U14003 (N_14003,N_13629,N_13934);
or U14004 (N_14004,N_13523,N_13648);
or U14005 (N_14005,N_13829,N_13951);
and U14006 (N_14006,N_13790,N_13977);
or U14007 (N_14007,N_13631,N_13872);
or U14008 (N_14008,N_13873,N_13999);
xnor U14009 (N_14009,N_13541,N_13616);
nand U14010 (N_14010,N_13695,N_13991);
xnor U14011 (N_14011,N_13861,N_13653);
nor U14012 (N_14012,N_13601,N_13634);
nor U14013 (N_14013,N_13887,N_13516);
and U14014 (N_14014,N_13835,N_13947);
nor U14015 (N_14015,N_13569,N_13850);
or U14016 (N_14016,N_13591,N_13785);
and U14017 (N_14017,N_13617,N_13903);
xnor U14018 (N_14018,N_13997,N_13874);
or U14019 (N_14019,N_13500,N_13960);
nand U14020 (N_14020,N_13556,N_13981);
nor U14021 (N_14021,N_13988,N_13729);
nor U14022 (N_14022,N_13654,N_13526);
nor U14023 (N_14023,N_13712,N_13703);
xor U14024 (N_14024,N_13986,N_13843);
xor U14025 (N_14025,N_13832,N_13839);
and U14026 (N_14026,N_13989,N_13805);
and U14027 (N_14027,N_13700,N_13678);
xor U14028 (N_14028,N_13708,N_13920);
nor U14029 (N_14029,N_13932,N_13704);
or U14030 (N_14030,N_13975,N_13530);
and U14031 (N_14031,N_13775,N_13661);
xnor U14032 (N_14032,N_13950,N_13618);
nand U14033 (N_14033,N_13944,N_13595);
nor U14034 (N_14034,N_13600,N_13558);
or U14035 (N_14035,N_13713,N_13881);
nor U14036 (N_14036,N_13817,N_13980);
and U14037 (N_14037,N_13707,N_13894);
or U14038 (N_14038,N_13779,N_13875);
nand U14039 (N_14039,N_13592,N_13889);
xnor U14040 (N_14040,N_13580,N_13773);
xnor U14041 (N_14041,N_13705,N_13974);
nor U14042 (N_14042,N_13992,N_13725);
and U14043 (N_14043,N_13590,N_13723);
nand U14044 (N_14044,N_13660,N_13597);
nand U14045 (N_14045,N_13701,N_13818);
xor U14046 (N_14046,N_13858,N_13761);
and U14047 (N_14047,N_13519,N_13689);
and U14048 (N_14048,N_13985,N_13630);
nor U14049 (N_14049,N_13942,N_13533);
nor U14050 (N_14050,N_13971,N_13706);
nand U14051 (N_14051,N_13902,N_13876);
or U14052 (N_14052,N_13594,N_13559);
nand U14053 (N_14053,N_13691,N_13882);
or U14054 (N_14054,N_13938,N_13751);
or U14055 (N_14055,N_13690,N_13928);
nor U14056 (N_14056,N_13615,N_13565);
nor U14057 (N_14057,N_13510,N_13680);
nand U14058 (N_14058,N_13633,N_13528);
nand U14059 (N_14059,N_13984,N_13681);
and U14060 (N_14060,N_13604,N_13531);
nor U14061 (N_14061,N_13507,N_13748);
nor U14062 (N_14062,N_13863,N_13855);
or U14063 (N_14063,N_13926,N_13912);
xor U14064 (N_14064,N_13682,N_13943);
nor U14065 (N_14065,N_13906,N_13793);
xor U14066 (N_14066,N_13904,N_13983);
xnor U14067 (N_14067,N_13513,N_13965);
nor U14068 (N_14068,N_13849,N_13717);
or U14069 (N_14069,N_13537,N_13599);
xor U14070 (N_14070,N_13791,N_13727);
xor U14071 (N_14071,N_13968,N_13796);
nand U14072 (N_14072,N_13508,N_13588);
nand U14073 (N_14073,N_13792,N_13525);
xor U14074 (N_14074,N_13870,N_13871);
nand U14075 (N_14075,N_13637,N_13766);
and U14076 (N_14076,N_13841,N_13685);
or U14077 (N_14077,N_13645,N_13834);
nor U14078 (N_14078,N_13758,N_13854);
nor U14079 (N_14079,N_13621,N_13784);
nand U14080 (N_14080,N_13866,N_13990);
xor U14081 (N_14081,N_13774,N_13995);
nand U14082 (N_14082,N_13750,N_13955);
and U14083 (N_14083,N_13860,N_13816);
or U14084 (N_14084,N_13852,N_13612);
nor U14085 (N_14085,N_13998,N_13524);
nor U14086 (N_14086,N_13715,N_13551);
or U14087 (N_14087,N_13540,N_13908);
nand U14088 (N_14088,N_13949,N_13940);
nor U14089 (N_14089,N_13552,N_13976);
and U14090 (N_14090,N_13546,N_13676);
and U14091 (N_14091,N_13845,N_13584);
xor U14092 (N_14092,N_13710,N_13824);
or U14093 (N_14093,N_13574,N_13665);
or U14094 (N_14094,N_13857,N_13963);
nor U14095 (N_14095,N_13564,N_13547);
and U14096 (N_14096,N_13570,N_13898);
nand U14097 (N_14097,N_13730,N_13573);
xor U14098 (N_14098,N_13699,N_13804);
nor U14099 (N_14099,N_13840,N_13820);
nand U14100 (N_14100,N_13673,N_13786);
nand U14101 (N_14101,N_13776,N_13884);
nor U14102 (N_14102,N_13671,N_13716);
nand U14103 (N_14103,N_13522,N_13821);
xor U14104 (N_14104,N_13709,N_13521);
xnor U14105 (N_14105,N_13783,N_13607);
nor U14106 (N_14106,N_13994,N_13736);
nand U14107 (N_14107,N_13737,N_13862);
nand U14108 (N_14108,N_13627,N_13649);
or U14109 (N_14109,N_13668,N_13836);
or U14110 (N_14110,N_13927,N_13954);
or U14111 (N_14111,N_13602,N_13911);
nor U14112 (N_14112,N_13828,N_13534);
and U14113 (N_14113,N_13823,N_13568);
nand U14114 (N_14114,N_13501,N_13837);
nor U14115 (N_14115,N_13657,N_13684);
nor U14116 (N_14116,N_13585,N_13868);
and U14117 (N_14117,N_13907,N_13925);
xor U14118 (N_14118,N_13806,N_13979);
xnor U14119 (N_14119,N_13683,N_13663);
nand U14120 (N_14120,N_13575,N_13762);
nor U14121 (N_14121,N_13972,N_13745);
nor U14122 (N_14122,N_13509,N_13800);
nand U14123 (N_14123,N_13587,N_13964);
nor U14124 (N_14124,N_13919,N_13635);
nand U14125 (N_14125,N_13619,N_13686);
or U14126 (N_14126,N_13505,N_13877);
or U14127 (N_14127,N_13656,N_13923);
or U14128 (N_14128,N_13694,N_13545);
nor U14129 (N_14129,N_13777,N_13644);
nand U14130 (N_14130,N_13543,N_13740);
xnor U14131 (N_14131,N_13566,N_13603);
nand U14132 (N_14132,N_13572,N_13935);
xnor U14133 (N_14133,N_13847,N_13856);
and U14134 (N_14134,N_13813,N_13810);
xnor U14135 (N_14135,N_13918,N_13909);
nand U14136 (N_14136,N_13562,N_13728);
or U14137 (N_14137,N_13605,N_13807);
or U14138 (N_14138,N_13953,N_13878);
nor U14139 (N_14139,N_13970,N_13899);
or U14140 (N_14140,N_13937,N_13833);
nand U14141 (N_14141,N_13846,N_13815);
or U14142 (N_14142,N_13544,N_13842);
nor U14143 (N_14143,N_13733,N_13711);
xor U14144 (N_14144,N_13739,N_13945);
nand U14145 (N_14145,N_13827,N_13931);
nand U14146 (N_14146,N_13620,N_13814);
nand U14147 (N_14147,N_13622,N_13515);
and U14148 (N_14148,N_13623,N_13808);
xnor U14149 (N_14149,N_13798,N_13672);
or U14150 (N_14150,N_13771,N_13638);
nor U14151 (N_14151,N_13581,N_13778);
nor U14152 (N_14152,N_13651,N_13799);
and U14153 (N_14153,N_13688,N_13670);
and U14154 (N_14154,N_13922,N_13744);
or U14155 (N_14155,N_13606,N_13532);
or U14156 (N_14156,N_13917,N_13936);
xor U14157 (N_14157,N_13851,N_13809);
and U14158 (N_14158,N_13896,N_13741);
and U14159 (N_14159,N_13993,N_13734);
xnor U14160 (N_14160,N_13687,N_13642);
nor U14161 (N_14161,N_13844,N_13848);
nor U14162 (N_14162,N_13789,N_13914);
nor U14163 (N_14163,N_13735,N_13826);
xnor U14164 (N_14164,N_13941,N_13760);
and U14165 (N_14165,N_13697,N_13853);
and U14166 (N_14166,N_13946,N_13752);
and U14167 (N_14167,N_13512,N_13679);
and U14168 (N_14168,N_13548,N_13747);
xor U14169 (N_14169,N_13967,N_13555);
and U14170 (N_14170,N_13506,N_13962);
nor U14171 (N_14171,N_13763,N_13770);
nand U14172 (N_14172,N_13830,N_13535);
xnor U14173 (N_14173,N_13557,N_13502);
nand U14174 (N_14174,N_13886,N_13859);
or U14175 (N_14175,N_13561,N_13738);
and U14176 (N_14176,N_13759,N_13518);
or U14177 (N_14177,N_13757,N_13529);
and U14178 (N_14178,N_13520,N_13794);
or U14179 (N_14179,N_13958,N_13582);
nand U14180 (N_14180,N_13702,N_13674);
xnor U14181 (N_14181,N_13662,N_13869);
nand U14182 (N_14182,N_13822,N_13571);
or U14183 (N_14183,N_13504,N_13879);
nand U14184 (N_14184,N_13732,N_13693);
or U14185 (N_14185,N_13891,N_13767);
nand U14186 (N_14186,N_13895,N_13567);
xnor U14187 (N_14187,N_13628,N_13838);
nor U14188 (N_14188,N_13596,N_13583);
nand U14189 (N_14189,N_13900,N_13659);
or U14190 (N_14190,N_13915,N_13652);
and U14191 (N_14191,N_13764,N_13643);
nor U14192 (N_14192,N_13867,N_13577);
or U14193 (N_14193,N_13973,N_13749);
xnor U14194 (N_14194,N_13880,N_13517);
and U14195 (N_14195,N_13801,N_13669);
or U14196 (N_14196,N_13905,N_13718);
nand U14197 (N_14197,N_13831,N_13610);
xnor U14198 (N_14198,N_13769,N_13677);
and U14199 (N_14199,N_13795,N_13812);
and U14200 (N_14200,N_13576,N_13890);
or U14201 (N_14201,N_13781,N_13536);
nand U14202 (N_14202,N_13768,N_13726);
nand U14203 (N_14203,N_13655,N_13626);
and U14204 (N_14204,N_13819,N_13948);
and U14205 (N_14205,N_13743,N_13957);
xnor U14206 (N_14206,N_13797,N_13924);
nor U14207 (N_14207,N_13641,N_13930);
nand U14208 (N_14208,N_13647,N_13746);
and U14209 (N_14209,N_13579,N_13916);
nor U14210 (N_14210,N_13611,N_13742);
and U14211 (N_14211,N_13666,N_13753);
or U14212 (N_14212,N_13696,N_13811);
nand U14213 (N_14213,N_13714,N_13724);
nand U14214 (N_14214,N_13553,N_13956);
nor U14215 (N_14215,N_13969,N_13639);
nand U14216 (N_14216,N_13772,N_13542);
and U14217 (N_14217,N_13632,N_13608);
nor U14218 (N_14218,N_13756,N_13609);
and U14219 (N_14219,N_13692,N_13614);
and U14220 (N_14220,N_13721,N_13549);
xor U14221 (N_14221,N_13921,N_13987);
xnor U14222 (N_14222,N_13802,N_13586);
nor U14223 (N_14223,N_13720,N_13765);
xor U14224 (N_14224,N_13982,N_13503);
and U14225 (N_14225,N_13825,N_13885);
or U14226 (N_14226,N_13787,N_13554);
and U14227 (N_14227,N_13754,N_13613);
or U14228 (N_14228,N_13624,N_13550);
or U14229 (N_14229,N_13646,N_13782);
and U14230 (N_14230,N_13722,N_13664);
xnor U14231 (N_14231,N_13719,N_13539);
nor U14232 (N_14232,N_13563,N_13514);
and U14233 (N_14233,N_13780,N_13731);
nand U14234 (N_14234,N_13667,N_13913);
and U14235 (N_14235,N_13966,N_13939);
nand U14236 (N_14236,N_13598,N_13883);
xor U14237 (N_14237,N_13897,N_13910);
nor U14238 (N_14238,N_13996,N_13527);
nand U14239 (N_14239,N_13952,N_13933);
nor U14240 (N_14240,N_13901,N_13675);
and U14241 (N_14241,N_13959,N_13961);
nand U14242 (N_14242,N_13864,N_13560);
nand U14243 (N_14243,N_13650,N_13892);
nand U14244 (N_14244,N_13589,N_13578);
nor U14245 (N_14245,N_13893,N_13755);
nand U14246 (N_14246,N_13636,N_13865);
nor U14247 (N_14247,N_13788,N_13929);
nand U14248 (N_14248,N_13978,N_13625);
and U14249 (N_14249,N_13538,N_13888);
xor U14250 (N_14250,N_13931,N_13754);
xnor U14251 (N_14251,N_13768,N_13634);
xor U14252 (N_14252,N_13652,N_13823);
and U14253 (N_14253,N_13816,N_13949);
and U14254 (N_14254,N_13685,N_13780);
nand U14255 (N_14255,N_13688,N_13852);
nand U14256 (N_14256,N_13890,N_13758);
nor U14257 (N_14257,N_13910,N_13671);
or U14258 (N_14258,N_13654,N_13609);
or U14259 (N_14259,N_13897,N_13808);
or U14260 (N_14260,N_13889,N_13568);
nor U14261 (N_14261,N_13668,N_13571);
nand U14262 (N_14262,N_13904,N_13966);
and U14263 (N_14263,N_13748,N_13781);
and U14264 (N_14264,N_13558,N_13757);
and U14265 (N_14265,N_13862,N_13912);
or U14266 (N_14266,N_13906,N_13818);
or U14267 (N_14267,N_13745,N_13867);
nand U14268 (N_14268,N_13686,N_13910);
and U14269 (N_14269,N_13704,N_13740);
nand U14270 (N_14270,N_13804,N_13553);
nor U14271 (N_14271,N_13573,N_13553);
and U14272 (N_14272,N_13960,N_13857);
and U14273 (N_14273,N_13595,N_13862);
xor U14274 (N_14274,N_13959,N_13548);
nor U14275 (N_14275,N_13545,N_13790);
or U14276 (N_14276,N_13808,N_13721);
xnor U14277 (N_14277,N_13572,N_13691);
and U14278 (N_14278,N_13861,N_13820);
nand U14279 (N_14279,N_13678,N_13758);
and U14280 (N_14280,N_13940,N_13681);
and U14281 (N_14281,N_13968,N_13834);
xor U14282 (N_14282,N_13902,N_13566);
or U14283 (N_14283,N_13880,N_13681);
or U14284 (N_14284,N_13881,N_13594);
xor U14285 (N_14285,N_13892,N_13698);
and U14286 (N_14286,N_13762,N_13560);
and U14287 (N_14287,N_13913,N_13603);
and U14288 (N_14288,N_13571,N_13637);
or U14289 (N_14289,N_13924,N_13921);
or U14290 (N_14290,N_13691,N_13501);
xor U14291 (N_14291,N_13633,N_13703);
and U14292 (N_14292,N_13915,N_13598);
xor U14293 (N_14293,N_13570,N_13706);
xnor U14294 (N_14294,N_13922,N_13631);
and U14295 (N_14295,N_13759,N_13674);
nor U14296 (N_14296,N_13819,N_13822);
nor U14297 (N_14297,N_13639,N_13941);
nand U14298 (N_14298,N_13579,N_13880);
nand U14299 (N_14299,N_13886,N_13660);
or U14300 (N_14300,N_13616,N_13571);
and U14301 (N_14301,N_13762,N_13884);
and U14302 (N_14302,N_13949,N_13765);
and U14303 (N_14303,N_13929,N_13645);
nor U14304 (N_14304,N_13849,N_13706);
nand U14305 (N_14305,N_13578,N_13518);
and U14306 (N_14306,N_13883,N_13908);
nor U14307 (N_14307,N_13805,N_13791);
and U14308 (N_14308,N_13801,N_13745);
nand U14309 (N_14309,N_13969,N_13908);
or U14310 (N_14310,N_13860,N_13983);
or U14311 (N_14311,N_13972,N_13707);
nor U14312 (N_14312,N_13707,N_13798);
and U14313 (N_14313,N_13833,N_13641);
xor U14314 (N_14314,N_13502,N_13563);
and U14315 (N_14315,N_13895,N_13815);
or U14316 (N_14316,N_13998,N_13678);
or U14317 (N_14317,N_13993,N_13600);
nor U14318 (N_14318,N_13683,N_13574);
and U14319 (N_14319,N_13556,N_13713);
and U14320 (N_14320,N_13525,N_13819);
and U14321 (N_14321,N_13939,N_13858);
nor U14322 (N_14322,N_13990,N_13683);
nor U14323 (N_14323,N_13538,N_13515);
and U14324 (N_14324,N_13898,N_13790);
nand U14325 (N_14325,N_13501,N_13953);
nor U14326 (N_14326,N_13862,N_13841);
nand U14327 (N_14327,N_13793,N_13983);
nand U14328 (N_14328,N_13533,N_13945);
nand U14329 (N_14329,N_13563,N_13608);
nor U14330 (N_14330,N_13942,N_13564);
xnor U14331 (N_14331,N_13840,N_13587);
nor U14332 (N_14332,N_13590,N_13604);
nor U14333 (N_14333,N_13792,N_13601);
or U14334 (N_14334,N_13657,N_13981);
and U14335 (N_14335,N_13600,N_13800);
and U14336 (N_14336,N_13835,N_13528);
xor U14337 (N_14337,N_13691,N_13963);
and U14338 (N_14338,N_13568,N_13851);
and U14339 (N_14339,N_13833,N_13845);
or U14340 (N_14340,N_13942,N_13934);
and U14341 (N_14341,N_13732,N_13739);
or U14342 (N_14342,N_13541,N_13547);
or U14343 (N_14343,N_13921,N_13507);
and U14344 (N_14344,N_13712,N_13633);
nor U14345 (N_14345,N_13583,N_13533);
nor U14346 (N_14346,N_13871,N_13745);
nand U14347 (N_14347,N_13765,N_13938);
or U14348 (N_14348,N_13964,N_13704);
or U14349 (N_14349,N_13986,N_13709);
and U14350 (N_14350,N_13799,N_13895);
xnor U14351 (N_14351,N_13941,N_13513);
or U14352 (N_14352,N_13529,N_13964);
or U14353 (N_14353,N_13921,N_13721);
xor U14354 (N_14354,N_13998,N_13896);
nor U14355 (N_14355,N_13563,N_13902);
or U14356 (N_14356,N_13561,N_13822);
nand U14357 (N_14357,N_13616,N_13735);
or U14358 (N_14358,N_13796,N_13891);
xor U14359 (N_14359,N_13509,N_13955);
and U14360 (N_14360,N_13534,N_13764);
xor U14361 (N_14361,N_13742,N_13990);
or U14362 (N_14362,N_13812,N_13536);
nand U14363 (N_14363,N_13967,N_13667);
and U14364 (N_14364,N_13721,N_13576);
nor U14365 (N_14365,N_13910,N_13954);
xnor U14366 (N_14366,N_13985,N_13782);
and U14367 (N_14367,N_13909,N_13711);
nor U14368 (N_14368,N_13949,N_13997);
xor U14369 (N_14369,N_13541,N_13524);
or U14370 (N_14370,N_13767,N_13942);
nand U14371 (N_14371,N_13766,N_13800);
xnor U14372 (N_14372,N_13705,N_13932);
or U14373 (N_14373,N_13536,N_13838);
nand U14374 (N_14374,N_13970,N_13595);
nand U14375 (N_14375,N_13916,N_13793);
xor U14376 (N_14376,N_13944,N_13574);
xnor U14377 (N_14377,N_13724,N_13936);
nor U14378 (N_14378,N_13978,N_13556);
xnor U14379 (N_14379,N_13768,N_13530);
and U14380 (N_14380,N_13573,N_13649);
and U14381 (N_14381,N_13692,N_13634);
xor U14382 (N_14382,N_13968,N_13991);
nand U14383 (N_14383,N_13936,N_13932);
nand U14384 (N_14384,N_13991,N_13553);
or U14385 (N_14385,N_13707,N_13955);
nand U14386 (N_14386,N_13620,N_13611);
nor U14387 (N_14387,N_13650,N_13932);
nand U14388 (N_14388,N_13594,N_13609);
or U14389 (N_14389,N_13543,N_13773);
nand U14390 (N_14390,N_13537,N_13627);
nor U14391 (N_14391,N_13970,N_13924);
or U14392 (N_14392,N_13891,N_13868);
or U14393 (N_14393,N_13540,N_13850);
or U14394 (N_14394,N_13994,N_13661);
nor U14395 (N_14395,N_13597,N_13964);
and U14396 (N_14396,N_13536,N_13696);
and U14397 (N_14397,N_13588,N_13794);
or U14398 (N_14398,N_13659,N_13827);
nand U14399 (N_14399,N_13565,N_13829);
nor U14400 (N_14400,N_13583,N_13784);
and U14401 (N_14401,N_13638,N_13731);
or U14402 (N_14402,N_13903,N_13962);
xor U14403 (N_14403,N_13529,N_13649);
or U14404 (N_14404,N_13585,N_13980);
nor U14405 (N_14405,N_13546,N_13970);
nand U14406 (N_14406,N_13583,N_13585);
xor U14407 (N_14407,N_13993,N_13938);
and U14408 (N_14408,N_13765,N_13827);
or U14409 (N_14409,N_13553,N_13687);
or U14410 (N_14410,N_13947,N_13536);
nand U14411 (N_14411,N_13733,N_13672);
nand U14412 (N_14412,N_13530,N_13692);
and U14413 (N_14413,N_13897,N_13919);
or U14414 (N_14414,N_13824,N_13692);
and U14415 (N_14415,N_13949,N_13525);
and U14416 (N_14416,N_13655,N_13686);
nor U14417 (N_14417,N_13551,N_13803);
nand U14418 (N_14418,N_13961,N_13930);
xnor U14419 (N_14419,N_13593,N_13893);
nor U14420 (N_14420,N_13526,N_13858);
and U14421 (N_14421,N_13711,N_13970);
xnor U14422 (N_14422,N_13948,N_13532);
nand U14423 (N_14423,N_13847,N_13641);
or U14424 (N_14424,N_13623,N_13638);
xnor U14425 (N_14425,N_13509,N_13784);
xnor U14426 (N_14426,N_13552,N_13932);
and U14427 (N_14427,N_13728,N_13648);
xor U14428 (N_14428,N_13877,N_13862);
xnor U14429 (N_14429,N_13735,N_13925);
nand U14430 (N_14430,N_13955,N_13595);
nand U14431 (N_14431,N_13812,N_13826);
nor U14432 (N_14432,N_13706,N_13740);
nor U14433 (N_14433,N_13921,N_13820);
nor U14434 (N_14434,N_13716,N_13773);
or U14435 (N_14435,N_13917,N_13518);
nand U14436 (N_14436,N_13630,N_13709);
nand U14437 (N_14437,N_13701,N_13774);
and U14438 (N_14438,N_13517,N_13797);
and U14439 (N_14439,N_13918,N_13571);
or U14440 (N_14440,N_13834,N_13596);
and U14441 (N_14441,N_13543,N_13528);
and U14442 (N_14442,N_13917,N_13640);
nor U14443 (N_14443,N_13596,N_13811);
nand U14444 (N_14444,N_13777,N_13959);
or U14445 (N_14445,N_13836,N_13536);
or U14446 (N_14446,N_13623,N_13941);
xnor U14447 (N_14447,N_13530,N_13897);
nand U14448 (N_14448,N_13711,N_13559);
nand U14449 (N_14449,N_13650,N_13505);
nor U14450 (N_14450,N_13895,N_13995);
nand U14451 (N_14451,N_13921,N_13800);
nand U14452 (N_14452,N_13979,N_13661);
xnor U14453 (N_14453,N_13934,N_13803);
xnor U14454 (N_14454,N_13876,N_13688);
or U14455 (N_14455,N_13537,N_13901);
and U14456 (N_14456,N_13827,N_13777);
xor U14457 (N_14457,N_13997,N_13985);
xor U14458 (N_14458,N_13583,N_13913);
xor U14459 (N_14459,N_13874,N_13983);
nand U14460 (N_14460,N_13838,N_13948);
xnor U14461 (N_14461,N_13728,N_13694);
nor U14462 (N_14462,N_13716,N_13741);
nor U14463 (N_14463,N_13543,N_13578);
or U14464 (N_14464,N_13551,N_13858);
or U14465 (N_14465,N_13694,N_13943);
or U14466 (N_14466,N_13731,N_13536);
xnor U14467 (N_14467,N_13646,N_13516);
nand U14468 (N_14468,N_13843,N_13582);
nor U14469 (N_14469,N_13585,N_13764);
nand U14470 (N_14470,N_13905,N_13860);
and U14471 (N_14471,N_13642,N_13605);
nand U14472 (N_14472,N_13941,N_13643);
nor U14473 (N_14473,N_13788,N_13902);
and U14474 (N_14474,N_13808,N_13530);
or U14475 (N_14475,N_13523,N_13908);
xor U14476 (N_14476,N_13842,N_13533);
and U14477 (N_14477,N_13836,N_13727);
or U14478 (N_14478,N_13860,N_13706);
and U14479 (N_14479,N_13542,N_13684);
nor U14480 (N_14480,N_13865,N_13903);
and U14481 (N_14481,N_13955,N_13846);
xor U14482 (N_14482,N_13950,N_13722);
xnor U14483 (N_14483,N_13594,N_13840);
xor U14484 (N_14484,N_13831,N_13755);
and U14485 (N_14485,N_13658,N_13539);
or U14486 (N_14486,N_13764,N_13861);
nand U14487 (N_14487,N_13607,N_13731);
nor U14488 (N_14488,N_13899,N_13724);
or U14489 (N_14489,N_13687,N_13915);
or U14490 (N_14490,N_13654,N_13547);
nor U14491 (N_14491,N_13795,N_13825);
nand U14492 (N_14492,N_13510,N_13810);
nor U14493 (N_14493,N_13820,N_13737);
and U14494 (N_14494,N_13972,N_13871);
xor U14495 (N_14495,N_13728,N_13817);
and U14496 (N_14496,N_13536,N_13777);
nand U14497 (N_14497,N_13705,N_13880);
nor U14498 (N_14498,N_13590,N_13621);
nand U14499 (N_14499,N_13658,N_13909);
and U14500 (N_14500,N_14127,N_14222);
xor U14501 (N_14501,N_14173,N_14408);
nor U14502 (N_14502,N_14297,N_14451);
or U14503 (N_14503,N_14402,N_14470);
nand U14504 (N_14504,N_14101,N_14434);
xor U14505 (N_14505,N_14036,N_14360);
or U14506 (N_14506,N_14387,N_14287);
nor U14507 (N_14507,N_14060,N_14311);
xnor U14508 (N_14508,N_14213,N_14370);
xnor U14509 (N_14509,N_14167,N_14467);
nor U14510 (N_14510,N_14437,N_14054);
xnor U14511 (N_14511,N_14483,N_14420);
or U14512 (N_14512,N_14361,N_14244);
xor U14513 (N_14513,N_14132,N_14091);
and U14514 (N_14514,N_14455,N_14495);
or U14515 (N_14515,N_14024,N_14089);
xnor U14516 (N_14516,N_14022,N_14034);
nand U14517 (N_14517,N_14227,N_14102);
nor U14518 (N_14518,N_14226,N_14413);
nor U14519 (N_14519,N_14010,N_14358);
nand U14520 (N_14520,N_14302,N_14114);
nand U14521 (N_14521,N_14189,N_14088);
nand U14522 (N_14522,N_14428,N_14400);
nor U14523 (N_14523,N_14016,N_14490);
and U14524 (N_14524,N_14053,N_14169);
or U14525 (N_14525,N_14144,N_14115);
xnor U14526 (N_14526,N_14085,N_14070);
xor U14527 (N_14527,N_14033,N_14039);
nand U14528 (N_14528,N_14069,N_14212);
and U14529 (N_14529,N_14469,N_14136);
and U14530 (N_14530,N_14366,N_14492);
nor U14531 (N_14531,N_14109,N_14152);
and U14532 (N_14532,N_14250,N_14350);
nand U14533 (N_14533,N_14165,N_14186);
nor U14534 (N_14534,N_14268,N_14232);
nor U14535 (N_14535,N_14418,N_14179);
xnor U14536 (N_14536,N_14139,N_14288);
and U14537 (N_14537,N_14267,N_14170);
xor U14538 (N_14538,N_14425,N_14049);
or U14539 (N_14539,N_14454,N_14386);
nand U14540 (N_14540,N_14011,N_14457);
nor U14541 (N_14541,N_14005,N_14471);
and U14542 (N_14542,N_14347,N_14309);
and U14543 (N_14543,N_14100,N_14310);
nor U14544 (N_14544,N_14151,N_14007);
xor U14545 (N_14545,N_14092,N_14211);
xnor U14546 (N_14546,N_14240,N_14415);
xor U14547 (N_14547,N_14161,N_14337);
and U14548 (N_14548,N_14048,N_14018);
nand U14549 (N_14549,N_14369,N_14112);
or U14550 (N_14550,N_14407,N_14330);
or U14551 (N_14551,N_14215,N_14453);
nor U14552 (N_14552,N_14015,N_14285);
or U14553 (N_14553,N_14148,N_14163);
nor U14554 (N_14554,N_14017,N_14234);
nor U14555 (N_14555,N_14411,N_14439);
xnor U14556 (N_14556,N_14318,N_14432);
or U14557 (N_14557,N_14328,N_14294);
or U14558 (N_14558,N_14476,N_14339);
and U14559 (N_14559,N_14023,N_14159);
or U14560 (N_14560,N_14441,N_14198);
nor U14561 (N_14561,N_14459,N_14208);
xnor U14562 (N_14562,N_14394,N_14141);
or U14563 (N_14563,N_14436,N_14218);
or U14564 (N_14564,N_14051,N_14095);
or U14565 (N_14565,N_14303,N_14317);
and U14566 (N_14566,N_14245,N_14143);
nor U14567 (N_14567,N_14073,N_14435);
xnor U14568 (N_14568,N_14351,N_14078);
xor U14569 (N_14569,N_14182,N_14031);
nor U14570 (N_14570,N_14345,N_14364);
nor U14571 (N_14571,N_14375,N_14314);
or U14572 (N_14572,N_14390,N_14162);
xor U14573 (N_14573,N_14461,N_14123);
and U14574 (N_14574,N_14153,N_14188);
or U14575 (N_14575,N_14075,N_14259);
nand U14576 (N_14576,N_14064,N_14154);
xnor U14577 (N_14577,N_14093,N_14325);
nand U14578 (N_14578,N_14197,N_14378);
xnor U14579 (N_14579,N_14032,N_14084);
and U14580 (N_14580,N_14072,N_14142);
or U14581 (N_14581,N_14265,N_14097);
or U14582 (N_14582,N_14104,N_14284);
xnor U14583 (N_14583,N_14125,N_14134);
nand U14584 (N_14584,N_14037,N_14140);
nand U14585 (N_14585,N_14313,N_14487);
or U14586 (N_14586,N_14111,N_14430);
nor U14587 (N_14587,N_14178,N_14044);
nor U14588 (N_14588,N_14449,N_14171);
or U14589 (N_14589,N_14191,N_14296);
or U14590 (N_14590,N_14074,N_14058);
nor U14591 (N_14591,N_14393,N_14399);
nand U14592 (N_14592,N_14202,N_14282);
xor U14593 (N_14593,N_14035,N_14025);
or U14594 (N_14594,N_14298,N_14083);
or U14595 (N_14595,N_14427,N_14331);
nand U14596 (N_14596,N_14175,N_14172);
or U14597 (N_14597,N_14359,N_14086);
or U14598 (N_14598,N_14126,N_14426);
xnor U14599 (N_14599,N_14237,N_14315);
or U14600 (N_14600,N_14105,N_14196);
and U14601 (N_14601,N_14263,N_14241);
and U14602 (N_14602,N_14447,N_14190);
nor U14603 (N_14603,N_14249,N_14365);
and U14604 (N_14604,N_14486,N_14261);
xnor U14605 (N_14605,N_14295,N_14379);
or U14606 (N_14606,N_14368,N_14329);
nor U14607 (N_14607,N_14305,N_14055);
or U14608 (N_14608,N_14343,N_14384);
or U14609 (N_14609,N_14193,N_14248);
nand U14610 (N_14610,N_14019,N_14038);
nand U14611 (N_14611,N_14204,N_14238);
and U14612 (N_14612,N_14416,N_14410);
and U14613 (N_14613,N_14417,N_14401);
nor U14614 (N_14614,N_14405,N_14306);
xor U14615 (N_14615,N_14004,N_14009);
and U14616 (N_14616,N_14499,N_14260);
nand U14617 (N_14617,N_14233,N_14185);
or U14618 (N_14618,N_14342,N_14160);
or U14619 (N_14619,N_14320,N_14409);
xnor U14620 (N_14620,N_14040,N_14349);
xor U14621 (N_14621,N_14258,N_14209);
nor U14622 (N_14622,N_14388,N_14026);
or U14623 (N_14623,N_14485,N_14020);
or U14624 (N_14624,N_14493,N_14116);
xor U14625 (N_14625,N_14444,N_14230);
and U14626 (N_14626,N_14027,N_14062);
or U14627 (N_14627,N_14326,N_14414);
xor U14628 (N_14628,N_14338,N_14164);
and U14629 (N_14629,N_14061,N_14251);
nand U14630 (N_14630,N_14274,N_14276);
or U14631 (N_14631,N_14442,N_14081);
and U14632 (N_14632,N_14429,N_14452);
nand U14633 (N_14633,N_14236,N_14319);
nor U14634 (N_14634,N_14146,N_14045);
nand U14635 (N_14635,N_14067,N_14458);
and U14636 (N_14636,N_14168,N_14118);
or U14637 (N_14637,N_14080,N_14203);
and U14638 (N_14638,N_14356,N_14277);
nor U14639 (N_14639,N_14176,N_14396);
or U14640 (N_14640,N_14113,N_14421);
xor U14641 (N_14641,N_14398,N_14255);
or U14642 (N_14642,N_14281,N_14120);
nor U14643 (N_14643,N_14214,N_14147);
xor U14644 (N_14644,N_14333,N_14316);
and U14645 (N_14645,N_14041,N_14419);
nor U14646 (N_14646,N_14477,N_14353);
xnor U14647 (N_14647,N_14275,N_14014);
xnor U14648 (N_14648,N_14341,N_14229);
xnor U14649 (N_14649,N_14029,N_14108);
and U14650 (N_14650,N_14488,N_14382);
or U14651 (N_14651,N_14256,N_14242);
or U14652 (N_14652,N_14362,N_14464);
and U14653 (N_14653,N_14082,N_14423);
nand U14654 (N_14654,N_14252,N_14050);
nor U14655 (N_14655,N_14220,N_14206);
xnor U14656 (N_14656,N_14231,N_14332);
or U14657 (N_14657,N_14389,N_14498);
xor U14658 (N_14658,N_14106,N_14210);
nand U14659 (N_14659,N_14225,N_14327);
or U14660 (N_14660,N_14395,N_14367);
or U14661 (N_14661,N_14056,N_14481);
xnor U14662 (N_14662,N_14128,N_14119);
nand U14663 (N_14663,N_14266,N_14304);
or U14664 (N_14664,N_14087,N_14107);
or U14665 (N_14665,N_14472,N_14246);
nand U14666 (N_14666,N_14363,N_14181);
or U14667 (N_14667,N_14257,N_14177);
nand U14668 (N_14668,N_14076,N_14496);
or U14669 (N_14669,N_14223,N_14028);
nand U14670 (N_14670,N_14079,N_14059);
nand U14671 (N_14671,N_14494,N_14006);
and U14672 (N_14672,N_14448,N_14099);
or U14673 (N_14673,N_14474,N_14334);
nand U14674 (N_14674,N_14012,N_14003);
or U14675 (N_14675,N_14155,N_14068);
and U14676 (N_14676,N_14446,N_14336);
or U14677 (N_14677,N_14312,N_14270);
nand U14678 (N_14678,N_14480,N_14096);
or U14679 (N_14679,N_14269,N_14090);
xnor U14680 (N_14680,N_14475,N_14158);
nor U14681 (N_14681,N_14385,N_14466);
xor U14682 (N_14682,N_14183,N_14290);
nor U14683 (N_14683,N_14124,N_14219);
and U14684 (N_14684,N_14440,N_14346);
xnor U14685 (N_14685,N_14254,N_14289);
or U14686 (N_14686,N_14323,N_14271);
nor U14687 (N_14687,N_14180,N_14205);
and U14688 (N_14688,N_14130,N_14324);
xor U14689 (N_14689,N_14392,N_14468);
nand U14690 (N_14690,N_14216,N_14235);
xor U14691 (N_14691,N_14431,N_14354);
nor U14692 (N_14692,N_14239,N_14192);
nand U14693 (N_14693,N_14371,N_14133);
and U14694 (N_14694,N_14121,N_14137);
and U14695 (N_14695,N_14110,N_14046);
nor U14696 (N_14696,N_14098,N_14103);
and U14697 (N_14697,N_14057,N_14463);
nand U14698 (N_14698,N_14299,N_14157);
nand U14699 (N_14699,N_14403,N_14000);
and U14700 (N_14700,N_14491,N_14122);
nor U14701 (N_14701,N_14077,N_14465);
nand U14702 (N_14702,N_14307,N_14001);
or U14703 (N_14703,N_14348,N_14042);
and U14704 (N_14704,N_14199,N_14335);
nor U14705 (N_14705,N_14445,N_14300);
or U14706 (N_14706,N_14221,N_14065);
nand U14707 (N_14707,N_14184,N_14374);
xnor U14708 (N_14708,N_14322,N_14352);
nor U14709 (N_14709,N_14373,N_14355);
nand U14710 (N_14710,N_14283,N_14243);
nand U14711 (N_14711,N_14484,N_14482);
xor U14712 (N_14712,N_14145,N_14253);
or U14713 (N_14713,N_14149,N_14383);
xnor U14714 (N_14714,N_14207,N_14397);
or U14715 (N_14715,N_14264,N_14135);
nor U14716 (N_14716,N_14292,N_14456);
nor U14717 (N_14717,N_14412,N_14424);
xnor U14718 (N_14718,N_14344,N_14150);
xnor U14719 (N_14719,N_14247,N_14021);
nand U14720 (N_14720,N_14047,N_14406);
or U14721 (N_14721,N_14478,N_14422);
nand U14722 (N_14722,N_14030,N_14301);
and U14723 (N_14723,N_14156,N_14278);
nor U14724 (N_14724,N_14200,N_14224);
and U14725 (N_14725,N_14450,N_14194);
and U14726 (N_14726,N_14262,N_14201);
xnor U14727 (N_14727,N_14443,N_14228);
nor U14728 (N_14728,N_14340,N_14291);
nor U14729 (N_14729,N_14286,N_14372);
nand U14730 (N_14730,N_14002,N_14166);
or U14731 (N_14731,N_14380,N_14308);
nand U14732 (N_14732,N_14195,N_14489);
nor U14733 (N_14733,N_14217,N_14131);
xnor U14734 (N_14734,N_14008,N_14460);
nand U14735 (N_14735,N_14052,N_14187);
nor U14736 (N_14736,N_14433,N_14381);
nand U14737 (N_14737,N_14043,N_14013);
nor U14738 (N_14738,N_14377,N_14280);
and U14739 (N_14739,N_14293,N_14479);
or U14740 (N_14740,N_14066,N_14438);
nor U14741 (N_14741,N_14497,N_14279);
or U14742 (N_14742,N_14391,N_14063);
nand U14743 (N_14743,N_14462,N_14272);
and U14744 (N_14744,N_14174,N_14473);
xor U14745 (N_14745,N_14071,N_14404);
nand U14746 (N_14746,N_14129,N_14357);
or U14747 (N_14747,N_14094,N_14321);
and U14748 (N_14748,N_14273,N_14376);
xor U14749 (N_14749,N_14138,N_14117);
and U14750 (N_14750,N_14454,N_14145);
nor U14751 (N_14751,N_14016,N_14129);
or U14752 (N_14752,N_14083,N_14481);
or U14753 (N_14753,N_14100,N_14217);
nor U14754 (N_14754,N_14366,N_14405);
and U14755 (N_14755,N_14078,N_14095);
nand U14756 (N_14756,N_14011,N_14055);
nor U14757 (N_14757,N_14212,N_14314);
and U14758 (N_14758,N_14337,N_14432);
nand U14759 (N_14759,N_14242,N_14481);
and U14760 (N_14760,N_14043,N_14483);
nand U14761 (N_14761,N_14268,N_14348);
nor U14762 (N_14762,N_14398,N_14075);
xor U14763 (N_14763,N_14159,N_14286);
or U14764 (N_14764,N_14371,N_14475);
or U14765 (N_14765,N_14111,N_14078);
nor U14766 (N_14766,N_14045,N_14328);
nand U14767 (N_14767,N_14335,N_14260);
or U14768 (N_14768,N_14324,N_14297);
xor U14769 (N_14769,N_14054,N_14002);
nand U14770 (N_14770,N_14395,N_14021);
or U14771 (N_14771,N_14440,N_14168);
nor U14772 (N_14772,N_14436,N_14068);
xnor U14773 (N_14773,N_14342,N_14051);
nand U14774 (N_14774,N_14294,N_14492);
and U14775 (N_14775,N_14245,N_14110);
and U14776 (N_14776,N_14365,N_14306);
nor U14777 (N_14777,N_14138,N_14262);
or U14778 (N_14778,N_14342,N_14462);
nor U14779 (N_14779,N_14151,N_14257);
nand U14780 (N_14780,N_14096,N_14397);
or U14781 (N_14781,N_14028,N_14094);
xor U14782 (N_14782,N_14140,N_14025);
nor U14783 (N_14783,N_14040,N_14045);
and U14784 (N_14784,N_14427,N_14320);
or U14785 (N_14785,N_14190,N_14035);
nor U14786 (N_14786,N_14156,N_14252);
nor U14787 (N_14787,N_14293,N_14120);
and U14788 (N_14788,N_14291,N_14490);
and U14789 (N_14789,N_14304,N_14223);
nand U14790 (N_14790,N_14263,N_14205);
nand U14791 (N_14791,N_14363,N_14404);
nand U14792 (N_14792,N_14083,N_14079);
or U14793 (N_14793,N_14074,N_14448);
xor U14794 (N_14794,N_14474,N_14252);
or U14795 (N_14795,N_14467,N_14113);
xnor U14796 (N_14796,N_14219,N_14095);
nor U14797 (N_14797,N_14468,N_14272);
or U14798 (N_14798,N_14163,N_14052);
nor U14799 (N_14799,N_14102,N_14153);
nor U14800 (N_14800,N_14100,N_14136);
nor U14801 (N_14801,N_14127,N_14223);
nor U14802 (N_14802,N_14076,N_14155);
and U14803 (N_14803,N_14324,N_14087);
xor U14804 (N_14804,N_14161,N_14460);
or U14805 (N_14805,N_14052,N_14249);
nor U14806 (N_14806,N_14064,N_14417);
xnor U14807 (N_14807,N_14438,N_14411);
xnor U14808 (N_14808,N_14366,N_14393);
xnor U14809 (N_14809,N_14188,N_14222);
or U14810 (N_14810,N_14442,N_14400);
and U14811 (N_14811,N_14153,N_14103);
or U14812 (N_14812,N_14268,N_14193);
and U14813 (N_14813,N_14075,N_14241);
and U14814 (N_14814,N_14466,N_14278);
or U14815 (N_14815,N_14338,N_14119);
or U14816 (N_14816,N_14457,N_14246);
nand U14817 (N_14817,N_14436,N_14178);
nand U14818 (N_14818,N_14447,N_14000);
nor U14819 (N_14819,N_14349,N_14305);
and U14820 (N_14820,N_14058,N_14363);
or U14821 (N_14821,N_14418,N_14306);
or U14822 (N_14822,N_14281,N_14006);
and U14823 (N_14823,N_14358,N_14070);
nor U14824 (N_14824,N_14226,N_14235);
or U14825 (N_14825,N_14291,N_14377);
and U14826 (N_14826,N_14409,N_14211);
nand U14827 (N_14827,N_14456,N_14196);
and U14828 (N_14828,N_14424,N_14366);
nand U14829 (N_14829,N_14355,N_14103);
and U14830 (N_14830,N_14435,N_14033);
and U14831 (N_14831,N_14283,N_14438);
xor U14832 (N_14832,N_14146,N_14097);
and U14833 (N_14833,N_14474,N_14201);
nor U14834 (N_14834,N_14160,N_14156);
nand U14835 (N_14835,N_14164,N_14313);
xnor U14836 (N_14836,N_14052,N_14373);
nand U14837 (N_14837,N_14258,N_14485);
nor U14838 (N_14838,N_14070,N_14315);
nand U14839 (N_14839,N_14052,N_14297);
and U14840 (N_14840,N_14271,N_14206);
xnor U14841 (N_14841,N_14247,N_14389);
or U14842 (N_14842,N_14244,N_14389);
and U14843 (N_14843,N_14235,N_14240);
nor U14844 (N_14844,N_14073,N_14272);
nand U14845 (N_14845,N_14116,N_14085);
nand U14846 (N_14846,N_14291,N_14076);
or U14847 (N_14847,N_14422,N_14086);
nand U14848 (N_14848,N_14416,N_14483);
and U14849 (N_14849,N_14495,N_14485);
and U14850 (N_14850,N_14400,N_14305);
xnor U14851 (N_14851,N_14303,N_14105);
xnor U14852 (N_14852,N_14347,N_14174);
or U14853 (N_14853,N_14439,N_14417);
or U14854 (N_14854,N_14023,N_14339);
and U14855 (N_14855,N_14126,N_14127);
and U14856 (N_14856,N_14183,N_14122);
nor U14857 (N_14857,N_14411,N_14409);
and U14858 (N_14858,N_14307,N_14438);
or U14859 (N_14859,N_14444,N_14301);
and U14860 (N_14860,N_14109,N_14051);
nand U14861 (N_14861,N_14036,N_14290);
and U14862 (N_14862,N_14064,N_14133);
xnor U14863 (N_14863,N_14111,N_14063);
nand U14864 (N_14864,N_14161,N_14225);
or U14865 (N_14865,N_14011,N_14156);
nor U14866 (N_14866,N_14226,N_14072);
nor U14867 (N_14867,N_14397,N_14289);
and U14868 (N_14868,N_14481,N_14176);
or U14869 (N_14869,N_14315,N_14185);
nor U14870 (N_14870,N_14122,N_14431);
and U14871 (N_14871,N_14142,N_14217);
and U14872 (N_14872,N_14313,N_14462);
nor U14873 (N_14873,N_14055,N_14332);
nor U14874 (N_14874,N_14368,N_14470);
xnor U14875 (N_14875,N_14341,N_14414);
xnor U14876 (N_14876,N_14279,N_14367);
nor U14877 (N_14877,N_14363,N_14393);
nand U14878 (N_14878,N_14240,N_14184);
nor U14879 (N_14879,N_14271,N_14048);
nand U14880 (N_14880,N_14273,N_14371);
and U14881 (N_14881,N_14220,N_14403);
or U14882 (N_14882,N_14032,N_14072);
nor U14883 (N_14883,N_14463,N_14405);
or U14884 (N_14884,N_14056,N_14132);
nor U14885 (N_14885,N_14247,N_14468);
nand U14886 (N_14886,N_14363,N_14374);
nand U14887 (N_14887,N_14132,N_14073);
or U14888 (N_14888,N_14498,N_14217);
nand U14889 (N_14889,N_14257,N_14279);
xnor U14890 (N_14890,N_14250,N_14208);
nand U14891 (N_14891,N_14139,N_14444);
nand U14892 (N_14892,N_14433,N_14397);
and U14893 (N_14893,N_14087,N_14304);
or U14894 (N_14894,N_14220,N_14175);
nand U14895 (N_14895,N_14050,N_14378);
and U14896 (N_14896,N_14065,N_14363);
and U14897 (N_14897,N_14258,N_14251);
nor U14898 (N_14898,N_14378,N_14370);
nor U14899 (N_14899,N_14321,N_14292);
xor U14900 (N_14900,N_14461,N_14418);
xor U14901 (N_14901,N_14289,N_14017);
nor U14902 (N_14902,N_14489,N_14068);
and U14903 (N_14903,N_14438,N_14349);
and U14904 (N_14904,N_14296,N_14294);
nand U14905 (N_14905,N_14167,N_14349);
or U14906 (N_14906,N_14481,N_14486);
xor U14907 (N_14907,N_14386,N_14139);
nand U14908 (N_14908,N_14494,N_14097);
or U14909 (N_14909,N_14099,N_14430);
and U14910 (N_14910,N_14039,N_14435);
nor U14911 (N_14911,N_14075,N_14332);
nand U14912 (N_14912,N_14056,N_14384);
xor U14913 (N_14913,N_14269,N_14259);
nor U14914 (N_14914,N_14391,N_14364);
and U14915 (N_14915,N_14306,N_14210);
or U14916 (N_14916,N_14217,N_14389);
or U14917 (N_14917,N_14052,N_14303);
and U14918 (N_14918,N_14497,N_14119);
and U14919 (N_14919,N_14378,N_14266);
xor U14920 (N_14920,N_14343,N_14222);
and U14921 (N_14921,N_14093,N_14283);
and U14922 (N_14922,N_14339,N_14248);
xor U14923 (N_14923,N_14168,N_14276);
or U14924 (N_14924,N_14135,N_14452);
nand U14925 (N_14925,N_14158,N_14066);
and U14926 (N_14926,N_14139,N_14248);
and U14927 (N_14927,N_14169,N_14346);
xor U14928 (N_14928,N_14056,N_14354);
or U14929 (N_14929,N_14082,N_14415);
nor U14930 (N_14930,N_14448,N_14239);
and U14931 (N_14931,N_14323,N_14263);
xnor U14932 (N_14932,N_14345,N_14342);
nor U14933 (N_14933,N_14089,N_14407);
xor U14934 (N_14934,N_14100,N_14097);
xor U14935 (N_14935,N_14497,N_14428);
or U14936 (N_14936,N_14009,N_14024);
and U14937 (N_14937,N_14058,N_14462);
nor U14938 (N_14938,N_14064,N_14362);
or U14939 (N_14939,N_14074,N_14196);
xor U14940 (N_14940,N_14223,N_14436);
or U14941 (N_14941,N_14369,N_14045);
and U14942 (N_14942,N_14300,N_14291);
and U14943 (N_14943,N_14112,N_14363);
and U14944 (N_14944,N_14284,N_14286);
xor U14945 (N_14945,N_14469,N_14075);
nand U14946 (N_14946,N_14423,N_14119);
nand U14947 (N_14947,N_14166,N_14467);
nor U14948 (N_14948,N_14084,N_14013);
xnor U14949 (N_14949,N_14225,N_14428);
or U14950 (N_14950,N_14252,N_14075);
or U14951 (N_14951,N_14419,N_14240);
or U14952 (N_14952,N_14179,N_14312);
nand U14953 (N_14953,N_14167,N_14221);
xor U14954 (N_14954,N_14409,N_14125);
nor U14955 (N_14955,N_14032,N_14068);
or U14956 (N_14956,N_14456,N_14478);
and U14957 (N_14957,N_14034,N_14020);
or U14958 (N_14958,N_14444,N_14051);
xor U14959 (N_14959,N_14090,N_14137);
and U14960 (N_14960,N_14395,N_14447);
or U14961 (N_14961,N_14268,N_14427);
nand U14962 (N_14962,N_14489,N_14174);
nor U14963 (N_14963,N_14129,N_14315);
nand U14964 (N_14964,N_14323,N_14388);
xor U14965 (N_14965,N_14314,N_14202);
or U14966 (N_14966,N_14256,N_14363);
and U14967 (N_14967,N_14175,N_14176);
and U14968 (N_14968,N_14177,N_14105);
nor U14969 (N_14969,N_14447,N_14084);
nand U14970 (N_14970,N_14140,N_14197);
xor U14971 (N_14971,N_14280,N_14109);
xor U14972 (N_14972,N_14173,N_14397);
nand U14973 (N_14973,N_14227,N_14036);
and U14974 (N_14974,N_14042,N_14015);
or U14975 (N_14975,N_14174,N_14456);
or U14976 (N_14976,N_14464,N_14201);
nand U14977 (N_14977,N_14291,N_14494);
nand U14978 (N_14978,N_14354,N_14043);
or U14979 (N_14979,N_14407,N_14041);
and U14980 (N_14980,N_14484,N_14091);
xnor U14981 (N_14981,N_14363,N_14101);
or U14982 (N_14982,N_14402,N_14111);
and U14983 (N_14983,N_14088,N_14196);
and U14984 (N_14984,N_14436,N_14394);
xnor U14985 (N_14985,N_14233,N_14144);
or U14986 (N_14986,N_14234,N_14011);
xor U14987 (N_14987,N_14286,N_14024);
xor U14988 (N_14988,N_14129,N_14419);
xnor U14989 (N_14989,N_14446,N_14025);
nor U14990 (N_14990,N_14404,N_14089);
and U14991 (N_14991,N_14009,N_14019);
or U14992 (N_14992,N_14300,N_14315);
and U14993 (N_14993,N_14347,N_14436);
and U14994 (N_14994,N_14393,N_14018);
nor U14995 (N_14995,N_14235,N_14412);
and U14996 (N_14996,N_14080,N_14377);
nand U14997 (N_14997,N_14338,N_14418);
nor U14998 (N_14998,N_14172,N_14107);
nor U14999 (N_14999,N_14167,N_14341);
and U15000 (N_15000,N_14622,N_14852);
nor U15001 (N_15001,N_14587,N_14659);
xnor U15002 (N_15002,N_14706,N_14891);
nand U15003 (N_15003,N_14855,N_14901);
and U15004 (N_15004,N_14524,N_14859);
nor U15005 (N_15005,N_14800,N_14988);
nand U15006 (N_15006,N_14872,N_14608);
or U15007 (N_15007,N_14580,N_14658);
nor U15008 (N_15008,N_14983,N_14644);
nand U15009 (N_15009,N_14812,N_14536);
nand U15010 (N_15010,N_14705,N_14760);
or U15011 (N_15011,N_14992,N_14876);
and U15012 (N_15012,N_14703,N_14900);
nor U15013 (N_15013,N_14878,N_14778);
nor U15014 (N_15014,N_14953,N_14591);
nand U15015 (N_15015,N_14964,N_14578);
nand U15016 (N_15016,N_14875,N_14813);
nor U15017 (N_15017,N_14736,N_14694);
and U15018 (N_15018,N_14827,N_14600);
or U15019 (N_15019,N_14885,N_14848);
and U15020 (N_15020,N_14929,N_14503);
nor U15021 (N_15021,N_14502,N_14850);
xor U15022 (N_15022,N_14571,N_14533);
xor U15023 (N_15023,N_14621,N_14595);
nor U15024 (N_15024,N_14635,N_14923);
nor U15025 (N_15025,N_14755,N_14687);
xnor U15026 (N_15026,N_14742,N_14551);
nand U15027 (N_15027,N_14728,N_14548);
nand U15028 (N_15028,N_14828,N_14961);
nand U15029 (N_15029,N_14904,N_14699);
nand U15030 (N_15030,N_14683,N_14797);
and U15031 (N_15031,N_14604,N_14973);
or U15032 (N_15032,N_14881,N_14997);
and U15033 (N_15033,N_14836,N_14814);
nand U15034 (N_15034,N_14761,N_14725);
or U15035 (N_15035,N_14739,N_14529);
xor U15036 (N_15036,N_14652,N_14949);
nor U15037 (N_15037,N_14523,N_14669);
and U15038 (N_15038,N_14612,N_14646);
xor U15039 (N_15039,N_14528,N_14806);
and U15040 (N_15040,N_14897,N_14856);
and U15041 (N_15041,N_14803,N_14557);
xnor U15042 (N_15042,N_14584,N_14666);
or U15043 (N_15043,N_14989,N_14768);
nor U15044 (N_15044,N_14990,N_14713);
nor U15045 (N_15045,N_14624,N_14509);
nand U15046 (N_15046,N_14746,N_14723);
and U15047 (N_15047,N_14782,N_14642);
xor U15048 (N_15048,N_14999,N_14516);
nor U15049 (N_15049,N_14701,N_14920);
xnor U15050 (N_15050,N_14545,N_14847);
xor U15051 (N_15051,N_14838,N_14960);
xnor U15052 (N_15052,N_14686,N_14977);
and U15053 (N_15053,N_14511,N_14741);
or U15054 (N_15054,N_14914,N_14919);
nor U15055 (N_15055,N_14765,N_14996);
nor U15056 (N_15056,N_14559,N_14573);
nand U15057 (N_15057,N_14508,N_14944);
xnor U15058 (N_15058,N_14500,N_14849);
xnor U15059 (N_15059,N_14611,N_14665);
nor U15060 (N_15060,N_14909,N_14517);
nor U15061 (N_15061,N_14547,N_14718);
nor U15062 (N_15062,N_14958,N_14799);
nand U15063 (N_15063,N_14592,N_14921);
xor U15064 (N_15064,N_14777,N_14530);
nor U15065 (N_15065,N_14829,N_14796);
xor U15066 (N_15066,N_14966,N_14771);
nor U15067 (N_15067,N_14939,N_14752);
nor U15068 (N_15068,N_14609,N_14926);
nor U15069 (N_15069,N_14776,N_14884);
nand U15070 (N_15070,N_14772,N_14626);
xnor U15071 (N_15071,N_14844,N_14916);
nor U15072 (N_15072,N_14714,N_14896);
or U15073 (N_15073,N_14678,N_14541);
xnor U15074 (N_15074,N_14815,N_14750);
or U15075 (N_15075,N_14676,N_14662);
or U15076 (N_15076,N_14864,N_14861);
nand U15077 (N_15077,N_14915,N_14586);
xor U15078 (N_15078,N_14906,N_14791);
or U15079 (N_15079,N_14538,N_14846);
nand U15080 (N_15080,N_14629,N_14692);
or U15081 (N_15081,N_14860,N_14719);
and U15082 (N_15082,N_14954,N_14691);
xnor U15083 (N_15083,N_14959,N_14733);
xnor U15084 (N_15084,N_14637,N_14638);
and U15085 (N_15085,N_14531,N_14950);
nand U15086 (N_15086,N_14756,N_14636);
nor U15087 (N_15087,N_14851,N_14552);
and U15088 (N_15088,N_14596,N_14873);
xor U15089 (N_15089,N_14895,N_14730);
and U15090 (N_15090,N_14729,N_14534);
or U15091 (N_15091,N_14822,N_14633);
nor U15092 (N_15092,N_14764,N_14722);
nand U15093 (N_15093,N_14708,N_14887);
nor U15094 (N_15094,N_14841,N_14918);
xnor U15095 (N_15095,N_14689,N_14734);
and U15096 (N_15096,N_14598,N_14537);
nor U15097 (N_15097,N_14707,N_14933);
and U15098 (N_15098,N_14677,N_14525);
nand U15099 (N_15099,N_14518,N_14858);
nand U15100 (N_15100,N_14780,N_14601);
and U15101 (N_15101,N_14630,N_14614);
nand U15102 (N_15102,N_14668,N_14819);
or U15103 (N_15103,N_14942,N_14656);
xor U15104 (N_15104,N_14971,N_14737);
and U15105 (N_15105,N_14907,N_14807);
nor U15106 (N_15106,N_14721,N_14912);
and U15107 (N_15107,N_14540,N_14744);
or U15108 (N_15108,N_14974,N_14899);
nor U15109 (N_15109,N_14978,N_14618);
xnor U15110 (N_15110,N_14790,N_14615);
or U15111 (N_15111,N_14902,N_14663);
nor U15112 (N_15112,N_14634,N_14697);
nor U15113 (N_15113,N_14947,N_14786);
nor U15114 (N_15114,N_14987,N_14565);
or U15115 (N_15115,N_14743,N_14857);
and U15116 (N_15116,N_14882,N_14564);
nor U15117 (N_15117,N_14754,N_14930);
nand U15118 (N_15118,N_14785,N_14970);
and U15119 (N_15119,N_14879,N_14821);
nand U15120 (N_15120,N_14962,N_14566);
xnor U15121 (N_15121,N_14763,N_14616);
or U15122 (N_15122,N_14769,N_14554);
xor U15123 (N_15123,N_14753,N_14766);
xor U15124 (N_15124,N_14539,N_14917);
nand U15125 (N_15125,N_14910,N_14787);
nand U15126 (N_15126,N_14886,N_14575);
nor U15127 (N_15127,N_14675,N_14762);
xnor U15128 (N_15128,N_14567,N_14967);
xnor U15129 (N_15129,N_14613,N_14617);
nand U15130 (N_15130,N_14653,N_14643);
or U15131 (N_15131,N_14840,N_14507);
and U15132 (N_15132,N_14550,N_14681);
nand U15133 (N_15133,N_14660,N_14811);
and U15134 (N_15134,N_14673,N_14981);
nand U15135 (N_15135,N_14808,N_14968);
and U15136 (N_15136,N_14732,N_14506);
nor U15137 (N_15137,N_14903,N_14986);
xor U15138 (N_15138,N_14854,N_14976);
nor U15139 (N_15139,N_14957,N_14560);
or U15140 (N_15140,N_14735,N_14520);
nand U15141 (N_15141,N_14757,N_14670);
nand U15142 (N_15142,N_14955,N_14985);
nand U15143 (N_15143,N_14579,N_14831);
nand U15144 (N_15144,N_14883,N_14843);
nand U15145 (N_15145,N_14606,N_14969);
and U15146 (N_15146,N_14866,N_14794);
and U15147 (N_15147,N_14783,N_14809);
or U15148 (N_15148,N_14569,N_14948);
xnor U15149 (N_15149,N_14504,N_14823);
or U15150 (N_15150,N_14519,N_14710);
nand U15151 (N_15151,N_14908,N_14758);
and U15152 (N_15152,N_14943,N_14995);
and U15153 (N_15153,N_14647,N_14830);
and U15154 (N_15154,N_14817,N_14927);
xor U15155 (N_15155,N_14684,N_14574);
xor U15156 (N_15156,N_14898,N_14657);
nor U15157 (N_15157,N_14980,N_14583);
and U15158 (N_15158,N_14543,N_14698);
and U15159 (N_15159,N_14610,N_14640);
and U15160 (N_15160,N_14715,N_14568);
and U15161 (N_15161,N_14946,N_14824);
nor U15162 (N_15162,N_14702,N_14625);
and U15163 (N_15163,N_14514,N_14655);
and U15164 (N_15164,N_14816,N_14561);
or U15165 (N_15165,N_14804,N_14679);
and U15166 (N_15166,N_14521,N_14795);
nand U15167 (N_15167,N_14720,N_14553);
nor U15168 (N_15168,N_14863,N_14928);
nand U15169 (N_15169,N_14745,N_14805);
nor U15170 (N_15170,N_14938,N_14682);
nand U15171 (N_15171,N_14798,N_14749);
or U15172 (N_15172,N_14667,N_14770);
nand U15173 (N_15173,N_14818,N_14724);
and U15174 (N_15174,N_14738,N_14716);
and U15175 (N_15175,N_14650,N_14802);
nor U15176 (N_15176,N_14842,N_14501);
nor U15177 (N_15177,N_14853,N_14688);
nor U15178 (N_15178,N_14868,N_14651);
or U15179 (N_15179,N_14700,N_14839);
nor U15180 (N_15180,N_14513,N_14696);
nand U15181 (N_15181,N_14972,N_14890);
or U15182 (N_15182,N_14727,N_14937);
or U15183 (N_15183,N_14620,N_14825);
or U15184 (N_15184,N_14639,N_14789);
nand U15185 (N_15185,N_14894,N_14993);
xnor U15186 (N_15186,N_14632,N_14645);
nor U15187 (N_15187,N_14712,N_14674);
and U15188 (N_15188,N_14704,N_14747);
nand U15189 (N_15189,N_14685,N_14549);
nand U15190 (N_15190,N_14963,N_14784);
nand U15191 (N_15191,N_14711,N_14982);
or U15192 (N_15192,N_14767,N_14588);
nand U15193 (N_15193,N_14623,N_14690);
xor U15194 (N_15194,N_14631,N_14932);
xor U15195 (N_15195,N_14751,N_14865);
nor U15196 (N_15196,N_14781,N_14922);
nor U15197 (N_15197,N_14563,N_14542);
or U15198 (N_15198,N_14773,N_14979);
xnor U15199 (N_15199,N_14582,N_14880);
xor U15200 (N_15200,N_14867,N_14505);
or U15201 (N_15201,N_14834,N_14936);
nand U15202 (N_15202,N_14759,N_14991);
xor U15203 (N_15203,N_14510,N_14585);
xnor U15204 (N_15204,N_14562,N_14941);
and U15205 (N_15205,N_14810,N_14717);
nor U15206 (N_15206,N_14820,N_14654);
nor U15207 (N_15207,N_14874,N_14593);
or U15208 (N_15208,N_14792,N_14998);
or U15209 (N_15209,N_14905,N_14925);
xnor U15210 (N_15210,N_14913,N_14793);
and U15211 (N_15211,N_14649,N_14862);
and U15212 (N_15212,N_14602,N_14581);
xnor U15213 (N_15213,N_14779,N_14870);
nor U15214 (N_15214,N_14788,N_14837);
xor U15215 (N_15215,N_14695,N_14731);
or U15216 (N_15216,N_14774,N_14556);
and U15217 (N_15217,N_14570,N_14603);
xor U15218 (N_15218,N_14835,N_14871);
and U15219 (N_15219,N_14893,N_14619);
and U15220 (N_15220,N_14911,N_14589);
xor U15221 (N_15221,N_14597,N_14672);
nor U15222 (N_15222,N_14935,N_14693);
nand U15223 (N_15223,N_14877,N_14522);
and U15224 (N_15224,N_14975,N_14576);
nor U15225 (N_15225,N_14648,N_14607);
xor U15226 (N_15226,N_14984,N_14605);
nor U15227 (N_15227,N_14572,N_14546);
nor U15228 (N_15228,N_14709,N_14931);
nand U15229 (N_15229,N_14740,N_14832);
or U15230 (N_15230,N_14934,N_14532);
and U15231 (N_15231,N_14775,N_14994);
and U15232 (N_15232,N_14952,N_14527);
xor U15233 (N_15233,N_14833,N_14535);
nor U15234 (N_15234,N_14555,N_14594);
xor U15235 (N_15235,N_14845,N_14515);
and U15236 (N_15236,N_14641,N_14924);
xnor U15237 (N_15237,N_14590,N_14544);
or U15238 (N_15238,N_14748,N_14558);
xnor U15239 (N_15239,N_14965,N_14869);
nor U15240 (N_15240,N_14661,N_14726);
xor U15241 (N_15241,N_14680,N_14512);
nor U15242 (N_15242,N_14888,N_14951);
and U15243 (N_15243,N_14627,N_14801);
or U15244 (N_15244,N_14956,N_14892);
or U15245 (N_15245,N_14577,N_14628);
and U15246 (N_15246,N_14826,N_14671);
nand U15247 (N_15247,N_14889,N_14945);
xor U15248 (N_15248,N_14940,N_14599);
or U15249 (N_15249,N_14664,N_14526);
xnor U15250 (N_15250,N_14855,N_14958);
nor U15251 (N_15251,N_14641,N_14945);
or U15252 (N_15252,N_14589,N_14705);
and U15253 (N_15253,N_14765,N_14718);
nand U15254 (N_15254,N_14526,N_14590);
nor U15255 (N_15255,N_14994,N_14604);
and U15256 (N_15256,N_14648,N_14750);
nand U15257 (N_15257,N_14784,N_14806);
or U15258 (N_15258,N_14942,N_14664);
xor U15259 (N_15259,N_14935,N_14835);
nor U15260 (N_15260,N_14914,N_14888);
and U15261 (N_15261,N_14558,N_14607);
nand U15262 (N_15262,N_14964,N_14953);
nor U15263 (N_15263,N_14838,N_14970);
or U15264 (N_15264,N_14588,N_14692);
and U15265 (N_15265,N_14894,N_14562);
or U15266 (N_15266,N_14727,N_14525);
xor U15267 (N_15267,N_14544,N_14594);
and U15268 (N_15268,N_14860,N_14762);
or U15269 (N_15269,N_14936,N_14663);
nor U15270 (N_15270,N_14508,N_14846);
or U15271 (N_15271,N_14811,N_14711);
nand U15272 (N_15272,N_14603,N_14961);
and U15273 (N_15273,N_14567,N_14820);
and U15274 (N_15274,N_14865,N_14631);
nor U15275 (N_15275,N_14793,N_14847);
or U15276 (N_15276,N_14852,N_14564);
xnor U15277 (N_15277,N_14783,N_14971);
nor U15278 (N_15278,N_14615,N_14943);
or U15279 (N_15279,N_14778,N_14663);
xor U15280 (N_15280,N_14975,N_14663);
and U15281 (N_15281,N_14613,N_14971);
xor U15282 (N_15282,N_14599,N_14539);
and U15283 (N_15283,N_14739,N_14988);
nand U15284 (N_15284,N_14988,N_14573);
nand U15285 (N_15285,N_14521,N_14724);
nor U15286 (N_15286,N_14901,N_14920);
nor U15287 (N_15287,N_14835,N_14777);
or U15288 (N_15288,N_14585,N_14501);
xnor U15289 (N_15289,N_14672,N_14917);
and U15290 (N_15290,N_14864,N_14823);
and U15291 (N_15291,N_14687,N_14839);
nand U15292 (N_15292,N_14792,N_14844);
nor U15293 (N_15293,N_14513,N_14518);
xnor U15294 (N_15294,N_14986,N_14736);
nor U15295 (N_15295,N_14526,N_14925);
or U15296 (N_15296,N_14923,N_14876);
or U15297 (N_15297,N_14559,N_14643);
or U15298 (N_15298,N_14513,N_14576);
nor U15299 (N_15299,N_14576,N_14595);
nor U15300 (N_15300,N_14955,N_14878);
xnor U15301 (N_15301,N_14798,N_14733);
nand U15302 (N_15302,N_14730,N_14744);
nand U15303 (N_15303,N_14683,N_14702);
xor U15304 (N_15304,N_14912,N_14904);
or U15305 (N_15305,N_14895,N_14953);
or U15306 (N_15306,N_14616,N_14544);
nor U15307 (N_15307,N_14745,N_14677);
xor U15308 (N_15308,N_14796,N_14965);
nand U15309 (N_15309,N_14573,N_14793);
or U15310 (N_15310,N_14784,N_14592);
xor U15311 (N_15311,N_14958,N_14587);
or U15312 (N_15312,N_14819,N_14936);
and U15313 (N_15313,N_14917,N_14719);
nand U15314 (N_15314,N_14817,N_14699);
xnor U15315 (N_15315,N_14974,N_14548);
xor U15316 (N_15316,N_14587,N_14644);
nor U15317 (N_15317,N_14576,N_14800);
and U15318 (N_15318,N_14767,N_14699);
xor U15319 (N_15319,N_14807,N_14770);
or U15320 (N_15320,N_14664,N_14966);
xor U15321 (N_15321,N_14822,N_14891);
nor U15322 (N_15322,N_14531,N_14941);
and U15323 (N_15323,N_14800,N_14898);
and U15324 (N_15324,N_14554,N_14529);
and U15325 (N_15325,N_14672,N_14566);
and U15326 (N_15326,N_14689,N_14770);
or U15327 (N_15327,N_14619,N_14916);
and U15328 (N_15328,N_14930,N_14511);
xor U15329 (N_15329,N_14625,N_14780);
nor U15330 (N_15330,N_14534,N_14907);
nand U15331 (N_15331,N_14759,N_14952);
nor U15332 (N_15332,N_14876,N_14971);
xnor U15333 (N_15333,N_14767,N_14688);
nor U15334 (N_15334,N_14866,N_14646);
xor U15335 (N_15335,N_14765,N_14860);
xnor U15336 (N_15336,N_14574,N_14946);
and U15337 (N_15337,N_14690,N_14687);
or U15338 (N_15338,N_14818,N_14863);
nor U15339 (N_15339,N_14618,N_14921);
and U15340 (N_15340,N_14736,N_14578);
and U15341 (N_15341,N_14560,N_14606);
and U15342 (N_15342,N_14916,N_14693);
nand U15343 (N_15343,N_14824,N_14767);
nand U15344 (N_15344,N_14670,N_14846);
and U15345 (N_15345,N_14600,N_14940);
and U15346 (N_15346,N_14992,N_14819);
and U15347 (N_15347,N_14860,N_14518);
and U15348 (N_15348,N_14880,N_14668);
nor U15349 (N_15349,N_14915,N_14906);
and U15350 (N_15350,N_14909,N_14573);
and U15351 (N_15351,N_14569,N_14762);
nand U15352 (N_15352,N_14965,N_14636);
and U15353 (N_15353,N_14714,N_14507);
nor U15354 (N_15354,N_14971,N_14577);
nor U15355 (N_15355,N_14788,N_14846);
xor U15356 (N_15356,N_14680,N_14984);
nand U15357 (N_15357,N_14696,N_14738);
nor U15358 (N_15358,N_14856,N_14952);
or U15359 (N_15359,N_14893,N_14548);
or U15360 (N_15360,N_14565,N_14503);
or U15361 (N_15361,N_14797,N_14899);
or U15362 (N_15362,N_14805,N_14513);
nand U15363 (N_15363,N_14830,N_14786);
or U15364 (N_15364,N_14752,N_14868);
xnor U15365 (N_15365,N_14552,N_14867);
and U15366 (N_15366,N_14909,N_14695);
xnor U15367 (N_15367,N_14794,N_14740);
or U15368 (N_15368,N_14884,N_14943);
or U15369 (N_15369,N_14687,N_14589);
nand U15370 (N_15370,N_14959,N_14711);
xnor U15371 (N_15371,N_14689,N_14706);
xor U15372 (N_15372,N_14910,N_14974);
and U15373 (N_15373,N_14762,N_14728);
or U15374 (N_15374,N_14709,N_14832);
and U15375 (N_15375,N_14950,N_14976);
and U15376 (N_15376,N_14731,N_14875);
or U15377 (N_15377,N_14569,N_14809);
nand U15378 (N_15378,N_14572,N_14761);
xor U15379 (N_15379,N_14555,N_14581);
xnor U15380 (N_15380,N_14559,N_14690);
nand U15381 (N_15381,N_14744,N_14844);
nand U15382 (N_15382,N_14801,N_14968);
nor U15383 (N_15383,N_14624,N_14852);
nor U15384 (N_15384,N_14780,N_14592);
or U15385 (N_15385,N_14545,N_14578);
or U15386 (N_15386,N_14642,N_14707);
xor U15387 (N_15387,N_14653,N_14574);
nor U15388 (N_15388,N_14528,N_14755);
or U15389 (N_15389,N_14882,N_14553);
nand U15390 (N_15390,N_14722,N_14828);
xor U15391 (N_15391,N_14664,N_14910);
nand U15392 (N_15392,N_14618,N_14808);
xor U15393 (N_15393,N_14981,N_14828);
or U15394 (N_15394,N_14902,N_14940);
or U15395 (N_15395,N_14757,N_14725);
nand U15396 (N_15396,N_14569,N_14660);
xnor U15397 (N_15397,N_14639,N_14865);
xnor U15398 (N_15398,N_14750,N_14850);
or U15399 (N_15399,N_14883,N_14624);
xnor U15400 (N_15400,N_14779,N_14702);
nor U15401 (N_15401,N_14545,N_14947);
or U15402 (N_15402,N_14610,N_14573);
and U15403 (N_15403,N_14740,N_14749);
xor U15404 (N_15404,N_14591,N_14912);
nor U15405 (N_15405,N_14964,N_14823);
nor U15406 (N_15406,N_14767,N_14750);
nand U15407 (N_15407,N_14601,N_14750);
or U15408 (N_15408,N_14799,N_14695);
xnor U15409 (N_15409,N_14851,N_14731);
or U15410 (N_15410,N_14573,N_14628);
nor U15411 (N_15411,N_14535,N_14528);
and U15412 (N_15412,N_14736,N_14690);
nor U15413 (N_15413,N_14788,N_14508);
and U15414 (N_15414,N_14697,N_14685);
xnor U15415 (N_15415,N_14513,N_14586);
xor U15416 (N_15416,N_14987,N_14729);
nor U15417 (N_15417,N_14558,N_14676);
nand U15418 (N_15418,N_14971,N_14675);
or U15419 (N_15419,N_14565,N_14722);
nor U15420 (N_15420,N_14886,N_14670);
nor U15421 (N_15421,N_14721,N_14948);
nor U15422 (N_15422,N_14792,N_14866);
and U15423 (N_15423,N_14952,N_14771);
and U15424 (N_15424,N_14659,N_14795);
xnor U15425 (N_15425,N_14712,N_14810);
nand U15426 (N_15426,N_14921,N_14992);
or U15427 (N_15427,N_14952,N_14700);
xor U15428 (N_15428,N_14530,N_14880);
nor U15429 (N_15429,N_14594,N_14801);
or U15430 (N_15430,N_14594,N_14810);
xnor U15431 (N_15431,N_14780,N_14725);
nand U15432 (N_15432,N_14961,N_14980);
nor U15433 (N_15433,N_14553,N_14898);
and U15434 (N_15434,N_14832,N_14821);
nor U15435 (N_15435,N_14693,N_14957);
or U15436 (N_15436,N_14636,N_14521);
nand U15437 (N_15437,N_14780,N_14977);
nor U15438 (N_15438,N_14506,N_14798);
nor U15439 (N_15439,N_14638,N_14904);
and U15440 (N_15440,N_14690,N_14871);
and U15441 (N_15441,N_14770,N_14700);
nand U15442 (N_15442,N_14819,N_14804);
xnor U15443 (N_15443,N_14804,N_14898);
nor U15444 (N_15444,N_14900,N_14904);
and U15445 (N_15445,N_14761,N_14940);
xor U15446 (N_15446,N_14988,N_14608);
xnor U15447 (N_15447,N_14965,N_14547);
and U15448 (N_15448,N_14940,N_14950);
xnor U15449 (N_15449,N_14649,N_14929);
nand U15450 (N_15450,N_14929,N_14911);
and U15451 (N_15451,N_14595,N_14783);
nor U15452 (N_15452,N_14620,N_14748);
nand U15453 (N_15453,N_14531,N_14543);
xnor U15454 (N_15454,N_14506,N_14927);
nor U15455 (N_15455,N_14737,N_14852);
xor U15456 (N_15456,N_14712,N_14867);
xor U15457 (N_15457,N_14988,N_14954);
xnor U15458 (N_15458,N_14716,N_14811);
xor U15459 (N_15459,N_14982,N_14536);
and U15460 (N_15460,N_14848,N_14999);
nand U15461 (N_15461,N_14847,N_14515);
xor U15462 (N_15462,N_14761,N_14835);
nand U15463 (N_15463,N_14686,N_14661);
xnor U15464 (N_15464,N_14810,N_14658);
nor U15465 (N_15465,N_14947,N_14823);
or U15466 (N_15466,N_14593,N_14923);
or U15467 (N_15467,N_14830,N_14568);
and U15468 (N_15468,N_14795,N_14513);
nor U15469 (N_15469,N_14670,N_14566);
nor U15470 (N_15470,N_14917,N_14741);
xor U15471 (N_15471,N_14819,N_14685);
xor U15472 (N_15472,N_14726,N_14649);
nor U15473 (N_15473,N_14932,N_14989);
xor U15474 (N_15474,N_14532,N_14945);
nand U15475 (N_15475,N_14926,N_14986);
xnor U15476 (N_15476,N_14545,N_14932);
and U15477 (N_15477,N_14718,N_14859);
and U15478 (N_15478,N_14833,N_14857);
and U15479 (N_15479,N_14959,N_14625);
and U15480 (N_15480,N_14630,N_14813);
and U15481 (N_15481,N_14610,N_14647);
nor U15482 (N_15482,N_14814,N_14566);
nor U15483 (N_15483,N_14888,N_14820);
and U15484 (N_15484,N_14597,N_14666);
xnor U15485 (N_15485,N_14556,N_14913);
xor U15486 (N_15486,N_14647,N_14757);
xor U15487 (N_15487,N_14945,N_14592);
or U15488 (N_15488,N_14804,N_14799);
and U15489 (N_15489,N_14875,N_14520);
nand U15490 (N_15490,N_14796,N_14647);
nand U15491 (N_15491,N_14591,N_14922);
or U15492 (N_15492,N_14816,N_14804);
or U15493 (N_15493,N_14868,N_14729);
nor U15494 (N_15494,N_14587,N_14722);
and U15495 (N_15495,N_14640,N_14577);
and U15496 (N_15496,N_14797,N_14721);
xor U15497 (N_15497,N_14860,N_14922);
nor U15498 (N_15498,N_14985,N_14506);
nor U15499 (N_15499,N_14886,N_14754);
nand U15500 (N_15500,N_15050,N_15189);
and U15501 (N_15501,N_15122,N_15120);
xnor U15502 (N_15502,N_15184,N_15239);
xnor U15503 (N_15503,N_15023,N_15195);
nand U15504 (N_15504,N_15290,N_15046);
nand U15505 (N_15505,N_15430,N_15223);
and U15506 (N_15506,N_15498,N_15291);
nand U15507 (N_15507,N_15328,N_15325);
or U15508 (N_15508,N_15116,N_15049);
and U15509 (N_15509,N_15481,N_15053);
or U15510 (N_15510,N_15034,N_15105);
and U15511 (N_15511,N_15370,N_15406);
or U15512 (N_15512,N_15231,N_15271);
and U15513 (N_15513,N_15044,N_15383);
xnor U15514 (N_15514,N_15075,N_15155);
nor U15515 (N_15515,N_15003,N_15356);
nand U15516 (N_15516,N_15019,N_15115);
or U15517 (N_15517,N_15061,N_15359);
nor U15518 (N_15518,N_15489,N_15079);
or U15519 (N_15519,N_15149,N_15274);
xor U15520 (N_15520,N_15399,N_15418);
nor U15521 (N_15521,N_15107,N_15211);
and U15522 (N_15522,N_15166,N_15277);
nor U15523 (N_15523,N_15371,N_15192);
and U15524 (N_15524,N_15462,N_15222);
or U15525 (N_15525,N_15386,N_15276);
nand U15526 (N_15526,N_15013,N_15329);
and U15527 (N_15527,N_15187,N_15445);
and U15528 (N_15528,N_15012,N_15497);
nand U15529 (N_15529,N_15146,N_15089);
and U15530 (N_15530,N_15478,N_15472);
or U15531 (N_15531,N_15473,N_15190);
and U15532 (N_15532,N_15315,N_15269);
and U15533 (N_15533,N_15167,N_15141);
or U15534 (N_15534,N_15416,N_15470);
nor U15535 (N_15535,N_15303,N_15310);
nand U15536 (N_15536,N_15449,N_15298);
xnor U15537 (N_15537,N_15273,N_15227);
xor U15538 (N_15538,N_15048,N_15431);
nand U15539 (N_15539,N_15495,N_15127);
xnor U15540 (N_15540,N_15461,N_15330);
xnor U15541 (N_15541,N_15086,N_15217);
and U15542 (N_15542,N_15186,N_15073);
or U15543 (N_15543,N_15218,N_15492);
nand U15544 (N_15544,N_15448,N_15459);
nor U15545 (N_15545,N_15027,N_15382);
or U15546 (N_15546,N_15368,N_15069);
nor U15547 (N_15547,N_15327,N_15425);
or U15548 (N_15548,N_15389,N_15142);
xor U15549 (N_15549,N_15214,N_15245);
xnor U15550 (N_15550,N_15018,N_15159);
or U15551 (N_15551,N_15098,N_15407);
xor U15552 (N_15552,N_15280,N_15204);
xnor U15553 (N_15553,N_15283,N_15347);
xnor U15554 (N_15554,N_15236,N_15056);
and U15555 (N_15555,N_15196,N_15096);
or U15556 (N_15556,N_15343,N_15080);
xnor U15557 (N_15557,N_15051,N_15188);
or U15558 (N_15558,N_15243,N_15033);
and U15559 (N_15559,N_15409,N_15474);
nor U15560 (N_15560,N_15026,N_15207);
and U15561 (N_15561,N_15494,N_15248);
and U15562 (N_15562,N_15471,N_15008);
nand U15563 (N_15563,N_15464,N_15309);
nand U15564 (N_15564,N_15452,N_15446);
or U15565 (N_15565,N_15077,N_15094);
nand U15566 (N_15566,N_15466,N_15060);
or U15567 (N_15567,N_15138,N_15366);
or U15568 (N_15568,N_15337,N_15191);
or U15569 (N_15569,N_15093,N_15154);
and U15570 (N_15570,N_15261,N_15219);
or U15571 (N_15571,N_15180,N_15288);
or U15572 (N_15572,N_15287,N_15254);
and U15573 (N_15573,N_15450,N_15110);
nor U15574 (N_15574,N_15394,N_15365);
or U15575 (N_15575,N_15139,N_15112);
xnor U15576 (N_15576,N_15106,N_15224);
nor U15577 (N_15577,N_15091,N_15314);
xnor U15578 (N_15578,N_15342,N_15028);
xor U15579 (N_15579,N_15210,N_15170);
nand U15580 (N_15580,N_15125,N_15379);
or U15581 (N_15581,N_15378,N_15304);
and U15582 (N_15582,N_15320,N_15117);
xor U15583 (N_15583,N_15296,N_15083);
and U15584 (N_15584,N_15024,N_15424);
nand U15585 (N_15585,N_15221,N_15468);
nor U15586 (N_15586,N_15388,N_15144);
xnor U15587 (N_15587,N_15369,N_15259);
or U15588 (N_15588,N_15066,N_15151);
nor U15589 (N_15589,N_15133,N_15163);
xor U15590 (N_15590,N_15410,N_15247);
xor U15591 (N_15591,N_15148,N_15453);
nor U15592 (N_15592,N_15006,N_15486);
nand U15593 (N_15593,N_15145,N_15490);
nand U15594 (N_15594,N_15266,N_15316);
nor U15595 (N_15595,N_15414,N_15264);
xnor U15596 (N_15596,N_15252,N_15121);
or U15597 (N_15597,N_15438,N_15011);
nand U15598 (N_15598,N_15367,N_15174);
and U15599 (N_15599,N_15401,N_15415);
nor U15600 (N_15600,N_15479,N_15268);
xnor U15601 (N_15601,N_15043,N_15391);
or U15602 (N_15602,N_15020,N_15016);
and U15603 (N_15603,N_15162,N_15040);
nor U15604 (N_15604,N_15168,N_15052);
xnor U15605 (N_15605,N_15226,N_15015);
or U15606 (N_15606,N_15228,N_15114);
nand U15607 (N_15607,N_15467,N_15358);
and U15608 (N_15608,N_15351,N_15451);
nand U15609 (N_15609,N_15436,N_15035);
xnor U15610 (N_15610,N_15156,N_15045);
or U15611 (N_15611,N_15336,N_15143);
and U15612 (N_15612,N_15477,N_15411);
nand U15613 (N_15613,N_15179,N_15463);
or U15614 (N_15614,N_15305,N_15161);
and U15615 (N_15615,N_15055,N_15341);
and U15616 (N_15616,N_15130,N_15102);
nand U15617 (N_15617,N_15443,N_15281);
nor U15618 (N_15618,N_15334,N_15126);
xor U15619 (N_15619,N_15289,N_15491);
nor U15620 (N_15620,N_15284,N_15308);
xor U15621 (N_15621,N_15128,N_15447);
or U15622 (N_15622,N_15256,N_15054);
nand U15623 (N_15623,N_15201,N_15230);
xor U15624 (N_15624,N_15009,N_15482);
xnor U15625 (N_15625,N_15483,N_15339);
and U15626 (N_15626,N_15119,N_15381);
nor U15627 (N_15627,N_15025,N_15345);
nor U15628 (N_15628,N_15004,N_15360);
nor U15629 (N_15629,N_15299,N_15353);
or U15630 (N_15630,N_15213,N_15272);
xnor U15631 (N_15631,N_15387,N_15169);
nor U15632 (N_15632,N_15235,N_15318);
nor U15633 (N_15633,N_15460,N_15307);
nand U15634 (N_15634,N_15417,N_15469);
nor U15635 (N_15635,N_15402,N_15253);
nand U15636 (N_15636,N_15263,N_15331);
nand U15637 (N_15637,N_15042,N_15076);
nor U15638 (N_15638,N_15302,N_15319);
nand U15639 (N_15639,N_15136,N_15005);
nand U15640 (N_15640,N_15442,N_15282);
nor U15641 (N_15641,N_15275,N_15301);
and U15642 (N_15642,N_15420,N_15255);
and U15643 (N_15643,N_15181,N_15123);
nor U15644 (N_15644,N_15002,N_15432);
or U15645 (N_15645,N_15278,N_15140);
nor U15646 (N_15646,N_15375,N_15017);
nand U15647 (N_15647,N_15022,N_15398);
nor U15648 (N_15648,N_15074,N_15376);
nor U15649 (N_15649,N_15109,N_15380);
xor U15650 (N_15650,N_15242,N_15030);
nand U15651 (N_15651,N_15372,N_15182);
nor U15652 (N_15652,N_15465,N_15000);
xnor U15653 (N_15653,N_15279,N_15158);
and U15654 (N_15654,N_15374,N_15185);
nand U15655 (N_15655,N_15476,N_15362);
nand U15656 (N_15656,N_15010,N_15039);
or U15657 (N_15657,N_15260,N_15103);
and U15658 (N_15658,N_15232,N_15496);
nand U15659 (N_15659,N_15108,N_15499);
or U15660 (N_15660,N_15220,N_15404);
xnor U15661 (N_15661,N_15295,N_15234);
xor U15662 (N_15662,N_15064,N_15072);
and U15663 (N_15663,N_15292,N_15286);
or U15664 (N_15664,N_15317,N_15062);
and U15665 (N_15665,N_15240,N_15193);
nor U15666 (N_15666,N_15421,N_15036);
nand U15667 (N_15667,N_15311,N_15238);
and U15668 (N_15668,N_15124,N_15338);
nand U15669 (N_15669,N_15428,N_15225);
xnor U15670 (N_15670,N_15396,N_15400);
nand U15671 (N_15671,N_15206,N_15194);
nor U15672 (N_15672,N_15348,N_15087);
nor U15673 (N_15673,N_15095,N_15029);
or U15674 (N_15674,N_15397,N_15198);
or U15675 (N_15675,N_15200,N_15419);
nand U15676 (N_15676,N_15135,N_15427);
or U15677 (N_15677,N_15067,N_15097);
and U15678 (N_15678,N_15444,N_15147);
nand U15679 (N_15679,N_15199,N_15249);
and U15680 (N_15680,N_15059,N_15405);
nor U15681 (N_15681,N_15165,N_15300);
nand U15682 (N_15682,N_15364,N_15433);
or U15683 (N_15683,N_15031,N_15014);
or U15684 (N_15684,N_15333,N_15313);
xor U15685 (N_15685,N_15392,N_15173);
or U15686 (N_15686,N_15340,N_15384);
nor U15687 (N_15687,N_15423,N_15251);
xor U15688 (N_15688,N_15244,N_15084);
or U15689 (N_15689,N_15395,N_15480);
or U15690 (N_15690,N_15385,N_15457);
and U15691 (N_15691,N_15322,N_15434);
nor U15692 (N_15692,N_15326,N_15485);
nand U15693 (N_15693,N_15041,N_15032);
or U15694 (N_15694,N_15101,N_15373);
xor U15695 (N_15695,N_15203,N_15175);
xnor U15696 (N_15696,N_15306,N_15357);
nand U15697 (N_15697,N_15354,N_15335);
and U15698 (N_15698,N_15177,N_15440);
or U15699 (N_15699,N_15202,N_15323);
xnor U15700 (N_15700,N_15007,N_15346);
nand U15701 (N_15701,N_15349,N_15350);
or U15702 (N_15702,N_15090,N_15352);
xnor U15703 (N_15703,N_15257,N_15171);
and U15704 (N_15704,N_15137,N_15412);
and U15705 (N_15705,N_15312,N_15092);
xnor U15706 (N_15706,N_15267,N_15437);
xnor U15707 (N_15707,N_15429,N_15355);
nand U15708 (N_15708,N_15152,N_15081);
nor U15709 (N_15709,N_15229,N_15160);
nand U15710 (N_15710,N_15250,N_15332);
or U15711 (N_15711,N_15361,N_15068);
xor U15712 (N_15712,N_15393,N_15297);
nor U15713 (N_15713,N_15208,N_15403);
nand U15714 (N_15714,N_15455,N_15293);
xnor U15715 (N_15715,N_15088,N_15183);
nor U15716 (N_15716,N_15426,N_15484);
and U15717 (N_15717,N_15265,N_15413);
xor U15718 (N_15718,N_15001,N_15065);
xnor U15719 (N_15719,N_15131,N_15132);
or U15720 (N_15720,N_15111,N_15258);
nand U15721 (N_15721,N_15118,N_15233);
nor U15722 (N_15722,N_15104,N_15172);
nor U15723 (N_15723,N_15197,N_15176);
xor U15724 (N_15724,N_15205,N_15129);
or U15725 (N_15725,N_15237,N_15475);
xor U15726 (N_15726,N_15082,N_15441);
nand U15727 (N_15727,N_15408,N_15134);
xnor U15728 (N_15728,N_15100,N_15270);
and U15729 (N_15729,N_15324,N_15078);
nand U15730 (N_15730,N_15458,N_15456);
or U15731 (N_15731,N_15212,N_15215);
nor U15732 (N_15732,N_15285,N_15153);
xor U15733 (N_15733,N_15363,N_15262);
nor U15734 (N_15734,N_15157,N_15099);
and U15735 (N_15735,N_15294,N_15085);
or U15736 (N_15736,N_15241,N_15487);
nor U15737 (N_15737,N_15377,N_15164);
and U15738 (N_15738,N_15493,N_15038);
nand U15739 (N_15739,N_15209,N_15390);
and U15740 (N_15740,N_15037,N_15435);
nand U15741 (N_15741,N_15021,N_15454);
xnor U15742 (N_15742,N_15216,N_15439);
nor U15743 (N_15743,N_15057,N_15071);
nor U15744 (N_15744,N_15070,N_15422);
nor U15745 (N_15745,N_15321,N_15178);
xor U15746 (N_15746,N_15113,N_15344);
or U15747 (N_15747,N_15488,N_15047);
nor U15748 (N_15748,N_15063,N_15150);
nor U15749 (N_15749,N_15246,N_15058);
xnor U15750 (N_15750,N_15471,N_15452);
nand U15751 (N_15751,N_15406,N_15222);
or U15752 (N_15752,N_15330,N_15321);
nand U15753 (N_15753,N_15413,N_15350);
and U15754 (N_15754,N_15144,N_15471);
and U15755 (N_15755,N_15065,N_15092);
and U15756 (N_15756,N_15474,N_15280);
and U15757 (N_15757,N_15296,N_15010);
or U15758 (N_15758,N_15292,N_15167);
or U15759 (N_15759,N_15040,N_15019);
or U15760 (N_15760,N_15441,N_15102);
and U15761 (N_15761,N_15345,N_15145);
nand U15762 (N_15762,N_15441,N_15440);
xor U15763 (N_15763,N_15026,N_15140);
nor U15764 (N_15764,N_15348,N_15044);
xnor U15765 (N_15765,N_15200,N_15376);
and U15766 (N_15766,N_15227,N_15328);
xor U15767 (N_15767,N_15471,N_15010);
and U15768 (N_15768,N_15148,N_15447);
xnor U15769 (N_15769,N_15420,N_15016);
xnor U15770 (N_15770,N_15193,N_15235);
xor U15771 (N_15771,N_15436,N_15232);
or U15772 (N_15772,N_15122,N_15085);
xnor U15773 (N_15773,N_15182,N_15106);
xnor U15774 (N_15774,N_15249,N_15172);
and U15775 (N_15775,N_15378,N_15435);
and U15776 (N_15776,N_15114,N_15414);
xnor U15777 (N_15777,N_15251,N_15010);
nor U15778 (N_15778,N_15019,N_15084);
and U15779 (N_15779,N_15342,N_15012);
nand U15780 (N_15780,N_15000,N_15306);
or U15781 (N_15781,N_15048,N_15350);
xor U15782 (N_15782,N_15258,N_15342);
or U15783 (N_15783,N_15320,N_15149);
and U15784 (N_15784,N_15246,N_15006);
nor U15785 (N_15785,N_15456,N_15415);
xor U15786 (N_15786,N_15047,N_15128);
and U15787 (N_15787,N_15358,N_15029);
or U15788 (N_15788,N_15122,N_15030);
and U15789 (N_15789,N_15216,N_15212);
xnor U15790 (N_15790,N_15348,N_15123);
xnor U15791 (N_15791,N_15167,N_15218);
xor U15792 (N_15792,N_15043,N_15493);
or U15793 (N_15793,N_15375,N_15178);
nand U15794 (N_15794,N_15038,N_15150);
and U15795 (N_15795,N_15097,N_15113);
xnor U15796 (N_15796,N_15370,N_15044);
and U15797 (N_15797,N_15116,N_15308);
nor U15798 (N_15798,N_15431,N_15142);
or U15799 (N_15799,N_15067,N_15025);
or U15800 (N_15800,N_15451,N_15058);
xnor U15801 (N_15801,N_15374,N_15397);
or U15802 (N_15802,N_15464,N_15440);
or U15803 (N_15803,N_15043,N_15479);
nor U15804 (N_15804,N_15299,N_15101);
xor U15805 (N_15805,N_15207,N_15397);
nand U15806 (N_15806,N_15304,N_15416);
and U15807 (N_15807,N_15129,N_15234);
and U15808 (N_15808,N_15137,N_15333);
xor U15809 (N_15809,N_15379,N_15332);
xnor U15810 (N_15810,N_15094,N_15345);
or U15811 (N_15811,N_15197,N_15280);
and U15812 (N_15812,N_15029,N_15233);
nand U15813 (N_15813,N_15322,N_15044);
and U15814 (N_15814,N_15261,N_15083);
nor U15815 (N_15815,N_15327,N_15256);
and U15816 (N_15816,N_15483,N_15070);
nand U15817 (N_15817,N_15343,N_15103);
and U15818 (N_15818,N_15289,N_15201);
xnor U15819 (N_15819,N_15488,N_15327);
xnor U15820 (N_15820,N_15065,N_15426);
and U15821 (N_15821,N_15498,N_15383);
nor U15822 (N_15822,N_15068,N_15436);
or U15823 (N_15823,N_15115,N_15235);
nand U15824 (N_15824,N_15332,N_15173);
and U15825 (N_15825,N_15318,N_15183);
or U15826 (N_15826,N_15412,N_15087);
nor U15827 (N_15827,N_15150,N_15032);
xor U15828 (N_15828,N_15266,N_15242);
nand U15829 (N_15829,N_15188,N_15334);
nor U15830 (N_15830,N_15354,N_15020);
nor U15831 (N_15831,N_15350,N_15432);
xnor U15832 (N_15832,N_15153,N_15452);
xor U15833 (N_15833,N_15258,N_15144);
nor U15834 (N_15834,N_15265,N_15461);
nand U15835 (N_15835,N_15389,N_15382);
nand U15836 (N_15836,N_15430,N_15447);
nor U15837 (N_15837,N_15364,N_15483);
and U15838 (N_15838,N_15343,N_15330);
nor U15839 (N_15839,N_15464,N_15199);
nand U15840 (N_15840,N_15011,N_15177);
xor U15841 (N_15841,N_15132,N_15316);
xor U15842 (N_15842,N_15343,N_15133);
nand U15843 (N_15843,N_15080,N_15359);
xor U15844 (N_15844,N_15388,N_15056);
nand U15845 (N_15845,N_15310,N_15106);
or U15846 (N_15846,N_15071,N_15378);
and U15847 (N_15847,N_15131,N_15096);
or U15848 (N_15848,N_15406,N_15211);
or U15849 (N_15849,N_15470,N_15140);
nor U15850 (N_15850,N_15282,N_15250);
xor U15851 (N_15851,N_15345,N_15481);
or U15852 (N_15852,N_15457,N_15496);
nand U15853 (N_15853,N_15283,N_15239);
or U15854 (N_15854,N_15228,N_15277);
and U15855 (N_15855,N_15314,N_15155);
nand U15856 (N_15856,N_15088,N_15242);
nand U15857 (N_15857,N_15042,N_15087);
xnor U15858 (N_15858,N_15134,N_15016);
or U15859 (N_15859,N_15007,N_15442);
nand U15860 (N_15860,N_15442,N_15037);
xor U15861 (N_15861,N_15384,N_15198);
xnor U15862 (N_15862,N_15290,N_15159);
nand U15863 (N_15863,N_15241,N_15481);
nor U15864 (N_15864,N_15142,N_15174);
or U15865 (N_15865,N_15046,N_15339);
and U15866 (N_15866,N_15077,N_15013);
nor U15867 (N_15867,N_15230,N_15032);
nand U15868 (N_15868,N_15490,N_15395);
or U15869 (N_15869,N_15039,N_15237);
and U15870 (N_15870,N_15226,N_15332);
and U15871 (N_15871,N_15198,N_15104);
xor U15872 (N_15872,N_15126,N_15464);
xnor U15873 (N_15873,N_15317,N_15345);
and U15874 (N_15874,N_15229,N_15034);
xor U15875 (N_15875,N_15207,N_15233);
or U15876 (N_15876,N_15077,N_15335);
xnor U15877 (N_15877,N_15320,N_15284);
and U15878 (N_15878,N_15203,N_15337);
nand U15879 (N_15879,N_15108,N_15290);
and U15880 (N_15880,N_15060,N_15107);
xor U15881 (N_15881,N_15390,N_15329);
and U15882 (N_15882,N_15338,N_15045);
nand U15883 (N_15883,N_15374,N_15388);
nor U15884 (N_15884,N_15124,N_15214);
or U15885 (N_15885,N_15043,N_15112);
and U15886 (N_15886,N_15434,N_15425);
nor U15887 (N_15887,N_15118,N_15023);
and U15888 (N_15888,N_15253,N_15287);
nor U15889 (N_15889,N_15081,N_15145);
xor U15890 (N_15890,N_15256,N_15446);
and U15891 (N_15891,N_15405,N_15252);
nand U15892 (N_15892,N_15097,N_15374);
xnor U15893 (N_15893,N_15340,N_15344);
and U15894 (N_15894,N_15244,N_15321);
nor U15895 (N_15895,N_15481,N_15117);
nor U15896 (N_15896,N_15109,N_15034);
xnor U15897 (N_15897,N_15217,N_15199);
nor U15898 (N_15898,N_15365,N_15400);
nor U15899 (N_15899,N_15070,N_15445);
nand U15900 (N_15900,N_15083,N_15176);
nand U15901 (N_15901,N_15415,N_15017);
nand U15902 (N_15902,N_15304,N_15051);
or U15903 (N_15903,N_15106,N_15280);
and U15904 (N_15904,N_15155,N_15312);
or U15905 (N_15905,N_15459,N_15386);
and U15906 (N_15906,N_15086,N_15339);
xnor U15907 (N_15907,N_15024,N_15416);
nor U15908 (N_15908,N_15391,N_15477);
xnor U15909 (N_15909,N_15242,N_15317);
or U15910 (N_15910,N_15026,N_15401);
nand U15911 (N_15911,N_15235,N_15356);
nor U15912 (N_15912,N_15454,N_15102);
nand U15913 (N_15913,N_15380,N_15226);
nor U15914 (N_15914,N_15342,N_15061);
xor U15915 (N_15915,N_15315,N_15388);
or U15916 (N_15916,N_15328,N_15137);
xor U15917 (N_15917,N_15195,N_15484);
xor U15918 (N_15918,N_15005,N_15343);
xnor U15919 (N_15919,N_15072,N_15326);
or U15920 (N_15920,N_15284,N_15271);
nor U15921 (N_15921,N_15199,N_15116);
xnor U15922 (N_15922,N_15381,N_15267);
nor U15923 (N_15923,N_15215,N_15408);
and U15924 (N_15924,N_15027,N_15291);
xor U15925 (N_15925,N_15415,N_15469);
xnor U15926 (N_15926,N_15435,N_15002);
xor U15927 (N_15927,N_15131,N_15216);
xnor U15928 (N_15928,N_15471,N_15281);
or U15929 (N_15929,N_15144,N_15262);
xor U15930 (N_15930,N_15407,N_15241);
nor U15931 (N_15931,N_15322,N_15215);
nor U15932 (N_15932,N_15227,N_15234);
xnor U15933 (N_15933,N_15140,N_15041);
nand U15934 (N_15934,N_15025,N_15087);
nor U15935 (N_15935,N_15002,N_15171);
or U15936 (N_15936,N_15134,N_15234);
and U15937 (N_15937,N_15128,N_15205);
nand U15938 (N_15938,N_15167,N_15192);
or U15939 (N_15939,N_15470,N_15195);
xnor U15940 (N_15940,N_15195,N_15372);
or U15941 (N_15941,N_15475,N_15005);
xnor U15942 (N_15942,N_15059,N_15478);
or U15943 (N_15943,N_15347,N_15300);
nor U15944 (N_15944,N_15070,N_15220);
nand U15945 (N_15945,N_15209,N_15167);
xor U15946 (N_15946,N_15334,N_15336);
nand U15947 (N_15947,N_15303,N_15426);
nor U15948 (N_15948,N_15476,N_15333);
nand U15949 (N_15949,N_15375,N_15072);
xor U15950 (N_15950,N_15220,N_15045);
nand U15951 (N_15951,N_15271,N_15021);
xnor U15952 (N_15952,N_15227,N_15441);
nand U15953 (N_15953,N_15483,N_15015);
and U15954 (N_15954,N_15416,N_15045);
nor U15955 (N_15955,N_15355,N_15335);
and U15956 (N_15956,N_15352,N_15426);
nand U15957 (N_15957,N_15027,N_15253);
nor U15958 (N_15958,N_15287,N_15433);
nand U15959 (N_15959,N_15202,N_15096);
or U15960 (N_15960,N_15233,N_15362);
xnor U15961 (N_15961,N_15400,N_15075);
and U15962 (N_15962,N_15368,N_15424);
or U15963 (N_15963,N_15117,N_15467);
and U15964 (N_15964,N_15073,N_15074);
nand U15965 (N_15965,N_15360,N_15060);
nand U15966 (N_15966,N_15033,N_15059);
or U15967 (N_15967,N_15401,N_15369);
and U15968 (N_15968,N_15004,N_15484);
or U15969 (N_15969,N_15093,N_15491);
xor U15970 (N_15970,N_15406,N_15408);
and U15971 (N_15971,N_15254,N_15491);
nand U15972 (N_15972,N_15210,N_15418);
or U15973 (N_15973,N_15268,N_15476);
nand U15974 (N_15974,N_15096,N_15188);
or U15975 (N_15975,N_15201,N_15212);
nor U15976 (N_15976,N_15228,N_15102);
and U15977 (N_15977,N_15134,N_15482);
xnor U15978 (N_15978,N_15198,N_15478);
nand U15979 (N_15979,N_15131,N_15006);
nand U15980 (N_15980,N_15496,N_15257);
nor U15981 (N_15981,N_15279,N_15076);
or U15982 (N_15982,N_15394,N_15100);
and U15983 (N_15983,N_15305,N_15190);
xor U15984 (N_15984,N_15222,N_15022);
nor U15985 (N_15985,N_15297,N_15269);
xor U15986 (N_15986,N_15368,N_15358);
or U15987 (N_15987,N_15114,N_15446);
xor U15988 (N_15988,N_15343,N_15050);
and U15989 (N_15989,N_15224,N_15322);
nor U15990 (N_15990,N_15289,N_15299);
nor U15991 (N_15991,N_15331,N_15365);
or U15992 (N_15992,N_15204,N_15003);
nand U15993 (N_15993,N_15480,N_15398);
or U15994 (N_15994,N_15450,N_15189);
xnor U15995 (N_15995,N_15414,N_15373);
nand U15996 (N_15996,N_15269,N_15258);
xnor U15997 (N_15997,N_15251,N_15074);
or U15998 (N_15998,N_15245,N_15464);
nor U15999 (N_15999,N_15327,N_15090);
and U16000 (N_16000,N_15988,N_15820);
or U16001 (N_16001,N_15792,N_15670);
or U16002 (N_16002,N_15680,N_15803);
xor U16003 (N_16003,N_15991,N_15763);
nor U16004 (N_16004,N_15566,N_15855);
nand U16005 (N_16005,N_15709,N_15989);
xor U16006 (N_16006,N_15722,N_15664);
nand U16007 (N_16007,N_15537,N_15922);
xnor U16008 (N_16008,N_15714,N_15668);
xnor U16009 (N_16009,N_15758,N_15913);
xor U16010 (N_16010,N_15757,N_15928);
nor U16011 (N_16011,N_15572,N_15614);
or U16012 (N_16012,N_15765,N_15834);
nand U16013 (N_16013,N_15607,N_15675);
or U16014 (N_16014,N_15587,N_15511);
xor U16015 (N_16015,N_15947,N_15903);
or U16016 (N_16016,N_15900,N_15643);
nor U16017 (N_16017,N_15731,N_15919);
nand U16018 (N_16018,N_15997,N_15770);
and U16019 (N_16019,N_15801,N_15743);
nand U16020 (N_16020,N_15817,N_15759);
nor U16021 (N_16021,N_15767,N_15982);
or U16022 (N_16022,N_15964,N_15550);
xnor U16023 (N_16023,N_15619,N_15836);
and U16024 (N_16024,N_15823,N_15569);
nand U16025 (N_16025,N_15527,N_15628);
and U16026 (N_16026,N_15910,N_15993);
nor U16027 (N_16027,N_15760,N_15916);
nor U16028 (N_16028,N_15719,N_15673);
and U16029 (N_16029,N_15662,N_15521);
nor U16030 (N_16030,N_15963,N_15816);
nand U16031 (N_16031,N_15694,N_15589);
or U16032 (N_16032,N_15700,N_15808);
or U16033 (N_16033,N_15917,N_15854);
nor U16034 (N_16034,N_15889,N_15898);
nor U16035 (N_16035,N_15818,N_15725);
nand U16036 (N_16036,N_15639,N_15815);
and U16037 (N_16037,N_15807,N_15875);
or U16038 (N_16038,N_15755,N_15789);
nand U16039 (N_16039,N_15519,N_15548);
xor U16040 (N_16040,N_15772,N_15973);
xnor U16041 (N_16041,N_15575,N_15790);
and U16042 (N_16042,N_15682,N_15976);
nand U16043 (N_16043,N_15800,N_15959);
nor U16044 (N_16044,N_15515,N_15971);
xor U16045 (N_16045,N_15653,N_15857);
or U16046 (N_16046,N_15661,N_15779);
nor U16047 (N_16047,N_15736,N_15509);
nand U16048 (N_16048,N_15631,N_15549);
xnor U16049 (N_16049,N_15874,N_15970);
nor U16050 (N_16050,N_15992,N_15825);
or U16051 (N_16051,N_15565,N_15996);
xnor U16052 (N_16052,N_15564,N_15932);
nor U16053 (N_16053,N_15858,N_15873);
nor U16054 (N_16054,N_15708,N_15877);
nand U16055 (N_16055,N_15711,N_15588);
nand U16056 (N_16056,N_15697,N_15707);
nor U16057 (N_16057,N_15824,N_15597);
xnor U16058 (N_16058,N_15863,N_15543);
xnor U16059 (N_16059,N_15615,N_15741);
nand U16060 (N_16060,N_15925,N_15582);
xor U16061 (N_16061,N_15799,N_15721);
nand U16062 (N_16062,N_15848,N_15654);
or U16063 (N_16063,N_15897,N_15881);
xnor U16064 (N_16064,N_15752,N_15906);
xor U16065 (N_16065,N_15835,N_15526);
and U16066 (N_16066,N_15570,N_15787);
nand U16067 (N_16067,N_15936,N_15567);
nor U16068 (N_16068,N_15551,N_15583);
nor U16069 (N_16069,N_15649,N_15638);
and U16070 (N_16070,N_15500,N_15561);
nor U16071 (N_16071,N_15702,N_15621);
and U16072 (N_16072,N_15609,N_15893);
nand U16073 (N_16073,N_15821,N_15958);
or U16074 (N_16074,N_15861,N_15876);
nand U16075 (N_16075,N_15555,N_15987);
nand U16076 (N_16076,N_15746,N_15655);
and U16077 (N_16077,N_15745,N_15592);
xnor U16078 (N_16078,N_15979,N_15882);
or U16079 (N_16079,N_15930,N_15980);
or U16080 (N_16080,N_15749,N_15831);
nor U16081 (N_16081,N_15774,N_15556);
nor U16082 (N_16082,N_15810,N_15802);
xor U16083 (N_16083,N_15524,N_15623);
nand U16084 (N_16084,N_15689,N_15942);
nor U16085 (N_16085,N_15776,N_15921);
nand U16086 (N_16086,N_15690,N_15571);
or U16087 (N_16087,N_15616,N_15613);
and U16088 (N_16088,N_15778,N_15813);
xnor U16089 (N_16089,N_15832,N_15775);
nand U16090 (N_16090,N_15842,N_15559);
or U16091 (N_16091,N_15819,N_15657);
or U16092 (N_16092,N_15594,N_15918);
or U16093 (N_16093,N_15652,N_15599);
or U16094 (N_16094,N_15705,N_15733);
xnor U16095 (N_16095,N_15972,N_15637);
xnor U16096 (N_16096,N_15867,N_15520);
or U16097 (N_16097,N_15901,N_15978);
nor U16098 (N_16098,N_15797,N_15927);
xor U16099 (N_16099,N_15905,N_15953);
xnor U16100 (N_16100,N_15961,N_15766);
nand U16101 (N_16101,N_15887,N_15811);
nor U16102 (N_16102,N_15620,N_15782);
nand U16103 (N_16103,N_15560,N_15517);
or U16104 (N_16104,N_15686,N_15502);
xor U16105 (N_16105,N_15986,N_15838);
nor U16106 (N_16106,N_15777,N_15920);
xor U16107 (N_16107,N_15915,N_15586);
nand U16108 (N_16108,N_15955,N_15850);
xor U16109 (N_16109,N_15510,N_15658);
or U16110 (N_16110,N_15839,N_15847);
and U16111 (N_16111,N_15868,N_15641);
or U16112 (N_16112,N_15600,N_15798);
xor U16113 (N_16113,N_15683,N_15533);
xnor U16114 (N_16114,N_15843,N_15523);
nand U16115 (N_16115,N_15626,N_15738);
nand U16116 (N_16116,N_15596,N_15895);
nor U16117 (N_16117,N_15879,N_15773);
and U16118 (N_16118,N_15914,N_15814);
nor U16119 (N_16119,N_15706,N_15644);
and U16120 (N_16120,N_15896,N_15562);
xnor U16121 (N_16121,N_15636,N_15545);
xnor U16122 (N_16122,N_15812,N_15912);
nor U16123 (N_16123,N_15977,N_15941);
nor U16124 (N_16124,N_15764,N_15679);
nor U16125 (N_16125,N_15627,N_15704);
and U16126 (N_16126,N_15531,N_15806);
or U16127 (N_16127,N_15625,N_15888);
or U16128 (N_16128,N_15975,N_15610);
or U16129 (N_16129,N_15650,N_15529);
xor U16130 (N_16130,N_15535,N_15886);
xnor U16131 (N_16131,N_15518,N_15909);
and U16132 (N_16132,N_15606,N_15576);
and U16133 (N_16133,N_15585,N_15591);
or U16134 (N_16134,N_15581,N_15715);
xnor U16135 (N_16135,N_15720,N_15751);
nand U16136 (N_16136,N_15956,N_15929);
or U16137 (N_16137,N_15859,N_15534);
or U16138 (N_16138,N_15783,N_15923);
and U16139 (N_16139,N_15701,N_15739);
nand U16140 (N_16140,N_15633,N_15530);
nor U16141 (N_16141,N_15660,N_15748);
nand U16142 (N_16142,N_15618,N_15860);
nand U16143 (N_16143,N_15864,N_15999);
xnor U16144 (N_16144,N_15578,N_15998);
nor U16145 (N_16145,N_15516,N_15937);
nor U16146 (N_16146,N_15703,N_15866);
xnor U16147 (N_16147,N_15786,N_15856);
and U16148 (N_16148,N_15883,N_15954);
nor U16149 (N_16149,N_15536,N_15781);
nor U16150 (N_16150,N_15553,N_15667);
nor U16151 (N_16151,N_15501,N_15846);
and U16152 (N_16152,N_15931,N_15995);
nor U16153 (N_16153,N_15890,N_15837);
xor U16154 (N_16154,N_15513,N_15841);
nor U16155 (N_16155,N_15984,N_15852);
and U16156 (N_16156,N_15730,N_15681);
nand U16157 (N_16157,N_15669,N_15943);
and U16158 (N_16158,N_15754,N_15648);
xnor U16159 (N_16159,N_15762,N_15547);
nor U16160 (N_16160,N_15962,N_15678);
xnor U16161 (N_16161,N_15632,N_15872);
nand U16162 (N_16162,N_15692,N_15784);
nand U16163 (N_16163,N_15870,N_15729);
nor U16164 (N_16164,N_15671,N_15590);
and U16165 (N_16165,N_15805,N_15769);
and U16166 (N_16166,N_15622,N_15528);
nor U16167 (N_16167,N_15880,N_15829);
and U16168 (N_16168,N_15505,N_15552);
xor U16169 (N_16169,N_15885,N_15716);
xnor U16170 (N_16170,N_15663,N_15538);
nand U16171 (N_16171,N_15794,N_15926);
or U16172 (N_16172,N_15574,N_15957);
or U16173 (N_16173,N_15611,N_15845);
or U16174 (N_16174,N_15568,N_15666);
and U16175 (N_16175,N_15532,N_15557);
nand U16176 (N_16176,N_15635,N_15742);
and U16177 (N_16177,N_15974,N_15788);
nor U16178 (N_16178,N_15747,N_15945);
nor U16179 (N_16179,N_15833,N_15983);
xnor U16180 (N_16180,N_15504,N_15944);
or U16181 (N_16181,N_15967,N_15617);
nand U16182 (N_16182,N_15907,N_15862);
nand U16183 (N_16183,N_15608,N_15699);
xor U16184 (N_16184,N_15891,N_15985);
xnor U16185 (N_16185,N_15573,N_15732);
nand U16186 (N_16186,N_15826,N_15950);
or U16187 (N_16187,N_15712,N_15698);
nand U16188 (N_16188,N_15563,N_15672);
and U16189 (N_16189,N_15791,N_15940);
nor U16190 (N_16190,N_15640,N_15541);
and U16191 (N_16191,N_15522,N_15849);
or U16192 (N_16192,N_15924,N_15908);
and U16193 (N_16193,N_15629,N_15934);
nor U16194 (N_16194,N_15994,N_15865);
nand U16195 (N_16195,N_15894,N_15965);
and U16196 (N_16196,N_15771,N_15804);
and U16197 (N_16197,N_15990,N_15761);
or U16198 (N_16198,N_15634,N_15539);
xor U16199 (N_16199,N_15981,N_15584);
xnor U16200 (N_16200,N_15737,N_15540);
nor U16201 (N_16201,N_15710,N_15809);
xnor U16202 (N_16202,N_15659,N_15795);
nand U16203 (N_16203,N_15851,N_15601);
nand U16204 (N_16204,N_15688,N_15726);
or U16205 (N_16205,N_15735,N_15844);
and U16206 (N_16206,N_15828,N_15827);
and U16207 (N_16207,N_15580,N_15948);
nor U16208 (N_16208,N_15605,N_15656);
nor U16209 (N_16209,N_15651,N_15951);
or U16210 (N_16210,N_15750,N_15684);
or U16211 (N_16211,N_15830,N_15546);
nand U16212 (N_16212,N_15691,N_15598);
nor U16213 (N_16213,N_15612,N_15554);
xor U16214 (N_16214,N_15577,N_15911);
and U16215 (N_16215,N_15946,N_15677);
nor U16216 (N_16216,N_15780,N_15718);
nor U16217 (N_16217,N_15674,N_15902);
xnor U16218 (N_16218,N_15740,N_15579);
nand U16219 (N_16219,N_15904,N_15507);
and U16220 (N_16220,N_15693,N_15933);
xnor U16221 (N_16221,N_15595,N_15878);
xnor U16222 (N_16222,N_15512,N_15899);
xor U16223 (N_16223,N_15645,N_15602);
xor U16224 (N_16224,N_15685,N_15952);
or U16225 (N_16225,N_15869,N_15728);
xor U16226 (N_16226,N_15796,N_15785);
nor U16227 (N_16227,N_15822,N_15724);
nor U16228 (N_16228,N_15676,N_15542);
and U16229 (N_16229,N_15647,N_15723);
and U16230 (N_16230,N_15884,N_15713);
or U16231 (N_16231,N_15727,N_15695);
and U16232 (N_16232,N_15558,N_15503);
or U16233 (N_16233,N_15938,N_15935);
nor U16234 (N_16234,N_15603,N_15514);
and U16235 (N_16235,N_15960,N_15696);
nor U16236 (N_16236,N_15753,N_15508);
nor U16237 (N_16237,N_15949,N_15630);
or U16238 (N_16238,N_15717,N_15840);
nor U16239 (N_16239,N_15646,N_15687);
nor U16240 (N_16240,N_15966,N_15793);
and U16241 (N_16241,N_15642,N_15969);
and U16242 (N_16242,N_15734,N_15768);
or U16243 (N_16243,N_15853,N_15968);
nor U16244 (N_16244,N_15593,N_15624);
xnor U16245 (N_16245,N_15544,N_15871);
nor U16246 (N_16246,N_15506,N_15892);
nand U16247 (N_16247,N_15939,N_15665);
nand U16248 (N_16248,N_15744,N_15756);
xnor U16249 (N_16249,N_15604,N_15525);
or U16250 (N_16250,N_15887,N_15572);
xnor U16251 (N_16251,N_15802,N_15749);
and U16252 (N_16252,N_15891,N_15731);
and U16253 (N_16253,N_15908,N_15552);
or U16254 (N_16254,N_15590,N_15686);
nand U16255 (N_16255,N_15665,N_15681);
or U16256 (N_16256,N_15787,N_15708);
and U16257 (N_16257,N_15881,N_15914);
nand U16258 (N_16258,N_15936,N_15937);
nand U16259 (N_16259,N_15788,N_15694);
xnor U16260 (N_16260,N_15650,N_15791);
xnor U16261 (N_16261,N_15801,N_15773);
nor U16262 (N_16262,N_15778,N_15889);
and U16263 (N_16263,N_15976,N_15999);
nor U16264 (N_16264,N_15877,N_15695);
xnor U16265 (N_16265,N_15881,N_15723);
and U16266 (N_16266,N_15613,N_15513);
xnor U16267 (N_16267,N_15517,N_15670);
or U16268 (N_16268,N_15705,N_15762);
xor U16269 (N_16269,N_15762,N_15837);
and U16270 (N_16270,N_15512,N_15750);
and U16271 (N_16271,N_15659,N_15775);
and U16272 (N_16272,N_15666,N_15601);
or U16273 (N_16273,N_15980,N_15566);
and U16274 (N_16274,N_15838,N_15741);
nor U16275 (N_16275,N_15632,N_15577);
xor U16276 (N_16276,N_15728,N_15642);
xor U16277 (N_16277,N_15734,N_15628);
xor U16278 (N_16278,N_15761,N_15845);
nand U16279 (N_16279,N_15907,N_15719);
xor U16280 (N_16280,N_15723,N_15756);
nor U16281 (N_16281,N_15860,N_15861);
nand U16282 (N_16282,N_15958,N_15787);
and U16283 (N_16283,N_15665,N_15784);
xor U16284 (N_16284,N_15708,N_15567);
and U16285 (N_16285,N_15819,N_15994);
and U16286 (N_16286,N_15538,N_15550);
nor U16287 (N_16287,N_15610,N_15925);
nor U16288 (N_16288,N_15983,N_15890);
nand U16289 (N_16289,N_15898,N_15578);
or U16290 (N_16290,N_15914,N_15616);
nand U16291 (N_16291,N_15821,N_15760);
or U16292 (N_16292,N_15968,N_15966);
or U16293 (N_16293,N_15968,N_15617);
nand U16294 (N_16294,N_15532,N_15648);
nand U16295 (N_16295,N_15959,N_15844);
nor U16296 (N_16296,N_15954,N_15923);
xor U16297 (N_16297,N_15863,N_15682);
and U16298 (N_16298,N_15939,N_15546);
or U16299 (N_16299,N_15541,N_15861);
nand U16300 (N_16300,N_15594,N_15870);
nor U16301 (N_16301,N_15753,N_15787);
and U16302 (N_16302,N_15707,N_15686);
or U16303 (N_16303,N_15969,N_15925);
and U16304 (N_16304,N_15859,N_15681);
and U16305 (N_16305,N_15867,N_15960);
and U16306 (N_16306,N_15512,N_15567);
xnor U16307 (N_16307,N_15634,N_15834);
or U16308 (N_16308,N_15655,N_15985);
xor U16309 (N_16309,N_15738,N_15504);
and U16310 (N_16310,N_15929,N_15654);
xor U16311 (N_16311,N_15724,N_15888);
or U16312 (N_16312,N_15674,N_15562);
nor U16313 (N_16313,N_15520,N_15572);
nor U16314 (N_16314,N_15674,N_15806);
nor U16315 (N_16315,N_15802,N_15518);
xor U16316 (N_16316,N_15656,N_15799);
nand U16317 (N_16317,N_15598,N_15546);
or U16318 (N_16318,N_15955,N_15936);
or U16319 (N_16319,N_15568,N_15708);
and U16320 (N_16320,N_15810,N_15534);
and U16321 (N_16321,N_15767,N_15954);
nand U16322 (N_16322,N_15788,N_15505);
nand U16323 (N_16323,N_15663,N_15912);
or U16324 (N_16324,N_15963,N_15641);
nand U16325 (N_16325,N_15816,N_15549);
xnor U16326 (N_16326,N_15650,N_15563);
xnor U16327 (N_16327,N_15564,N_15693);
xor U16328 (N_16328,N_15561,N_15956);
xor U16329 (N_16329,N_15943,N_15766);
nand U16330 (N_16330,N_15866,N_15628);
nand U16331 (N_16331,N_15940,N_15899);
or U16332 (N_16332,N_15515,N_15842);
nand U16333 (N_16333,N_15691,N_15704);
nand U16334 (N_16334,N_15883,N_15621);
and U16335 (N_16335,N_15556,N_15908);
xnor U16336 (N_16336,N_15580,N_15583);
and U16337 (N_16337,N_15527,N_15676);
nor U16338 (N_16338,N_15977,N_15522);
nor U16339 (N_16339,N_15912,N_15518);
nor U16340 (N_16340,N_15603,N_15866);
and U16341 (N_16341,N_15642,N_15841);
or U16342 (N_16342,N_15689,N_15507);
nand U16343 (N_16343,N_15962,N_15870);
nand U16344 (N_16344,N_15619,N_15975);
or U16345 (N_16345,N_15993,N_15914);
xnor U16346 (N_16346,N_15604,N_15745);
nand U16347 (N_16347,N_15509,N_15850);
nand U16348 (N_16348,N_15540,N_15883);
nor U16349 (N_16349,N_15718,N_15846);
xnor U16350 (N_16350,N_15772,N_15842);
nor U16351 (N_16351,N_15743,N_15611);
nor U16352 (N_16352,N_15646,N_15784);
nand U16353 (N_16353,N_15686,N_15605);
or U16354 (N_16354,N_15964,N_15516);
and U16355 (N_16355,N_15518,N_15946);
or U16356 (N_16356,N_15770,N_15905);
or U16357 (N_16357,N_15912,N_15641);
and U16358 (N_16358,N_15725,N_15871);
xnor U16359 (N_16359,N_15810,N_15942);
and U16360 (N_16360,N_15674,N_15822);
and U16361 (N_16361,N_15503,N_15999);
or U16362 (N_16362,N_15626,N_15741);
xor U16363 (N_16363,N_15589,N_15647);
xnor U16364 (N_16364,N_15951,N_15937);
nor U16365 (N_16365,N_15793,N_15944);
nand U16366 (N_16366,N_15802,N_15540);
nand U16367 (N_16367,N_15927,N_15621);
nand U16368 (N_16368,N_15536,N_15647);
or U16369 (N_16369,N_15786,N_15596);
xor U16370 (N_16370,N_15837,N_15726);
and U16371 (N_16371,N_15814,N_15727);
xor U16372 (N_16372,N_15893,N_15749);
xor U16373 (N_16373,N_15804,N_15727);
and U16374 (N_16374,N_15574,N_15861);
nand U16375 (N_16375,N_15588,N_15861);
or U16376 (N_16376,N_15567,N_15820);
nor U16377 (N_16377,N_15970,N_15593);
nor U16378 (N_16378,N_15878,N_15713);
and U16379 (N_16379,N_15928,N_15897);
xor U16380 (N_16380,N_15555,N_15623);
and U16381 (N_16381,N_15895,N_15829);
xor U16382 (N_16382,N_15547,N_15672);
or U16383 (N_16383,N_15580,N_15807);
xor U16384 (N_16384,N_15618,N_15895);
xnor U16385 (N_16385,N_15579,N_15586);
nor U16386 (N_16386,N_15876,N_15818);
and U16387 (N_16387,N_15949,N_15547);
or U16388 (N_16388,N_15740,N_15624);
nand U16389 (N_16389,N_15622,N_15830);
and U16390 (N_16390,N_15912,N_15525);
xnor U16391 (N_16391,N_15898,N_15691);
nor U16392 (N_16392,N_15909,N_15706);
and U16393 (N_16393,N_15955,N_15710);
and U16394 (N_16394,N_15515,N_15683);
or U16395 (N_16395,N_15871,N_15671);
or U16396 (N_16396,N_15504,N_15812);
xnor U16397 (N_16397,N_15845,N_15945);
xor U16398 (N_16398,N_15804,N_15908);
nor U16399 (N_16399,N_15997,N_15511);
and U16400 (N_16400,N_15832,N_15743);
xor U16401 (N_16401,N_15717,N_15943);
and U16402 (N_16402,N_15707,N_15808);
or U16403 (N_16403,N_15641,N_15815);
or U16404 (N_16404,N_15795,N_15744);
and U16405 (N_16405,N_15531,N_15891);
xor U16406 (N_16406,N_15516,N_15641);
or U16407 (N_16407,N_15832,N_15788);
nor U16408 (N_16408,N_15799,N_15956);
and U16409 (N_16409,N_15835,N_15599);
or U16410 (N_16410,N_15595,N_15894);
xnor U16411 (N_16411,N_15830,N_15905);
nand U16412 (N_16412,N_15731,N_15644);
and U16413 (N_16413,N_15779,N_15649);
nor U16414 (N_16414,N_15942,N_15642);
and U16415 (N_16415,N_15629,N_15639);
and U16416 (N_16416,N_15732,N_15689);
nand U16417 (N_16417,N_15970,N_15612);
or U16418 (N_16418,N_15983,N_15799);
and U16419 (N_16419,N_15979,N_15687);
and U16420 (N_16420,N_15789,N_15583);
nor U16421 (N_16421,N_15670,N_15980);
or U16422 (N_16422,N_15665,N_15868);
nand U16423 (N_16423,N_15701,N_15649);
nor U16424 (N_16424,N_15639,N_15741);
or U16425 (N_16425,N_15531,N_15745);
nor U16426 (N_16426,N_15666,N_15535);
nor U16427 (N_16427,N_15953,N_15605);
xor U16428 (N_16428,N_15717,N_15990);
xor U16429 (N_16429,N_15560,N_15708);
nor U16430 (N_16430,N_15579,N_15923);
xor U16431 (N_16431,N_15560,N_15908);
and U16432 (N_16432,N_15917,N_15524);
xor U16433 (N_16433,N_15928,N_15532);
nand U16434 (N_16434,N_15986,N_15672);
nor U16435 (N_16435,N_15867,N_15838);
or U16436 (N_16436,N_15973,N_15982);
nand U16437 (N_16437,N_15681,N_15722);
and U16438 (N_16438,N_15885,N_15687);
or U16439 (N_16439,N_15624,N_15698);
and U16440 (N_16440,N_15930,N_15788);
xnor U16441 (N_16441,N_15843,N_15705);
or U16442 (N_16442,N_15933,N_15664);
nand U16443 (N_16443,N_15575,N_15739);
nor U16444 (N_16444,N_15802,N_15531);
nand U16445 (N_16445,N_15993,N_15959);
nand U16446 (N_16446,N_15683,N_15789);
or U16447 (N_16447,N_15838,N_15784);
nand U16448 (N_16448,N_15760,N_15739);
and U16449 (N_16449,N_15533,N_15967);
nor U16450 (N_16450,N_15705,N_15545);
and U16451 (N_16451,N_15596,N_15699);
xor U16452 (N_16452,N_15692,N_15557);
and U16453 (N_16453,N_15942,N_15580);
xor U16454 (N_16454,N_15568,N_15624);
nor U16455 (N_16455,N_15764,N_15760);
and U16456 (N_16456,N_15564,N_15530);
or U16457 (N_16457,N_15767,N_15508);
xnor U16458 (N_16458,N_15800,N_15527);
nor U16459 (N_16459,N_15542,N_15837);
and U16460 (N_16460,N_15819,N_15719);
nand U16461 (N_16461,N_15866,N_15802);
and U16462 (N_16462,N_15922,N_15982);
nand U16463 (N_16463,N_15766,N_15688);
nor U16464 (N_16464,N_15712,N_15726);
xor U16465 (N_16465,N_15819,N_15972);
or U16466 (N_16466,N_15695,N_15607);
nand U16467 (N_16467,N_15597,N_15841);
xnor U16468 (N_16468,N_15875,N_15615);
or U16469 (N_16469,N_15845,N_15770);
nand U16470 (N_16470,N_15885,N_15962);
xor U16471 (N_16471,N_15691,N_15674);
nand U16472 (N_16472,N_15937,N_15927);
and U16473 (N_16473,N_15694,N_15578);
xor U16474 (N_16474,N_15649,N_15751);
and U16475 (N_16475,N_15704,N_15736);
nor U16476 (N_16476,N_15886,N_15964);
or U16477 (N_16477,N_15592,N_15938);
xnor U16478 (N_16478,N_15933,N_15927);
and U16479 (N_16479,N_15982,N_15529);
xnor U16480 (N_16480,N_15954,N_15811);
and U16481 (N_16481,N_15620,N_15944);
nand U16482 (N_16482,N_15572,N_15842);
xor U16483 (N_16483,N_15788,N_15562);
xnor U16484 (N_16484,N_15767,N_15622);
xor U16485 (N_16485,N_15510,N_15611);
nand U16486 (N_16486,N_15953,N_15944);
nor U16487 (N_16487,N_15624,N_15706);
xnor U16488 (N_16488,N_15802,N_15829);
or U16489 (N_16489,N_15799,N_15751);
and U16490 (N_16490,N_15829,N_15555);
or U16491 (N_16491,N_15637,N_15735);
xnor U16492 (N_16492,N_15614,N_15542);
xnor U16493 (N_16493,N_15745,N_15797);
nand U16494 (N_16494,N_15876,N_15670);
nor U16495 (N_16495,N_15994,N_15987);
nor U16496 (N_16496,N_15664,N_15511);
and U16497 (N_16497,N_15719,N_15722);
xor U16498 (N_16498,N_15683,N_15687);
nand U16499 (N_16499,N_15797,N_15564);
nor U16500 (N_16500,N_16182,N_16360);
and U16501 (N_16501,N_16227,N_16122);
nand U16502 (N_16502,N_16251,N_16430);
nor U16503 (N_16503,N_16133,N_16248);
nor U16504 (N_16504,N_16381,N_16448);
xnor U16505 (N_16505,N_16282,N_16070);
or U16506 (N_16506,N_16319,N_16088);
nand U16507 (N_16507,N_16472,N_16329);
nor U16508 (N_16508,N_16264,N_16173);
or U16509 (N_16509,N_16275,N_16418);
nand U16510 (N_16510,N_16034,N_16243);
xor U16511 (N_16511,N_16374,N_16307);
and U16512 (N_16512,N_16195,N_16454);
nor U16513 (N_16513,N_16345,N_16179);
nor U16514 (N_16514,N_16138,N_16372);
nor U16515 (N_16515,N_16285,N_16224);
and U16516 (N_16516,N_16438,N_16115);
or U16517 (N_16517,N_16040,N_16229);
and U16518 (N_16518,N_16223,N_16164);
and U16519 (N_16519,N_16038,N_16333);
nand U16520 (N_16520,N_16490,N_16068);
xnor U16521 (N_16521,N_16405,N_16361);
xnor U16522 (N_16522,N_16254,N_16209);
nor U16523 (N_16523,N_16242,N_16047);
nand U16524 (N_16524,N_16002,N_16450);
xor U16525 (N_16525,N_16163,N_16286);
nor U16526 (N_16526,N_16222,N_16210);
nor U16527 (N_16527,N_16476,N_16279);
nor U16528 (N_16528,N_16150,N_16011);
and U16529 (N_16529,N_16260,N_16004);
and U16530 (N_16530,N_16406,N_16069);
nor U16531 (N_16531,N_16484,N_16300);
nand U16532 (N_16532,N_16111,N_16441);
xor U16533 (N_16533,N_16323,N_16487);
or U16534 (N_16534,N_16082,N_16241);
and U16535 (N_16535,N_16114,N_16410);
or U16536 (N_16536,N_16477,N_16013);
nand U16537 (N_16537,N_16053,N_16439);
nor U16538 (N_16538,N_16431,N_16186);
xor U16539 (N_16539,N_16095,N_16027);
nand U16540 (N_16540,N_16193,N_16204);
nor U16541 (N_16541,N_16428,N_16412);
or U16542 (N_16542,N_16312,N_16196);
nor U16543 (N_16543,N_16464,N_16245);
nor U16544 (N_16544,N_16432,N_16315);
xor U16545 (N_16545,N_16335,N_16313);
and U16546 (N_16546,N_16256,N_16469);
and U16547 (N_16547,N_16000,N_16126);
and U16548 (N_16548,N_16453,N_16375);
nand U16549 (N_16549,N_16420,N_16259);
nor U16550 (N_16550,N_16263,N_16029);
xnor U16551 (N_16551,N_16250,N_16455);
xor U16552 (N_16552,N_16211,N_16281);
and U16553 (N_16553,N_16155,N_16079);
or U16554 (N_16554,N_16178,N_16142);
nor U16555 (N_16555,N_16239,N_16203);
nor U16556 (N_16556,N_16192,N_16035);
and U16557 (N_16557,N_16143,N_16039);
nand U16558 (N_16558,N_16328,N_16347);
nand U16559 (N_16559,N_16475,N_16368);
and U16560 (N_16560,N_16171,N_16465);
xnor U16561 (N_16561,N_16378,N_16495);
nor U16562 (N_16562,N_16184,N_16308);
and U16563 (N_16563,N_16467,N_16444);
xnor U16564 (N_16564,N_16409,N_16459);
and U16565 (N_16565,N_16385,N_16481);
nand U16566 (N_16566,N_16370,N_16299);
or U16567 (N_16567,N_16435,N_16161);
nand U16568 (N_16568,N_16205,N_16208);
nor U16569 (N_16569,N_16283,N_16147);
or U16570 (N_16570,N_16080,N_16094);
nand U16571 (N_16571,N_16221,N_16235);
nor U16572 (N_16572,N_16261,N_16181);
or U16573 (N_16573,N_16197,N_16064);
and U16574 (N_16574,N_16072,N_16436);
nor U16575 (N_16575,N_16493,N_16124);
and U16576 (N_16576,N_16343,N_16295);
nand U16577 (N_16577,N_16103,N_16445);
xor U16578 (N_16578,N_16463,N_16189);
and U16579 (N_16579,N_16066,N_16451);
and U16580 (N_16580,N_16429,N_16137);
or U16581 (N_16581,N_16046,N_16305);
and U16582 (N_16582,N_16352,N_16353);
nor U16583 (N_16583,N_16398,N_16019);
nand U16584 (N_16584,N_16212,N_16015);
nor U16585 (N_16585,N_16177,N_16421);
nor U16586 (N_16586,N_16234,N_16311);
and U16587 (N_16587,N_16157,N_16321);
or U16588 (N_16588,N_16437,N_16231);
nand U16589 (N_16589,N_16310,N_16393);
nor U16590 (N_16590,N_16244,N_16379);
nand U16591 (N_16591,N_16036,N_16434);
nor U16592 (N_16592,N_16402,N_16257);
xnor U16593 (N_16593,N_16292,N_16032);
and U16594 (N_16594,N_16166,N_16277);
and U16595 (N_16595,N_16109,N_16258);
xnor U16596 (N_16596,N_16492,N_16377);
nand U16597 (N_16597,N_16014,N_16020);
or U16598 (N_16598,N_16373,N_16468);
and U16599 (N_16599,N_16121,N_16217);
nor U16600 (N_16600,N_16132,N_16376);
and U16601 (N_16601,N_16201,N_16025);
or U16602 (N_16602,N_16386,N_16494);
or U16603 (N_16603,N_16271,N_16059);
or U16604 (N_16604,N_16380,N_16425);
nor U16605 (N_16605,N_16449,N_16165);
and U16606 (N_16606,N_16306,N_16270);
and U16607 (N_16607,N_16022,N_16233);
nor U16608 (N_16608,N_16348,N_16424);
nand U16609 (N_16609,N_16188,N_16466);
nor U16610 (N_16610,N_16098,N_16317);
and U16611 (N_16611,N_16009,N_16175);
and U16612 (N_16612,N_16216,N_16006);
or U16613 (N_16613,N_16062,N_16156);
nor U16614 (N_16614,N_16470,N_16099);
nor U16615 (N_16615,N_16028,N_16240);
nor U16616 (N_16616,N_16169,N_16461);
or U16617 (N_16617,N_16400,N_16276);
nor U16618 (N_16618,N_16303,N_16010);
or U16619 (N_16619,N_16050,N_16289);
xnor U16620 (N_16620,N_16489,N_16273);
xnor U16621 (N_16621,N_16026,N_16265);
nand U16622 (N_16622,N_16052,N_16226);
nor U16623 (N_16623,N_16391,N_16005);
xor U16624 (N_16624,N_16351,N_16284);
nand U16625 (N_16625,N_16012,N_16093);
and U16626 (N_16626,N_16364,N_16118);
or U16627 (N_16627,N_16214,N_16411);
or U16628 (N_16628,N_16366,N_16389);
and U16629 (N_16629,N_16344,N_16051);
nor U16630 (N_16630,N_16322,N_16457);
nor U16631 (N_16631,N_16349,N_16120);
nand U16632 (N_16632,N_16443,N_16037);
or U16633 (N_16633,N_16117,N_16061);
and U16634 (N_16634,N_16479,N_16304);
xnor U16635 (N_16635,N_16294,N_16136);
nand U16636 (N_16636,N_16365,N_16355);
nor U16637 (N_16637,N_16255,N_16269);
nand U16638 (N_16638,N_16357,N_16225);
or U16639 (N_16639,N_16408,N_16413);
and U16640 (N_16640,N_16427,N_16054);
and U16641 (N_16641,N_16041,N_16280);
xnor U16642 (N_16642,N_16316,N_16085);
or U16643 (N_16643,N_16397,N_16102);
xor U16644 (N_16644,N_16392,N_16452);
nand U16645 (N_16645,N_16268,N_16339);
nand U16646 (N_16646,N_16314,N_16262);
nor U16647 (N_16647,N_16350,N_16325);
and U16648 (N_16648,N_16087,N_16309);
nand U16649 (N_16649,N_16119,N_16185);
nor U16650 (N_16650,N_16458,N_16423);
nand U16651 (N_16651,N_16499,N_16297);
or U16652 (N_16652,N_16340,N_16151);
or U16653 (N_16653,N_16125,N_16191);
nand U16654 (N_16654,N_16030,N_16354);
nor U16655 (N_16655,N_16123,N_16154);
and U16656 (N_16656,N_16100,N_16485);
or U16657 (N_16657,N_16336,N_16198);
nor U16658 (N_16658,N_16176,N_16332);
and U16659 (N_16659,N_16130,N_16358);
or U16660 (N_16660,N_16440,N_16482);
or U16661 (N_16661,N_16016,N_16327);
nor U16662 (N_16662,N_16042,N_16288);
nand U16663 (N_16663,N_16091,N_16159);
nand U16664 (N_16664,N_16394,N_16077);
nand U16665 (N_16665,N_16152,N_16302);
or U16666 (N_16666,N_16416,N_16456);
and U16667 (N_16667,N_16384,N_16168);
nand U16668 (N_16668,N_16135,N_16274);
and U16669 (N_16669,N_16346,N_16110);
or U16670 (N_16670,N_16447,N_16287);
nand U16671 (N_16671,N_16218,N_16096);
and U16672 (N_16672,N_16442,N_16215);
nand U16673 (N_16673,N_16049,N_16362);
nand U16674 (N_16674,N_16141,N_16158);
and U16675 (N_16675,N_16160,N_16057);
or U16676 (N_16676,N_16063,N_16106);
and U16677 (N_16677,N_16101,N_16140);
nand U16678 (N_16678,N_16206,N_16090);
nand U16679 (N_16679,N_16474,N_16471);
nand U16680 (N_16680,N_16324,N_16200);
and U16681 (N_16681,N_16105,N_16334);
nand U16682 (N_16682,N_16071,N_16407);
nand U16683 (N_16683,N_16056,N_16480);
nor U16684 (N_16684,N_16033,N_16075);
xnor U16685 (N_16685,N_16228,N_16084);
nand U16686 (N_16686,N_16083,N_16395);
nor U16687 (N_16687,N_16170,N_16266);
and U16688 (N_16688,N_16048,N_16067);
nor U16689 (N_16689,N_16043,N_16017);
nor U16690 (N_16690,N_16296,N_16318);
xor U16691 (N_16691,N_16001,N_16247);
xnor U16692 (N_16692,N_16237,N_16253);
nand U16693 (N_16693,N_16387,N_16183);
and U16694 (N_16694,N_16399,N_16278);
xor U16695 (N_16695,N_16076,N_16008);
xor U16696 (N_16696,N_16129,N_16446);
nor U16697 (N_16697,N_16162,N_16403);
nand U16698 (N_16698,N_16473,N_16496);
xor U16699 (N_16699,N_16415,N_16326);
nor U16700 (N_16700,N_16153,N_16107);
nand U16701 (N_16701,N_16128,N_16127);
nor U16702 (N_16702,N_16003,N_16272);
or U16703 (N_16703,N_16498,N_16422);
xnor U16704 (N_16704,N_16230,N_16058);
nor U16705 (N_16705,N_16097,N_16116);
xor U16706 (N_16706,N_16220,N_16383);
or U16707 (N_16707,N_16460,N_16359);
xnor U16708 (N_16708,N_16060,N_16246);
nand U16709 (N_16709,N_16131,N_16139);
and U16710 (N_16710,N_16108,N_16024);
xor U16711 (N_16711,N_16190,N_16187);
xnor U16712 (N_16712,N_16018,N_16007);
nor U16713 (N_16713,N_16371,N_16031);
nand U16714 (N_16714,N_16369,N_16236);
nand U16715 (N_16715,N_16074,N_16044);
and U16716 (N_16716,N_16396,N_16199);
or U16717 (N_16717,N_16382,N_16172);
or U16718 (N_16718,N_16113,N_16149);
nand U16719 (N_16719,N_16073,N_16104);
and U16720 (N_16720,N_16249,N_16144);
nand U16721 (N_16721,N_16419,N_16367);
xor U16722 (N_16722,N_16078,N_16426);
or U16723 (N_16723,N_16267,N_16338);
xnor U16724 (N_16724,N_16342,N_16433);
nand U16725 (N_16725,N_16194,N_16337);
nand U16726 (N_16726,N_16390,N_16401);
nor U16727 (N_16727,N_16112,N_16356);
and U16728 (N_16728,N_16086,N_16483);
and U16729 (N_16729,N_16167,N_16145);
nor U16730 (N_16730,N_16298,N_16331);
nand U16731 (N_16731,N_16238,N_16363);
nor U16732 (N_16732,N_16301,N_16486);
xnor U16733 (N_16733,N_16081,N_16488);
nand U16734 (N_16734,N_16092,N_16293);
nand U16735 (N_16735,N_16089,N_16320);
xnor U16736 (N_16736,N_16219,N_16388);
or U16737 (N_16737,N_16180,N_16045);
nand U16738 (N_16738,N_16213,N_16330);
or U16739 (N_16739,N_16404,N_16146);
xor U16740 (N_16740,N_16055,N_16341);
and U16741 (N_16741,N_16414,N_16291);
nor U16742 (N_16742,N_16207,N_16023);
and U16743 (N_16743,N_16065,N_16148);
nor U16744 (N_16744,N_16462,N_16290);
xnor U16745 (N_16745,N_16417,N_16174);
or U16746 (N_16746,N_16497,N_16232);
nor U16747 (N_16747,N_16134,N_16021);
xor U16748 (N_16748,N_16491,N_16202);
nand U16749 (N_16749,N_16252,N_16478);
xnor U16750 (N_16750,N_16085,N_16267);
xnor U16751 (N_16751,N_16496,N_16146);
nor U16752 (N_16752,N_16116,N_16138);
nor U16753 (N_16753,N_16384,N_16434);
or U16754 (N_16754,N_16392,N_16398);
nor U16755 (N_16755,N_16418,N_16056);
or U16756 (N_16756,N_16003,N_16346);
or U16757 (N_16757,N_16164,N_16411);
nand U16758 (N_16758,N_16364,N_16425);
or U16759 (N_16759,N_16076,N_16446);
nand U16760 (N_16760,N_16346,N_16314);
or U16761 (N_16761,N_16252,N_16332);
and U16762 (N_16762,N_16391,N_16372);
or U16763 (N_16763,N_16106,N_16485);
nand U16764 (N_16764,N_16046,N_16281);
nor U16765 (N_16765,N_16466,N_16080);
or U16766 (N_16766,N_16212,N_16030);
and U16767 (N_16767,N_16093,N_16404);
and U16768 (N_16768,N_16216,N_16309);
nand U16769 (N_16769,N_16339,N_16078);
nor U16770 (N_16770,N_16295,N_16182);
nand U16771 (N_16771,N_16032,N_16127);
nor U16772 (N_16772,N_16436,N_16258);
nand U16773 (N_16773,N_16088,N_16052);
nand U16774 (N_16774,N_16207,N_16376);
xnor U16775 (N_16775,N_16400,N_16076);
nand U16776 (N_16776,N_16046,N_16082);
xor U16777 (N_16777,N_16020,N_16249);
nand U16778 (N_16778,N_16344,N_16249);
nor U16779 (N_16779,N_16015,N_16250);
xor U16780 (N_16780,N_16230,N_16120);
nand U16781 (N_16781,N_16145,N_16328);
or U16782 (N_16782,N_16093,N_16224);
and U16783 (N_16783,N_16452,N_16275);
nand U16784 (N_16784,N_16386,N_16222);
and U16785 (N_16785,N_16173,N_16101);
and U16786 (N_16786,N_16071,N_16078);
nor U16787 (N_16787,N_16382,N_16318);
or U16788 (N_16788,N_16060,N_16291);
nor U16789 (N_16789,N_16171,N_16065);
nand U16790 (N_16790,N_16341,N_16402);
xnor U16791 (N_16791,N_16038,N_16335);
nand U16792 (N_16792,N_16276,N_16151);
xor U16793 (N_16793,N_16012,N_16241);
and U16794 (N_16794,N_16048,N_16045);
nor U16795 (N_16795,N_16464,N_16158);
or U16796 (N_16796,N_16251,N_16468);
nor U16797 (N_16797,N_16237,N_16138);
nand U16798 (N_16798,N_16074,N_16355);
or U16799 (N_16799,N_16466,N_16067);
nor U16800 (N_16800,N_16108,N_16386);
and U16801 (N_16801,N_16051,N_16442);
xor U16802 (N_16802,N_16460,N_16447);
nor U16803 (N_16803,N_16096,N_16125);
or U16804 (N_16804,N_16370,N_16490);
and U16805 (N_16805,N_16356,N_16188);
nor U16806 (N_16806,N_16219,N_16217);
and U16807 (N_16807,N_16118,N_16480);
nand U16808 (N_16808,N_16316,N_16315);
nand U16809 (N_16809,N_16399,N_16467);
xor U16810 (N_16810,N_16237,N_16325);
and U16811 (N_16811,N_16461,N_16121);
xor U16812 (N_16812,N_16020,N_16152);
xnor U16813 (N_16813,N_16224,N_16328);
xnor U16814 (N_16814,N_16108,N_16391);
xor U16815 (N_16815,N_16184,N_16229);
nand U16816 (N_16816,N_16270,N_16258);
or U16817 (N_16817,N_16313,N_16132);
or U16818 (N_16818,N_16354,N_16107);
and U16819 (N_16819,N_16003,N_16015);
nand U16820 (N_16820,N_16250,N_16296);
nand U16821 (N_16821,N_16027,N_16498);
xor U16822 (N_16822,N_16436,N_16182);
nor U16823 (N_16823,N_16401,N_16472);
nor U16824 (N_16824,N_16304,N_16131);
nand U16825 (N_16825,N_16062,N_16004);
nor U16826 (N_16826,N_16398,N_16298);
nand U16827 (N_16827,N_16006,N_16429);
nor U16828 (N_16828,N_16229,N_16422);
or U16829 (N_16829,N_16464,N_16021);
xnor U16830 (N_16830,N_16116,N_16411);
or U16831 (N_16831,N_16355,N_16433);
or U16832 (N_16832,N_16133,N_16138);
xnor U16833 (N_16833,N_16065,N_16361);
xnor U16834 (N_16834,N_16170,N_16389);
or U16835 (N_16835,N_16248,N_16057);
xnor U16836 (N_16836,N_16434,N_16489);
xor U16837 (N_16837,N_16352,N_16407);
or U16838 (N_16838,N_16134,N_16456);
and U16839 (N_16839,N_16087,N_16196);
xnor U16840 (N_16840,N_16133,N_16168);
nor U16841 (N_16841,N_16172,N_16312);
and U16842 (N_16842,N_16311,N_16295);
or U16843 (N_16843,N_16387,N_16047);
nor U16844 (N_16844,N_16132,N_16202);
xor U16845 (N_16845,N_16426,N_16229);
nor U16846 (N_16846,N_16097,N_16328);
nor U16847 (N_16847,N_16082,N_16014);
nand U16848 (N_16848,N_16022,N_16371);
nor U16849 (N_16849,N_16433,N_16260);
and U16850 (N_16850,N_16325,N_16475);
or U16851 (N_16851,N_16116,N_16142);
or U16852 (N_16852,N_16027,N_16399);
xnor U16853 (N_16853,N_16434,N_16300);
or U16854 (N_16854,N_16180,N_16303);
and U16855 (N_16855,N_16015,N_16127);
nand U16856 (N_16856,N_16479,N_16262);
or U16857 (N_16857,N_16015,N_16387);
and U16858 (N_16858,N_16223,N_16043);
or U16859 (N_16859,N_16432,N_16324);
or U16860 (N_16860,N_16253,N_16013);
xnor U16861 (N_16861,N_16041,N_16338);
and U16862 (N_16862,N_16163,N_16362);
nand U16863 (N_16863,N_16144,N_16167);
nor U16864 (N_16864,N_16441,N_16498);
and U16865 (N_16865,N_16284,N_16337);
xor U16866 (N_16866,N_16088,N_16318);
nor U16867 (N_16867,N_16151,N_16014);
nor U16868 (N_16868,N_16396,N_16245);
xor U16869 (N_16869,N_16022,N_16204);
xnor U16870 (N_16870,N_16239,N_16305);
xnor U16871 (N_16871,N_16447,N_16331);
and U16872 (N_16872,N_16151,N_16071);
nor U16873 (N_16873,N_16313,N_16038);
nor U16874 (N_16874,N_16475,N_16088);
xor U16875 (N_16875,N_16459,N_16045);
nand U16876 (N_16876,N_16062,N_16224);
and U16877 (N_16877,N_16477,N_16057);
nand U16878 (N_16878,N_16294,N_16327);
nor U16879 (N_16879,N_16397,N_16248);
xor U16880 (N_16880,N_16310,N_16051);
nor U16881 (N_16881,N_16369,N_16160);
and U16882 (N_16882,N_16132,N_16330);
nand U16883 (N_16883,N_16446,N_16046);
nand U16884 (N_16884,N_16151,N_16108);
xnor U16885 (N_16885,N_16018,N_16099);
and U16886 (N_16886,N_16182,N_16310);
or U16887 (N_16887,N_16147,N_16148);
nor U16888 (N_16888,N_16254,N_16260);
nand U16889 (N_16889,N_16309,N_16080);
xnor U16890 (N_16890,N_16307,N_16401);
nand U16891 (N_16891,N_16484,N_16102);
nor U16892 (N_16892,N_16376,N_16499);
and U16893 (N_16893,N_16289,N_16114);
nand U16894 (N_16894,N_16080,N_16197);
and U16895 (N_16895,N_16182,N_16409);
nor U16896 (N_16896,N_16155,N_16385);
xnor U16897 (N_16897,N_16394,N_16126);
xnor U16898 (N_16898,N_16250,N_16343);
and U16899 (N_16899,N_16395,N_16175);
nor U16900 (N_16900,N_16251,N_16189);
xor U16901 (N_16901,N_16322,N_16454);
nor U16902 (N_16902,N_16414,N_16403);
or U16903 (N_16903,N_16203,N_16000);
or U16904 (N_16904,N_16350,N_16265);
xnor U16905 (N_16905,N_16133,N_16435);
xor U16906 (N_16906,N_16383,N_16264);
nand U16907 (N_16907,N_16163,N_16224);
nand U16908 (N_16908,N_16187,N_16178);
or U16909 (N_16909,N_16012,N_16046);
nand U16910 (N_16910,N_16143,N_16078);
nor U16911 (N_16911,N_16008,N_16454);
nor U16912 (N_16912,N_16429,N_16480);
nor U16913 (N_16913,N_16255,N_16027);
nor U16914 (N_16914,N_16169,N_16368);
nand U16915 (N_16915,N_16336,N_16382);
nor U16916 (N_16916,N_16235,N_16188);
nor U16917 (N_16917,N_16229,N_16161);
and U16918 (N_16918,N_16010,N_16285);
nand U16919 (N_16919,N_16318,N_16070);
xor U16920 (N_16920,N_16000,N_16263);
nor U16921 (N_16921,N_16231,N_16477);
or U16922 (N_16922,N_16371,N_16279);
nor U16923 (N_16923,N_16036,N_16381);
xor U16924 (N_16924,N_16442,N_16267);
nor U16925 (N_16925,N_16158,N_16100);
and U16926 (N_16926,N_16127,N_16205);
nand U16927 (N_16927,N_16395,N_16065);
nand U16928 (N_16928,N_16174,N_16410);
and U16929 (N_16929,N_16471,N_16100);
or U16930 (N_16930,N_16359,N_16241);
nor U16931 (N_16931,N_16404,N_16354);
or U16932 (N_16932,N_16366,N_16030);
or U16933 (N_16933,N_16061,N_16049);
nor U16934 (N_16934,N_16217,N_16287);
nand U16935 (N_16935,N_16216,N_16478);
or U16936 (N_16936,N_16139,N_16065);
nor U16937 (N_16937,N_16386,N_16215);
nor U16938 (N_16938,N_16073,N_16148);
or U16939 (N_16939,N_16110,N_16212);
and U16940 (N_16940,N_16490,N_16092);
or U16941 (N_16941,N_16252,N_16108);
xnor U16942 (N_16942,N_16481,N_16014);
nand U16943 (N_16943,N_16450,N_16369);
or U16944 (N_16944,N_16407,N_16051);
and U16945 (N_16945,N_16150,N_16087);
and U16946 (N_16946,N_16361,N_16180);
or U16947 (N_16947,N_16208,N_16474);
and U16948 (N_16948,N_16252,N_16033);
xor U16949 (N_16949,N_16249,N_16254);
xnor U16950 (N_16950,N_16055,N_16017);
xor U16951 (N_16951,N_16340,N_16493);
xnor U16952 (N_16952,N_16390,N_16250);
nand U16953 (N_16953,N_16384,N_16466);
or U16954 (N_16954,N_16167,N_16138);
nor U16955 (N_16955,N_16423,N_16465);
nand U16956 (N_16956,N_16298,N_16363);
and U16957 (N_16957,N_16027,N_16489);
nor U16958 (N_16958,N_16206,N_16305);
or U16959 (N_16959,N_16366,N_16231);
or U16960 (N_16960,N_16226,N_16085);
nor U16961 (N_16961,N_16426,N_16135);
and U16962 (N_16962,N_16411,N_16402);
or U16963 (N_16963,N_16338,N_16142);
and U16964 (N_16964,N_16027,N_16104);
nor U16965 (N_16965,N_16096,N_16415);
nand U16966 (N_16966,N_16194,N_16015);
xor U16967 (N_16967,N_16394,N_16010);
xor U16968 (N_16968,N_16096,N_16216);
nor U16969 (N_16969,N_16099,N_16060);
nor U16970 (N_16970,N_16424,N_16016);
nand U16971 (N_16971,N_16361,N_16232);
nand U16972 (N_16972,N_16139,N_16384);
or U16973 (N_16973,N_16270,N_16218);
nand U16974 (N_16974,N_16094,N_16498);
and U16975 (N_16975,N_16285,N_16051);
or U16976 (N_16976,N_16318,N_16434);
or U16977 (N_16977,N_16319,N_16229);
nand U16978 (N_16978,N_16384,N_16203);
nand U16979 (N_16979,N_16218,N_16138);
nor U16980 (N_16980,N_16424,N_16061);
or U16981 (N_16981,N_16437,N_16188);
xor U16982 (N_16982,N_16379,N_16320);
nand U16983 (N_16983,N_16362,N_16323);
nor U16984 (N_16984,N_16019,N_16430);
and U16985 (N_16985,N_16457,N_16336);
nand U16986 (N_16986,N_16207,N_16465);
and U16987 (N_16987,N_16475,N_16149);
nor U16988 (N_16988,N_16438,N_16002);
and U16989 (N_16989,N_16275,N_16186);
nand U16990 (N_16990,N_16451,N_16419);
nand U16991 (N_16991,N_16274,N_16464);
xnor U16992 (N_16992,N_16409,N_16002);
xor U16993 (N_16993,N_16292,N_16280);
or U16994 (N_16994,N_16159,N_16064);
nor U16995 (N_16995,N_16092,N_16190);
nor U16996 (N_16996,N_16029,N_16490);
nor U16997 (N_16997,N_16392,N_16457);
nor U16998 (N_16998,N_16460,N_16324);
xor U16999 (N_16999,N_16490,N_16062);
or U17000 (N_17000,N_16832,N_16673);
or U17001 (N_17001,N_16845,N_16955);
or U17002 (N_17002,N_16609,N_16577);
or U17003 (N_17003,N_16793,N_16707);
or U17004 (N_17004,N_16555,N_16620);
nor U17005 (N_17005,N_16676,N_16571);
and U17006 (N_17006,N_16970,N_16792);
and U17007 (N_17007,N_16783,N_16551);
xnor U17008 (N_17008,N_16935,N_16947);
nand U17009 (N_17009,N_16627,N_16718);
xor U17010 (N_17010,N_16769,N_16693);
and U17011 (N_17011,N_16597,N_16547);
nand U17012 (N_17012,N_16573,N_16840);
and U17013 (N_17013,N_16869,N_16533);
and U17014 (N_17014,N_16923,N_16613);
xor U17015 (N_17015,N_16595,N_16511);
or U17016 (N_17016,N_16959,N_16744);
nor U17017 (N_17017,N_16558,N_16716);
and U17018 (N_17018,N_16748,N_16619);
or U17019 (N_17019,N_16807,N_16733);
xnor U17020 (N_17020,N_16683,N_16844);
and U17021 (N_17021,N_16896,N_16757);
nand U17022 (N_17022,N_16870,N_16981);
or U17023 (N_17023,N_16696,N_16752);
and U17024 (N_17024,N_16580,N_16822);
and U17025 (N_17025,N_16809,N_16552);
nor U17026 (N_17026,N_16690,N_16908);
nor U17027 (N_17027,N_16904,N_16637);
nor U17028 (N_17028,N_16501,N_16841);
xnor U17029 (N_17029,N_16785,N_16991);
nor U17030 (N_17030,N_16916,N_16529);
nand U17031 (N_17031,N_16817,N_16521);
nand U17032 (N_17032,N_16838,N_16852);
nor U17033 (N_17033,N_16761,N_16576);
nand U17034 (N_17034,N_16814,N_16711);
or U17035 (N_17035,N_16585,N_16980);
or U17036 (N_17036,N_16952,N_16650);
or U17037 (N_17037,N_16633,N_16999);
nor U17038 (N_17038,N_16868,N_16765);
nor U17039 (N_17039,N_16767,N_16941);
or U17040 (N_17040,N_16678,N_16588);
nand U17041 (N_17041,N_16608,N_16988);
xor U17042 (N_17042,N_16976,N_16641);
or U17043 (N_17043,N_16928,N_16975);
nand U17044 (N_17044,N_16973,N_16788);
nand U17045 (N_17045,N_16979,N_16758);
and U17046 (N_17046,N_16601,N_16879);
or U17047 (N_17047,N_16987,N_16557);
and U17048 (N_17048,N_16566,N_16517);
nand U17049 (N_17049,N_16962,N_16539);
or U17050 (N_17050,N_16631,N_16944);
or U17051 (N_17051,N_16741,N_16713);
or U17052 (N_17052,N_16874,N_16569);
xor U17053 (N_17053,N_16885,N_16871);
nor U17054 (N_17054,N_16554,N_16528);
nand U17055 (N_17055,N_16544,N_16684);
nor U17056 (N_17056,N_16836,N_16509);
xnor U17057 (N_17057,N_16724,N_16854);
and U17058 (N_17058,N_16961,N_16968);
nand U17059 (N_17059,N_16589,N_16815);
and U17060 (N_17060,N_16727,N_16930);
and U17061 (N_17061,N_16773,N_16903);
nor U17062 (N_17062,N_16634,N_16686);
and U17063 (N_17063,N_16656,N_16820);
nand U17064 (N_17064,N_16695,N_16992);
nand U17065 (N_17065,N_16680,N_16804);
or U17066 (N_17066,N_16594,N_16969);
nand U17067 (N_17067,N_16786,N_16519);
or U17068 (N_17068,N_16805,N_16772);
or U17069 (N_17069,N_16721,N_16787);
or U17070 (N_17070,N_16742,N_16892);
nor U17071 (N_17071,N_16922,N_16636);
nand U17072 (N_17072,N_16598,N_16685);
or U17073 (N_17073,N_16500,N_16993);
and U17074 (N_17074,N_16888,N_16645);
or U17075 (N_17075,N_16689,N_16971);
or U17076 (N_17076,N_16704,N_16654);
and U17077 (N_17077,N_16965,N_16910);
nor U17078 (N_17078,N_16556,N_16953);
and U17079 (N_17079,N_16861,N_16801);
or U17080 (N_17080,N_16644,N_16775);
xor U17081 (N_17081,N_16766,N_16846);
xor U17082 (N_17082,N_16682,N_16812);
or U17083 (N_17083,N_16790,N_16729);
and U17084 (N_17084,N_16702,N_16628);
xnor U17085 (N_17085,N_16894,N_16646);
and U17086 (N_17086,N_16675,N_16966);
and U17087 (N_17087,N_16756,N_16564);
and U17088 (N_17088,N_16937,N_16622);
nand U17089 (N_17089,N_16829,N_16859);
xnor U17090 (N_17090,N_16826,N_16698);
xnor U17091 (N_17091,N_16850,N_16599);
nor U17092 (N_17092,N_16606,N_16535);
nand U17093 (N_17093,N_16912,N_16915);
xor U17094 (N_17094,N_16731,N_16866);
xor U17095 (N_17095,N_16816,N_16653);
and U17096 (N_17096,N_16990,N_16843);
xnor U17097 (N_17097,N_16661,N_16768);
or U17098 (N_17098,N_16590,N_16545);
and U17099 (N_17099,N_16819,N_16638);
nor U17100 (N_17100,N_16818,N_16899);
or U17101 (N_17101,N_16506,N_16940);
nand U17102 (N_17102,N_16668,N_16643);
nor U17103 (N_17103,N_16909,N_16746);
and U17104 (N_17104,N_16747,N_16934);
and U17105 (N_17105,N_16679,N_16808);
xor U17106 (N_17106,N_16640,N_16745);
xor U17107 (N_17107,N_16699,N_16967);
nor U17108 (N_17108,N_16945,N_16583);
nand U17109 (N_17109,N_16985,N_16732);
nor U17110 (N_17110,N_16880,N_16738);
nand U17111 (N_17111,N_16612,N_16740);
xnor U17112 (N_17112,N_16881,N_16532);
and U17113 (N_17113,N_16578,N_16712);
or U17114 (N_17114,N_16760,N_16642);
xnor U17115 (N_17115,N_16784,N_16505);
nor U17116 (N_17116,N_16582,N_16651);
or U17117 (N_17117,N_16925,N_16914);
nor U17118 (N_17118,N_16847,N_16964);
or U17119 (N_17119,N_16700,N_16614);
nor U17120 (N_17120,N_16708,N_16677);
xor U17121 (N_17121,N_16887,N_16986);
nand U17122 (N_17122,N_16921,N_16743);
nand U17123 (N_17123,N_16994,N_16665);
or U17124 (N_17124,N_16895,N_16978);
nand U17125 (N_17125,N_16575,N_16974);
or U17126 (N_17126,N_16891,N_16779);
and U17127 (N_17127,N_16722,N_16701);
nor U17128 (N_17128,N_16797,N_16860);
or U17129 (N_17129,N_16581,N_16504);
and U17130 (N_17130,N_16719,N_16503);
nor U17131 (N_17131,N_16662,N_16893);
nor U17132 (N_17132,N_16763,N_16536);
or U17133 (N_17133,N_16605,N_16806);
or U17134 (N_17134,N_16919,N_16548);
or U17135 (N_17135,N_16877,N_16534);
nor U17136 (N_17136,N_16728,N_16853);
nand U17137 (N_17137,N_16659,N_16939);
or U17138 (N_17138,N_16512,N_16996);
nand U17139 (N_17139,N_16810,N_16824);
nor U17140 (N_17140,N_16574,N_16794);
nand U17141 (N_17141,N_16562,N_16825);
xor U17142 (N_17142,N_16688,N_16956);
nor U17143 (N_17143,N_16586,N_16717);
xor U17144 (N_17144,N_16750,N_16603);
and U17145 (N_17145,N_16592,N_16540);
xor U17146 (N_17146,N_16621,N_16697);
and U17147 (N_17147,N_16560,N_16543);
or U17148 (N_17148,N_16570,N_16649);
xor U17149 (N_17149,N_16671,N_16776);
xor U17150 (N_17150,N_16883,N_16559);
nand U17151 (N_17151,N_16591,N_16856);
or U17152 (N_17152,N_16799,N_16872);
nor U17153 (N_17153,N_16672,N_16957);
nor U17154 (N_17154,N_16751,N_16943);
nor U17155 (N_17155,N_16889,N_16998);
nand U17156 (N_17156,N_16584,N_16706);
and U17157 (N_17157,N_16873,N_16827);
nor U17158 (N_17158,N_16647,N_16924);
and U17159 (N_17159,N_16753,N_16884);
and U17160 (N_17160,N_16663,N_16681);
xnor U17161 (N_17161,N_16513,N_16596);
or U17162 (N_17162,N_16674,N_16795);
nand U17163 (N_17163,N_16897,N_16878);
nand U17164 (N_17164,N_16813,N_16625);
xnor U17165 (N_17165,N_16936,N_16780);
nor U17166 (N_17166,N_16531,N_16714);
and U17167 (N_17167,N_16648,N_16542);
or U17168 (N_17168,N_16762,N_16525);
xnor U17169 (N_17169,N_16932,N_16926);
xnor U17170 (N_17170,N_16906,N_16726);
or U17171 (N_17171,N_16777,N_16720);
nor U17172 (N_17172,N_16803,N_16725);
xor U17173 (N_17173,N_16593,N_16837);
or U17174 (N_17174,N_16755,N_16929);
nor U17175 (N_17175,N_16567,N_16565);
and U17176 (N_17176,N_16823,N_16905);
and U17177 (N_17177,N_16778,N_16670);
or U17178 (N_17178,N_16516,N_16520);
and U17179 (N_17179,N_16624,N_16710);
nand U17180 (N_17180,N_16918,N_16983);
and U17181 (N_17181,N_16735,N_16931);
nand U17182 (N_17182,N_16913,N_16617);
and U17183 (N_17183,N_16629,N_16610);
or U17184 (N_17184,N_16691,N_16858);
nand U17185 (N_17185,N_16611,N_16876);
nor U17186 (N_17186,N_16754,N_16972);
xnor U17187 (N_17187,N_16655,N_16657);
or U17188 (N_17188,N_16951,N_16607);
nor U17189 (N_17189,N_16736,N_16958);
and U17190 (N_17190,N_16508,N_16639);
nor U17191 (N_17191,N_16984,N_16802);
xor U17192 (N_17192,N_16835,N_16664);
nand U17193 (N_17193,N_16911,N_16821);
nor U17194 (N_17194,N_16524,N_16523);
and U17195 (N_17195,N_16800,N_16687);
nor U17196 (N_17196,N_16515,N_16946);
nor U17197 (N_17197,N_16770,N_16938);
xor U17198 (N_17198,N_16848,N_16907);
and U17199 (N_17199,N_16537,N_16730);
or U17200 (N_17200,N_16997,N_16660);
nor U17201 (N_17201,N_16982,N_16635);
nor U17202 (N_17202,N_16587,N_16715);
xor U17203 (N_17203,N_16789,N_16563);
xnor U17204 (N_17204,N_16867,N_16527);
nand U17205 (N_17205,N_16995,N_16759);
nand U17206 (N_17206,N_16632,N_16549);
or U17207 (N_17207,N_16694,N_16550);
and U17208 (N_17208,N_16749,N_16703);
nor U17209 (N_17209,N_16890,N_16842);
nor U17210 (N_17210,N_16602,N_16898);
nor U17211 (N_17211,N_16862,N_16546);
xnor U17212 (N_17212,N_16510,N_16933);
or U17213 (N_17213,N_16798,N_16530);
nand U17214 (N_17214,N_16830,N_16849);
xnor U17215 (N_17215,N_16901,N_16781);
and U17216 (N_17216,N_16954,N_16865);
and U17217 (N_17217,N_16518,N_16658);
nand U17218 (N_17218,N_16737,N_16709);
and U17219 (N_17219,N_16833,N_16839);
nor U17220 (N_17220,N_16630,N_16723);
xnor U17221 (N_17221,N_16831,N_16950);
or U17222 (N_17222,N_16902,N_16572);
or U17223 (N_17223,N_16791,N_16600);
nand U17224 (N_17224,N_16949,N_16811);
nor U17225 (N_17225,N_16538,N_16764);
nand U17226 (N_17226,N_16652,N_16875);
nor U17227 (N_17227,N_16692,N_16828);
and U17228 (N_17228,N_16514,N_16526);
nor U17229 (N_17229,N_16623,N_16616);
nand U17230 (N_17230,N_16851,N_16942);
xnor U17231 (N_17231,N_16900,N_16739);
nand U17232 (N_17232,N_16948,N_16507);
and U17233 (N_17233,N_16782,N_16579);
xnor U17234 (N_17234,N_16522,N_16920);
or U17235 (N_17235,N_16977,N_16834);
xnor U17236 (N_17236,N_16989,N_16604);
xor U17237 (N_17237,N_16618,N_16855);
nand U17238 (N_17238,N_16882,N_16666);
xor U17239 (N_17239,N_16541,N_16917);
or U17240 (N_17240,N_16771,N_16705);
or U17241 (N_17241,N_16667,N_16615);
nor U17242 (N_17242,N_16553,N_16669);
xor U17243 (N_17243,N_16864,N_16568);
xor U17244 (N_17244,N_16960,N_16863);
and U17245 (N_17245,N_16857,N_16502);
or U17246 (N_17246,N_16963,N_16561);
xor U17247 (N_17247,N_16774,N_16886);
nand U17248 (N_17248,N_16734,N_16796);
nand U17249 (N_17249,N_16626,N_16927);
or U17250 (N_17250,N_16631,N_16814);
nor U17251 (N_17251,N_16561,N_16508);
or U17252 (N_17252,N_16707,N_16958);
and U17253 (N_17253,N_16567,N_16812);
xor U17254 (N_17254,N_16991,N_16734);
nand U17255 (N_17255,N_16520,N_16941);
xor U17256 (N_17256,N_16521,N_16974);
xor U17257 (N_17257,N_16688,N_16547);
nor U17258 (N_17258,N_16643,N_16589);
or U17259 (N_17259,N_16679,N_16655);
nor U17260 (N_17260,N_16836,N_16756);
nor U17261 (N_17261,N_16638,N_16730);
nor U17262 (N_17262,N_16778,N_16731);
nor U17263 (N_17263,N_16752,N_16961);
or U17264 (N_17264,N_16915,N_16523);
xnor U17265 (N_17265,N_16885,N_16540);
or U17266 (N_17266,N_16540,N_16909);
nor U17267 (N_17267,N_16688,N_16912);
or U17268 (N_17268,N_16943,N_16915);
and U17269 (N_17269,N_16553,N_16652);
or U17270 (N_17270,N_16937,N_16912);
nor U17271 (N_17271,N_16704,N_16864);
nor U17272 (N_17272,N_16724,N_16984);
nand U17273 (N_17273,N_16809,N_16976);
nand U17274 (N_17274,N_16797,N_16952);
and U17275 (N_17275,N_16552,N_16872);
nor U17276 (N_17276,N_16803,N_16509);
or U17277 (N_17277,N_16583,N_16838);
nand U17278 (N_17278,N_16562,N_16667);
and U17279 (N_17279,N_16705,N_16633);
nor U17280 (N_17280,N_16589,N_16682);
and U17281 (N_17281,N_16633,N_16694);
xnor U17282 (N_17282,N_16751,N_16681);
nor U17283 (N_17283,N_16975,N_16712);
xnor U17284 (N_17284,N_16882,N_16693);
and U17285 (N_17285,N_16639,N_16613);
xnor U17286 (N_17286,N_16975,N_16739);
or U17287 (N_17287,N_16945,N_16734);
and U17288 (N_17288,N_16978,N_16635);
xor U17289 (N_17289,N_16671,N_16754);
xor U17290 (N_17290,N_16737,N_16728);
or U17291 (N_17291,N_16793,N_16786);
xnor U17292 (N_17292,N_16560,N_16871);
or U17293 (N_17293,N_16563,N_16686);
or U17294 (N_17294,N_16684,N_16562);
and U17295 (N_17295,N_16664,N_16651);
nor U17296 (N_17296,N_16776,N_16508);
and U17297 (N_17297,N_16791,N_16577);
nand U17298 (N_17298,N_16528,N_16852);
and U17299 (N_17299,N_16930,N_16904);
nor U17300 (N_17300,N_16787,N_16606);
xor U17301 (N_17301,N_16836,N_16895);
xor U17302 (N_17302,N_16506,N_16976);
and U17303 (N_17303,N_16737,N_16870);
xnor U17304 (N_17304,N_16627,N_16780);
and U17305 (N_17305,N_16535,N_16532);
xnor U17306 (N_17306,N_16741,N_16969);
nor U17307 (N_17307,N_16769,N_16989);
xor U17308 (N_17308,N_16613,N_16953);
nor U17309 (N_17309,N_16833,N_16598);
and U17310 (N_17310,N_16935,N_16668);
nor U17311 (N_17311,N_16558,N_16909);
nand U17312 (N_17312,N_16722,N_16682);
nor U17313 (N_17313,N_16650,N_16959);
nor U17314 (N_17314,N_16826,N_16656);
or U17315 (N_17315,N_16679,N_16725);
or U17316 (N_17316,N_16564,N_16691);
nand U17317 (N_17317,N_16976,N_16545);
or U17318 (N_17318,N_16767,N_16650);
nor U17319 (N_17319,N_16502,N_16796);
and U17320 (N_17320,N_16614,N_16582);
xor U17321 (N_17321,N_16503,N_16847);
xnor U17322 (N_17322,N_16595,N_16732);
and U17323 (N_17323,N_16643,N_16824);
nor U17324 (N_17324,N_16756,N_16673);
xnor U17325 (N_17325,N_16602,N_16612);
or U17326 (N_17326,N_16754,N_16716);
nand U17327 (N_17327,N_16637,N_16602);
nor U17328 (N_17328,N_16764,N_16967);
xnor U17329 (N_17329,N_16929,N_16728);
nor U17330 (N_17330,N_16860,N_16714);
or U17331 (N_17331,N_16560,N_16916);
nand U17332 (N_17332,N_16876,N_16518);
xor U17333 (N_17333,N_16525,N_16774);
and U17334 (N_17334,N_16532,N_16738);
nand U17335 (N_17335,N_16923,N_16836);
xnor U17336 (N_17336,N_16876,N_16921);
and U17337 (N_17337,N_16746,N_16551);
xor U17338 (N_17338,N_16911,N_16958);
xnor U17339 (N_17339,N_16537,N_16756);
nor U17340 (N_17340,N_16747,N_16933);
nor U17341 (N_17341,N_16543,N_16715);
nand U17342 (N_17342,N_16942,N_16829);
or U17343 (N_17343,N_16974,N_16922);
or U17344 (N_17344,N_16958,N_16771);
xor U17345 (N_17345,N_16923,N_16577);
xor U17346 (N_17346,N_16517,N_16775);
nor U17347 (N_17347,N_16897,N_16648);
and U17348 (N_17348,N_16638,N_16884);
xnor U17349 (N_17349,N_16886,N_16651);
nor U17350 (N_17350,N_16895,N_16977);
or U17351 (N_17351,N_16506,N_16950);
or U17352 (N_17352,N_16694,N_16965);
and U17353 (N_17353,N_16970,N_16658);
and U17354 (N_17354,N_16950,N_16932);
or U17355 (N_17355,N_16854,N_16864);
xnor U17356 (N_17356,N_16836,N_16735);
xor U17357 (N_17357,N_16735,N_16859);
nand U17358 (N_17358,N_16553,N_16675);
nor U17359 (N_17359,N_16639,N_16618);
or U17360 (N_17360,N_16625,N_16788);
nand U17361 (N_17361,N_16856,N_16510);
or U17362 (N_17362,N_16975,N_16656);
and U17363 (N_17363,N_16936,N_16949);
or U17364 (N_17364,N_16765,N_16535);
and U17365 (N_17365,N_16727,N_16934);
and U17366 (N_17366,N_16743,N_16608);
xor U17367 (N_17367,N_16914,N_16855);
and U17368 (N_17368,N_16680,N_16690);
or U17369 (N_17369,N_16708,N_16950);
nand U17370 (N_17370,N_16922,N_16906);
nand U17371 (N_17371,N_16632,N_16967);
and U17372 (N_17372,N_16957,N_16668);
and U17373 (N_17373,N_16771,N_16928);
nand U17374 (N_17374,N_16889,N_16507);
nand U17375 (N_17375,N_16663,N_16578);
nor U17376 (N_17376,N_16964,N_16591);
xnor U17377 (N_17377,N_16880,N_16984);
or U17378 (N_17378,N_16989,N_16592);
nand U17379 (N_17379,N_16959,N_16858);
or U17380 (N_17380,N_16725,N_16941);
and U17381 (N_17381,N_16927,N_16636);
or U17382 (N_17382,N_16820,N_16743);
or U17383 (N_17383,N_16875,N_16870);
nand U17384 (N_17384,N_16726,N_16750);
nand U17385 (N_17385,N_16628,N_16641);
nor U17386 (N_17386,N_16802,N_16844);
or U17387 (N_17387,N_16923,N_16884);
nand U17388 (N_17388,N_16532,N_16922);
or U17389 (N_17389,N_16907,N_16539);
nor U17390 (N_17390,N_16818,N_16831);
nor U17391 (N_17391,N_16877,N_16942);
xnor U17392 (N_17392,N_16617,N_16920);
xnor U17393 (N_17393,N_16954,N_16710);
nor U17394 (N_17394,N_16708,N_16605);
nand U17395 (N_17395,N_16550,N_16767);
nand U17396 (N_17396,N_16588,N_16558);
nor U17397 (N_17397,N_16935,N_16627);
and U17398 (N_17398,N_16842,N_16986);
and U17399 (N_17399,N_16653,N_16933);
nor U17400 (N_17400,N_16558,N_16707);
xor U17401 (N_17401,N_16629,N_16763);
nor U17402 (N_17402,N_16650,N_16917);
nand U17403 (N_17403,N_16801,N_16877);
nor U17404 (N_17404,N_16675,N_16843);
nor U17405 (N_17405,N_16734,N_16702);
nand U17406 (N_17406,N_16899,N_16805);
nor U17407 (N_17407,N_16611,N_16649);
or U17408 (N_17408,N_16979,N_16933);
nor U17409 (N_17409,N_16910,N_16751);
or U17410 (N_17410,N_16644,N_16817);
and U17411 (N_17411,N_16601,N_16502);
and U17412 (N_17412,N_16873,N_16670);
nor U17413 (N_17413,N_16814,N_16967);
nor U17414 (N_17414,N_16698,N_16646);
or U17415 (N_17415,N_16740,N_16964);
xnor U17416 (N_17416,N_16731,N_16981);
and U17417 (N_17417,N_16974,N_16564);
xor U17418 (N_17418,N_16724,N_16917);
xor U17419 (N_17419,N_16976,N_16995);
xnor U17420 (N_17420,N_16709,N_16941);
nor U17421 (N_17421,N_16524,N_16501);
xor U17422 (N_17422,N_16849,N_16789);
and U17423 (N_17423,N_16802,N_16819);
or U17424 (N_17424,N_16791,N_16738);
or U17425 (N_17425,N_16585,N_16964);
nor U17426 (N_17426,N_16844,N_16501);
and U17427 (N_17427,N_16614,N_16738);
or U17428 (N_17428,N_16530,N_16714);
or U17429 (N_17429,N_16524,N_16791);
and U17430 (N_17430,N_16585,N_16574);
or U17431 (N_17431,N_16887,N_16812);
or U17432 (N_17432,N_16989,N_16930);
nand U17433 (N_17433,N_16739,N_16747);
nand U17434 (N_17434,N_16879,N_16606);
or U17435 (N_17435,N_16675,N_16618);
nand U17436 (N_17436,N_16568,N_16896);
nor U17437 (N_17437,N_16948,N_16513);
or U17438 (N_17438,N_16501,N_16811);
nor U17439 (N_17439,N_16698,N_16534);
and U17440 (N_17440,N_16886,N_16928);
or U17441 (N_17441,N_16672,N_16927);
nand U17442 (N_17442,N_16636,N_16953);
or U17443 (N_17443,N_16821,N_16699);
or U17444 (N_17444,N_16627,N_16912);
nand U17445 (N_17445,N_16559,N_16517);
xnor U17446 (N_17446,N_16808,N_16841);
and U17447 (N_17447,N_16909,N_16725);
and U17448 (N_17448,N_16843,N_16627);
and U17449 (N_17449,N_16995,N_16713);
or U17450 (N_17450,N_16704,N_16942);
xnor U17451 (N_17451,N_16959,N_16895);
nand U17452 (N_17452,N_16600,N_16558);
xnor U17453 (N_17453,N_16528,N_16513);
or U17454 (N_17454,N_16630,N_16754);
xnor U17455 (N_17455,N_16512,N_16826);
xnor U17456 (N_17456,N_16976,N_16945);
and U17457 (N_17457,N_16926,N_16645);
nor U17458 (N_17458,N_16591,N_16576);
or U17459 (N_17459,N_16847,N_16732);
nor U17460 (N_17460,N_16828,N_16929);
or U17461 (N_17461,N_16589,N_16588);
nor U17462 (N_17462,N_16706,N_16725);
xnor U17463 (N_17463,N_16736,N_16881);
nand U17464 (N_17464,N_16653,N_16710);
xnor U17465 (N_17465,N_16800,N_16851);
or U17466 (N_17466,N_16929,N_16901);
or U17467 (N_17467,N_16707,N_16601);
and U17468 (N_17468,N_16756,N_16719);
xnor U17469 (N_17469,N_16522,N_16660);
xnor U17470 (N_17470,N_16802,N_16631);
and U17471 (N_17471,N_16586,N_16579);
and U17472 (N_17472,N_16923,N_16573);
nand U17473 (N_17473,N_16700,N_16719);
nand U17474 (N_17474,N_16539,N_16655);
nor U17475 (N_17475,N_16614,N_16938);
xnor U17476 (N_17476,N_16956,N_16523);
nor U17477 (N_17477,N_16931,N_16528);
nor U17478 (N_17478,N_16898,N_16664);
xnor U17479 (N_17479,N_16888,N_16664);
xnor U17480 (N_17480,N_16639,N_16864);
and U17481 (N_17481,N_16500,N_16654);
nor U17482 (N_17482,N_16832,N_16682);
or U17483 (N_17483,N_16565,N_16706);
and U17484 (N_17484,N_16695,N_16659);
nand U17485 (N_17485,N_16850,N_16870);
or U17486 (N_17486,N_16894,N_16932);
or U17487 (N_17487,N_16567,N_16658);
xor U17488 (N_17488,N_16598,N_16885);
or U17489 (N_17489,N_16556,N_16668);
or U17490 (N_17490,N_16884,N_16708);
nor U17491 (N_17491,N_16503,N_16756);
nand U17492 (N_17492,N_16844,N_16982);
nand U17493 (N_17493,N_16907,N_16612);
nor U17494 (N_17494,N_16832,N_16528);
nand U17495 (N_17495,N_16953,N_16958);
or U17496 (N_17496,N_16674,N_16649);
nor U17497 (N_17497,N_16915,N_16542);
xor U17498 (N_17498,N_16768,N_16917);
or U17499 (N_17499,N_16710,N_16884);
or U17500 (N_17500,N_17198,N_17383);
nand U17501 (N_17501,N_17202,N_17475);
or U17502 (N_17502,N_17128,N_17416);
and U17503 (N_17503,N_17478,N_17459);
or U17504 (N_17504,N_17207,N_17238);
and U17505 (N_17505,N_17010,N_17485);
nand U17506 (N_17506,N_17012,N_17251);
and U17507 (N_17507,N_17394,N_17448);
nand U17508 (N_17508,N_17280,N_17480);
xnor U17509 (N_17509,N_17494,N_17147);
or U17510 (N_17510,N_17036,N_17337);
and U17511 (N_17511,N_17250,N_17163);
nand U17512 (N_17512,N_17189,N_17232);
xnor U17513 (N_17513,N_17275,N_17146);
nor U17514 (N_17514,N_17242,N_17328);
nor U17515 (N_17515,N_17210,N_17068);
and U17516 (N_17516,N_17150,N_17365);
nor U17517 (N_17517,N_17083,N_17355);
or U17518 (N_17518,N_17130,N_17339);
xor U17519 (N_17519,N_17477,N_17199);
nor U17520 (N_17520,N_17118,N_17284);
and U17521 (N_17521,N_17079,N_17161);
or U17522 (N_17522,N_17447,N_17122);
nand U17523 (N_17523,N_17126,N_17315);
xor U17524 (N_17524,N_17261,N_17100);
xnor U17525 (N_17525,N_17353,N_17341);
and U17526 (N_17526,N_17316,N_17167);
or U17527 (N_17527,N_17295,N_17006);
nand U17528 (N_17528,N_17352,N_17392);
nand U17529 (N_17529,N_17183,N_17466);
or U17530 (N_17530,N_17299,N_17443);
xor U17531 (N_17531,N_17450,N_17446);
nor U17532 (N_17532,N_17347,N_17405);
nor U17533 (N_17533,N_17029,N_17180);
xor U17534 (N_17534,N_17170,N_17211);
or U17535 (N_17535,N_17219,N_17402);
nor U17536 (N_17536,N_17041,N_17194);
xnor U17537 (N_17537,N_17488,N_17433);
and U17538 (N_17538,N_17314,N_17472);
or U17539 (N_17539,N_17473,N_17438);
nand U17540 (N_17540,N_17022,N_17270);
and U17541 (N_17541,N_17111,N_17437);
xor U17542 (N_17542,N_17268,N_17432);
nand U17543 (N_17543,N_17181,N_17252);
and U17544 (N_17544,N_17296,N_17186);
nor U17545 (N_17545,N_17049,N_17423);
or U17546 (N_17546,N_17227,N_17411);
nor U17547 (N_17547,N_17135,N_17336);
or U17548 (N_17548,N_17214,N_17212);
xor U17549 (N_17549,N_17182,N_17192);
or U17550 (N_17550,N_17326,N_17149);
or U17551 (N_17551,N_17322,N_17174);
or U17552 (N_17552,N_17230,N_17441);
nand U17553 (N_17553,N_17308,N_17412);
nor U17554 (N_17554,N_17101,N_17329);
and U17555 (N_17555,N_17074,N_17004);
xor U17556 (N_17556,N_17116,N_17358);
and U17557 (N_17557,N_17440,N_17203);
nand U17558 (N_17558,N_17027,N_17060);
and U17559 (N_17559,N_17063,N_17046);
xnor U17560 (N_17560,N_17240,N_17127);
nor U17561 (N_17561,N_17095,N_17094);
nor U17562 (N_17562,N_17221,N_17097);
and U17563 (N_17563,N_17385,N_17499);
nor U17564 (N_17564,N_17318,N_17469);
nor U17565 (N_17565,N_17445,N_17265);
nand U17566 (N_17566,N_17037,N_17114);
nor U17567 (N_17567,N_17082,N_17279);
xnor U17568 (N_17568,N_17248,N_17197);
xnor U17569 (N_17569,N_17388,N_17136);
and U17570 (N_17570,N_17398,N_17104);
nor U17571 (N_17571,N_17382,N_17304);
nor U17572 (N_17572,N_17056,N_17014);
nor U17573 (N_17573,N_17334,N_17332);
nor U17574 (N_17574,N_17307,N_17093);
or U17575 (N_17575,N_17498,N_17073);
and U17576 (N_17576,N_17138,N_17312);
and U17577 (N_17577,N_17455,N_17291);
xnor U17578 (N_17578,N_17044,N_17461);
and U17579 (N_17579,N_17324,N_17195);
and U17580 (N_17580,N_17397,N_17487);
nand U17581 (N_17581,N_17452,N_17172);
and U17582 (N_17582,N_17470,N_17298);
xnor U17583 (N_17583,N_17401,N_17017);
nand U17584 (N_17584,N_17076,N_17342);
and U17585 (N_17585,N_17178,N_17200);
or U17586 (N_17586,N_17369,N_17255);
or U17587 (N_17587,N_17370,N_17368);
or U17588 (N_17588,N_17393,N_17306);
nand U17589 (N_17589,N_17495,N_17463);
nor U17590 (N_17590,N_17436,N_17099);
or U17591 (N_17591,N_17035,N_17143);
nand U17592 (N_17592,N_17069,N_17429);
nand U17593 (N_17593,N_17077,N_17206);
nor U17594 (N_17594,N_17263,N_17154);
or U17595 (N_17595,N_17327,N_17223);
nor U17596 (N_17596,N_17415,N_17427);
or U17597 (N_17597,N_17108,N_17439);
nor U17598 (N_17598,N_17343,N_17051);
nor U17599 (N_17599,N_17335,N_17374);
nand U17600 (N_17600,N_17000,N_17205);
or U17601 (N_17601,N_17493,N_17396);
xor U17602 (N_17602,N_17460,N_17020);
xnor U17603 (N_17603,N_17271,N_17153);
or U17604 (N_17604,N_17418,N_17058);
nor U17605 (N_17605,N_17325,N_17377);
or U17606 (N_17606,N_17344,N_17399);
xnor U17607 (N_17607,N_17317,N_17254);
nand U17608 (N_17608,N_17474,N_17176);
nor U17609 (N_17609,N_17030,N_17257);
nand U17610 (N_17610,N_17262,N_17145);
nor U17611 (N_17611,N_17103,N_17237);
nor U17612 (N_17612,N_17018,N_17115);
nor U17613 (N_17613,N_17346,N_17430);
and U17614 (N_17614,N_17349,N_17410);
xor U17615 (N_17615,N_17162,N_17239);
or U17616 (N_17616,N_17244,N_17323);
xor U17617 (N_17617,N_17387,N_17464);
nand U17618 (N_17618,N_17084,N_17390);
nand U17619 (N_17619,N_17380,N_17266);
or U17620 (N_17620,N_17013,N_17067);
nor U17621 (N_17621,N_17444,N_17070);
xor U17622 (N_17622,N_17208,N_17276);
nand U17623 (N_17623,N_17120,N_17098);
nor U17624 (N_17624,N_17096,N_17129);
nand U17625 (N_17625,N_17362,N_17021);
and U17626 (N_17626,N_17081,N_17222);
or U17627 (N_17627,N_17497,N_17159);
xnor U17628 (N_17628,N_17483,N_17330);
nand U17629 (N_17629,N_17391,N_17031);
nand U17630 (N_17630,N_17338,N_17139);
nand U17631 (N_17631,N_17288,N_17264);
xnor U17632 (N_17632,N_17491,N_17476);
or U17633 (N_17633,N_17413,N_17121);
nand U17634 (N_17634,N_17196,N_17218);
nor U17635 (N_17635,N_17309,N_17340);
xnor U17636 (N_17636,N_17231,N_17356);
and U17637 (N_17637,N_17300,N_17033);
or U17638 (N_17638,N_17320,N_17061);
and U17639 (N_17639,N_17243,N_17331);
or U17640 (N_17640,N_17064,N_17071);
nand U17641 (N_17641,N_17204,N_17019);
and U17642 (N_17642,N_17354,N_17384);
xor U17643 (N_17643,N_17420,N_17386);
and U17644 (N_17644,N_17190,N_17363);
xnor U17645 (N_17645,N_17481,N_17102);
and U17646 (N_17646,N_17241,N_17175);
nor U17647 (N_17647,N_17419,N_17272);
nor U17648 (N_17648,N_17187,N_17152);
and U17649 (N_17649,N_17245,N_17267);
and U17650 (N_17650,N_17080,N_17158);
nor U17651 (N_17651,N_17132,N_17213);
nor U17652 (N_17652,N_17305,N_17414);
xor U17653 (N_17653,N_17372,N_17140);
nor U17654 (N_17654,N_17313,N_17112);
xnor U17655 (N_17655,N_17085,N_17297);
xor U17656 (N_17656,N_17148,N_17028);
nor U17657 (N_17657,N_17089,N_17424);
nor U17658 (N_17658,N_17292,N_17294);
xnor U17659 (N_17659,N_17364,N_17426);
nor U17660 (N_17660,N_17359,N_17421);
xnor U17661 (N_17661,N_17404,N_17425);
and U17662 (N_17662,N_17256,N_17042);
nand U17663 (N_17663,N_17075,N_17293);
nand U17664 (N_17664,N_17166,N_17220);
nor U17665 (N_17665,N_17034,N_17348);
and U17666 (N_17666,N_17065,N_17216);
or U17667 (N_17667,N_17005,N_17050);
xor U17668 (N_17668,N_17133,N_17273);
and U17669 (N_17669,N_17465,N_17072);
nand U17670 (N_17670,N_17281,N_17278);
and U17671 (N_17671,N_17454,N_17226);
nor U17672 (N_17672,N_17259,N_17224);
or U17673 (N_17673,N_17078,N_17052);
nand U17674 (N_17674,N_17131,N_17428);
or U17675 (N_17675,N_17225,N_17449);
nor U17676 (N_17676,N_17236,N_17124);
nor U17677 (N_17677,N_17045,N_17389);
and U17678 (N_17678,N_17177,N_17422);
or U17679 (N_17679,N_17468,N_17467);
nand U17680 (N_17680,N_17302,N_17016);
nor U17681 (N_17681,N_17253,N_17217);
and U17682 (N_17682,N_17451,N_17185);
nor U17683 (N_17683,N_17179,N_17490);
nor U17684 (N_17684,N_17001,N_17274);
nand U17685 (N_17685,N_17173,N_17113);
nor U17686 (N_17686,N_17417,N_17053);
and U17687 (N_17687,N_17289,N_17011);
xor U17688 (N_17688,N_17040,N_17310);
xor U17689 (N_17689,N_17039,N_17457);
xor U17690 (N_17690,N_17168,N_17286);
xor U17691 (N_17691,N_17290,N_17048);
nand U17692 (N_17692,N_17025,N_17106);
xnor U17693 (N_17693,N_17054,N_17376);
and U17694 (N_17694,N_17165,N_17090);
or U17695 (N_17695,N_17109,N_17350);
and U17696 (N_17696,N_17169,N_17191);
xnor U17697 (N_17697,N_17373,N_17247);
xnor U17698 (N_17698,N_17458,N_17351);
nor U17699 (N_17699,N_17395,N_17026);
xor U17700 (N_17700,N_17269,N_17151);
and U17701 (N_17701,N_17201,N_17091);
xor U17702 (N_17702,N_17233,N_17141);
nand U17703 (N_17703,N_17489,N_17249);
xnor U17704 (N_17704,N_17345,N_17366);
or U17705 (N_17705,N_17038,N_17007);
nor U17706 (N_17706,N_17333,N_17406);
and U17707 (N_17707,N_17055,N_17367);
nand U17708 (N_17708,N_17215,N_17285);
and U17709 (N_17709,N_17434,N_17024);
nand U17710 (N_17710,N_17456,N_17125);
nand U17711 (N_17711,N_17319,N_17379);
nor U17712 (N_17712,N_17375,N_17229);
xor U17713 (N_17713,N_17142,N_17408);
or U17714 (N_17714,N_17403,N_17287);
xor U17715 (N_17715,N_17087,N_17107);
nor U17716 (N_17716,N_17479,N_17407);
or U17717 (N_17717,N_17371,N_17110);
nand U17718 (N_17718,N_17357,N_17134);
and U17719 (N_17719,N_17435,N_17193);
or U17720 (N_17720,N_17160,N_17361);
nand U17721 (N_17721,N_17023,N_17409);
or U17722 (N_17722,N_17144,N_17117);
xnor U17723 (N_17723,N_17066,N_17360);
xor U17724 (N_17724,N_17486,N_17171);
or U17725 (N_17725,N_17188,N_17484);
nor U17726 (N_17726,N_17492,N_17156);
or U17727 (N_17727,N_17453,N_17260);
or U17728 (N_17728,N_17311,N_17471);
xor U17729 (N_17729,N_17209,N_17228);
and U17730 (N_17730,N_17009,N_17431);
nor U17731 (N_17731,N_17282,N_17496);
nor U17732 (N_17732,N_17157,N_17283);
nand U17733 (N_17733,N_17378,N_17105);
nor U17734 (N_17734,N_17442,N_17303);
nor U17735 (N_17735,N_17015,N_17092);
or U17736 (N_17736,N_17062,N_17137);
xnor U17737 (N_17737,N_17462,N_17277);
nand U17738 (N_17738,N_17088,N_17301);
nor U17739 (N_17739,N_17482,N_17032);
xnor U17740 (N_17740,N_17002,N_17246);
nor U17741 (N_17741,N_17258,N_17003);
and U17742 (N_17742,N_17123,N_17164);
or U17743 (N_17743,N_17008,N_17043);
nor U17744 (N_17744,N_17234,N_17086);
and U17745 (N_17745,N_17235,N_17155);
nand U17746 (N_17746,N_17400,N_17381);
xor U17747 (N_17747,N_17059,N_17119);
nand U17748 (N_17748,N_17321,N_17057);
xnor U17749 (N_17749,N_17047,N_17184);
xor U17750 (N_17750,N_17399,N_17442);
nor U17751 (N_17751,N_17474,N_17305);
or U17752 (N_17752,N_17337,N_17107);
nor U17753 (N_17753,N_17398,N_17392);
xor U17754 (N_17754,N_17179,N_17471);
nor U17755 (N_17755,N_17230,N_17126);
or U17756 (N_17756,N_17179,N_17047);
and U17757 (N_17757,N_17216,N_17329);
xnor U17758 (N_17758,N_17205,N_17467);
xnor U17759 (N_17759,N_17468,N_17007);
and U17760 (N_17760,N_17047,N_17045);
xnor U17761 (N_17761,N_17029,N_17427);
xor U17762 (N_17762,N_17105,N_17162);
or U17763 (N_17763,N_17331,N_17093);
nor U17764 (N_17764,N_17236,N_17352);
xor U17765 (N_17765,N_17026,N_17019);
or U17766 (N_17766,N_17028,N_17036);
xnor U17767 (N_17767,N_17452,N_17003);
nand U17768 (N_17768,N_17305,N_17437);
nand U17769 (N_17769,N_17262,N_17169);
and U17770 (N_17770,N_17286,N_17116);
nand U17771 (N_17771,N_17227,N_17144);
or U17772 (N_17772,N_17351,N_17359);
nand U17773 (N_17773,N_17141,N_17119);
and U17774 (N_17774,N_17018,N_17405);
nand U17775 (N_17775,N_17247,N_17263);
or U17776 (N_17776,N_17408,N_17472);
nor U17777 (N_17777,N_17338,N_17028);
or U17778 (N_17778,N_17479,N_17260);
and U17779 (N_17779,N_17010,N_17126);
nor U17780 (N_17780,N_17371,N_17349);
xnor U17781 (N_17781,N_17009,N_17324);
nand U17782 (N_17782,N_17140,N_17317);
or U17783 (N_17783,N_17065,N_17319);
or U17784 (N_17784,N_17072,N_17452);
nor U17785 (N_17785,N_17254,N_17151);
and U17786 (N_17786,N_17317,N_17177);
xnor U17787 (N_17787,N_17104,N_17089);
nor U17788 (N_17788,N_17441,N_17416);
and U17789 (N_17789,N_17292,N_17298);
nand U17790 (N_17790,N_17106,N_17089);
and U17791 (N_17791,N_17403,N_17232);
nor U17792 (N_17792,N_17411,N_17110);
nor U17793 (N_17793,N_17489,N_17328);
or U17794 (N_17794,N_17050,N_17460);
and U17795 (N_17795,N_17299,N_17005);
nor U17796 (N_17796,N_17256,N_17112);
nor U17797 (N_17797,N_17241,N_17132);
and U17798 (N_17798,N_17441,N_17478);
nor U17799 (N_17799,N_17130,N_17139);
xor U17800 (N_17800,N_17216,N_17400);
and U17801 (N_17801,N_17240,N_17290);
nand U17802 (N_17802,N_17379,N_17420);
or U17803 (N_17803,N_17072,N_17458);
and U17804 (N_17804,N_17418,N_17378);
and U17805 (N_17805,N_17330,N_17051);
or U17806 (N_17806,N_17255,N_17290);
xnor U17807 (N_17807,N_17214,N_17272);
or U17808 (N_17808,N_17382,N_17392);
xnor U17809 (N_17809,N_17498,N_17402);
and U17810 (N_17810,N_17194,N_17267);
and U17811 (N_17811,N_17394,N_17366);
xor U17812 (N_17812,N_17064,N_17146);
and U17813 (N_17813,N_17368,N_17250);
or U17814 (N_17814,N_17292,N_17268);
xnor U17815 (N_17815,N_17276,N_17300);
nand U17816 (N_17816,N_17124,N_17209);
and U17817 (N_17817,N_17345,N_17041);
xor U17818 (N_17818,N_17310,N_17441);
and U17819 (N_17819,N_17464,N_17161);
xnor U17820 (N_17820,N_17234,N_17470);
xor U17821 (N_17821,N_17098,N_17061);
nor U17822 (N_17822,N_17317,N_17222);
and U17823 (N_17823,N_17068,N_17027);
nand U17824 (N_17824,N_17278,N_17250);
xor U17825 (N_17825,N_17292,N_17315);
or U17826 (N_17826,N_17217,N_17290);
nor U17827 (N_17827,N_17273,N_17373);
xnor U17828 (N_17828,N_17359,N_17168);
nor U17829 (N_17829,N_17307,N_17089);
xnor U17830 (N_17830,N_17462,N_17265);
nor U17831 (N_17831,N_17170,N_17338);
nor U17832 (N_17832,N_17417,N_17233);
nor U17833 (N_17833,N_17219,N_17035);
nor U17834 (N_17834,N_17208,N_17488);
and U17835 (N_17835,N_17391,N_17349);
nand U17836 (N_17836,N_17420,N_17080);
nor U17837 (N_17837,N_17377,N_17278);
or U17838 (N_17838,N_17096,N_17147);
nor U17839 (N_17839,N_17467,N_17096);
or U17840 (N_17840,N_17333,N_17432);
nand U17841 (N_17841,N_17098,N_17100);
nand U17842 (N_17842,N_17009,N_17382);
and U17843 (N_17843,N_17047,N_17349);
and U17844 (N_17844,N_17109,N_17345);
xor U17845 (N_17845,N_17343,N_17076);
nand U17846 (N_17846,N_17473,N_17229);
xnor U17847 (N_17847,N_17367,N_17102);
xor U17848 (N_17848,N_17481,N_17129);
nand U17849 (N_17849,N_17001,N_17195);
and U17850 (N_17850,N_17040,N_17404);
or U17851 (N_17851,N_17413,N_17386);
nor U17852 (N_17852,N_17081,N_17164);
or U17853 (N_17853,N_17007,N_17411);
or U17854 (N_17854,N_17432,N_17119);
nand U17855 (N_17855,N_17386,N_17279);
nand U17856 (N_17856,N_17394,N_17458);
nor U17857 (N_17857,N_17417,N_17113);
or U17858 (N_17858,N_17494,N_17302);
and U17859 (N_17859,N_17465,N_17045);
or U17860 (N_17860,N_17040,N_17069);
xor U17861 (N_17861,N_17402,N_17215);
or U17862 (N_17862,N_17356,N_17025);
or U17863 (N_17863,N_17027,N_17361);
and U17864 (N_17864,N_17124,N_17347);
nand U17865 (N_17865,N_17217,N_17292);
or U17866 (N_17866,N_17274,N_17461);
and U17867 (N_17867,N_17135,N_17199);
nand U17868 (N_17868,N_17498,N_17188);
xor U17869 (N_17869,N_17483,N_17192);
xnor U17870 (N_17870,N_17017,N_17364);
nand U17871 (N_17871,N_17130,N_17096);
nor U17872 (N_17872,N_17045,N_17335);
and U17873 (N_17873,N_17263,N_17290);
or U17874 (N_17874,N_17459,N_17048);
xor U17875 (N_17875,N_17313,N_17491);
or U17876 (N_17876,N_17000,N_17233);
nor U17877 (N_17877,N_17471,N_17159);
or U17878 (N_17878,N_17008,N_17082);
xnor U17879 (N_17879,N_17128,N_17250);
and U17880 (N_17880,N_17132,N_17197);
xor U17881 (N_17881,N_17299,N_17211);
nand U17882 (N_17882,N_17183,N_17174);
nand U17883 (N_17883,N_17311,N_17063);
and U17884 (N_17884,N_17292,N_17280);
and U17885 (N_17885,N_17128,N_17016);
and U17886 (N_17886,N_17184,N_17005);
xnor U17887 (N_17887,N_17140,N_17168);
nor U17888 (N_17888,N_17228,N_17080);
and U17889 (N_17889,N_17195,N_17058);
xor U17890 (N_17890,N_17136,N_17289);
or U17891 (N_17891,N_17186,N_17332);
xor U17892 (N_17892,N_17299,N_17354);
or U17893 (N_17893,N_17287,N_17453);
and U17894 (N_17894,N_17403,N_17219);
nand U17895 (N_17895,N_17005,N_17321);
nor U17896 (N_17896,N_17014,N_17226);
and U17897 (N_17897,N_17171,N_17058);
nor U17898 (N_17898,N_17292,N_17308);
and U17899 (N_17899,N_17022,N_17472);
nor U17900 (N_17900,N_17440,N_17043);
and U17901 (N_17901,N_17135,N_17203);
or U17902 (N_17902,N_17072,N_17499);
nor U17903 (N_17903,N_17121,N_17046);
nor U17904 (N_17904,N_17179,N_17253);
and U17905 (N_17905,N_17490,N_17222);
xnor U17906 (N_17906,N_17031,N_17056);
xor U17907 (N_17907,N_17005,N_17337);
or U17908 (N_17908,N_17486,N_17066);
nor U17909 (N_17909,N_17099,N_17299);
nor U17910 (N_17910,N_17449,N_17404);
or U17911 (N_17911,N_17112,N_17108);
nor U17912 (N_17912,N_17058,N_17088);
nor U17913 (N_17913,N_17098,N_17222);
or U17914 (N_17914,N_17305,N_17043);
or U17915 (N_17915,N_17126,N_17088);
or U17916 (N_17916,N_17394,N_17263);
and U17917 (N_17917,N_17042,N_17196);
xnor U17918 (N_17918,N_17278,N_17400);
or U17919 (N_17919,N_17096,N_17323);
or U17920 (N_17920,N_17141,N_17481);
nand U17921 (N_17921,N_17085,N_17027);
and U17922 (N_17922,N_17199,N_17296);
xnor U17923 (N_17923,N_17351,N_17335);
and U17924 (N_17924,N_17048,N_17134);
nand U17925 (N_17925,N_17148,N_17393);
nand U17926 (N_17926,N_17145,N_17094);
xnor U17927 (N_17927,N_17116,N_17423);
nand U17928 (N_17928,N_17038,N_17389);
and U17929 (N_17929,N_17046,N_17055);
nand U17930 (N_17930,N_17422,N_17345);
xnor U17931 (N_17931,N_17401,N_17456);
or U17932 (N_17932,N_17474,N_17446);
or U17933 (N_17933,N_17321,N_17244);
and U17934 (N_17934,N_17395,N_17340);
and U17935 (N_17935,N_17310,N_17194);
xor U17936 (N_17936,N_17009,N_17071);
xnor U17937 (N_17937,N_17291,N_17461);
nand U17938 (N_17938,N_17287,N_17156);
nor U17939 (N_17939,N_17262,N_17155);
nor U17940 (N_17940,N_17064,N_17022);
nor U17941 (N_17941,N_17072,N_17200);
nand U17942 (N_17942,N_17268,N_17403);
or U17943 (N_17943,N_17429,N_17423);
xnor U17944 (N_17944,N_17096,N_17195);
and U17945 (N_17945,N_17338,N_17254);
nor U17946 (N_17946,N_17167,N_17192);
or U17947 (N_17947,N_17281,N_17019);
nor U17948 (N_17948,N_17152,N_17477);
nand U17949 (N_17949,N_17447,N_17213);
and U17950 (N_17950,N_17454,N_17099);
nor U17951 (N_17951,N_17465,N_17044);
nor U17952 (N_17952,N_17481,N_17054);
nor U17953 (N_17953,N_17424,N_17154);
xor U17954 (N_17954,N_17297,N_17090);
nand U17955 (N_17955,N_17397,N_17089);
or U17956 (N_17956,N_17024,N_17168);
xnor U17957 (N_17957,N_17427,N_17432);
and U17958 (N_17958,N_17440,N_17238);
nor U17959 (N_17959,N_17358,N_17429);
nor U17960 (N_17960,N_17186,N_17494);
or U17961 (N_17961,N_17164,N_17254);
or U17962 (N_17962,N_17387,N_17114);
xor U17963 (N_17963,N_17402,N_17394);
nand U17964 (N_17964,N_17327,N_17433);
or U17965 (N_17965,N_17296,N_17482);
nand U17966 (N_17966,N_17153,N_17326);
nand U17967 (N_17967,N_17091,N_17351);
or U17968 (N_17968,N_17259,N_17234);
nand U17969 (N_17969,N_17353,N_17080);
nand U17970 (N_17970,N_17213,N_17229);
and U17971 (N_17971,N_17492,N_17032);
or U17972 (N_17972,N_17413,N_17111);
or U17973 (N_17973,N_17410,N_17426);
or U17974 (N_17974,N_17332,N_17101);
nor U17975 (N_17975,N_17317,N_17347);
nand U17976 (N_17976,N_17460,N_17198);
nand U17977 (N_17977,N_17443,N_17360);
nor U17978 (N_17978,N_17377,N_17424);
or U17979 (N_17979,N_17040,N_17230);
xnor U17980 (N_17980,N_17156,N_17044);
nand U17981 (N_17981,N_17039,N_17225);
and U17982 (N_17982,N_17336,N_17411);
nand U17983 (N_17983,N_17342,N_17171);
and U17984 (N_17984,N_17096,N_17339);
nor U17985 (N_17985,N_17091,N_17317);
nand U17986 (N_17986,N_17404,N_17287);
xnor U17987 (N_17987,N_17424,N_17251);
and U17988 (N_17988,N_17323,N_17179);
xnor U17989 (N_17989,N_17451,N_17210);
or U17990 (N_17990,N_17100,N_17387);
nor U17991 (N_17991,N_17181,N_17328);
nand U17992 (N_17992,N_17319,N_17078);
or U17993 (N_17993,N_17221,N_17354);
or U17994 (N_17994,N_17102,N_17211);
and U17995 (N_17995,N_17422,N_17247);
nor U17996 (N_17996,N_17443,N_17047);
or U17997 (N_17997,N_17425,N_17349);
nor U17998 (N_17998,N_17099,N_17311);
or U17999 (N_17999,N_17035,N_17329);
nor U18000 (N_18000,N_17870,N_17505);
nor U18001 (N_18001,N_17747,N_17941);
and U18002 (N_18002,N_17990,N_17985);
nor U18003 (N_18003,N_17520,N_17576);
xor U18004 (N_18004,N_17541,N_17709);
or U18005 (N_18005,N_17866,N_17641);
or U18006 (N_18006,N_17906,N_17827);
or U18007 (N_18007,N_17713,N_17819);
xnor U18008 (N_18008,N_17804,N_17968);
and U18009 (N_18009,N_17569,N_17605);
or U18010 (N_18010,N_17835,N_17892);
or U18011 (N_18011,N_17664,N_17663);
or U18012 (N_18012,N_17573,N_17696);
nand U18013 (N_18013,N_17585,N_17869);
nand U18014 (N_18014,N_17519,N_17853);
and U18015 (N_18015,N_17679,N_17843);
nand U18016 (N_18016,N_17547,N_17572);
and U18017 (N_18017,N_17518,N_17983);
or U18018 (N_18018,N_17535,N_17953);
nand U18019 (N_18019,N_17807,N_17739);
nand U18020 (N_18020,N_17741,N_17684);
nand U18021 (N_18021,N_17754,N_17859);
xnor U18022 (N_18022,N_17829,N_17860);
xnor U18023 (N_18023,N_17513,N_17634);
xnor U18024 (N_18024,N_17961,N_17975);
nor U18025 (N_18025,N_17994,N_17918);
xor U18026 (N_18026,N_17948,N_17742);
nor U18027 (N_18027,N_17915,N_17920);
nand U18028 (N_18028,N_17735,N_17743);
xor U18029 (N_18029,N_17856,N_17562);
and U18030 (N_18030,N_17897,N_17740);
xnor U18031 (N_18031,N_17933,N_17507);
or U18032 (N_18032,N_17607,N_17960);
xnor U18033 (N_18033,N_17723,N_17658);
nand U18034 (N_18034,N_17724,N_17595);
or U18035 (N_18035,N_17616,N_17511);
xnor U18036 (N_18036,N_17579,N_17707);
xor U18037 (N_18037,N_17722,N_17534);
or U18038 (N_18038,N_17670,N_17524);
nor U18039 (N_18039,N_17622,N_17639);
nor U18040 (N_18040,N_17976,N_17563);
and U18041 (N_18041,N_17659,N_17732);
xor U18042 (N_18042,N_17868,N_17863);
xnor U18043 (N_18043,N_17940,N_17686);
and U18044 (N_18044,N_17700,N_17597);
xnor U18045 (N_18045,N_17927,N_17858);
and U18046 (N_18046,N_17554,N_17956);
or U18047 (N_18047,N_17556,N_17626);
nor U18048 (N_18048,N_17662,N_17525);
xor U18049 (N_18049,N_17553,N_17677);
xnor U18050 (N_18050,N_17673,N_17877);
nand U18051 (N_18051,N_17533,N_17705);
nand U18052 (N_18052,N_17529,N_17881);
xnor U18053 (N_18053,N_17545,N_17672);
nand U18054 (N_18054,N_17586,N_17760);
nand U18055 (N_18055,N_17795,N_17557);
nor U18056 (N_18056,N_17652,N_17980);
and U18057 (N_18057,N_17773,N_17687);
nand U18058 (N_18058,N_17911,N_17901);
and U18059 (N_18059,N_17884,N_17781);
nand U18060 (N_18060,N_17988,N_17594);
xnor U18061 (N_18061,N_17889,N_17637);
and U18062 (N_18062,N_17744,N_17548);
or U18063 (N_18063,N_17671,N_17708);
nor U18064 (N_18064,N_17631,N_17796);
and U18065 (N_18065,N_17717,N_17864);
and U18066 (N_18066,N_17890,N_17522);
nand U18067 (N_18067,N_17598,N_17971);
or U18068 (N_18068,N_17674,N_17935);
xor U18069 (N_18069,N_17734,N_17720);
or U18070 (N_18070,N_17582,N_17934);
nor U18071 (N_18071,N_17831,N_17731);
xor U18072 (N_18072,N_17632,N_17846);
nand U18073 (N_18073,N_17924,N_17624);
nand U18074 (N_18074,N_17617,N_17521);
nand U18075 (N_18075,N_17504,N_17957);
nand U18076 (N_18076,N_17803,N_17715);
nor U18077 (N_18077,N_17840,N_17876);
xor U18078 (N_18078,N_17822,N_17502);
and U18079 (N_18079,N_17602,N_17613);
nor U18080 (N_18080,N_17660,N_17729);
and U18081 (N_18081,N_17748,N_17694);
and U18082 (N_18082,N_17818,N_17949);
and U18083 (N_18083,N_17759,N_17922);
or U18084 (N_18084,N_17931,N_17647);
nand U18085 (N_18085,N_17855,N_17575);
xor U18086 (N_18086,N_17643,N_17566);
nor U18087 (N_18087,N_17791,N_17805);
nor U18088 (N_18088,N_17978,N_17973);
nand U18089 (N_18089,N_17813,N_17873);
or U18090 (N_18090,N_17792,N_17947);
or U18091 (N_18091,N_17746,N_17838);
xnor U18092 (N_18092,N_17712,N_17645);
nor U18093 (N_18093,N_17536,N_17900);
and U18094 (N_18094,N_17955,N_17825);
and U18095 (N_18095,N_17726,N_17691);
xnor U18096 (N_18096,N_17560,N_17779);
xnor U18097 (N_18097,N_17527,N_17736);
and U18098 (N_18098,N_17550,N_17703);
or U18099 (N_18099,N_17806,N_17763);
nand U18100 (N_18100,N_17718,N_17991);
nand U18101 (N_18101,N_17689,N_17730);
and U18102 (N_18102,N_17903,N_17714);
nor U18103 (N_18103,N_17651,N_17638);
nand U18104 (N_18104,N_17826,N_17999);
and U18105 (N_18105,N_17800,N_17907);
nor U18106 (N_18106,N_17783,N_17894);
and U18107 (N_18107,N_17899,N_17842);
nand U18108 (N_18108,N_17830,N_17503);
and U18109 (N_18109,N_17644,N_17697);
or U18110 (N_18110,N_17762,N_17501);
nand U18111 (N_18111,N_17801,N_17775);
nand U18112 (N_18112,N_17623,N_17681);
or U18113 (N_18113,N_17666,N_17844);
and U18114 (N_18114,N_17725,N_17516);
and U18115 (N_18115,N_17621,N_17833);
nand U18116 (N_18116,N_17539,N_17642);
and U18117 (N_18117,N_17929,N_17570);
nand U18118 (N_18118,N_17625,N_17802);
nor U18119 (N_18119,N_17909,N_17517);
nand U18120 (N_18120,N_17727,N_17815);
nor U18121 (N_18121,N_17981,N_17510);
nor U18122 (N_18122,N_17657,N_17636);
xnor U18123 (N_18123,N_17710,N_17782);
or U18124 (N_18124,N_17883,N_17698);
nand U18125 (N_18125,N_17584,N_17982);
xor U18126 (N_18126,N_17794,N_17635);
nor U18127 (N_18127,N_17919,N_17808);
xor U18128 (N_18128,N_17962,N_17603);
or U18129 (N_18129,N_17615,N_17926);
nor U18130 (N_18130,N_17544,N_17841);
nand U18131 (N_18131,N_17568,N_17711);
xnor U18132 (N_18132,N_17606,N_17506);
and U18133 (N_18133,N_17737,N_17761);
and U18134 (N_18134,N_17852,N_17910);
xnor U18135 (N_18135,N_17704,N_17969);
nor U18136 (N_18136,N_17649,N_17977);
and U18137 (N_18137,N_17604,N_17619);
and U18138 (N_18138,N_17882,N_17862);
nand U18139 (N_18139,N_17596,N_17721);
or U18140 (N_18140,N_17942,N_17778);
xnor U18141 (N_18141,N_17581,N_17787);
and U18142 (N_18142,N_17656,N_17592);
nand U18143 (N_18143,N_17848,N_17850);
nand U18144 (N_18144,N_17515,N_17546);
nand U18145 (N_18145,N_17701,N_17967);
nand U18146 (N_18146,N_17667,N_17514);
or U18147 (N_18147,N_17765,N_17610);
or U18148 (N_18148,N_17512,N_17893);
xor U18149 (N_18149,N_17790,N_17532);
xnor U18150 (N_18150,N_17683,N_17758);
or U18151 (N_18151,N_17950,N_17832);
and U18152 (N_18152,N_17680,N_17745);
or U18153 (N_18153,N_17963,N_17688);
xnor U18154 (N_18154,N_17865,N_17574);
or U18155 (N_18155,N_17665,N_17542);
and U18156 (N_18156,N_17784,N_17912);
xnor U18157 (N_18157,N_17676,N_17917);
and U18158 (N_18158,N_17526,N_17706);
xnor U18159 (N_18159,N_17809,N_17530);
and U18160 (N_18160,N_17549,N_17836);
or U18161 (N_18161,N_17875,N_17757);
or U18162 (N_18162,N_17943,N_17817);
and U18163 (N_18163,N_17690,N_17814);
xor U18164 (N_18164,N_17799,N_17620);
nor U18165 (N_18165,N_17768,N_17888);
or U18166 (N_18166,N_17733,N_17611);
xnor U18167 (N_18167,N_17945,N_17678);
nor U18168 (N_18168,N_17798,N_17923);
nor U18169 (N_18169,N_17954,N_17989);
nor U18170 (N_18170,N_17577,N_17552);
xnor U18171 (N_18171,N_17788,N_17880);
or U18172 (N_18172,N_17693,N_17685);
nor U18173 (N_18173,N_17851,N_17640);
and U18174 (N_18174,N_17908,N_17951);
or U18175 (N_18175,N_17528,N_17719);
and U18176 (N_18176,N_17543,N_17921);
nor U18177 (N_18177,N_17810,N_17992);
xor U18178 (N_18178,N_17823,N_17655);
or U18179 (N_18179,N_17555,N_17564);
or U18180 (N_18180,N_17902,N_17904);
and U18181 (N_18181,N_17702,N_17932);
xnor U18182 (N_18182,N_17580,N_17630);
nand U18183 (N_18183,N_17633,N_17936);
xor U18184 (N_18184,N_17692,N_17756);
or U18185 (N_18185,N_17561,N_17571);
nand U18186 (N_18186,N_17590,N_17699);
nand U18187 (N_18187,N_17587,N_17668);
nor U18188 (N_18188,N_17966,N_17793);
and U18189 (N_18189,N_17669,N_17627);
xnor U18190 (N_18190,N_17837,N_17872);
nand U18191 (N_18191,N_17772,N_17895);
nor U18192 (N_18192,N_17523,N_17970);
xor U18193 (N_18193,N_17538,N_17834);
xnor U18194 (N_18194,N_17599,N_17608);
nor U18195 (N_18195,N_17753,N_17738);
nor U18196 (N_18196,N_17774,N_17540);
nor U18197 (N_18197,N_17972,N_17885);
and U18198 (N_18198,N_17979,N_17612);
xnor U18199 (N_18199,N_17776,N_17589);
nor U18200 (N_18200,N_17618,N_17786);
nand U18201 (N_18201,N_17509,N_17845);
or U18202 (N_18202,N_17661,N_17591);
and U18203 (N_18203,N_17946,N_17769);
and U18204 (N_18204,N_17752,N_17937);
and U18205 (N_18205,N_17887,N_17986);
or U18206 (N_18206,N_17916,N_17789);
xnor U18207 (N_18207,N_17811,N_17764);
nor U18208 (N_18208,N_17886,N_17675);
and U18209 (N_18209,N_17938,N_17770);
nand U18210 (N_18210,N_17974,N_17609);
xor U18211 (N_18211,N_17531,N_17558);
or U18212 (N_18212,N_17821,N_17614);
xor U18213 (N_18213,N_17998,N_17628);
nand U18214 (N_18214,N_17650,N_17785);
nand U18215 (N_18215,N_17944,N_17767);
nor U18216 (N_18216,N_17755,N_17648);
xor U18217 (N_18217,N_17993,N_17820);
or U18218 (N_18218,N_17849,N_17750);
nand U18219 (N_18219,N_17871,N_17824);
and U18220 (N_18220,N_17898,N_17896);
and U18221 (N_18221,N_17952,N_17984);
or U18222 (N_18222,N_17874,N_17653);
and U18223 (N_18223,N_17551,N_17600);
xnor U18224 (N_18224,N_17780,N_17508);
nand U18225 (N_18225,N_17925,N_17751);
nor U18226 (N_18226,N_17987,N_17559);
or U18227 (N_18227,N_17958,N_17995);
nor U18228 (N_18228,N_17861,N_17500);
nand U18229 (N_18229,N_17777,N_17965);
xor U18230 (N_18230,N_17928,N_17537);
and U18231 (N_18231,N_17867,N_17997);
xnor U18232 (N_18232,N_17749,N_17567);
and U18233 (N_18233,N_17695,N_17905);
nand U18234 (N_18234,N_17646,N_17914);
xnor U18235 (N_18235,N_17959,N_17879);
nor U18236 (N_18236,N_17878,N_17654);
xor U18237 (N_18237,N_17812,N_17939);
or U18238 (N_18238,N_17629,N_17728);
or U18239 (N_18239,N_17771,N_17716);
xor U18240 (N_18240,N_17797,N_17565);
or U18241 (N_18241,N_17601,N_17857);
xor U18242 (N_18242,N_17913,N_17847);
nor U18243 (N_18243,N_17588,N_17828);
and U18244 (N_18244,N_17854,N_17682);
nor U18245 (N_18245,N_17996,N_17816);
nor U18246 (N_18246,N_17583,N_17593);
or U18247 (N_18247,N_17766,N_17891);
and U18248 (N_18248,N_17578,N_17964);
and U18249 (N_18249,N_17930,N_17839);
or U18250 (N_18250,N_17562,N_17979);
or U18251 (N_18251,N_17769,N_17743);
nand U18252 (N_18252,N_17848,N_17839);
and U18253 (N_18253,N_17636,N_17917);
or U18254 (N_18254,N_17977,N_17948);
nor U18255 (N_18255,N_17990,N_17679);
nand U18256 (N_18256,N_17802,N_17518);
nor U18257 (N_18257,N_17874,N_17614);
nand U18258 (N_18258,N_17824,N_17583);
nand U18259 (N_18259,N_17965,N_17932);
xor U18260 (N_18260,N_17656,N_17914);
nor U18261 (N_18261,N_17722,N_17997);
xor U18262 (N_18262,N_17596,N_17558);
and U18263 (N_18263,N_17583,N_17708);
nand U18264 (N_18264,N_17926,N_17546);
and U18265 (N_18265,N_17838,N_17645);
or U18266 (N_18266,N_17996,N_17528);
or U18267 (N_18267,N_17965,N_17869);
xor U18268 (N_18268,N_17664,N_17768);
xor U18269 (N_18269,N_17927,N_17936);
nor U18270 (N_18270,N_17661,N_17756);
nand U18271 (N_18271,N_17853,N_17878);
or U18272 (N_18272,N_17657,N_17672);
xnor U18273 (N_18273,N_17525,N_17576);
nand U18274 (N_18274,N_17808,N_17620);
and U18275 (N_18275,N_17559,N_17867);
nand U18276 (N_18276,N_17750,N_17933);
nand U18277 (N_18277,N_17556,N_17719);
nor U18278 (N_18278,N_17874,N_17918);
or U18279 (N_18279,N_17661,N_17534);
nor U18280 (N_18280,N_17976,N_17784);
and U18281 (N_18281,N_17904,N_17966);
nand U18282 (N_18282,N_17592,N_17820);
or U18283 (N_18283,N_17728,N_17662);
xnor U18284 (N_18284,N_17982,N_17905);
xor U18285 (N_18285,N_17648,N_17868);
nor U18286 (N_18286,N_17962,N_17722);
xor U18287 (N_18287,N_17515,N_17795);
xor U18288 (N_18288,N_17535,N_17874);
or U18289 (N_18289,N_17667,N_17785);
nand U18290 (N_18290,N_17667,N_17787);
or U18291 (N_18291,N_17589,N_17822);
and U18292 (N_18292,N_17863,N_17581);
xnor U18293 (N_18293,N_17896,N_17717);
nand U18294 (N_18294,N_17879,N_17571);
or U18295 (N_18295,N_17704,N_17557);
or U18296 (N_18296,N_17711,N_17935);
nand U18297 (N_18297,N_17802,N_17952);
and U18298 (N_18298,N_17787,N_17738);
nor U18299 (N_18299,N_17916,N_17956);
and U18300 (N_18300,N_17511,N_17792);
or U18301 (N_18301,N_17960,N_17994);
nand U18302 (N_18302,N_17778,N_17691);
or U18303 (N_18303,N_17699,N_17712);
or U18304 (N_18304,N_17613,N_17900);
xnor U18305 (N_18305,N_17912,N_17857);
and U18306 (N_18306,N_17505,N_17696);
nor U18307 (N_18307,N_17949,N_17858);
and U18308 (N_18308,N_17708,N_17659);
nor U18309 (N_18309,N_17978,N_17886);
and U18310 (N_18310,N_17634,N_17651);
and U18311 (N_18311,N_17611,N_17667);
nand U18312 (N_18312,N_17969,N_17840);
or U18313 (N_18313,N_17636,N_17884);
xor U18314 (N_18314,N_17668,N_17841);
and U18315 (N_18315,N_17804,N_17720);
nor U18316 (N_18316,N_17921,N_17825);
nor U18317 (N_18317,N_17775,N_17914);
and U18318 (N_18318,N_17576,N_17906);
xor U18319 (N_18319,N_17672,N_17504);
nand U18320 (N_18320,N_17934,N_17608);
nor U18321 (N_18321,N_17718,N_17571);
xor U18322 (N_18322,N_17759,N_17527);
nand U18323 (N_18323,N_17614,N_17535);
nor U18324 (N_18324,N_17649,N_17768);
or U18325 (N_18325,N_17620,N_17741);
nand U18326 (N_18326,N_17889,N_17551);
xnor U18327 (N_18327,N_17899,N_17592);
nand U18328 (N_18328,N_17822,N_17718);
nand U18329 (N_18329,N_17886,N_17582);
nor U18330 (N_18330,N_17896,N_17653);
xor U18331 (N_18331,N_17786,N_17970);
nor U18332 (N_18332,N_17568,N_17917);
nor U18333 (N_18333,N_17960,N_17990);
nand U18334 (N_18334,N_17749,N_17711);
and U18335 (N_18335,N_17647,N_17603);
and U18336 (N_18336,N_17784,N_17524);
nor U18337 (N_18337,N_17693,N_17766);
xnor U18338 (N_18338,N_17939,N_17806);
nor U18339 (N_18339,N_17782,N_17818);
xor U18340 (N_18340,N_17534,N_17521);
and U18341 (N_18341,N_17710,N_17967);
nor U18342 (N_18342,N_17513,N_17749);
nor U18343 (N_18343,N_17780,N_17715);
nor U18344 (N_18344,N_17897,N_17913);
xnor U18345 (N_18345,N_17883,N_17739);
and U18346 (N_18346,N_17811,N_17665);
nor U18347 (N_18347,N_17784,N_17635);
or U18348 (N_18348,N_17784,N_17858);
and U18349 (N_18349,N_17842,N_17784);
and U18350 (N_18350,N_17555,N_17625);
nor U18351 (N_18351,N_17642,N_17862);
xnor U18352 (N_18352,N_17967,N_17979);
xnor U18353 (N_18353,N_17764,N_17895);
or U18354 (N_18354,N_17550,N_17662);
nand U18355 (N_18355,N_17635,N_17906);
or U18356 (N_18356,N_17787,N_17597);
and U18357 (N_18357,N_17833,N_17629);
xor U18358 (N_18358,N_17521,N_17728);
xor U18359 (N_18359,N_17629,N_17653);
or U18360 (N_18360,N_17735,N_17643);
nor U18361 (N_18361,N_17950,N_17959);
nor U18362 (N_18362,N_17707,N_17656);
or U18363 (N_18363,N_17679,N_17609);
nor U18364 (N_18364,N_17942,N_17535);
nand U18365 (N_18365,N_17814,N_17510);
nor U18366 (N_18366,N_17693,N_17914);
and U18367 (N_18367,N_17503,N_17629);
or U18368 (N_18368,N_17995,N_17913);
and U18369 (N_18369,N_17873,N_17505);
nand U18370 (N_18370,N_17833,N_17995);
xnor U18371 (N_18371,N_17958,N_17534);
and U18372 (N_18372,N_17788,N_17791);
nor U18373 (N_18373,N_17776,N_17542);
or U18374 (N_18374,N_17716,N_17537);
or U18375 (N_18375,N_17673,N_17634);
xor U18376 (N_18376,N_17637,N_17947);
nor U18377 (N_18377,N_17666,N_17978);
and U18378 (N_18378,N_17752,N_17909);
nor U18379 (N_18379,N_17767,N_17929);
nor U18380 (N_18380,N_17743,N_17943);
and U18381 (N_18381,N_17561,N_17933);
or U18382 (N_18382,N_17876,N_17746);
and U18383 (N_18383,N_17568,N_17894);
nand U18384 (N_18384,N_17736,N_17876);
xor U18385 (N_18385,N_17591,N_17761);
or U18386 (N_18386,N_17742,N_17555);
and U18387 (N_18387,N_17700,N_17611);
and U18388 (N_18388,N_17799,N_17511);
xnor U18389 (N_18389,N_17774,N_17521);
and U18390 (N_18390,N_17547,N_17921);
nor U18391 (N_18391,N_17811,N_17776);
nand U18392 (N_18392,N_17906,N_17640);
nand U18393 (N_18393,N_17550,N_17680);
nor U18394 (N_18394,N_17734,N_17586);
nand U18395 (N_18395,N_17742,N_17979);
nor U18396 (N_18396,N_17720,N_17929);
xor U18397 (N_18397,N_17897,N_17688);
nor U18398 (N_18398,N_17990,N_17839);
xnor U18399 (N_18399,N_17617,N_17832);
and U18400 (N_18400,N_17953,N_17921);
nor U18401 (N_18401,N_17774,N_17543);
xnor U18402 (N_18402,N_17828,N_17808);
and U18403 (N_18403,N_17758,N_17978);
or U18404 (N_18404,N_17879,N_17794);
nor U18405 (N_18405,N_17875,N_17761);
xnor U18406 (N_18406,N_17614,N_17563);
and U18407 (N_18407,N_17889,N_17812);
xnor U18408 (N_18408,N_17991,N_17840);
nand U18409 (N_18409,N_17669,N_17584);
nand U18410 (N_18410,N_17558,N_17524);
and U18411 (N_18411,N_17812,N_17716);
and U18412 (N_18412,N_17760,N_17862);
and U18413 (N_18413,N_17599,N_17615);
nand U18414 (N_18414,N_17705,N_17831);
nand U18415 (N_18415,N_17547,N_17579);
and U18416 (N_18416,N_17704,N_17844);
and U18417 (N_18417,N_17675,N_17609);
nand U18418 (N_18418,N_17571,N_17956);
nor U18419 (N_18419,N_17704,N_17508);
xnor U18420 (N_18420,N_17663,N_17543);
or U18421 (N_18421,N_17609,N_17793);
xnor U18422 (N_18422,N_17519,N_17609);
xor U18423 (N_18423,N_17527,N_17639);
nor U18424 (N_18424,N_17730,N_17657);
nor U18425 (N_18425,N_17616,N_17673);
or U18426 (N_18426,N_17965,N_17723);
nor U18427 (N_18427,N_17753,N_17518);
and U18428 (N_18428,N_17926,N_17985);
and U18429 (N_18429,N_17832,N_17926);
or U18430 (N_18430,N_17609,N_17977);
and U18431 (N_18431,N_17623,N_17737);
xor U18432 (N_18432,N_17763,N_17914);
and U18433 (N_18433,N_17645,N_17964);
nor U18434 (N_18434,N_17974,N_17502);
xor U18435 (N_18435,N_17562,N_17983);
and U18436 (N_18436,N_17580,N_17548);
or U18437 (N_18437,N_17611,N_17897);
or U18438 (N_18438,N_17757,N_17888);
or U18439 (N_18439,N_17516,N_17639);
nand U18440 (N_18440,N_17711,N_17744);
or U18441 (N_18441,N_17993,N_17702);
or U18442 (N_18442,N_17680,N_17835);
nor U18443 (N_18443,N_17710,N_17847);
xor U18444 (N_18444,N_17595,N_17934);
nand U18445 (N_18445,N_17951,N_17845);
nor U18446 (N_18446,N_17516,N_17535);
or U18447 (N_18447,N_17541,N_17824);
and U18448 (N_18448,N_17719,N_17858);
or U18449 (N_18449,N_17786,N_17680);
nor U18450 (N_18450,N_17944,N_17760);
and U18451 (N_18451,N_17656,N_17815);
and U18452 (N_18452,N_17772,N_17936);
nor U18453 (N_18453,N_17846,N_17727);
xor U18454 (N_18454,N_17700,N_17673);
xnor U18455 (N_18455,N_17651,N_17763);
or U18456 (N_18456,N_17859,N_17692);
or U18457 (N_18457,N_17810,N_17827);
nor U18458 (N_18458,N_17949,N_17926);
nor U18459 (N_18459,N_17641,N_17832);
xor U18460 (N_18460,N_17512,N_17748);
and U18461 (N_18461,N_17993,N_17596);
xor U18462 (N_18462,N_17663,N_17755);
and U18463 (N_18463,N_17607,N_17740);
or U18464 (N_18464,N_17704,N_17919);
nor U18465 (N_18465,N_17647,N_17830);
xnor U18466 (N_18466,N_17663,N_17935);
and U18467 (N_18467,N_17593,N_17508);
nand U18468 (N_18468,N_17703,N_17567);
nand U18469 (N_18469,N_17850,N_17962);
nand U18470 (N_18470,N_17850,N_17918);
xor U18471 (N_18471,N_17583,N_17780);
nand U18472 (N_18472,N_17880,N_17592);
and U18473 (N_18473,N_17542,N_17863);
or U18474 (N_18474,N_17837,N_17718);
and U18475 (N_18475,N_17635,N_17668);
and U18476 (N_18476,N_17840,N_17537);
nand U18477 (N_18477,N_17694,N_17988);
and U18478 (N_18478,N_17617,N_17911);
nor U18479 (N_18479,N_17640,N_17691);
and U18480 (N_18480,N_17563,N_17946);
and U18481 (N_18481,N_17753,N_17763);
or U18482 (N_18482,N_17727,N_17587);
xnor U18483 (N_18483,N_17838,N_17845);
xnor U18484 (N_18484,N_17936,N_17588);
or U18485 (N_18485,N_17733,N_17594);
nand U18486 (N_18486,N_17512,N_17574);
xor U18487 (N_18487,N_17922,N_17854);
xor U18488 (N_18488,N_17721,N_17896);
nor U18489 (N_18489,N_17656,N_17509);
or U18490 (N_18490,N_17658,N_17922);
xor U18491 (N_18491,N_17601,N_17591);
nand U18492 (N_18492,N_17881,N_17915);
nand U18493 (N_18493,N_17503,N_17739);
nand U18494 (N_18494,N_17814,N_17816);
or U18495 (N_18495,N_17861,N_17905);
or U18496 (N_18496,N_17544,N_17925);
or U18497 (N_18497,N_17652,N_17561);
and U18498 (N_18498,N_17738,N_17964);
or U18499 (N_18499,N_17829,N_17500);
and U18500 (N_18500,N_18456,N_18159);
or U18501 (N_18501,N_18006,N_18360);
nand U18502 (N_18502,N_18478,N_18134);
nand U18503 (N_18503,N_18171,N_18352);
nand U18504 (N_18504,N_18147,N_18344);
nor U18505 (N_18505,N_18135,N_18066);
or U18506 (N_18506,N_18272,N_18407);
nor U18507 (N_18507,N_18174,N_18454);
xnor U18508 (N_18508,N_18137,N_18323);
nand U18509 (N_18509,N_18379,N_18363);
and U18510 (N_18510,N_18370,N_18394);
and U18511 (N_18511,N_18179,N_18103);
and U18512 (N_18512,N_18414,N_18030);
xnor U18513 (N_18513,N_18497,N_18464);
and U18514 (N_18514,N_18098,N_18012);
nor U18515 (N_18515,N_18243,N_18242);
xnor U18516 (N_18516,N_18383,N_18452);
nand U18517 (N_18517,N_18451,N_18225);
nor U18518 (N_18518,N_18120,N_18266);
xnor U18519 (N_18519,N_18300,N_18298);
nand U18520 (N_18520,N_18093,N_18447);
nor U18521 (N_18521,N_18201,N_18138);
nor U18522 (N_18522,N_18273,N_18020);
nand U18523 (N_18523,N_18484,N_18355);
nand U18524 (N_18524,N_18269,N_18264);
xnor U18525 (N_18525,N_18037,N_18393);
xnor U18526 (N_18526,N_18167,N_18359);
and U18527 (N_18527,N_18309,N_18153);
xnor U18528 (N_18528,N_18458,N_18079);
or U18529 (N_18529,N_18113,N_18307);
or U18530 (N_18530,N_18249,N_18475);
nand U18531 (N_18531,N_18114,N_18165);
nand U18532 (N_18532,N_18178,N_18241);
and U18533 (N_18533,N_18354,N_18263);
nand U18534 (N_18534,N_18110,N_18317);
and U18535 (N_18535,N_18450,N_18202);
nand U18536 (N_18536,N_18122,N_18372);
nand U18537 (N_18537,N_18169,N_18400);
xor U18538 (N_18538,N_18074,N_18423);
nand U18539 (N_18539,N_18205,N_18286);
xor U18540 (N_18540,N_18231,N_18189);
or U18541 (N_18541,N_18401,N_18318);
xor U18542 (N_18542,N_18373,N_18163);
nand U18543 (N_18543,N_18488,N_18190);
xnor U18544 (N_18544,N_18402,N_18118);
nor U18545 (N_18545,N_18059,N_18463);
nand U18546 (N_18546,N_18109,N_18397);
xnor U18547 (N_18547,N_18365,N_18092);
nor U18548 (N_18548,N_18084,N_18388);
xnor U18549 (N_18549,N_18429,N_18026);
and U18550 (N_18550,N_18117,N_18290);
or U18551 (N_18551,N_18455,N_18405);
nor U18552 (N_18552,N_18005,N_18196);
nand U18553 (N_18553,N_18029,N_18040);
or U18554 (N_18554,N_18177,N_18068);
nand U18555 (N_18555,N_18374,N_18157);
and U18556 (N_18556,N_18016,N_18297);
xor U18557 (N_18557,N_18268,N_18440);
nor U18558 (N_18558,N_18461,N_18391);
nand U18559 (N_18559,N_18337,N_18238);
nand U18560 (N_18560,N_18237,N_18282);
and U18561 (N_18561,N_18426,N_18121);
or U18562 (N_18562,N_18472,N_18421);
xor U18563 (N_18563,N_18413,N_18267);
nand U18564 (N_18564,N_18041,N_18380);
nand U18565 (N_18565,N_18403,N_18050);
nand U18566 (N_18566,N_18070,N_18442);
and U18567 (N_18567,N_18180,N_18351);
or U18568 (N_18568,N_18244,N_18090);
nand U18569 (N_18569,N_18141,N_18449);
nand U18570 (N_18570,N_18161,N_18187);
nor U18571 (N_18571,N_18197,N_18411);
and U18572 (N_18572,N_18001,N_18130);
xor U18573 (N_18573,N_18253,N_18132);
nor U18574 (N_18574,N_18233,N_18228);
xor U18575 (N_18575,N_18462,N_18281);
nor U18576 (N_18576,N_18493,N_18014);
xnor U18577 (N_18577,N_18047,N_18367);
or U18578 (N_18578,N_18437,N_18473);
nor U18579 (N_18579,N_18482,N_18034);
xor U18580 (N_18580,N_18312,N_18203);
nand U18581 (N_18581,N_18129,N_18075);
nand U18582 (N_18582,N_18369,N_18191);
nor U18583 (N_18583,N_18424,N_18319);
xor U18584 (N_18584,N_18051,N_18025);
or U18585 (N_18585,N_18055,N_18158);
and U18586 (N_18586,N_18427,N_18305);
xnor U18587 (N_18587,N_18230,N_18096);
or U18588 (N_18588,N_18459,N_18448);
and U18589 (N_18589,N_18313,N_18303);
xnor U18590 (N_18590,N_18322,N_18293);
xor U18591 (N_18591,N_18353,N_18058);
nor U18592 (N_18592,N_18328,N_18087);
or U18593 (N_18593,N_18152,N_18491);
nand U18594 (N_18594,N_18222,N_18049);
nor U18595 (N_18595,N_18010,N_18035);
and U18596 (N_18596,N_18236,N_18387);
or U18597 (N_18597,N_18218,N_18311);
xor U18598 (N_18598,N_18435,N_18284);
and U18599 (N_18599,N_18494,N_18368);
and U18600 (N_18600,N_18386,N_18061);
and U18601 (N_18601,N_18406,N_18127);
nand U18602 (N_18602,N_18036,N_18358);
nor U18603 (N_18603,N_18404,N_18495);
and U18604 (N_18604,N_18211,N_18065);
and U18605 (N_18605,N_18457,N_18162);
and U18606 (N_18606,N_18071,N_18396);
nor U18607 (N_18607,N_18057,N_18033);
nor U18608 (N_18608,N_18215,N_18356);
nor U18609 (N_18609,N_18166,N_18257);
nand U18610 (N_18610,N_18335,N_18466);
or U18611 (N_18611,N_18198,N_18206);
or U18612 (N_18612,N_18314,N_18086);
nand U18613 (N_18613,N_18479,N_18143);
nand U18614 (N_18614,N_18334,N_18106);
nand U18615 (N_18615,N_18139,N_18185);
or U18616 (N_18616,N_18279,N_18056);
or U18617 (N_18617,N_18195,N_18155);
nor U18618 (N_18618,N_18046,N_18333);
nor U18619 (N_18619,N_18390,N_18348);
or U18620 (N_18620,N_18140,N_18392);
xnor U18621 (N_18621,N_18389,N_18436);
or U18622 (N_18622,N_18486,N_18149);
and U18623 (N_18623,N_18219,N_18043);
xor U18624 (N_18624,N_18485,N_18200);
xor U18625 (N_18625,N_18376,N_18441);
and U18626 (N_18626,N_18416,N_18271);
nand U18627 (N_18627,N_18326,N_18146);
and U18628 (N_18628,N_18007,N_18095);
nor U18629 (N_18629,N_18002,N_18277);
nor U18630 (N_18630,N_18256,N_18038);
nor U18631 (N_18631,N_18013,N_18168);
nor U18632 (N_18632,N_18192,N_18476);
or U18633 (N_18633,N_18347,N_18213);
or U18634 (N_18634,N_18062,N_18338);
or U18635 (N_18635,N_18142,N_18252);
or U18636 (N_18636,N_18063,N_18151);
xor U18637 (N_18637,N_18060,N_18112);
xnor U18638 (N_18638,N_18176,N_18115);
nor U18639 (N_18639,N_18227,N_18150);
nor U18640 (N_18640,N_18052,N_18496);
nand U18641 (N_18641,N_18069,N_18193);
or U18642 (N_18642,N_18255,N_18321);
and U18643 (N_18643,N_18144,N_18015);
or U18644 (N_18644,N_18415,N_18164);
nand U18645 (N_18645,N_18432,N_18209);
nand U18646 (N_18646,N_18417,N_18245);
nand U18647 (N_18647,N_18409,N_18136);
nand U18648 (N_18648,N_18100,N_18102);
or U18649 (N_18649,N_18097,N_18310);
or U18650 (N_18650,N_18430,N_18124);
xor U18651 (N_18651,N_18184,N_18294);
xor U18652 (N_18652,N_18011,N_18316);
nor U18653 (N_18653,N_18287,N_18104);
and U18654 (N_18654,N_18131,N_18123);
xor U18655 (N_18655,N_18031,N_18304);
nor U18656 (N_18656,N_18042,N_18341);
nand U18657 (N_18657,N_18172,N_18289);
nand U18658 (N_18658,N_18003,N_18082);
or U18659 (N_18659,N_18221,N_18385);
nand U18660 (N_18660,N_18039,N_18072);
and U18661 (N_18661,N_18296,N_18081);
xor U18662 (N_18662,N_18349,N_18258);
xor U18663 (N_18663,N_18381,N_18499);
xor U18664 (N_18664,N_18412,N_18028);
nand U18665 (N_18665,N_18160,N_18469);
xor U18666 (N_18666,N_18226,N_18019);
xnor U18667 (N_18667,N_18073,N_18308);
xnor U18668 (N_18668,N_18483,N_18364);
or U18669 (N_18669,N_18302,N_18023);
or U18670 (N_18670,N_18301,N_18418);
nor U18671 (N_18671,N_18467,N_18422);
or U18672 (N_18672,N_18292,N_18306);
nand U18673 (N_18673,N_18325,N_18280);
nor U18674 (N_18674,N_18453,N_18246);
nand U18675 (N_18675,N_18339,N_18145);
or U18676 (N_18676,N_18021,N_18017);
and U18677 (N_18677,N_18089,N_18235);
and U18678 (N_18678,N_18384,N_18077);
or U18679 (N_18679,N_18288,N_18199);
nor U18680 (N_18680,N_18125,N_18000);
and U18681 (N_18681,N_18234,N_18446);
nor U18682 (N_18682,N_18330,N_18259);
xnor U18683 (N_18683,N_18399,N_18324);
nand U18684 (N_18684,N_18091,N_18439);
nand U18685 (N_18685,N_18067,N_18248);
nand U18686 (N_18686,N_18471,N_18220);
or U18687 (N_18687,N_18343,N_18101);
xor U18688 (N_18688,N_18395,N_18420);
xnor U18689 (N_18689,N_18076,N_18480);
or U18690 (N_18690,N_18044,N_18156);
nand U18691 (N_18691,N_18239,N_18275);
nor U18692 (N_18692,N_18377,N_18444);
xnor U18693 (N_18693,N_18329,N_18299);
or U18694 (N_18694,N_18240,N_18274);
or U18695 (N_18695,N_18465,N_18229);
nand U18696 (N_18696,N_18004,N_18080);
xnor U18697 (N_18697,N_18489,N_18078);
xor U18698 (N_18698,N_18382,N_18018);
and U18699 (N_18699,N_18265,N_18278);
and U18700 (N_18700,N_18408,N_18182);
or U18701 (N_18701,N_18350,N_18470);
nor U18702 (N_18702,N_18260,N_18434);
nor U18703 (N_18703,N_18154,N_18232);
xor U18704 (N_18704,N_18094,N_18361);
or U18705 (N_18705,N_18492,N_18291);
nor U18706 (N_18706,N_18216,N_18487);
xnor U18707 (N_18707,N_18208,N_18194);
and U18708 (N_18708,N_18261,N_18445);
or U18709 (N_18709,N_18099,N_18210);
nor U18710 (N_18710,N_18217,N_18204);
nor U18711 (N_18711,N_18214,N_18477);
and U18712 (N_18712,N_18188,N_18468);
nand U18713 (N_18713,N_18366,N_18064);
xor U18714 (N_18714,N_18250,N_18024);
nand U18715 (N_18715,N_18083,N_18419);
nand U18716 (N_18716,N_18223,N_18254);
and U18717 (N_18717,N_18285,N_18276);
xor U18718 (N_18718,N_18342,N_18170);
xnor U18719 (N_18719,N_18148,N_18357);
nand U18720 (N_18720,N_18498,N_18048);
or U18721 (N_18721,N_18022,N_18428);
or U18722 (N_18722,N_18331,N_18362);
and U18723 (N_18723,N_18398,N_18105);
and U18724 (N_18724,N_18175,N_18490);
or U18725 (N_18725,N_18433,N_18128);
and U18726 (N_18726,N_18460,N_18481);
or U18727 (N_18727,N_18346,N_18251);
xnor U18728 (N_18728,N_18410,N_18053);
or U18729 (N_18729,N_18207,N_18247);
nor U18730 (N_18730,N_18371,N_18133);
and U18731 (N_18731,N_18332,N_18181);
or U18732 (N_18732,N_18425,N_18431);
and U18733 (N_18733,N_18224,N_18111);
nand U18734 (N_18734,N_18262,N_18126);
and U18735 (N_18735,N_18088,N_18008);
or U18736 (N_18736,N_18045,N_18378);
or U18737 (N_18737,N_18027,N_18032);
and U18738 (N_18738,N_18054,N_18212);
xnor U18739 (N_18739,N_18116,N_18336);
nor U18740 (N_18740,N_18085,N_18438);
xor U18741 (N_18741,N_18345,N_18009);
or U18742 (N_18742,N_18327,N_18186);
nand U18743 (N_18743,N_18283,N_18474);
and U18744 (N_18744,N_18119,N_18270);
xor U18745 (N_18745,N_18315,N_18107);
and U18746 (N_18746,N_18183,N_18295);
nor U18747 (N_18747,N_18340,N_18173);
xor U18748 (N_18748,N_18443,N_18320);
and U18749 (N_18749,N_18108,N_18375);
xnor U18750 (N_18750,N_18032,N_18146);
nor U18751 (N_18751,N_18178,N_18085);
or U18752 (N_18752,N_18377,N_18127);
xor U18753 (N_18753,N_18266,N_18319);
and U18754 (N_18754,N_18341,N_18405);
or U18755 (N_18755,N_18239,N_18475);
or U18756 (N_18756,N_18125,N_18466);
or U18757 (N_18757,N_18407,N_18362);
and U18758 (N_18758,N_18391,N_18337);
nor U18759 (N_18759,N_18147,N_18419);
nand U18760 (N_18760,N_18035,N_18112);
or U18761 (N_18761,N_18157,N_18072);
xor U18762 (N_18762,N_18166,N_18476);
xor U18763 (N_18763,N_18378,N_18383);
nor U18764 (N_18764,N_18068,N_18231);
and U18765 (N_18765,N_18147,N_18452);
nor U18766 (N_18766,N_18232,N_18119);
xnor U18767 (N_18767,N_18480,N_18349);
nor U18768 (N_18768,N_18007,N_18253);
nand U18769 (N_18769,N_18292,N_18282);
xor U18770 (N_18770,N_18343,N_18032);
nand U18771 (N_18771,N_18249,N_18323);
xor U18772 (N_18772,N_18055,N_18418);
and U18773 (N_18773,N_18414,N_18096);
nand U18774 (N_18774,N_18471,N_18200);
nor U18775 (N_18775,N_18407,N_18337);
nand U18776 (N_18776,N_18335,N_18247);
or U18777 (N_18777,N_18315,N_18266);
nand U18778 (N_18778,N_18068,N_18028);
or U18779 (N_18779,N_18018,N_18238);
xor U18780 (N_18780,N_18383,N_18322);
or U18781 (N_18781,N_18268,N_18023);
or U18782 (N_18782,N_18324,N_18047);
and U18783 (N_18783,N_18249,N_18151);
xor U18784 (N_18784,N_18421,N_18145);
nand U18785 (N_18785,N_18287,N_18203);
nor U18786 (N_18786,N_18326,N_18411);
nand U18787 (N_18787,N_18481,N_18196);
nand U18788 (N_18788,N_18325,N_18360);
and U18789 (N_18789,N_18479,N_18343);
xor U18790 (N_18790,N_18314,N_18486);
nand U18791 (N_18791,N_18380,N_18179);
xor U18792 (N_18792,N_18151,N_18174);
and U18793 (N_18793,N_18061,N_18107);
xor U18794 (N_18794,N_18409,N_18189);
or U18795 (N_18795,N_18025,N_18248);
xor U18796 (N_18796,N_18097,N_18419);
xor U18797 (N_18797,N_18063,N_18266);
xor U18798 (N_18798,N_18058,N_18376);
nand U18799 (N_18799,N_18312,N_18309);
and U18800 (N_18800,N_18131,N_18354);
or U18801 (N_18801,N_18077,N_18498);
nand U18802 (N_18802,N_18198,N_18360);
or U18803 (N_18803,N_18003,N_18381);
or U18804 (N_18804,N_18080,N_18495);
and U18805 (N_18805,N_18330,N_18106);
nor U18806 (N_18806,N_18309,N_18307);
and U18807 (N_18807,N_18062,N_18461);
xnor U18808 (N_18808,N_18145,N_18252);
nor U18809 (N_18809,N_18040,N_18080);
nor U18810 (N_18810,N_18187,N_18090);
nor U18811 (N_18811,N_18033,N_18301);
and U18812 (N_18812,N_18016,N_18296);
nand U18813 (N_18813,N_18462,N_18155);
and U18814 (N_18814,N_18390,N_18213);
and U18815 (N_18815,N_18290,N_18353);
xor U18816 (N_18816,N_18328,N_18132);
xnor U18817 (N_18817,N_18486,N_18435);
nand U18818 (N_18818,N_18493,N_18166);
nand U18819 (N_18819,N_18256,N_18416);
nand U18820 (N_18820,N_18252,N_18428);
xor U18821 (N_18821,N_18303,N_18043);
and U18822 (N_18822,N_18490,N_18173);
xnor U18823 (N_18823,N_18341,N_18097);
or U18824 (N_18824,N_18196,N_18369);
nand U18825 (N_18825,N_18476,N_18205);
and U18826 (N_18826,N_18103,N_18478);
nand U18827 (N_18827,N_18357,N_18334);
or U18828 (N_18828,N_18018,N_18399);
nand U18829 (N_18829,N_18169,N_18367);
nand U18830 (N_18830,N_18206,N_18055);
and U18831 (N_18831,N_18057,N_18492);
nor U18832 (N_18832,N_18303,N_18062);
nand U18833 (N_18833,N_18348,N_18041);
xnor U18834 (N_18834,N_18219,N_18028);
and U18835 (N_18835,N_18233,N_18264);
and U18836 (N_18836,N_18102,N_18057);
nor U18837 (N_18837,N_18056,N_18409);
nor U18838 (N_18838,N_18144,N_18121);
and U18839 (N_18839,N_18046,N_18135);
nand U18840 (N_18840,N_18221,N_18493);
and U18841 (N_18841,N_18371,N_18375);
xnor U18842 (N_18842,N_18121,N_18196);
xor U18843 (N_18843,N_18295,N_18419);
nor U18844 (N_18844,N_18321,N_18305);
and U18845 (N_18845,N_18002,N_18000);
and U18846 (N_18846,N_18477,N_18147);
or U18847 (N_18847,N_18158,N_18130);
and U18848 (N_18848,N_18210,N_18188);
and U18849 (N_18849,N_18459,N_18100);
and U18850 (N_18850,N_18204,N_18117);
or U18851 (N_18851,N_18351,N_18310);
nand U18852 (N_18852,N_18138,N_18092);
nand U18853 (N_18853,N_18283,N_18039);
xor U18854 (N_18854,N_18272,N_18241);
or U18855 (N_18855,N_18256,N_18410);
nor U18856 (N_18856,N_18126,N_18281);
or U18857 (N_18857,N_18116,N_18192);
or U18858 (N_18858,N_18124,N_18303);
nor U18859 (N_18859,N_18443,N_18258);
or U18860 (N_18860,N_18081,N_18138);
and U18861 (N_18861,N_18402,N_18384);
nand U18862 (N_18862,N_18395,N_18362);
nand U18863 (N_18863,N_18467,N_18326);
nand U18864 (N_18864,N_18416,N_18094);
xnor U18865 (N_18865,N_18118,N_18442);
nor U18866 (N_18866,N_18183,N_18466);
nand U18867 (N_18867,N_18334,N_18111);
nand U18868 (N_18868,N_18426,N_18169);
nor U18869 (N_18869,N_18342,N_18358);
nand U18870 (N_18870,N_18159,N_18413);
or U18871 (N_18871,N_18011,N_18360);
and U18872 (N_18872,N_18097,N_18259);
and U18873 (N_18873,N_18416,N_18211);
nor U18874 (N_18874,N_18233,N_18241);
nor U18875 (N_18875,N_18085,N_18202);
nor U18876 (N_18876,N_18455,N_18198);
and U18877 (N_18877,N_18221,N_18367);
xor U18878 (N_18878,N_18455,N_18287);
nand U18879 (N_18879,N_18472,N_18387);
xor U18880 (N_18880,N_18454,N_18120);
and U18881 (N_18881,N_18440,N_18141);
nor U18882 (N_18882,N_18421,N_18465);
nor U18883 (N_18883,N_18270,N_18096);
nand U18884 (N_18884,N_18481,N_18058);
nand U18885 (N_18885,N_18345,N_18380);
nand U18886 (N_18886,N_18321,N_18267);
or U18887 (N_18887,N_18229,N_18486);
and U18888 (N_18888,N_18223,N_18024);
nand U18889 (N_18889,N_18000,N_18411);
or U18890 (N_18890,N_18363,N_18219);
and U18891 (N_18891,N_18230,N_18116);
xor U18892 (N_18892,N_18157,N_18257);
and U18893 (N_18893,N_18003,N_18442);
nor U18894 (N_18894,N_18218,N_18074);
nor U18895 (N_18895,N_18124,N_18351);
nand U18896 (N_18896,N_18463,N_18118);
nand U18897 (N_18897,N_18192,N_18295);
nand U18898 (N_18898,N_18339,N_18022);
and U18899 (N_18899,N_18438,N_18488);
nor U18900 (N_18900,N_18211,N_18139);
or U18901 (N_18901,N_18171,N_18497);
xnor U18902 (N_18902,N_18403,N_18341);
and U18903 (N_18903,N_18033,N_18336);
and U18904 (N_18904,N_18389,N_18499);
xnor U18905 (N_18905,N_18245,N_18281);
nor U18906 (N_18906,N_18087,N_18043);
nor U18907 (N_18907,N_18021,N_18272);
nand U18908 (N_18908,N_18416,N_18021);
and U18909 (N_18909,N_18259,N_18263);
nor U18910 (N_18910,N_18217,N_18219);
or U18911 (N_18911,N_18010,N_18327);
nand U18912 (N_18912,N_18245,N_18482);
nand U18913 (N_18913,N_18432,N_18391);
and U18914 (N_18914,N_18291,N_18087);
nor U18915 (N_18915,N_18296,N_18411);
xnor U18916 (N_18916,N_18117,N_18055);
xnor U18917 (N_18917,N_18299,N_18477);
or U18918 (N_18918,N_18217,N_18084);
and U18919 (N_18919,N_18171,N_18140);
nand U18920 (N_18920,N_18148,N_18035);
or U18921 (N_18921,N_18148,N_18431);
or U18922 (N_18922,N_18351,N_18003);
nor U18923 (N_18923,N_18289,N_18208);
xnor U18924 (N_18924,N_18037,N_18111);
or U18925 (N_18925,N_18097,N_18387);
and U18926 (N_18926,N_18045,N_18417);
or U18927 (N_18927,N_18027,N_18151);
nor U18928 (N_18928,N_18343,N_18440);
and U18929 (N_18929,N_18161,N_18378);
xor U18930 (N_18930,N_18291,N_18022);
or U18931 (N_18931,N_18126,N_18490);
or U18932 (N_18932,N_18328,N_18071);
nand U18933 (N_18933,N_18028,N_18161);
nand U18934 (N_18934,N_18260,N_18469);
and U18935 (N_18935,N_18300,N_18437);
and U18936 (N_18936,N_18171,N_18094);
nand U18937 (N_18937,N_18321,N_18440);
xnor U18938 (N_18938,N_18411,N_18015);
and U18939 (N_18939,N_18090,N_18362);
or U18940 (N_18940,N_18132,N_18227);
nor U18941 (N_18941,N_18245,N_18293);
or U18942 (N_18942,N_18416,N_18275);
nor U18943 (N_18943,N_18085,N_18485);
nor U18944 (N_18944,N_18331,N_18174);
xor U18945 (N_18945,N_18194,N_18053);
or U18946 (N_18946,N_18157,N_18250);
or U18947 (N_18947,N_18003,N_18303);
or U18948 (N_18948,N_18497,N_18453);
xor U18949 (N_18949,N_18368,N_18269);
nand U18950 (N_18950,N_18381,N_18200);
nand U18951 (N_18951,N_18007,N_18187);
nand U18952 (N_18952,N_18436,N_18349);
nand U18953 (N_18953,N_18334,N_18385);
xnor U18954 (N_18954,N_18472,N_18307);
and U18955 (N_18955,N_18069,N_18171);
xnor U18956 (N_18956,N_18074,N_18016);
or U18957 (N_18957,N_18109,N_18211);
or U18958 (N_18958,N_18020,N_18080);
and U18959 (N_18959,N_18293,N_18069);
or U18960 (N_18960,N_18284,N_18132);
or U18961 (N_18961,N_18495,N_18378);
nand U18962 (N_18962,N_18091,N_18147);
or U18963 (N_18963,N_18286,N_18202);
nor U18964 (N_18964,N_18214,N_18091);
nand U18965 (N_18965,N_18180,N_18340);
xnor U18966 (N_18966,N_18298,N_18264);
and U18967 (N_18967,N_18460,N_18406);
and U18968 (N_18968,N_18059,N_18264);
and U18969 (N_18969,N_18001,N_18415);
xor U18970 (N_18970,N_18244,N_18461);
nor U18971 (N_18971,N_18028,N_18259);
xor U18972 (N_18972,N_18087,N_18387);
or U18973 (N_18973,N_18313,N_18328);
and U18974 (N_18974,N_18481,N_18013);
nor U18975 (N_18975,N_18111,N_18181);
nor U18976 (N_18976,N_18089,N_18393);
and U18977 (N_18977,N_18045,N_18312);
nor U18978 (N_18978,N_18115,N_18199);
and U18979 (N_18979,N_18333,N_18456);
xor U18980 (N_18980,N_18150,N_18073);
and U18981 (N_18981,N_18180,N_18200);
nor U18982 (N_18982,N_18144,N_18238);
nand U18983 (N_18983,N_18234,N_18424);
nand U18984 (N_18984,N_18140,N_18021);
nor U18985 (N_18985,N_18271,N_18009);
or U18986 (N_18986,N_18162,N_18428);
nand U18987 (N_18987,N_18392,N_18133);
nor U18988 (N_18988,N_18402,N_18219);
or U18989 (N_18989,N_18483,N_18162);
and U18990 (N_18990,N_18292,N_18453);
and U18991 (N_18991,N_18382,N_18468);
or U18992 (N_18992,N_18275,N_18250);
and U18993 (N_18993,N_18061,N_18325);
and U18994 (N_18994,N_18233,N_18272);
nor U18995 (N_18995,N_18050,N_18211);
xnor U18996 (N_18996,N_18399,N_18390);
nor U18997 (N_18997,N_18200,N_18453);
xor U18998 (N_18998,N_18190,N_18099);
or U18999 (N_18999,N_18047,N_18284);
or U19000 (N_19000,N_18565,N_18774);
nand U19001 (N_19001,N_18708,N_18698);
nor U19002 (N_19002,N_18938,N_18559);
and U19003 (N_19003,N_18600,N_18736);
and U19004 (N_19004,N_18739,N_18597);
xor U19005 (N_19005,N_18725,N_18504);
nand U19006 (N_19006,N_18624,N_18956);
nand U19007 (N_19007,N_18680,N_18834);
or U19008 (N_19008,N_18779,N_18733);
and U19009 (N_19009,N_18825,N_18584);
nand U19010 (N_19010,N_18931,N_18943);
nand U19011 (N_19011,N_18686,N_18660);
nand U19012 (N_19012,N_18722,N_18959);
or U19013 (N_19013,N_18861,N_18901);
xnor U19014 (N_19014,N_18630,N_18681);
xor U19015 (N_19015,N_18862,N_18812);
or U19016 (N_19016,N_18976,N_18509);
nor U19017 (N_19017,N_18541,N_18591);
nor U19018 (N_19018,N_18513,N_18616);
and U19019 (N_19019,N_18868,N_18993);
or U19020 (N_19020,N_18973,N_18989);
xnor U19021 (N_19021,N_18794,N_18639);
nor U19022 (N_19022,N_18870,N_18661);
xor U19023 (N_19023,N_18685,N_18902);
nor U19024 (N_19024,N_18614,N_18878);
or U19025 (N_19025,N_18699,N_18998);
nor U19026 (N_19026,N_18879,N_18545);
nand U19027 (N_19027,N_18816,N_18835);
xnor U19028 (N_19028,N_18824,N_18622);
or U19029 (N_19029,N_18766,N_18845);
xnor U19030 (N_19030,N_18769,N_18970);
and U19031 (N_19031,N_18690,N_18795);
nor U19032 (N_19032,N_18646,N_18991);
nor U19033 (N_19033,N_18642,N_18873);
nand U19034 (N_19034,N_18728,N_18745);
xnor U19035 (N_19035,N_18720,N_18631);
and U19036 (N_19036,N_18582,N_18884);
and U19037 (N_19037,N_18760,N_18992);
nand U19038 (N_19038,N_18536,N_18838);
nand U19039 (N_19039,N_18633,N_18542);
or U19040 (N_19040,N_18714,N_18859);
nor U19041 (N_19041,N_18598,N_18529);
nor U19042 (N_19042,N_18549,N_18819);
nor U19043 (N_19043,N_18653,N_18744);
nor U19044 (N_19044,N_18514,N_18923);
nor U19045 (N_19045,N_18520,N_18789);
xor U19046 (N_19046,N_18511,N_18572);
or U19047 (N_19047,N_18710,N_18783);
nand U19048 (N_19048,N_18735,N_18594);
and U19049 (N_19049,N_18727,N_18562);
and U19050 (N_19050,N_18945,N_18953);
nor U19051 (N_19051,N_18926,N_18811);
nor U19052 (N_19052,N_18921,N_18900);
or U19053 (N_19053,N_18607,N_18571);
nor U19054 (N_19054,N_18941,N_18895);
or U19055 (N_19055,N_18979,N_18502);
and U19056 (N_19056,N_18846,N_18674);
and U19057 (N_19057,N_18601,N_18781);
and U19058 (N_19058,N_18826,N_18822);
nor U19059 (N_19059,N_18623,N_18737);
nand U19060 (N_19060,N_18919,N_18673);
nand U19061 (N_19061,N_18537,N_18620);
nand U19062 (N_19062,N_18758,N_18797);
and U19063 (N_19063,N_18823,N_18915);
and U19064 (N_19064,N_18543,N_18899);
and U19065 (N_19065,N_18944,N_18629);
or U19066 (N_19066,N_18531,N_18867);
nor U19067 (N_19067,N_18679,N_18750);
xnor U19068 (N_19068,N_18648,N_18837);
nor U19069 (N_19069,N_18687,N_18676);
or U19070 (N_19070,N_18765,N_18599);
and U19071 (N_19071,N_18881,N_18592);
nor U19072 (N_19072,N_18694,N_18732);
nand U19073 (N_19073,N_18688,N_18922);
nor U19074 (N_19074,N_18856,N_18668);
xor U19075 (N_19075,N_18869,N_18820);
nand U19076 (N_19076,N_18626,N_18930);
nor U19077 (N_19077,N_18999,N_18875);
nand U19078 (N_19078,N_18790,N_18920);
or U19079 (N_19079,N_18664,N_18530);
xor U19080 (N_19080,N_18854,N_18711);
nand U19081 (N_19081,N_18963,N_18683);
and U19082 (N_19082,N_18833,N_18928);
and U19083 (N_19083,N_18893,N_18780);
nor U19084 (N_19084,N_18666,N_18756);
nor U19085 (N_19085,N_18505,N_18877);
xor U19086 (N_19086,N_18715,N_18508);
nor U19087 (N_19087,N_18843,N_18525);
nor U19088 (N_19088,N_18964,N_18975);
nor U19089 (N_19089,N_18995,N_18815);
or U19090 (N_19090,N_18813,N_18649);
nor U19091 (N_19091,N_18883,N_18782);
or U19092 (N_19092,N_18585,N_18654);
or U19093 (N_19093,N_18526,N_18994);
or U19094 (N_19094,N_18593,N_18717);
and U19095 (N_19095,N_18675,N_18768);
and U19096 (N_19096,N_18942,N_18982);
and U19097 (N_19097,N_18665,N_18621);
nor U19098 (N_19098,N_18932,N_18645);
xor U19099 (N_19099,N_18880,N_18772);
nand U19100 (N_19100,N_18552,N_18821);
xnor U19101 (N_19101,N_18535,N_18644);
nand U19102 (N_19102,N_18850,N_18532);
nor U19103 (N_19103,N_18831,N_18807);
nand U19104 (N_19104,N_18934,N_18734);
and U19105 (N_19105,N_18810,N_18596);
xnor U19106 (N_19106,N_18703,N_18684);
or U19107 (N_19107,N_18561,N_18628);
xnor U19108 (N_19108,N_18830,N_18551);
nand U19109 (N_19109,N_18839,N_18857);
and U19110 (N_19110,N_18985,N_18707);
and U19111 (N_19111,N_18962,N_18609);
nor U19112 (N_19112,N_18652,N_18618);
nor U19113 (N_19113,N_18983,N_18738);
nor U19114 (N_19114,N_18635,N_18967);
nor U19115 (N_19115,N_18527,N_18517);
xor U19116 (N_19116,N_18605,N_18540);
or U19117 (N_19117,N_18558,N_18887);
and U19118 (N_19118,N_18557,N_18897);
xnor U19119 (N_19119,N_18602,N_18863);
nand U19120 (N_19120,N_18556,N_18796);
or U19121 (N_19121,N_18905,N_18791);
and U19122 (N_19122,N_18961,N_18625);
and U19123 (N_19123,N_18809,N_18589);
xor U19124 (N_19124,N_18718,N_18578);
nand U19125 (N_19125,N_18904,N_18776);
nand U19126 (N_19126,N_18808,N_18671);
and U19127 (N_19127,N_18990,N_18672);
nor U19128 (N_19128,N_18757,N_18615);
nor U19129 (N_19129,N_18632,N_18740);
and U19130 (N_19130,N_18896,N_18603);
and U19131 (N_19131,N_18641,N_18951);
nand U19132 (N_19132,N_18909,N_18709);
and U19133 (N_19133,N_18748,N_18519);
and U19134 (N_19134,N_18954,N_18804);
and U19135 (N_19135,N_18871,N_18606);
or U19136 (N_19136,N_18534,N_18829);
and U19137 (N_19137,N_18784,N_18640);
or U19138 (N_19138,N_18972,N_18658);
xor U19139 (N_19139,N_18764,N_18981);
or U19140 (N_19140,N_18693,N_18637);
nand U19141 (N_19141,N_18864,N_18729);
nand U19142 (N_19142,N_18917,N_18827);
xor U19143 (N_19143,N_18980,N_18918);
nor U19144 (N_19144,N_18876,N_18761);
nand U19145 (N_19145,N_18691,N_18955);
nand U19146 (N_19146,N_18818,N_18988);
and U19147 (N_19147,N_18762,N_18885);
xor U19148 (N_19148,N_18908,N_18701);
xor U19149 (N_19149,N_18848,N_18528);
nand U19150 (N_19150,N_18771,N_18828);
nor U19151 (N_19151,N_18841,N_18907);
or U19152 (N_19152,N_18716,N_18849);
nand U19153 (N_19153,N_18759,N_18803);
or U19154 (N_19154,N_18925,N_18872);
xor U19155 (N_19155,N_18777,N_18906);
nand U19156 (N_19156,N_18501,N_18832);
or U19157 (N_19157,N_18563,N_18523);
or U19158 (N_19158,N_18507,N_18538);
or U19159 (N_19159,N_18987,N_18946);
xor U19160 (N_19160,N_18533,N_18705);
or U19161 (N_19161,N_18984,N_18889);
nand U19162 (N_19162,N_18965,N_18700);
or U19163 (N_19163,N_18969,N_18663);
xnor U19164 (N_19164,N_18677,N_18793);
or U19165 (N_19165,N_18997,N_18888);
nand U19166 (N_19166,N_18719,N_18912);
and U19167 (N_19167,N_18583,N_18546);
xnor U19168 (N_19168,N_18590,N_18595);
nor U19169 (N_19169,N_18555,N_18503);
nor U19170 (N_19170,N_18657,N_18911);
xor U19171 (N_19171,N_18860,N_18662);
or U19172 (N_19172,N_18891,N_18724);
or U19173 (N_19173,N_18682,N_18773);
and U19174 (N_19174,N_18580,N_18886);
nor U19175 (N_19175,N_18586,N_18712);
xor U19176 (N_19176,N_18512,N_18894);
nand U19177 (N_19177,N_18763,N_18619);
xnor U19178 (N_19178,N_18892,N_18650);
and U19179 (N_19179,N_18842,N_18550);
nand U19180 (N_19180,N_18933,N_18858);
and U19181 (N_19181,N_18806,N_18882);
and U19182 (N_19182,N_18966,N_18996);
nor U19183 (N_19183,N_18655,N_18567);
and U19184 (N_19184,N_18627,N_18643);
xnor U19185 (N_19185,N_18576,N_18890);
or U19186 (N_19186,N_18952,N_18566);
nor U19187 (N_19187,N_18554,N_18689);
nor U19188 (N_19188,N_18788,N_18678);
xor U19189 (N_19189,N_18852,N_18778);
and U19190 (N_19190,N_18634,N_18579);
or U19191 (N_19191,N_18787,N_18581);
and U19192 (N_19192,N_18948,N_18723);
or U19193 (N_19193,N_18617,N_18741);
or U19194 (N_19194,N_18770,N_18924);
nand U19195 (N_19195,N_18721,N_18805);
nand U19196 (N_19196,N_18754,N_18939);
and U19197 (N_19197,N_18817,N_18749);
or U19198 (N_19198,N_18751,N_18574);
nand U19199 (N_19199,N_18874,N_18799);
nor U19200 (N_19200,N_18713,N_18516);
nand U19201 (N_19201,N_18974,N_18611);
and U19202 (N_19202,N_18950,N_18553);
nand U19203 (N_19203,N_18914,N_18604);
xnor U19204 (N_19204,N_18753,N_18743);
xor U19205 (N_19205,N_18569,N_18865);
xnor U19206 (N_19206,N_18986,N_18669);
and U19207 (N_19207,N_18610,N_18903);
nand U19208 (N_19208,N_18692,N_18667);
nor U19209 (N_19209,N_18706,N_18971);
and U19210 (N_19210,N_18500,N_18847);
nand U19211 (N_19211,N_18851,N_18522);
nor U19212 (N_19212,N_18855,N_18651);
nand U19213 (N_19213,N_18746,N_18656);
nand U19214 (N_19214,N_18747,N_18844);
xor U19215 (N_19215,N_18853,N_18978);
or U19216 (N_19216,N_18929,N_18947);
and U19217 (N_19217,N_18564,N_18957);
and U19218 (N_19218,N_18659,N_18587);
or U19219 (N_19219,N_18937,N_18785);
nand U19220 (N_19220,N_18521,N_18731);
nor U19221 (N_19221,N_18840,N_18767);
xor U19222 (N_19222,N_18968,N_18786);
and U19223 (N_19223,N_18612,N_18548);
and U19224 (N_19224,N_18742,N_18958);
xor U19225 (N_19225,N_18670,N_18575);
nand U19226 (N_19226,N_18518,N_18524);
nand U19227 (N_19227,N_18696,N_18801);
nor U19228 (N_19228,N_18730,N_18539);
nor U19229 (N_19229,N_18573,N_18936);
nor U19230 (N_19230,N_18506,N_18916);
xnor U19231 (N_19231,N_18608,N_18977);
xnor U19232 (N_19232,N_18697,N_18910);
nor U19233 (N_19233,N_18613,N_18836);
and U19234 (N_19234,N_18898,N_18752);
and U19235 (N_19235,N_18798,N_18726);
nand U19236 (N_19236,N_18510,N_18940);
nor U19237 (N_19237,N_18814,N_18802);
and U19238 (N_19238,N_18560,N_18927);
and U19239 (N_19239,N_18702,N_18935);
nand U19240 (N_19240,N_18588,N_18638);
xnor U19241 (N_19241,N_18960,N_18636);
or U19242 (N_19242,N_18647,N_18913);
nor U19243 (N_19243,N_18695,N_18866);
or U19244 (N_19244,N_18755,N_18949);
nor U19245 (N_19245,N_18704,N_18775);
nand U19246 (N_19246,N_18792,N_18570);
and U19247 (N_19247,N_18800,N_18544);
or U19248 (N_19248,N_18547,N_18577);
or U19249 (N_19249,N_18515,N_18568);
nor U19250 (N_19250,N_18668,N_18542);
xnor U19251 (N_19251,N_18968,N_18679);
xor U19252 (N_19252,N_18860,N_18921);
nor U19253 (N_19253,N_18785,N_18733);
or U19254 (N_19254,N_18990,N_18557);
xnor U19255 (N_19255,N_18856,N_18645);
nand U19256 (N_19256,N_18507,N_18522);
or U19257 (N_19257,N_18565,N_18842);
nand U19258 (N_19258,N_18683,N_18871);
or U19259 (N_19259,N_18883,N_18534);
and U19260 (N_19260,N_18967,N_18783);
nand U19261 (N_19261,N_18940,N_18614);
and U19262 (N_19262,N_18685,N_18819);
nand U19263 (N_19263,N_18500,N_18593);
nand U19264 (N_19264,N_18749,N_18577);
nor U19265 (N_19265,N_18860,N_18582);
or U19266 (N_19266,N_18980,N_18665);
and U19267 (N_19267,N_18838,N_18784);
nor U19268 (N_19268,N_18763,N_18583);
or U19269 (N_19269,N_18571,N_18633);
or U19270 (N_19270,N_18918,N_18640);
nor U19271 (N_19271,N_18921,N_18952);
nor U19272 (N_19272,N_18528,N_18936);
nor U19273 (N_19273,N_18906,N_18513);
nor U19274 (N_19274,N_18581,N_18504);
nand U19275 (N_19275,N_18817,N_18735);
or U19276 (N_19276,N_18636,N_18527);
xor U19277 (N_19277,N_18664,N_18705);
nor U19278 (N_19278,N_18553,N_18641);
and U19279 (N_19279,N_18734,N_18664);
xnor U19280 (N_19280,N_18833,N_18891);
and U19281 (N_19281,N_18941,N_18860);
nor U19282 (N_19282,N_18744,N_18725);
or U19283 (N_19283,N_18958,N_18929);
and U19284 (N_19284,N_18547,N_18626);
and U19285 (N_19285,N_18559,N_18770);
xnor U19286 (N_19286,N_18538,N_18782);
nand U19287 (N_19287,N_18511,N_18663);
nor U19288 (N_19288,N_18555,N_18523);
or U19289 (N_19289,N_18597,N_18621);
nand U19290 (N_19290,N_18526,N_18910);
xnor U19291 (N_19291,N_18770,N_18841);
or U19292 (N_19292,N_18664,N_18555);
xnor U19293 (N_19293,N_18515,N_18971);
xor U19294 (N_19294,N_18550,N_18739);
nor U19295 (N_19295,N_18618,N_18987);
xnor U19296 (N_19296,N_18856,N_18628);
nand U19297 (N_19297,N_18886,N_18743);
or U19298 (N_19298,N_18648,N_18950);
xnor U19299 (N_19299,N_18881,N_18751);
and U19300 (N_19300,N_18669,N_18958);
nor U19301 (N_19301,N_18910,N_18859);
and U19302 (N_19302,N_18624,N_18710);
and U19303 (N_19303,N_18818,N_18870);
nand U19304 (N_19304,N_18716,N_18870);
nor U19305 (N_19305,N_18506,N_18957);
or U19306 (N_19306,N_18531,N_18960);
and U19307 (N_19307,N_18993,N_18966);
nor U19308 (N_19308,N_18652,N_18641);
and U19309 (N_19309,N_18581,N_18697);
or U19310 (N_19310,N_18531,N_18737);
nor U19311 (N_19311,N_18641,N_18863);
nand U19312 (N_19312,N_18850,N_18577);
nor U19313 (N_19313,N_18806,N_18748);
or U19314 (N_19314,N_18593,N_18600);
xor U19315 (N_19315,N_18986,N_18740);
nor U19316 (N_19316,N_18912,N_18694);
nand U19317 (N_19317,N_18636,N_18830);
or U19318 (N_19318,N_18515,N_18744);
xor U19319 (N_19319,N_18863,N_18700);
nand U19320 (N_19320,N_18954,N_18960);
nand U19321 (N_19321,N_18852,N_18753);
or U19322 (N_19322,N_18687,N_18756);
xor U19323 (N_19323,N_18846,N_18964);
xnor U19324 (N_19324,N_18857,N_18567);
xnor U19325 (N_19325,N_18943,N_18890);
or U19326 (N_19326,N_18926,N_18776);
and U19327 (N_19327,N_18689,N_18938);
and U19328 (N_19328,N_18623,N_18790);
and U19329 (N_19329,N_18984,N_18854);
xor U19330 (N_19330,N_18852,N_18553);
xnor U19331 (N_19331,N_18544,N_18939);
nand U19332 (N_19332,N_18758,N_18894);
and U19333 (N_19333,N_18631,N_18670);
or U19334 (N_19334,N_18509,N_18943);
nand U19335 (N_19335,N_18724,N_18848);
nand U19336 (N_19336,N_18570,N_18627);
or U19337 (N_19337,N_18853,N_18933);
and U19338 (N_19338,N_18835,N_18736);
nor U19339 (N_19339,N_18505,N_18537);
or U19340 (N_19340,N_18522,N_18744);
nor U19341 (N_19341,N_18650,N_18724);
nand U19342 (N_19342,N_18735,N_18963);
nand U19343 (N_19343,N_18656,N_18573);
or U19344 (N_19344,N_18832,N_18954);
nand U19345 (N_19345,N_18969,N_18569);
nor U19346 (N_19346,N_18550,N_18639);
nor U19347 (N_19347,N_18896,N_18857);
xor U19348 (N_19348,N_18726,N_18615);
and U19349 (N_19349,N_18584,N_18984);
nor U19350 (N_19350,N_18965,N_18703);
and U19351 (N_19351,N_18998,N_18920);
or U19352 (N_19352,N_18820,N_18530);
xnor U19353 (N_19353,N_18561,N_18674);
and U19354 (N_19354,N_18874,N_18563);
xnor U19355 (N_19355,N_18705,N_18861);
nand U19356 (N_19356,N_18673,N_18694);
xnor U19357 (N_19357,N_18628,N_18877);
nand U19358 (N_19358,N_18867,N_18747);
nor U19359 (N_19359,N_18955,N_18914);
or U19360 (N_19360,N_18577,N_18663);
and U19361 (N_19361,N_18607,N_18744);
nand U19362 (N_19362,N_18837,N_18818);
nor U19363 (N_19363,N_18704,N_18972);
nand U19364 (N_19364,N_18902,N_18533);
xnor U19365 (N_19365,N_18621,N_18976);
nand U19366 (N_19366,N_18903,N_18731);
and U19367 (N_19367,N_18786,N_18823);
xor U19368 (N_19368,N_18551,N_18719);
xor U19369 (N_19369,N_18997,N_18932);
and U19370 (N_19370,N_18736,N_18561);
and U19371 (N_19371,N_18755,N_18584);
nand U19372 (N_19372,N_18525,N_18996);
nor U19373 (N_19373,N_18895,N_18882);
or U19374 (N_19374,N_18779,N_18833);
nand U19375 (N_19375,N_18719,N_18527);
and U19376 (N_19376,N_18959,N_18833);
or U19377 (N_19377,N_18846,N_18640);
xnor U19378 (N_19378,N_18665,N_18712);
and U19379 (N_19379,N_18634,N_18903);
nand U19380 (N_19380,N_18694,N_18804);
and U19381 (N_19381,N_18863,N_18570);
nor U19382 (N_19382,N_18730,N_18931);
nand U19383 (N_19383,N_18774,N_18986);
xnor U19384 (N_19384,N_18942,N_18869);
nor U19385 (N_19385,N_18733,N_18718);
or U19386 (N_19386,N_18839,N_18833);
xor U19387 (N_19387,N_18940,N_18739);
or U19388 (N_19388,N_18886,N_18844);
nor U19389 (N_19389,N_18687,N_18820);
and U19390 (N_19390,N_18542,N_18757);
and U19391 (N_19391,N_18568,N_18541);
xor U19392 (N_19392,N_18824,N_18682);
nor U19393 (N_19393,N_18518,N_18632);
and U19394 (N_19394,N_18621,N_18881);
nor U19395 (N_19395,N_18956,N_18608);
xor U19396 (N_19396,N_18938,N_18648);
xnor U19397 (N_19397,N_18546,N_18524);
xor U19398 (N_19398,N_18536,N_18933);
and U19399 (N_19399,N_18811,N_18777);
and U19400 (N_19400,N_18798,N_18780);
nor U19401 (N_19401,N_18933,N_18753);
nor U19402 (N_19402,N_18752,N_18915);
xnor U19403 (N_19403,N_18904,N_18745);
xor U19404 (N_19404,N_18970,N_18708);
and U19405 (N_19405,N_18897,N_18822);
nand U19406 (N_19406,N_18618,N_18710);
or U19407 (N_19407,N_18647,N_18674);
and U19408 (N_19408,N_18915,N_18670);
nor U19409 (N_19409,N_18534,N_18690);
and U19410 (N_19410,N_18593,N_18803);
and U19411 (N_19411,N_18727,N_18548);
or U19412 (N_19412,N_18571,N_18564);
or U19413 (N_19413,N_18652,N_18946);
or U19414 (N_19414,N_18567,N_18744);
or U19415 (N_19415,N_18940,N_18692);
nor U19416 (N_19416,N_18935,N_18556);
or U19417 (N_19417,N_18962,N_18554);
or U19418 (N_19418,N_18806,N_18618);
nand U19419 (N_19419,N_18768,N_18505);
or U19420 (N_19420,N_18779,N_18760);
and U19421 (N_19421,N_18816,N_18760);
nand U19422 (N_19422,N_18594,N_18909);
and U19423 (N_19423,N_18848,N_18529);
xor U19424 (N_19424,N_18745,N_18919);
xnor U19425 (N_19425,N_18793,N_18684);
xnor U19426 (N_19426,N_18548,N_18896);
or U19427 (N_19427,N_18947,N_18843);
xnor U19428 (N_19428,N_18944,N_18717);
and U19429 (N_19429,N_18815,N_18785);
xor U19430 (N_19430,N_18538,N_18959);
nor U19431 (N_19431,N_18986,N_18715);
and U19432 (N_19432,N_18654,N_18622);
xnor U19433 (N_19433,N_18967,N_18728);
nand U19434 (N_19434,N_18629,N_18662);
xor U19435 (N_19435,N_18877,N_18910);
nand U19436 (N_19436,N_18504,N_18823);
or U19437 (N_19437,N_18739,N_18990);
and U19438 (N_19438,N_18923,N_18592);
nand U19439 (N_19439,N_18785,N_18831);
and U19440 (N_19440,N_18775,N_18943);
or U19441 (N_19441,N_18599,N_18542);
xnor U19442 (N_19442,N_18785,N_18701);
nand U19443 (N_19443,N_18780,N_18932);
and U19444 (N_19444,N_18700,N_18592);
nand U19445 (N_19445,N_18828,N_18777);
xnor U19446 (N_19446,N_18922,N_18967);
xor U19447 (N_19447,N_18616,N_18659);
xnor U19448 (N_19448,N_18834,N_18771);
and U19449 (N_19449,N_18573,N_18626);
and U19450 (N_19450,N_18508,N_18966);
nor U19451 (N_19451,N_18663,N_18602);
or U19452 (N_19452,N_18966,N_18761);
xnor U19453 (N_19453,N_18562,N_18986);
and U19454 (N_19454,N_18921,N_18675);
nand U19455 (N_19455,N_18969,N_18575);
nand U19456 (N_19456,N_18612,N_18988);
or U19457 (N_19457,N_18698,N_18881);
nand U19458 (N_19458,N_18698,N_18778);
nor U19459 (N_19459,N_18520,N_18824);
xnor U19460 (N_19460,N_18783,N_18512);
or U19461 (N_19461,N_18871,N_18769);
nor U19462 (N_19462,N_18671,N_18773);
nor U19463 (N_19463,N_18795,N_18941);
xnor U19464 (N_19464,N_18602,N_18891);
or U19465 (N_19465,N_18944,N_18725);
and U19466 (N_19466,N_18671,N_18960);
and U19467 (N_19467,N_18804,N_18921);
nor U19468 (N_19468,N_18845,N_18877);
or U19469 (N_19469,N_18676,N_18832);
or U19470 (N_19470,N_18517,N_18741);
and U19471 (N_19471,N_18917,N_18543);
nand U19472 (N_19472,N_18775,N_18520);
or U19473 (N_19473,N_18590,N_18904);
xor U19474 (N_19474,N_18535,N_18663);
xor U19475 (N_19475,N_18840,N_18922);
and U19476 (N_19476,N_18555,N_18999);
nor U19477 (N_19477,N_18853,N_18656);
xnor U19478 (N_19478,N_18732,N_18621);
nor U19479 (N_19479,N_18646,N_18903);
or U19480 (N_19480,N_18513,N_18715);
or U19481 (N_19481,N_18849,N_18647);
nor U19482 (N_19482,N_18621,N_18527);
and U19483 (N_19483,N_18620,N_18749);
nor U19484 (N_19484,N_18854,N_18709);
nor U19485 (N_19485,N_18777,N_18504);
or U19486 (N_19486,N_18883,N_18913);
xor U19487 (N_19487,N_18668,N_18742);
xnor U19488 (N_19488,N_18875,N_18697);
or U19489 (N_19489,N_18747,N_18949);
and U19490 (N_19490,N_18548,N_18850);
nand U19491 (N_19491,N_18757,N_18930);
or U19492 (N_19492,N_18872,N_18701);
xnor U19493 (N_19493,N_18553,N_18978);
and U19494 (N_19494,N_18757,N_18648);
nor U19495 (N_19495,N_18908,N_18942);
nor U19496 (N_19496,N_18575,N_18660);
xor U19497 (N_19497,N_18975,N_18868);
nor U19498 (N_19498,N_18611,N_18631);
nand U19499 (N_19499,N_18940,N_18791);
or U19500 (N_19500,N_19102,N_19313);
and U19501 (N_19501,N_19376,N_19497);
or U19502 (N_19502,N_19067,N_19339);
nor U19503 (N_19503,N_19066,N_19487);
xor U19504 (N_19504,N_19476,N_19143);
xor U19505 (N_19505,N_19494,N_19443);
nor U19506 (N_19506,N_19464,N_19237);
xor U19507 (N_19507,N_19206,N_19417);
and U19508 (N_19508,N_19056,N_19113);
nand U19509 (N_19509,N_19086,N_19352);
nand U19510 (N_19510,N_19452,N_19117);
xnor U19511 (N_19511,N_19266,N_19481);
or U19512 (N_19512,N_19164,N_19049);
nor U19513 (N_19513,N_19478,N_19027);
or U19514 (N_19514,N_19420,N_19083);
nand U19515 (N_19515,N_19069,N_19387);
xor U19516 (N_19516,N_19071,N_19465);
and U19517 (N_19517,N_19236,N_19114);
and U19518 (N_19518,N_19227,N_19292);
and U19519 (N_19519,N_19344,N_19447);
and U19520 (N_19520,N_19010,N_19409);
xnor U19521 (N_19521,N_19419,N_19490);
nand U19522 (N_19522,N_19239,N_19274);
nand U19523 (N_19523,N_19097,N_19343);
nor U19524 (N_19524,N_19238,N_19278);
nor U19525 (N_19525,N_19231,N_19175);
and U19526 (N_19526,N_19248,N_19099);
or U19527 (N_19527,N_19299,N_19311);
or U19528 (N_19528,N_19110,N_19005);
or U19529 (N_19529,N_19435,N_19403);
or U19530 (N_19530,N_19170,N_19038);
nor U19531 (N_19531,N_19275,N_19264);
and U19532 (N_19532,N_19093,N_19061);
nand U19533 (N_19533,N_19151,N_19324);
xor U19534 (N_19534,N_19378,N_19199);
or U19535 (N_19535,N_19309,N_19335);
or U19536 (N_19536,N_19222,N_19136);
nor U19537 (N_19537,N_19156,N_19214);
or U19538 (N_19538,N_19054,N_19233);
nand U19539 (N_19539,N_19124,N_19258);
and U19540 (N_19540,N_19127,N_19342);
and U19541 (N_19541,N_19004,N_19101);
xor U19542 (N_19542,N_19259,N_19123);
and U19543 (N_19543,N_19215,N_19469);
or U19544 (N_19544,N_19091,N_19297);
and U19545 (N_19545,N_19483,N_19211);
and U19546 (N_19546,N_19012,N_19319);
nand U19547 (N_19547,N_19493,N_19455);
xor U19548 (N_19548,N_19131,N_19281);
and U19549 (N_19549,N_19208,N_19267);
nand U19550 (N_19550,N_19158,N_19461);
nor U19551 (N_19551,N_19090,N_19060);
and U19552 (N_19552,N_19265,N_19251);
or U19553 (N_19553,N_19043,N_19022);
nand U19554 (N_19554,N_19453,N_19449);
nand U19555 (N_19555,N_19047,N_19003);
nand U19556 (N_19556,N_19210,N_19159);
nand U19557 (N_19557,N_19169,N_19139);
or U19558 (N_19558,N_19482,N_19219);
nor U19559 (N_19559,N_19204,N_19141);
or U19560 (N_19560,N_19293,N_19374);
xnor U19561 (N_19561,N_19314,N_19044);
nand U19562 (N_19562,N_19031,N_19082);
xnor U19563 (N_19563,N_19250,N_19023);
xnor U19564 (N_19564,N_19485,N_19228);
or U19565 (N_19565,N_19371,N_19207);
nor U19566 (N_19566,N_19225,N_19213);
nand U19567 (N_19567,N_19496,N_19077);
xor U19568 (N_19568,N_19221,N_19499);
and U19569 (N_19569,N_19039,N_19389);
or U19570 (N_19570,N_19130,N_19401);
nand U19571 (N_19571,N_19104,N_19326);
xnor U19572 (N_19572,N_19379,N_19394);
or U19573 (N_19573,N_19224,N_19057);
xor U19574 (N_19574,N_19122,N_19115);
or U19575 (N_19575,N_19128,N_19477);
nand U19576 (N_19576,N_19323,N_19303);
or U19577 (N_19577,N_19253,N_19018);
nor U19578 (N_19578,N_19171,N_19080);
and U19579 (N_19579,N_19386,N_19075);
and U19580 (N_19580,N_19334,N_19355);
and U19581 (N_19581,N_19486,N_19137);
and U19582 (N_19582,N_19246,N_19406);
xnor U19583 (N_19583,N_19349,N_19340);
nor U19584 (N_19584,N_19329,N_19306);
or U19585 (N_19585,N_19016,N_19445);
nor U19586 (N_19586,N_19242,N_19256);
xor U19587 (N_19587,N_19384,N_19184);
xnor U19588 (N_19588,N_19190,N_19350);
nor U19589 (N_19589,N_19468,N_19098);
or U19590 (N_19590,N_19072,N_19226);
or U19591 (N_19591,N_19084,N_19149);
xnor U19592 (N_19592,N_19300,N_19397);
nor U19593 (N_19593,N_19120,N_19174);
nand U19594 (N_19594,N_19491,N_19173);
nand U19595 (N_19595,N_19034,N_19446);
or U19596 (N_19596,N_19422,N_19232);
or U19597 (N_19597,N_19390,N_19112);
nor U19598 (N_19598,N_19229,N_19235);
nor U19599 (N_19599,N_19172,N_19459);
or U19600 (N_19600,N_19456,N_19203);
nor U19601 (N_19601,N_19198,N_19263);
and U19602 (N_19602,N_19051,N_19310);
nand U19603 (N_19603,N_19341,N_19188);
xnor U19604 (N_19604,N_19357,N_19183);
nand U19605 (N_19605,N_19289,N_19367);
nand U19606 (N_19606,N_19138,N_19145);
or U19607 (N_19607,N_19092,N_19282);
or U19608 (N_19608,N_19404,N_19019);
nand U19609 (N_19609,N_19327,N_19121);
nor U19610 (N_19610,N_19048,N_19166);
nor U19611 (N_19611,N_19347,N_19398);
and U19612 (N_19612,N_19070,N_19234);
nand U19613 (N_19613,N_19358,N_19372);
or U19614 (N_19614,N_19073,N_19150);
nand U19615 (N_19615,N_19094,N_19261);
and U19616 (N_19616,N_19200,N_19157);
xor U19617 (N_19617,N_19142,N_19365);
and U19618 (N_19618,N_19416,N_19277);
nand U19619 (N_19619,N_19153,N_19103);
nor U19620 (N_19620,N_19035,N_19014);
and U19621 (N_19621,N_19193,N_19212);
nor U19622 (N_19622,N_19382,N_19205);
or U19623 (N_19623,N_19163,N_19432);
nand U19624 (N_19624,N_19360,N_19021);
nor U19625 (N_19625,N_19036,N_19336);
or U19626 (N_19626,N_19498,N_19223);
or U19627 (N_19627,N_19279,N_19108);
and U19628 (N_19628,N_19029,N_19195);
xor U19629 (N_19629,N_19146,N_19002);
or U19630 (N_19630,N_19162,N_19053);
nor U19631 (N_19631,N_19454,N_19176);
xnor U19632 (N_19632,N_19272,N_19241);
nor U19633 (N_19633,N_19167,N_19421);
and U19634 (N_19634,N_19105,N_19074);
nand U19635 (N_19635,N_19148,N_19413);
or U19636 (N_19636,N_19109,N_19252);
and U19637 (N_19637,N_19424,N_19429);
or U19638 (N_19638,N_19011,N_19026);
and U19639 (N_19639,N_19007,N_19305);
and U19640 (N_19640,N_19088,N_19437);
or U19641 (N_19641,N_19196,N_19436);
nor U19642 (N_19642,N_19479,N_19194);
and U19643 (N_19643,N_19373,N_19472);
and U19644 (N_19644,N_19442,N_19187);
nand U19645 (N_19645,N_19189,N_19107);
xor U19646 (N_19646,N_19366,N_19134);
nor U19647 (N_19647,N_19216,N_19154);
xor U19648 (N_19648,N_19271,N_19249);
xor U19649 (N_19649,N_19359,N_19316);
nor U19650 (N_19650,N_19030,N_19155);
xnor U19651 (N_19651,N_19434,N_19475);
xnor U19652 (N_19652,N_19257,N_19337);
or U19653 (N_19653,N_19045,N_19202);
and U19654 (N_19654,N_19474,N_19106);
or U19655 (N_19655,N_19433,N_19348);
xor U19656 (N_19656,N_19118,N_19050);
nor U19657 (N_19657,N_19059,N_19430);
or U19658 (N_19658,N_19458,N_19388);
xor U19659 (N_19659,N_19492,N_19407);
nand U19660 (N_19660,N_19414,N_19197);
or U19661 (N_19661,N_19370,N_19353);
nor U19662 (N_19662,N_19361,N_19042);
nand U19663 (N_19663,N_19381,N_19046);
nand U19664 (N_19664,N_19439,N_19063);
and U19665 (N_19665,N_19395,N_19220);
and U19666 (N_19666,N_19408,N_19135);
nand U19667 (N_19667,N_19426,N_19296);
nor U19668 (N_19668,N_19418,N_19160);
or U19669 (N_19669,N_19470,N_19133);
nor U19670 (N_19670,N_19402,N_19178);
nand U19671 (N_19671,N_19444,N_19037);
and U19672 (N_19672,N_19346,N_19144);
xnor U19673 (N_19673,N_19025,N_19116);
xnor U19674 (N_19674,N_19192,N_19280);
nand U19675 (N_19675,N_19308,N_19254);
nor U19676 (N_19676,N_19191,N_19412);
xnor U19677 (N_19677,N_19177,N_19325);
nor U19678 (N_19678,N_19377,N_19298);
nor U19679 (N_19679,N_19119,N_19284);
or U19680 (N_19680,N_19307,N_19368);
xor U19681 (N_19681,N_19286,N_19000);
nor U19682 (N_19682,N_19268,N_19065);
nand U19683 (N_19683,N_19338,N_19245);
and U19684 (N_19684,N_19399,N_19321);
xnor U19685 (N_19685,N_19008,N_19312);
xnor U19686 (N_19686,N_19383,N_19425);
nor U19687 (N_19687,N_19411,N_19017);
nor U19688 (N_19688,N_19428,N_19400);
nand U19689 (N_19689,N_19255,N_19218);
xor U19690 (N_19690,N_19240,N_19333);
xor U19691 (N_19691,N_19457,N_19095);
and U19692 (N_19692,N_19362,N_19262);
and U19693 (N_19693,N_19427,N_19363);
nor U19694 (N_19694,N_19460,N_19466);
or U19695 (N_19695,N_19096,N_19396);
nor U19696 (N_19696,N_19354,N_19078);
and U19697 (N_19697,N_19140,N_19315);
or U19698 (N_19698,N_19283,N_19009);
nand U19699 (N_19699,N_19186,N_19369);
xor U19700 (N_19700,N_19168,N_19209);
or U19701 (N_19701,N_19380,N_19364);
xor U19702 (N_19702,N_19161,N_19230);
or U19703 (N_19703,N_19330,N_19495);
nand U19704 (N_19704,N_19129,N_19013);
and U19705 (N_19705,N_19290,N_19285);
nand U19706 (N_19706,N_19015,N_19032);
and U19707 (N_19707,N_19273,N_19181);
and U19708 (N_19708,N_19385,N_19270);
nor U19709 (N_19709,N_19462,N_19322);
xor U19710 (N_19710,N_19081,N_19302);
and U19711 (N_19711,N_19185,N_19179);
xnor U19712 (N_19712,N_19448,N_19295);
nor U19713 (N_19713,N_19058,N_19331);
nor U19714 (N_19714,N_19431,N_19087);
nand U19715 (N_19715,N_19438,N_19041);
nand U19716 (N_19716,N_19304,N_19276);
or U19717 (N_19717,N_19345,N_19180);
xor U19718 (N_19718,N_19111,N_19076);
nand U19719 (N_19719,N_19320,N_19217);
xor U19720 (N_19720,N_19126,N_19484);
and U19721 (N_19721,N_19440,N_19028);
xnor U19722 (N_19722,N_19165,N_19288);
or U19723 (N_19723,N_19467,N_19125);
xor U19724 (N_19724,N_19488,N_19244);
xor U19725 (N_19725,N_19040,N_19147);
nand U19726 (N_19726,N_19375,N_19328);
nor U19727 (N_19727,N_19085,N_19356);
nor U19728 (N_19728,N_19318,N_19463);
or U19729 (N_19729,N_19415,N_19393);
nor U19730 (N_19730,N_19064,N_19489);
nor U19731 (N_19731,N_19201,N_19423);
and U19732 (N_19732,N_19052,N_19079);
nand U19733 (N_19733,N_19450,N_19068);
and U19734 (N_19734,N_19480,N_19024);
xor U19735 (N_19735,N_19089,N_19006);
and U19736 (N_19736,N_19152,N_19287);
and U19737 (N_19737,N_19182,N_19441);
nand U19738 (N_19738,N_19269,N_19291);
nor U19739 (N_19739,N_19243,N_19301);
nor U19740 (N_19740,N_19260,N_19332);
xor U19741 (N_19741,N_19294,N_19391);
or U19742 (N_19742,N_19055,N_19033);
nand U19743 (N_19743,N_19351,N_19100);
nor U19744 (N_19744,N_19001,N_19471);
and U19745 (N_19745,N_19317,N_19020);
nand U19746 (N_19746,N_19473,N_19247);
xnor U19747 (N_19747,N_19062,N_19405);
or U19748 (N_19748,N_19410,N_19132);
or U19749 (N_19749,N_19451,N_19392);
nand U19750 (N_19750,N_19424,N_19382);
or U19751 (N_19751,N_19260,N_19063);
or U19752 (N_19752,N_19445,N_19323);
nor U19753 (N_19753,N_19281,N_19376);
nand U19754 (N_19754,N_19384,N_19159);
nand U19755 (N_19755,N_19462,N_19182);
or U19756 (N_19756,N_19021,N_19328);
nand U19757 (N_19757,N_19170,N_19096);
nor U19758 (N_19758,N_19099,N_19019);
nor U19759 (N_19759,N_19106,N_19244);
nand U19760 (N_19760,N_19263,N_19201);
xnor U19761 (N_19761,N_19063,N_19116);
or U19762 (N_19762,N_19021,N_19370);
nand U19763 (N_19763,N_19200,N_19288);
or U19764 (N_19764,N_19166,N_19056);
nor U19765 (N_19765,N_19471,N_19099);
or U19766 (N_19766,N_19047,N_19444);
or U19767 (N_19767,N_19140,N_19452);
or U19768 (N_19768,N_19220,N_19055);
nor U19769 (N_19769,N_19277,N_19301);
xnor U19770 (N_19770,N_19093,N_19216);
nand U19771 (N_19771,N_19230,N_19150);
nand U19772 (N_19772,N_19264,N_19258);
or U19773 (N_19773,N_19352,N_19381);
xor U19774 (N_19774,N_19206,N_19109);
nand U19775 (N_19775,N_19311,N_19087);
xor U19776 (N_19776,N_19009,N_19250);
and U19777 (N_19777,N_19292,N_19044);
or U19778 (N_19778,N_19473,N_19390);
xor U19779 (N_19779,N_19415,N_19271);
or U19780 (N_19780,N_19235,N_19078);
and U19781 (N_19781,N_19471,N_19152);
nand U19782 (N_19782,N_19013,N_19115);
xor U19783 (N_19783,N_19409,N_19024);
or U19784 (N_19784,N_19274,N_19172);
and U19785 (N_19785,N_19348,N_19041);
nand U19786 (N_19786,N_19458,N_19143);
nor U19787 (N_19787,N_19057,N_19072);
and U19788 (N_19788,N_19336,N_19070);
nor U19789 (N_19789,N_19393,N_19094);
or U19790 (N_19790,N_19358,N_19207);
and U19791 (N_19791,N_19355,N_19001);
or U19792 (N_19792,N_19241,N_19259);
and U19793 (N_19793,N_19077,N_19278);
or U19794 (N_19794,N_19259,N_19314);
or U19795 (N_19795,N_19306,N_19256);
xor U19796 (N_19796,N_19319,N_19156);
and U19797 (N_19797,N_19467,N_19170);
or U19798 (N_19798,N_19335,N_19237);
xor U19799 (N_19799,N_19387,N_19359);
nor U19800 (N_19800,N_19459,N_19493);
or U19801 (N_19801,N_19297,N_19264);
xnor U19802 (N_19802,N_19080,N_19101);
xnor U19803 (N_19803,N_19000,N_19013);
nand U19804 (N_19804,N_19472,N_19103);
xor U19805 (N_19805,N_19421,N_19414);
nand U19806 (N_19806,N_19447,N_19126);
xnor U19807 (N_19807,N_19421,N_19102);
xor U19808 (N_19808,N_19418,N_19486);
nor U19809 (N_19809,N_19439,N_19387);
and U19810 (N_19810,N_19259,N_19297);
nand U19811 (N_19811,N_19179,N_19359);
xor U19812 (N_19812,N_19095,N_19081);
nand U19813 (N_19813,N_19186,N_19319);
nor U19814 (N_19814,N_19408,N_19160);
nor U19815 (N_19815,N_19467,N_19375);
nand U19816 (N_19816,N_19077,N_19258);
nand U19817 (N_19817,N_19019,N_19001);
xnor U19818 (N_19818,N_19239,N_19362);
nor U19819 (N_19819,N_19116,N_19361);
and U19820 (N_19820,N_19082,N_19401);
or U19821 (N_19821,N_19194,N_19070);
xnor U19822 (N_19822,N_19148,N_19459);
or U19823 (N_19823,N_19202,N_19119);
and U19824 (N_19824,N_19142,N_19178);
nor U19825 (N_19825,N_19162,N_19410);
or U19826 (N_19826,N_19068,N_19286);
nor U19827 (N_19827,N_19016,N_19440);
nand U19828 (N_19828,N_19217,N_19499);
nand U19829 (N_19829,N_19223,N_19490);
nor U19830 (N_19830,N_19301,N_19153);
and U19831 (N_19831,N_19399,N_19278);
nand U19832 (N_19832,N_19309,N_19150);
or U19833 (N_19833,N_19256,N_19444);
nand U19834 (N_19834,N_19000,N_19034);
nand U19835 (N_19835,N_19058,N_19173);
nor U19836 (N_19836,N_19182,N_19301);
xor U19837 (N_19837,N_19112,N_19097);
nor U19838 (N_19838,N_19177,N_19342);
or U19839 (N_19839,N_19245,N_19213);
xnor U19840 (N_19840,N_19030,N_19452);
xnor U19841 (N_19841,N_19377,N_19416);
xnor U19842 (N_19842,N_19483,N_19455);
or U19843 (N_19843,N_19102,N_19294);
xnor U19844 (N_19844,N_19421,N_19024);
and U19845 (N_19845,N_19429,N_19240);
xor U19846 (N_19846,N_19274,N_19247);
xor U19847 (N_19847,N_19455,N_19095);
and U19848 (N_19848,N_19006,N_19132);
or U19849 (N_19849,N_19483,N_19329);
and U19850 (N_19850,N_19001,N_19124);
nor U19851 (N_19851,N_19235,N_19093);
or U19852 (N_19852,N_19271,N_19050);
or U19853 (N_19853,N_19185,N_19093);
and U19854 (N_19854,N_19016,N_19323);
nor U19855 (N_19855,N_19063,N_19068);
xnor U19856 (N_19856,N_19339,N_19087);
xnor U19857 (N_19857,N_19035,N_19345);
nand U19858 (N_19858,N_19336,N_19286);
and U19859 (N_19859,N_19216,N_19230);
nor U19860 (N_19860,N_19237,N_19388);
nor U19861 (N_19861,N_19302,N_19036);
nor U19862 (N_19862,N_19416,N_19296);
nand U19863 (N_19863,N_19119,N_19240);
nor U19864 (N_19864,N_19171,N_19350);
xor U19865 (N_19865,N_19349,N_19219);
nor U19866 (N_19866,N_19122,N_19421);
nand U19867 (N_19867,N_19095,N_19250);
xnor U19868 (N_19868,N_19177,N_19210);
or U19869 (N_19869,N_19393,N_19202);
nand U19870 (N_19870,N_19278,N_19485);
xnor U19871 (N_19871,N_19170,N_19471);
and U19872 (N_19872,N_19162,N_19114);
or U19873 (N_19873,N_19463,N_19315);
nand U19874 (N_19874,N_19005,N_19497);
nand U19875 (N_19875,N_19013,N_19392);
nand U19876 (N_19876,N_19050,N_19426);
or U19877 (N_19877,N_19118,N_19235);
or U19878 (N_19878,N_19470,N_19093);
nor U19879 (N_19879,N_19344,N_19234);
xor U19880 (N_19880,N_19337,N_19186);
and U19881 (N_19881,N_19401,N_19017);
and U19882 (N_19882,N_19380,N_19461);
and U19883 (N_19883,N_19327,N_19449);
xnor U19884 (N_19884,N_19337,N_19476);
or U19885 (N_19885,N_19256,N_19054);
nor U19886 (N_19886,N_19193,N_19211);
nor U19887 (N_19887,N_19016,N_19267);
or U19888 (N_19888,N_19202,N_19080);
nand U19889 (N_19889,N_19393,N_19248);
and U19890 (N_19890,N_19219,N_19285);
nand U19891 (N_19891,N_19065,N_19258);
nand U19892 (N_19892,N_19340,N_19321);
nor U19893 (N_19893,N_19024,N_19045);
xor U19894 (N_19894,N_19231,N_19318);
nor U19895 (N_19895,N_19492,N_19325);
nor U19896 (N_19896,N_19475,N_19165);
or U19897 (N_19897,N_19361,N_19201);
xnor U19898 (N_19898,N_19133,N_19269);
or U19899 (N_19899,N_19403,N_19110);
or U19900 (N_19900,N_19184,N_19151);
or U19901 (N_19901,N_19062,N_19204);
xnor U19902 (N_19902,N_19438,N_19268);
nand U19903 (N_19903,N_19197,N_19313);
or U19904 (N_19904,N_19477,N_19070);
xnor U19905 (N_19905,N_19017,N_19157);
nand U19906 (N_19906,N_19159,N_19297);
nand U19907 (N_19907,N_19396,N_19389);
xnor U19908 (N_19908,N_19375,N_19061);
or U19909 (N_19909,N_19298,N_19482);
nor U19910 (N_19910,N_19005,N_19026);
or U19911 (N_19911,N_19274,N_19076);
or U19912 (N_19912,N_19313,N_19190);
or U19913 (N_19913,N_19022,N_19319);
xor U19914 (N_19914,N_19463,N_19017);
or U19915 (N_19915,N_19287,N_19125);
xnor U19916 (N_19916,N_19029,N_19449);
and U19917 (N_19917,N_19476,N_19435);
and U19918 (N_19918,N_19420,N_19344);
nor U19919 (N_19919,N_19216,N_19069);
and U19920 (N_19920,N_19067,N_19094);
nor U19921 (N_19921,N_19194,N_19131);
xnor U19922 (N_19922,N_19008,N_19426);
or U19923 (N_19923,N_19044,N_19392);
nand U19924 (N_19924,N_19066,N_19357);
or U19925 (N_19925,N_19142,N_19418);
and U19926 (N_19926,N_19287,N_19020);
and U19927 (N_19927,N_19365,N_19065);
nand U19928 (N_19928,N_19392,N_19468);
nor U19929 (N_19929,N_19236,N_19002);
and U19930 (N_19930,N_19488,N_19486);
nor U19931 (N_19931,N_19415,N_19237);
nor U19932 (N_19932,N_19007,N_19001);
or U19933 (N_19933,N_19265,N_19223);
and U19934 (N_19934,N_19300,N_19496);
or U19935 (N_19935,N_19343,N_19311);
or U19936 (N_19936,N_19195,N_19432);
nand U19937 (N_19937,N_19432,N_19312);
nand U19938 (N_19938,N_19398,N_19236);
xor U19939 (N_19939,N_19290,N_19122);
xor U19940 (N_19940,N_19302,N_19473);
nand U19941 (N_19941,N_19458,N_19329);
xor U19942 (N_19942,N_19047,N_19385);
xor U19943 (N_19943,N_19106,N_19232);
or U19944 (N_19944,N_19188,N_19241);
and U19945 (N_19945,N_19287,N_19432);
or U19946 (N_19946,N_19184,N_19227);
or U19947 (N_19947,N_19326,N_19282);
and U19948 (N_19948,N_19098,N_19137);
and U19949 (N_19949,N_19473,N_19236);
nand U19950 (N_19950,N_19043,N_19149);
and U19951 (N_19951,N_19210,N_19185);
nand U19952 (N_19952,N_19468,N_19211);
or U19953 (N_19953,N_19040,N_19003);
nor U19954 (N_19954,N_19367,N_19183);
and U19955 (N_19955,N_19392,N_19374);
nor U19956 (N_19956,N_19230,N_19157);
xor U19957 (N_19957,N_19045,N_19174);
nor U19958 (N_19958,N_19216,N_19275);
and U19959 (N_19959,N_19441,N_19112);
nand U19960 (N_19960,N_19220,N_19481);
and U19961 (N_19961,N_19029,N_19111);
xor U19962 (N_19962,N_19126,N_19348);
or U19963 (N_19963,N_19038,N_19217);
xor U19964 (N_19964,N_19149,N_19346);
nand U19965 (N_19965,N_19352,N_19361);
xor U19966 (N_19966,N_19199,N_19385);
and U19967 (N_19967,N_19079,N_19319);
xor U19968 (N_19968,N_19459,N_19102);
xor U19969 (N_19969,N_19335,N_19450);
nor U19970 (N_19970,N_19014,N_19419);
and U19971 (N_19971,N_19046,N_19195);
and U19972 (N_19972,N_19130,N_19199);
or U19973 (N_19973,N_19140,N_19251);
or U19974 (N_19974,N_19101,N_19354);
xor U19975 (N_19975,N_19064,N_19160);
nor U19976 (N_19976,N_19358,N_19201);
or U19977 (N_19977,N_19109,N_19138);
nor U19978 (N_19978,N_19216,N_19352);
xor U19979 (N_19979,N_19224,N_19431);
and U19980 (N_19980,N_19199,N_19472);
nor U19981 (N_19981,N_19235,N_19346);
and U19982 (N_19982,N_19366,N_19275);
xor U19983 (N_19983,N_19190,N_19244);
or U19984 (N_19984,N_19318,N_19336);
nand U19985 (N_19985,N_19303,N_19074);
or U19986 (N_19986,N_19022,N_19377);
and U19987 (N_19987,N_19412,N_19005);
and U19988 (N_19988,N_19254,N_19030);
or U19989 (N_19989,N_19455,N_19363);
and U19990 (N_19990,N_19340,N_19024);
or U19991 (N_19991,N_19053,N_19026);
and U19992 (N_19992,N_19002,N_19497);
or U19993 (N_19993,N_19028,N_19442);
nand U19994 (N_19994,N_19039,N_19084);
or U19995 (N_19995,N_19167,N_19090);
nand U19996 (N_19996,N_19354,N_19362);
nand U19997 (N_19997,N_19051,N_19203);
or U19998 (N_19998,N_19138,N_19424);
or U19999 (N_19999,N_19196,N_19447);
or UO_0 (O_0,N_19500,N_19992);
nor UO_1 (O_1,N_19727,N_19893);
or UO_2 (O_2,N_19879,N_19999);
nand UO_3 (O_3,N_19663,N_19506);
nor UO_4 (O_4,N_19628,N_19864);
and UO_5 (O_5,N_19741,N_19674);
nand UO_6 (O_6,N_19671,N_19836);
and UO_7 (O_7,N_19722,N_19941);
nand UO_8 (O_8,N_19818,N_19988);
xor UO_9 (O_9,N_19853,N_19954);
nor UO_10 (O_10,N_19655,N_19750);
and UO_11 (O_11,N_19822,N_19636);
or UO_12 (O_12,N_19967,N_19933);
or UO_13 (O_13,N_19591,N_19813);
xor UO_14 (O_14,N_19584,N_19731);
nor UO_15 (O_15,N_19590,N_19672);
and UO_16 (O_16,N_19502,N_19667);
xor UO_17 (O_17,N_19985,N_19969);
and UO_18 (O_18,N_19754,N_19517);
nand UO_19 (O_19,N_19695,N_19610);
or UO_20 (O_20,N_19598,N_19603);
xnor UO_21 (O_21,N_19611,N_19530);
xor UO_22 (O_22,N_19850,N_19563);
nand UO_23 (O_23,N_19989,N_19842);
or UO_24 (O_24,N_19849,N_19622);
and UO_25 (O_25,N_19793,N_19659);
nor UO_26 (O_26,N_19957,N_19561);
nor UO_27 (O_27,N_19649,N_19846);
or UO_28 (O_28,N_19608,N_19788);
nor UO_29 (O_29,N_19553,N_19617);
nor UO_30 (O_30,N_19535,N_19587);
or UO_31 (O_31,N_19520,N_19632);
xor UO_32 (O_32,N_19812,N_19810);
or UO_33 (O_33,N_19872,N_19523);
nand UO_34 (O_34,N_19567,N_19800);
nand UO_35 (O_35,N_19748,N_19665);
and UO_36 (O_36,N_19658,N_19994);
nor UO_37 (O_37,N_19844,N_19537);
nand UO_38 (O_38,N_19582,N_19915);
or UO_39 (O_39,N_19943,N_19743);
nand UO_40 (O_40,N_19705,N_19538);
nor UO_41 (O_41,N_19634,N_19828);
and UO_42 (O_42,N_19605,N_19935);
and UO_43 (O_43,N_19918,N_19669);
nand UO_44 (O_44,N_19895,N_19834);
xnor UO_45 (O_45,N_19703,N_19757);
or UO_46 (O_46,N_19824,N_19951);
and UO_47 (O_47,N_19599,N_19675);
nand UO_48 (O_48,N_19522,N_19960);
or UO_49 (O_49,N_19620,N_19513);
and UO_50 (O_50,N_19845,N_19977);
or UO_51 (O_51,N_19693,N_19886);
nand UO_52 (O_52,N_19556,N_19959);
nor UO_53 (O_53,N_19607,N_19682);
nor UO_54 (O_54,N_19714,N_19884);
and UO_55 (O_55,N_19863,N_19949);
and UO_56 (O_56,N_19709,N_19580);
nand UO_57 (O_57,N_19568,N_19692);
and UO_58 (O_58,N_19830,N_19630);
or UO_59 (O_59,N_19880,N_19588);
nand UO_60 (O_60,N_19546,N_19737);
or UO_61 (O_61,N_19916,N_19572);
or UO_62 (O_62,N_19971,N_19753);
xor UO_63 (O_63,N_19772,N_19797);
or UO_64 (O_64,N_19527,N_19545);
or UO_65 (O_65,N_19579,N_19765);
or UO_66 (O_66,N_19679,N_19504);
nor UO_67 (O_67,N_19621,N_19725);
nor UO_68 (O_68,N_19681,N_19982);
and UO_69 (O_69,N_19816,N_19633);
nand UO_70 (O_70,N_19713,N_19647);
nor UO_71 (O_71,N_19564,N_19749);
xor UO_72 (O_72,N_19688,N_19648);
xor UO_73 (O_73,N_19791,N_19548);
or UO_74 (O_74,N_19926,N_19883);
nand UO_75 (O_75,N_19928,N_19939);
xor UO_76 (O_76,N_19711,N_19676);
nor UO_77 (O_77,N_19925,N_19904);
nand UO_78 (O_78,N_19593,N_19787);
or UO_79 (O_79,N_19790,N_19931);
nand UO_80 (O_80,N_19877,N_19920);
or UO_81 (O_81,N_19697,N_19825);
or UO_82 (O_82,N_19917,N_19644);
or UO_83 (O_83,N_19616,N_19874);
nor UO_84 (O_84,N_19574,N_19759);
xor UO_85 (O_85,N_19801,N_19963);
nor UO_86 (O_86,N_19910,N_19751);
and UO_87 (O_87,N_19706,N_19595);
nand UO_88 (O_88,N_19654,N_19514);
nor UO_89 (O_89,N_19639,N_19686);
or UO_90 (O_90,N_19726,N_19701);
xor UO_91 (O_91,N_19745,N_19638);
nand UO_92 (O_92,N_19898,N_19902);
nor UO_93 (O_93,N_19889,N_19764);
xnor UO_94 (O_94,N_19600,N_19577);
and UO_95 (O_95,N_19852,N_19859);
or UO_96 (O_96,N_19952,N_19687);
or UO_97 (O_97,N_19732,N_19948);
xnor UO_98 (O_98,N_19717,N_19507);
nand UO_99 (O_99,N_19871,N_19562);
or UO_100 (O_100,N_19673,N_19823);
and UO_101 (O_101,N_19905,N_19991);
or UO_102 (O_102,N_19606,N_19503);
or UO_103 (O_103,N_19569,N_19981);
nand UO_104 (O_104,N_19715,N_19998);
and UO_105 (O_105,N_19642,N_19766);
or UO_106 (O_106,N_19792,N_19592);
or UO_107 (O_107,N_19885,N_19856);
xor UO_108 (O_108,N_19913,N_19937);
nand UO_109 (O_109,N_19733,N_19704);
or UO_110 (O_110,N_19909,N_19651);
nor UO_111 (O_111,N_19511,N_19668);
and UO_112 (O_112,N_19785,N_19940);
xor UO_113 (O_113,N_19804,N_19558);
and UO_114 (O_114,N_19983,N_19597);
or UO_115 (O_115,N_19854,N_19515);
or UO_116 (O_116,N_19964,N_19526);
nor UO_117 (O_117,N_19547,N_19802);
nand UO_118 (O_118,N_19867,N_19696);
nor UO_119 (O_119,N_19542,N_19589);
xor UO_120 (O_120,N_19795,N_19510);
and UO_121 (O_121,N_19770,N_19829);
and UO_122 (O_122,N_19736,N_19640);
nor UO_123 (O_123,N_19549,N_19805);
nor UO_124 (O_124,N_19919,N_19936);
nand UO_125 (O_125,N_19891,N_19763);
nand UO_126 (O_126,N_19664,N_19873);
and UO_127 (O_127,N_19811,N_19708);
nand UO_128 (O_128,N_19557,N_19956);
xor UO_129 (O_129,N_19888,N_19831);
nand UO_130 (O_130,N_19942,N_19907);
nor UO_131 (O_131,N_19626,N_19923);
and UO_132 (O_132,N_19718,N_19614);
or UO_133 (O_133,N_19968,N_19570);
and UO_134 (O_134,N_19966,N_19972);
or UO_135 (O_135,N_19958,N_19758);
xor UO_136 (O_136,N_19820,N_19650);
nand UO_137 (O_137,N_19979,N_19914);
and UO_138 (O_138,N_19906,N_19911);
and UO_139 (O_139,N_19821,N_19560);
or UO_140 (O_140,N_19631,N_19550);
nor UO_141 (O_141,N_19762,N_19990);
nand UO_142 (O_142,N_19728,N_19827);
nor UO_143 (O_143,N_19833,N_19625);
or UO_144 (O_144,N_19996,N_19719);
or UO_145 (O_145,N_19987,N_19694);
nor UO_146 (O_146,N_19809,N_19735);
nand UO_147 (O_147,N_19720,N_19578);
and UO_148 (O_148,N_19865,N_19922);
and UO_149 (O_149,N_19629,N_19585);
nor UO_150 (O_150,N_19678,N_19738);
xor UO_151 (O_151,N_19938,N_19861);
and UO_152 (O_152,N_19835,N_19552);
nor UO_153 (O_153,N_19531,N_19803);
xor UO_154 (O_154,N_19615,N_19740);
xor UO_155 (O_155,N_19768,N_19601);
nand UO_156 (O_156,N_19868,N_19583);
nor UO_157 (O_157,N_19912,N_19734);
and UO_158 (O_158,N_19784,N_19635);
and UO_159 (O_159,N_19993,N_19858);
or UO_160 (O_160,N_19742,N_19571);
or UO_161 (O_161,N_19586,N_19783);
xnor UO_162 (O_162,N_19519,N_19539);
xnor UO_163 (O_163,N_19817,N_19932);
xor UO_164 (O_164,N_19995,N_19899);
nand UO_165 (O_165,N_19984,N_19525);
nor UO_166 (O_166,N_19613,N_19755);
xnor UO_167 (O_167,N_19536,N_19826);
nand UO_168 (O_168,N_19712,N_19739);
or UO_169 (O_169,N_19646,N_19662);
nor UO_170 (O_170,N_19953,N_19819);
nor UO_171 (O_171,N_19660,N_19851);
or UO_172 (O_172,N_19908,N_19661);
or UO_173 (O_173,N_19776,N_19573);
nand UO_174 (O_174,N_19534,N_19976);
and UO_175 (O_175,N_19707,N_19652);
xnor UO_176 (O_176,N_19690,N_19848);
or UO_177 (O_177,N_19778,N_19729);
nand UO_178 (O_178,N_19961,N_19575);
xnor UO_179 (O_179,N_19841,N_19934);
nor UO_180 (O_180,N_19855,N_19698);
xor UO_181 (O_181,N_19799,N_19689);
nor UO_182 (O_182,N_19806,N_19807);
and UO_183 (O_183,N_19878,N_19594);
nand UO_184 (O_184,N_19767,N_19945);
and UO_185 (O_185,N_19840,N_19724);
or UO_186 (O_186,N_19779,N_19847);
or UO_187 (O_187,N_19540,N_19860);
nand UO_188 (O_188,N_19666,N_19814);
nor UO_189 (O_189,N_19524,N_19516);
xor UO_190 (O_190,N_19716,N_19896);
xor UO_191 (O_191,N_19508,N_19839);
xnor UO_192 (O_192,N_19700,N_19653);
nand UO_193 (O_193,N_19950,N_19837);
or UO_194 (O_194,N_19897,N_19930);
xor UO_195 (O_195,N_19887,N_19890);
and UO_196 (O_196,N_19532,N_19533);
nand UO_197 (O_197,N_19843,N_19760);
nand UO_198 (O_198,N_19955,N_19946);
and UO_199 (O_199,N_19645,N_19794);
xnor UO_200 (O_200,N_19541,N_19773);
nand UO_201 (O_201,N_19882,N_19554);
or UO_202 (O_202,N_19744,N_19619);
or UO_203 (O_203,N_19774,N_19602);
or UO_204 (O_204,N_19747,N_19509);
xnor UO_205 (O_205,N_19986,N_19980);
nand UO_206 (O_206,N_19832,N_19680);
xnor UO_207 (O_207,N_19881,N_19677);
xnor UO_208 (O_208,N_19710,N_19746);
and UO_209 (O_209,N_19944,N_19657);
and UO_210 (O_210,N_19781,N_19780);
or UO_211 (O_211,N_19974,N_19643);
and UO_212 (O_212,N_19894,N_19518);
nor UO_213 (O_213,N_19771,N_19581);
xnor UO_214 (O_214,N_19559,N_19875);
nor UO_215 (O_215,N_19900,N_19786);
and UO_216 (O_216,N_19612,N_19921);
nand UO_217 (O_217,N_19604,N_19808);
or UO_218 (O_218,N_19528,N_19866);
or UO_219 (O_219,N_19596,N_19975);
nor UO_220 (O_220,N_19551,N_19857);
and UO_221 (O_221,N_19566,N_19512);
nor UO_222 (O_222,N_19702,N_19685);
nand UO_223 (O_223,N_19501,N_19947);
nor UO_224 (O_224,N_19627,N_19761);
xnor UO_225 (O_225,N_19901,N_19965);
and UO_226 (O_226,N_19699,N_19838);
nor UO_227 (O_227,N_19623,N_19789);
and UO_228 (O_228,N_19618,N_19609);
xnor UO_229 (O_229,N_19555,N_19927);
nand UO_230 (O_230,N_19752,N_19769);
or UO_231 (O_231,N_19730,N_19815);
nand UO_232 (O_232,N_19798,N_19641);
or UO_233 (O_233,N_19544,N_19683);
nand UO_234 (O_234,N_19997,N_19862);
nand UO_235 (O_235,N_19576,N_19684);
xnor UO_236 (O_236,N_19929,N_19721);
nand UO_237 (O_237,N_19777,N_19691);
nor UO_238 (O_238,N_19892,N_19656);
nand UO_239 (O_239,N_19521,N_19637);
nand UO_240 (O_240,N_19870,N_19962);
or UO_241 (O_241,N_19624,N_19756);
xor UO_242 (O_242,N_19529,N_19796);
and UO_243 (O_243,N_19924,N_19775);
or UO_244 (O_244,N_19903,N_19505);
and UO_245 (O_245,N_19876,N_19670);
nand UO_246 (O_246,N_19973,N_19543);
and UO_247 (O_247,N_19565,N_19970);
nand UO_248 (O_248,N_19978,N_19782);
xnor UO_249 (O_249,N_19723,N_19869);
and UO_250 (O_250,N_19531,N_19630);
nor UO_251 (O_251,N_19919,N_19604);
nand UO_252 (O_252,N_19972,N_19750);
and UO_253 (O_253,N_19966,N_19634);
nor UO_254 (O_254,N_19599,N_19752);
and UO_255 (O_255,N_19505,N_19948);
or UO_256 (O_256,N_19974,N_19501);
xnor UO_257 (O_257,N_19932,N_19777);
or UO_258 (O_258,N_19645,N_19733);
xor UO_259 (O_259,N_19627,N_19619);
xnor UO_260 (O_260,N_19807,N_19540);
xor UO_261 (O_261,N_19587,N_19895);
or UO_262 (O_262,N_19862,N_19881);
or UO_263 (O_263,N_19841,N_19892);
nand UO_264 (O_264,N_19747,N_19759);
nand UO_265 (O_265,N_19798,N_19909);
xor UO_266 (O_266,N_19810,N_19643);
xnor UO_267 (O_267,N_19697,N_19773);
nor UO_268 (O_268,N_19553,N_19704);
nor UO_269 (O_269,N_19711,N_19786);
or UO_270 (O_270,N_19782,N_19873);
or UO_271 (O_271,N_19756,N_19637);
xor UO_272 (O_272,N_19664,N_19785);
xor UO_273 (O_273,N_19653,N_19677);
xor UO_274 (O_274,N_19788,N_19651);
xor UO_275 (O_275,N_19882,N_19598);
xor UO_276 (O_276,N_19578,N_19957);
nand UO_277 (O_277,N_19663,N_19779);
or UO_278 (O_278,N_19551,N_19800);
or UO_279 (O_279,N_19895,N_19639);
or UO_280 (O_280,N_19608,N_19686);
and UO_281 (O_281,N_19730,N_19994);
and UO_282 (O_282,N_19978,N_19654);
and UO_283 (O_283,N_19525,N_19911);
or UO_284 (O_284,N_19792,N_19926);
nand UO_285 (O_285,N_19815,N_19977);
nand UO_286 (O_286,N_19595,N_19778);
nor UO_287 (O_287,N_19743,N_19578);
nand UO_288 (O_288,N_19921,N_19834);
nand UO_289 (O_289,N_19966,N_19834);
and UO_290 (O_290,N_19602,N_19556);
or UO_291 (O_291,N_19931,N_19736);
xor UO_292 (O_292,N_19842,N_19687);
or UO_293 (O_293,N_19582,N_19635);
or UO_294 (O_294,N_19645,N_19796);
or UO_295 (O_295,N_19960,N_19838);
xor UO_296 (O_296,N_19692,N_19638);
or UO_297 (O_297,N_19970,N_19837);
and UO_298 (O_298,N_19825,N_19646);
nand UO_299 (O_299,N_19936,N_19532);
and UO_300 (O_300,N_19978,N_19816);
or UO_301 (O_301,N_19776,N_19631);
nor UO_302 (O_302,N_19730,N_19887);
or UO_303 (O_303,N_19996,N_19698);
nand UO_304 (O_304,N_19715,N_19914);
nand UO_305 (O_305,N_19565,N_19676);
nor UO_306 (O_306,N_19765,N_19743);
xnor UO_307 (O_307,N_19770,N_19555);
nand UO_308 (O_308,N_19702,N_19757);
or UO_309 (O_309,N_19644,N_19568);
xnor UO_310 (O_310,N_19779,N_19920);
or UO_311 (O_311,N_19708,N_19971);
nor UO_312 (O_312,N_19669,N_19572);
nand UO_313 (O_313,N_19941,N_19669);
nand UO_314 (O_314,N_19976,N_19520);
or UO_315 (O_315,N_19917,N_19529);
and UO_316 (O_316,N_19556,N_19671);
and UO_317 (O_317,N_19940,N_19795);
and UO_318 (O_318,N_19503,N_19710);
or UO_319 (O_319,N_19940,N_19508);
nor UO_320 (O_320,N_19663,N_19835);
and UO_321 (O_321,N_19974,N_19745);
and UO_322 (O_322,N_19719,N_19889);
nand UO_323 (O_323,N_19684,N_19578);
nand UO_324 (O_324,N_19528,N_19826);
xnor UO_325 (O_325,N_19621,N_19988);
nor UO_326 (O_326,N_19846,N_19766);
and UO_327 (O_327,N_19821,N_19667);
or UO_328 (O_328,N_19664,N_19565);
nor UO_329 (O_329,N_19582,N_19748);
or UO_330 (O_330,N_19963,N_19717);
or UO_331 (O_331,N_19564,N_19704);
or UO_332 (O_332,N_19786,N_19954);
or UO_333 (O_333,N_19685,N_19737);
or UO_334 (O_334,N_19801,N_19735);
or UO_335 (O_335,N_19560,N_19696);
nor UO_336 (O_336,N_19993,N_19998);
xnor UO_337 (O_337,N_19853,N_19566);
or UO_338 (O_338,N_19758,N_19621);
and UO_339 (O_339,N_19649,N_19785);
xnor UO_340 (O_340,N_19991,N_19914);
xor UO_341 (O_341,N_19718,N_19588);
nand UO_342 (O_342,N_19952,N_19737);
and UO_343 (O_343,N_19873,N_19813);
xor UO_344 (O_344,N_19771,N_19704);
or UO_345 (O_345,N_19980,N_19696);
nand UO_346 (O_346,N_19911,N_19674);
xnor UO_347 (O_347,N_19525,N_19544);
xnor UO_348 (O_348,N_19991,N_19922);
and UO_349 (O_349,N_19858,N_19839);
nor UO_350 (O_350,N_19623,N_19959);
xor UO_351 (O_351,N_19847,N_19677);
or UO_352 (O_352,N_19725,N_19748);
xnor UO_353 (O_353,N_19850,N_19600);
nor UO_354 (O_354,N_19663,N_19675);
or UO_355 (O_355,N_19606,N_19824);
nor UO_356 (O_356,N_19803,N_19691);
and UO_357 (O_357,N_19804,N_19912);
nor UO_358 (O_358,N_19696,N_19858);
or UO_359 (O_359,N_19792,N_19560);
nand UO_360 (O_360,N_19939,N_19625);
nand UO_361 (O_361,N_19969,N_19885);
xor UO_362 (O_362,N_19564,N_19592);
nor UO_363 (O_363,N_19920,N_19952);
nor UO_364 (O_364,N_19519,N_19602);
nor UO_365 (O_365,N_19528,N_19988);
or UO_366 (O_366,N_19512,N_19730);
nor UO_367 (O_367,N_19842,N_19997);
xor UO_368 (O_368,N_19951,N_19777);
and UO_369 (O_369,N_19851,N_19532);
xnor UO_370 (O_370,N_19669,N_19979);
nor UO_371 (O_371,N_19938,N_19989);
nor UO_372 (O_372,N_19924,N_19887);
nand UO_373 (O_373,N_19747,N_19658);
and UO_374 (O_374,N_19923,N_19651);
nor UO_375 (O_375,N_19942,N_19912);
nor UO_376 (O_376,N_19917,N_19502);
nand UO_377 (O_377,N_19840,N_19623);
nor UO_378 (O_378,N_19946,N_19924);
xor UO_379 (O_379,N_19601,N_19980);
nor UO_380 (O_380,N_19905,N_19685);
nor UO_381 (O_381,N_19829,N_19606);
or UO_382 (O_382,N_19592,N_19638);
xor UO_383 (O_383,N_19925,N_19523);
xor UO_384 (O_384,N_19805,N_19524);
or UO_385 (O_385,N_19935,N_19914);
nor UO_386 (O_386,N_19581,N_19500);
xor UO_387 (O_387,N_19828,N_19632);
nand UO_388 (O_388,N_19501,N_19658);
and UO_389 (O_389,N_19620,N_19964);
and UO_390 (O_390,N_19812,N_19718);
xnor UO_391 (O_391,N_19657,N_19907);
nand UO_392 (O_392,N_19893,N_19673);
and UO_393 (O_393,N_19539,N_19977);
and UO_394 (O_394,N_19531,N_19629);
nor UO_395 (O_395,N_19959,N_19922);
or UO_396 (O_396,N_19923,N_19890);
and UO_397 (O_397,N_19641,N_19944);
xor UO_398 (O_398,N_19996,N_19526);
nand UO_399 (O_399,N_19971,N_19670);
nor UO_400 (O_400,N_19540,N_19552);
nand UO_401 (O_401,N_19688,N_19545);
nand UO_402 (O_402,N_19938,N_19707);
xor UO_403 (O_403,N_19934,N_19776);
and UO_404 (O_404,N_19832,N_19753);
or UO_405 (O_405,N_19949,N_19839);
nand UO_406 (O_406,N_19720,N_19830);
nor UO_407 (O_407,N_19940,N_19641);
and UO_408 (O_408,N_19795,N_19613);
and UO_409 (O_409,N_19799,N_19869);
nor UO_410 (O_410,N_19992,N_19538);
nand UO_411 (O_411,N_19959,N_19996);
xnor UO_412 (O_412,N_19907,N_19725);
nand UO_413 (O_413,N_19508,N_19825);
or UO_414 (O_414,N_19894,N_19674);
or UO_415 (O_415,N_19929,N_19842);
and UO_416 (O_416,N_19625,N_19984);
xor UO_417 (O_417,N_19705,N_19698);
and UO_418 (O_418,N_19539,N_19647);
xnor UO_419 (O_419,N_19549,N_19843);
nor UO_420 (O_420,N_19669,N_19883);
and UO_421 (O_421,N_19807,N_19662);
xnor UO_422 (O_422,N_19835,N_19572);
and UO_423 (O_423,N_19811,N_19572);
or UO_424 (O_424,N_19763,N_19595);
nor UO_425 (O_425,N_19982,N_19748);
and UO_426 (O_426,N_19805,N_19955);
nand UO_427 (O_427,N_19651,N_19775);
or UO_428 (O_428,N_19500,N_19961);
or UO_429 (O_429,N_19739,N_19513);
nor UO_430 (O_430,N_19937,N_19971);
nor UO_431 (O_431,N_19651,N_19697);
and UO_432 (O_432,N_19814,N_19859);
and UO_433 (O_433,N_19904,N_19513);
and UO_434 (O_434,N_19957,N_19832);
and UO_435 (O_435,N_19793,N_19562);
or UO_436 (O_436,N_19624,N_19574);
nand UO_437 (O_437,N_19970,N_19505);
xor UO_438 (O_438,N_19745,N_19806);
nand UO_439 (O_439,N_19526,N_19889);
nand UO_440 (O_440,N_19862,N_19630);
nand UO_441 (O_441,N_19880,N_19599);
nand UO_442 (O_442,N_19556,N_19929);
or UO_443 (O_443,N_19742,N_19995);
or UO_444 (O_444,N_19521,N_19638);
and UO_445 (O_445,N_19865,N_19589);
and UO_446 (O_446,N_19630,N_19941);
nand UO_447 (O_447,N_19774,N_19606);
and UO_448 (O_448,N_19895,N_19788);
nand UO_449 (O_449,N_19602,N_19881);
or UO_450 (O_450,N_19805,N_19511);
and UO_451 (O_451,N_19868,N_19551);
nor UO_452 (O_452,N_19707,N_19575);
nand UO_453 (O_453,N_19621,N_19812);
or UO_454 (O_454,N_19691,N_19570);
xnor UO_455 (O_455,N_19979,N_19755);
or UO_456 (O_456,N_19706,N_19936);
or UO_457 (O_457,N_19560,N_19919);
and UO_458 (O_458,N_19926,N_19823);
xor UO_459 (O_459,N_19791,N_19860);
nand UO_460 (O_460,N_19842,N_19933);
nor UO_461 (O_461,N_19812,N_19857);
nand UO_462 (O_462,N_19515,N_19882);
xnor UO_463 (O_463,N_19745,N_19534);
nand UO_464 (O_464,N_19784,N_19983);
nand UO_465 (O_465,N_19534,N_19623);
or UO_466 (O_466,N_19774,N_19949);
or UO_467 (O_467,N_19942,N_19783);
and UO_468 (O_468,N_19628,N_19915);
and UO_469 (O_469,N_19907,N_19787);
and UO_470 (O_470,N_19846,N_19519);
and UO_471 (O_471,N_19955,N_19697);
nand UO_472 (O_472,N_19508,N_19553);
nand UO_473 (O_473,N_19833,N_19927);
xnor UO_474 (O_474,N_19887,N_19665);
nand UO_475 (O_475,N_19708,N_19753);
nand UO_476 (O_476,N_19860,N_19613);
or UO_477 (O_477,N_19777,N_19975);
nor UO_478 (O_478,N_19882,N_19794);
and UO_479 (O_479,N_19816,N_19704);
and UO_480 (O_480,N_19556,N_19909);
nand UO_481 (O_481,N_19936,N_19898);
xnor UO_482 (O_482,N_19913,N_19810);
xnor UO_483 (O_483,N_19541,N_19655);
or UO_484 (O_484,N_19668,N_19586);
or UO_485 (O_485,N_19848,N_19803);
and UO_486 (O_486,N_19794,N_19900);
xnor UO_487 (O_487,N_19876,N_19901);
nand UO_488 (O_488,N_19843,N_19517);
or UO_489 (O_489,N_19613,N_19586);
xnor UO_490 (O_490,N_19684,N_19889);
nand UO_491 (O_491,N_19821,N_19752);
nor UO_492 (O_492,N_19621,N_19975);
and UO_493 (O_493,N_19670,N_19985);
xnor UO_494 (O_494,N_19588,N_19647);
xor UO_495 (O_495,N_19933,N_19556);
or UO_496 (O_496,N_19839,N_19578);
xnor UO_497 (O_497,N_19630,N_19519);
nand UO_498 (O_498,N_19922,N_19660);
nor UO_499 (O_499,N_19554,N_19976);
nand UO_500 (O_500,N_19855,N_19927);
or UO_501 (O_501,N_19880,N_19726);
and UO_502 (O_502,N_19729,N_19929);
and UO_503 (O_503,N_19969,N_19829);
nand UO_504 (O_504,N_19973,N_19787);
xnor UO_505 (O_505,N_19881,N_19924);
and UO_506 (O_506,N_19846,N_19889);
or UO_507 (O_507,N_19562,N_19929);
xnor UO_508 (O_508,N_19529,N_19513);
xor UO_509 (O_509,N_19500,N_19993);
xor UO_510 (O_510,N_19859,N_19886);
and UO_511 (O_511,N_19839,N_19699);
xnor UO_512 (O_512,N_19604,N_19661);
and UO_513 (O_513,N_19563,N_19503);
or UO_514 (O_514,N_19917,N_19711);
and UO_515 (O_515,N_19782,N_19720);
nor UO_516 (O_516,N_19570,N_19958);
nand UO_517 (O_517,N_19982,N_19990);
or UO_518 (O_518,N_19982,N_19635);
nand UO_519 (O_519,N_19724,N_19675);
or UO_520 (O_520,N_19733,N_19900);
or UO_521 (O_521,N_19782,N_19684);
xor UO_522 (O_522,N_19785,N_19551);
nand UO_523 (O_523,N_19691,N_19629);
nand UO_524 (O_524,N_19592,N_19922);
xnor UO_525 (O_525,N_19928,N_19650);
xor UO_526 (O_526,N_19922,N_19757);
xnor UO_527 (O_527,N_19593,N_19838);
xnor UO_528 (O_528,N_19819,N_19849);
nand UO_529 (O_529,N_19512,N_19969);
nand UO_530 (O_530,N_19825,N_19918);
or UO_531 (O_531,N_19929,N_19538);
xnor UO_532 (O_532,N_19553,N_19871);
xnor UO_533 (O_533,N_19799,N_19904);
nand UO_534 (O_534,N_19577,N_19812);
xnor UO_535 (O_535,N_19783,N_19718);
nand UO_536 (O_536,N_19936,N_19703);
xnor UO_537 (O_537,N_19962,N_19840);
nor UO_538 (O_538,N_19766,N_19954);
nor UO_539 (O_539,N_19736,N_19867);
or UO_540 (O_540,N_19752,N_19961);
nor UO_541 (O_541,N_19864,N_19730);
or UO_542 (O_542,N_19937,N_19845);
nand UO_543 (O_543,N_19544,N_19871);
nor UO_544 (O_544,N_19738,N_19757);
nand UO_545 (O_545,N_19669,N_19700);
and UO_546 (O_546,N_19723,N_19516);
nand UO_547 (O_547,N_19720,N_19729);
and UO_548 (O_548,N_19597,N_19646);
and UO_549 (O_549,N_19769,N_19511);
nor UO_550 (O_550,N_19979,N_19535);
and UO_551 (O_551,N_19694,N_19509);
nor UO_552 (O_552,N_19736,N_19757);
nand UO_553 (O_553,N_19895,N_19955);
nand UO_554 (O_554,N_19861,N_19834);
xor UO_555 (O_555,N_19652,N_19929);
nand UO_556 (O_556,N_19897,N_19799);
or UO_557 (O_557,N_19970,N_19766);
and UO_558 (O_558,N_19725,N_19913);
xnor UO_559 (O_559,N_19753,N_19720);
xnor UO_560 (O_560,N_19757,N_19508);
and UO_561 (O_561,N_19749,N_19554);
xor UO_562 (O_562,N_19630,N_19528);
nor UO_563 (O_563,N_19896,N_19935);
nand UO_564 (O_564,N_19801,N_19540);
nor UO_565 (O_565,N_19687,N_19771);
nor UO_566 (O_566,N_19583,N_19578);
nor UO_567 (O_567,N_19742,N_19578);
xnor UO_568 (O_568,N_19527,N_19570);
or UO_569 (O_569,N_19551,N_19699);
and UO_570 (O_570,N_19841,N_19927);
xor UO_571 (O_571,N_19856,N_19846);
xnor UO_572 (O_572,N_19503,N_19719);
nor UO_573 (O_573,N_19849,N_19890);
nor UO_574 (O_574,N_19715,N_19645);
and UO_575 (O_575,N_19808,N_19569);
nand UO_576 (O_576,N_19686,N_19860);
xor UO_577 (O_577,N_19621,N_19618);
nand UO_578 (O_578,N_19614,N_19503);
and UO_579 (O_579,N_19998,N_19975);
or UO_580 (O_580,N_19559,N_19949);
nand UO_581 (O_581,N_19845,N_19617);
xnor UO_582 (O_582,N_19548,N_19853);
xnor UO_583 (O_583,N_19960,N_19965);
xor UO_584 (O_584,N_19540,N_19526);
and UO_585 (O_585,N_19713,N_19792);
or UO_586 (O_586,N_19774,N_19997);
or UO_587 (O_587,N_19838,N_19519);
or UO_588 (O_588,N_19651,N_19882);
and UO_589 (O_589,N_19818,N_19596);
and UO_590 (O_590,N_19954,N_19563);
xnor UO_591 (O_591,N_19960,N_19579);
nor UO_592 (O_592,N_19859,N_19971);
or UO_593 (O_593,N_19542,N_19625);
nand UO_594 (O_594,N_19728,N_19908);
xnor UO_595 (O_595,N_19807,N_19960);
and UO_596 (O_596,N_19638,N_19667);
and UO_597 (O_597,N_19955,N_19833);
xor UO_598 (O_598,N_19651,N_19905);
xnor UO_599 (O_599,N_19752,N_19836);
or UO_600 (O_600,N_19698,N_19971);
nor UO_601 (O_601,N_19673,N_19879);
nor UO_602 (O_602,N_19801,N_19587);
and UO_603 (O_603,N_19537,N_19763);
or UO_604 (O_604,N_19567,N_19919);
and UO_605 (O_605,N_19915,N_19554);
xor UO_606 (O_606,N_19774,N_19814);
and UO_607 (O_607,N_19708,N_19524);
xnor UO_608 (O_608,N_19976,N_19667);
and UO_609 (O_609,N_19710,N_19580);
and UO_610 (O_610,N_19913,N_19551);
nor UO_611 (O_611,N_19946,N_19890);
nor UO_612 (O_612,N_19897,N_19510);
or UO_613 (O_613,N_19707,N_19796);
and UO_614 (O_614,N_19757,N_19714);
nor UO_615 (O_615,N_19546,N_19762);
nor UO_616 (O_616,N_19671,N_19772);
xor UO_617 (O_617,N_19840,N_19785);
xor UO_618 (O_618,N_19820,N_19770);
xor UO_619 (O_619,N_19526,N_19747);
and UO_620 (O_620,N_19822,N_19961);
nor UO_621 (O_621,N_19892,N_19964);
nor UO_622 (O_622,N_19529,N_19869);
and UO_623 (O_623,N_19857,N_19609);
nor UO_624 (O_624,N_19643,N_19612);
nor UO_625 (O_625,N_19554,N_19969);
nand UO_626 (O_626,N_19665,N_19597);
xor UO_627 (O_627,N_19750,N_19658);
and UO_628 (O_628,N_19661,N_19570);
xor UO_629 (O_629,N_19590,N_19765);
nor UO_630 (O_630,N_19728,N_19636);
or UO_631 (O_631,N_19587,N_19797);
xor UO_632 (O_632,N_19619,N_19663);
or UO_633 (O_633,N_19990,N_19712);
nand UO_634 (O_634,N_19962,N_19775);
xnor UO_635 (O_635,N_19660,N_19969);
nand UO_636 (O_636,N_19684,N_19605);
nor UO_637 (O_637,N_19845,N_19809);
and UO_638 (O_638,N_19546,N_19945);
nor UO_639 (O_639,N_19708,N_19618);
and UO_640 (O_640,N_19609,N_19830);
and UO_641 (O_641,N_19965,N_19534);
and UO_642 (O_642,N_19790,N_19784);
xor UO_643 (O_643,N_19923,N_19942);
or UO_644 (O_644,N_19547,N_19900);
nor UO_645 (O_645,N_19891,N_19621);
or UO_646 (O_646,N_19783,N_19757);
nor UO_647 (O_647,N_19799,N_19775);
nor UO_648 (O_648,N_19615,N_19929);
nor UO_649 (O_649,N_19858,N_19682);
xnor UO_650 (O_650,N_19979,N_19751);
and UO_651 (O_651,N_19949,N_19718);
and UO_652 (O_652,N_19772,N_19784);
and UO_653 (O_653,N_19933,N_19833);
nor UO_654 (O_654,N_19500,N_19879);
nor UO_655 (O_655,N_19687,N_19659);
nor UO_656 (O_656,N_19914,N_19821);
xor UO_657 (O_657,N_19707,N_19639);
and UO_658 (O_658,N_19957,N_19650);
or UO_659 (O_659,N_19722,N_19533);
and UO_660 (O_660,N_19591,N_19858);
or UO_661 (O_661,N_19629,N_19729);
xor UO_662 (O_662,N_19743,N_19701);
nand UO_663 (O_663,N_19962,N_19677);
xnor UO_664 (O_664,N_19548,N_19511);
or UO_665 (O_665,N_19559,N_19604);
and UO_666 (O_666,N_19730,N_19837);
and UO_667 (O_667,N_19865,N_19551);
nand UO_668 (O_668,N_19895,N_19581);
nand UO_669 (O_669,N_19551,N_19970);
or UO_670 (O_670,N_19940,N_19936);
nor UO_671 (O_671,N_19957,N_19515);
or UO_672 (O_672,N_19916,N_19659);
and UO_673 (O_673,N_19674,N_19927);
or UO_674 (O_674,N_19949,N_19824);
or UO_675 (O_675,N_19646,N_19977);
nor UO_676 (O_676,N_19569,N_19850);
nor UO_677 (O_677,N_19738,N_19798);
xor UO_678 (O_678,N_19592,N_19860);
and UO_679 (O_679,N_19705,N_19878);
xor UO_680 (O_680,N_19591,N_19889);
or UO_681 (O_681,N_19886,N_19651);
nor UO_682 (O_682,N_19969,N_19645);
nand UO_683 (O_683,N_19881,N_19841);
and UO_684 (O_684,N_19510,N_19599);
nand UO_685 (O_685,N_19867,N_19841);
or UO_686 (O_686,N_19776,N_19967);
nor UO_687 (O_687,N_19860,N_19772);
and UO_688 (O_688,N_19566,N_19664);
xnor UO_689 (O_689,N_19587,N_19844);
and UO_690 (O_690,N_19624,N_19536);
nand UO_691 (O_691,N_19587,N_19735);
nand UO_692 (O_692,N_19784,N_19639);
nor UO_693 (O_693,N_19685,N_19537);
and UO_694 (O_694,N_19640,N_19959);
nor UO_695 (O_695,N_19508,N_19501);
and UO_696 (O_696,N_19894,N_19617);
and UO_697 (O_697,N_19754,N_19919);
and UO_698 (O_698,N_19561,N_19780);
nor UO_699 (O_699,N_19900,N_19911);
xor UO_700 (O_700,N_19801,N_19740);
and UO_701 (O_701,N_19781,N_19606);
nor UO_702 (O_702,N_19884,N_19892);
and UO_703 (O_703,N_19932,N_19730);
or UO_704 (O_704,N_19504,N_19842);
or UO_705 (O_705,N_19791,N_19950);
nand UO_706 (O_706,N_19784,N_19591);
xnor UO_707 (O_707,N_19981,N_19661);
nor UO_708 (O_708,N_19983,N_19839);
nand UO_709 (O_709,N_19998,N_19844);
and UO_710 (O_710,N_19969,N_19614);
nor UO_711 (O_711,N_19536,N_19825);
xnor UO_712 (O_712,N_19648,N_19846);
nor UO_713 (O_713,N_19991,N_19973);
or UO_714 (O_714,N_19716,N_19614);
xor UO_715 (O_715,N_19659,N_19769);
nor UO_716 (O_716,N_19620,N_19908);
nor UO_717 (O_717,N_19865,N_19682);
and UO_718 (O_718,N_19534,N_19622);
nor UO_719 (O_719,N_19559,N_19959);
xnor UO_720 (O_720,N_19647,N_19560);
and UO_721 (O_721,N_19953,N_19587);
nor UO_722 (O_722,N_19855,N_19613);
xnor UO_723 (O_723,N_19542,N_19964);
nand UO_724 (O_724,N_19811,N_19587);
or UO_725 (O_725,N_19563,N_19615);
nand UO_726 (O_726,N_19922,N_19821);
xor UO_727 (O_727,N_19855,N_19710);
or UO_728 (O_728,N_19904,N_19658);
or UO_729 (O_729,N_19648,N_19727);
and UO_730 (O_730,N_19798,N_19850);
xor UO_731 (O_731,N_19901,N_19513);
or UO_732 (O_732,N_19570,N_19725);
and UO_733 (O_733,N_19627,N_19871);
nand UO_734 (O_734,N_19529,N_19948);
and UO_735 (O_735,N_19525,N_19784);
nand UO_736 (O_736,N_19840,N_19603);
and UO_737 (O_737,N_19620,N_19653);
nor UO_738 (O_738,N_19959,N_19572);
nand UO_739 (O_739,N_19627,N_19984);
or UO_740 (O_740,N_19664,N_19997);
and UO_741 (O_741,N_19752,N_19963);
and UO_742 (O_742,N_19893,N_19714);
xnor UO_743 (O_743,N_19752,N_19848);
and UO_744 (O_744,N_19585,N_19654);
nand UO_745 (O_745,N_19896,N_19519);
nand UO_746 (O_746,N_19672,N_19504);
or UO_747 (O_747,N_19808,N_19606);
nand UO_748 (O_748,N_19519,N_19545);
nor UO_749 (O_749,N_19637,N_19969);
or UO_750 (O_750,N_19984,N_19638);
or UO_751 (O_751,N_19678,N_19579);
or UO_752 (O_752,N_19781,N_19575);
nand UO_753 (O_753,N_19975,N_19568);
xor UO_754 (O_754,N_19674,N_19837);
or UO_755 (O_755,N_19714,N_19750);
nor UO_756 (O_756,N_19609,N_19919);
nand UO_757 (O_757,N_19785,N_19887);
or UO_758 (O_758,N_19729,N_19915);
nor UO_759 (O_759,N_19791,N_19744);
and UO_760 (O_760,N_19892,N_19790);
or UO_761 (O_761,N_19603,N_19639);
or UO_762 (O_762,N_19549,N_19514);
and UO_763 (O_763,N_19601,N_19704);
nand UO_764 (O_764,N_19579,N_19580);
and UO_765 (O_765,N_19717,N_19743);
or UO_766 (O_766,N_19578,N_19948);
and UO_767 (O_767,N_19977,N_19740);
nor UO_768 (O_768,N_19501,N_19569);
nand UO_769 (O_769,N_19665,N_19842);
xnor UO_770 (O_770,N_19510,N_19527);
nand UO_771 (O_771,N_19761,N_19578);
xor UO_772 (O_772,N_19520,N_19726);
or UO_773 (O_773,N_19622,N_19777);
and UO_774 (O_774,N_19715,N_19850);
nor UO_775 (O_775,N_19714,N_19959);
nor UO_776 (O_776,N_19979,N_19548);
xor UO_777 (O_777,N_19654,N_19718);
nand UO_778 (O_778,N_19652,N_19873);
and UO_779 (O_779,N_19803,N_19690);
and UO_780 (O_780,N_19707,N_19680);
xor UO_781 (O_781,N_19515,N_19652);
xnor UO_782 (O_782,N_19662,N_19680);
nor UO_783 (O_783,N_19990,N_19543);
nand UO_784 (O_784,N_19926,N_19625);
and UO_785 (O_785,N_19580,N_19741);
nor UO_786 (O_786,N_19577,N_19759);
nor UO_787 (O_787,N_19859,N_19965);
nor UO_788 (O_788,N_19893,N_19915);
xnor UO_789 (O_789,N_19914,N_19614);
or UO_790 (O_790,N_19776,N_19715);
or UO_791 (O_791,N_19707,N_19659);
xor UO_792 (O_792,N_19530,N_19566);
or UO_793 (O_793,N_19587,N_19537);
and UO_794 (O_794,N_19581,N_19921);
nor UO_795 (O_795,N_19778,N_19984);
or UO_796 (O_796,N_19910,N_19654);
and UO_797 (O_797,N_19755,N_19602);
and UO_798 (O_798,N_19511,N_19966);
xnor UO_799 (O_799,N_19644,N_19545);
nand UO_800 (O_800,N_19581,N_19586);
or UO_801 (O_801,N_19746,N_19845);
nand UO_802 (O_802,N_19961,N_19617);
nor UO_803 (O_803,N_19829,N_19516);
or UO_804 (O_804,N_19602,N_19964);
and UO_805 (O_805,N_19511,N_19877);
nand UO_806 (O_806,N_19725,N_19613);
and UO_807 (O_807,N_19766,N_19533);
nor UO_808 (O_808,N_19626,N_19973);
nand UO_809 (O_809,N_19725,N_19631);
nand UO_810 (O_810,N_19908,N_19925);
nor UO_811 (O_811,N_19537,N_19689);
nand UO_812 (O_812,N_19956,N_19580);
nor UO_813 (O_813,N_19554,N_19512);
and UO_814 (O_814,N_19892,N_19529);
or UO_815 (O_815,N_19868,N_19825);
nor UO_816 (O_816,N_19529,N_19530);
nand UO_817 (O_817,N_19541,N_19933);
and UO_818 (O_818,N_19978,N_19884);
and UO_819 (O_819,N_19939,N_19705);
nor UO_820 (O_820,N_19578,N_19705);
or UO_821 (O_821,N_19530,N_19852);
nand UO_822 (O_822,N_19800,N_19879);
nor UO_823 (O_823,N_19897,N_19813);
xor UO_824 (O_824,N_19769,N_19616);
or UO_825 (O_825,N_19508,N_19862);
xor UO_826 (O_826,N_19654,N_19891);
xor UO_827 (O_827,N_19979,N_19818);
xor UO_828 (O_828,N_19888,N_19537);
xnor UO_829 (O_829,N_19920,N_19701);
xnor UO_830 (O_830,N_19982,N_19873);
nor UO_831 (O_831,N_19872,N_19948);
and UO_832 (O_832,N_19711,N_19890);
xnor UO_833 (O_833,N_19547,N_19552);
nand UO_834 (O_834,N_19990,N_19997);
nand UO_835 (O_835,N_19928,N_19712);
nand UO_836 (O_836,N_19989,N_19575);
and UO_837 (O_837,N_19722,N_19865);
or UO_838 (O_838,N_19562,N_19763);
xnor UO_839 (O_839,N_19969,N_19628);
or UO_840 (O_840,N_19781,N_19854);
xnor UO_841 (O_841,N_19809,N_19980);
or UO_842 (O_842,N_19981,N_19725);
nor UO_843 (O_843,N_19841,N_19680);
nand UO_844 (O_844,N_19961,N_19840);
xnor UO_845 (O_845,N_19601,N_19911);
nand UO_846 (O_846,N_19820,N_19630);
xnor UO_847 (O_847,N_19801,N_19759);
nand UO_848 (O_848,N_19804,N_19773);
nor UO_849 (O_849,N_19804,N_19530);
nand UO_850 (O_850,N_19708,N_19638);
and UO_851 (O_851,N_19512,N_19623);
xor UO_852 (O_852,N_19948,N_19816);
or UO_853 (O_853,N_19782,N_19821);
nor UO_854 (O_854,N_19733,N_19901);
or UO_855 (O_855,N_19913,N_19727);
nor UO_856 (O_856,N_19859,N_19658);
and UO_857 (O_857,N_19562,N_19950);
nor UO_858 (O_858,N_19984,N_19820);
nand UO_859 (O_859,N_19784,N_19845);
nor UO_860 (O_860,N_19687,N_19947);
xnor UO_861 (O_861,N_19521,N_19939);
nor UO_862 (O_862,N_19669,N_19666);
or UO_863 (O_863,N_19671,N_19820);
nor UO_864 (O_864,N_19878,N_19632);
nor UO_865 (O_865,N_19822,N_19793);
or UO_866 (O_866,N_19717,N_19872);
nand UO_867 (O_867,N_19504,N_19555);
xnor UO_868 (O_868,N_19894,N_19696);
and UO_869 (O_869,N_19532,N_19771);
nor UO_870 (O_870,N_19674,N_19919);
nor UO_871 (O_871,N_19558,N_19838);
nand UO_872 (O_872,N_19752,N_19875);
nor UO_873 (O_873,N_19606,N_19587);
or UO_874 (O_874,N_19555,N_19805);
and UO_875 (O_875,N_19710,N_19609);
nand UO_876 (O_876,N_19610,N_19599);
xnor UO_877 (O_877,N_19817,N_19954);
and UO_878 (O_878,N_19605,N_19662);
nand UO_879 (O_879,N_19944,N_19756);
or UO_880 (O_880,N_19986,N_19746);
xnor UO_881 (O_881,N_19589,N_19682);
xor UO_882 (O_882,N_19951,N_19517);
or UO_883 (O_883,N_19552,N_19692);
xnor UO_884 (O_884,N_19979,N_19917);
and UO_885 (O_885,N_19668,N_19691);
and UO_886 (O_886,N_19945,N_19689);
and UO_887 (O_887,N_19954,N_19752);
or UO_888 (O_888,N_19757,N_19786);
nand UO_889 (O_889,N_19729,N_19567);
and UO_890 (O_890,N_19853,N_19869);
and UO_891 (O_891,N_19909,N_19538);
nor UO_892 (O_892,N_19984,N_19953);
nor UO_893 (O_893,N_19579,N_19662);
xor UO_894 (O_894,N_19781,N_19579);
xnor UO_895 (O_895,N_19876,N_19724);
nand UO_896 (O_896,N_19554,N_19662);
nor UO_897 (O_897,N_19645,N_19604);
nor UO_898 (O_898,N_19998,N_19911);
and UO_899 (O_899,N_19631,N_19800);
or UO_900 (O_900,N_19697,N_19787);
nand UO_901 (O_901,N_19597,N_19549);
xnor UO_902 (O_902,N_19852,N_19507);
nand UO_903 (O_903,N_19625,N_19832);
or UO_904 (O_904,N_19745,N_19753);
nor UO_905 (O_905,N_19849,N_19645);
nor UO_906 (O_906,N_19648,N_19597);
xor UO_907 (O_907,N_19626,N_19531);
nor UO_908 (O_908,N_19645,N_19563);
nor UO_909 (O_909,N_19816,N_19935);
nand UO_910 (O_910,N_19724,N_19548);
and UO_911 (O_911,N_19525,N_19861);
or UO_912 (O_912,N_19843,N_19501);
xnor UO_913 (O_913,N_19786,N_19615);
nand UO_914 (O_914,N_19846,N_19572);
nand UO_915 (O_915,N_19831,N_19735);
or UO_916 (O_916,N_19880,N_19584);
and UO_917 (O_917,N_19757,N_19828);
xnor UO_918 (O_918,N_19530,N_19673);
or UO_919 (O_919,N_19814,N_19897);
nor UO_920 (O_920,N_19975,N_19872);
xor UO_921 (O_921,N_19862,N_19996);
and UO_922 (O_922,N_19634,N_19783);
or UO_923 (O_923,N_19889,N_19810);
xnor UO_924 (O_924,N_19557,N_19584);
nor UO_925 (O_925,N_19898,N_19759);
or UO_926 (O_926,N_19865,N_19931);
nand UO_927 (O_927,N_19704,N_19966);
xnor UO_928 (O_928,N_19981,N_19670);
nand UO_929 (O_929,N_19733,N_19974);
or UO_930 (O_930,N_19820,N_19512);
and UO_931 (O_931,N_19651,N_19701);
and UO_932 (O_932,N_19611,N_19963);
or UO_933 (O_933,N_19525,N_19753);
or UO_934 (O_934,N_19761,N_19827);
or UO_935 (O_935,N_19552,N_19775);
or UO_936 (O_936,N_19849,N_19558);
nor UO_937 (O_937,N_19747,N_19985);
nand UO_938 (O_938,N_19678,N_19573);
or UO_939 (O_939,N_19586,N_19899);
or UO_940 (O_940,N_19730,N_19993);
nand UO_941 (O_941,N_19719,N_19795);
or UO_942 (O_942,N_19625,N_19644);
nor UO_943 (O_943,N_19916,N_19690);
nor UO_944 (O_944,N_19801,N_19704);
and UO_945 (O_945,N_19874,N_19966);
and UO_946 (O_946,N_19687,N_19758);
nor UO_947 (O_947,N_19771,N_19721);
nor UO_948 (O_948,N_19826,N_19967);
and UO_949 (O_949,N_19644,N_19860);
or UO_950 (O_950,N_19698,N_19599);
xor UO_951 (O_951,N_19687,N_19977);
or UO_952 (O_952,N_19609,N_19522);
and UO_953 (O_953,N_19691,N_19597);
nand UO_954 (O_954,N_19874,N_19814);
and UO_955 (O_955,N_19664,N_19948);
or UO_956 (O_956,N_19665,N_19829);
and UO_957 (O_957,N_19506,N_19979);
nor UO_958 (O_958,N_19505,N_19963);
nor UO_959 (O_959,N_19972,N_19764);
nand UO_960 (O_960,N_19986,N_19987);
nand UO_961 (O_961,N_19723,N_19570);
nor UO_962 (O_962,N_19640,N_19770);
or UO_963 (O_963,N_19655,N_19946);
or UO_964 (O_964,N_19528,N_19757);
xnor UO_965 (O_965,N_19621,N_19685);
nand UO_966 (O_966,N_19563,N_19959);
and UO_967 (O_967,N_19941,N_19763);
nand UO_968 (O_968,N_19658,N_19669);
nand UO_969 (O_969,N_19521,N_19921);
xor UO_970 (O_970,N_19892,N_19791);
xor UO_971 (O_971,N_19613,N_19743);
and UO_972 (O_972,N_19958,N_19550);
nand UO_973 (O_973,N_19959,N_19605);
nand UO_974 (O_974,N_19796,N_19950);
nand UO_975 (O_975,N_19639,N_19738);
and UO_976 (O_976,N_19686,N_19825);
xor UO_977 (O_977,N_19572,N_19605);
nand UO_978 (O_978,N_19996,N_19958);
and UO_979 (O_979,N_19943,N_19990);
xnor UO_980 (O_980,N_19970,N_19831);
and UO_981 (O_981,N_19577,N_19562);
and UO_982 (O_982,N_19753,N_19817);
or UO_983 (O_983,N_19850,N_19548);
nor UO_984 (O_984,N_19514,N_19598);
and UO_985 (O_985,N_19950,N_19934);
nand UO_986 (O_986,N_19502,N_19859);
and UO_987 (O_987,N_19945,N_19825);
nand UO_988 (O_988,N_19860,N_19892);
xor UO_989 (O_989,N_19615,N_19612);
and UO_990 (O_990,N_19634,N_19651);
or UO_991 (O_991,N_19983,N_19888);
nand UO_992 (O_992,N_19940,N_19697);
nor UO_993 (O_993,N_19745,N_19774);
xnor UO_994 (O_994,N_19671,N_19754);
and UO_995 (O_995,N_19639,N_19679);
or UO_996 (O_996,N_19740,N_19868);
xor UO_997 (O_997,N_19729,N_19882);
or UO_998 (O_998,N_19853,N_19634);
nand UO_999 (O_999,N_19675,N_19997);
or UO_1000 (O_1000,N_19579,N_19796);
nor UO_1001 (O_1001,N_19903,N_19673);
nor UO_1002 (O_1002,N_19921,N_19886);
xnor UO_1003 (O_1003,N_19549,N_19939);
xor UO_1004 (O_1004,N_19828,N_19756);
and UO_1005 (O_1005,N_19925,N_19736);
nor UO_1006 (O_1006,N_19825,N_19816);
or UO_1007 (O_1007,N_19708,N_19511);
nor UO_1008 (O_1008,N_19587,N_19767);
and UO_1009 (O_1009,N_19887,N_19688);
xnor UO_1010 (O_1010,N_19582,N_19949);
nor UO_1011 (O_1011,N_19893,N_19656);
nor UO_1012 (O_1012,N_19802,N_19545);
nand UO_1013 (O_1013,N_19536,N_19961);
xor UO_1014 (O_1014,N_19764,N_19528);
xnor UO_1015 (O_1015,N_19535,N_19622);
xnor UO_1016 (O_1016,N_19663,N_19531);
xnor UO_1017 (O_1017,N_19509,N_19693);
or UO_1018 (O_1018,N_19732,N_19666);
nor UO_1019 (O_1019,N_19677,N_19874);
nor UO_1020 (O_1020,N_19975,N_19706);
nor UO_1021 (O_1021,N_19921,N_19603);
and UO_1022 (O_1022,N_19553,N_19928);
xor UO_1023 (O_1023,N_19560,N_19881);
nand UO_1024 (O_1024,N_19722,N_19999);
xor UO_1025 (O_1025,N_19710,N_19964);
or UO_1026 (O_1026,N_19813,N_19807);
nand UO_1027 (O_1027,N_19731,N_19553);
nor UO_1028 (O_1028,N_19788,N_19813);
xor UO_1029 (O_1029,N_19667,N_19807);
nor UO_1030 (O_1030,N_19576,N_19812);
nor UO_1031 (O_1031,N_19543,N_19930);
and UO_1032 (O_1032,N_19966,N_19519);
and UO_1033 (O_1033,N_19655,N_19755);
xor UO_1034 (O_1034,N_19960,N_19687);
and UO_1035 (O_1035,N_19738,N_19990);
nand UO_1036 (O_1036,N_19951,N_19861);
nor UO_1037 (O_1037,N_19588,N_19707);
xnor UO_1038 (O_1038,N_19629,N_19714);
nor UO_1039 (O_1039,N_19540,N_19741);
nor UO_1040 (O_1040,N_19702,N_19876);
nand UO_1041 (O_1041,N_19716,N_19879);
xnor UO_1042 (O_1042,N_19904,N_19699);
and UO_1043 (O_1043,N_19891,N_19510);
nor UO_1044 (O_1044,N_19603,N_19569);
or UO_1045 (O_1045,N_19629,N_19528);
and UO_1046 (O_1046,N_19715,N_19802);
and UO_1047 (O_1047,N_19546,N_19657);
xor UO_1048 (O_1048,N_19592,N_19682);
nor UO_1049 (O_1049,N_19615,N_19735);
or UO_1050 (O_1050,N_19749,N_19729);
nor UO_1051 (O_1051,N_19729,N_19928);
xor UO_1052 (O_1052,N_19829,N_19914);
nor UO_1053 (O_1053,N_19804,N_19754);
or UO_1054 (O_1054,N_19737,N_19989);
xor UO_1055 (O_1055,N_19786,N_19655);
or UO_1056 (O_1056,N_19964,N_19879);
nand UO_1057 (O_1057,N_19680,N_19552);
nor UO_1058 (O_1058,N_19611,N_19886);
nand UO_1059 (O_1059,N_19674,N_19747);
or UO_1060 (O_1060,N_19877,N_19757);
xor UO_1061 (O_1061,N_19884,N_19920);
xor UO_1062 (O_1062,N_19636,N_19500);
and UO_1063 (O_1063,N_19622,N_19780);
nor UO_1064 (O_1064,N_19847,N_19866);
nand UO_1065 (O_1065,N_19605,N_19797);
nor UO_1066 (O_1066,N_19637,N_19875);
nor UO_1067 (O_1067,N_19693,N_19665);
and UO_1068 (O_1068,N_19822,N_19577);
nor UO_1069 (O_1069,N_19963,N_19690);
nor UO_1070 (O_1070,N_19902,N_19687);
and UO_1071 (O_1071,N_19949,N_19671);
nand UO_1072 (O_1072,N_19515,N_19797);
and UO_1073 (O_1073,N_19536,N_19589);
xor UO_1074 (O_1074,N_19588,N_19578);
nor UO_1075 (O_1075,N_19965,N_19923);
xor UO_1076 (O_1076,N_19586,N_19715);
and UO_1077 (O_1077,N_19561,N_19641);
and UO_1078 (O_1078,N_19542,N_19648);
and UO_1079 (O_1079,N_19958,N_19893);
xnor UO_1080 (O_1080,N_19835,N_19780);
xor UO_1081 (O_1081,N_19542,N_19909);
and UO_1082 (O_1082,N_19607,N_19719);
nand UO_1083 (O_1083,N_19791,N_19665);
xnor UO_1084 (O_1084,N_19787,N_19549);
nor UO_1085 (O_1085,N_19936,N_19956);
or UO_1086 (O_1086,N_19568,N_19822);
xnor UO_1087 (O_1087,N_19955,N_19719);
and UO_1088 (O_1088,N_19733,N_19515);
and UO_1089 (O_1089,N_19856,N_19736);
nor UO_1090 (O_1090,N_19655,N_19607);
or UO_1091 (O_1091,N_19870,N_19700);
and UO_1092 (O_1092,N_19996,N_19653);
nor UO_1093 (O_1093,N_19580,N_19880);
xor UO_1094 (O_1094,N_19665,N_19801);
and UO_1095 (O_1095,N_19829,N_19546);
xor UO_1096 (O_1096,N_19800,N_19994);
nor UO_1097 (O_1097,N_19780,N_19741);
xnor UO_1098 (O_1098,N_19570,N_19756);
nand UO_1099 (O_1099,N_19847,N_19938);
nand UO_1100 (O_1100,N_19825,N_19538);
and UO_1101 (O_1101,N_19666,N_19942);
or UO_1102 (O_1102,N_19503,N_19810);
or UO_1103 (O_1103,N_19822,N_19606);
nor UO_1104 (O_1104,N_19890,N_19812);
nor UO_1105 (O_1105,N_19724,N_19743);
or UO_1106 (O_1106,N_19665,N_19979);
xor UO_1107 (O_1107,N_19870,N_19740);
and UO_1108 (O_1108,N_19680,N_19514);
xnor UO_1109 (O_1109,N_19500,N_19741);
or UO_1110 (O_1110,N_19575,N_19732);
xnor UO_1111 (O_1111,N_19983,N_19502);
xor UO_1112 (O_1112,N_19558,N_19716);
or UO_1113 (O_1113,N_19818,N_19636);
nand UO_1114 (O_1114,N_19787,N_19609);
nor UO_1115 (O_1115,N_19950,N_19517);
nor UO_1116 (O_1116,N_19804,N_19956);
or UO_1117 (O_1117,N_19736,N_19501);
or UO_1118 (O_1118,N_19861,N_19711);
nor UO_1119 (O_1119,N_19569,N_19823);
and UO_1120 (O_1120,N_19902,N_19976);
xor UO_1121 (O_1121,N_19663,N_19929);
nor UO_1122 (O_1122,N_19841,N_19503);
or UO_1123 (O_1123,N_19786,N_19512);
nand UO_1124 (O_1124,N_19631,N_19639);
xor UO_1125 (O_1125,N_19791,N_19750);
nand UO_1126 (O_1126,N_19676,N_19765);
or UO_1127 (O_1127,N_19959,N_19533);
or UO_1128 (O_1128,N_19819,N_19724);
xnor UO_1129 (O_1129,N_19865,N_19871);
or UO_1130 (O_1130,N_19758,N_19838);
nor UO_1131 (O_1131,N_19771,N_19604);
and UO_1132 (O_1132,N_19652,N_19891);
and UO_1133 (O_1133,N_19708,N_19810);
nor UO_1134 (O_1134,N_19820,N_19929);
nor UO_1135 (O_1135,N_19517,N_19816);
nand UO_1136 (O_1136,N_19879,N_19931);
and UO_1137 (O_1137,N_19500,N_19597);
nor UO_1138 (O_1138,N_19719,N_19940);
nand UO_1139 (O_1139,N_19761,N_19743);
nor UO_1140 (O_1140,N_19588,N_19599);
xor UO_1141 (O_1141,N_19922,N_19774);
and UO_1142 (O_1142,N_19534,N_19651);
or UO_1143 (O_1143,N_19639,N_19557);
xnor UO_1144 (O_1144,N_19702,N_19849);
nand UO_1145 (O_1145,N_19604,N_19636);
nand UO_1146 (O_1146,N_19806,N_19965);
nand UO_1147 (O_1147,N_19977,N_19645);
or UO_1148 (O_1148,N_19590,N_19753);
xnor UO_1149 (O_1149,N_19814,N_19872);
xnor UO_1150 (O_1150,N_19678,N_19767);
nor UO_1151 (O_1151,N_19619,N_19668);
or UO_1152 (O_1152,N_19640,N_19729);
or UO_1153 (O_1153,N_19962,N_19697);
nand UO_1154 (O_1154,N_19741,N_19692);
xor UO_1155 (O_1155,N_19885,N_19513);
xor UO_1156 (O_1156,N_19930,N_19697);
or UO_1157 (O_1157,N_19668,N_19649);
and UO_1158 (O_1158,N_19566,N_19550);
and UO_1159 (O_1159,N_19840,N_19862);
nand UO_1160 (O_1160,N_19830,N_19939);
nor UO_1161 (O_1161,N_19659,N_19722);
or UO_1162 (O_1162,N_19935,N_19558);
and UO_1163 (O_1163,N_19780,N_19737);
nor UO_1164 (O_1164,N_19981,N_19830);
or UO_1165 (O_1165,N_19653,N_19550);
xor UO_1166 (O_1166,N_19528,N_19948);
nand UO_1167 (O_1167,N_19723,N_19865);
nor UO_1168 (O_1168,N_19557,N_19610);
nor UO_1169 (O_1169,N_19804,N_19588);
or UO_1170 (O_1170,N_19567,N_19601);
or UO_1171 (O_1171,N_19726,N_19944);
or UO_1172 (O_1172,N_19690,N_19598);
xnor UO_1173 (O_1173,N_19601,N_19542);
nor UO_1174 (O_1174,N_19572,N_19739);
or UO_1175 (O_1175,N_19862,N_19605);
nand UO_1176 (O_1176,N_19877,N_19738);
nand UO_1177 (O_1177,N_19598,N_19991);
nand UO_1178 (O_1178,N_19720,N_19622);
and UO_1179 (O_1179,N_19709,N_19564);
and UO_1180 (O_1180,N_19617,N_19880);
xnor UO_1181 (O_1181,N_19690,N_19535);
or UO_1182 (O_1182,N_19622,N_19650);
xor UO_1183 (O_1183,N_19872,N_19854);
and UO_1184 (O_1184,N_19571,N_19629);
nor UO_1185 (O_1185,N_19889,N_19659);
and UO_1186 (O_1186,N_19518,N_19541);
xnor UO_1187 (O_1187,N_19875,N_19912);
nand UO_1188 (O_1188,N_19540,N_19974);
nor UO_1189 (O_1189,N_19505,N_19943);
nand UO_1190 (O_1190,N_19607,N_19553);
nand UO_1191 (O_1191,N_19570,N_19744);
nor UO_1192 (O_1192,N_19933,N_19815);
and UO_1193 (O_1193,N_19678,N_19532);
xnor UO_1194 (O_1194,N_19710,N_19627);
or UO_1195 (O_1195,N_19979,N_19508);
and UO_1196 (O_1196,N_19709,N_19517);
nand UO_1197 (O_1197,N_19858,N_19750);
nand UO_1198 (O_1198,N_19995,N_19552);
nand UO_1199 (O_1199,N_19534,N_19628);
nand UO_1200 (O_1200,N_19919,N_19922);
xnor UO_1201 (O_1201,N_19634,N_19760);
or UO_1202 (O_1202,N_19858,N_19708);
xnor UO_1203 (O_1203,N_19604,N_19662);
and UO_1204 (O_1204,N_19672,N_19884);
or UO_1205 (O_1205,N_19982,N_19576);
xor UO_1206 (O_1206,N_19924,N_19867);
or UO_1207 (O_1207,N_19788,N_19629);
nand UO_1208 (O_1208,N_19826,N_19954);
xnor UO_1209 (O_1209,N_19925,N_19593);
or UO_1210 (O_1210,N_19594,N_19758);
nand UO_1211 (O_1211,N_19974,N_19897);
nand UO_1212 (O_1212,N_19757,N_19803);
and UO_1213 (O_1213,N_19782,N_19942);
or UO_1214 (O_1214,N_19976,N_19845);
xnor UO_1215 (O_1215,N_19612,N_19512);
nand UO_1216 (O_1216,N_19943,N_19775);
and UO_1217 (O_1217,N_19825,N_19813);
nor UO_1218 (O_1218,N_19712,N_19933);
or UO_1219 (O_1219,N_19923,N_19693);
and UO_1220 (O_1220,N_19665,N_19681);
nand UO_1221 (O_1221,N_19887,N_19616);
or UO_1222 (O_1222,N_19994,N_19630);
or UO_1223 (O_1223,N_19794,N_19896);
xor UO_1224 (O_1224,N_19915,N_19857);
and UO_1225 (O_1225,N_19821,N_19762);
or UO_1226 (O_1226,N_19948,N_19920);
xnor UO_1227 (O_1227,N_19945,N_19714);
and UO_1228 (O_1228,N_19664,N_19518);
xnor UO_1229 (O_1229,N_19960,N_19679);
or UO_1230 (O_1230,N_19891,N_19555);
nor UO_1231 (O_1231,N_19507,N_19729);
or UO_1232 (O_1232,N_19910,N_19875);
nor UO_1233 (O_1233,N_19852,N_19506);
xor UO_1234 (O_1234,N_19566,N_19529);
or UO_1235 (O_1235,N_19711,N_19744);
and UO_1236 (O_1236,N_19877,N_19847);
nor UO_1237 (O_1237,N_19773,N_19598);
or UO_1238 (O_1238,N_19599,N_19873);
or UO_1239 (O_1239,N_19507,N_19518);
or UO_1240 (O_1240,N_19626,N_19651);
nor UO_1241 (O_1241,N_19986,N_19672);
and UO_1242 (O_1242,N_19577,N_19669);
nand UO_1243 (O_1243,N_19833,N_19938);
nor UO_1244 (O_1244,N_19950,N_19597);
or UO_1245 (O_1245,N_19513,N_19694);
nand UO_1246 (O_1246,N_19522,N_19869);
or UO_1247 (O_1247,N_19938,N_19911);
and UO_1248 (O_1248,N_19794,N_19835);
and UO_1249 (O_1249,N_19737,N_19789);
nor UO_1250 (O_1250,N_19728,N_19865);
nand UO_1251 (O_1251,N_19980,N_19988);
or UO_1252 (O_1252,N_19986,N_19846);
xnor UO_1253 (O_1253,N_19822,N_19708);
xnor UO_1254 (O_1254,N_19740,N_19555);
or UO_1255 (O_1255,N_19559,N_19520);
nand UO_1256 (O_1256,N_19724,N_19964);
nand UO_1257 (O_1257,N_19660,N_19507);
nand UO_1258 (O_1258,N_19794,N_19697);
and UO_1259 (O_1259,N_19812,N_19619);
nor UO_1260 (O_1260,N_19839,N_19771);
xnor UO_1261 (O_1261,N_19606,N_19789);
or UO_1262 (O_1262,N_19993,N_19957);
nand UO_1263 (O_1263,N_19536,N_19741);
and UO_1264 (O_1264,N_19701,N_19806);
nor UO_1265 (O_1265,N_19776,N_19547);
nor UO_1266 (O_1266,N_19881,N_19622);
nor UO_1267 (O_1267,N_19815,N_19643);
nand UO_1268 (O_1268,N_19998,N_19653);
nand UO_1269 (O_1269,N_19636,N_19944);
and UO_1270 (O_1270,N_19532,N_19671);
and UO_1271 (O_1271,N_19973,N_19713);
xor UO_1272 (O_1272,N_19839,N_19505);
nand UO_1273 (O_1273,N_19973,N_19943);
and UO_1274 (O_1274,N_19706,N_19913);
and UO_1275 (O_1275,N_19987,N_19674);
or UO_1276 (O_1276,N_19877,N_19973);
or UO_1277 (O_1277,N_19691,N_19897);
nand UO_1278 (O_1278,N_19841,N_19546);
nand UO_1279 (O_1279,N_19722,N_19755);
nor UO_1280 (O_1280,N_19693,N_19960);
xor UO_1281 (O_1281,N_19586,N_19602);
and UO_1282 (O_1282,N_19694,N_19971);
or UO_1283 (O_1283,N_19708,N_19619);
or UO_1284 (O_1284,N_19610,N_19854);
nor UO_1285 (O_1285,N_19611,N_19659);
xor UO_1286 (O_1286,N_19570,N_19911);
xor UO_1287 (O_1287,N_19583,N_19771);
and UO_1288 (O_1288,N_19850,N_19673);
and UO_1289 (O_1289,N_19834,N_19725);
and UO_1290 (O_1290,N_19826,N_19636);
nor UO_1291 (O_1291,N_19774,N_19663);
and UO_1292 (O_1292,N_19915,N_19774);
or UO_1293 (O_1293,N_19735,N_19577);
and UO_1294 (O_1294,N_19895,N_19577);
xor UO_1295 (O_1295,N_19811,N_19544);
xnor UO_1296 (O_1296,N_19669,N_19988);
and UO_1297 (O_1297,N_19897,N_19600);
nand UO_1298 (O_1298,N_19822,N_19671);
and UO_1299 (O_1299,N_19744,N_19710);
or UO_1300 (O_1300,N_19747,N_19917);
xnor UO_1301 (O_1301,N_19938,N_19748);
xor UO_1302 (O_1302,N_19589,N_19880);
xnor UO_1303 (O_1303,N_19888,N_19802);
nor UO_1304 (O_1304,N_19929,N_19756);
or UO_1305 (O_1305,N_19519,N_19744);
and UO_1306 (O_1306,N_19975,N_19510);
or UO_1307 (O_1307,N_19988,N_19709);
or UO_1308 (O_1308,N_19834,N_19651);
nor UO_1309 (O_1309,N_19571,N_19802);
nor UO_1310 (O_1310,N_19652,N_19583);
and UO_1311 (O_1311,N_19594,N_19728);
or UO_1312 (O_1312,N_19599,N_19642);
xor UO_1313 (O_1313,N_19827,N_19816);
nand UO_1314 (O_1314,N_19941,N_19621);
and UO_1315 (O_1315,N_19935,N_19875);
and UO_1316 (O_1316,N_19926,N_19998);
or UO_1317 (O_1317,N_19572,N_19509);
or UO_1318 (O_1318,N_19651,N_19510);
nor UO_1319 (O_1319,N_19892,N_19504);
xor UO_1320 (O_1320,N_19626,N_19590);
nor UO_1321 (O_1321,N_19846,N_19712);
nor UO_1322 (O_1322,N_19806,N_19795);
or UO_1323 (O_1323,N_19854,N_19701);
xnor UO_1324 (O_1324,N_19887,N_19540);
nor UO_1325 (O_1325,N_19810,N_19557);
xor UO_1326 (O_1326,N_19609,N_19855);
xor UO_1327 (O_1327,N_19740,N_19586);
nor UO_1328 (O_1328,N_19626,N_19933);
xnor UO_1329 (O_1329,N_19670,N_19579);
xnor UO_1330 (O_1330,N_19522,N_19590);
nor UO_1331 (O_1331,N_19637,N_19730);
nand UO_1332 (O_1332,N_19852,N_19592);
xnor UO_1333 (O_1333,N_19578,N_19989);
or UO_1334 (O_1334,N_19613,N_19911);
or UO_1335 (O_1335,N_19900,N_19937);
nand UO_1336 (O_1336,N_19955,N_19978);
or UO_1337 (O_1337,N_19749,N_19844);
nor UO_1338 (O_1338,N_19932,N_19515);
or UO_1339 (O_1339,N_19930,N_19923);
nand UO_1340 (O_1340,N_19772,N_19799);
xor UO_1341 (O_1341,N_19821,N_19941);
or UO_1342 (O_1342,N_19761,N_19837);
or UO_1343 (O_1343,N_19710,N_19537);
xnor UO_1344 (O_1344,N_19532,N_19735);
or UO_1345 (O_1345,N_19579,N_19525);
nor UO_1346 (O_1346,N_19938,N_19671);
nand UO_1347 (O_1347,N_19900,N_19709);
and UO_1348 (O_1348,N_19634,N_19998);
or UO_1349 (O_1349,N_19871,N_19995);
and UO_1350 (O_1350,N_19537,N_19854);
nor UO_1351 (O_1351,N_19902,N_19592);
nand UO_1352 (O_1352,N_19663,N_19816);
nor UO_1353 (O_1353,N_19689,N_19870);
nor UO_1354 (O_1354,N_19568,N_19564);
or UO_1355 (O_1355,N_19738,N_19894);
and UO_1356 (O_1356,N_19755,N_19527);
or UO_1357 (O_1357,N_19649,N_19939);
nand UO_1358 (O_1358,N_19657,N_19692);
and UO_1359 (O_1359,N_19578,N_19508);
or UO_1360 (O_1360,N_19526,N_19591);
xor UO_1361 (O_1361,N_19735,N_19638);
xnor UO_1362 (O_1362,N_19833,N_19702);
or UO_1363 (O_1363,N_19782,N_19621);
nand UO_1364 (O_1364,N_19685,N_19754);
nor UO_1365 (O_1365,N_19894,N_19523);
xnor UO_1366 (O_1366,N_19531,N_19859);
or UO_1367 (O_1367,N_19742,N_19599);
and UO_1368 (O_1368,N_19669,N_19506);
and UO_1369 (O_1369,N_19965,N_19845);
or UO_1370 (O_1370,N_19701,N_19569);
and UO_1371 (O_1371,N_19685,N_19599);
and UO_1372 (O_1372,N_19617,N_19821);
or UO_1373 (O_1373,N_19607,N_19827);
xor UO_1374 (O_1374,N_19708,N_19973);
and UO_1375 (O_1375,N_19673,N_19575);
xnor UO_1376 (O_1376,N_19873,N_19581);
or UO_1377 (O_1377,N_19554,N_19853);
xnor UO_1378 (O_1378,N_19975,N_19586);
xor UO_1379 (O_1379,N_19777,N_19683);
nor UO_1380 (O_1380,N_19528,N_19961);
nand UO_1381 (O_1381,N_19910,N_19812);
or UO_1382 (O_1382,N_19748,N_19696);
or UO_1383 (O_1383,N_19831,N_19993);
and UO_1384 (O_1384,N_19596,N_19686);
or UO_1385 (O_1385,N_19839,N_19864);
nand UO_1386 (O_1386,N_19975,N_19876);
nand UO_1387 (O_1387,N_19972,N_19930);
or UO_1388 (O_1388,N_19592,N_19927);
or UO_1389 (O_1389,N_19788,N_19843);
xor UO_1390 (O_1390,N_19993,N_19749);
nand UO_1391 (O_1391,N_19852,N_19720);
nor UO_1392 (O_1392,N_19523,N_19877);
nand UO_1393 (O_1393,N_19639,N_19722);
xnor UO_1394 (O_1394,N_19603,N_19990);
or UO_1395 (O_1395,N_19954,N_19531);
nor UO_1396 (O_1396,N_19675,N_19896);
nor UO_1397 (O_1397,N_19939,N_19596);
nand UO_1398 (O_1398,N_19870,N_19818);
xnor UO_1399 (O_1399,N_19773,N_19601);
and UO_1400 (O_1400,N_19543,N_19995);
or UO_1401 (O_1401,N_19747,N_19821);
nor UO_1402 (O_1402,N_19815,N_19619);
nand UO_1403 (O_1403,N_19708,N_19964);
nand UO_1404 (O_1404,N_19890,N_19829);
xor UO_1405 (O_1405,N_19934,N_19579);
or UO_1406 (O_1406,N_19960,N_19545);
nor UO_1407 (O_1407,N_19716,N_19733);
nand UO_1408 (O_1408,N_19834,N_19859);
and UO_1409 (O_1409,N_19604,N_19652);
and UO_1410 (O_1410,N_19969,N_19724);
xnor UO_1411 (O_1411,N_19824,N_19574);
nor UO_1412 (O_1412,N_19940,N_19671);
and UO_1413 (O_1413,N_19644,N_19719);
nor UO_1414 (O_1414,N_19723,N_19894);
and UO_1415 (O_1415,N_19698,N_19883);
nor UO_1416 (O_1416,N_19599,N_19755);
nand UO_1417 (O_1417,N_19563,N_19828);
and UO_1418 (O_1418,N_19996,N_19539);
or UO_1419 (O_1419,N_19851,N_19531);
or UO_1420 (O_1420,N_19945,N_19713);
nor UO_1421 (O_1421,N_19553,N_19821);
nor UO_1422 (O_1422,N_19917,N_19723);
and UO_1423 (O_1423,N_19729,N_19597);
and UO_1424 (O_1424,N_19662,N_19905);
xor UO_1425 (O_1425,N_19880,N_19984);
nor UO_1426 (O_1426,N_19856,N_19710);
nor UO_1427 (O_1427,N_19928,N_19571);
or UO_1428 (O_1428,N_19816,N_19965);
nor UO_1429 (O_1429,N_19831,N_19593);
and UO_1430 (O_1430,N_19573,N_19999);
xnor UO_1431 (O_1431,N_19722,N_19727);
nor UO_1432 (O_1432,N_19834,N_19908);
nor UO_1433 (O_1433,N_19907,N_19519);
nand UO_1434 (O_1434,N_19683,N_19871);
and UO_1435 (O_1435,N_19886,N_19889);
or UO_1436 (O_1436,N_19981,N_19787);
or UO_1437 (O_1437,N_19685,N_19838);
and UO_1438 (O_1438,N_19558,N_19714);
nor UO_1439 (O_1439,N_19721,N_19607);
nor UO_1440 (O_1440,N_19851,N_19616);
nand UO_1441 (O_1441,N_19584,N_19965);
and UO_1442 (O_1442,N_19682,N_19544);
or UO_1443 (O_1443,N_19676,N_19996);
xor UO_1444 (O_1444,N_19719,N_19571);
and UO_1445 (O_1445,N_19834,N_19710);
xor UO_1446 (O_1446,N_19548,N_19813);
or UO_1447 (O_1447,N_19907,N_19516);
or UO_1448 (O_1448,N_19748,N_19807);
nor UO_1449 (O_1449,N_19938,N_19729);
and UO_1450 (O_1450,N_19826,N_19905);
and UO_1451 (O_1451,N_19740,N_19716);
nor UO_1452 (O_1452,N_19888,N_19903);
and UO_1453 (O_1453,N_19612,N_19596);
nand UO_1454 (O_1454,N_19901,N_19730);
nand UO_1455 (O_1455,N_19727,N_19716);
nand UO_1456 (O_1456,N_19634,N_19985);
nand UO_1457 (O_1457,N_19962,N_19921);
xnor UO_1458 (O_1458,N_19528,N_19789);
xor UO_1459 (O_1459,N_19677,N_19846);
xor UO_1460 (O_1460,N_19878,N_19829);
and UO_1461 (O_1461,N_19978,N_19581);
or UO_1462 (O_1462,N_19536,N_19905);
nor UO_1463 (O_1463,N_19986,N_19794);
nand UO_1464 (O_1464,N_19585,N_19851);
nor UO_1465 (O_1465,N_19765,N_19888);
nand UO_1466 (O_1466,N_19900,N_19502);
or UO_1467 (O_1467,N_19801,N_19778);
or UO_1468 (O_1468,N_19693,N_19768);
xor UO_1469 (O_1469,N_19591,N_19973);
nand UO_1470 (O_1470,N_19512,N_19643);
nor UO_1471 (O_1471,N_19909,N_19745);
and UO_1472 (O_1472,N_19856,N_19907);
nand UO_1473 (O_1473,N_19555,N_19918);
nand UO_1474 (O_1474,N_19746,N_19922);
nor UO_1475 (O_1475,N_19907,N_19724);
or UO_1476 (O_1476,N_19754,N_19809);
xnor UO_1477 (O_1477,N_19602,N_19544);
or UO_1478 (O_1478,N_19952,N_19740);
nand UO_1479 (O_1479,N_19535,N_19985);
and UO_1480 (O_1480,N_19661,N_19722);
and UO_1481 (O_1481,N_19951,N_19993);
or UO_1482 (O_1482,N_19792,N_19738);
and UO_1483 (O_1483,N_19512,N_19500);
or UO_1484 (O_1484,N_19910,N_19706);
nor UO_1485 (O_1485,N_19653,N_19775);
and UO_1486 (O_1486,N_19864,N_19909);
nor UO_1487 (O_1487,N_19662,N_19981);
xor UO_1488 (O_1488,N_19731,N_19672);
nor UO_1489 (O_1489,N_19538,N_19955);
nand UO_1490 (O_1490,N_19592,N_19900);
or UO_1491 (O_1491,N_19633,N_19730);
nand UO_1492 (O_1492,N_19601,N_19720);
nand UO_1493 (O_1493,N_19765,N_19874);
and UO_1494 (O_1494,N_19756,N_19859);
or UO_1495 (O_1495,N_19897,N_19999);
nor UO_1496 (O_1496,N_19668,N_19989);
or UO_1497 (O_1497,N_19770,N_19811);
and UO_1498 (O_1498,N_19619,N_19584);
nor UO_1499 (O_1499,N_19641,N_19780);
xnor UO_1500 (O_1500,N_19750,N_19756);
or UO_1501 (O_1501,N_19701,N_19521);
xnor UO_1502 (O_1502,N_19712,N_19772);
or UO_1503 (O_1503,N_19507,N_19523);
nor UO_1504 (O_1504,N_19996,N_19928);
or UO_1505 (O_1505,N_19578,N_19689);
nand UO_1506 (O_1506,N_19717,N_19580);
and UO_1507 (O_1507,N_19782,N_19952);
and UO_1508 (O_1508,N_19989,N_19637);
nand UO_1509 (O_1509,N_19534,N_19786);
nand UO_1510 (O_1510,N_19803,N_19586);
nand UO_1511 (O_1511,N_19929,N_19667);
xor UO_1512 (O_1512,N_19915,N_19527);
and UO_1513 (O_1513,N_19950,N_19889);
xnor UO_1514 (O_1514,N_19810,N_19844);
or UO_1515 (O_1515,N_19694,N_19740);
xnor UO_1516 (O_1516,N_19574,N_19782);
and UO_1517 (O_1517,N_19969,N_19727);
nand UO_1518 (O_1518,N_19719,N_19530);
nor UO_1519 (O_1519,N_19560,N_19777);
nor UO_1520 (O_1520,N_19809,N_19871);
nand UO_1521 (O_1521,N_19800,N_19877);
or UO_1522 (O_1522,N_19953,N_19571);
nand UO_1523 (O_1523,N_19602,N_19637);
and UO_1524 (O_1524,N_19645,N_19605);
nor UO_1525 (O_1525,N_19828,N_19690);
and UO_1526 (O_1526,N_19968,N_19768);
xor UO_1527 (O_1527,N_19719,N_19917);
nor UO_1528 (O_1528,N_19648,N_19671);
xnor UO_1529 (O_1529,N_19602,N_19716);
xor UO_1530 (O_1530,N_19671,N_19591);
and UO_1531 (O_1531,N_19651,N_19600);
nand UO_1532 (O_1532,N_19510,N_19547);
nand UO_1533 (O_1533,N_19921,N_19761);
nor UO_1534 (O_1534,N_19943,N_19812);
nand UO_1535 (O_1535,N_19655,N_19620);
and UO_1536 (O_1536,N_19727,N_19576);
nand UO_1537 (O_1537,N_19646,N_19538);
nor UO_1538 (O_1538,N_19571,N_19579);
xor UO_1539 (O_1539,N_19612,N_19550);
nand UO_1540 (O_1540,N_19693,N_19794);
or UO_1541 (O_1541,N_19880,N_19549);
or UO_1542 (O_1542,N_19526,N_19575);
xor UO_1543 (O_1543,N_19647,N_19739);
xor UO_1544 (O_1544,N_19773,N_19904);
nor UO_1545 (O_1545,N_19698,N_19529);
nor UO_1546 (O_1546,N_19913,N_19597);
and UO_1547 (O_1547,N_19774,N_19573);
or UO_1548 (O_1548,N_19658,N_19684);
or UO_1549 (O_1549,N_19739,N_19814);
nor UO_1550 (O_1550,N_19827,N_19521);
nand UO_1551 (O_1551,N_19634,N_19795);
xnor UO_1552 (O_1552,N_19652,N_19837);
nand UO_1553 (O_1553,N_19903,N_19889);
and UO_1554 (O_1554,N_19898,N_19909);
xnor UO_1555 (O_1555,N_19602,N_19831);
or UO_1556 (O_1556,N_19507,N_19889);
nor UO_1557 (O_1557,N_19639,N_19717);
nand UO_1558 (O_1558,N_19975,N_19875);
and UO_1559 (O_1559,N_19504,N_19627);
nand UO_1560 (O_1560,N_19792,N_19908);
xor UO_1561 (O_1561,N_19591,N_19543);
nand UO_1562 (O_1562,N_19532,N_19599);
and UO_1563 (O_1563,N_19690,N_19814);
and UO_1564 (O_1564,N_19566,N_19688);
nor UO_1565 (O_1565,N_19708,N_19614);
xor UO_1566 (O_1566,N_19543,N_19823);
nor UO_1567 (O_1567,N_19990,N_19507);
or UO_1568 (O_1568,N_19712,N_19560);
xnor UO_1569 (O_1569,N_19754,N_19832);
nor UO_1570 (O_1570,N_19950,N_19994);
xor UO_1571 (O_1571,N_19986,N_19978);
nor UO_1572 (O_1572,N_19813,N_19842);
nand UO_1573 (O_1573,N_19524,N_19552);
and UO_1574 (O_1574,N_19759,N_19523);
xnor UO_1575 (O_1575,N_19856,N_19750);
xor UO_1576 (O_1576,N_19894,N_19768);
xor UO_1577 (O_1577,N_19968,N_19619);
nand UO_1578 (O_1578,N_19700,N_19734);
nor UO_1579 (O_1579,N_19791,N_19529);
nor UO_1580 (O_1580,N_19625,N_19539);
and UO_1581 (O_1581,N_19816,N_19863);
and UO_1582 (O_1582,N_19851,N_19890);
and UO_1583 (O_1583,N_19603,N_19811);
nand UO_1584 (O_1584,N_19898,N_19740);
nor UO_1585 (O_1585,N_19573,N_19520);
and UO_1586 (O_1586,N_19770,N_19869);
or UO_1587 (O_1587,N_19775,N_19806);
nand UO_1588 (O_1588,N_19579,N_19982);
and UO_1589 (O_1589,N_19528,N_19858);
and UO_1590 (O_1590,N_19738,N_19518);
xor UO_1591 (O_1591,N_19665,N_19691);
xnor UO_1592 (O_1592,N_19994,N_19531);
and UO_1593 (O_1593,N_19587,N_19964);
nor UO_1594 (O_1594,N_19842,N_19956);
or UO_1595 (O_1595,N_19872,N_19525);
and UO_1596 (O_1596,N_19911,N_19715);
nor UO_1597 (O_1597,N_19637,N_19965);
nand UO_1598 (O_1598,N_19849,N_19721);
nor UO_1599 (O_1599,N_19633,N_19870);
or UO_1600 (O_1600,N_19616,N_19591);
nor UO_1601 (O_1601,N_19669,N_19853);
xor UO_1602 (O_1602,N_19937,N_19979);
and UO_1603 (O_1603,N_19532,N_19819);
nor UO_1604 (O_1604,N_19841,N_19957);
or UO_1605 (O_1605,N_19927,N_19588);
nand UO_1606 (O_1606,N_19932,N_19860);
nor UO_1607 (O_1607,N_19794,N_19798);
nor UO_1608 (O_1608,N_19789,N_19795);
or UO_1609 (O_1609,N_19820,N_19935);
and UO_1610 (O_1610,N_19728,N_19514);
xnor UO_1611 (O_1611,N_19687,N_19775);
xor UO_1612 (O_1612,N_19870,N_19763);
nand UO_1613 (O_1613,N_19920,N_19675);
nand UO_1614 (O_1614,N_19622,N_19645);
and UO_1615 (O_1615,N_19884,N_19612);
nand UO_1616 (O_1616,N_19962,N_19978);
nand UO_1617 (O_1617,N_19579,N_19998);
and UO_1618 (O_1618,N_19923,N_19528);
or UO_1619 (O_1619,N_19870,N_19542);
and UO_1620 (O_1620,N_19758,N_19819);
or UO_1621 (O_1621,N_19707,N_19672);
nand UO_1622 (O_1622,N_19604,N_19562);
xnor UO_1623 (O_1623,N_19729,N_19845);
nor UO_1624 (O_1624,N_19820,N_19500);
nand UO_1625 (O_1625,N_19506,N_19623);
and UO_1626 (O_1626,N_19616,N_19896);
or UO_1627 (O_1627,N_19860,N_19689);
and UO_1628 (O_1628,N_19856,N_19979);
or UO_1629 (O_1629,N_19811,N_19927);
and UO_1630 (O_1630,N_19989,N_19854);
or UO_1631 (O_1631,N_19930,N_19689);
and UO_1632 (O_1632,N_19845,N_19831);
nand UO_1633 (O_1633,N_19646,N_19692);
xnor UO_1634 (O_1634,N_19831,N_19808);
nand UO_1635 (O_1635,N_19529,N_19745);
and UO_1636 (O_1636,N_19896,N_19538);
xor UO_1637 (O_1637,N_19741,N_19712);
nand UO_1638 (O_1638,N_19633,N_19529);
or UO_1639 (O_1639,N_19922,N_19854);
xnor UO_1640 (O_1640,N_19615,N_19944);
and UO_1641 (O_1641,N_19596,N_19505);
and UO_1642 (O_1642,N_19832,N_19916);
xor UO_1643 (O_1643,N_19766,N_19800);
nor UO_1644 (O_1644,N_19667,N_19886);
or UO_1645 (O_1645,N_19808,N_19883);
or UO_1646 (O_1646,N_19829,N_19744);
and UO_1647 (O_1647,N_19587,N_19654);
nor UO_1648 (O_1648,N_19527,N_19637);
nor UO_1649 (O_1649,N_19918,N_19860);
xor UO_1650 (O_1650,N_19996,N_19825);
or UO_1651 (O_1651,N_19586,N_19764);
and UO_1652 (O_1652,N_19617,N_19754);
nand UO_1653 (O_1653,N_19511,N_19927);
xor UO_1654 (O_1654,N_19833,N_19659);
nor UO_1655 (O_1655,N_19790,N_19791);
nand UO_1656 (O_1656,N_19894,N_19625);
or UO_1657 (O_1657,N_19746,N_19931);
xor UO_1658 (O_1658,N_19911,N_19978);
and UO_1659 (O_1659,N_19980,N_19815);
or UO_1660 (O_1660,N_19807,N_19589);
nand UO_1661 (O_1661,N_19757,N_19698);
nand UO_1662 (O_1662,N_19662,N_19526);
nand UO_1663 (O_1663,N_19569,N_19833);
xnor UO_1664 (O_1664,N_19519,N_19769);
or UO_1665 (O_1665,N_19566,N_19794);
or UO_1666 (O_1666,N_19901,N_19621);
nor UO_1667 (O_1667,N_19508,N_19755);
nor UO_1668 (O_1668,N_19520,N_19575);
or UO_1669 (O_1669,N_19512,N_19950);
nand UO_1670 (O_1670,N_19658,N_19833);
or UO_1671 (O_1671,N_19982,N_19847);
or UO_1672 (O_1672,N_19848,N_19949);
nor UO_1673 (O_1673,N_19691,N_19630);
or UO_1674 (O_1674,N_19871,N_19895);
and UO_1675 (O_1675,N_19596,N_19745);
nor UO_1676 (O_1676,N_19734,N_19548);
and UO_1677 (O_1677,N_19833,N_19685);
nor UO_1678 (O_1678,N_19956,N_19986);
nor UO_1679 (O_1679,N_19569,N_19574);
xnor UO_1680 (O_1680,N_19549,N_19972);
xor UO_1681 (O_1681,N_19823,N_19687);
nor UO_1682 (O_1682,N_19637,N_19504);
nand UO_1683 (O_1683,N_19501,N_19839);
xor UO_1684 (O_1684,N_19998,N_19628);
and UO_1685 (O_1685,N_19995,N_19725);
or UO_1686 (O_1686,N_19637,N_19535);
and UO_1687 (O_1687,N_19581,N_19537);
xnor UO_1688 (O_1688,N_19857,N_19586);
xnor UO_1689 (O_1689,N_19629,N_19887);
xnor UO_1690 (O_1690,N_19565,N_19543);
nand UO_1691 (O_1691,N_19806,N_19861);
nand UO_1692 (O_1692,N_19872,N_19728);
and UO_1693 (O_1693,N_19593,N_19872);
and UO_1694 (O_1694,N_19717,N_19932);
and UO_1695 (O_1695,N_19587,N_19753);
or UO_1696 (O_1696,N_19700,N_19757);
xnor UO_1697 (O_1697,N_19515,N_19518);
or UO_1698 (O_1698,N_19917,N_19788);
and UO_1699 (O_1699,N_19841,N_19865);
xor UO_1700 (O_1700,N_19709,N_19762);
nor UO_1701 (O_1701,N_19644,N_19599);
or UO_1702 (O_1702,N_19574,N_19662);
or UO_1703 (O_1703,N_19693,N_19976);
and UO_1704 (O_1704,N_19867,N_19821);
and UO_1705 (O_1705,N_19678,N_19920);
and UO_1706 (O_1706,N_19627,N_19825);
or UO_1707 (O_1707,N_19961,N_19545);
nand UO_1708 (O_1708,N_19882,N_19621);
nand UO_1709 (O_1709,N_19942,N_19945);
nor UO_1710 (O_1710,N_19854,N_19616);
or UO_1711 (O_1711,N_19771,N_19886);
xor UO_1712 (O_1712,N_19659,N_19751);
nor UO_1713 (O_1713,N_19896,N_19919);
nand UO_1714 (O_1714,N_19575,N_19860);
nor UO_1715 (O_1715,N_19875,N_19976);
xor UO_1716 (O_1716,N_19874,N_19703);
xor UO_1717 (O_1717,N_19828,N_19653);
nor UO_1718 (O_1718,N_19801,N_19851);
xnor UO_1719 (O_1719,N_19535,N_19725);
nor UO_1720 (O_1720,N_19607,N_19927);
and UO_1721 (O_1721,N_19822,N_19843);
nor UO_1722 (O_1722,N_19553,N_19662);
xnor UO_1723 (O_1723,N_19764,N_19648);
xor UO_1724 (O_1724,N_19623,N_19515);
xnor UO_1725 (O_1725,N_19573,N_19667);
nor UO_1726 (O_1726,N_19974,N_19730);
or UO_1727 (O_1727,N_19795,N_19959);
nor UO_1728 (O_1728,N_19528,N_19513);
nor UO_1729 (O_1729,N_19542,N_19818);
and UO_1730 (O_1730,N_19815,N_19752);
and UO_1731 (O_1731,N_19811,N_19583);
nor UO_1732 (O_1732,N_19578,N_19825);
nor UO_1733 (O_1733,N_19749,N_19557);
xnor UO_1734 (O_1734,N_19850,N_19785);
xor UO_1735 (O_1735,N_19656,N_19745);
or UO_1736 (O_1736,N_19596,N_19735);
nor UO_1737 (O_1737,N_19858,N_19636);
xor UO_1738 (O_1738,N_19729,N_19994);
xor UO_1739 (O_1739,N_19524,N_19929);
and UO_1740 (O_1740,N_19706,N_19862);
or UO_1741 (O_1741,N_19868,N_19588);
nor UO_1742 (O_1742,N_19778,N_19893);
nand UO_1743 (O_1743,N_19534,N_19527);
and UO_1744 (O_1744,N_19921,N_19702);
or UO_1745 (O_1745,N_19805,N_19716);
nor UO_1746 (O_1746,N_19598,N_19961);
nand UO_1747 (O_1747,N_19619,N_19624);
or UO_1748 (O_1748,N_19609,N_19693);
and UO_1749 (O_1749,N_19586,N_19839);
nor UO_1750 (O_1750,N_19854,N_19798);
or UO_1751 (O_1751,N_19994,N_19888);
xor UO_1752 (O_1752,N_19785,N_19630);
nor UO_1753 (O_1753,N_19650,N_19711);
nor UO_1754 (O_1754,N_19743,N_19791);
and UO_1755 (O_1755,N_19868,N_19905);
or UO_1756 (O_1756,N_19862,N_19571);
or UO_1757 (O_1757,N_19735,N_19968);
xor UO_1758 (O_1758,N_19856,N_19849);
nor UO_1759 (O_1759,N_19939,N_19697);
nor UO_1760 (O_1760,N_19602,N_19913);
xor UO_1761 (O_1761,N_19801,N_19904);
nor UO_1762 (O_1762,N_19768,N_19822);
nor UO_1763 (O_1763,N_19776,N_19652);
and UO_1764 (O_1764,N_19970,N_19820);
xor UO_1765 (O_1765,N_19623,N_19880);
xnor UO_1766 (O_1766,N_19635,N_19544);
nand UO_1767 (O_1767,N_19543,N_19696);
nand UO_1768 (O_1768,N_19803,N_19874);
xor UO_1769 (O_1769,N_19557,N_19876);
nor UO_1770 (O_1770,N_19668,N_19613);
nor UO_1771 (O_1771,N_19892,N_19540);
nand UO_1772 (O_1772,N_19698,N_19512);
and UO_1773 (O_1773,N_19769,N_19604);
nor UO_1774 (O_1774,N_19951,N_19869);
xor UO_1775 (O_1775,N_19967,N_19833);
nor UO_1776 (O_1776,N_19542,N_19763);
xor UO_1777 (O_1777,N_19628,N_19620);
nor UO_1778 (O_1778,N_19830,N_19614);
xor UO_1779 (O_1779,N_19801,N_19966);
xnor UO_1780 (O_1780,N_19879,N_19617);
and UO_1781 (O_1781,N_19973,N_19606);
nor UO_1782 (O_1782,N_19905,N_19965);
xnor UO_1783 (O_1783,N_19619,N_19525);
nand UO_1784 (O_1784,N_19821,N_19574);
or UO_1785 (O_1785,N_19784,N_19826);
nor UO_1786 (O_1786,N_19945,N_19570);
xor UO_1787 (O_1787,N_19869,N_19943);
and UO_1788 (O_1788,N_19681,N_19993);
and UO_1789 (O_1789,N_19817,N_19540);
xor UO_1790 (O_1790,N_19586,N_19758);
nor UO_1791 (O_1791,N_19828,N_19700);
nand UO_1792 (O_1792,N_19529,N_19678);
nor UO_1793 (O_1793,N_19949,N_19513);
xor UO_1794 (O_1794,N_19593,N_19997);
and UO_1795 (O_1795,N_19610,N_19773);
or UO_1796 (O_1796,N_19914,N_19781);
nor UO_1797 (O_1797,N_19756,N_19968);
and UO_1798 (O_1798,N_19883,N_19722);
nor UO_1799 (O_1799,N_19965,N_19795);
and UO_1800 (O_1800,N_19895,N_19853);
or UO_1801 (O_1801,N_19766,N_19967);
nor UO_1802 (O_1802,N_19634,N_19967);
nand UO_1803 (O_1803,N_19568,N_19957);
and UO_1804 (O_1804,N_19634,N_19971);
nor UO_1805 (O_1805,N_19942,N_19890);
and UO_1806 (O_1806,N_19967,N_19789);
or UO_1807 (O_1807,N_19711,N_19935);
or UO_1808 (O_1808,N_19597,N_19564);
nor UO_1809 (O_1809,N_19723,N_19989);
and UO_1810 (O_1810,N_19608,N_19790);
nand UO_1811 (O_1811,N_19604,N_19638);
xor UO_1812 (O_1812,N_19767,N_19632);
and UO_1813 (O_1813,N_19922,N_19837);
or UO_1814 (O_1814,N_19950,N_19717);
nor UO_1815 (O_1815,N_19658,N_19891);
nand UO_1816 (O_1816,N_19948,N_19992);
or UO_1817 (O_1817,N_19985,N_19579);
nor UO_1818 (O_1818,N_19603,N_19889);
or UO_1819 (O_1819,N_19712,N_19677);
or UO_1820 (O_1820,N_19820,N_19720);
or UO_1821 (O_1821,N_19613,N_19807);
or UO_1822 (O_1822,N_19627,N_19980);
or UO_1823 (O_1823,N_19775,N_19895);
and UO_1824 (O_1824,N_19837,N_19834);
xnor UO_1825 (O_1825,N_19611,N_19639);
or UO_1826 (O_1826,N_19921,N_19923);
and UO_1827 (O_1827,N_19942,N_19553);
xnor UO_1828 (O_1828,N_19673,N_19800);
xnor UO_1829 (O_1829,N_19608,N_19900);
xor UO_1830 (O_1830,N_19819,N_19782);
or UO_1831 (O_1831,N_19514,N_19625);
nand UO_1832 (O_1832,N_19924,N_19541);
nor UO_1833 (O_1833,N_19904,N_19949);
and UO_1834 (O_1834,N_19715,N_19843);
nor UO_1835 (O_1835,N_19801,N_19773);
and UO_1836 (O_1836,N_19837,N_19555);
nand UO_1837 (O_1837,N_19719,N_19612);
nor UO_1838 (O_1838,N_19555,N_19687);
or UO_1839 (O_1839,N_19983,N_19613);
and UO_1840 (O_1840,N_19807,N_19512);
and UO_1841 (O_1841,N_19511,N_19757);
or UO_1842 (O_1842,N_19544,N_19783);
or UO_1843 (O_1843,N_19524,N_19661);
or UO_1844 (O_1844,N_19560,N_19536);
nand UO_1845 (O_1845,N_19938,N_19968);
xnor UO_1846 (O_1846,N_19805,N_19685);
nand UO_1847 (O_1847,N_19565,N_19621);
xnor UO_1848 (O_1848,N_19698,N_19753);
and UO_1849 (O_1849,N_19657,N_19521);
or UO_1850 (O_1850,N_19921,N_19944);
and UO_1851 (O_1851,N_19918,N_19823);
xnor UO_1852 (O_1852,N_19504,N_19660);
or UO_1853 (O_1853,N_19673,N_19668);
xnor UO_1854 (O_1854,N_19519,N_19989);
nor UO_1855 (O_1855,N_19843,N_19586);
or UO_1856 (O_1856,N_19735,N_19601);
or UO_1857 (O_1857,N_19582,N_19846);
nor UO_1858 (O_1858,N_19816,N_19636);
or UO_1859 (O_1859,N_19899,N_19901);
and UO_1860 (O_1860,N_19800,N_19934);
and UO_1861 (O_1861,N_19991,N_19651);
nor UO_1862 (O_1862,N_19735,N_19768);
nand UO_1863 (O_1863,N_19634,N_19583);
or UO_1864 (O_1864,N_19805,N_19972);
and UO_1865 (O_1865,N_19855,N_19993);
or UO_1866 (O_1866,N_19811,N_19952);
xnor UO_1867 (O_1867,N_19736,N_19702);
nand UO_1868 (O_1868,N_19906,N_19636);
nand UO_1869 (O_1869,N_19763,N_19614);
xor UO_1870 (O_1870,N_19840,N_19891);
nor UO_1871 (O_1871,N_19717,N_19706);
nor UO_1872 (O_1872,N_19724,N_19552);
xnor UO_1873 (O_1873,N_19834,N_19636);
nand UO_1874 (O_1874,N_19764,N_19624);
nand UO_1875 (O_1875,N_19657,N_19999);
nor UO_1876 (O_1876,N_19570,N_19900);
nor UO_1877 (O_1877,N_19858,N_19746);
nor UO_1878 (O_1878,N_19974,N_19614);
and UO_1879 (O_1879,N_19640,N_19692);
or UO_1880 (O_1880,N_19517,N_19791);
nand UO_1881 (O_1881,N_19902,N_19863);
nand UO_1882 (O_1882,N_19532,N_19888);
nand UO_1883 (O_1883,N_19647,N_19877);
xnor UO_1884 (O_1884,N_19931,N_19979);
and UO_1885 (O_1885,N_19727,N_19631);
and UO_1886 (O_1886,N_19982,N_19737);
xnor UO_1887 (O_1887,N_19796,N_19652);
nand UO_1888 (O_1888,N_19656,N_19741);
and UO_1889 (O_1889,N_19991,N_19686);
and UO_1890 (O_1890,N_19812,N_19650);
and UO_1891 (O_1891,N_19933,N_19881);
xnor UO_1892 (O_1892,N_19967,N_19948);
nor UO_1893 (O_1893,N_19829,N_19855);
and UO_1894 (O_1894,N_19526,N_19699);
nand UO_1895 (O_1895,N_19634,N_19798);
and UO_1896 (O_1896,N_19772,N_19783);
nand UO_1897 (O_1897,N_19869,N_19584);
nand UO_1898 (O_1898,N_19825,N_19787);
and UO_1899 (O_1899,N_19887,N_19918);
and UO_1900 (O_1900,N_19611,N_19723);
nand UO_1901 (O_1901,N_19638,N_19744);
or UO_1902 (O_1902,N_19591,N_19971);
or UO_1903 (O_1903,N_19670,N_19986);
nor UO_1904 (O_1904,N_19542,N_19778);
or UO_1905 (O_1905,N_19745,N_19556);
nor UO_1906 (O_1906,N_19814,N_19504);
nor UO_1907 (O_1907,N_19623,N_19608);
nor UO_1908 (O_1908,N_19927,N_19706);
nand UO_1909 (O_1909,N_19900,N_19935);
xor UO_1910 (O_1910,N_19618,N_19706);
nor UO_1911 (O_1911,N_19621,N_19894);
and UO_1912 (O_1912,N_19917,N_19954);
nor UO_1913 (O_1913,N_19910,N_19705);
nand UO_1914 (O_1914,N_19710,N_19776);
xor UO_1915 (O_1915,N_19757,N_19886);
xor UO_1916 (O_1916,N_19764,N_19952);
or UO_1917 (O_1917,N_19514,N_19727);
nand UO_1918 (O_1918,N_19653,N_19763);
nand UO_1919 (O_1919,N_19747,N_19954);
xnor UO_1920 (O_1920,N_19889,N_19562);
nand UO_1921 (O_1921,N_19556,N_19713);
nand UO_1922 (O_1922,N_19795,N_19989);
nand UO_1923 (O_1923,N_19582,N_19799);
or UO_1924 (O_1924,N_19580,N_19828);
or UO_1925 (O_1925,N_19808,N_19847);
nand UO_1926 (O_1926,N_19804,N_19819);
and UO_1927 (O_1927,N_19561,N_19627);
and UO_1928 (O_1928,N_19935,N_19755);
and UO_1929 (O_1929,N_19763,N_19576);
and UO_1930 (O_1930,N_19867,N_19893);
or UO_1931 (O_1931,N_19500,N_19951);
nand UO_1932 (O_1932,N_19913,N_19591);
nor UO_1933 (O_1933,N_19913,N_19713);
and UO_1934 (O_1934,N_19864,N_19783);
and UO_1935 (O_1935,N_19796,N_19948);
xnor UO_1936 (O_1936,N_19522,N_19508);
xnor UO_1937 (O_1937,N_19522,N_19681);
xor UO_1938 (O_1938,N_19890,N_19513);
and UO_1939 (O_1939,N_19627,N_19713);
nor UO_1940 (O_1940,N_19729,N_19923);
or UO_1941 (O_1941,N_19749,N_19902);
or UO_1942 (O_1942,N_19867,N_19955);
and UO_1943 (O_1943,N_19709,N_19758);
xor UO_1944 (O_1944,N_19574,N_19708);
or UO_1945 (O_1945,N_19935,N_19882);
nor UO_1946 (O_1946,N_19591,N_19733);
nand UO_1947 (O_1947,N_19782,N_19523);
xnor UO_1948 (O_1948,N_19802,N_19895);
xor UO_1949 (O_1949,N_19963,N_19636);
or UO_1950 (O_1950,N_19500,N_19584);
nor UO_1951 (O_1951,N_19602,N_19801);
nand UO_1952 (O_1952,N_19867,N_19933);
or UO_1953 (O_1953,N_19715,N_19738);
or UO_1954 (O_1954,N_19623,N_19693);
and UO_1955 (O_1955,N_19608,N_19658);
and UO_1956 (O_1956,N_19849,N_19809);
xor UO_1957 (O_1957,N_19854,N_19955);
nor UO_1958 (O_1958,N_19935,N_19822);
or UO_1959 (O_1959,N_19858,N_19640);
nor UO_1960 (O_1960,N_19670,N_19839);
nor UO_1961 (O_1961,N_19743,N_19731);
and UO_1962 (O_1962,N_19770,N_19699);
or UO_1963 (O_1963,N_19510,N_19855);
or UO_1964 (O_1964,N_19926,N_19655);
and UO_1965 (O_1965,N_19601,N_19621);
and UO_1966 (O_1966,N_19906,N_19681);
or UO_1967 (O_1967,N_19550,N_19855);
nand UO_1968 (O_1968,N_19537,N_19667);
nand UO_1969 (O_1969,N_19989,N_19814);
and UO_1970 (O_1970,N_19553,N_19669);
nand UO_1971 (O_1971,N_19863,N_19503);
nand UO_1972 (O_1972,N_19746,N_19666);
and UO_1973 (O_1973,N_19834,N_19971);
or UO_1974 (O_1974,N_19909,N_19676);
and UO_1975 (O_1975,N_19761,N_19755);
xnor UO_1976 (O_1976,N_19946,N_19735);
and UO_1977 (O_1977,N_19754,N_19764);
nand UO_1978 (O_1978,N_19817,N_19842);
or UO_1979 (O_1979,N_19523,N_19909);
nand UO_1980 (O_1980,N_19734,N_19631);
and UO_1981 (O_1981,N_19542,N_19567);
xor UO_1982 (O_1982,N_19996,N_19594);
or UO_1983 (O_1983,N_19619,N_19696);
and UO_1984 (O_1984,N_19589,N_19693);
nand UO_1985 (O_1985,N_19992,N_19563);
nor UO_1986 (O_1986,N_19631,N_19879);
or UO_1987 (O_1987,N_19530,N_19985);
xor UO_1988 (O_1988,N_19967,N_19760);
xnor UO_1989 (O_1989,N_19825,N_19662);
nor UO_1990 (O_1990,N_19939,N_19595);
or UO_1991 (O_1991,N_19518,N_19967);
nand UO_1992 (O_1992,N_19516,N_19538);
and UO_1993 (O_1993,N_19608,N_19578);
nor UO_1994 (O_1994,N_19835,N_19791);
xor UO_1995 (O_1995,N_19701,N_19584);
nand UO_1996 (O_1996,N_19646,N_19764);
or UO_1997 (O_1997,N_19949,N_19698);
or UO_1998 (O_1998,N_19826,N_19766);
and UO_1999 (O_1999,N_19600,N_19629);
or UO_2000 (O_2000,N_19901,N_19528);
nand UO_2001 (O_2001,N_19868,N_19762);
xor UO_2002 (O_2002,N_19661,N_19571);
or UO_2003 (O_2003,N_19873,N_19753);
nor UO_2004 (O_2004,N_19644,N_19732);
and UO_2005 (O_2005,N_19974,N_19815);
nand UO_2006 (O_2006,N_19738,N_19783);
or UO_2007 (O_2007,N_19993,N_19510);
nand UO_2008 (O_2008,N_19938,N_19803);
or UO_2009 (O_2009,N_19943,N_19961);
nor UO_2010 (O_2010,N_19823,N_19628);
and UO_2011 (O_2011,N_19560,N_19715);
xor UO_2012 (O_2012,N_19596,N_19992);
and UO_2013 (O_2013,N_19607,N_19596);
xor UO_2014 (O_2014,N_19507,N_19903);
and UO_2015 (O_2015,N_19848,N_19923);
and UO_2016 (O_2016,N_19922,N_19723);
and UO_2017 (O_2017,N_19917,N_19801);
and UO_2018 (O_2018,N_19530,N_19833);
xnor UO_2019 (O_2019,N_19594,N_19546);
and UO_2020 (O_2020,N_19993,N_19683);
xnor UO_2021 (O_2021,N_19999,N_19550);
or UO_2022 (O_2022,N_19705,N_19971);
nand UO_2023 (O_2023,N_19538,N_19524);
nor UO_2024 (O_2024,N_19984,N_19936);
or UO_2025 (O_2025,N_19582,N_19741);
and UO_2026 (O_2026,N_19790,N_19769);
nor UO_2027 (O_2027,N_19881,N_19767);
xnor UO_2028 (O_2028,N_19519,N_19670);
nor UO_2029 (O_2029,N_19932,N_19714);
nor UO_2030 (O_2030,N_19687,N_19722);
or UO_2031 (O_2031,N_19791,N_19568);
and UO_2032 (O_2032,N_19716,N_19709);
nand UO_2033 (O_2033,N_19672,N_19934);
nor UO_2034 (O_2034,N_19732,N_19545);
or UO_2035 (O_2035,N_19910,N_19824);
or UO_2036 (O_2036,N_19999,N_19631);
nor UO_2037 (O_2037,N_19901,N_19861);
xor UO_2038 (O_2038,N_19852,N_19739);
and UO_2039 (O_2039,N_19609,N_19905);
and UO_2040 (O_2040,N_19544,N_19590);
and UO_2041 (O_2041,N_19618,N_19528);
or UO_2042 (O_2042,N_19756,N_19747);
xnor UO_2043 (O_2043,N_19783,N_19912);
or UO_2044 (O_2044,N_19652,N_19927);
or UO_2045 (O_2045,N_19868,N_19605);
nand UO_2046 (O_2046,N_19679,N_19706);
nand UO_2047 (O_2047,N_19511,N_19998);
nand UO_2048 (O_2048,N_19820,N_19614);
nor UO_2049 (O_2049,N_19619,N_19872);
and UO_2050 (O_2050,N_19887,N_19693);
xor UO_2051 (O_2051,N_19938,N_19788);
xor UO_2052 (O_2052,N_19514,N_19655);
nand UO_2053 (O_2053,N_19961,N_19684);
nand UO_2054 (O_2054,N_19543,N_19952);
and UO_2055 (O_2055,N_19620,N_19528);
and UO_2056 (O_2056,N_19904,N_19899);
nand UO_2057 (O_2057,N_19924,N_19546);
and UO_2058 (O_2058,N_19935,N_19752);
or UO_2059 (O_2059,N_19705,N_19702);
and UO_2060 (O_2060,N_19627,N_19548);
nor UO_2061 (O_2061,N_19732,N_19718);
nor UO_2062 (O_2062,N_19822,N_19762);
nand UO_2063 (O_2063,N_19889,N_19632);
and UO_2064 (O_2064,N_19798,N_19605);
and UO_2065 (O_2065,N_19848,N_19879);
nor UO_2066 (O_2066,N_19864,N_19612);
and UO_2067 (O_2067,N_19683,N_19672);
nor UO_2068 (O_2068,N_19665,N_19550);
nand UO_2069 (O_2069,N_19989,N_19750);
nor UO_2070 (O_2070,N_19768,N_19755);
nand UO_2071 (O_2071,N_19692,N_19572);
and UO_2072 (O_2072,N_19546,N_19868);
or UO_2073 (O_2073,N_19586,N_19513);
xnor UO_2074 (O_2074,N_19876,N_19887);
nor UO_2075 (O_2075,N_19885,N_19774);
or UO_2076 (O_2076,N_19663,N_19744);
or UO_2077 (O_2077,N_19711,N_19882);
nand UO_2078 (O_2078,N_19613,N_19718);
nand UO_2079 (O_2079,N_19809,N_19501);
or UO_2080 (O_2080,N_19959,N_19943);
nand UO_2081 (O_2081,N_19574,N_19896);
nand UO_2082 (O_2082,N_19583,N_19844);
nand UO_2083 (O_2083,N_19762,N_19979);
nor UO_2084 (O_2084,N_19742,N_19970);
xnor UO_2085 (O_2085,N_19577,N_19796);
nor UO_2086 (O_2086,N_19864,N_19891);
nor UO_2087 (O_2087,N_19502,N_19610);
nor UO_2088 (O_2088,N_19808,N_19895);
and UO_2089 (O_2089,N_19718,N_19629);
nand UO_2090 (O_2090,N_19723,N_19839);
and UO_2091 (O_2091,N_19626,N_19744);
xnor UO_2092 (O_2092,N_19947,N_19520);
and UO_2093 (O_2093,N_19685,N_19528);
xor UO_2094 (O_2094,N_19526,N_19624);
or UO_2095 (O_2095,N_19691,N_19937);
nor UO_2096 (O_2096,N_19620,N_19867);
and UO_2097 (O_2097,N_19915,N_19652);
xnor UO_2098 (O_2098,N_19738,N_19627);
nor UO_2099 (O_2099,N_19588,N_19645);
or UO_2100 (O_2100,N_19644,N_19512);
nor UO_2101 (O_2101,N_19859,N_19838);
nand UO_2102 (O_2102,N_19551,N_19710);
or UO_2103 (O_2103,N_19512,N_19592);
and UO_2104 (O_2104,N_19505,N_19744);
nor UO_2105 (O_2105,N_19926,N_19944);
nand UO_2106 (O_2106,N_19977,N_19744);
xnor UO_2107 (O_2107,N_19609,N_19606);
or UO_2108 (O_2108,N_19559,N_19952);
or UO_2109 (O_2109,N_19678,N_19715);
nor UO_2110 (O_2110,N_19721,N_19828);
and UO_2111 (O_2111,N_19957,N_19973);
or UO_2112 (O_2112,N_19585,N_19798);
and UO_2113 (O_2113,N_19954,N_19527);
nand UO_2114 (O_2114,N_19718,N_19685);
and UO_2115 (O_2115,N_19799,N_19583);
nand UO_2116 (O_2116,N_19833,N_19939);
and UO_2117 (O_2117,N_19696,N_19837);
nand UO_2118 (O_2118,N_19719,N_19883);
or UO_2119 (O_2119,N_19895,N_19700);
and UO_2120 (O_2120,N_19850,N_19623);
xnor UO_2121 (O_2121,N_19944,N_19770);
nand UO_2122 (O_2122,N_19996,N_19687);
nand UO_2123 (O_2123,N_19649,N_19751);
nor UO_2124 (O_2124,N_19959,N_19911);
nand UO_2125 (O_2125,N_19632,N_19946);
xor UO_2126 (O_2126,N_19850,N_19515);
nand UO_2127 (O_2127,N_19865,N_19508);
nor UO_2128 (O_2128,N_19891,N_19919);
xnor UO_2129 (O_2129,N_19830,N_19766);
or UO_2130 (O_2130,N_19758,N_19566);
or UO_2131 (O_2131,N_19550,N_19581);
or UO_2132 (O_2132,N_19889,N_19803);
and UO_2133 (O_2133,N_19665,N_19990);
nor UO_2134 (O_2134,N_19673,N_19918);
xor UO_2135 (O_2135,N_19835,N_19979);
and UO_2136 (O_2136,N_19785,N_19642);
nand UO_2137 (O_2137,N_19548,N_19942);
or UO_2138 (O_2138,N_19641,N_19717);
nor UO_2139 (O_2139,N_19980,N_19875);
and UO_2140 (O_2140,N_19643,N_19533);
nor UO_2141 (O_2141,N_19572,N_19729);
and UO_2142 (O_2142,N_19785,N_19714);
or UO_2143 (O_2143,N_19578,N_19728);
nor UO_2144 (O_2144,N_19784,N_19876);
nor UO_2145 (O_2145,N_19884,N_19822);
and UO_2146 (O_2146,N_19982,N_19549);
nor UO_2147 (O_2147,N_19955,N_19905);
nand UO_2148 (O_2148,N_19565,N_19528);
xnor UO_2149 (O_2149,N_19881,N_19838);
or UO_2150 (O_2150,N_19918,N_19744);
xnor UO_2151 (O_2151,N_19709,N_19647);
nand UO_2152 (O_2152,N_19676,N_19766);
nor UO_2153 (O_2153,N_19650,N_19854);
and UO_2154 (O_2154,N_19619,N_19707);
nor UO_2155 (O_2155,N_19866,N_19660);
or UO_2156 (O_2156,N_19903,N_19694);
nor UO_2157 (O_2157,N_19862,N_19912);
xor UO_2158 (O_2158,N_19628,N_19588);
or UO_2159 (O_2159,N_19875,N_19892);
nand UO_2160 (O_2160,N_19598,N_19975);
nor UO_2161 (O_2161,N_19565,N_19554);
nor UO_2162 (O_2162,N_19558,N_19686);
or UO_2163 (O_2163,N_19575,N_19576);
or UO_2164 (O_2164,N_19955,N_19546);
or UO_2165 (O_2165,N_19990,N_19967);
or UO_2166 (O_2166,N_19828,N_19641);
nand UO_2167 (O_2167,N_19833,N_19793);
nand UO_2168 (O_2168,N_19530,N_19710);
nand UO_2169 (O_2169,N_19938,N_19777);
xor UO_2170 (O_2170,N_19580,N_19644);
nand UO_2171 (O_2171,N_19607,N_19786);
nand UO_2172 (O_2172,N_19992,N_19773);
or UO_2173 (O_2173,N_19775,N_19753);
nor UO_2174 (O_2174,N_19512,N_19588);
and UO_2175 (O_2175,N_19644,N_19975);
xor UO_2176 (O_2176,N_19566,N_19698);
nand UO_2177 (O_2177,N_19725,N_19611);
or UO_2178 (O_2178,N_19871,N_19766);
xor UO_2179 (O_2179,N_19848,N_19681);
nand UO_2180 (O_2180,N_19926,N_19527);
nand UO_2181 (O_2181,N_19600,N_19830);
and UO_2182 (O_2182,N_19519,N_19613);
or UO_2183 (O_2183,N_19604,N_19629);
or UO_2184 (O_2184,N_19873,N_19805);
xnor UO_2185 (O_2185,N_19748,N_19606);
xnor UO_2186 (O_2186,N_19783,N_19550);
and UO_2187 (O_2187,N_19632,N_19807);
and UO_2188 (O_2188,N_19558,N_19520);
xor UO_2189 (O_2189,N_19789,N_19892);
xor UO_2190 (O_2190,N_19890,N_19659);
xnor UO_2191 (O_2191,N_19912,N_19686);
and UO_2192 (O_2192,N_19927,N_19777);
xor UO_2193 (O_2193,N_19520,N_19659);
nand UO_2194 (O_2194,N_19666,N_19600);
and UO_2195 (O_2195,N_19802,N_19665);
and UO_2196 (O_2196,N_19638,N_19826);
nor UO_2197 (O_2197,N_19791,N_19894);
or UO_2198 (O_2198,N_19914,N_19787);
nor UO_2199 (O_2199,N_19841,N_19861);
nor UO_2200 (O_2200,N_19975,N_19707);
xor UO_2201 (O_2201,N_19781,N_19550);
xnor UO_2202 (O_2202,N_19988,N_19952);
or UO_2203 (O_2203,N_19798,N_19956);
or UO_2204 (O_2204,N_19745,N_19693);
nor UO_2205 (O_2205,N_19748,N_19569);
and UO_2206 (O_2206,N_19607,N_19569);
xor UO_2207 (O_2207,N_19755,N_19983);
nor UO_2208 (O_2208,N_19806,N_19670);
nand UO_2209 (O_2209,N_19810,N_19533);
nor UO_2210 (O_2210,N_19825,N_19635);
nand UO_2211 (O_2211,N_19740,N_19556);
nor UO_2212 (O_2212,N_19952,N_19643);
nand UO_2213 (O_2213,N_19589,N_19981);
or UO_2214 (O_2214,N_19912,N_19611);
or UO_2215 (O_2215,N_19656,N_19972);
nand UO_2216 (O_2216,N_19614,N_19769);
nor UO_2217 (O_2217,N_19813,N_19794);
nand UO_2218 (O_2218,N_19604,N_19581);
nand UO_2219 (O_2219,N_19686,N_19505);
nor UO_2220 (O_2220,N_19986,N_19928);
nor UO_2221 (O_2221,N_19870,N_19835);
or UO_2222 (O_2222,N_19700,N_19851);
nor UO_2223 (O_2223,N_19848,N_19768);
xor UO_2224 (O_2224,N_19513,N_19816);
nand UO_2225 (O_2225,N_19699,N_19777);
nand UO_2226 (O_2226,N_19583,N_19990);
xnor UO_2227 (O_2227,N_19624,N_19933);
and UO_2228 (O_2228,N_19807,N_19713);
nor UO_2229 (O_2229,N_19773,N_19885);
or UO_2230 (O_2230,N_19611,N_19899);
nand UO_2231 (O_2231,N_19546,N_19891);
or UO_2232 (O_2232,N_19708,N_19972);
and UO_2233 (O_2233,N_19594,N_19781);
xnor UO_2234 (O_2234,N_19628,N_19949);
and UO_2235 (O_2235,N_19924,N_19535);
or UO_2236 (O_2236,N_19527,N_19778);
xor UO_2237 (O_2237,N_19627,N_19708);
xor UO_2238 (O_2238,N_19986,N_19510);
nor UO_2239 (O_2239,N_19858,N_19924);
nand UO_2240 (O_2240,N_19569,N_19890);
and UO_2241 (O_2241,N_19683,N_19809);
nor UO_2242 (O_2242,N_19728,N_19824);
nand UO_2243 (O_2243,N_19794,N_19775);
nand UO_2244 (O_2244,N_19877,N_19876);
nor UO_2245 (O_2245,N_19902,N_19628);
xnor UO_2246 (O_2246,N_19803,N_19932);
or UO_2247 (O_2247,N_19841,N_19591);
and UO_2248 (O_2248,N_19596,N_19697);
nand UO_2249 (O_2249,N_19961,N_19702);
and UO_2250 (O_2250,N_19585,N_19972);
nand UO_2251 (O_2251,N_19796,N_19537);
and UO_2252 (O_2252,N_19860,N_19694);
nor UO_2253 (O_2253,N_19848,N_19770);
nand UO_2254 (O_2254,N_19922,N_19941);
or UO_2255 (O_2255,N_19911,N_19833);
nand UO_2256 (O_2256,N_19531,N_19928);
and UO_2257 (O_2257,N_19951,N_19699);
xnor UO_2258 (O_2258,N_19883,N_19683);
or UO_2259 (O_2259,N_19977,N_19950);
nand UO_2260 (O_2260,N_19515,N_19788);
and UO_2261 (O_2261,N_19798,N_19990);
xnor UO_2262 (O_2262,N_19891,N_19587);
and UO_2263 (O_2263,N_19749,N_19917);
nor UO_2264 (O_2264,N_19881,N_19898);
nand UO_2265 (O_2265,N_19645,N_19924);
nand UO_2266 (O_2266,N_19549,N_19574);
or UO_2267 (O_2267,N_19982,N_19668);
nor UO_2268 (O_2268,N_19858,N_19771);
and UO_2269 (O_2269,N_19608,N_19525);
and UO_2270 (O_2270,N_19798,N_19925);
or UO_2271 (O_2271,N_19753,N_19694);
or UO_2272 (O_2272,N_19678,N_19998);
nand UO_2273 (O_2273,N_19503,N_19932);
and UO_2274 (O_2274,N_19602,N_19687);
xnor UO_2275 (O_2275,N_19543,N_19663);
xor UO_2276 (O_2276,N_19640,N_19584);
nand UO_2277 (O_2277,N_19719,N_19716);
and UO_2278 (O_2278,N_19650,N_19661);
nor UO_2279 (O_2279,N_19791,N_19775);
or UO_2280 (O_2280,N_19703,N_19637);
or UO_2281 (O_2281,N_19843,N_19971);
nor UO_2282 (O_2282,N_19583,N_19687);
and UO_2283 (O_2283,N_19827,N_19527);
nand UO_2284 (O_2284,N_19693,N_19788);
xnor UO_2285 (O_2285,N_19565,N_19792);
nand UO_2286 (O_2286,N_19964,N_19946);
or UO_2287 (O_2287,N_19611,N_19928);
nand UO_2288 (O_2288,N_19800,N_19840);
or UO_2289 (O_2289,N_19556,N_19814);
nor UO_2290 (O_2290,N_19515,N_19924);
nand UO_2291 (O_2291,N_19568,N_19922);
xnor UO_2292 (O_2292,N_19796,N_19566);
xor UO_2293 (O_2293,N_19506,N_19830);
nand UO_2294 (O_2294,N_19923,N_19551);
nand UO_2295 (O_2295,N_19567,N_19721);
xor UO_2296 (O_2296,N_19784,N_19958);
or UO_2297 (O_2297,N_19955,N_19617);
xor UO_2298 (O_2298,N_19572,N_19723);
and UO_2299 (O_2299,N_19776,N_19730);
and UO_2300 (O_2300,N_19584,N_19970);
or UO_2301 (O_2301,N_19876,N_19978);
xnor UO_2302 (O_2302,N_19912,N_19595);
and UO_2303 (O_2303,N_19728,N_19948);
nor UO_2304 (O_2304,N_19824,N_19664);
xnor UO_2305 (O_2305,N_19766,N_19839);
or UO_2306 (O_2306,N_19721,N_19708);
nor UO_2307 (O_2307,N_19556,N_19605);
and UO_2308 (O_2308,N_19716,N_19893);
nor UO_2309 (O_2309,N_19537,N_19828);
and UO_2310 (O_2310,N_19846,N_19764);
and UO_2311 (O_2311,N_19572,N_19734);
or UO_2312 (O_2312,N_19920,N_19628);
and UO_2313 (O_2313,N_19881,N_19892);
or UO_2314 (O_2314,N_19882,N_19947);
nor UO_2315 (O_2315,N_19708,N_19697);
nand UO_2316 (O_2316,N_19807,N_19615);
or UO_2317 (O_2317,N_19995,N_19638);
and UO_2318 (O_2318,N_19616,N_19628);
nand UO_2319 (O_2319,N_19718,N_19892);
nor UO_2320 (O_2320,N_19784,N_19731);
nand UO_2321 (O_2321,N_19826,N_19594);
nor UO_2322 (O_2322,N_19672,N_19735);
nand UO_2323 (O_2323,N_19807,N_19968);
or UO_2324 (O_2324,N_19934,N_19653);
or UO_2325 (O_2325,N_19650,N_19729);
nand UO_2326 (O_2326,N_19643,N_19697);
nor UO_2327 (O_2327,N_19874,N_19512);
or UO_2328 (O_2328,N_19775,N_19694);
xor UO_2329 (O_2329,N_19811,N_19975);
and UO_2330 (O_2330,N_19579,N_19526);
nor UO_2331 (O_2331,N_19939,N_19749);
xnor UO_2332 (O_2332,N_19650,N_19886);
xnor UO_2333 (O_2333,N_19616,N_19825);
and UO_2334 (O_2334,N_19901,N_19752);
and UO_2335 (O_2335,N_19547,N_19814);
nor UO_2336 (O_2336,N_19507,N_19510);
or UO_2337 (O_2337,N_19505,N_19896);
nor UO_2338 (O_2338,N_19519,N_19637);
nand UO_2339 (O_2339,N_19590,N_19527);
xnor UO_2340 (O_2340,N_19767,N_19706);
nand UO_2341 (O_2341,N_19936,N_19764);
and UO_2342 (O_2342,N_19699,N_19525);
nor UO_2343 (O_2343,N_19927,N_19802);
nor UO_2344 (O_2344,N_19532,N_19786);
nand UO_2345 (O_2345,N_19598,N_19786);
and UO_2346 (O_2346,N_19944,N_19952);
xor UO_2347 (O_2347,N_19672,N_19973);
nor UO_2348 (O_2348,N_19781,N_19624);
and UO_2349 (O_2349,N_19775,N_19994);
nand UO_2350 (O_2350,N_19713,N_19555);
nor UO_2351 (O_2351,N_19647,N_19750);
xnor UO_2352 (O_2352,N_19672,N_19758);
nor UO_2353 (O_2353,N_19710,N_19944);
xnor UO_2354 (O_2354,N_19806,N_19856);
or UO_2355 (O_2355,N_19625,N_19714);
and UO_2356 (O_2356,N_19800,N_19894);
nand UO_2357 (O_2357,N_19925,N_19940);
and UO_2358 (O_2358,N_19982,N_19700);
and UO_2359 (O_2359,N_19819,N_19977);
xnor UO_2360 (O_2360,N_19744,N_19745);
or UO_2361 (O_2361,N_19545,N_19885);
xor UO_2362 (O_2362,N_19900,N_19987);
nor UO_2363 (O_2363,N_19501,N_19823);
nand UO_2364 (O_2364,N_19622,N_19770);
nor UO_2365 (O_2365,N_19831,N_19677);
and UO_2366 (O_2366,N_19739,N_19711);
nand UO_2367 (O_2367,N_19559,N_19761);
and UO_2368 (O_2368,N_19795,N_19675);
or UO_2369 (O_2369,N_19925,N_19639);
and UO_2370 (O_2370,N_19528,N_19639);
nand UO_2371 (O_2371,N_19944,N_19586);
or UO_2372 (O_2372,N_19761,N_19629);
nor UO_2373 (O_2373,N_19849,N_19740);
or UO_2374 (O_2374,N_19895,N_19839);
xnor UO_2375 (O_2375,N_19746,N_19919);
nor UO_2376 (O_2376,N_19521,N_19778);
and UO_2377 (O_2377,N_19674,N_19998);
nor UO_2378 (O_2378,N_19518,N_19900);
nand UO_2379 (O_2379,N_19774,N_19728);
and UO_2380 (O_2380,N_19940,N_19786);
or UO_2381 (O_2381,N_19825,N_19746);
nor UO_2382 (O_2382,N_19867,N_19546);
nor UO_2383 (O_2383,N_19541,N_19505);
nand UO_2384 (O_2384,N_19652,N_19549);
nor UO_2385 (O_2385,N_19833,N_19853);
and UO_2386 (O_2386,N_19723,N_19810);
or UO_2387 (O_2387,N_19545,N_19755);
or UO_2388 (O_2388,N_19619,N_19863);
or UO_2389 (O_2389,N_19590,N_19692);
nor UO_2390 (O_2390,N_19826,N_19748);
nand UO_2391 (O_2391,N_19676,N_19758);
nand UO_2392 (O_2392,N_19722,N_19812);
or UO_2393 (O_2393,N_19533,N_19718);
nor UO_2394 (O_2394,N_19641,N_19618);
or UO_2395 (O_2395,N_19515,N_19532);
nor UO_2396 (O_2396,N_19957,N_19955);
xnor UO_2397 (O_2397,N_19851,N_19736);
xor UO_2398 (O_2398,N_19875,N_19828);
or UO_2399 (O_2399,N_19703,N_19938);
nand UO_2400 (O_2400,N_19720,N_19792);
and UO_2401 (O_2401,N_19677,N_19679);
xnor UO_2402 (O_2402,N_19699,N_19713);
nor UO_2403 (O_2403,N_19812,N_19922);
nor UO_2404 (O_2404,N_19542,N_19638);
xnor UO_2405 (O_2405,N_19510,N_19816);
nand UO_2406 (O_2406,N_19968,N_19632);
nand UO_2407 (O_2407,N_19507,N_19572);
xor UO_2408 (O_2408,N_19644,N_19726);
or UO_2409 (O_2409,N_19877,N_19868);
and UO_2410 (O_2410,N_19503,N_19968);
xnor UO_2411 (O_2411,N_19868,N_19977);
and UO_2412 (O_2412,N_19988,N_19566);
or UO_2413 (O_2413,N_19572,N_19718);
nor UO_2414 (O_2414,N_19542,N_19653);
nand UO_2415 (O_2415,N_19859,N_19742);
xnor UO_2416 (O_2416,N_19951,N_19893);
xnor UO_2417 (O_2417,N_19545,N_19537);
xnor UO_2418 (O_2418,N_19672,N_19639);
xor UO_2419 (O_2419,N_19906,N_19528);
nor UO_2420 (O_2420,N_19862,N_19587);
and UO_2421 (O_2421,N_19687,N_19697);
and UO_2422 (O_2422,N_19741,N_19898);
and UO_2423 (O_2423,N_19600,N_19847);
nor UO_2424 (O_2424,N_19982,N_19814);
nor UO_2425 (O_2425,N_19582,N_19767);
and UO_2426 (O_2426,N_19506,N_19612);
xnor UO_2427 (O_2427,N_19632,N_19703);
nor UO_2428 (O_2428,N_19992,N_19831);
nand UO_2429 (O_2429,N_19661,N_19550);
and UO_2430 (O_2430,N_19915,N_19881);
and UO_2431 (O_2431,N_19887,N_19690);
nand UO_2432 (O_2432,N_19718,N_19515);
and UO_2433 (O_2433,N_19798,N_19985);
nand UO_2434 (O_2434,N_19729,N_19951);
nand UO_2435 (O_2435,N_19585,N_19904);
xor UO_2436 (O_2436,N_19980,N_19852);
xnor UO_2437 (O_2437,N_19693,N_19922);
nor UO_2438 (O_2438,N_19844,N_19752);
and UO_2439 (O_2439,N_19516,N_19617);
nor UO_2440 (O_2440,N_19561,N_19628);
xor UO_2441 (O_2441,N_19593,N_19678);
nor UO_2442 (O_2442,N_19920,N_19719);
nor UO_2443 (O_2443,N_19883,N_19558);
and UO_2444 (O_2444,N_19836,N_19848);
nor UO_2445 (O_2445,N_19937,N_19982);
nand UO_2446 (O_2446,N_19948,N_19979);
nor UO_2447 (O_2447,N_19562,N_19818);
nand UO_2448 (O_2448,N_19873,N_19572);
nand UO_2449 (O_2449,N_19500,N_19892);
xor UO_2450 (O_2450,N_19687,N_19595);
xnor UO_2451 (O_2451,N_19919,N_19857);
and UO_2452 (O_2452,N_19776,N_19951);
and UO_2453 (O_2453,N_19562,N_19596);
xnor UO_2454 (O_2454,N_19960,N_19984);
nor UO_2455 (O_2455,N_19529,N_19540);
nand UO_2456 (O_2456,N_19693,N_19603);
or UO_2457 (O_2457,N_19854,N_19561);
or UO_2458 (O_2458,N_19836,N_19888);
and UO_2459 (O_2459,N_19797,N_19529);
xnor UO_2460 (O_2460,N_19689,N_19587);
xor UO_2461 (O_2461,N_19556,N_19613);
nor UO_2462 (O_2462,N_19801,N_19990);
nand UO_2463 (O_2463,N_19844,N_19671);
nand UO_2464 (O_2464,N_19993,N_19963);
or UO_2465 (O_2465,N_19607,N_19741);
nor UO_2466 (O_2466,N_19823,N_19795);
or UO_2467 (O_2467,N_19804,N_19597);
xor UO_2468 (O_2468,N_19605,N_19711);
xnor UO_2469 (O_2469,N_19595,N_19843);
nor UO_2470 (O_2470,N_19603,N_19929);
and UO_2471 (O_2471,N_19767,N_19988);
and UO_2472 (O_2472,N_19673,N_19551);
nand UO_2473 (O_2473,N_19642,N_19879);
nand UO_2474 (O_2474,N_19906,N_19837);
nand UO_2475 (O_2475,N_19556,N_19618);
and UO_2476 (O_2476,N_19821,N_19960);
xnor UO_2477 (O_2477,N_19815,N_19510);
nor UO_2478 (O_2478,N_19938,N_19515);
nor UO_2479 (O_2479,N_19568,N_19570);
nand UO_2480 (O_2480,N_19836,N_19521);
and UO_2481 (O_2481,N_19947,N_19908);
or UO_2482 (O_2482,N_19738,N_19600);
nor UO_2483 (O_2483,N_19959,N_19574);
or UO_2484 (O_2484,N_19709,N_19721);
or UO_2485 (O_2485,N_19603,N_19670);
nor UO_2486 (O_2486,N_19529,N_19942);
xor UO_2487 (O_2487,N_19818,N_19628);
nor UO_2488 (O_2488,N_19679,N_19994);
xnor UO_2489 (O_2489,N_19829,N_19596);
nor UO_2490 (O_2490,N_19533,N_19730);
xnor UO_2491 (O_2491,N_19636,N_19729);
nand UO_2492 (O_2492,N_19825,N_19733);
and UO_2493 (O_2493,N_19619,N_19929);
xor UO_2494 (O_2494,N_19638,N_19764);
or UO_2495 (O_2495,N_19877,N_19581);
nand UO_2496 (O_2496,N_19732,N_19947);
nor UO_2497 (O_2497,N_19880,N_19649);
or UO_2498 (O_2498,N_19731,N_19901);
or UO_2499 (O_2499,N_19584,N_19806);
endmodule