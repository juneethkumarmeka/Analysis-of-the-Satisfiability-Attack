module basic_1000_10000_1500_50_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_802,In_397);
and U1 (N_1,In_708,In_516);
and U2 (N_2,In_995,In_206);
nor U3 (N_3,In_421,In_104);
nor U4 (N_4,In_161,In_909);
xor U5 (N_5,In_902,In_150);
and U6 (N_6,In_843,In_575);
and U7 (N_7,In_712,In_438);
and U8 (N_8,In_619,In_588);
or U9 (N_9,In_638,In_68);
and U10 (N_10,In_842,In_817);
nor U11 (N_11,In_243,In_634);
nand U12 (N_12,In_128,In_30);
nor U13 (N_13,In_444,In_349);
nor U14 (N_14,In_747,In_761);
xnor U15 (N_15,In_798,In_484);
xnor U16 (N_16,In_207,In_671);
or U17 (N_17,In_137,In_94);
nand U18 (N_18,In_470,In_83);
nor U19 (N_19,In_544,In_821);
xnor U20 (N_20,In_403,In_317);
and U21 (N_21,In_606,In_256);
nor U22 (N_22,In_139,In_687);
and U23 (N_23,In_229,In_209);
or U24 (N_24,In_330,In_432);
nand U25 (N_25,In_290,In_399);
and U26 (N_26,In_368,In_551);
nor U27 (N_27,In_834,In_13);
nand U28 (N_28,In_78,In_953);
or U29 (N_29,In_491,In_408);
or U30 (N_30,In_333,In_98);
xnor U31 (N_31,In_298,In_54);
and U32 (N_32,In_149,In_210);
nor U33 (N_33,In_646,In_85);
and U34 (N_34,In_156,In_1);
nor U35 (N_35,In_503,In_932);
xnor U36 (N_36,In_598,In_748);
xor U37 (N_37,In_215,In_966);
and U38 (N_38,In_433,In_88);
or U39 (N_39,In_65,In_682);
nor U40 (N_40,In_859,In_372);
nand U41 (N_41,In_416,In_93);
xnor U42 (N_42,In_487,In_246);
and U43 (N_43,In_986,In_188);
nor U44 (N_44,In_311,In_732);
and U45 (N_45,In_160,In_570);
nor U46 (N_46,In_861,In_445);
and U47 (N_47,In_291,In_528);
and U48 (N_48,In_559,In_144);
nor U49 (N_49,In_522,In_205);
xor U50 (N_50,In_504,In_300);
xnor U51 (N_51,In_576,In_9);
nor U52 (N_52,In_459,In_364);
xor U53 (N_53,In_868,In_158);
xnor U54 (N_54,In_879,In_579);
nand U55 (N_55,In_546,In_976);
nor U56 (N_56,In_766,In_120);
or U57 (N_57,In_335,In_635);
or U58 (N_58,In_531,In_412);
and U59 (N_59,In_686,In_954);
nor U60 (N_60,In_739,In_552);
nand U61 (N_61,In_299,In_911);
or U62 (N_62,In_376,In_782);
and U63 (N_63,In_788,In_6);
nor U64 (N_64,In_829,In_18);
or U65 (N_65,In_770,In_3);
nand U66 (N_66,In_910,In_948);
nand U67 (N_67,In_200,In_230);
nand U68 (N_68,In_138,In_266);
nand U69 (N_69,In_702,In_988);
and U70 (N_70,In_167,In_39);
xor U71 (N_71,In_680,In_42);
or U72 (N_72,In_107,In_480);
nor U73 (N_73,In_250,In_591);
and U74 (N_74,In_697,In_382);
and U75 (N_75,In_675,In_74);
nand U76 (N_76,In_142,In_305);
xnor U77 (N_77,In_58,In_858);
and U78 (N_78,In_924,In_771);
and U79 (N_79,In_884,In_287);
nand U80 (N_80,In_14,In_886);
xnor U81 (N_81,In_939,In_975);
or U82 (N_82,In_991,In_707);
xor U83 (N_83,In_791,In_961);
xnor U84 (N_84,In_37,In_688);
or U85 (N_85,In_235,In_239);
nand U86 (N_86,In_768,In_50);
or U87 (N_87,In_944,In_965);
nand U88 (N_88,In_226,In_353);
and U89 (N_89,In_454,In_324);
nand U90 (N_90,In_222,In_783);
xnor U91 (N_91,In_340,In_560);
or U92 (N_92,In_611,In_900);
nand U93 (N_93,In_295,In_224);
nor U94 (N_94,In_34,In_864);
nand U95 (N_95,In_694,In_862);
or U96 (N_96,In_386,In_418);
nand U97 (N_97,In_187,In_826);
or U98 (N_98,In_375,In_539);
xnor U99 (N_99,In_153,In_390);
and U100 (N_100,In_781,In_987);
nand U101 (N_101,In_269,In_586);
nand U102 (N_102,In_283,In_973);
or U103 (N_103,In_587,In_679);
xnor U104 (N_104,In_323,In_322);
xnor U105 (N_105,In_562,In_247);
nor U106 (N_106,In_971,In_468);
xnor U107 (N_107,In_609,In_213);
nor U108 (N_108,In_492,In_925);
nand U109 (N_109,In_281,In_564);
or U110 (N_110,In_148,In_84);
and U111 (N_111,In_760,In_392);
nand U112 (N_112,In_106,In_721);
nor U113 (N_113,In_898,In_354);
nor U114 (N_114,In_286,In_846);
or U115 (N_115,In_371,In_453);
or U116 (N_116,In_92,In_267);
nand U117 (N_117,In_271,In_97);
nor U118 (N_118,In_379,In_66);
or U119 (N_119,In_102,In_828);
or U120 (N_120,In_912,In_596);
nand U121 (N_121,In_437,In_532);
xnor U122 (N_122,In_268,In_279);
or U123 (N_123,In_75,In_358);
xnor U124 (N_124,In_57,In_530);
xor U125 (N_125,In_240,In_296);
xor U126 (N_126,In_729,In_652);
and U127 (N_127,In_162,In_461);
or U128 (N_128,In_977,In_822);
and U129 (N_129,In_872,In_816);
xor U130 (N_130,In_832,In_719);
nor U131 (N_131,In_601,In_630);
nor U132 (N_132,In_310,In_409);
nand U133 (N_133,In_417,In_327);
xnor U134 (N_134,In_775,In_893);
nand U135 (N_135,In_677,In_391);
xor U136 (N_136,In_543,In_815);
and U137 (N_137,In_952,In_590);
nor U138 (N_138,In_151,In_881);
and U139 (N_139,In_664,In_380);
nand U140 (N_140,In_969,In_479);
nand U141 (N_141,In_608,In_238);
nand U142 (N_142,In_593,In_644);
nand U143 (N_143,In_398,In_607);
nor U144 (N_144,In_850,In_177);
xor U145 (N_145,In_393,In_508);
nand U146 (N_146,In_101,In_655);
or U147 (N_147,In_347,In_293);
nor U148 (N_148,In_981,In_61);
or U149 (N_149,In_550,In_494);
nand U150 (N_150,In_254,In_159);
nand U151 (N_151,In_571,In_110);
and U152 (N_152,In_517,In_204);
xnor U153 (N_153,In_157,In_521);
nor U154 (N_154,In_15,In_183);
xnor U155 (N_155,In_535,In_998);
xor U156 (N_156,In_124,In_242);
xnor U157 (N_157,In_363,In_117);
nor U158 (N_158,In_477,In_373);
or U159 (N_159,In_26,In_661);
nor U160 (N_160,In_272,In_860);
xor U161 (N_161,In_169,In_374);
nor U162 (N_162,In_663,In_665);
and U163 (N_163,In_48,In_915);
nand U164 (N_164,In_573,In_733);
nand U165 (N_165,In_584,In_624);
or U166 (N_166,In_352,In_930);
and U167 (N_167,In_429,In_219);
xor U168 (N_168,In_152,In_599);
nor U169 (N_169,In_166,In_105);
or U170 (N_170,In_838,In_650);
xor U171 (N_171,In_264,In_325);
nand U172 (N_172,In_285,In_536);
nor U173 (N_173,In_116,In_90);
nand U174 (N_174,In_651,In_994);
nor U175 (N_175,In_113,In_131);
nand U176 (N_176,In_478,In_795);
and U177 (N_177,In_649,In_474);
xnor U178 (N_178,In_427,In_304);
xor U179 (N_179,In_818,In_849);
or U180 (N_180,In_441,In_690);
nor U181 (N_181,In_863,In_890);
and U182 (N_182,In_819,In_431);
and U183 (N_183,In_689,In_672);
and U184 (N_184,In_307,In_471);
or U185 (N_185,In_643,In_520);
nor U186 (N_186,In_22,In_907);
or U187 (N_187,In_647,In_796);
nand U188 (N_188,In_752,In_955);
or U189 (N_189,In_683,In_178);
or U190 (N_190,In_141,In_855);
or U191 (N_191,In_615,In_904);
or U192 (N_192,In_145,In_874);
nand U193 (N_193,In_125,In_114);
or U194 (N_194,In_198,In_289);
xor U195 (N_195,In_227,In_847);
nand U196 (N_196,In_742,In_997);
and U197 (N_197,In_595,In_823);
nor U198 (N_198,In_339,In_937);
xor U199 (N_199,In_184,In_983);
nor U200 (N_200,N_5,In_119);
nor U201 (N_201,In_121,In_764);
xor U202 (N_202,In_11,In_972);
and U203 (N_203,In_866,In_55);
nor U204 (N_204,N_42,In_133);
or U205 (N_205,N_26,In_563);
or U206 (N_206,In_274,In_830);
xnor U207 (N_207,In_197,In_684);
xor U208 (N_208,N_125,In_331);
nor U209 (N_209,In_5,N_198);
nor U210 (N_210,In_28,In_597);
xnor U211 (N_211,N_86,In_540);
and U212 (N_212,In_980,In_696);
nor U213 (N_213,In_542,In_958);
and U214 (N_214,In_334,In_583);
or U215 (N_215,In_414,N_112);
xor U216 (N_216,N_178,In_118);
xnor U217 (N_217,N_54,In_67);
xor U218 (N_218,N_185,In_348);
and U219 (N_219,N_53,In_518);
nor U220 (N_220,In_734,In_610);
nor U221 (N_221,In_612,N_192);
nand U222 (N_222,In_824,N_186);
or U223 (N_223,In_440,N_93);
nor U224 (N_224,N_197,In_985);
or U225 (N_225,In_234,N_149);
nand U226 (N_226,N_3,In_888);
nor U227 (N_227,In_103,In_422);
nand U228 (N_228,In_553,N_156);
nand U229 (N_229,In_578,In_73);
nor U230 (N_230,In_45,In_365);
xor U231 (N_231,In_848,In_957);
xor U232 (N_232,In_992,In_814);
nand U233 (N_233,In_653,In_308);
or U234 (N_234,In_901,In_434);
xor U235 (N_235,N_126,In_202);
nor U236 (N_236,In_882,In_337);
xor U237 (N_237,In_548,In_275);
xnor U238 (N_238,N_72,In_797);
or U239 (N_239,In_614,In_574);
xor U240 (N_240,In_931,In_786);
nor U241 (N_241,In_514,In_41);
nor U242 (N_242,In_767,In_329);
nor U243 (N_243,In_996,N_159);
nand U244 (N_244,N_7,In_716);
or U245 (N_245,In_490,In_918);
xnor U246 (N_246,N_92,N_67);
nand U247 (N_247,N_199,In_35);
nand U248 (N_248,In_755,N_1);
and U249 (N_249,In_450,In_255);
and U250 (N_250,N_13,N_21);
xnor U251 (N_251,In_703,In_314);
nor U252 (N_252,In_537,N_61);
or U253 (N_253,In_633,In_244);
or U254 (N_254,N_32,In_749);
nor U255 (N_255,In_385,In_731);
and U256 (N_256,In_582,In_396);
xor U257 (N_257,In_592,N_194);
xnor U258 (N_258,In_344,In_746);
or U259 (N_259,In_715,In_189);
and U260 (N_260,In_251,In_8);
nor U261 (N_261,In_640,In_475);
or U262 (N_262,N_123,In_942);
xnor U263 (N_263,N_116,N_157);
xnor U264 (N_264,In_132,In_613);
and U265 (N_265,In_741,In_0);
nor U266 (N_266,N_152,In_660);
xnor U267 (N_267,In_130,In_538);
and U268 (N_268,In_765,In_343);
nor U269 (N_269,In_632,In_485);
xor U270 (N_270,N_82,N_147);
nor U271 (N_271,In_248,In_439);
or U272 (N_272,In_273,In_637);
nand U273 (N_273,In_501,In_799);
nand U274 (N_274,In_4,In_351);
and U275 (N_275,In_297,N_31);
and U276 (N_276,In_217,N_153);
nand U277 (N_277,In_69,In_678);
nor U278 (N_278,In_109,In_367);
nand U279 (N_279,In_772,In_81);
xor U280 (N_280,N_155,N_184);
or U281 (N_281,In_498,N_45);
xnor U282 (N_282,N_140,In_629);
nor U283 (N_283,In_713,In_261);
nor U284 (N_284,N_73,N_34);
and U285 (N_285,N_10,In_100);
nor U286 (N_286,N_113,In_443);
xnor U287 (N_287,In_369,N_130);
xor U288 (N_288,N_11,In_357);
xor U289 (N_289,In_943,In_306);
nand U290 (N_290,N_6,In_525);
nand U291 (N_291,In_482,In_497);
xor U292 (N_292,In_727,N_107);
nor U293 (N_293,In_112,In_174);
nand U294 (N_294,In_500,In_76);
and U295 (N_295,N_191,In_89);
and U296 (N_296,N_35,In_59);
or U297 (N_297,N_135,In_515);
nor U298 (N_298,In_303,In_29);
or U299 (N_299,In_777,N_90);
nand U300 (N_300,In_143,In_430);
nand U301 (N_301,In_963,N_151);
nand U302 (N_302,In_916,In_63);
nand U303 (N_303,In_714,In_173);
and U304 (N_304,In_870,In_603);
xor U305 (N_305,In_435,In_56);
xnor U306 (N_306,In_617,In_917);
and U307 (N_307,In_914,In_956);
and U308 (N_308,N_8,In_705);
nand U309 (N_309,In_171,In_700);
and U310 (N_310,In_837,In_389);
nor U311 (N_311,In_753,In_654);
and U312 (N_312,In_362,In_99);
nand U313 (N_313,In_127,In_180);
nand U314 (N_314,In_43,N_170);
nor U315 (N_315,In_577,In_561);
and U316 (N_316,N_9,In_221);
or U317 (N_317,N_17,N_83);
nor U318 (N_318,In_964,In_556);
nor U319 (N_319,N_88,In_758);
xor U320 (N_320,In_185,In_449);
and U321 (N_321,In_827,In_669);
xor U322 (N_322,N_59,N_58);
xnor U323 (N_323,In_395,In_704);
or U324 (N_324,N_142,In_452);
or U325 (N_325,In_86,N_91);
xnor U326 (N_326,In_620,N_84);
nand U327 (N_327,In_628,In_877);
nor U328 (N_328,In_941,In_388);
and U329 (N_329,N_23,N_37);
xnor U330 (N_330,In_962,In_203);
nor U331 (N_331,In_659,N_75);
or U332 (N_332,In_420,In_233);
and U333 (N_333,N_109,In_841);
nor U334 (N_334,In_164,In_903);
and U335 (N_335,N_96,N_110);
nand U336 (N_336,N_137,In_807);
and U337 (N_337,In_892,In_621);
nand U338 (N_338,N_71,In_968);
nor U339 (N_339,In_737,In_147);
nor U340 (N_340,In_257,N_79);
nand U341 (N_341,In_726,In_448);
xnor U342 (N_342,In_639,In_618);
xor U343 (N_343,In_735,In_20);
nand U344 (N_344,In_80,In_249);
nand U345 (N_345,In_208,In_605);
or U346 (N_346,In_883,N_36);
or U347 (N_347,In_260,In_813);
nor U348 (N_348,N_179,N_27);
nor U349 (N_349,In_446,In_889);
nand U350 (N_350,In_122,In_524);
nand U351 (N_351,In_346,In_320);
and U352 (N_352,In_790,In_554);
or U353 (N_353,In_60,In_568);
xor U354 (N_354,In_53,In_216);
xor U355 (N_355,In_51,In_64);
and U356 (N_356,In_865,In_722);
xnor U357 (N_357,In_871,N_50);
nand U358 (N_358,N_99,N_145);
xnor U359 (N_359,In_318,In_938);
nor U360 (N_360,In_87,In_545);
or U361 (N_361,In_466,N_160);
or U362 (N_362,In_825,In_673);
nor U363 (N_363,In_259,N_63);
nand U364 (N_364,N_136,In_24);
xnor U365 (N_365,In_464,In_425);
nor U366 (N_366,In_626,In_840);
nor U367 (N_367,In_359,In_897);
or U368 (N_368,In_856,In_17);
nor U369 (N_369,N_133,In_967);
and U370 (N_370,In_241,In_277);
xor U371 (N_371,In_990,In_456);
or U372 (N_372,In_111,In_214);
nor U373 (N_373,N_174,In_736);
xnor U374 (N_374,N_144,In_361);
nand U375 (N_375,In_294,In_175);
xor U376 (N_376,N_128,In_585);
nor U377 (N_377,In_176,In_873);
or U378 (N_378,In_282,N_77);
and U379 (N_379,In_489,In_820);
nor U380 (N_380,In_47,In_895);
nor U381 (N_381,In_885,In_541);
and U382 (N_382,N_129,In_555);
nand U383 (N_383,In_776,In_225);
xnor U384 (N_384,N_158,N_18);
nand U385 (N_385,In_38,In_745);
and U386 (N_386,In_999,In_666);
nand U387 (N_387,In_301,N_193);
or U388 (N_388,In_79,In_12);
nor U389 (N_389,In_253,In_465);
xnor U390 (N_390,In_648,In_123);
nor U391 (N_391,N_166,In_321);
and U392 (N_392,In_581,In_940);
and U393 (N_393,In_738,In_336);
or U394 (N_394,N_122,In_52);
and U395 (N_395,In_905,N_29);
and U396 (N_396,In_523,N_66);
nand U397 (N_397,In_342,N_188);
or U398 (N_398,N_55,In_622);
and U399 (N_399,N_138,In_165);
nor U400 (N_400,In_82,N_373);
and U401 (N_401,N_187,In_922);
or U402 (N_402,N_294,N_350);
nor U403 (N_403,N_183,In_692);
and U404 (N_404,In_676,N_215);
nand U405 (N_405,N_148,In_258);
nand U406 (N_406,N_180,N_229);
nor U407 (N_407,In_631,N_65);
and U408 (N_408,N_127,In_706);
and U409 (N_409,N_0,N_312);
nand U410 (N_410,In_645,N_47);
and U411 (N_411,N_70,In_656);
and U412 (N_412,N_169,N_393);
or U413 (N_413,In_407,N_276);
xnor U414 (N_414,In_723,In_237);
nand U415 (N_415,N_356,In_218);
or U416 (N_416,N_218,N_94);
nand U417 (N_417,N_318,In_428);
or U418 (N_418,N_234,In_77);
nor U419 (N_419,In_91,In_921);
and U420 (N_420,In_978,N_323);
and U421 (N_421,In_442,N_352);
and U422 (N_422,N_263,N_48);
xnor U423 (N_423,In_356,N_134);
or U424 (N_424,In_779,N_375);
and U425 (N_425,In_46,In_70);
xnor U426 (N_426,N_372,N_300);
xnor U427 (N_427,N_365,In_979);
and U428 (N_428,In_836,In_400);
xor U429 (N_429,In_891,N_33);
xnor U430 (N_430,In_332,N_98);
or U431 (N_431,In_744,In_804);
nor U432 (N_432,In_168,N_251);
and U433 (N_433,N_173,In_693);
and U434 (N_434,In_72,N_101);
nor U435 (N_435,In_698,In_220);
nand U436 (N_436,N_383,N_217);
nor U437 (N_437,In_670,In_701);
nor U438 (N_438,N_319,N_246);
nand U439 (N_439,In_928,N_120);
nor U440 (N_440,N_282,N_222);
xnor U441 (N_441,In_44,N_115);
xor U442 (N_442,In_462,N_390);
and U443 (N_443,N_57,In_276);
and U444 (N_444,In_750,N_230);
or U445 (N_445,In_580,N_195);
nand U446 (N_446,In_394,In_831);
nand U447 (N_447,In_457,N_235);
or U448 (N_448,N_85,In_288);
xnor U449 (N_449,N_271,N_146);
and U450 (N_450,In_424,In_572);
nand U451 (N_451,N_286,N_207);
or U452 (N_452,In_801,In_387);
or U453 (N_453,In_472,N_231);
and U454 (N_454,N_384,In_181);
and U455 (N_455,In_887,In_129);
nand U456 (N_456,N_297,N_81);
nand U457 (N_457,N_68,In_923);
and U458 (N_458,N_267,In_383);
or U459 (N_459,N_287,In_510);
xor U460 (N_460,In_191,N_292);
and U461 (N_461,N_346,In_642);
nand U462 (N_462,In_96,N_4);
nand U463 (N_463,In_451,N_103);
or U464 (N_464,In_341,In_201);
nor U465 (N_465,In_960,In_547);
or U466 (N_466,In_481,N_302);
nand U467 (N_467,In_163,In_236);
nand U468 (N_468,In_778,In_728);
nor U469 (N_469,N_24,N_228);
nor U470 (N_470,In_496,In_616);
nor U471 (N_471,N_366,N_280);
xnor U472 (N_472,N_278,N_76);
and U473 (N_473,N_254,In_993);
nand U474 (N_474,N_196,N_22);
xnor U475 (N_475,N_259,N_248);
and U476 (N_476,N_38,In_906);
and U477 (N_477,N_106,In_695);
xnor U478 (N_478,N_209,N_293);
or U479 (N_479,In_720,N_387);
nor U480 (N_480,In_401,N_182);
nor U481 (N_481,In_447,In_787);
xnor U482 (N_482,N_380,In_808);
xnor U483 (N_483,In_455,N_370);
xor U484 (N_484,N_397,In_926);
nor U485 (N_485,In_108,In_529);
nor U486 (N_486,In_488,N_317);
and U487 (N_487,N_386,In_486);
or U488 (N_488,In_627,N_349);
nand U489 (N_489,In_774,N_143);
or U490 (N_490,In_366,In_23);
nand U491 (N_491,N_398,N_273);
nor U492 (N_492,In_405,N_200);
and U493 (N_493,In_402,N_216);
and U494 (N_494,N_303,N_52);
xor U495 (N_495,N_224,In_193);
or U496 (N_496,In_513,In_231);
xnor U497 (N_497,N_80,N_260);
nand U498 (N_498,In_833,N_379);
xor U499 (N_499,N_270,N_311);
or U500 (N_500,In_668,In_803);
nand U501 (N_501,N_330,In_284);
nand U502 (N_502,N_308,In_950);
xnor U503 (N_503,N_343,N_244);
xor U504 (N_504,N_14,In_929);
and U505 (N_505,In_896,N_43);
and U506 (N_506,In_970,N_12);
nor U507 (N_507,In_725,N_225);
and U508 (N_508,N_392,N_334);
and U509 (N_509,N_291,In_869);
xnor U510 (N_510,In_519,N_290);
xnor U511 (N_511,N_304,N_306);
or U512 (N_512,N_118,In_567);
or U513 (N_513,In_566,In_699);
nor U514 (N_514,N_227,N_313);
nand U515 (N_515,N_320,N_131);
nor U516 (N_516,N_121,In_549);
xnor U517 (N_517,In_558,In_36);
nor U518 (N_518,In_328,In_436);
nand U519 (N_519,In_867,N_223);
and U520 (N_520,N_335,N_213);
and U521 (N_521,In_270,In_534);
nand U522 (N_522,N_351,N_226);
nand U523 (N_523,In_384,In_179);
or U524 (N_524,N_374,In_604);
or U525 (N_525,N_395,N_172);
xor U526 (N_526,N_279,In_854);
nand U527 (N_527,N_295,In_934);
xor U528 (N_528,N_333,In_805);
nand U529 (N_529,N_132,In_740);
nor U530 (N_530,In_406,N_382);
nor U531 (N_531,In_155,In_146);
nand U532 (N_532,In_674,In_315);
or U533 (N_533,In_190,In_754);
xor U534 (N_534,N_255,N_16);
nor U535 (N_535,In_32,N_208);
and U536 (N_536,In_410,N_277);
nand U537 (N_537,In_469,In_426);
nor U538 (N_538,In_913,N_385);
xnor U539 (N_539,In_809,N_249);
nor U540 (N_540,N_325,N_236);
and U541 (N_541,In_350,In_423);
nor U542 (N_542,N_348,N_378);
and U543 (N_543,In_839,In_681);
nor U544 (N_544,In_467,In_381);
nand U545 (N_545,In_769,N_190);
xnor U546 (N_546,N_298,In_710);
xor U547 (N_547,In_312,N_210);
or U548 (N_548,In_691,In_507);
xnor U549 (N_549,In_493,N_275);
nand U550 (N_550,In_594,N_391);
xor U551 (N_551,N_124,In_223);
nor U552 (N_552,In_899,N_338);
and U553 (N_553,In_527,N_321);
nor U554 (N_554,N_388,In_533);
or U555 (N_555,In_313,N_344);
nand U556 (N_556,In_730,In_936);
nor U557 (N_557,N_367,In_589);
xnor U558 (N_558,In_724,In_989);
and U559 (N_559,In_851,In_811);
nor U560 (N_560,In_134,In_140);
nand U561 (N_561,N_212,N_40);
nor U562 (N_562,N_327,N_331);
nor U563 (N_563,N_301,N_205);
and U564 (N_564,In_316,N_240);
nand U565 (N_565,In_569,In_262);
nand U566 (N_566,N_39,In_404);
nor U567 (N_567,N_15,In_959);
nand U568 (N_568,In_458,N_353);
and U569 (N_569,In_115,In_845);
nand U570 (N_570,N_307,In_800);
nor U571 (N_571,In_717,N_141);
xnor U572 (N_572,In_565,N_371);
xor U573 (N_573,In_326,N_60);
or U574 (N_574,N_332,In_502);
nor U575 (N_575,In_945,N_309);
nand U576 (N_576,In_345,N_322);
xnor U577 (N_577,In_946,N_161);
xor U578 (N_578,In_360,N_239);
nor U579 (N_579,N_62,N_176);
nor U580 (N_580,In_794,In_170);
and U581 (N_581,N_283,In_623);
and U582 (N_582,N_203,In_483);
nand U583 (N_583,N_233,N_256);
xnor U584 (N_584,N_368,In_196);
nand U585 (N_585,In_853,In_658);
nor U586 (N_586,N_264,N_167);
xor U587 (N_587,In_878,In_25);
or U588 (N_588,N_269,In_263);
xnor U589 (N_589,N_214,N_87);
nand U590 (N_590,In_499,In_21);
nor U591 (N_591,In_473,In_602);
and U592 (N_592,In_835,In_186);
nand U593 (N_593,N_339,N_108);
and U594 (N_594,In_280,N_201);
and U595 (N_595,N_150,N_296);
or U596 (N_596,N_377,N_51);
nand U597 (N_597,In_415,In_784);
and U598 (N_598,In_154,In_927);
or U599 (N_599,N_104,In_278);
xor U600 (N_600,N_539,In_935);
nand U601 (N_601,N_419,In_657);
xnor U602 (N_602,N_516,N_253);
or U603 (N_603,N_457,N_437);
or U604 (N_604,In_557,N_288);
xnor U605 (N_605,N_447,N_329);
or U606 (N_606,N_451,N_97);
nand U607 (N_607,N_546,N_458);
xor U608 (N_608,N_164,N_399);
xnor U609 (N_609,N_114,In_411);
or U610 (N_610,In_309,N_410);
or U611 (N_611,N_525,N_243);
and U612 (N_612,In_780,N_314);
and U613 (N_613,In_195,N_432);
nand U614 (N_614,N_587,N_404);
xor U615 (N_615,N_247,In_16);
and U616 (N_616,In_757,N_521);
nor U617 (N_617,N_324,N_547);
nor U618 (N_618,N_534,N_44);
xor U619 (N_619,In_27,In_711);
or U620 (N_620,N_500,N_430);
or U621 (N_621,In_600,N_497);
xnor U622 (N_622,In_920,N_464);
and U623 (N_623,N_581,In_662);
xnor U624 (N_624,N_412,In_667);
xor U625 (N_625,N_100,In_49);
nand U626 (N_626,In_476,N_411);
or U627 (N_627,N_206,N_56);
or U628 (N_628,N_502,N_438);
nor U629 (N_629,N_363,N_477);
nand U630 (N_630,In_509,N_445);
nor U631 (N_631,N_30,N_559);
xnor U632 (N_632,N_511,N_396);
nor U633 (N_633,N_274,N_310);
nand U634 (N_634,In_265,In_806);
xor U635 (N_635,N_266,N_20);
and U636 (N_636,N_460,N_95);
and U637 (N_637,In_793,N_455);
xor U638 (N_638,N_337,N_488);
nor U639 (N_639,N_316,N_598);
nor U640 (N_640,In_908,N_541);
nand U641 (N_641,N_484,N_553);
nand U642 (N_642,N_165,N_499);
and U643 (N_643,N_524,N_485);
nor U644 (N_644,N_417,In_495);
or U645 (N_645,In_182,N_119);
or U646 (N_646,N_507,N_468);
and U647 (N_647,In_377,N_328);
or U648 (N_648,N_268,N_509);
nand U649 (N_649,In_31,In_982);
and U650 (N_650,N_505,N_503);
or U651 (N_651,N_394,N_362);
nand U652 (N_652,N_381,N_582);
xnor U653 (N_653,In_751,N_326);
nor U654 (N_654,In_228,N_592);
nand U655 (N_655,N_429,N_245);
and U656 (N_656,N_232,N_416);
and U657 (N_657,In_625,N_237);
nand U658 (N_658,N_550,In_172);
nor U659 (N_659,N_551,In_245);
and U660 (N_660,N_357,In_933);
nand U661 (N_661,N_443,In_974);
xnor U662 (N_662,N_428,N_421);
or U663 (N_663,N_436,N_487);
xor U664 (N_664,N_359,N_486);
and U665 (N_665,N_555,In_880);
nand U666 (N_666,In_370,N_250);
nor U667 (N_667,In_506,N_105);
nand U668 (N_668,N_426,N_354);
or U669 (N_669,N_513,N_469);
and U670 (N_670,N_575,In_894);
or U671 (N_671,N_567,N_219);
nand U672 (N_672,N_496,In_33);
nand U673 (N_673,In_810,N_448);
nand U674 (N_674,In_252,In_763);
nor U675 (N_675,N_483,N_342);
nand U676 (N_676,N_424,N_529);
xor U677 (N_677,N_252,N_538);
or U678 (N_678,In_136,N_591);
nand U679 (N_679,N_489,N_431);
nand U680 (N_680,N_465,N_532);
or U681 (N_681,N_238,N_573);
xor U682 (N_682,In_949,N_498);
xor U683 (N_683,N_470,N_540);
nand U684 (N_684,N_450,N_41);
nor U685 (N_685,N_336,In_743);
xor U686 (N_686,In_947,N_542);
xnor U687 (N_687,N_537,In_789);
nor U688 (N_688,N_117,N_544);
and U689 (N_689,N_568,N_501);
or U690 (N_690,N_520,N_177);
or U691 (N_691,N_401,In_792);
or U692 (N_692,N_413,N_74);
nand U693 (N_693,N_369,N_442);
or U694 (N_694,N_479,N_163);
or U695 (N_695,N_358,In_762);
and U696 (N_696,N_242,N_548);
nor U697 (N_697,N_449,In_192);
nor U698 (N_698,N_418,N_459);
nor U699 (N_699,N_528,N_590);
and U700 (N_700,In_685,In_773);
and U701 (N_701,N_444,N_204);
or U702 (N_702,In_199,N_506);
and U703 (N_703,N_284,N_583);
nor U704 (N_704,In_984,N_355);
nor U705 (N_705,N_361,N_589);
nand U706 (N_706,In_95,N_565);
nand U707 (N_707,N_561,In_135);
and U708 (N_708,N_305,N_425);
nor U709 (N_709,N_466,N_299);
and U710 (N_710,In_919,N_272);
and U711 (N_711,In_463,N_536);
or U712 (N_712,In_126,N_476);
xor U713 (N_713,N_409,N_474);
and U714 (N_714,In_212,N_552);
and U715 (N_715,N_162,In_419);
and U716 (N_716,N_28,N_475);
nand U717 (N_717,N_452,N_480);
xnor U718 (N_718,N_49,N_490);
nor U719 (N_719,N_154,N_533);
xnor U720 (N_720,N_376,N_554);
xor U721 (N_721,N_478,In_512);
nand U722 (N_722,N_512,In_71);
xor U723 (N_723,N_46,N_473);
or U724 (N_724,N_221,N_420);
nand U725 (N_725,N_168,N_440);
nand U726 (N_726,In_40,N_515);
nor U727 (N_727,In_718,In_876);
nor U728 (N_728,N_595,N_523);
or U729 (N_729,N_414,N_171);
xnor U730 (N_730,In_302,N_422);
xor U731 (N_731,In_857,N_570);
nor U732 (N_732,N_588,N_341);
nor U733 (N_733,N_558,N_406);
xnor U734 (N_734,N_405,N_563);
nor U735 (N_735,N_556,N_389);
or U736 (N_736,N_285,In_338);
and U737 (N_737,N_456,In_844);
and U738 (N_738,N_202,In_460);
or U739 (N_739,In_875,N_69);
nand U740 (N_740,N_364,N_89);
or U741 (N_741,N_261,N_102);
nand U742 (N_742,In_355,N_579);
or U743 (N_743,N_19,N_577);
and U744 (N_744,N_522,N_530);
and U745 (N_745,N_434,N_481);
or U746 (N_746,N_531,In_2);
or U747 (N_747,In_378,N_564);
or U748 (N_748,N_211,In_526);
and U749 (N_749,N_111,N_64);
or U750 (N_750,N_574,In_232);
and U751 (N_751,N_175,N_543);
nor U752 (N_752,N_599,N_433);
and U753 (N_753,In_951,In_194);
nand U754 (N_754,N_495,N_494);
or U755 (N_755,N_527,N_78);
and U756 (N_756,N_569,In_413);
and U757 (N_757,N_580,In_785);
nor U758 (N_758,In_7,N_571);
and U759 (N_759,In_292,In_812);
nor U760 (N_760,N_491,In_852);
and U761 (N_761,N_281,N_514);
xor U762 (N_762,In_709,In_19);
nor U763 (N_763,N_407,N_25);
nand U764 (N_764,N_576,N_493);
and U765 (N_765,N_400,N_517);
or U766 (N_766,N_545,N_423);
xnor U767 (N_767,N_572,N_189);
xor U768 (N_768,N_2,N_462);
and U769 (N_769,N_596,N_578);
xnor U770 (N_770,N_472,N_258);
and U771 (N_771,N_345,N_510);
nor U772 (N_772,N_562,N_467);
nor U773 (N_773,N_594,N_262);
nor U774 (N_774,N_526,N_508);
nand U775 (N_775,N_415,N_403);
or U776 (N_776,In_10,N_446);
nor U777 (N_777,In_636,N_549);
nand U778 (N_778,N_519,N_504);
nor U779 (N_779,N_220,In_759);
nand U780 (N_780,N_597,N_535);
nand U781 (N_781,N_585,N_518);
nand U782 (N_782,In_511,In_641);
or U783 (N_783,N_439,N_593);
and U784 (N_784,N_453,N_265);
and U785 (N_785,In_62,N_257);
nand U786 (N_786,N_584,N_471);
xor U787 (N_787,In_505,N_181);
or U788 (N_788,N_435,N_454);
nand U789 (N_789,N_340,In_211);
or U790 (N_790,N_139,N_557);
and U791 (N_791,N_427,In_319);
nand U792 (N_792,In_756,N_241);
xnor U793 (N_793,N_586,N_402);
or U794 (N_794,N_441,N_360);
or U795 (N_795,N_566,N_461);
nand U796 (N_796,N_347,N_492);
xor U797 (N_797,N_408,N_289);
or U798 (N_798,N_315,N_482);
xnor U799 (N_799,N_560,N_463);
or U800 (N_800,N_782,N_721);
nor U801 (N_801,N_749,N_776);
nand U802 (N_802,N_674,N_797);
or U803 (N_803,N_730,N_763);
xor U804 (N_804,N_625,N_619);
nand U805 (N_805,N_767,N_793);
xor U806 (N_806,N_626,N_709);
or U807 (N_807,N_781,N_644);
nor U808 (N_808,N_702,N_613);
nand U809 (N_809,N_679,N_663);
nand U810 (N_810,N_632,N_636);
or U811 (N_811,N_764,N_690);
or U812 (N_812,N_637,N_734);
or U813 (N_813,N_680,N_718);
xor U814 (N_814,N_726,N_668);
nor U815 (N_815,N_617,N_707);
nand U816 (N_816,N_785,N_758);
nand U817 (N_817,N_684,N_645);
nand U818 (N_818,N_760,N_659);
xnor U819 (N_819,N_724,N_687);
xnor U820 (N_820,N_685,N_783);
and U821 (N_821,N_701,N_608);
nand U822 (N_822,N_662,N_729);
nand U823 (N_823,N_683,N_706);
nand U824 (N_824,N_694,N_735);
nand U825 (N_825,N_642,N_635);
and U826 (N_826,N_720,N_631);
and U827 (N_827,N_745,N_778);
nand U828 (N_828,N_689,N_751);
nand U829 (N_829,N_603,N_743);
and U830 (N_830,N_670,N_789);
and U831 (N_831,N_601,N_747);
nor U832 (N_832,N_616,N_657);
nor U833 (N_833,N_630,N_736);
and U834 (N_834,N_737,N_739);
and U835 (N_835,N_667,N_704);
and U836 (N_836,N_646,N_725);
or U837 (N_837,N_634,N_715);
and U838 (N_838,N_777,N_699);
or U839 (N_839,N_703,N_688);
and U840 (N_840,N_677,N_748);
and U841 (N_841,N_757,N_710);
or U842 (N_842,N_638,N_744);
nor U843 (N_843,N_798,N_605);
nand U844 (N_844,N_666,N_711);
nor U845 (N_845,N_772,N_686);
nor U846 (N_846,N_697,N_600);
nand U847 (N_847,N_787,N_672);
nor U848 (N_848,N_713,N_673);
nor U849 (N_849,N_615,N_682);
and U850 (N_850,N_692,N_658);
nor U851 (N_851,N_602,N_746);
and U852 (N_852,N_653,N_648);
or U853 (N_853,N_728,N_780);
or U854 (N_854,N_762,N_795);
nor U855 (N_855,N_705,N_671);
or U856 (N_856,N_651,N_611);
and U857 (N_857,N_622,N_714);
xnor U858 (N_858,N_652,N_691);
and U859 (N_859,N_627,N_738);
or U860 (N_860,N_770,N_765);
and U861 (N_861,N_769,N_761);
nand U862 (N_862,N_722,N_607);
and U863 (N_863,N_784,N_654);
nor U864 (N_864,N_773,N_639);
xnor U865 (N_865,N_733,N_731);
or U866 (N_866,N_609,N_664);
nand U867 (N_867,N_641,N_640);
xor U868 (N_868,N_768,N_693);
and U869 (N_869,N_796,N_792);
or U870 (N_870,N_698,N_650);
and U871 (N_871,N_620,N_759);
and U872 (N_872,N_696,N_661);
and U873 (N_873,N_604,N_771);
and U874 (N_874,N_755,N_676);
xor U875 (N_875,N_712,N_628);
nand U876 (N_876,N_788,N_756);
xor U877 (N_877,N_790,N_695);
nand U878 (N_878,N_754,N_669);
and U879 (N_879,N_752,N_675);
xnor U880 (N_880,N_629,N_612);
and U881 (N_881,N_740,N_621);
nor U882 (N_882,N_723,N_775);
or U883 (N_883,N_649,N_610);
nand U884 (N_884,N_779,N_624);
xnor U885 (N_885,N_606,N_647);
or U886 (N_886,N_660,N_623);
nor U887 (N_887,N_633,N_716);
nand U888 (N_888,N_766,N_727);
or U889 (N_889,N_786,N_732);
or U890 (N_890,N_708,N_717);
nor U891 (N_891,N_741,N_794);
or U892 (N_892,N_665,N_742);
or U893 (N_893,N_791,N_700);
xnor U894 (N_894,N_681,N_719);
nor U895 (N_895,N_655,N_614);
and U896 (N_896,N_656,N_678);
xnor U897 (N_897,N_750,N_799);
nor U898 (N_898,N_643,N_774);
and U899 (N_899,N_618,N_753);
xnor U900 (N_900,N_711,N_717);
xnor U901 (N_901,N_748,N_788);
nand U902 (N_902,N_653,N_796);
nor U903 (N_903,N_609,N_792);
xor U904 (N_904,N_636,N_796);
nand U905 (N_905,N_704,N_749);
nand U906 (N_906,N_678,N_708);
nor U907 (N_907,N_615,N_760);
xnor U908 (N_908,N_675,N_605);
or U909 (N_909,N_755,N_649);
nand U910 (N_910,N_719,N_790);
xor U911 (N_911,N_702,N_686);
and U912 (N_912,N_742,N_628);
and U913 (N_913,N_769,N_665);
and U914 (N_914,N_613,N_799);
and U915 (N_915,N_691,N_711);
and U916 (N_916,N_793,N_666);
nand U917 (N_917,N_756,N_650);
and U918 (N_918,N_799,N_798);
nand U919 (N_919,N_676,N_770);
and U920 (N_920,N_699,N_687);
and U921 (N_921,N_655,N_777);
nand U922 (N_922,N_666,N_651);
and U923 (N_923,N_766,N_770);
nand U924 (N_924,N_682,N_601);
nand U925 (N_925,N_672,N_619);
nand U926 (N_926,N_716,N_778);
and U927 (N_927,N_616,N_770);
xor U928 (N_928,N_756,N_711);
xor U929 (N_929,N_779,N_787);
nand U930 (N_930,N_753,N_754);
or U931 (N_931,N_728,N_783);
and U932 (N_932,N_748,N_671);
or U933 (N_933,N_668,N_646);
nor U934 (N_934,N_608,N_639);
nor U935 (N_935,N_668,N_622);
nor U936 (N_936,N_685,N_790);
nand U937 (N_937,N_696,N_703);
or U938 (N_938,N_714,N_780);
or U939 (N_939,N_673,N_652);
nand U940 (N_940,N_721,N_615);
xor U941 (N_941,N_643,N_726);
xor U942 (N_942,N_627,N_639);
nor U943 (N_943,N_658,N_677);
or U944 (N_944,N_687,N_746);
nand U945 (N_945,N_755,N_785);
xor U946 (N_946,N_611,N_783);
and U947 (N_947,N_793,N_691);
nor U948 (N_948,N_691,N_621);
nor U949 (N_949,N_724,N_768);
nor U950 (N_950,N_711,N_767);
nand U951 (N_951,N_612,N_698);
xnor U952 (N_952,N_689,N_675);
or U953 (N_953,N_679,N_686);
and U954 (N_954,N_714,N_682);
or U955 (N_955,N_790,N_736);
and U956 (N_956,N_682,N_715);
nand U957 (N_957,N_675,N_660);
nor U958 (N_958,N_672,N_638);
nand U959 (N_959,N_666,N_618);
and U960 (N_960,N_637,N_634);
or U961 (N_961,N_761,N_741);
and U962 (N_962,N_770,N_741);
or U963 (N_963,N_651,N_778);
nand U964 (N_964,N_610,N_719);
and U965 (N_965,N_654,N_636);
nand U966 (N_966,N_744,N_673);
and U967 (N_967,N_789,N_622);
nand U968 (N_968,N_738,N_786);
xor U969 (N_969,N_799,N_796);
or U970 (N_970,N_784,N_630);
xor U971 (N_971,N_791,N_652);
nor U972 (N_972,N_786,N_603);
xnor U973 (N_973,N_645,N_679);
or U974 (N_974,N_714,N_786);
and U975 (N_975,N_630,N_770);
nor U976 (N_976,N_659,N_666);
nand U977 (N_977,N_644,N_638);
xnor U978 (N_978,N_790,N_766);
nand U979 (N_979,N_751,N_759);
nor U980 (N_980,N_662,N_718);
nor U981 (N_981,N_731,N_779);
nor U982 (N_982,N_707,N_717);
and U983 (N_983,N_643,N_624);
or U984 (N_984,N_686,N_642);
nor U985 (N_985,N_644,N_607);
or U986 (N_986,N_715,N_621);
xor U987 (N_987,N_635,N_731);
xnor U988 (N_988,N_628,N_648);
or U989 (N_989,N_645,N_697);
and U990 (N_990,N_761,N_757);
nand U991 (N_991,N_712,N_765);
xor U992 (N_992,N_733,N_728);
nand U993 (N_993,N_762,N_775);
nor U994 (N_994,N_725,N_773);
nor U995 (N_995,N_733,N_626);
nor U996 (N_996,N_742,N_705);
nand U997 (N_997,N_730,N_628);
and U998 (N_998,N_720,N_759);
nand U999 (N_999,N_724,N_658);
and U1000 (N_1000,N_986,N_817);
or U1001 (N_1001,N_931,N_849);
nand U1002 (N_1002,N_956,N_848);
xor U1003 (N_1003,N_900,N_871);
and U1004 (N_1004,N_930,N_832);
xnor U1005 (N_1005,N_807,N_912);
nand U1006 (N_1006,N_854,N_915);
or U1007 (N_1007,N_935,N_815);
or U1008 (N_1008,N_914,N_934);
and U1009 (N_1009,N_928,N_949);
nand U1010 (N_1010,N_992,N_951);
or U1011 (N_1011,N_975,N_824);
nor U1012 (N_1012,N_836,N_963);
nor U1013 (N_1013,N_907,N_864);
nor U1014 (N_1014,N_853,N_976);
nand U1015 (N_1015,N_978,N_991);
xor U1016 (N_1016,N_879,N_926);
and U1017 (N_1017,N_958,N_985);
and U1018 (N_1018,N_881,N_882);
xor U1019 (N_1019,N_897,N_938);
or U1020 (N_1020,N_954,N_970);
nand U1021 (N_1021,N_961,N_920);
xnor U1022 (N_1022,N_875,N_862);
or U1023 (N_1023,N_910,N_966);
or U1024 (N_1024,N_837,N_982);
nor U1025 (N_1025,N_808,N_813);
or U1026 (N_1026,N_841,N_932);
xnor U1027 (N_1027,N_923,N_916);
nand U1028 (N_1028,N_867,N_964);
nor U1029 (N_1029,N_884,N_904);
nor U1030 (N_1030,N_840,N_901);
xor U1031 (N_1031,N_973,N_895);
or U1032 (N_1032,N_859,N_857);
or U1033 (N_1033,N_947,N_936);
and U1034 (N_1034,N_816,N_814);
or U1035 (N_1035,N_998,N_869);
nor U1036 (N_1036,N_967,N_969);
xnor U1037 (N_1037,N_908,N_903);
or U1038 (N_1038,N_996,N_819);
nand U1039 (N_1039,N_922,N_870);
nor U1040 (N_1040,N_833,N_863);
or U1041 (N_1041,N_825,N_890);
xor U1042 (N_1042,N_979,N_925);
xnor U1043 (N_1043,N_866,N_946);
or U1044 (N_1044,N_858,N_850);
or U1045 (N_1045,N_942,N_803);
nand U1046 (N_1046,N_905,N_885);
and U1047 (N_1047,N_899,N_945);
nand U1048 (N_1048,N_812,N_893);
or U1049 (N_1049,N_980,N_820);
xor U1050 (N_1050,N_906,N_948);
or U1051 (N_1051,N_886,N_801);
or U1052 (N_1052,N_944,N_883);
nor U1053 (N_1053,N_913,N_962);
nor U1054 (N_1054,N_918,N_984);
and U1055 (N_1055,N_878,N_983);
or U1056 (N_1056,N_818,N_810);
nor U1057 (N_1057,N_995,N_826);
nor U1058 (N_1058,N_856,N_887);
nand U1059 (N_1059,N_929,N_873);
xor U1060 (N_1060,N_872,N_909);
or U1061 (N_1061,N_874,N_927);
nor U1062 (N_1062,N_971,N_894);
nor U1063 (N_1063,N_835,N_999);
or U1064 (N_1064,N_804,N_851);
nand U1065 (N_1065,N_843,N_953);
nor U1066 (N_1066,N_993,N_952);
or U1067 (N_1067,N_990,N_941);
and U1068 (N_1068,N_827,N_981);
xor U1069 (N_1069,N_888,N_809);
nand U1070 (N_1070,N_823,N_847);
nand U1071 (N_1071,N_891,N_852);
nand U1072 (N_1072,N_940,N_974);
nand U1073 (N_1073,N_805,N_800);
nand U1074 (N_1074,N_831,N_917);
xor U1075 (N_1075,N_844,N_834);
nor U1076 (N_1076,N_939,N_911);
nand U1077 (N_1077,N_921,N_902);
xnor U1078 (N_1078,N_898,N_937);
and U1079 (N_1079,N_968,N_806);
nand U1080 (N_1080,N_988,N_959);
and U1081 (N_1081,N_924,N_802);
xor U1082 (N_1082,N_994,N_839);
nor U1083 (N_1083,N_829,N_861);
and U1084 (N_1084,N_972,N_828);
nand U1085 (N_1085,N_846,N_860);
nor U1086 (N_1086,N_877,N_977);
and U1087 (N_1087,N_943,N_868);
xor U1088 (N_1088,N_842,N_960);
or U1089 (N_1089,N_880,N_955);
xor U1090 (N_1090,N_855,N_950);
nand U1091 (N_1091,N_876,N_987);
xnor U1092 (N_1092,N_821,N_965);
or U1093 (N_1093,N_889,N_845);
and U1094 (N_1094,N_989,N_957);
or U1095 (N_1095,N_892,N_997);
and U1096 (N_1096,N_896,N_838);
xor U1097 (N_1097,N_830,N_811);
nor U1098 (N_1098,N_822,N_865);
and U1099 (N_1099,N_919,N_933);
and U1100 (N_1100,N_935,N_893);
nand U1101 (N_1101,N_872,N_807);
or U1102 (N_1102,N_939,N_895);
nand U1103 (N_1103,N_813,N_845);
nor U1104 (N_1104,N_996,N_903);
and U1105 (N_1105,N_840,N_801);
xor U1106 (N_1106,N_958,N_887);
xor U1107 (N_1107,N_954,N_984);
nor U1108 (N_1108,N_863,N_837);
and U1109 (N_1109,N_990,N_898);
xnor U1110 (N_1110,N_948,N_890);
nor U1111 (N_1111,N_843,N_990);
nand U1112 (N_1112,N_980,N_828);
xnor U1113 (N_1113,N_848,N_913);
and U1114 (N_1114,N_897,N_850);
nor U1115 (N_1115,N_813,N_937);
nand U1116 (N_1116,N_980,N_972);
nor U1117 (N_1117,N_897,N_876);
or U1118 (N_1118,N_841,N_919);
or U1119 (N_1119,N_932,N_966);
and U1120 (N_1120,N_958,N_827);
nand U1121 (N_1121,N_936,N_826);
or U1122 (N_1122,N_841,N_856);
nor U1123 (N_1123,N_830,N_955);
nand U1124 (N_1124,N_940,N_899);
nand U1125 (N_1125,N_978,N_954);
or U1126 (N_1126,N_939,N_986);
nand U1127 (N_1127,N_815,N_824);
nand U1128 (N_1128,N_825,N_820);
nand U1129 (N_1129,N_847,N_874);
nand U1130 (N_1130,N_804,N_971);
xnor U1131 (N_1131,N_884,N_867);
or U1132 (N_1132,N_991,N_886);
and U1133 (N_1133,N_853,N_802);
nand U1134 (N_1134,N_821,N_973);
xor U1135 (N_1135,N_961,N_905);
xor U1136 (N_1136,N_943,N_902);
and U1137 (N_1137,N_872,N_947);
nor U1138 (N_1138,N_847,N_873);
nor U1139 (N_1139,N_975,N_835);
nor U1140 (N_1140,N_890,N_906);
nor U1141 (N_1141,N_965,N_942);
nand U1142 (N_1142,N_924,N_800);
nor U1143 (N_1143,N_916,N_921);
xnor U1144 (N_1144,N_833,N_955);
nand U1145 (N_1145,N_826,N_955);
and U1146 (N_1146,N_845,N_863);
xor U1147 (N_1147,N_958,N_910);
nand U1148 (N_1148,N_919,N_802);
nor U1149 (N_1149,N_881,N_861);
nand U1150 (N_1150,N_959,N_814);
or U1151 (N_1151,N_965,N_847);
or U1152 (N_1152,N_817,N_892);
and U1153 (N_1153,N_831,N_836);
nor U1154 (N_1154,N_962,N_858);
nor U1155 (N_1155,N_807,N_941);
nand U1156 (N_1156,N_825,N_979);
nand U1157 (N_1157,N_943,N_989);
and U1158 (N_1158,N_840,N_804);
nor U1159 (N_1159,N_855,N_817);
xor U1160 (N_1160,N_990,N_841);
nor U1161 (N_1161,N_940,N_891);
nand U1162 (N_1162,N_963,N_848);
and U1163 (N_1163,N_994,N_867);
nand U1164 (N_1164,N_858,N_960);
or U1165 (N_1165,N_843,N_824);
and U1166 (N_1166,N_818,N_814);
xnor U1167 (N_1167,N_877,N_810);
nand U1168 (N_1168,N_808,N_946);
or U1169 (N_1169,N_962,N_908);
nor U1170 (N_1170,N_997,N_866);
nand U1171 (N_1171,N_883,N_881);
nand U1172 (N_1172,N_862,N_908);
or U1173 (N_1173,N_841,N_884);
and U1174 (N_1174,N_912,N_907);
nor U1175 (N_1175,N_828,N_865);
nand U1176 (N_1176,N_998,N_862);
nand U1177 (N_1177,N_819,N_867);
nand U1178 (N_1178,N_962,N_911);
and U1179 (N_1179,N_820,N_864);
nand U1180 (N_1180,N_968,N_985);
nor U1181 (N_1181,N_883,N_870);
nand U1182 (N_1182,N_906,N_957);
and U1183 (N_1183,N_910,N_906);
xnor U1184 (N_1184,N_869,N_854);
xor U1185 (N_1185,N_873,N_960);
xor U1186 (N_1186,N_992,N_872);
nor U1187 (N_1187,N_920,N_895);
nor U1188 (N_1188,N_843,N_878);
nand U1189 (N_1189,N_919,N_996);
nor U1190 (N_1190,N_997,N_834);
nor U1191 (N_1191,N_994,N_882);
or U1192 (N_1192,N_952,N_926);
nor U1193 (N_1193,N_920,N_930);
nand U1194 (N_1194,N_868,N_951);
nor U1195 (N_1195,N_900,N_849);
or U1196 (N_1196,N_959,N_991);
or U1197 (N_1197,N_866,N_899);
xnor U1198 (N_1198,N_959,N_864);
nand U1199 (N_1199,N_965,N_851);
nor U1200 (N_1200,N_1156,N_1075);
or U1201 (N_1201,N_1071,N_1130);
nor U1202 (N_1202,N_1103,N_1064);
nand U1203 (N_1203,N_1134,N_1050);
nor U1204 (N_1204,N_1089,N_1128);
nand U1205 (N_1205,N_1013,N_1179);
xor U1206 (N_1206,N_1092,N_1026);
nor U1207 (N_1207,N_1029,N_1042);
nor U1208 (N_1208,N_1030,N_1043);
or U1209 (N_1209,N_1052,N_1021);
nand U1210 (N_1210,N_1153,N_1188);
or U1211 (N_1211,N_1184,N_1161);
nand U1212 (N_1212,N_1139,N_1058);
and U1213 (N_1213,N_1081,N_1023);
xnor U1214 (N_1214,N_1121,N_1066);
nand U1215 (N_1215,N_1119,N_1025);
nand U1216 (N_1216,N_1088,N_1004);
nor U1217 (N_1217,N_1093,N_1032);
and U1218 (N_1218,N_1149,N_1138);
or U1219 (N_1219,N_1125,N_1067);
or U1220 (N_1220,N_1057,N_1129);
nor U1221 (N_1221,N_1082,N_1054);
nand U1222 (N_1222,N_1018,N_1123);
or U1223 (N_1223,N_1173,N_1022);
or U1224 (N_1224,N_1199,N_1051);
and U1225 (N_1225,N_1176,N_1187);
and U1226 (N_1226,N_1024,N_1132);
or U1227 (N_1227,N_1001,N_1116);
xor U1228 (N_1228,N_1078,N_1014);
and U1229 (N_1229,N_1155,N_1069);
and U1230 (N_1230,N_1056,N_1095);
and U1231 (N_1231,N_1037,N_1118);
and U1232 (N_1232,N_1099,N_1146);
nand U1233 (N_1233,N_1106,N_1198);
or U1234 (N_1234,N_1062,N_1005);
and U1235 (N_1235,N_1133,N_1197);
xor U1236 (N_1236,N_1105,N_1060);
xor U1237 (N_1237,N_1152,N_1114);
nand U1238 (N_1238,N_1080,N_1124);
nand U1239 (N_1239,N_1148,N_1035);
nand U1240 (N_1240,N_1034,N_1158);
and U1241 (N_1241,N_1190,N_1140);
and U1242 (N_1242,N_1175,N_1151);
or U1243 (N_1243,N_1010,N_1192);
and U1244 (N_1244,N_1097,N_1015);
xor U1245 (N_1245,N_1036,N_1061);
xnor U1246 (N_1246,N_1104,N_1033);
and U1247 (N_1247,N_1112,N_1055);
xnor U1248 (N_1248,N_1186,N_1193);
or U1249 (N_1249,N_1012,N_1028);
and U1250 (N_1250,N_1086,N_1181);
nand U1251 (N_1251,N_1145,N_1059);
or U1252 (N_1252,N_1006,N_1084);
and U1253 (N_1253,N_1044,N_1194);
nor U1254 (N_1254,N_1142,N_1031);
nand U1255 (N_1255,N_1111,N_1045);
nand U1256 (N_1256,N_1027,N_1016);
xor U1257 (N_1257,N_1000,N_1127);
and U1258 (N_1258,N_1172,N_1048);
xor U1259 (N_1259,N_1040,N_1191);
and U1260 (N_1260,N_1136,N_1108);
nor U1261 (N_1261,N_1195,N_1115);
or U1262 (N_1262,N_1068,N_1094);
or U1263 (N_1263,N_1019,N_1162);
nand U1264 (N_1264,N_1180,N_1144);
nor U1265 (N_1265,N_1167,N_1120);
or U1266 (N_1266,N_1169,N_1003);
xor U1267 (N_1267,N_1131,N_1185);
xor U1268 (N_1268,N_1159,N_1090);
xor U1269 (N_1269,N_1072,N_1171);
or U1270 (N_1270,N_1110,N_1076);
or U1271 (N_1271,N_1007,N_1137);
and U1272 (N_1272,N_1098,N_1083);
or U1273 (N_1273,N_1135,N_1147);
nand U1274 (N_1274,N_1070,N_1168);
nand U1275 (N_1275,N_1107,N_1164);
xor U1276 (N_1276,N_1174,N_1177);
and U1277 (N_1277,N_1183,N_1087);
or U1278 (N_1278,N_1063,N_1038);
and U1279 (N_1279,N_1160,N_1178);
and U1280 (N_1280,N_1143,N_1020);
xor U1281 (N_1281,N_1085,N_1182);
nand U1282 (N_1282,N_1041,N_1196);
nand U1283 (N_1283,N_1073,N_1049);
or U1284 (N_1284,N_1122,N_1079);
or U1285 (N_1285,N_1150,N_1113);
or U1286 (N_1286,N_1002,N_1065);
and U1287 (N_1287,N_1102,N_1096);
xor U1288 (N_1288,N_1077,N_1047);
and U1289 (N_1289,N_1101,N_1141);
nor U1290 (N_1290,N_1074,N_1009);
or U1291 (N_1291,N_1163,N_1166);
and U1292 (N_1292,N_1109,N_1100);
xor U1293 (N_1293,N_1053,N_1039);
nor U1294 (N_1294,N_1011,N_1170);
nor U1295 (N_1295,N_1017,N_1189);
and U1296 (N_1296,N_1117,N_1008);
and U1297 (N_1297,N_1165,N_1154);
xor U1298 (N_1298,N_1091,N_1126);
and U1299 (N_1299,N_1157,N_1046);
nand U1300 (N_1300,N_1010,N_1197);
nor U1301 (N_1301,N_1168,N_1165);
nor U1302 (N_1302,N_1083,N_1081);
xnor U1303 (N_1303,N_1130,N_1079);
nand U1304 (N_1304,N_1159,N_1033);
nor U1305 (N_1305,N_1134,N_1183);
nand U1306 (N_1306,N_1005,N_1041);
and U1307 (N_1307,N_1182,N_1016);
nand U1308 (N_1308,N_1029,N_1101);
and U1309 (N_1309,N_1114,N_1153);
and U1310 (N_1310,N_1030,N_1102);
xnor U1311 (N_1311,N_1174,N_1199);
xor U1312 (N_1312,N_1076,N_1126);
or U1313 (N_1313,N_1132,N_1047);
or U1314 (N_1314,N_1181,N_1164);
nand U1315 (N_1315,N_1148,N_1107);
nor U1316 (N_1316,N_1154,N_1186);
and U1317 (N_1317,N_1129,N_1132);
xnor U1318 (N_1318,N_1164,N_1154);
or U1319 (N_1319,N_1196,N_1116);
xnor U1320 (N_1320,N_1169,N_1012);
xnor U1321 (N_1321,N_1068,N_1180);
nor U1322 (N_1322,N_1140,N_1068);
xor U1323 (N_1323,N_1052,N_1029);
nand U1324 (N_1324,N_1197,N_1042);
nand U1325 (N_1325,N_1163,N_1012);
and U1326 (N_1326,N_1124,N_1034);
or U1327 (N_1327,N_1029,N_1188);
or U1328 (N_1328,N_1044,N_1024);
or U1329 (N_1329,N_1170,N_1062);
or U1330 (N_1330,N_1010,N_1017);
nor U1331 (N_1331,N_1124,N_1078);
nor U1332 (N_1332,N_1037,N_1188);
and U1333 (N_1333,N_1047,N_1061);
or U1334 (N_1334,N_1179,N_1159);
or U1335 (N_1335,N_1030,N_1169);
or U1336 (N_1336,N_1089,N_1182);
or U1337 (N_1337,N_1090,N_1145);
xnor U1338 (N_1338,N_1169,N_1109);
nand U1339 (N_1339,N_1119,N_1139);
and U1340 (N_1340,N_1007,N_1198);
nand U1341 (N_1341,N_1030,N_1113);
nand U1342 (N_1342,N_1088,N_1101);
xnor U1343 (N_1343,N_1197,N_1108);
nand U1344 (N_1344,N_1004,N_1059);
or U1345 (N_1345,N_1174,N_1118);
nand U1346 (N_1346,N_1124,N_1151);
nor U1347 (N_1347,N_1196,N_1001);
and U1348 (N_1348,N_1110,N_1129);
xor U1349 (N_1349,N_1117,N_1068);
and U1350 (N_1350,N_1104,N_1026);
and U1351 (N_1351,N_1087,N_1196);
and U1352 (N_1352,N_1076,N_1146);
and U1353 (N_1353,N_1009,N_1069);
or U1354 (N_1354,N_1180,N_1028);
xor U1355 (N_1355,N_1029,N_1127);
and U1356 (N_1356,N_1093,N_1008);
nand U1357 (N_1357,N_1015,N_1187);
nor U1358 (N_1358,N_1187,N_1198);
nor U1359 (N_1359,N_1003,N_1053);
xnor U1360 (N_1360,N_1156,N_1068);
nor U1361 (N_1361,N_1011,N_1186);
xor U1362 (N_1362,N_1103,N_1080);
nand U1363 (N_1363,N_1100,N_1092);
xor U1364 (N_1364,N_1174,N_1098);
or U1365 (N_1365,N_1017,N_1045);
nor U1366 (N_1366,N_1003,N_1122);
or U1367 (N_1367,N_1066,N_1178);
nand U1368 (N_1368,N_1075,N_1032);
nor U1369 (N_1369,N_1184,N_1086);
xor U1370 (N_1370,N_1135,N_1098);
xor U1371 (N_1371,N_1038,N_1073);
or U1372 (N_1372,N_1142,N_1160);
or U1373 (N_1373,N_1061,N_1115);
xnor U1374 (N_1374,N_1084,N_1115);
nor U1375 (N_1375,N_1077,N_1072);
nand U1376 (N_1376,N_1114,N_1155);
xnor U1377 (N_1377,N_1121,N_1027);
nor U1378 (N_1378,N_1050,N_1031);
or U1379 (N_1379,N_1189,N_1053);
nand U1380 (N_1380,N_1048,N_1184);
xor U1381 (N_1381,N_1115,N_1138);
nor U1382 (N_1382,N_1194,N_1149);
nor U1383 (N_1383,N_1047,N_1011);
nor U1384 (N_1384,N_1139,N_1117);
or U1385 (N_1385,N_1102,N_1078);
nand U1386 (N_1386,N_1135,N_1165);
nor U1387 (N_1387,N_1010,N_1133);
nand U1388 (N_1388,N_1115,N_1167);
nand U1389 (N_1389,N_1081,N_1067);
nand U1390 (N_1390,N_1184,N_1078);
and U1391 (N_1391,N_1114,N_1008);
nor U1392 (N_1392,N_1103,N_1075);
and U1393 (N_1393,N_1087,N_1106);
nand U1394 (N_1394,N_1045,N_1057);
xor U1395 (N_1395,N_1100,N_1170);
nand U1396 (N_1396,N_1015,N_1115);
nand U1397 (N_1397,N_1023,N_1176);
xor U1398 (N_1398,N_1144,N_1199);
xnor U1399 (N_1399,N_1183,N_1151);
or U1400 (N_1400,N_1322,N_1250);
and U1401 (N_1401,N_1303,N_1383);
or U1402 (N_1402,N_1293,N_1287);
or U1403 (N_1403,N_1291,N_1331);
and U1404 (N_1404,N_1329,N_1355);
nor U1405 (N_1405,N_1392,N_1320);
xor U1406 (N_1406,N_1248,N_1267);
and U1407 (N_1407,N_1274,N_1339);
nor U1408 (N_1408,N_1321,N_1237);
xor U1409 (N_1409,N_1273,N_1368);
nor U1410 (N_1410,N_1288,N_1387);
xor U1411 (N_1411,N_1280,N_1292);
and U1412 (N_1412,N_1359,N_1312);
xor U1413 (N_1413,N_1294,N_1212);
and U1414 (N_1414,N_1390,N_1367);
and U1415 (N_1415,N_1342,N_1268);
nor U1416 (N_1416,N_1344,N_1300);
nand U1417 (N_1417,N_1297,N_1253);
xnor U1418 (N_1418,N_1216,N_1333);
nand U1419 (N_1419,N_1286,N_1228);
xor U1420 (N_1420,N_1346,N_1213);
nand U1421 (N_1421,N_1371,N_1307);
nand U1422 (N_1422,N_1222,N_1337);
nor U1423 (N_1423,N_1356,N_1374);
xnor U1424 (N_1424,N_1334,N_1317);
nand U1425 (N_1425,N_1323,N_1231);
nor U1426 (N_1426,N_1394,N_1330);
and U1427 (N_1427,N_1207,N_1245);
nand U1428 (N_1428,N_1380,N_1397);
nor U1429 (N_1429,N_1360,N_1296);
nor U1430 (N_1430,N_1234,N_1233);
nand U1431 (N_1431,N_1388,N_1350);
nand U1432 (N_1432,N_1332,N_1217);
or U1433 (N_1433,N_1283,N_1271);
nor U1434 (N_1434,N_1252,N_1313);
nor U1435 (N_1435,N_1247,N_1362);
or U1436 (N_1436,N_1364,N_1395);
and U1437 (N_1437,N_1311,N_1206);
nor U1438 (N_1438,N_1304,N_1200);
nor U1439 (N_1439,N_1255,N_1325);
nor U1440 (N_1440,N_1351,N_1336);
xnor U1441 (N_1441,N_1232,N_1315);
nor U1442 (N_1442,N_1279,N_1347);
nand U1443 (N_1443,N_1257,N_1201);
or U1444 (N_1444,N_1378,N_1377);
and U1445 (N_1445,N_1361,N_1215);
nor U1446 (N_1446,N_1272,N_1246);
xnor U1447 (N_1447,N_1389,N_1306);
and U1448 (N_1448,N_1264,N_1308);
nor U1449 (N_1449,N_1240,N_1370);
or U1450 (N_1450,N_1352,N_1243);
and U1451 (N_1451,N_1261,N_1372);
xor U1452 (N_1452,N_1242,N_1373);
or U1453 (N_1453,N_1358,N_1230);
nand U1454 (N_1454,N_1276,N_1254);
and U1455 (N_1455,N_1298,N_1365);
nor U1456 (N_1456,N_1284,N_1341);
nor U1457 (N_1457,N_1345,N_1326);
and U1458 (N_1458,N_1316,N_1393);
nor U1459 (N_1459,N_1302,N_1309);
and U1460 (N_1460,N_1295,N_1369);
nor U1461 (N_1461,N_1266,N_1241);
nor U1462 (N_1462,N_1310,N_1275);
and U1463 (N_1463,N_1260,N_1343);
nand U1464 (N_1464,N_1204,N_1210);
and U1465 (N_1465,N_1375,N_1376);
nor U1466 (N_1466,N_1269,N_1229);
nor U1467 (N_1467,N_1396,N_1220);
and U1468 (N_1468,N_1305,N_1219);
and U1469 (N_1469,N_1244,N_1224);
nand U1470 (N_1470,N_1235,N_1209);
xor U1471 (N_1471,N_1270,N_1236);
or U1472 (N_1472,N_1357,N_1382);
nor U1473 (N_1473,N_1262,N_1314);
nand U1474 (N_1474,N_1214,N_1223);
nor U1475 (N_1475,N_1328,N_1354);
nor U1476 (N_1476,N_1281,N_1318);
xnor U1477 (N_1477,N_1258,N_1208);
nor U1478 (N_1478,N_1239,N_1265);
xnor U1479 (N_1479,N_1301,N_1340);
or U1480 (N_1480,N_1227,N_1327);
xnor U1481 (N_1481,N_1259,N_1353);
and U1482 (N_1482,N_1384,N_1290);
and U1483 (N_1483,N_1319,N_1203);
nand U1484 (N_1484,N_1205,N_1277);
nand U1485 (N_1485,N_1381,N_1289);
and U1486 (N_1486,N_1226,N_1249);
and U1487 (N_1487,N_1335,N_1386);
or U1488 (N_1488,N_1202,N_1366);
or U1489 (N_1489,N_1238,N_1349);
xnor U1490 (N_1490,N_1385,N_1218);
or U1491 (N_1491,N_1221,N_1379);
xor U1492 (N_1492,N_1225,N_1211);
nand U1493 (N_1493,N_1256,N_1348);
nand U1494 (N_1494,N_1399,N_1251);
or U1495 (N_1495,N_1299,N_1338);
nor U1496 (N_1496,N_1398,N_1278);
nand U1497 (N_1497,N_1263,N_1282);
nand U1498 (N_1498,N_1363,N_1391);
or U1499 (N_1499,N_1324,N_1285);
nor U1500 (N_1500,N_1306,N_1235);
nand U1501 (N_1501,N_1398,N_1211);
or U1502 (N_1502,N_1320,N_1350);
xnor U1503 (N_1503,N_1269,N_1207);
and U1504 (N_1504,N_1275,N_1393);
and U1505 (N_1505,N_1206,N_1260);
or U1506 (N_1506,N_1376,N_1342);
nand U1507 (N_1507,N_1348,N_1293);
and U1508 (N_1508,N_1288,N_1343);
xnor U1509 (N_1509,N_1257,N_1373);
and U1510 (N_1510,N_1358,N_1245);
nand U1511 (N_1511,N_1343,N_1372);
nor U1512 (N_1512,N_1250,N_1361);
nor U1513 (N_1513,N_1316,N_1338);
or U1514 (N_1514,N_1292,N_1306);
or U1515 (N_1515,N_1336,N_1268);
or U1516 (N_1516,N_1245,N_1219);
xor U1517 (N_1517,N_1398,N_1259);
nand U1518 (N_1518,N_1355,N_1303);
nand U1519 (N_1519,N_1310,N_1364);
nand U1520 (N_1520,N_1228,N_1217);
and U1521 (N_1521,N_1313,N_1381);
xnor U1522 (N_1522,N_1322,N_1218);
nor U1523 (N_1523,N_1351,N_1267);
xnor U1524 (N_1524,N_1213,N_1370);
or U1525 (N_1525,N_1379,N_1389);
nand U1526 (N_1526,N_1263,N_1224);
xnor U1527 (N_1527,N_1201,N_1301);
nor U1528 (N_1528,N_1382,N_1212);
and U1529 (N_1529,N_1330,N_1240);
and U1530 (N_1530,N_1274,N_1322);
or U1531 (N_1531,N_1387,N_1268);
xnor U1532 (N_1532,N_1302,N_1260);
nor U1533 (N_1533,N_1273,N_1256);
or U1534 (N_1534,N_1303,N_1227);
xor U1535 (N_1535,N_1281,N_1200);
and U1536 (N_1536,N_1203,N_1315);
and U1537 (N_1537,N_1399,N_1307);
or U1538 (N_1538,N_1318,N_1337);
or U1539 (N_1539,N_1310,N_1313);
nor U1540 (N_1540,N_1312,N_1276);
xnor U1541 (N_1541,N_1273,N_1319);
and U1542 (N_1542,N_1250,N_1210);
and U1543 (N_1543,N_1240,N_1231);
nor U1544 (N_1544,N_1241,N_1243);
nand U1545 (N_1545,N_1256,N_1293);
or U1546 (N_1546,N_1229,N_1365);
nor U1547 (N_1547,N_1241,N_1289);
or U1548 (N_1548,N_1257,N_1275);
xnor U1549 (N_1549,N_1205,N_1326);
xor U1550 (N_1550,N_1284,N_1345);
nor U1551 (N_1551,N_1392,N_1360);
or U1552 (N_1552,N_1375,N_1229);
and U1553 (N_1553,N_1348,N_1217);
xor U1554 (N_1554,N_1372,N_1274);
or U1555 (N_1555,N_1236,N_1203);
nor U1556 (N_1556,N_1360,N_1377);
or U1557 (N_1557,N_1267,N_1377);
nand U1558 (N_1558,N_1213,N_1361);
nor U1559 (N_1559,N_1245,N_1238);
and U1560 (N_1560,N_1202,N_1257);
xor U1561 (N_1561,N_1252,N_1270);
and U1562 (N_1562,N_1328,N_1267);
nand U1563 (N_1563,N_1375,N_1393);
nand U1564 (N_1564,N_1318,N_1217);
or U1565 (N_1565,N_1214,N_1342);
nor U1566 (N_1566,N_1339,N_1208);
xor U1567 (N_1567,N_1394,N_1264);
nand U1568 (N_1568,N_1235,N_1286);
xor U1569 (N_1569,N_1290,N_1313);
and U1570 (N_1570,N_1331,N_1300);
xor U1571 (N_1571,N_1263,N_1235);
or U1572 (N_1572,N_1307,N_1326);
and U1573 (N_1573,N_1236,N_1391);
and U1574 (N_1574,N_1226,N_1280);
xor U1575 (N_1575,N_1333,N_1267);
or U1576 (N_1576,N_1384,N_1214);
or U1577 (N_1577,N_1254,N_1281);
nor U1578 (N_1578,N_1289,N_1263);
nor U1579 (N_1579,N_1274,N_1341);
and U1580 (N_1580,N_1202,N_1316);
nor U1581 (N_1581,N_1253,N_1323);
and U1582 (N_1582,N_1266,N_1267);
or U1583 (N_1583,N_1232,N_1356);
and U1584 (N_1584,N_1339,N_1238);
xor U1585 (N_1585,N_1394,N_1321);
and U1586 (N_1586,N_1345,N_1270);
and U1587 (N_1587,N_1361,N_1224);
nor U1588 (N_1588,N_1399,N_1324);
nor U1589 (N_1589,N_1268,N_1206);
or U1590 (N_1590,N_1343,N_1254);
xnor U1591 (N_1591,N_1398,N_1383);
xnor U1592 (N_1592,N_1382,N_1208);
xor U1593 (N_1593,N_1281,N_1306);
or U1594 (N_1594,N_1383,N_1312);
xor U1595 (N_1595,N_1266,N_1314);
or U1596 (N_1596,N_1253,N_1333);
nand U1597 (N_1597,N_1334,N_1225);
or U1598 (N_1598,N_1289,N_1313);
or U1599 (N_1599,N_1204,N_1242);
nand U1600 (N_1600,N_1565,N_1578);
nand U1601 (N_1601,N_1594,N_1439);
or U1602 (N_1602,N_1413,N_1417);
and U1603 (N_1603,N_1421,N_1472);
nor U1604 (N_1604,N_1525,N_1542);
or U1605 (N_1605,N_1489,N_1593);
or U1606 (N_1606,N_1552,N_1587);
and U1607 (N_1607,N_1474,N_1524);
xnor U1608 (N_1608,N_1546,N_1558);
nand U1609 (N_1609,N_1400,N_1501);
or U1610 (N_1610,N_1586,N_1547);
xor U1611 (N_1611,N_1584,N_1485);
or U1612 (N_1612,N_1479,N_1585);
nor U1613 (N_1613,N_1564,N_1486);
and U1614 (N_1614,N_1441,N_1581);
or U1615 (N_1615,N_1409,N_1466);
nand U1616 (N_1616,N_1462,N_1561);
xor U1617 (N_1617,N_1530,N_1495);
xnor U1618 (N_1618,N_1509,N_1595);
xnor U1619 (N_1619,N_1599,N_1438);
or U1620 (N_1620,N_1568,N_1478);
and U1621 (N_1621,N_1414,N_1433);
or U1622 (N_1622,N_1569,N_1492);
nand U1623 (N_1623,N_1420,N_1523);
xor U1624 (N_1624,N_1498,N_1536);
nand U1625 (N_1625,N_1480,N_1473);
or U1626 (N_1626,N_1511,N_1598);
and U1627 (N_1627,N_1502,N_1477);
and U1628 (N_1628,N_1447,N_1468);
nand U1629 (N_1629,N_1455,N_1482);
nand U1630 (N_1630,N_1562,N_1431);
or U1631 (N_1631,N_1465,N_1419);
and U1632 (N_1632,N_1460,N_1550);
nor U1633 (N_1633,N_1567,N_1458);
nand U1634 (N_1634,N_1582,N_1405);
or U1635 (N_1635,N_1583,N_1496);
xor U1636 (N_1636,N_1461,N_1519);
and U1637 (N_1637,N_1450,N_1463);
or U1638 (N_1638,N_1580,N_1505);
nor U1639 (N_1639,N_1516,N_1551);
xor U1640 (N_1640,N_1408,N_1481);
nand U1641 (N_1641,N_1576,N_1410);
xor U1642 (N_1642,N_1435,N_1402);
nand U1643 (N_1643,N_1467,N_1557);
and U1644 (N_1644,N_1437,N_1520);
nand U1645 (N_1645,N_1416,N_1573);
nor U1646 (N_1646,N_1436,N_1471);
nor U1647 (N_1647,N_1539,N_1488);
or U1648 (N_1648,N_1529,N_1574);
nand U1649 (N_1649,N_1434,N_1483);
nor U1650 (N_1650,N_1428,N_1588);
and U1651 (N_1651,N_1401,N_1545);
xor U1652 (N_1652,N_1544,N_1423);
nor U1653 (N_1653,N_1476,N_1560);
xnor U1654 (N_1654,N_1592,N_1540);
nor U1655 (N_1655,N_1493,N_1490);
xnor U1656 (N_1656,N_1521,N_1541);
or U1657 (N_1657,N_1532,N_1444);
nor U1658 (N_1658,N_1499,N_1445);
xor U1659 (N_1659,N_1448,N_1470);
and U1660 (N_1660,N_1548,N_1554);
and U1661 (N_1661,N_1589,N_1454);
xnor U1662 (N_1662,N_1559,N_1512);
nand U1663 (N_1663,N_1456,N_1407);
xor U1664 (N_1664,N_1526,N_1491);
nand U1665 (N_1665,N_1459,N_1534);
xor U1666 (N_1666,N_1570,N_1590);
nor U1667 (N_1667,N_1572,N_1591);
xor U1668 (N_1668,N_1555,N_1549);
and U1669 (N_1669,N_1411,N_1429);
or U1670 (N_1670,N_1571,N_1563);
nor U1671 (N_1671,N_1553,N_1537);
nand U1672 (N_1672,N_1504,N_1566);
nor U1673 (N_1673,N_1418,N_1517);
xor U1674 (N_1674,N_1475,N_1415);
and U1675 (N_1675,N_1507,N_1597);
and U1676 (N_1676,N_1531,N_1451);
nand U1677 (N_1677,N_1446,N_1443);
or U1678 (N_1678,N_1426,N_1440);
and U1679 (N_1679,N_1575,N_1457);
xor U1680 (N_1680,N_1533,N_1596);
or U1681 (N_1681,N_1464,N_1494);
xnor U1682 (N_1682,N_1403,N_1556);
nor U1683 (N_1683,N_1453,N_1500);
and U1684 (N_1684,N_1577,N_1449);
and U1685 (N_1685,N_1432,N_1510);
and U1686 (N_1686,N_1518,N_1412);
nand U1687 (N_1687,N_1497,N_1514);
nand U1688 (N_1688,N_1513,N_1487);
nor U1689 (N_1689,N_1430,N_1424);
nand U1690 (N_1690,N_1543,N_1484);
nor U1691 (N_1691,N_1528,N_1538);
or U1692 (N_1692,N_1425,N_1508);
and U1693 (N_1693,N_1503,N_1406);
xnor U1694 (N_1694,N_1527,N_1515);
or U1695 (N_1695,N_1506,N_1535);
nand U1696 (N_1696,N_1579,N_1469);
and U1697 (N_1697,N_1427,N_1422);
nor U1698 (N_1698,N_1404,N_1452);
xor U1699 (N_1699,N_1442,N_1522);
and U1700 (N_1700,N_1474,N_1550);
xor U1701 (N_1701,N_1509,N_1591);
nor U1702 (N_1702,N_1413,N_1567);
nor U1703 (N_1703,N_1577,N_1448);
nand U1704 (N_1704,N_1486,N_1465);
xnor U1705 (N_1705,N_1461,N_1492);
and U1706 (N_1706,N_1523,N_1434);
nor U1707 (N_1707,N_1516,N_1459);
xor U1708 (N_1708,N_1457,N_1553);
and U1709 (N_1709,N_1579,N_1545);
nand U1710 (N_1710,N_1519,N_1545);
or U1711 (N_1711,N_1473,N_1448);
nand U1712 (N_1712,N_1438,N_1524);
nor U1713 (N_1713,N_1571,N_1524);
or U1714 (N_1714,N_1527,N_1447);
and U1715 (N_1715,N_1461,N_1526);
nand U1716 (N_1716,N_1559,N_1492);
nor U1717 (N_1717,N_1429,N_1445);
xor U1718 (N_1718,N_1544,N_1515);
nand U1719 (N_1719,N_1454,N_1552);
and U1720 (N_1720,N_1565,N_1480);
and U1721 (N_1721,N_1423,N_1552);
or U1722 (N_1722,N_1413,N_1593);
xnor U1723 (N_1723,N_1597,N_1413);
or U1724 (N_1724,N_1506,N_1471);
and U1725 (N_1725,N_1481,N_1432);
or U1726 (N_1726,N_1522,N_1546);
nor U1727 (N_1727,N_1535,N_1538);
or U1728 (N_1728,N_1425,N_1465);
xor U1729 (N_1729,N_1586,N_1504);
nand U1730 (N_1730,N_1457,N_1545);
nand U1731 (N_1731,N_1472,N_1485);
and U1732 (N_1732,N_1481,N_1419);
xor U1733 (N_1733,N_1534,N_1520);
nand U1734 (N_1734,N_1578,N_1541);
xnor U1735 (N_1735,N_1429,N_1496);
and U1736 (N_1736,N_1411,N_1571);
nand U1737 (N_1737,N_1489,N_1493);
nor U1738 (N_1738,N_1502,N_1515);
nor U1739 (N_1739,N_1598,N_1505);
nor U1740 (N_1740,N_1521,N_1574);
xnor U1741 (N_1741,N_1420,N_1474);
nor U1742 (N_1742,N_1543,N_1514);
and U1743 (N_1743,N_1497,N_1587);
nand U1744 (N_1744,N_1582,N_1501);
xnor U1745 (N_1745,N_1449,N_1575);
nor U1746 (N_1746,N_1440,N_1442);
and U1747 (N_1747,N_1480,N_1518);
or U1748 (N_1748,N_1536,N_1407);
nor U1749 (N_1749,N_1489,N_1419);
nand U1750 (N_1750,N_1528,N_1559);
and U1751 (N_1751,N_1540,N_1466);
and U1752 (N_1752,N_1559,N_1459);
nand U1753 (N_1753,N_1582,N_1565);
nor U1754 (N_1754,N_1579,N_1555);
xor U1755 (N_1755,N_1473,N_1418);
nand U1756 (N_1756,N_1479,N_1417);
xor U1757 (N_1757,N_1572,N_1554);
or U1758 (N_1758,N_1547,N_1455);
nor U1759 (N_1759,N_1586,N_1451);
or U1760 (N_1760,N_1554,N_1510);
nor U1761 (N_1761,N_1561,N_1572);
nand U1762 (N_1762,N_1407,N_1481);
and U1763 (N_1763,N_1414,N_1459);
nand U1764 (N_1764,N_1595,N_1402);
or U1765 (N_1765,N_1496,N_1545);
and U1766 (N_1766,N_1401,N_1556);
and U1767 (N_1767,N_1535,N_1509);
and U1768 (N_1768,N_1431,N_1503);
nand U1769 (N_1769,N_1586,N_1571);
and U1770 (N_1770,N_1592,N_1470);
or U1771 (N_1771,N_1485,N_1531);
nand U1772 (N_1772,N_1511,N_1475);
and U1773 (N_1773,N_1463,N_1492);
nor U1774 (N_1774,N_1418,N_1458);
and U1775 (N_1775,N_1413,N_1466);
nand U1776 (N_1776,N_1432,N_1428);
or U1777 (N_1777,N_1592,N_1411);
and U1778 (N_1778,N_1571,N_1469);
or U1779 (N_1779,N_1496,N_1591);
or U1780 (N_1780,N_1483,N_1578);
xnor U1781 (N_1781,N_1562,N_1465);
xnor U1782 (N_1782,N_1542,N_1464);
xor U1783 (N_1783,N_1545,N_1422);
or U1784 (N_1784,N_1489,N_1578);
or U1785 (N_1785,N_1587,N_1565);
and U1786 (N_1786,N_1541,N_1450);
or U1787 (N_1787,N_1400,N_1472);
and U1788 (N_1788,N_1566,N_1489);
xor U1789 (N_1789,N_1409,N_1557);
and U1790 (N_1790,N_1546,N_1534);
or U1791 (N_1791,N_1423,N_1556);
or U1792 (N_1792,N_1511,N_1590);
or U1793 (N_1793,N_1416,N_1571);
and U1794 (N_1794,N_1400,N_1514);
and U1795 (N_1795,N_1531,N_1583);
nand U1796 (N_1796,N_1538,N_1492);
and U1797 (N_1797,N_1506,N_1524);
nand U1798 (N_1798,N_1527,N_1408);
nand U1799 (N_1799,N_1514,N_1499);
and U1800 (N_1800,N_1764,N_1603);
xnor U1801 (N_1801,N_1798,N_1792);
xnor U1802 (N_1802,N_1742,N_1775);
or U1803 (N_1803,N_1679,N_1674);
or U1804 (N_1804,N_1678,N_1776);
nor U1805 (N_1805,N_1602,N_1777);
and U1806 (N_1806,N_1624,N_1688);
or U1807 (N_1807,N_1715,N_1714);
nand U1808 (N_1808,N_1720,N_1628);
nor U1809 (N_1809,N_1605,N_1762);
nand U1810 (N_1810,N_1672,N_1658);
and U1811 (N_1811,N_1627,N_1645);
nand U1812 (N_1812,N_1657,N_1612);
xor U1813 (N_1813,N_1693,N_1640);
or U1814 (N_1814,N_1769,N_1621);
and U1815 (N_1815,N_1610,N_1699);
nor U1816 (N_1816,N_1730,N_1702);
xnor U1817 (N_1817,N_1726,N_1709);
xnor U1818 (N_1818,N_1751,N_1670);
and U1819 (N_1819,N_1689,N_1719);
nor U1820 (N_1820,N_1782,N_1634);
xnor U1821 (N_1821,N_1653,N_1647);
nor U1822 (N_1822,N_1677,N_1739);
nor U1823 (N_1823,N_1606,N_1607);
and U1824 (N_1824,N_1745,N_1698);
nor U1825 (N_1825,N_1660,N_1754);
and U1826 (N_1826,N_1744,N_1622);
nand U1827 (N_1827,N_1737,N_1664);
or U1828 (N_1828,N_1601,N_1700);
nor U1829 (N_1829,N_1789,N_1671);
nand U1830 (N_1830,N_1774,N_1799);
and U1831 (N_1831,N_1625,N_1747);
xnor U1832 (N_1832,N_1796,N_1659);
nand U1833 (N_1833,N_1649,N_1770);
xor U1834 (N_1834,N_1691,N_1680);
and U1835 (N_1835,N_1790,N_1686);
and U1836 (N_1836,N_1685,N_1692);
or U1837 (N_1837,N_1723,N_1633);
nor U1838 (N_1838,N_1760,N_1636);
nor U1839 (N_1839,N_1684,N_1614);
nand U1840 (N_1840,N_1787,N_1683);
or U1841 (N_1841,N_1718,N_1663);
xor U1842 (N_1842,N_1785,N_1611);
and U1843 (N_1843,N_1757,N_1665);
or U1844 (N_1844,N_1646,N_1741);
and U1845 (N_1845,N_1711,N_1701);
nand U1846 (N_1846,N_1766,N_1629);
nand U1847 (N_1847,N_1626,N_1619);
nor U1848 (N_1848,N_1681,N_1731);
and U1849 (N_1849,N_1673,N_1650);
nand U1850 (N_1850,N_1729,N_1662);
and U1851 (N_1851,N_1748,N_1779);
nand U1852 (N_1852,N_1716,N_1791);
xnor U1853 (N_1853,N_1758,N_1753);
xor U1854 (N_1854,N_1765,N_1604);
and U1855 (N_1855,N_1778,N_1661);
nor U1856 (N_1856,N_1797,N_1704);
xor U1857 (N_1857,N_1732,N_1793);
and U1858 (N_1858,N_1690,N_1608);
or U1859 (N_1859,N_1675,N_1786);
nand U1860 (N_1860,N_1752,N_1722);
and U1861 (N_1861,N_1727,N_1746);
or U1862 (N_1862,N_1721,N_1725);
nor U1863 (N_1863,N_1710,N_1713);
nand U1864 (N_1864,N_1697,N_1794);
nor U1865 (N_1865,N_1728,N_1617);
nand U1866 (N_1866,N_1620,N_1652);
or U1867 (N_1867,N_1687,N_1733);
nor U1868 (N_1868,N_1736,N_1638);
nand U1869 (N_1869,N_1717,N_1756);
nor U1870 (N_1870,N_1631,N_1767);
xnor U1871 (N_1871,N_1761,N_1784);
and U1872 (N_1872,N_1676,N_1771);
nor U1873 (N_1873,N_1648,N_1696);
xor U1874 (N_1874,N_1632,N_1668);
and U1875 (N_1875,N_1639,N_1695);
and U1876 (N_1876,N_1609,N_1763);
nand U1877 (N_1877,N_1705,N_1615);
or U1878 (N_1878,N_1616,N_1734);
and U1879 (N_1879,N_1750,N_1795);
nor U1880 (N_1880,N_1768,N_1735);
or U1881 (N_1881,N_1788,N_1759);
nor U1882 (N_1882,N_1740,N_1781);
xor U1883 (N_1883,N_1706,N_1637);
nor U1884 (N_1884,N_1635,N_1654);
and U1885 (N_1885,N_1707,N_1643);
nand U1886 (N_1886,N_1749,N_1682);
and U1887 (N_1887,N_1655,N_1667);
and U1888 (N_1888,N_1600,N_1724);
or U1889 (N_1889,N_1613,N_1755);
or U1890 (N_1890,N_1641,N_1669);
and U1891 (N_1891,N_1630,N_1642);
nand U1892 (N_1892,N_1666,N_1780);
nand U1893 (N_1893,N_1773,N_1694);
nor U1894 (N_1894,N_1703,N_1783);
or U1895 (N_1895,N_1644,N_1656);
nor U1896 (N_1896,N_1618,N_1712);
and U1897 (N_1897,N_1708,N_1743);
nand U1898 (N_1898,N_1623,N_1738);
xnor U1899 (N_1899,N_1651,N_1772);
or U1900 (N_1900,N_1787,N_1662);
nor U1901 (N_1901,N_1604,N_1618);
xnor U1902 (N_1902,N_1626,N_1752);
nor U1903 (N_1903,N_1635,N_1736);
or U1904 (N_1904,N_1700,N_1684);
nand U1905 (N_1905,N_1690,N_1785);
or U1906 (N_1906,N_1764,N_1628);
or U1907 (N_1907,N_1682,N_1742);
xor U1908 (N_1908,N_1688,N_1615);
or U1909 (N_1909,N_1742,N_1727);
nand U1910 (N_1910,N_1644,N_1705);
or U1911 (N_1911,N_1766,N_1718);
and U1912 (N_1912,N_1682,N_1743);
and U1913 (N_1913,N_1685,N_1760);
nor U1914 (N_1914,N_1795,N_1721);
and U1915 (N_1915,N_1678,N_1786);
nand U1916 (N_1916,N_1779,N_1662);
nor U1917 (N_1917,N_1706,N_1658);
xnor U1918 (N_1918,N_1673,N_1712);
and U1919 (N_1919,N_1764,N_1718);
nand U1920 (N_1920,N_1769,N_1788);
nor U1921 (N_1921,N_1771,N_1726);
and U1922 (N_1922,N_1600,N_1676);
nor U1923 (N_1923,N_1604,N_1721);
and U1924 (N_1924,N_1743,N_1613);
or U1925 (N_1925,N_1776,N_1653);
nand U1926 (N_1926,N_1632,N_1711);
and U1927 (N_1927,N_1653,N_1760);
and U1928 (N_1928,N_1799,N_1628);
nand U1929 (N_1929,N_1634,N_1650);
nand U1930 (N_1930,N_1780,N_1796);
nand U1931 (N_1931,N_1640,N_1739);
nand U1932 (N_1932,N_1693,N_1645);
nor U1933 (N_1933,N_1752,N_1727);
and U1934 (N_1934,N_1704,N_1691);
nor U1935 (N_1935,N_1657,N_1700);
or U1936 (N_1936,N_1619,N_1676);
and U1937 (N_1937,N_1793,N_1603);
and U1938 (N_1938,N_1698,N_1650);
and U1939 (N_1939,N_1668,N_1766);
or U1940 (N_1940,N_1793,N_1602);
xor U1941 (N_1941,N_1611,N_1745);
or U1942 (N_1942,N_1651,N_1751);
or U1943 (N_1943,N_1687,N_1677);
or U1944 (N_1944,N_1767,N_1634);
nor U1945 (N_1945,N_1706,N_1715);
nor U1946 (N_1946,N_1785,N_1773);
or U1947 (N_1947,N_1637,N_1786);
xnor U1948 (N_1948,N_1631,N_1648);
nand U1949 (N_1949,N_1761,N_1731);
xnor U1950 (N_1950,N_1720,N_1666);
nand U1951 (N_1951,N_1688,N_1646);
and U1952 (N_1952,N_1606,N_1652);
nand U1953 (N_1953,N_1703,N_1780);
nor U1954 (N_1954,N_1670,N_1608);
and U1955 (N_1955,N_1700,N_1608);
xor U1956 (N_1956,N_1719,N_1701);
nand U1957 (N_1957,N_1726,N_1723);
and U1958 (N_1958,N_1707,N_1718);
nor U1959 (N_1959,N_1665,N_1603);
and U1960 (N_1960,N_1771,N_1765);
or U1961 (N_1961,N_1622,N_1770);
nand U1962 (N_1962,N_1605,N_1688);
and U1963 (N_1963,N_1699,N_1773);
or U1964 (N_1964,N_1726,N_1716);
xnor U1965 (N_1965,N_1782,N_1709);
xor U1966 (N_1966,N_1632,N_1726);
nor U1967 (N_1967,N_1666,N_1636);
nor U1968 (N_1968,N_1771,N_1721);
xnor U1969 (N_1969,N_1790,N_1770);
nand U1970 (N_1970,N_1780,N_1635);
nand U1971 (N_1971,N_1774,N_1663);
nor U1972 (N_1972,N_1669,N_1654);
or U1973 (N_1973,N_1670,N_1754);
xnor U1974 (N_1974,N_1749,N_1759);
nand U1975 (N_1975,N_1720,N_1740);
nor U1976 (N_1976,N_1739,N_1703);
and U1977 (N_1977,N_1774,N_1717);
nand U1978 (N_1978,N_1764,N_1663);
and U1979 (N_1979,N_1649,N_1664);
or U1980 (N_1980,N_1772,N_1666);
nand U1981 (N_1981,N_1664,N_1692);
nor U1982 (N_1982,N_1631,N_1669);
xor U1983 (N_1983,N_1700,N_1654);
nand U1984 (N_1984,N_1752,N_1664);
xnor U1985 (N_1985,N_1719,N_1781);
xor U1986 (N_1986,N_1769,N_1781);
and U1987 (N_1987,N_1610,N_1650);
and U1988 (N_1988,N_1748,N_1600);
nand U1989 (N_1989,N_1642,N_1619);
nor U1990 (N_1990,N_1755,N_1705);
or U1991 (N_1991,N_1658,N_1630);
or U1992 (N_1992,N_1781,N_1611);
or U1993 (N_1993,N_1783,N_1644);
nor U1994 (N_1994,N_1711,N_1736);
or U1995 (N_1995,N_1708,N_1671);
nor U1996 (N_1996,N_1638,N_1716);
xnor U1997 (N_1997,N_1694,N_1772);
nor U1998 (N_1998,N_1689,N_1605);
nor U1999 (N_1999,N_1692,N_1607);
or U2000 (N_2000,N_1802,N_1975);
nand U2001 (N_2001,N_1835,N_1893);
nand U2002 (N_2002,N_1963,N_1988);
nor U2003 (N_2003,N_1932,N_1845);
nor U2004 (N_2004,N_1927,N_1926);
or U2005 (N_2005,N_1892,N_1933);
nor U2006 (N_2006,N_1951,N_1948);
and U2007 (N_2007,N_1969,N_1978);
nor U2008 (N_2008,N_1847,N_1928);
xor U2009 (N_2009,N_1889,N_1959);
nand U2010 (N_2010,N_1877,N_1849);
nand U2011 (N_2011,N_1878,N_1866);
xnor U2012 (N_2012,N_1905,N_1828);
or U2013 (N_2013,N_1834,N_1820);
or U2014 (N_2014,N_1996,N_1865);
nand U2015 (N_2015,N_1982,N_1950);
nor U2016 (N_2016,N_1929,N_1987);
nand U2017 (N_2017,N_1887,N_1954);
nand U2018 (N_2018,N_1995,N_1985);
nor U2019 (N_2019,N_1984,N_1962);
nor U2020 (N_2020,N_1943,N_1825);
nand U2021 (N_2021,N_1971,N_1821);
nor U2022 (N_2022,N_1871,N_1942);
nand U2023 (N_2023,N_1886,N_1851);
and U2024 (N_2024,N_1953,N_1961);
and U2025 (N_2025,N_1937,N_1890);
xnor U2026 (N_2026,N_1999,N_1966);
and U2027 (N_2027,N_1908,N_1850);
and U2028 (N_2028,N_1891,N_1980);
xnor U2029 (N_2029,N_1819,N_1918);
and U2030 (N_2030,N_1842,N_1884);
nand U2031 (N_2031,N_1867,N_1925);
nand U2032 (N_2032,N_1843,N_1860);
or U2033 (N_2033,N_1862,N_1917);
nand U2034 (N_2034,N_1822,N_1832);
or U2035 (N_2035,N_1903,N_1906);
or U2036 (N_2036,N_1855,N_1934);
nand U2037 (N_2037,N_1976,N_1883);
nand U2038 (N_2038,N_1874,N_1900);
and U2039 (N_2039,N_1946,N_1808);
or U2040 (N_2040,N_1854,N_1936);
xnor U2041 (N_2041,N_1840,N_1833);
and U2042 (N_2042,N_1970,N_1997);
and U2043 (N_2043,N_1881,N_1872);
nand U2044 (N_2044,N_1967,N_1979);
nor U2045 (N_2045,N_1896,N_1879);
and U2046 (N_2046,N_1931,N_1955);
and U2047 (N_2047,N_1801,N_1809);
and U2048 (N_2048,N_1880,N_1895);
xor U2049 (N_2049,N_1869,N_1814);
nand U2050 (N_2050,N_1923,N_1816);
xnor U2051 (N_2051,N_1977,N_1910);
or U2052 (N_2052,N_1810,N_1993);
nand U2053 (N_2053,N_1817,N_1804);
xnor U2054 (N_2054,N_1830,N_1813);
nand U2055 (N_2055,N_1807,N_1841);
nand U2056 (N_2056,N_1897,N_1812);
xnor U2057 (N_2057,N_1998,N_1852);
nand U2058 (N_2058,N_1914,N_1912);
nand U2059 (N_2059,N_1831,N_1829);
or U2060 (N_2060,N_1894,N_1968);
xor U2061 (N_2061,N_1864,N_1972);
or U2062 (N_2062,N_1838,N_1935);
and U2063 (N_2063,N_1940,N_1876);
nor U2064 (N_2064,N_1882,N_1858);
or U2065 (N_2065,N_1919,N_1960);
or U2066 (N_2066,N_1921,N_1992);
nand U2067 (N_2067,N_1989,N_1907);
nor U2068 (N_2068,N_1949,N_1837);
xnor U2069 (N_2069,N_1957,N_1899);
and U2070 (N_2070,N_1856,N_1965);
nor U2071 (N_2071,N_1916,N_1904);
nor U2072 (N_2072,N_1956,N_1991);
nand U2073 (N_2073,N_1815,N_1836);
nor U2074 (N_2074,N_1915,N_1875);
nor U2075 (N_2075,N_1857,N_1939);
xnor U2076 (N_2076,N_1973,N_1994);
nand U2077 (N_2077,N_1848,N_1888);
nand U2078 (N_2078,N_1938,N_1922);
and U2079 (N_2079,N_1974,N_1909);
xnor U2080 (N_2080,N_1870,N_1827);
or U2081 (N_2081,N_1898,N_1902);
and U2082 (N_2082,N_1806,N_1885);
or U2083 (N_2083,N_1944,N_1800);
nand U2084 (N_2084,N_1868,N_1853);
and U2085 (N_2085,N_1986,N_1844);
and U2086 (N_2086,N_1818,N_1947);
xor U2087 (N_2087,N_1981,N_1824);
and U2088 (N_2088,N_1913,N_1805);
or U2089 (N_2089,N_1861,N_1911);
xor U2090 (N_2090,N_1873,N_1826);
nand U2091 (N_2091,N_1924,N_1823);
nand U2092 (N_2092,N_1930,N_1859);
nand U2093 (N_2093,N_1952,N_1920);
nand U2094 (N_2094,N_1863,N_1990);
xor U2095 (N_2095,N_1846,N_1803);
xor U2096 (N_2096,N_1945,N_1839);
or U2097 (N_2097,N_1958,N_1811);
nand U2098 (N_2098,N_1964,N_1941);
nor U2099 (N_2099,N_1901,N_1983);
nand U2100 (N_2100,N_1818,N_1915);
nor U2101 (N_2101,N_1976,N_1845);
nor U2102 (N_2102,N_1896,N_1831);
and U2103 (N_2103,N_1882,N_1908);
xnor U2104 (N_2104,N_1827,N_1835);
or U2105 (N_2105,N_1814,N_1866);
and U2106 (N_2106,N_1827,N_1831);
xor U2107 (N_2107,N_1935,N_1978);
or U2108 (N_2108,N_1990,N_1819);
xor U2109 (N_2109,N_1981,N_1879);
xor U2110 (N_2110,N_1938,N_1874);
or U2111 (N_2111,N_1888,N_1845);
nor U2112 (N_2112,N_1996,N_1890);
or U2113 (N_2113,N_1978,N_1812);
or U2114 (N_2114,N_1913,N_1861);
and U2115 (N_2115,N_1869,N_1948);
nand U2116 (N_2116,N_1897,N_1817);
xnor U2117 (N_2117,N_1943,N_1901);
xnor U2118 (N_2118,N_1936,N_1972);
and U2119 (N_2119,N_1980,N_1947);
and U2120 (N_2120,N_1948,N_1922);
or U2121 (N_2121,N_1963,N_1946);
xnor U2122 (N_2122,N_1978,N_1894);
nor U2123 (N_2123,N_1958,N_1875);
or U2124 (N_2124,N_1962,N_1865);
nor U2125 (N_2125,N_1836,N_1816);
xnor U2126 (N_2126,N_1896,N_1966);
or U2127 (N_2127,N_1885,N_1914);
or U2128 (N_2128,N_1848,N_1951);
nand U2129 (N_2129,N_1966,N_1854);
and U2130 (N_2130,N_1853,N_1962);
and U2131 (N_2131,N_1852,N_1963);
and U2132 (N_2132,N_1800,N_1834);
nand U2133 (N_2133,N_1898,N_1823);
nand U2134 (N_2134,N_1904,N_1961);
and U2135 (N_2135,N_1995,N_1847);
and U2136 (N_2136,N_1934,N_1868);
and U2137 (N_2137,N_1962,N_1876);
and U2138 (N_2138,N_1876,N_1968);
nor U2139 (N_2139,N_1836,N_1970);
xnor U2140 (N_2140,N_1967,N_1888);
nor U2141 (N_2141,N_1905,N_1823);
xnor U2142 (N_2142,N_1889,N_1926);
and U2143 (N_2143,N_1841,N_1889);
xnor U2144 (N_2144,N_1844,N_1943);
nand U2145 (N_2145,N_1924,N_1875);
nand U2146 (N_2146,N_1937,N_1805);
nor U2147 (N_2147,N_1907,N_1863);
nor U2148 (N_2148,N_1870,N_1832);
nand U2149 (N_2149,N_1998,N_1910);
or U2150 (N_2150,N_1957,N_1927);
nor U2151 (N_2151,N_1952,N_1841);
xor U2152 (N_2152,N_1842,N_1893);
and U2153 (N_2153,N_1873,N_1978);
xnor U2154 (N_2154,N_1934,N_1846);
xnor U2155 (N_2155,N_1970,N_1960);
and U2156 (N_2156,N_1855,N_1876);
nor U2157 (N_2157,N_1939,N_1942);
xor U2158 (N_2158,N_1865,N_1909);
xor U2159 (N_2159,N_1837,N_1879);
nor U2160 (N_2160,N_1823,N_1878);
nor U2161 (N_2161,N_1858,N_1804);
nand U2162 (N_2162,N_1802,N_1845);
nand U2163 (N_2163,N_1820,N_1880);
nor U2164 (N_2164,N_1858,N_1911);
nor U2165 (N_2165,N_1981,N_1848);
xor U2166 (N_2166,N_1999,N_1862);
nor U2167 (N_2167,N_1944,N_1857);
nor U2168 (N_2168,N_1945,N_1878);
and U2169 (N_2169,N_1956,N_1839);
or U2170 (N_2170,N_1916,N_1888);
nand U2171 (N_2171,N_1942,N_1902);
nand U2172 (N_2172,N_1821,N_1843);
nand U2173 (N_2173,N_1815,N_1990);
nand U2174 (N_2174,N_1898,N_1961);
nand U2175 (N_2175,N_1901,N_1860);
and U2176 (N_2176,N_1998,N_1927);
and U2177 (N_2177,N_1935,N_1915);
or U2178 (N_2178,N_1834,N_1959);
nand U2179 (N_2179,N_1866,N_1946);
nor U2180 (N_2180,N_1990,N_1932);
and U2181 (N_2181,N_1991,N_1960);
or U2182 (N_2182,N_1938,N_1856);
and U2183 (N_2183,N_1801,N_1938);
nand U2184 (N_2184,N_1817,N_1986);
and U2185 (N_2185,N_1898,N_1892);
or U2186 (N_2186,N_1820,N_1836);
nand U2187 (N_2187,N_1838,N_1885);
nand U2188 (N_2188,N_1860,N_1983);
xnor U2189 (N_2189,N_1997,N_1822);
xnor U2190 (N_2190,N_1881,N_1819);
nand U2191 (N_2191,N_1921,N_1908);
nand U2192 (N_2192,N_1913,N_1953);
and U2193 (N_2193,N_1883,N_1825);
or U2194 (N_2194,N_1858,N_1929);
nand U2195 (N_2195,N_1952,N_1929);
nand U2196 (N_2196,N_1861,N_1925);
nand U2197 (N_2197,N_1972,N_1907);
or U2198 (N_2198,N_1837,N_1870);
xor U2199 (N_2199,N_1937,N_1830);
or U2200 (N_2200,N_2055,N_2083);
nand U2201 (N_2201,N_2141,N_2198);
nor U2202 (N_2202,N_2041,N_2170);
xor U2203 (N_2203,N_2163,N_2032);
nand U2204 (N_2204,N_2002,N_2082);
xnor U2205 (N_2205,N_2023,N_2169);
nor U2206 (N_2206,N_2124,N_2053);
nand U2207 (N_2207,N_2021,N_2061);
xnor U2208 (N_2208,N_2133,N_2167);
xnor U2209 (N_2209,N_2050,N_2152);
xor U2210 (N_2210,N_2146,N_2057);
xnor U2211 (N_2211,N_2038,N_2070);
and U2212 (N_2212,N_2001,N_2086);
and U2213 (N_2213,N_2175,N_2077);
and U2214 (N_2214,N_2197,N_2068);
nor U2215 (N_2215,N_2059,N_2158);
nor U2216 (N_2216,N_2111,N_2015);
nand U2217 (N_2217,N_2026,N_2044);
xnor U2218 (N_2218,N_2101,N_2119);
xor U2219 (N_2219,N_2052,N_2143);
nand U2220 (N_2220,N_2154,N_2145);
or U2221 (N_2221,N_2153,N_2110);
and U2222 (N_2222,N_2131,N_2007);
and U2223 (N_2223,N_2012,N_2132);
nand U2224 (N_2224,N_2172,N_2051);
xnor U2225 (N_2225,N_2065,N_2164);
nand U2226 (N_2226,N_2004,N_2165);
nor U2227 (N_2227,N_2099,N_2171);
or U2228 (N_2228,N_2076,N_2089);
xor U2229 (N_2229,N_2036,N_2104);
and U2230 (N_2230,N_2182,N_2107);
nand U2231 (N_2231,N_2011,N_2162);
and U2232 (N_2232,N_2192,N_2116);
nand U2233 (N_2233,N_2195,N_2122);
xor U2234 (N_2234,N_2029,N_2084);
or U2235 (N_2235,N_2034,N_2081);
or U2236 (N_2236,N_2128,N_2048);
nand U2237 (N_2237,N_2114,N_2039);
nor U2238 (N_2238,N_2037,N_2091);
nand U2239 (N_2239,N_2071,N_2121);
nand U2240 (N_2240,N_2137,N_2060);
and U2241 (N_2241,N_2017,N_2035);
nand U2242 (N_2242,N_2100,N_2063);
xor U2243 (N_2243,N_2073,N_2180);
and U2244 (N_2244,N_2043,N_2087);
nand U2245 (N_2245,N_2189,N_2160);
or U2246 (N_2246,N_2097,N_2148);
nand U2247 (N_2247,N_2138,N_2078);
xnor U2248 (N_2248,N_2109,N_2126);
and U2249 (N_2249,N_2115,N_2067);
nand U2250 (N_2250,N_2177,N_2058);
or U2251 (N_2251,N_2150,N_2009);
and U2252 (N_2252,N_2056,N_2022);
and U2253 (N_2253,N_2120,N_2066);
nand U2254 (N_2254,N_2005,N_2003);
xor U2255 (N_2255,N_2016,N_2129);
and U2256 (N_2256,N_2117,N_2147);
nand U2257 (N_2257,N_2174,N_2185);
or U2258 (N_2258,N_2040,N_2157);
nor U2259 (N_2259,N_2062,N_2045);
nand U2260 (N_2260,N_2049,N_2173);
and U2261 (N_2261,N_2139,N_2074);
nor U2262 (N_2262,N_2151,N_2064);
nand U2263 (N_2263,N_2008,N_2191);
and U2264 (N_2264,N_2024,N_2176);
and U2265 (N_2265,N_2127,N_2098);
or U2266 (N_2266,N_2149,N_2069);
and U2267 (N_2267,N_2006,N_2010);
nor U2268 (N_2268,N_2135,N_2075);
nand U2269 (N_2269,N_2108,N_2161);
nand U2270 (N_2270,N_2095,N_2168);
or U2271 (N_2271,N_2125,N_2144);
or U2272 (N_2272,N_2103,N_2027);
xor U2273 (N_2273,N_2106,N_2030);
and U2274 (N_2274,N_2018,N_2196);
xor U2275 (N_2275,N_2080,N_2014);
nor U2276 (N_2276,N_2019,N_2092);
xnor U2277 (N_2277,N_2047,N_2042);
nor U2278 (N_2278,N_2166,N_2085);
nor U2279 (N_2279,N_2088,N_2184);
and U2280 (N_2280,N_2020,N_2186);
and U2281 (N_2281,N_2102,N_2178);
nor U2282 (N_2282,N_2046,N_2025);
xnor U2283 (N_2283,N_2013,N_2136);
and U2284 (N_2284,N_2190,N_2199);
nor U2285 (N_2285,N_2031,N_2033);
and U2286 (N_2286,N_2118,N_2194);
and U2287 (N_2287,N_2181,N_2000);
nor U2288 (N_2288,N_2140,N_2096);
or U2289 (N_2289,N_2130,N_2179);
or U2290 (N_2290,N_2142,N_2079);
nand U2291 (N_2291,N_2156,N_2054);
or U2292 (N_2292,N_2134,N_2105);
xor U2293 (N_2293,N_2028,N_2112);
xor U2294 (N_2294,N_2093,N_2094);
and U2295 (N_2295,N_2155,N_2123);
or U2296 (N_2296,N_2113,N_2072);
xnor U2297 (N_2297,N_2183,N_2159);
and U2298 (N_2298,N_2188,N_2187);
nor U2299 (N_2299,N_2193,N_2090);
nor U2300 (N_2300,N_2159,N_2106);
or U2301 (N_2301,N_2002,N_2034);
nor U2302 (N_2302,N_2038,N_2108);
and U2303 (N_2303,N_2025,N_2032);
or U2304 (N_2304,N_2033,N_2168);
or U2305 (N_2305,N_2112,N_2077);
and U2306 (N_2306,N_2087,N_2003);
nor U2307 (N_2307,N_2067,N_2074);
xnor U2308 (N_2308,N_2028,N_2037);
nand U2309 (N_2309,N_2153,N_2175);
xor U2310 (N_2310,N_2195,N_2073);
xnor U2311 (N_2311,N_2181,N_2180);
or U2312 (N_2312,N_2075,N_2086);
or U2313 (N_2313,N_2025,N_2178);
nor U2314 (N_2314,N_2110,N_2086);
nor U2315 (N_2315,N_2056,N_2115);
or U2316 (N_2316,N_2185,N_2083);
and U2317 (N_2317,N_2069,N_2099);
or U2318 (N_2318,N_2137,N_2075);
and U2319 (N_2319,N_2091,N_2198);
xor U2320 (N_2320,N_2070,N_2190);
or U2321 (N_2321,N_2189,N_2102);
or U2322 (N_2322,N_2132,N_2016);
xnor U2323 (N_2323,N_2136,N_2037);
and U2324 (N_2324,N_2095,N_2118);
nand U2325 (N_2325,N_2111,N_2002);
or U2326 (N_2326,N_2021,N_2185);
or U2327 (N_2327,N_2137,N_2013);
and U2328 (N_2328,N_2126,N_2115);
nand U2329 (N_2329,N_2086,N_2005);
nand U2330 (N_2330,N_2073,N_2021);
xor U2331 (N_2331,N_2102,N_2162);
and U2332 (N_2332,N_2137,N_2126);
xnor U2333 (N_2333,N_2064,N_2133);
xnor U2334 (N_2334,N_2070,N_2110);
xnor U2335 (N_2335,N_2126,N_2021);
xor U2336 (N_2336,N_2128,N_2041);
xnor U2337 (N_2337,N_2116,N_2094);
and U2338 (N_2338,N_2138,N_2021);
and U2339 (N_2339,N_2083,N_2183);
nand U2340 (N_2340,N_2158,N_2181);
nor U2341 (N_2341,N_2156,N_2157);
or U2342 (N_2342,N_2121,N_2078);
nand U2343 (N_2343,N_2146,N_2051);
nand U2344 (N_2344,N_2109,N_2148);
xor U2345 (N_2345,N_2060,N_2133);
xor U2346 (N_2346,N_2053,N_2168);
xnor U2347 (N_2347,N_2183,N_2111);
nor U2348 (N_2348,N_2003,N_2019);
nor U2349 (N_2349,N_2006,N_2025);
xor U2350 (N_2350,N_2062,N_2152);
nor U2351 (N_2351,N_2018,N_2126);
xnor U2352 (N_2352,N_2137,N_2182);
nor U2353 (N_2353,N_2159,N_2130);
xor U2354 (N_2354,N_2180,N_2144);
nor U2355 (N_2355,N_2109,N_2073);
nand U2356 (N_2356,N_2101,N_2076);
and U2357 (N_2357,N_2098,N_2010);
nand U2358 (N_2358,N_2005,N_2144);
xor U2359 (N_2359,N_2150,N_2148);
xor U2360 (N_2360,N_2036,N_2052);
nor U2361 (N_2361,N_2082,N_2133);
and U2362 (N_2362,N_2095,N_2159);
nand U2363 (N_2363,N_2086,N_2057);
xor U2364 (N_2364,N_2059,N_2019);
and U2365 (N_2365,N_2000,N_2051);
and U2366 (N_2366,N_2143,N_2156);
and U2367 (N_2367,N_2138,N_2032);
nor U2368 (N_2368,N_2044,N_2111);
or U2369 (N_2369,N_2172,N_2067);
and U2370 (N_2370,N_2107,N_2112);
nor U2371 (N_2371,N_2077,N_2189);
xor U2372 (N_2372,N_2046,N_2198);
xor U2373 (N_2373,N_2143,N_2037);
nand U2374 (N_2374,N_2024,N_2069);
nand U2375 (N_2375,N_2187,N_2086);
nand U2376 (N_2376,N_2062,N_2028);
nor U2377 (N_2377,N_2092,N_2173);
xor U2378 (N_2378,N_2139,N_2183);
and U2379 (N_2379,N_2183,N_2100);
and U2380 (N_2380,N_2030,N_2154);
xnor U2381 (N_2381,N_2199,N_2001);
xnor U2382 (N_2382,N_2050,N_2114);
and U2383 (N_2383,N_2142,N_2003);
and U2384 (N_2384,N_2037,N_2057);
nor U2385 (N_2385,N_2137,N_2035);
nand U2386 (N_2386,N_2037,N_2140);
and U2387 (N_2387,N_2159,N_2009);
and U2388 (N_2388,N_2135,N_2034);
xor U2389 (N_2389,N_2164,N_2111);
nor U2390 (N_2390,N_2062,N_2190);
nand U2391 (N_2391,N_2192,N_2018);
and U2392 (N_2392,N_2004,N_2162);
and U2393 (N_2393,N_2021,N_2063);
and U2394 (N_2394,N_2180,N_2063);
xor U2395 (N_2395,N_2140,N_2024);
and U2396 (N_2396,N_2196,N_2197);
xnor U2397 (N_2397,N_2001,N_2055);
or U2398 (N_2398,N_2145,N_2156);
nor U2399 (N_2399,N_2088,N_2161);
nand U2400 (N_2400,N_2335,N_2391);
xor U2401 (N_2401,N_2392,N_2217);
nor U2402 (N_2402,N_2272,N_2252);
nor U2403 (N_2403,N_2316,N_2220);
nor U2404 (N_2404,N_2326,N_2204);
nand U2405 (N_2405,N_2228,N_2355);
nor U2406 (N_2406,N_2352,N_2322);
nor U2407 (N_2407,N_2236,N_2376);
and U2408 (N_2408,N_2334,N_2203);
or U2409 (N_2409,N_2264,N_2336);
nor U2410 (N_2410,N_2240,N_2311);
nor U2411 (N_2411,N_2246,N_2370);
nor U2412 (N_2412,N_2274,N_2296);
or U2413 (N_2413,N_2314,N_2259);
and U2414 (N_2414,N_2306,N_2202);
and U2415 (N_2415,N_2292,N_2289);
xor U2416 (N_2416,N_2249,N_2210);
nand U2417 (N_2417,N_2318,N_2364);
xor U2418 (N_2418,N_2271,N_2331);
nor U2419 (N_2419,N_2341,N_2347);
nand U2420 (N_2420,N_2389,N_2224);
xnor U2421 (N_2421,N_2382,N_2215);
or U2422 (N_2422,N_2221,N_2354);
nand U2423 (N_2423,N_2283,N_2241);
or U2424 (N_2424,N_2287,N_2398);
or U2425 (N_2425,N_2397,N_2396);
nor U2426 (N_2426,N_2328,N_2369);
xnor U2427 (N_2427,N_2363,N_2325);
xor U2428 (N_2428,N_2226,N_2386);
and U2429 (N_2429,N_2279,N_2375);
nand U2430 (N_2430,N_2394,N_2372);
nor U2431 (N_2431,N_2267,N_2214);
or U2432 (N_2432,N_2356,N_2270);
xor U2433 (N_2433,N_2309,N_2348);
nor U2434 (N_2434,N_2345,N_2294);
nor U2435 (N_2435,N_2346,N_2280);
xor U2436 (N_2436,N_2303,N_2254);
xor U2437 (N_2437,N_2317,N_2366);
or U2438 (N_2438,N_2388,N_2358);
nor U2439 (N_2439,N_2208,N_2213);
xor U2440 (N_2440,N_2349,N_2378);
nand U2441 (N_2441,N_2269,N_2298);
or U2442 (N_2442,N_2357,N_2248);
xor U2443 (N_2443,N_2247,N_2360);
and U2444 (N_2444,N_2205,N_2286);
nor U2445 (N_2445,N_2302,N_2351);
xnor U2446 (N_2446,N_2327,N_2290);
nand U2447 (N_2447,N_2321,N_2277);
and U2448 (N_2448,N_2231,N_2230);
xnor U2449 (N_2449,N_2380,N_2340);
and U2450 (N_2450,N_2381,N_2361);
xor U2451 (N_2451,N_2206,N_2333);
or U2452 (N_2452,N_2374,N_2332);
xor U2453 (N_2453,N_2219,N_2265);
xnor U2454 (N_2454,N_2233,N_2330);
or U2455 (N_2455,N_2385,N_2201);
or U2456 (N_2456,N_2211,N_2266);
xor U2457 (N_2457,N_2310,N_2212);
or U2458 (N_2458,N_2229,N_2207);
and U2459 (N_2459,N_2305,N_2281);
nor U2460 (N_2460,N_2373,N_2261);
nor U2461 (N_2461,N_2238,N_2342);
nor U2462 (N_2462,N_2218,N_2390);
and U2463 (N_2463,N_2239,N_2242);
nand U2464 (N_2464,N_2350,N_2216);
xor U2465 (N_2465,N_2209,N_2234);
and U2466 (N_2466,N_2320,N_2288);
nor U2467 (N_2467,N_2395,N_2227);
xor U2468 (N_2468,N_2295,N_2256);
or U2469 (N_2469,N_2243,N_2235);
and U2470 (N_2470,N_2368,N_2225);
xor U2471 (N_2471,N_2285,N_2275);
or U2472 (N_2472,N_2237,N_2338);
and U2473 (N_2473,N_2251,N_2387);
nand U2474 (N_2474,N_2308,N_2324);
or U2475 (N_2475,N_2313,N_2276);
nand U2476 (N_2476,N_2323,N_2268);
nand U2477 (N_2477,N_2293,N_2371);
or U2478 (N_2478,N_2367,N_2278);
nor U2479 (N_2479,N_2223,N_2255);
xnor U2480 (N_2480,N_2260,N_2245);
and U2481 (N_2481,N_2377,N_2300);
xor U2482 (N_2482,N_2258,N_2257);
or U2483 (N_2483,N_2262,N_2304);
and U2484 (N_2484,N_2299,N_2315);
or U2485 (N_2485,N_2273,N_2284);
nand U2486 (N_2486,N_2344,N_2362);
nor U2487 (N_2487,N_2339,N_2383);
or U2488 (N_2488,N_2222,N_2263);
nand U2489 (N_2489,N_2319,N_2312);
nor U2490 (N_2490,N_2253,N_2343);
nor U2491 (N_2491,N_2365,N_2282);
or U2492 (N_2492,N_2359,N_2399);
nor U2493 (N_2493,N_2337,N_2384);
or U2494 (N_2494,N_2353,N_2393);
nor U2495 (N_2495,N_2329,N_2250);
nand U2496 (N_2496,N_2200,N_2291);
xnor U2497 (N_2497,N_2301,N_2379);
xnor U2498 (N_2498,N_2297,N_2232);
xor U2499 (N_2499,N_2307,N_2244);
xnor U2500 (N_2500,N_2256,N_2246);
and U2501 (N_2501,N_2311,N_2239);
or U2502 (N_2502,N_2248,N_2207);
nand U2503 (N_2503,N_2386,N_2352);
xor U2504 (N_2504,N_2253,N_2339);
xnor U2505 (N_2505,N_2226,N_2284);
and U2506 (N_2506,N_2375,N_2260);
and U2507 (N_2507,N_2319,N_2344);
nand U2508 (N_2508,N_2395,N_2295);
or U2509 (N_2509,N_2370,N_2317);
xor U2510 (N_2510,N_2217,N_2275);
xnor U2511 (N_2511,N_2220,N_2300);
xnor U2512 (N_2512,N_2289,N_2280);
and U2513 (N_2513,N_2371,N_2358);
xnor U2514 (N_2514,N_2270,N_2316);
or U2515 (N_2515,N_2388,N_2314);
xnor U2516 (N_2516,N_2222,N_2364);
xor U2517 (N_2517,N_2266,N_2344);
nand U2518 (N_2518,N_2201,N_2277);
nor U2519 (N_2519,N_2302,N_2263);
xor U2520 (N_2520,N_2277,N_2213);
and U2521 (N_2521,N_2215,N_2340);
and U2522 (N_2522,N_2249,N_2203);
and U2523 (N_2523,N_2279,N_2311);
xor U2524 (N_2524,N_2261,N_2213);
nand U2525 (N_2525,N_2241,N_2313);
and U2526 (N_2526,N_2254,N_2292);
or U2527 (N_2527,N_2293,N_2365);
nand U2528 (N_2528,N_2248,N_2225);
nor U2529 (N_2529,N_2342,N_2216);
or U2530 (N_2530,N_2310,N_2379);
and U2531 (N_2531,N_2251,N_2224);
and U2532 (N_2532,N_2334,N_2345);
and U2533 (N_2533,N_2235,N_2372);
nand U2534 (N_2534,N_2263,N_2280);
nor U2535 (N_2535,N_2231,N_2366);
or U2536 (N_2536,N_2314,N_2264);
xor U2537 (N_2537,N_2316,N_2213);
nand U2538 (N_2538,N_2379,N_2242);
and U2539 (N_2539,N_2342,N_2256);
xor U2540 (N_2540,N_2356,N_2341);
xnor U2541 (N_2541,N_2307,N_2257);
xor U2542 (N_2542,N_2201,N_2203);
xor U2543 (N_2543,N_2202,N_2341);
nor U2544 (N_2544,N_2205,N_2325);
xor U2545 (N_2545,N_2300,N_2272);
and U2546 (N_2546,N_2294,N_2329);
nand U2547 (N_2547,N_2202,N_2258);
and U2548 (N_2548,N_2235,N_2210);
nand U2549 (N_2549,N_2205,N_2203);
nand U2550 (N_2550,N_2320,N_2214);
or U2551 (N_2551,N_2231,N_2305);
nor U2552 (N_2552,N_2341,N_2216);
and U2553 (N_2553,N_2273,N_2335);
nor U2554 (N_2554,N_2278,N_2380);
nand U2555 (N_2555,N_2296,N_2254);
nor U2556 (N_2556,N_2282,N_2301);
or U2557 (N_2557,N_2211,N_2342);
and U2558 (N_2558,N_2280,N_2304);
or U2559 (N_2559,N_2332,N_2397);
nand U2560 (N_2560,N_2378,N_2331);
nor U2561 (N_2561,N_2216,N_2234);
and U2562 (N_2562,N_2235,N_2274);
nand U2563 (N_2563,N_2208,N_2375);
nand U2564 (N_2564,N_2273,N_2334);
or U2565 (N_2565,N_2334,N_2201);
nand U2566 (N_2566,N_2297,N_2380);
xnor U2567 (N_2567,N_2363,N_2257);
nand U2568 (N_2568,N_2224,N_2222);
xnor U2569 (N_2569,N_2217,N_2221);
or U2570 (N_2570,N_2216,N_2224);
or U2571 (N_2571,N_2243,N_2334);
and U2572 (N_2572,N_2220,N_2211);
or U2573 (N_2573,N_2316,N_2286);
or U2574 (N_2574,N_2395,N_2289);
xor U2575 (N_2575,N_2314,N_2201);
and U2576 (N_2576,N_2363,N_2367);
or U2577 (N_2577,N_2366,N_2341);
nand U2578 (N_2578,N_2209,N_2273);
nor U2579 (N_2579,N_2365,N_2393);
or U2580 (N_2580,N_2368,N_2286);
xnor U2581 (N_2581,N_2230,N_2224);
xor U2582 (N_2582,N_2204,N_2372);
nor U2583 (N_2583,N_2211,N_2226);
nand U2584 (N_2584,N_2345,N_2288);
or U2585 (N_2585,N_2351,N_2288);
nand U2586 (N_2586,N_2206,N_2205);
and U2587 (N_2587,N_2258,N_2327);
and U2588 (N_2588,N_2248,N_2208);
xnor U2589 (N_2589,N_2385,N_2231);
nand U2590 (N_2590,N_2208,N_2239);
nand U2591 (N_2591,N_2382,N_2228);
xnor U2592 (N_2592,N_2373,N_2298);
xor U2593 (N_2593,N_2307,N_2374);
nand U2594 (N_2594,N_2364,N_2250);
xor U2595 (N_2595,N_2329,N_2378);
and U2596 (N_2596,N_2393,N_2311);
and U2597 (N_2597,N_2394,N_2293);
or U2598 (N_2598,N_2349,N_2268);
nand U2599 (N_2599,N_2213,N_2231);
xnor U2600 (N_2600,N_2530,N_2456);
nand U2601 (N_2601,N_2413,N_2415);
or U2602 (N_2602,N_2560,N_2444);
nor U2603 (N_2603,N_2419,N_2402);
nor U2604 (N_2604,N_2541,N_2578);
nand U2605 (N_2605,N_2513,N_2511);
and U2606 (N_2606,N_2490,N_2499);
or U2607 (N_2607,N_2549,N_2569);
xor U2608 (N_2608,N_2586,N_2590);
nor U2609 (N_2609,N_2567,N_2529);
and U2610 (N_2610,N_2571,N_2598);
nand U2611 (N_2611,N_2426,N_2485);
and U2612 (N_2612,N_2554,N_2409);
xnor U2613 (N_2613,N_2400,N_2583);
xnor U2614 (N_2614,N_2568,N_2498);
nand U2615 (N_2615,N_2538,N_2421);
or U2616 (N_2616,N_2469,N_2570);
xor U2617 (N_2617,N_2536,N_2446);
nand U2618 (N_2618,N_2540,N_2427);
or U2619 (N_2619,N_2435,N_2489);
or U2620 (N_2620,N_2510,N_2585);
and U2621 (N_2621,N_2437,N_2448);
or U2622 (N_2622,N_2575,N_2597);
nor U2623 (N_2623,N_2423,N_2599);
or U2624 (N_2624,N_2522,N_2425);
or U2625 (N_2625,N_2500,N_2595);
and U2626 (N_2626,N_2493,N_2480);
or U2627 (N_2627,N_2520,N_2521);
or U2628 (N_2628,N_2534,N_2563);
xor U2629 (N_2629,N_2581,N_2557);
and U2630 (N_2630,N_2512,N_2436);
nor U2631 (N_2631,N_2532,N_2454);
xor U2632 (N_2632,N_2574,N_2483);
or U2633 (N_2633,N_2556,N_2466);
and U2634 (N_2634,N_2475,N_2408);
nor U2635 (N_2635,N_2507,N_2533);
or U2636 (N_2636,N_2539,N_2593);
or U2637 (N_2637,N_2438,N_2464);
nor U2638 (N_2638,N_2591,N_2531);
xnor U2639 (N_2639,N_2572,N_2473);
or U2640 (N_2640,N_2577,N_2451);
and U2641 (N_2641,N_2564,N_2524);
nand U2642 (N_2642,N_2516,N_2566);
or U2643 (N_2643,N_2501,N_2404);
or U2644 (N_2644,N_2503,N_2526);
nor U2645 (N_2645,N_2458,N_2420);
xor U2646 (N_2646,N_2552,N_2465);
nor U2647 (N_2647,N_2496,N_2472);
or U2648 (N_2648,N_2491,N_2481);
or U2649 (N_2649,N_2527,N_2582);
nor U2650 (N_2650,N_2514,N_2594);
or U2651 (N_2651,N_2478,N_2416);
xnor U2652 (N_2652,N_2449,N_2418);
or U2653 (N_2653,N_2525,N_2535);
and U2654 (N_2654,N_2589,N_2548);
xnor U2655 (N_2655,N_2544,N_2584);
xor U2656 (N_2656,N_2573,N_2445);
and U2657 (N_2657,N_2553,N_2441);
nand U2658 (N_2658,N_2509,N_2470);
nor U2659 (N_2659,N_2417,N_2440);
and U2660 (N_2660,N_2555,N_2488);
nand U2661 (N_2661,N_2407,N_2528);
xnor U2662 (N_2662,N_2433,N_2477);
and U2663 (N_2663,N_2580,N_2432);
nor U2664 (N_2664,N_2565,N_2474);
nor U2665 (N_2665,N_2547,N_2495);
xnor U2666 (N_2666,N_2486,N_2558);
and U2667 (N_2667,N_2411,N_2406);
or U2668 (N_2668,N_2403,N_2459);
or U2669 (N_2669,N_2588,N_2550);
nand U2670 (N_2670,N_2447,N_2596);
nor U2671 (N_2671,N_2471,N_2506);
and U2672 (N_2672,N_2523,N_2450);
nor U2673 (N_2673,N_2559,N_2587);
xor U2674 (N_2674,N_2479,N_2504);
nor U2675 (N_2675,N_2460,N_2546);
nand U2676 (N_2676,N_2517,N_2453);
nand U2677 (N_2677,N_2457,N_2461);
and U2678 (N_2678,N_2429,N_2428);
and U2679 (N_2679,N_2476,N_2442);
and U2680 (N_2680,N_2519,N_2542);
and U2681 (N_2681,N_2430,N_2494);
nor U2682 (N_2682,N_2537,N_2468);
xnor U2683 (N_2683,N_2434,N_2508);
xor U2684 (N_2684,N_2463,N_2561);
xnor U2685 (N_2685,N_2543,N_2422);
xnor U2686 (N_2686,N_2482,N_2518);
and U2687 (N_2687,N_2545,N_2484);
and U2688 (N_2688,N_2579,N_2497);
xnor U2689 (N_2689,N_2515,N_2443);
nor U2690 (N_2690,N_2439,N_2455);
xor U2691 (N_2691,N_2576,N_2492);
and U2692 (N_2692,N_2487,N_2424);
nand U2693 (N_2693,N_2410,N_2401);
nor U2694 (N_2694,N_2502,N_2431);
nor U2695 (N_2695,N_2551,N_2414);
xor U2696 (N_2696,N_2562,N_2452);
nand U2697 (N_2697,N_2467,N_2412);
or U2698 (N_2698,N_2462,N_2592);
xnor U2699 (N_2699,N_2405,N_2505);
and U2700 (N_2700,N_2562,N_2419);
and U2701 (N_2701,N_2564,N_2551);
xor U2702 (N_2702,N_2544,N_2427);
or U2703 (N_2703,N_2549,N_2512);
and U2704 (N_2704,N_2467,N_2503);
xnor U2705 (N_2705,N_2582,N_2485);
and U2706 (N_2706,N_2580,N_2469);
and U2707 (N_2707,N_2481,N_2420);
and U2708 (N_2708,N_2446,N_2585);
or U2709 (N_2709,N_2473,N_2540);
or U2710 (N_2710,N_2584,N_2483);
nand U2711 (N_2711,N_2466,N_2402);
xnor U2712 (N_2712,N_2427,N_2555);
nand U2713 (N_2713,N_2417,N_2536);
and U2714 (N_2714,N_2419,N_2498);
xnor U2715 (N_2715,N_2599,N_2509);
xnor U2716 (N_2716,N_2438,N_2597);
xor U2717 (N_2717,N_2519,N_2461);
nand U2718 (N_2718,N_2446,N_2576);
xnor U2719 (N_2719,N_2476,N_2568);
or U2720 (N_2720,N_2428,N_2500);
or U2721 (N_2721,N_2584,N_2458);
nor U2722 (N_2722,N_2591,N_2435);
nor U2723 (N_2723,N_2524,N_2491);
nand U2724 (N_2724,N_2531,N_2550);
or U2725 (N_2725,N_2510,N_2467);
xor U2726 (N_2726,N_2575,N_2503);
nor U2727 (N_2727,N_2597,N_2476);
xor U2728 (N_2728,N_2408,N_2499);
nor U2729 (N_2729,N_2593,N_2485);
nor U2730 (N_2730,N_2427,N_2558);
or U2731 (N_2731,N_2548,N_2487);
xor U2732 (N_2732,N_2515,N_2457);
nor U2733 (N_2733,N_2585,N_2450);
or U2734 (N_2734,N_2451,N_2489);
xnor U2735 (N_2735,N_2465,N_2481);
nand U2736 (N_2736,N_2493,N_2473);
nand U2737 (N_2737,N_2459,N_2488);
xor U2738 (N_2738,N_2537,N_2463);
nand U2739 (N_2739,N_2523,N_2501);
xor U2740 (N_2740,N_2475,N_2538);
or U2741 (N_2741,N_2509,N_2591);
or U2742 (N_2742,N_2409,N_2459);
and U2743 (N_2743,N_2576,N_2420);
nor U2744 (N_2744,N_2426,N_2425);
or U2745 (N_2745,N_2571,N_2501);
xnor U2746 (N_2746,N_2409,N_2457);
xnor U2747 (N_2747,N_2527,N_2496);
nand U2748 (N_2748,N_2401,N_2427);
or U2749 (N_2749,N_2453,N_2531);
xor U2750 (N_2750,N_2583,N_2565);
and U2751 (N_2751,N_2513,N_2410);
nand U2752 (N_2752,N_2504,N_2449);
nand U2753 (N_2753,N_2567,N_2592);
or U2754 (N_2754,N_2437,N_2584);
nor U2755 (N_2755,N_2491,N_2499);
nor U2756 (N_2756,N_2595,N_2505);
and U2757 (N_2757,N_2482,N_2448);
xor U2758 (N_2758,N_2575,N_2539);
nand U2759 (N_2759,N_2417,N_2405);
nand U2760 (N_2760,N_2451,N_2546);
or U2761 (N_2761,N_2515,N_2492);
nand U2762 (N_2762,N_2432,N_2481);
xor U2763 (N_2763,N_2471,N_2592);
and U2764 (N_2764,N_2495,N_2435);
nand U2765 (N_2765,N_2481,N_2422);
and U2766 (N_2766,N_2427,N_2523);
nor U2767 (N_2767,N_2560,N_2511);
nor U2768 (N_2768,N_2437,N_2433);
xor U2769 (N_2769,N_2444,N_2435);
xnor U2770 (N_2770,N_2470,N_2508);
nand U2771 (N_2771,N_2543,N_2456);
nand U2772 (N_2772,N_2548,N_2519);
and U2773 (N_2773,N_2444,N_2566);
and U2774 (N_2774,N_2506,N_2462);
xnor U2775 (N_2775,N_2470,N_2450);
and U2776 (N_2776,N_2441,N_2431);
and U2777 (N_2777,N_2480,N_2448);
or U2778 (N_2778,N_2510,N_2594);
nand U2779 (N_2779,N_2463,N_2594);
and U2780 (N_2780,N_2440,N_2523);
nor U2781 (N_2781,N_2438,N_2520);
or U2782 (N_2782,N_2440,N_2585);
nand U2783 (N_2783,N_2576,N_2487);
and U2784 (N_2784,N_2580,N_2452);
or U2785 (N_2785,N_2515,N_2589);
nand U2786 (N_2786,N_2412,N_2413);
xor U2787 (N_2787,N_2428,N_2537);
nand U2788 (N_2788,N_2480,N_2412);
nor U2789 (N_2789,N_2492,N_2545);
nor U2790 (N_2790,N_2451,N_2464);
or U2791 (N_2791,N_2559,N_2496);
or U2792 (N_2792,N_2420,N_2497);
or U2793 (N_2793,N_2586,N_2559);
xnor U2794 (N_2794,N_2530,N_2429);
nand U2795 (N_2795,N_2525,N_2590);
xor U2796 (N_2796,N_2486,N_2441);
nor U2797 (N_2797,N_2491,N_2453);
and U2798 (N_2798,N_2426,N_2449);
xnor U2799 (N_2799,N_2566,N_2438);
nor U2800 (N_2800,N_2756,N_2632);
nor U2801 (N_2801,N_2741,N_2710);
and U2802 (N_2802,N_2673,N_2616);
xnor U2803 (N_2803,N_2605,N_2725);
nand U2804 (N_2804,N_2682,N_2743);
or U2805 (N_2805,N_2792,N_2728);
and U2806 (N_2806,N_2630,N_2608);
xor U2807 (N_2807,N_2600,N_2647);
nand U2808 (N_2808,N_2736,N_2637);
or U2809 (N_2809,N_2612,N_2752);
nor U2810 (N_2810,N_2604,N_2702);
xor U2811 (N_2811,N_2690,N_2732);
xnor U2812 (N_2812,N_2731,N_2615);
nor U2813 (N_2813,N_2685,N_2622);
and U2814 (N_2814,N_2755,N_2699);
xnor U2815 (N_2815,N_2665,N_2761);
or U2816 (N_2816,N_2719,N_2705);
and U2817 (N_2817,N_2675,N_2652);
nor U2818 (N_2818,N_2687,N_2672);
nand U2819 (N_2819,N_2669,N_2763);
or U2820 (N_2820,N_2779,N_2644);
nor U2821 (N_2821,N_2711,N_2636);
and U2822 (N_2822,N_2631,N_2775);
and U2823 (N_2823,N_2733,N_2683);
nor U2824 (N_2824,N_2718,N_2772);
or U2825 (N_2825,N_2712,N_2714);
xnor U2826 (N_2826,N_2793,N_2701);
nor U2827 (N_2827,N_2740,N_2746);
nor U2828 (N_2828,N_2601,N_2767);
or U2829 (N_2829,N_2643,N_2610);
or U2830 (N_2830,N_2624,N_2656);
nand U2831 (N_2831,N_2694,N_2759);
and U2832 (N_2832,N_2771,N_2753);
or U2833 (N_2833,N_2639,N_2726);
and U2834 (N_2834,N_2789,N_2773);
nand U2835 (N_2835,N_2762,N_2623);
nor U2836 (N_2836,N_2655,N_2668);
xor U2837 (N_2837,N_2768,N_2620);
xnor U2838 (N_2838,N_2757,N_2716);
and U2839 (N_2839,N_2609,N_2654);
or U2840 (N_2840,N_2730,N_2723);
xor U2841 (N_2841,N_2602,N_2786);
xor U2842 (N_2842,N_2742,N_2765);
nand U2843 (N_2843,N_2778,N_2737);
xnor U2844 (N_2844,N_2735,N_2641);
nand U2845 (N_2845,N_2670,N_2770);
nand U2846 (N_2846,N_2780,N_2646);
or U2847 (N_2847,N_2677,N_2720);
nand U2848 (N_2848,N_2794,N_2783);
nand U2849 (N_2849,N_2662,N_2707);
nand U2850 (N_2850,N_2717,N_2729);
or U2851 (N_2851,N_2678,N_2661);
nor U2852 (N_2852,N_2634,N_2704);
nand U2853 (N_2853,N_2744,N_2784);
xor U2854 (N_2854,N_2769,N_2750);
or U2855 (N_2855,N_2798,N_2739);
nand U2856 (N_2856,N_2697,N_2617);
nor U2857 (N_2857,N_2679,N_2791);
nand U2858 (N_2858,N_2635,N_2727);
nor U2859 (N_2859,N_2666,N_2628);
nor U2860 (N_2860,N_2626,N_2689);
xnor U2861 (N_2861,N_2664,N_2788);
xor U2862 (N_2862,N_2703,N_2642);
nor U2863 (N_2863,N_2721,N_2696);
nand U2864 (N_2864,N_2629,N_2619);
and U2865 (N_2865,N_2766,N_2603);
nand U2866 (N_2866,N_2688,N_2651);
or U2867 (N_2867,N_2648,N_2782);
or U2868 (N_2868,N_2734,N_2691);
nor U2869 (N_2869,N_2745,N_2749);
and U2870 (N_2870,N_2650,N_2613);
or U2871 (N_2871,N_2645,N_2700);
and U2872 (N_2872,N_2611,N_2671);
or U2873 (N_2873,N_2738,N_2797);
and U2874 (N_2874,N_2649,N_2676);
xnor U2875 (N_2875,N_2795,N_2627);
xor U2876 (N_2876,N_2660,N_2633);
and U2877 (N_2877,N_2680,N_2667);
nor U2878 (N_2878,N_2692,N_2722);
or U2879 (N_2879,N_2748,N_2684);
or U2880 (N_2880,N_2658,N_2693);
and U2881 (N_2881,N_2663,N_2713);
and U2882 (N_2882,N_2724,N_2751);
xnor U2883 (N_2883,N_2686,N_2674);
xnor U2884 (N_2884,N_2747,N_2790);
and U2885 (N_2885,N_2638,N_2659);
and U2886 (N_2886,N_2695,N_2754);
xor U2887 (N_2887,N_2614,N_2709);
and U2888 (N_2888,N_2625,N_2657);
nand U2889 (N_2889,N_2715,N_2698);
nand U2890 (N_2890,N_2606,N_2777);
nor U2891 (N_2891,N_2774,N_2787);
nand U2892 (N_2892,N_2706,N_2640);
or U2893 (N_2893,N_2785,N_2776);
xor U2894 (N_2894,N_2760,N_2607);
nor U2895 (N_2895,N_2796,N_2653);
and U2896 (N_2896,N_2618,N_2758);
or U2897 (N_2897,N_2621,N_2764);
xor U2898 (N_2898,N_2781,N_2708);
nor U2899 (N_2899,N_2799,N_2681);
and U2900 (N_2900,N_2783,N_2678);
and U2901 (N_2901,N_2683,N_2639);
nand U2902 (N_2902,N_2618,N_2663);
or U2903 (N_2903,N_2662,N_2701);
xor U2904 (N_2904,N_2641,N_2794);
and U2905 (N_2905,N_2636,N_2764);
nand U2906 (N_2906,N_2776,N_2684);
nand U2907 (N_2907,N_2700,N_2708);
or U2908 (N_2908,N_2609,N_2709);
and U2909 (N_2909,N_2715,N_2794);
nor U2910 (N_2910,N_2612,N_2618);
nand U2911 (N_2911,N_2606,N_2749);
and U2912 (N_2912,N_2655,N_2627);
xor U2913 (N_2913,N_2707,N_2605);
or U2914 (N_2914,N_2657,N_2745);
or U2915 (N_2915,N_2734,N_2738);
xor U2916 (N_2916,N_2617,N_2606);
and U2917 (N_2917,N_2779,N_2788);
and U2918 (N_2918,N_2720,N_2683);
nand U2919 (N_2919,N_2726,N_2719);
and U2920 (N_2920,N_2789,N_2612);
nor U2921 (N_2921,N_2723,N_2691);
and U2922 (N_2922,N_2759,N_2727);
xnor U2923 (N_2923,N_2645,N_2622);
nor U2924 (N_2924,N_2758,N_2669);
xor U2925 (N_2925,N_2638,N_2676);
nor U2926 (N_2926,N_2666,N_2608);
and U2927 (N_2927,N_2714,N_2652);
or U2928 (N_2928,N_2651,N_2710);
xor U2929 (N_2929,N_2757,N_2636);
nor U2930 (N_2930,N_2618,N_2799);
nand U2931 (N_2931,N_2638,N_2655);
or U2932 (N_2932,N_2754,N_2645);
and U2933 (N_2933,N_2779,N_2700);
nand U2934 (N_2934,N_2735,N_2623);
nor U2935 (N_2935,N_2639,N_2711);
xor U2936 (N_2936,N_2680,N_2795);
and U2937 (N_2937,N_2789,N_2646);
nor U2938 (N_2938,N_2723,N_2701);
and U2939 (N_2939,N_2710,N_2770);
and U2940 (N_2940,N_2735,N_2631);
nand U2941 (N_2941,N_2692,N_2616);
nand U2942 (N_2942,N_2601,N_2663);
and U2943 (N_2943,N_2722,N_2792);
xnor U2944 (N_2944,N_2600,N_2785);
and U2945 (N_2945,N_2669,N_2604);
xnor U2946 (N_2946,N_2769,N_2654);
xnor U2947 (N_2947,N_2799,N_2684);
nor U2948 (N_2948,N_2605,N_2701);
nor U2949 (N_2949,N_2737,N_2731);
xor U2950 (N_2950,N_2704,N_2640);
xor U2951 (N_2951,N_2738,N_2624);
nor U2952 (N_2952,N_2661,N_2712);
xor U2953 (N_2953,N_2664,N_2608);
or U2954 (N_2954,N_2727,N_2644);
nor U2955 (N_2955,N_2610,N_2711);
or U2956 (N_2956,N_2728,N_2633);
nand U2957 (N_2957,N_2728,N_2623);
nor U2958 (N_2958,N_2624,N_2748);
nor U2959 (N_2959,N_2663,N_2653);
and U2960 (N_2960,N_2734,N_2733);
and U2961 (N_2961,N_2794,N_2633);
xnor U2962 (N_2962,N_2641,N_2700);
nor U2963 (N_2963,N_2710,N_2780);
nor U2964 (N_2964,N_2711,N_2776);
nor U2965 (N_2965,N_2675,N_2753);
and U2966 (N_2966,N_2771,N_2688);
or U2967 (N_2967,N_2762,N_2777);
or U2968 (N_2968,N_2715,N_2734);
and U2969 (N_2969,N_2717,N_2693);
or U2970 (N_2970,N_2605,N_2657);
and U2971 (N_2971,N_2695,N_2684);
or U2972 (N_2972,N_2679,N_2606);
nor U2973 (N_2973,N_2603,N_2768);
or U2974 (N_2974,N_2739,N_2679);
xor U2975 (N_2975,N_2671,N_2685);
nor U2976 (N_2976,N_2715,N_2626);
xnor U2977 (N_2977,N_2676,N_2776);
nor U2978 (N_2978,N_2694,N_2712);
nor U2979 (N_2979,N_2712,N_2609);
nand U2980 (N_2980,N_2666,N_2755);
nand U2981 (N_2981,N_2764,N_2780);
nor U2982 (N_2982,N_2713,N_2724);
and U2983 (N_2983,N_2796,N_2631);
nor U2984 (N_2984,N_2620,N_2715);
or U2985 (N_2985,N_2670,N_2653);
nor U2986 (N_2986,N_2690,N_2719);
nand U2987 (N_2987,N_2730,N_2681);
or U2988 (N_2988,N_2778,N_2762);
or U2989 (N_2989,N_2623,N_2761);
or U2990 (N_2990,N_2652,N_2745);
nand U2991 (N_2991,N_2633,N_2775);
nor U2992 (N_2992,N_2741,N_2711);
nand U2993 (N_2993,N_2768,N_2716);
or U2994 (N_2994,N_2796,N_2721);
or U2995 (N_2995,N_2658,N_2631);
or U2996 (N_2996,N_2661,N_2736);
nor U2997 (N_2997,N_2644,N_2634);
xor U2998 (N_2998,N_2727,N_2647);
nor U2999 (N_2999,N_2665,N_2618);
and U3000 (N_3000,N_2917,N_2839);
nand U3001 (N_3001,N_2869,N_2944);
xnor U3002 (N_3002,N_2885,N_2967);
nor U3003 (N_3003,N_2914,N_2861);
and U3004 (N_3004,N_2829,N_2964);
or U3005 (N_3005,N_2928,N_2808);
xor U3006 (N_3006,N_2905,N_2804);
nor U3007 (N_3007,N_2925,N_2986);
nand U3008 (N_3008,N_2880,N_2844);
xor U3009 (N_3009,N_2897,N_2823);
and U3010 (N_3010,N_2998,N_2939);
nand U3011 (N_3011,N_2913,N_2972);
and U3012 (N_3012,N_2990,N_2920);
nand U3013 (N_3013,N_2931,N_2958);
and U3014 (N_3014,N_2859,N_2973);
nand U3015 (N_3015,N_2989,N_2940);
xor U3016 (N_3016,N_2827,N_2802);
nand U3017 (N_3017,N_2966,N_2898);
and U3018 (N_3018,N_2965,N_2826);
xor U3019 (N_3019,N_2831,N_2975);
and U3020 (N_3020,N_2969,N_2924);
xnor U3021 (N_3021,N_2961,N_2891);
nand U3022 (N_3022,N_2968,N_2817);
nand U3023 (N_3023,N_2910,N_2999);
xor U3024 (N_3024,N_2919,N_2815);
nor U3025 (N_3025,N_2980,N_2946);
nor U3026 (N_3026,N_2899,N_2895);
nand U3027 (N_3027,N_2811,N_2801);
nor U3028 (N_3028,N_2997,N_2988);
xor U3029 (N_3029,N_2821,N_2872);
and U3030 (N_3030,N_2810,N_2971);
or U3031 (N_3031,N_2888,N_2955);
nor U3032 (N_3032,N_2870,N_2952);
xnor U3033 (N_3033,N_2894,N_2948);
xnor U3034 (N_3034,N_2868,N_2953);
nor U3035 (N_3035,N_2838,N_2837);
and U3036 (N_3036,N_2960,N_2835);
xnor U3037 (N_3037,N_2876,N_2949);
nor U3038 (N_3038,N_2904,N_2819);
or U3039 (N_3039,N_2865,N_2806);
nand U3040 (N_3040,N_2991,N_2995);
nor U3041 (N_3041,N_2881,N_2850);
or U3042 (N_3042,N_2916,N_2959);
nand U3043 (N_3043,N_2922,N_2884);
nand U3044 (N_3044,N_2851,N_2800);
or U3045 (N_3045,N_2987,N_2896);
nand U3046 (N_3046,N_2822,N_2882);
or U3047 (N_3047,N_2963,N_2954);
nand U3048 (N_3048,N_2974,N_2903);
xor U3049 (N_3049,N_2848,N_2845);
and U3050 (N_3050,N_2816,N_2849);
nand U3051 (N_3051,N_2942,N_2856);
or U3052 (N_3052,N_2812,N_2840);
xnor U3053 (N_3053,N_2814,N_2828);
xor U3054 (N_3054,N_2836,N_2858);
nor U3055 (N_3055,N_2996,N_2886);
xor U3056 (N_3056,N_2893,N_2824);
or U3057 (N_3057,N_2943,N_2956);
or U3058 (N_3058,N_2841,N_2833);
or U3059 (N_3059,N_2901,N_2879);
or U3060 (N_3060,N_2825,N_2979);
xor U3061 (N_3061,N_2809,N_2842);
xor U3062 (N_3062,N_2871,N_2992);
or U3063 (N_3063,N_2950,N_2981);
or U3064 (N_3064,N_2951,N_2935);
nand U3065 (N_3065,N_2873,N_2962);
xor U3066 (N_3066,N_2866,N_2985);
nor U3067 (N_3067,N_2957,N_2887);
and U3068 (N_3068,N_2921,N_2941);
xnor U3069 (N_3069,N_2923,N_2807);
or U3070 (N_3070,N_2993,N_2982);
and U3071 (N_3071,N_2853,N_2915);
nor U3072 (N_3072,N_2883,N_2854);
and U3073 (N_3073,N_2805,N_2994);
and U3074 (N_3074,N_2936,N_2857);
and U3075 (N_3075,N_2867,N_2830);
or U3076 (N_3076,N_2818,N_2878);
nor U3077 (N_3077,N_2820,N_2918);
nor U3078 (N_3078,N_2846,N_2908);
nor U3079 (N_3079,N_2947,N_2877);
or U3080 (N_3080,N_2900,N_2937);
nor U3081 (N_3081,N_2929,N_2911);
xor U3082 (N_3082,N_2926,N_2930);
or U3083 (N_3083,N_2890,N_2843);
or U3084 (N_3084,N_2852,N_2977);
nor U3085 (N_3085,N_2927,N_2983);
and U3086 (N_3086,N_2932,N_2874);
or U3087 (N_3087,N_2889,N_2984);
xnor U3088 (N_3088,N_2934,N_2945);
nand U3089 (N_3089,N_2907,N_2832);
or U3090 (N_3090,N_2909,N_2933);
xor U3091 (N_3091,N_2978,N_2906);
nor U3092 (N_3092,N_2855,N_2847);
and U3093 (N_3093,N_2912,N_2863);
and U3094 (N_3094,N_2976,N_2938);
and U3095 (N_3095,N_2803,N_2860);
and U3096 (N_3096,N_2970,N_2862);
nor U3097 (N_3097,N_2902,N_2864);
and U3098 (N_3098,N_2834,N_2892);
xnor U3099 (N_3099,N_2875,N_2813);
xor U3100 (N_3100,N_2966,N_2904);
or U3101 (N_3101,N_2875,N_2858);
or U3102 (N_3102,N_2827,N_2804);
nand U3103 (N_3103,N_2935,N_2838);
or U3104 (N_3104,N_2980,N_2864);
nand U3105 (N_3105,N_2876,N_2933);
nor U3106 (N_3106,N_2902,N_2801);
or U3107 (N_3107,N_2841,N_2939);
or U3108 (N_3108,N_2804,N_2987);
and U3109 (N_3109,N_2834,N_2850);
xnor U3110 (N_3110,N_2829,N_2916);
nand U3111 (N_3111,N_2932,N_2943);
or U3112 (N_3112,N_2846,N_2907);
and U3113 (N_3113,N_2867,N_2805);
or U3114 (N_3114,N_2880,N_2867);
nor U3115 (N_3115,N_2928,N_2998);
nor U3116 (N_3116,N_2968,N_2930);
or U3117 (N_3117,N_2964,N_2907);
or U3118 (N_3118,N_2942,N_2860);
and U3119 (N_3119,N_2961,N_2912);
xnor U3120 (N_3120,N_2936,N_2991);
nand U3121 (N_3121,N_2984,N_2901);
nand U3122 (N_3122,N_2980,N_2830);
or U3123 (N_3123,N_2951,N_2936);
and U3124 (N_3124,N_2814,N_2890);
and U3125 (N_3125,N_2965,N_2923);
xnor U3126 (N_3126,N_2901,N_2896);
xnor U3127 (N_3127,N_2874,N_2930);
xor U3128 (N_3128,N_2872,N_2852);
nand U3129 (N_3129,N_2949,N_2849);
or U3130 (N_3130,N_2958,N_2871);
and U3131 (N_3131,N_2954,N_2833);
nand U3132 (N_3132,N_2803,N_2812);
nand U3133 (N_3133,N_2960,N_2944);
xor U3134 (N_3134,N_2971,N_2857);
or U3135 (N_3135,N_2956,N_2812);
nand U3136 (N_3136,N_2966,N_2936);
nor U3137 (N_3137,N_2846,N_2854);
nand U3138 (N_3138,N_2919,N_2977);
xor U3139 (N_3139,N_2905,N_2997);
xnor U3140 (N_3140,N_2956,N_2997);
xor U3141 (N_3141,N_2893,N_2871);
and U3142 (N_3142,N_2908,N_2824);
or U3143 (N_3143,N_2958,N_2875);
nand U3144 (N_3144,N_2966,N_2946);
xnor U3145 (N_3145,N_2872,N_2937);
and U3146 (N_3146,N_2803,N_2952);
nand U3147 (N_3147,N_2873,N_2804);
and U3148 (N_3148,N_2981,N_2856);
nand U3149 (N_3149,N_2990,N_2895);
nand U3150 (N_3150,N_2966,N_2840);
or U3151 (N_3151,N_2839,N_2887);
and U3152 (N_3152,N_2953,N_2867);
or U3153 (N_3153,N_2875,N_2897);
xor U3154 (N_3154,N_2952,N_2891);
xnor U3155 (N_3155,N_2917,N_2826);
and U3156 (N_3156,N_2987,N_2862);
nor U3157 (N_3157,N_2951,N_2917);
and U3158 (N_3158,N_2822,N_2811);
xnor U3159 (N_3159,N_2999,N_2974);
xor U3160 (N_3160,N_2974,N_2814);
nand U3161 (N_3161,N_2882,N_2893);
nand U3162 (N_3162,N_2923,N_2930);
nand U3163 (N_3163,N_2922,N_2935);
and U3164 (N_3164,N_2848,N_2838);
nand U3165 (N_3165,N_2870,N_2934);
or U3166 (N_3166,N_2866,N_2895);
nand U3167 (N_3167,N_2894,N_2875);
and U3168 (N_3168,N_2844,N_2941);
or U3169 (N_3169,N_2871,N_2846);
nor U3170 (N_3170,N_2829,N_2811);
nand U3171 (N_3171,N_2923,N_2851);
or U3172 (N_3172,N_2912,N_2841);
nor U3173 (N_3173,N_2800,N_2954);
nor U3174 (N_3174,N_2813,N_2855);
nand U3175 (N_3175,N_2929,N_2947);
nor U3176 (N_3176,N_2974,N_2994);
xnor U3177 (N_3177,N_2914,N_2957);
or U3178 (N_3178,N_2872,N_2800);
nor U3179 (N_3179,N_2985,N_2940);
nor U3180 (N_3180,N_2812,N_2948);
nand U3181 (N_3181,N_2897,N_2984);
nand U3182 (N_3182,N_2919,N_2822);
xor U3183 (N_3183,N_2940,N_2869);
and U3184 (N_3184,N_2888,N_2991);
xor U3185 (N_3185,N_2840,N_2982);
nor U3186 (N_3186,N_2982,N_2874);
or U3187 (N_3187,N_2847,N_2871);
and U3188 (N_3188,N_2948,N_2813);
nor U3189 (N_3189,N_2967,N_2866);
nor U3190 (N_3190,N_2956,N_2838);
xnor U3191 (N_3191,N_2970,N_2916);
and U3192 (N_3192,N_2811,N_2850);
nor U3193 (N_3193,N_2927,N_2896);
nand U3194 (N_3194,N_2897,N_2849);
or U3195 (N_3195,N_2870,N_2988);
xnor U3196 (N_3196,N_2865,N_2950);
nand U3197 (N_3197,N_2960,N_2959);
and U3198 (N_3198,N_2902,N_2999);
nor U3199 (N_3199,N_2867,N_2850);
nor U3200 (N_3200,N_3021,N_3152);
nor U3201 (N_3201,N_3116,N_3065);
and U3202 (N_3202,N_3103,N_3167);
nand U3203 (N_3203,N_3113,N_3105);
or U3204 (N_3204,N_3177,N_3134);
and U3205 (N_3205,N_3074,N_3026);
nand U3206 (N_3206,N_3019,N_3030);
or U3207 (N_3207,N_3023,N_3137);
xor U3208 (N_3208,N_3064,N_3079);
nand U3209 (N_3209,N_3052,N_3133);
xnor U3210 (N_3210,N_3163,N_3087);
nor U3211 (N_3211,N_3169,N_3076);
or U3212 (N_3212,N_3162,N_3014);
nand U3213 (N_3213,N_3101,N_3082);
nor U3214 (N_3214,N_3010,N_3012);
nand U3215 (N_3215,N_3121,N_3047);
nor U3216 (N_3216,N_3093,N_3092);
xor U3217 (N_3217,N_3122,N_3127);
and U3218 (N_3218,N_3172,N_3187);
or U3219 (N_3219,N_3056,N_3181);
nand U3220 (N_3220,N_3000,N_3009);
nor U3221 (N_3221,N_3060,N_3164);
nor U3222 (N_3222,N_3085,N_3048);
nor U3223 (N_3223,N_3018,N_3110);
xor U3224 (N_3224,N_3128,N_3017);
and U3225 (N_3225,N_3183,N_3155);
and U3226 (N_3226,N_3198,N_3178);
and U3227 (N_3227,N_3096,N_3156);
xnor U3228 (N_3228,N_3095,N_3193);
xor U3229 (N_3229,N_3044,N_3022);
nor U3230 (N_3230,N_3180,N_3192);
xnor U3231 (N_3231,N_3150,N_3111);
nand U3232 (N_3232,N_3040,N_3147);
nor U3233 (N_3233,N_3153,N_3175);
nand U3234 (N_3234,N_3179,N_3077);
or U3235 (N_3235,N_3090,N_3188);
nor U3236 (N_3236,N_3028,N_3058);
or U3237 (N_3237,N_3125,N_3020);
or U3238 (N_3238,N_3114,N_3130);
and U3239 (N_3239,N_3142,N_3015);
and U3240 (N_3240,N_3034,N_3036);
or U3241 (N_3241,N_3124,N_3126);
nor U3242 (N_3242,N_3136,N_3051);
and U3243 (N_3243,N_3002,N_3099);
or U3244 (N_3244,N_3050,N_3118);
nor U3245 (N_3245,N_3158,N_3146);
or U3246 (N_3246,N_3184,N_3001);
nand U3247 (N_3247,N_3173,N_3185);
or U3248 (N_3248,N_3004,N_3145);
nor U3249 (N_3249,N_3117,N_3123);
nor U3250 (N_3250,N_3088,N_3013);
and U3251 (N_3251,N_3190,N_3038);
xnor U3252 (N_3252,N_3106,N_3005);
xnor U3253 (N_3253,N_3182,N_3032);
or U3254 (N_3254,N_3166,N_3072);
xor U3255 (N_3255,N_3140,N_3100);
or U3256 (N_3256,N_3160,N_3008);
xor U3257 (N_3257,N_3196,N_3068);
nand U3258 (N_3258,N_3104,N_3186);
nor U3259 (N_3259,N_3086,N_3097);
nand U3260 (N_3260,N_3066,N_3119);
or U3261 (N_3261,N_3171,N_3161);
xnor U3262 (N_3262,N_3141,N_3041);
or U3263 (N_3263,N_3091,N_3081);
or U3264 (N_3264,N_3073,N_3011);
nor U3265 (N_3265,N_3035,N_3176);
or U3266 (N_3266,N_3129,N_3078);
or U3267 (N_3267,N_3109,N_3159);
xnor U3268 (N_3268,N_3075,N_3049);
and U3269 (N_3269,N_3089,N_3157);
nor U3270 (N_3270,N_3107,N_3054);
nor U3271 (N_3271,N_3170,N_3042);
xor U3272 (N_3272,N_3053,N_3025);
and U3273 (N_3273,N_3098,N_3080);
and U3274 (N_3274,N_3059,N_3069);
and U3275 (N_3275,N_3131,N_3003);
and U3276 (N_3276,N_3191,N_3067);
xor U3277 (N_3277,N_3151,N_3148);
nand U3278 (N_3278,N_3149,N_3194);
and U3279 (N_3279,N_3165,N_3029);
and U3280 (N_3280,N_3046,N_3197);
xnor U3281 (N_3281,N_3062,N_3063);
nand U3282 (N_3282,N_3135,N_3061);
or U3283 (N_3283,N_3168,N_3115);
and U3284 (N_3284,N_3037,N_3094);
and U3285 (N_3285,N_3024,N_3084);
and U3286 (N_3286,N_3071,N_3027);
xnor U3287 (N_3287,N_3070,N_3033);
and U3288 (N_3288,N_3195,N_3174);
nand U3289 (N_3289,N_3138,N_3043);
nor U3290 (N_3290,N_3083,N_3045);
nand U3291 (N_3291,N_3039,N_3102);
nand U3292 (N_3292,N_3112,N_3144);
or U3293 (N_3293,N_3108,N_3139);
and U3294 (N_3294,N_3006,N_3016);
nor U3295 (N_3295,N_3007,N_3031);
xor U3296 (N_3296,N_3057,N_3055);
or U3297 (N_3297,N_3199,N_3132);
nand U3298 (N_3298,N_3189,N_3120);
or U3299 (N_3299,N_3143,N_3154);
nor U3300 (N_3300,N_3158,N_3035);
nor U3301 (N_3301,N_3161,N_3023);
and U3302 (N_3302,N_3095,N_3107);
nand U3303 (N_3303,N_3056,N_3176);
nor U3304 (N_3304,N_3081,N_3139);
nand U3305 (N_3305,N_3136,N_3064);
or U3306 (N_3306,N_3187,N_3081);
or U3307 (N_3307,N_3135,N_3073);
and U3308 (N_3308,N_3023,N_3132);
nand U3309 (N_3309,N_3090,N_3194);
nand U3310 (N_3310,N_3104,N_3172);
or U3311 (N_3311,N_3065,N_3063);
nor U3312 (N_3312,N_3187,N_3180);
xor U3313 (N_3313,N_3193,N_3096);
and U3314 (N_3314,N_3163,N_3084);
nand U3315 (N_3315,N_3051,N_3175);
and U3316 (N_3316,N_3197,N_3042);
and U3317 (N_3317,N_3184,N_3197);
nor U3318 (N_3318,N_3181,N_3193);
or U3319 (N_3319,N_3185,N_3199);
nor U3320 (N_3320,N_3155,N_3141);
nor U3321 (N_3321,N_3140,N_3160);
and U3322 (N_3322,N_3096,N_3183);
and U3323 (N_3323,N_3068,N_3180);
xnor U3324 (N_3324,N_3093,N_3190);
nor U3325 (N_3325,N_3043,N_3040);
xor U3326 (N_3326,N_3030,N_3191);
and U3327 (N_3327,N_3152,N_3150);
nor U3328 (N_3328,N_3197,N_3075);
or U3329 (N_3329,N_3052,N_3018);
and U3330 (N_3330,N_3088,N_3006);
and U3331 (N_3331,N_3052,N_3167);
or U3332 (N_3332,N_3125,N_3039);
and U3333 (N_3333,N_3060,N_3146);
nand U3334 (N_3334,N_3168,N_3076);
nand U3335 (N_3335,N_3078,N_3133);
nand U3336 (N_3336,N_3144,N_3015);
nor U3337 (N_3337,N_3160,N_3094);
and U3338 (N_3338,N_3100,N_3196);
nand U3339 (N_3339,N_3190,N_3066);
xor U3340 (N_3340,N_3183,N_3036);
xor U3341 (N_3341,N_3090,N_3158);
nand U3342 (N_3342,N_3121,N_3130);
nand U3343 (N_3343,N_3055,N_3072);
or U3344 (N_3344,N_3018,N_3123);
xnor U3345 (N_3345,N_3027,N_3125);
and U3346 (N_3346,N_3056,N_3137);
xor U3347 (N_3347,N_3107,N_3050);
xnor U3348 (N_3348,N_3112,N_3051);
xnor U3349 (N_3349,N_3111,N_3100);
nor U3350 (N_3350,N_3198,N_3150);
xnor U3351 (N_3351,N_3110,N_3114);
or U3352 (N_3352,N_3044,N_3144);
nand U3353 (N_3353,N_3094,N_3015);
or U3354 (N_3354,N_3102,N_3081);
nor U3355 (N_3355,N_3105,N_3114);
or U3356 (N_3356,N_3152,N_3098);
and U3357 (N_3357,N_3113,N_3133);
nor U3358 (N_3358,N_3017,N_3161);
nor U3359 (N_3359,N_3181,N_3099);
nand U3360 (N_3360,N_3021,N_3057);
and U3361 (N_3361,N_3032,N_3023);
nand U3362 (N_3362,N_3154,N_3186);
or U3363 (N_3363,N_3128,N_3195);
nand U3364 (N_3364,N_3007,N_3098);
or U3365 (N_3365,N_3009,N_3082);
nand U3366 (N_3366,N_3088,N_3068);
and U3367 (N_3367,N_3147,N_3066);
xnor U3368 (N_3368,N_3132,N_3012);
xnor U3369 (N_3369,N_3149,N_3199);
or U3370 (N_3370,N_3174,N_3061);
and U3371 (N_3371,N_3004,N_3152);
xnor U3372 (N_3372,N_3084,N_3042);
nor U3373 (N_3373,N_3094,N_3020);
nor U3374 (N_3374,N_3090,N_3064);
and U3375 (N_3375,N_3019,N_3027);
nand U3376 (N_3376,N_3097,N_3053);
nor U3377 (N_3377,N_3182,N_3177);
xnor U3378 (N_3378,N_3045,N_3128);
and U3379 (N_3379,N_3110,N_3139);
nand U3380 (N_3380,N_3010,N_3069);
and U3381 (N_3381,N_3112,N_3071);
and U3382 (N_3382,N_3173,N_3146);
nor U3383 (N_3383,N_3141,N_3142);
nand U3384 (N_3384,N_3186,N_3060);
nor U3385 (N_3385,N_3105,N_3059);
nor U3386 (N_3386,N_3167,N_3105);
or U3387 (N_3387,N_3068,N_3138);
and U3388 (N_3388,N_3134,N_3034);
and U3389 (N_3389,N_3181,N_3075);
nor U3390 (N_3390,N_3123,N_3080);
nor U3391 (N_3391,N_3056,N_3125);
or U3392 (N_3392,N_3151,N_3096);
nand U3393 (N_3393,N_3174,N_3067);
and U3394 (N_3394,N_3145,N_3023);
nand U3395 (N_3395,N_3186,N_3119);
nor U3396 (N_3396,N_3143,N_3170);
or U3397 (N_3397,N_3145,N_3153);
and U3398 (N_3398,N_3028,N_3159);
nand U3399 (N_3399,N_3110,N_3033);
nand U3400 (N_3400,N_3331,N_3314);
or U3401 (N_3401,N_3397,N_3286);
nor U3402 (N_3402,N_3366,N_3277);
and U3403 (N_3403,N_3399,N_3227);
nor U3404 (N_3404,N_3289,N_3212);
and U3405 (N_3405,N_3240,N_3288);
xnor U3406 (N_3406,N_3296,N_3283);
nor U3407 (N_3407,N_3217,N_3219);
and U3408 (N_3408,N_3231,N_3222);
nor U3409 (N_3409,N_3254,N_3360);
or U3410 (N_3410,N_3332,N_3259);
xor U3411 (N_3411,N_3234,N_3373);
or U3412 (N_3412,N_3301,N_3232);
or U3413 (N_3413,N_3356,N_3276);
xor U3414 (N_3414,N_3305,N_3316);
xnor U3415 (N_3415,N_3229,N_3261);
nand U3416 (N_3416,N_3355,N_3207);
nand U3417 (N_3417,N_3224,N_3327);
nor U3418 (N_3418,N_3392,N_3326);
xnor U3419 (N_3419,N_3223,N_3368);
or U3420 (N_3420,N_3202,N_3213);
nand U3421 (N_3421,N_3307,N_3270);
xnor U3422 (N_3422,N_3280,N_3258);
nor U3423 (N_3423,N_3386,N_3230);
xnor U3424 (N_3424,N_3244,N_3354);
nor U3425 (N_3425,N_3236,N_3242);
and U3426 (N_3426,N_3380,N_3334);
nand U3427 (N_3427,N_3214,N_3357);
xor U3428 (N_3428,N_3315,N_3274);
or U3429 (N_3429,N_3353,N_3374);
and U3430 (N_3430,N_3248,N_3204);
nor U3431 (N_3431,N_3279,N_3350);
and U3432 (N_3432,N_3383,N_3255);
nand U3433 (N_3433,N_3273,N_3284);
nand U3434 (N_3434,N_3239,N_3226);
or U3435 (N_3435,N_3395,N_3385);
and U3436 (N_3436,N_3343,N_3324);
xnor U3437 (N_3437,N_3361,N_3210);
and U3438 (N_3438,N_3206,N_3209);
xnor U3439 (N_3439,N_3338,N_3352);
and U3440 (N_3440,N_3396,N_3295);
xnor U3441 (N_3441,N_3225,N_3370);
or U3442 (N_3442,N_3318,N_3320);
xnor U3443 (N_3443,N_3233,N_3345);
and U3444 (N_3444,N_3387,N_3351);
xnor U3445 (N_3445,N_3391,N_3249);
and U3446 (N_3446,N_3294,N_3260);
or U3447 (N_3447,N_3247,N_3382);
nand U3448 (N_3448,N_3333,N_3252);
and U3449 (N_3449,N_3319,N_3265);
nor U3450 (N_3450,N_3359,N_3228);
nand U3451 (N_3451,N_3309,N_3300);
nand U3452 (N_3452,N_3215,N_3381);
xnor U3453 (N_3453,N_3310,N_3369);
nor U3454 (N_3454,N_3264,N_3275);
xnor U3455 (N_3455,N_3220,N_3358);
nor U3456 (N_3456,N_3313,N_3329);
xor U3457 (N_3457,N_3216,N_3297);
nand U3458 (N_3458,N_3347,N_3268);
or U3459 (N_3459,N_3367,N_3384);
nor U3460 (N_3460,N_3340,N_3290);
nand U3461 (N_3461,N_3371,N_3344);
nor U3462 (N_3462,N_3211,N_3263);
and U3463 (N_3463,N_3235,N_3237);
xnor U3464 (N_3464,N_3201,N_3308);
xnor U3465 (N_3465,N_3363,N_3218);
and U3466 (N_3466,N_3398,N_3266);
and U3467 (N_3467,N_3322,N_3200);
or U3468 (N_3468,N_3245,N_3271);
and U3469 (N_3469,N_3378,N_3349);
and U3470 (N_3470,N_3299,N_3241);
xnor U3471 (N_3471,N_3388,N_3282);
or U3472 (N_3472,N_3262,N_3250);
and U3473 (N_3473,N_3394,N_3330);
nor U3474 (N_3474,N_3304,N_3365);
or U3475 (N_3475,N_3272,N_3375);
nand U3476 (N_3476,N_3376,N_3253);
or U3477 (N_3477,N_3321,N_3205);
xor U3478 (N_3478,N_3302,N_3311);
or U3479 (N_3479,N_3298,N_3303);
nor U3480 (N_3480,N_3292,N_3203);
and U3481 (N_3481,N_3246,N_3328);
nand U3482 (N_3482,N_3393,N_3337);
nand U3483 (N_3483,N_3348,N_3287);
and U3484 (N_3484,N_3377,N_3267);
and U3485 (N_3485,N_3251,N_3278);
nand U3486 (N_3486,N_3346,N_3342);
nand U3487 (N_3487,N_3389,N_3281);
xnor U3488 (N_3488,N_3372,N_3341);
and U3489 (N_3489,N_3306,N_3390);
or U3490 (N_3490,N_3325,N_3293);
and U3491 (N_3491,N_3291,N_3257);
or U3492 (N_3492,N_3221,N_3243);
or U3493 (N_3493,N_3364,N_3285);
nand U3494 (N_3494,N_3238,N_3339);
xnor U3495 (N_3495,N_3362,N_3336);
nor U3496 (N_3496,N_3256,N_3379);
nor U3497 (N_3497,N_3208,N_3269);
nand U3498 (N_3498,N_3312,N_3323);
xnor U3499 (N_3499,N_3335,N_3317);
xnor U3500 (N_3500,N_3283,N_3223);
and U3501 (N_3501,N_3380,N_3351);
and U3502 (N_3502,N_3327,N_3392);
or U3503 (N_3503,N_3303,N_3344);
xor U3504 (N_3504,N_3282,N_3247);
or U3505 (N_3505,N_3284,N_3367);
and U3506 (N_3506,N_3370,N_3342);
nand U3507 (N_3507,N_3344,N_3293);
and U3508 (N_3508,N_3346,N_3230);
xnor U3509 (N_3509,N_3374,N_3384);
and U3510 (N_3510,N_3380,N_3303);
xnor U3511 (N_3511,N_3262,N_3264);
nor U3512 (N_3512,N_3390,N_3265);
nand U3513 (N_3513,N_3254,N_3275);
xnor U3514 (N_3514,N_3382,N_3356);
or U3515 (N_3515,N_3278,N_3230);
nor U3516 (N_3516,N_3397,N_3344);
nor U3517 (N_3517,N_3318,N_3235);
nor U3518 (N_3518,N_3336,N_3358);
or U3519 (N_3519,N_3243,N_3355);
or U3520 (N_3520,N_3380,N_3344);
nor U3521 (N_3521,N_3227,N_3286);
xnor U3522 (N_3522,N_3307,N_3309);
xnor U3523 (N_3523,N_3241,N_3258);
and U3524 (N_3524,N_3221,N_3241);
or U3525 (N_3525,N_3377,N_3232);
or U3526 (N_3526,N_3301,N_3201);
and U3527 (N_3527,N_3354,N_3378);
nor U3528 (N_3528,N_3335,N_3225);
xor U3529 (N_3529,N_3352,N_3382);
xor U3530 (N_3530,N_3208,N_3353);
nor U3531 (N_3531,N_3351,N_3213);
and U3532 (N_3532,N_3382,N_3284);
nor U3533 (N_3533,N_3204,N_3249);
and U3534 (N_3534,N_3281,N_3263);
xnor U3535 (N_3535,N_3356,N_3370);
or U3536 (N_3536,N_3308,N_3207);
nor U3537 (N_3537,N_3270,N_3222);
xor U3538 (N_3538,N_3310,N_3284);
xnor U3539 (N_3539,N_3357,N_3305);
xor U3540 (N_3540,N_3290,N_3394);
nand U3541 (N_3541,N_3371,N_3300);
xnor U3542 (N_3542,N_3289,N_3208);
or U3543 (N_3543,N_3236,N_3245);
xor U3544 (N_3544,N_3387,N_3259);
xnor U3545 (N_3545,N_3240,N_3203);
or U3546 (N_3546,N_3313,N_3353);
or U3547 (N_3547,N_3389,N_3268);
nor U3548 (N_3548,N_3306,N_3325);
or U3549 (N_3549,N_3360,N_3233);
nor U3550 (N_3550,N_3321,N_3278);
xnor U3551 (N_3551,N_3321,N_3244);
nor U3552 (N_3552,N_3232,N_3227);
nor U3553 (N_3553,N_3212,N_3288);
and U3554 (N_3554,N_3387,N_3222);
nor U3555 (N_3555,N_3323,N_3359);
or U3556 (N_3556,N_3390,N_3214);
nor U3557 (N_3557,N_3205,N_3305);
xnor U3558 (N_3558,N_3326,N_3386);
xnor U3559 (N_3559,N_3290,N_3329);
xor U3560 (N_3560,N_3379,N_3315);
xor U3561 (N_3561,N_3327,N_3256);
nand U3562 (N_3562,N_3314,N_3394);
nor U3563 (N_3563,N_3223,N_3390);
and U3564 (N_3564,N_3274,N_3238);
nand U3565 (N_3565,N_3262,N_3295);
or U3566 (N_3566,N_3310,N_3377);
xor U3567 (N_3567,N_3301,N_3250);
or U3568 (N_3568,N_3263,N_3364);
and U3569 (N_3569,N_3262,N_3376);
nand U3570 (N_3570,N_3387,N_3296);
nor U3571 (N_3571,N_3350,N_3325);
nor U3572 (N_3572,N_3232,N_3335);
nor U3573 (N_3573,N_3373,N_3283);
or U3574 (N_3574,N_3345,N_3202);
xnor U3575 (N_3575,N_3395,N_3340);
xor U3576 (N_3576,N_3336,N_3241);
xor U3577 (N_3577,N_3295,N_3217);
and U3578 (N_3578,N_3325,N_3210);
xnor U3579 (N_3579,N_3399,N_3237);
and U3580 (N_3580,N_3233,N_3319);
nand U3581 (N_3581,N_3327,N_3332);
or U3582 (N_3582,N_3369,N_3213);
nor U3583 (N_3583,N_3290,N_3291);
nand U3584 (N_3584,N_3272,N_3320);
xor U3585 (N_3585,N_3248,N_3380);
nor U3586 (N_3586,N_3396,N_3207);
xnor U3587 (N_3587,N_3241,N_3214);
nand U3588 (N_3588,N_3381,N_3313);
or U3589 (N_3589,N_3204,N_3239);
and U3590 (N_3590,N_3365,N_3343);
xor U3591 (N_3591,N_3234,N_3302);
nor U3592 (N_3592,N_3372,N_3384);
xnor U3593 (N_3593,N_3365,N_3337);
xor U3594 (N_3594,N_3327,N_3335);
and U3595 (N_3595,N_3345,N_3265);
or U3596 (N_3596,N_3368,N_3329);
or U3597 (N_3597,N_3217,N_3375);
xnor U3598 (N_3598,N_3297,N_3369);
xor U3599 (N_3599,N_3215,N_3370);
or U3600 (N_3600,N_3402,N_3439);
nand U3601 (N_3601,N_3546,N_3572);
and U3602 (N_3602,N_3500,N_3492);
nor U3603 (N_3603,N_3468,N_3537);
nand U3604 (N_3604,N_3476,N_3483);
or U3605 (N_3605,N_3542,N_3433);
and U3606 (N_3606,N_3455,N_3556);
nor U3607 (N_3607,N_3416,N_3449);
and U3608 (N_3608,N_3522,N_3495);
nor U3609 (N_3609,N_3502,N_3406);
xor U3610 (N_3610,N_3498,N_3504);
or U3611 (N_3611,N_3471,N_3530);
nand U3612 (N_3612,N_3536,N_3554);
nor U3613 (N_3613,N_3519,N_3539);
and U3614 (N_3614,N_3497,N_3426);
and U3615 (N_3615,N_3405,N_3501);
nor U3616 (N_3616,N_3525,N_3477);
nor U3617 (N_3617,N_3472,N_3538);
xnor U3618 (N_3618,N_3494,N_3496);
nand U3619 (N_3619,N_3430,N_3515);
and U3620 (N_3620,N_3568,N_3505);
or U3621 (N_3621,N_3541,N_3480);
or U3622 (N_3622,N_3548,N_3585);
nor U3623 (N_3623,N_3550,N_3418);
or U3624 (N_3624,N_3404,N_3493);
nand U3625 (N_3625,N_3532,N_3485);
or U3626 (N_3626,N_3429,N_3486);
and U3627 (N_3627,N_3436,N_3528);
xnor U3628 (N_3628,N_3407,N_3469);
nand U3629 (N_3629,N_3540,N_3591);
nand U3630 (N_3630,N_3558,N_3435);
and U3631 (N_3631,N_3434,N_3467);
xnor U3632 (N_3632,N_3456,N_3417);
nand U3633 (N_3633,N_3488,N_3578);
xnor U3634 (N_3634,N_3592,N_3461);
xnor U3635 (N_3635,N_3575,N_3589);
and U3636 (N_3636,N_3465,N_3574);
nor U3637 (N_3637,N_3441,N_3458);
xnor U3638 (N_3638,N_3450,N_3593);
nand U3639 (N_3639,N_3422,N_3424);
and U3640 (N_3640,N_3453,N_3508);
nor U3641 (N_3641,N_3503,N_3551);
or U3642 (N_3642,N_3527,N_3560);
and U3643 (N_3643,N_3466,N_3529);
nand U3644 (N_3644,N_3544,N_3577);
xor U3645 (N_3645,N_3506,N_3533);
or U3646 (N_3646,N_3526,N_3547);
and U3647 (N_3647,N_3470,N_3597);
xnor U3648 (N_3648,N_3510,N_3581);
or U3649 (N_3649,N_3516,N_3411);
xnor U3650 (N_3650,N_3576,N_3549);
and U3651 (N_3651,N_3473,N_3553);
or U3652 (N_3652,N_3415,N_3507);
nor U3653 (N_3653,N_3583,N_3440);
or U3654 (N_3654,N_3414,N_3552);
or U3655 (N_3655,N_3564,N_3535);
xnor U3656 (N_3656,N_3478,N_3484);
or U3657 (N_3657,N_3565,N_3587);
or U3658 (N_3658,N_3590,N_3409);
xnor U3659 (N_3659,N_3513,N_3517);
and U3660 (N_3660,N_3474,N_3566);
or U3661 (N_3661,N_3531,N_3445);
and U3662 (N_3662,N_3425,N_3448);
or U3663 (N_3663,N_3588,N_3462);
nand U3664 (N_3664,N_3569,N_3431);
nand U3665 (N_3665,N_3582,N_3584);
and U3666 (N_3666,N_3479,N_3571);
xor U3667 (N_3667,N_3490,N_3579);
and U3668 (N_3668,N_3447,N_3557);
and U3669 (N_3669,N_3487,N_3442);
and U3670 (N_3670,N_3460,N_3419);
and U3671 (N_3671,N_3412,N_3586);
and U3672 (N_3672,N_3401,N_3491);
nand U3673 (N_3673,N_3580,N_3443);
xor U3674 (N_3674,N_3410,N_3459);
nand U3675 (N_3675,N_3523,N_3559);
and U3676 (N_3676,N_3555,N_3423);
nor U3677 (N_3677,N_3432,N_3534);
xnor U3678 (N_3678,N_3545,N_3509);
nand U3679 (N_3679,N_3570,N_3514);
and U3680 (N_3680,N_3567,N_3428);
and U3681 (N_3681,N_3400,N_3518);
xor U3682 (N_3682,N_3454,N_3598);
xor U3683 (N_3683,N_3457,N_3499);
and U3684 (N_3684,N_3481,N_3446);
and U3685 (N_3685,N_3482,N_3427);
nor U3686 (N_3686,N_3438,N_3489);
or U3687 (N_3687,N_3420,N_3594);
nand U3688 (N_3688,N_3561,N_3563);
or U3689 (N_3689,N_3408,N_3512);
or U3690 (N_3690,N_3437,N_3596);
and U3691 (N_3691,N_3403,N_3599);
nor U3692 (N_3692,N_3520,N_3463);
nor U3693 (N_3693,N_3511,N_3451);
nand U3694 (N_3694,N_3444,N_3464);
and U3695 (N_3695,N_3521,N_3543);
xor U3696 (N_3696,N_3413,N_3524);
or U3697 (N_3697,N_3475,N_3562);
and U3698 (N_3698,N_3573,N_3595);
or U3699 (N_3699,N_3421,N_3452);
nand U3700 (N_3700,N_3557,N_3466);
xnor U3701 (N_3701,N_3460,N_3556);
or U3702 (N_3702,N_3496,N_3533);
nand U3703 (N_3703,N_3479,N_3410);
nor U3704 (N_3704,N_3523,N_3477);
and U3705 (N_3705,N_3526,N_3454);
and U3706 (N_3706,N_3426,N_3450);
and U3707 (N_3707,N_3474,N_3528);
and U3708 (N_3708,N_3561,N_3415);
nand U3709 (N_3709,N_3406,N_3413);
nor U3710 (N_3710,N_3555,N_3452);
and U3711 (N_3711,N_3526,N_3460);
nand U3712 (N_3712,N_3587,N_3477);
or U3713 (N_3713,N_3419,N_3420);
nor U3714 (N_3714,N_3598,N_3475);
and U3715 (N_3715,N_3549,N_3493);
or U3716 (N_3716,N_3435,N_3526);
and U3717 (N_3717,N_3468,N_3566);
nor U3718 (N_3718,N_3589,N_3484);
or U3719 (N_3719,N_3408,N_3496);
nand U3720 (N_3720,N_3531,N_3533);
xor U3721 (N_3721,N_3562,N_3445);
nor U3722 (N_3722,N_3508,N_3573);
nor U3723 (N_3723,N_3566,N_3462);
nand U3724 (N_3724,N_3544,N_3499);
xnor U3725 (N_3725,N_3435,N_3566);
nor U3726 (N_3726,N_3522,N_3405);
or U3727 (N_3727,N_3495,N_3559);
and U3728 (N_3728,N_3535,N_3498);
nor U3729 (N_3729,N_3431,N_3542);
xor U3730 (N_3730,N_3425,N_3429);
or U3731 (N_3731,N_3400,N_3448);
or U3732 (N_3732,N_3402,N_3401);
nor U3733 (N_3733,N_3507,N_3526);
nor U3734 (N_3734,N_3473,N_3409);
nor U3735 (N_3735,N_3458,N_3549);
nand U3736 (N_3736,N_3514,N_3568);
and U3737 (N_3737,N_3524,N_3526);
xnor U3738 (N_3738,N_3512,N_3414);
xor U3739 (N_3739,N_3469,N_3520);
and U3740 (N_3740,N_3581,N_3486);
nand U3741 (N_3741,N_3409,N_3504);
nor U3742 (N_3742,N_3469,N_3471);
nor U3743 (N_3743,N_3471,N_3543);
nor U3744 (N_3744,N_3433,N_3463);
or U3745 (N_3745,N_3464,N_3432);
xnor U3746 (N_3746,N_3400,N_3412);
or U3747 (N_3747,N_3466,N_3401);
nor U3748 (N_3748,N_3464,N_3437);
and U3749 (N_3749,N_3538,N_3400);
and U3750 (N_3750,N_3414,N_3571);
nor U3751 (N_3751,N_3488,N_3534);
or U3752 (N_3752,N_3556,N_3492);
nand U3753 (N_3753,N_3469,N_3470);
or U3754 (N_3754,N_3530,N_3482);
and U3755 (N_3755,N_3423,N_3458);
or U3756 (N_3756,N_3571,N_3443);
or U3757 (N_3757,N_3438,N_3576);
xnor U3758 (N_3758,N_3585,N_3583);
or U3759 (N_3759,N_3423,N_3480);
or U3760 (N_3760,N_3521,N_3580);
and U3761 (N_3761,N_3526,N_3573);
xor U3762 (N_3762,N_3468,N_3422);
nor U3763 (N_3763,N_3472,N_3528);
xnor U3764 (N_3764,N_3424,N_3585);
nand U3765 (N_3765,N_3433,N_3462);
xor U3766 (N_3766,N_3428,N_3519);
nor U3767 (N_3767,N_3442,N_3414);
nor U3768 (N_3768,N_3528,N_3500);
or U3769 (N_3769,N_3479,N_3427);
or U3770 (N_3770,N_3566,N_3443);
or U3771 (N_3771,N_3411,N_3587);
and U3772 (N_3772,N_3442,N_3569);
xnor U3773 (N_3773,N_3442,N_3424);
or U3774 (N_3774,N_3404,N_3556);
nand U3775 (N_3775,N_3568,N_3421);
and U3776 (N_3776,N_3567,N_3537);
nor U3777 (N_3777,N_3577,N_3479);
xnor U3778 (N_3778,N_3576,N_3448);
xor U3779 (N_3779,N_3470,N_3405);
nor U3780 (N_3780,N_3538,N_3412);
and U3781 (N_3781,N_3506,N_3565);
nand U3782 (N_3782,N_3527,N_3588);
xor U3783 (N_3783,N_3578,N_3533);
xor U3784 (N_3784,N_3591,N_3586);
nand U3785 (N_3785,N_3429,N_3475);
or U3786 (N_3786,N_3561,N_3556);
and U3787 (N_3787,N_3520,N_3448);
xnor U3788 (N_3788,N_3425,N_3540);
xnor U3789 (N_3789,N_3490,N_3533);
and U3790 (N_3790,N_3548,N_3570);
xnor U3791 (N_3791,N_3516,N_3551);
nand U3792 (N_3792,N_3517,N_3536);
or U3793 (N_3793,N_3574,N_3570);
or U3794 (N_3794,N_3483,N_3496);
xnor U3795 (N_3795,N_3418,N_3552);
and U3796 (N_3796,N_3467,N_3576);
nand U3797 (N_3797,N_3491,N_3563);
xor U3798 (N_3798,N_3500,N_3453);
and U3799 (N_3799,N_3429,N_3409);
or U3800 (N_3800,N_3720,N_3663);
or U3801 (N_3801,N_3760,N_3657);
or U3802 (N_3802,N_3776,N_3747);
xor U3803 (N_3803,N_3768,N_3717);
and U3804 (N_3804,N_3771,N_3721);
xor U3805 (N_3805,N_3614,N_3647);
or U3806 (N_3806,N_3687,N_3682);
nor U3807 (N_3807,N_3677,N_3696);
or U3808 (N_3808,N_3670,N_3659);
nand U3809 (N_3809,N_3683,N_3748);
nand U3810 (N_3810,N_3770,N_3788);
or U3811 (N_3811,N_3711,N_3627);
nor U3812 (N_3812,N_3634,N_3620);
and U3813 (N_3813,N_3666,N_3631);
nor U3814 (N_3814,N_3793,N_3654);
nand U3815 (N_3815,N_3616,N_3679);
nor U3816 (N_3816,N_3693,N_3727);
nand U3817 (N_3817,N_3678,N_3613);
nand U3818 (N_3818,N_3664,N_3769);
nand U3819 (N_3819,N_3705,N_3636);
and U3820 (N_3820,N_3629,N_3697);
or U3821 (N_3821,N_3645,N_3667);
xor U3822 (N_3822,N_3795,N_3798);
or U3823 (N_3823,N_3669,N_3623);
nand U3824 (N_3824,N_3619,N_3656);
or U3825 (N_3825,N_3751,N_3610);
and U3826 (N_3826,N_3780,N_3783);
nand U3827 (N_3827,N_3665,N_3655);
and U3828 (N_3828,N_3649,N_3699);
xnor U3829 (N_3829,N_3766,N_3733);
nand U3830 (N_3830,N_3618,N_3689);
nor U3831 (N_3831,N_3668,N_3648);
and U3832 (N_3832,N_3622,N_3764);
or U3833 (N_3833,N_3797,N_3672);
nor U3834 (N_3834,N_3782,N_3673);
nand U3835 (N_3835,N_3778,N_3617);
xor U3836 (N_3836,N_3671,N_3734);
nor U3837 (N_3837,N_3624,N_3713);
nand U3838 (N_3838,N_3730,N_3716);
nand U3839 (N_3839,N_3701,N_3792);
xor U3840 (N_3840,N_3628,N_3737);
or U3841 (N_3841,N_3741,N_3753);
nand U3842 (N_3842,N_3653,N_3743);
nor U3843 (N_3843,N_3725,N_3731);
nor U3844 (N_3844,N_3740,N_3691);
xnor U3845 (N_3845,N_3736,N_3643);
or U3846 (N_3846,N_3676,N_3723);
nand U3847 (N_3847,N_3763,N_3744);
nand U3848 (N_3848,N_3646,N_3715);
xnor U3849 (N_3849,N_3612,N_3794);
xnor U3850 (N_3850,N_3781,N_3718);
xnor U3851 (N_3851,N_3603,N_3785);
nand U3852 (N_3852,N_3692,N_3752);
and U3853 (N_3853,N_3735,N_3661);
xor U3854 (N_3854,N_3761,N_3680);
nor U3855 (N_3855,N_3660,N_3707);
and U3856 (N_3856,N_3704,N_3681);
and U3857 (N_3857,N_3708,N_3714);
nor U3858 (N_3858,N_3722,N_3605);
nand U3859 (N_3859,N_3652,N_3706);
nand U3860 (N_3860,N_3637,N_3772);
xnor U3861 (N_3861,N_3686,N_3710);
nand U3862 (N_3862,N_3675,N_3746);
nor U3863 (N_3863,N_3685,N_3719);
nand U3864 (N_3864,N_3602,N_3642);
nor U3865 (N_3865,N_3611,N_3674);
xnor U3866 (N_3866,N_3639,N_3688);
and U3867 (N_3867,N_3762,N_3742);
nor U3868 (N_3868,N_3786,N_3728);
nor U3869 (N_3869,N_3750,N_3774);
xnor U3870 (N_3870,N_3621,N_3626);
xor U3871 (N_3871,N_3745,N_3606);
and U3872 (N_3872,N_3630,N_3767);
nor U3873 (N_3873,N_3791,N_3601);
nor U3874 (N_3874,N_3695,N_3758);
and U3875 (N_3875,N_3690,N_3651);
and U3876 (N_3876,N_3739,N_3600);
nor U3877 (N_3877,N_3609,N_3738);
nand U3878 (N_3878,N_3755,N_3702);
or U3879 (N_3879,N_3724,N_3644);
nand U3880 (N_3880,N_3726,N_3635);
or U3881 (N_3881,N_3604,N_3633);
and U3882 (N_3882,N_3773,N_3796);
xor U3883 (N_3883,N_3698,N_3759);
xnor U3884 (N_3884,N_3615,N_3756);
xor U3885 (N_3885,N_3754,N_3625);
nor U3886 (N_3886,N_3638,N_3650);
or U3887 (N_3887,N_3775,N_3732);
xnor U3888 (N_3888,N_3607,N_3694);
nor U3889 (N_3889,N_3779,N_3777);
nor U3890 (N_3890,N_3789,N_3662);
xnor U3891 (N_3891,N_3765,N_3658);
and U3892 (N_3892,N_3790,N_3684);
and U3893 (N_3893,N_3787,N_3799);
nor U3894 (N_3894,N_3709,N_3749);
xnor U3895 (N_3895,N_3784,N_3757);
xnor U3896 (N_3896,N_3640,N_3703);
or U3897 (N_3897,N_3700,N_3641);
xnor U3898 (N_3898,N_3632,N_3712);
or U3899 (N_3899,N_3729,N_3608);
or U3900 (N_3900,N_3638,N_3726);
nor U3901 (N_3901,N_3637,N_3622);
or U3902 (N_3902,N_3620,N_3684);
and U3903 (N_3903,N_3680,N_3655);
xnor U3904 (N_3904,N_3637,N_3720);
nor U3905 (N_3905,N_3709,N_3664);
xnor U3906 (N_3906,N_3691,N_3675);
or U3907 (N_3907,N_3770,N_3631);
xnor U3908 (N_3908,N_3604,N_3671);
nor U3909 (N_3909,N_3690,N_3757);
nand U3910 (N_3910,N_3718,N_3771);
xor U3911 (N_3911,N_3750,N_3678);
and U3912 (N_3912,N_3747,N_3798);
nor U3913 (N_3913,N_3693,N_3679);
nand U3914 (N_3914,N_3661,N_3702);
and U3915 (N_3915,N_3755,N_3660);
nand U3916 (N_3916,N_3677,N_3638);
or U3917 (N_3917,N_3791,N_3661);
xnor U3918 (N_3918,N_3645,N_3625);
or U3919 (N_3919,N_3707,N_3745);
nor U3920 (N_3920,N_3669,N_3611);
nor U3921 (N_3921,N_3776,N_3637);
nand U3922 (N_3922,N_3761,N_3708);
xnor U3923 (N_3923,N_3790,N_3745);
or U3924 (N_3924,N_3650,N_3619);
or U3925 (N_3925,N_3645,N_3602);
and U3926 (N_3926,N_3682,N_3621);
nand U3927 (N_3927,N_3680,N_3674);
or U3928 (N_3928,N_3792,N_3750);
or U3929 (N_3929,N_3795,N_3650);
nor U3930 (N_3930,N_3762,N_3654);
xnor U3931 (N_3931,N_3742,N_3614);
nor U3932 (N_3932,N_3615,N_3614);
nand U3933 (N_3933,N_3638,N_3633);
xnor U3934 (N_3934,N_3692,N_3713);
nand U3935 (N_3935,N_3617,N_3672);
nand U3936 (N_3936,N_3657,N_3719);
and U3937 (N_3937,N_3784,N_3782);
xnor U3938 (N_3938,N_3621,N_3654);
or U3939 (N_3939,N_3643,N_3760);
nor U3940 (N_3940,N_3705,N_3763);
and U3941 (N_3941,N_3665,N_3768);
nand U3942 (N_3942,N_3654,N_3752);
xor U3943 (N_3943,N_3620,N_3683);
nor U3944 (N_3944,N_3724,N_3777);
xnor U3945 (N_3945,N_3699,N_3643);
or U3946 (N_3946,N_3748,N_3774);
or U3947 (N_3947,N_3605,N_3607);
nor U3948 (N_3948,N_3633,N_3632);
xnor U3949 (N_3949,N_3714,N_3770);
xor U3950 (N_3950,N_3614,N_3674);
xnor U3951 (N_3951,N_3796,N_3666);
nor U3952 (N_3952,N_3781,N_3684);
nor U3953 (N_3953,N_3676,N_3644);
nor U3954 (N_3954,N_3788,N_3637);
and U3955 (N_3955,N_3786,N_3629);
xor U3956 (N_3956,N_3793,N_3602);
nor U3957 (N_3957,N_3620,N_3628);
nand U3958 (N_3958,N_3751,N_3722);
xor U3959 (N_3959,N_3614,N_3734);
xnor U3960 (N_3960,N_3776,N_3741);
and U3961 (N_3961,N_3774,N_3777);
and U3962 (N_3962,N_3659,N_3673);
and U3963 (N_3963,N_3608,N_3735);
or U3964 (N_3964,N_3606,N_3643);
or U3965 (N_3965,N_3783,N_3724);
nor U3966 (N_3966,N_3759,N_3731);
nand U3967 (N_3967,N_3659,N_3617);
nor U3968 (N_3968,N_3631,N_3691);
xnor U3969 (N_3969,N_3609,N_3786);
nor U3970 (N_3970,N_3647,N_3702);
nor U3971 (N_3971,N_3794,N_3618);
and U3972 (N_3972,N_3678,N_3789);
and U3973 (N_3973,N_3726,N_3762);
nor U3974 (N_3974,N_3717,N_3755);
nand U3975 (N_3975,N_3691,N_3730);
or U3976 (N_3976,N_3650,N_3786);
or U3977 (N_3977,N_3767,N_3658);
xnor U3978 (N_3978,N_3701,N_3685);
or U3979 (N_3979,N_3689,N_3739);
and U3980 (N_3980,N_3603,N_3663);
or U3981 (N_3981,N_3646,N_3732);
nand U3982 (N_3982,N_3708,N_3757);
nand U3983 (N_3983,N_3619,N_3645);
and U3984 (N_3984,N_3663,N_3617);
xnor U3985 (N_3985,N_3660,N_3737);
nand U3986 (N_3986,N_3741,N_3757);
nand U3987 (N_3987,N_3760,N_3611);
or U3988 (N_3988,N_3651,N_3692);
nand U3989 (N_3989,N_3662,N_3644);
xnor U3990 (N_3990,N_3664,N_3663);
nor U3991 (N_3991,N_3655,N_3726);
nand U3992 (N_3992,N_3689,N_3667);
nor U3993 (N_3993,N_3738,N_3698);
or U3994 (N_3994,N_3622,N_3768);
nor U3995 (N_3995,N_3671,N_3771);
and U3996 (N_3996,N_3704,N_3753);
xnor U3997 (N_3997,N_3710,N_3799);
or U3998 (N_3998,N_3683,N_3762);
nor U3999 (N_3999,N_3658,N_3773);
or U4000 (N_4000,N_3876,N_3831);
or U4001 (N_4001,N_3962,N_3971);
and U4002 (N_4002,N_3823,N_3809);
or U4003 (N_4003,N_3916,N_3917);
and U4004 (N_4004,N_3841,N_3848);
or U4005 (N_4005,N_3896,N_3897);
nand U4006 (N_4006,N_3838,N_3937);
nand U4007 (N_4007,N_3961,N_3981);
xor U4008 (N_4008,N_3909,N_3949);
nor U4009 (N_4009,N_3807,N_3965);
or U4010 (N_4010,N_3969,N_3998);
and U4011 (N_4011,N_3936,N_3834);
xnor U4012 (N_4012,N_3932,N_3846);
nor U4013 (N_4013,N_3927,N_3803);
and U4014 (N_4014,N_3999,N_3817);
nor U4015 (N_4015,N_3914,N_3968);
or U4016 (N_4016,N_3913,N_3910);
nand U4017 (N_4017,N_3825,N_3938);
nor U4018 (N_4018,N_3901,N_3811);
and U4019 (N_4019,N_3862,N_3947);
xor U4020 (N_4020,N_3833,N_3902);
nor U4021 (N_4021,N_3898,N_3921);
xor U4022 (N_4022,N_3855,N_3836);
nand U4023 (N_4023,N_3959,N_3864);
nand U4024 (N_4024,N_3824,N_3943);
or U4025 (N_4025,N_3985,N_3977);
xnor U4026 (N_4026,N_3960,N_3890);
nand U4027 (N_4027,N_3858,N_3857);
or U4028 (N_4028,N_3972,N_3993);
xor U4029 (N_4029,N_3839,N_3870);
and U4030 (N_4030,N_3859,N_3970);
nand U4031 (N_4031,N_3941,N_3801);
and U4032 (N_4032,N_3905,N_3919);
nor U4033 (N_4033,N_3950,N_3895);
nand U4034 (N_4034,N_3966,N_3991);
or U4035 (N_4035,N_3967,N_3874);
nor U4036 (N_4036,N_3854,N_3875);
and U4037 (N_4037,N_3946,N_3948);
nand U4038 (N_4038,N_3812,N_3860);
xor U4039 (N_4039,N_3877,N_3867);
or U4040 (N_4040,N_3982,N_3911);
and U4041 (N_4041,N_3815,N_3879);
xnor U4042 (N_4042,N_3851,N_3926);
or U4043 (N_4043,N_3872,N_3931);
nor U4044 (N_4044,N_3954,N_3878);
or U4045 (N_4045,N_3808,N_3845);
nor U4046 (N_4046,N_3849,N_3853);
xor U4047 (N_4047,N_3928,N_3802);
nand U4048 (N_4048,N_3847,N_3925);
nand U4049 (N_4049,N_3816,N_3918);
xnor U4050 (N_4050,N_3976,N_3933);
nor U4051 (N_4051,N_3994,N_3873);
xor U4052 (N_4052,N_3881,N_3829);
nor U4053 (N_4053,N_3983,N_3894);
or U4054 (N_4054,N_3893,N_3830);
nand U4055 (N_4055,N_3863,N_3904);
nand U4056 (N_4056,N_3978,N_3922);
nor U4057 (N_4057,N_3889,N_3804);
and U4058 (N_4058,N_3975,N_3819);
xor U4059 (N_4059,N_3996,N_3835);
and U4060 (N_4060,N_3930,N_3837);
nor U4061 (N_4061,N_3821,N_3852);
and U4062 (N_4062,N_3887,N_3886);
or U4063 (N_4063,N_3974,N_3832);
nor U4064 (N_4064,N_3842,N_3843);
or U4065 (N_4065,N_3944,N_3912);
xor U4066 (N_4066,N_3953,N_3888);
and U4067 (N_4067,N_3973,N_3814);
nor U4068 (N_4068,N_3956,N_3957);
nor U4069 (N_4069,N_3891,N_3868);
nor U4070 (N_4070,N_3906,N_3892);
or U4071 (N_4071,N_3923,N_3987);
nor U4072 (N_4072,N_3856,N_3884);
nand U4073 (N_4073,N_3865,N_3979);
nand U4074 (N_4074,N_3951,N_3984);
nor U4075 (N_4075,N_3900,N_3997);
nor U4076 (N_4076,N_3882,N_3958);
nand U4077 (N_4077,N_3939,N_3840);
nor U4078 (N_4078,N_3963,N_3903);
or U4079 (N_4079,N_3942,N_3915);
or U4080 (N_4080,N_3990,N_3940);
or U4081 (N_4081,N_3866,N_3805);
xnor U4082 (N_4082,N_3964,N_3820);
or U4083 (N_4083,N_3934,N_3980);
xnor U4084 (N_4084,N_3899,N_3800);
nor U4085 (N_4085,N_3861,N_3813);
or U4086 (N_4086,N_3935,N_3920);
nand U4087 (N_4087,N_3885,N_3986);
nand U4088 (N_4088,N_3924,N_3908);
nor U4089 (N_4089,N_3871,N_3826);
and U4090 (N_4090,N_3822,N_3995);
xnor U4091 (N_4091,N_3989,N_3880);
nor U4092 (N_4092,N_3945,N_3929);
and U4093 (N_4093,N_3844,N_3827);
nand U4094 (N_4094,N_3850,N_3883);
nor U4095 (N_4095,N_3818,N_3869);
and U4096 (N_4096,N_3810,N_3907);
nand U4097 (N_4097,N_3955,N_3828);
and U4098 (N_4098,N_3988,N_3806);
xor U4099 (N_4099,N_3952,N_3992);
nand U4100 (N_4100,N_3971,N_3955);
nor U4101 (N_4101,N_3908,N_3931);
nand U4102 (N_4102,N_3941,N_3828);
or U4103 (N_4103,N_3900,N_3879);
or U4104 (N_4104,N_3962,N_3813);
nor U4105 (N_4105,N_3810,N_3857);
xnor U4106 (N_4106,N_3867,N_3876);
and U4107 (N_4107,N_3914,N_3928);
and U4108 (N_4108,N_3994,N_3808);
nor U4109 (N_4109,N_3872,N_3917);
nand U4110 (N_4110,N_3812,N_3902);
and U4111 (N_4111,N_3875,N_3958);
and U4112 (N_4112,N_3960,N_3857);
and U4113 (N_4113,N_3937,N_3806);
or U4114 (N_4114,N_3973,N_3991);
xor U4115 (N_4115,N_3928,N_3983);
nor U4116 (N_4116,N_3849,N_3990);
or U4117 (N_4117,N_3905,N_3944);
or U4118 (N_4118,N_3918,N_3847);
xnor U4119 (N_4119,N_3866,N_3916);
or U4120 (N_4120,N_3819,N_3876);
and U4121 (N_4121,N_3856,N_3804);
or U4122 (N_4122,N_3811,N_3817);
and U4123 (N_4123,N_3874,N_3979);
xnor U4124 (N_4124,N_3910,N_3911);
nor U4125 (N_4125,N_3976,N_3907);
nor U4126 (N_4126,N_3910,N_3866);
nand U4127 (N_4127,N_3820,N_3919);
or U4128 (N_4128,N_3993,N_3988);
and U4129 (N_4129,N_3851,N_3927);
nor U4130 (N_4130,N_3825,N_3928);
xor U4131 (N_4131,N_3816,N_3864);
and U4132 (N_4132,N_3875,N_3909);
xor U4133 (N_4133,N_3816,N_3965);
or U4134 (N_4134,N_3858,N_3828);
or U4135 (N_4135,N_3828,N_3908);
nand U4136 (N_4136,N_3905,N_3942);
nor U4137 (N_4137,N_3984,N_3889);
nand U4138 (N_4138,N_3812,N_3994);
or U4139 (N_4139,N_3987,N_3830);
and U4140 (N_4140,N_3834,N_3937);
nand U4141 (N_4141,N_3876,N_3843);
nor U4142 (N_4142,N_3871,N_3851);
nor U4143 (N_4143,N_3810,N_3944);
xor U4144 (N_4144,N_3994,N_3939);
xor U4145 (N_4145,N_3942,N_3958);
xor U4146 (N_4146,N_3968,N_3810);
and U4147 (N_4147,N_3845,N_3950);
xnor U4148 (N_4148,N_3804,N_3906);
xor U4149 (N_4149,N_3870,N_3828);
nor U4150 (N_4150,N_3985,N_3861);
nor U4151 (N_4151,N_3918,N_3997);
xor U4152 (N_4152,N_3887,N_3870);
xnor U4153 (N_4153,N_3938,N_3976);
nor U4154 (N_4154,N_3964,N_3944);
xor U4155 (N_4155,N_3839,N_3947);
nand U4156 (N_4156,N_3803,N_3907);
or U4157 (N_4157,N_3988,N_3825);
and U4158 (N_4158,N_3986,N_3872);
and U4159 (N_4159,N_3931,N_3823);
and U4160 (N_4160,N_3828,N_3976);
nand U4161 (N_4161,N_3964,N_3960);
nand U4162 (N_4162,N_3959,N_3851);
or U4163 (N_4163,N_3930,N_3903);
nor U4164 (N_4164,N_3909,N_3878);
nor U4165 (N_4165,N_3800,N_3894);
or U4166 (N_4166,N_3933,N_3975);
and U4167 (N_4167,N_3909,N_3910);
nor U4168 (N_4168,N_3961,N_3838);
or U4169 (N_4169,N_3997,N_3829);
xnor U4170 (N_4170,N_3830,N_3819);
xor U4171 (N_4171,N_3960,N_3953);
nand U4172 (N_4172,N_3987,N_3949);
or U4173 (N_4173,N_3813,N_3832);
nand U4174 (N_4174,N_3844,N_3975);
nand U4175 (N_4175,N_3871,N_3901);
xnor U4176 (N_4176,N_3835,N_3970);
or U4177 (N_4177,N_3973,N_3859);
and U4178 (N_4178,N_3957,N_3903);
and U4179 (N_4179,N_3887,N_3960);
nand U4180 (N_4180,N_3841,N_3941);
or U4181 (N_4181,N_3830,N_3936);
xor U4182 (N_4182,N_3960,N_3904);
and U4183 (N_4183,N_3975,N_3840);
and U4184 (N_4184,N_3953,N_3878);
nor U4185 (N_4185,N_3933,N_3998);
nand U4186 (N_4186,N_3845,N_3931);
or U4187 (N_4187,N_3987,N_3808);
nor U4188 (N_4188,N_3876,N_3863);
and U4189 (N_4189,N_3810,N_3929);
or U4190 (N_4190,N_3874,N_3873);
and U4191 (N_4191,N_3852,N_3949);
or U4192 (N_4192,N_3991,N_3933);
nor U4193 (N_4193,N_3874,N_3847);
xnor U4194 (N_4194,N_3853,N_3909);
xnor U4195 (N_4195,N_3884,N_3860);
nand U4196 (N_4196,N_3933,N_3851);
nor U4197 (N_4197,N_3899,N_3904);
xor U4198 (N_4198,N_3972,N_3877);
xor U4199 (N_4199,N_3830,N_3829);
or U4200 (N_4200,N_4076,N_4160);
xnor U4201 (N_4201,N_4174,N_4077);
or U4202 (N_4202,N_4082,N_4086);
and U4203 (N_4203,N_4012,N_4090);
and U4204 (N_4204,N_4168,N_4070);
xor U4205 (N_4205,N_4198,N_4091);
xnor U4206 (N_4206,N_4135,N_4154);
nor U4207 (N_4207,N_4013,N_4105);
nand U4208 (N_4208,N_4148,N_4040);
nand U4209 (N_4209,N_4062,N_4099);
xor U4210 (N_4210,N_4145,N_4189);
nand U4211 (N_4211,N_4184,N_4152);
nand U4212 (N_4212,N_4030,N_4196);
nor U4213 (N_4213,N_4016,N_4022);
or U4214 (N_4214,N_4035,N_4142);
xor U4215 (N_4215,N_4151,N_4079);
nand U4216 (N_4216,N_4129,N_4038);
or U4217 (N_4217,N_4139,N_4185);
and U4218 (N_4218,N_4072,N_4109);
or U4219 (N_4219,N_4164,N_4102);
xnor U4220 (N_4220,N_4060,N_4195);
nand U4221 (N_4221,N_4118,N_4071);
and U4222 (N_4222,N_4114,N_4179);
nor U4223 (N_4223,N_4026,N_4113);
xnor U4224 (N_4224,N_4094,N_4008);
nand U4225 (N_4225,N_4044,N_4107);
and U4226 (N_4226,N_4052,N_4036);
nor U4227 (N_4227,N_4178,N_4047);
nand U4228 (N_4228,N_4192,N_4006);
xnor U4229 (N_4229,N_4033,N_4001);
and U4230 (N_4230,N_4123,N_4059);
and U4231 (N_4231,N_4138,N_4180);
xnor U4232 (N_4232,N_4015,N_4106);
and U4233 (N_4233,N_4023,N_4014);
and U4234 (N_4234,N_4081,N_4197);
and U4235 (N_4235,N_4067,N_4009);
or U4236 (N_4236,N_4149,N_4066);
or U4237 (N_4237,N_4084,N_4085);
nand U4238 (N_4238,N_4005,N_4078);
xor U4239 (N_4239,N_4055,N_4186);
xor U4240 (N_4240,N_4157,N_4173);
nor U4241 (N_4241,N_4125,N_4108);
xnor U4242 (N_4242,N_4183,N_4159);
nor U4243 (N_4243,N_4115,N_4046);
nor U4244 (N_4244,N_4092,N_4171);
nor U4245 (N_4245,N_4073,N_4063);
and U4246 (N_4246,N_4111,N_4188);
or U4247 (N_4247,N_4025,N_4193);
or U4248 (N_4248,N_4065,N_4032);
nor U4249 (N_4249,N_4019,N_4042);
nor U4250 (N_4250,N_4098,N_4034);
and U4251 (N_4251,N_4083,N_4068);
or U4252 (N_4252,N_4002,N_4000);
nand U4253 (N_4253,N_4147,N_4003);
xnor U4254 (N_4254,N_4136,N_4161);
or U4255 (N_4255,N_4037,N_4130);
nor U4256 (N_4256,N_4170,N_4163);
and U4257 (N_4257,N_4177,N_4069);
and U4258 (N_4258,N_4112,N_4051);
nor U4259 (N_4259,N_4004,N_4126);
xor U4260 (N_4260,N_4156,N_4080);
or U4261 (N_4261,N_4074,N_4144);
nand U4262 (N_4262,N_4028,N_4120);
and U4263 (N_4263,N_4117,N_4191);
nand U4264 (N_4264,N_4021,N_4121);
nor U4265 (N_4265,N_4061,N_4140);
xor U4266 (N_4266,N_4043,N_4155);
nor U4267 (N_4267,N_4095,N_4064);
and U4268 (N_4268,N_4049,N_4176);
nand U4269 (N_4269,N_4075,N_4187);
nor U4270 (N_4270,N_4050,N_4131);
nor U4271 (N_4271,N_4018,N_4190);
or U4272 (N_4272,N_4045,N_4169);
and U4273 (N_4273,N_4089,N_4143);
and U4274 (N_4274,N_4011,N_4141);
xor U4275 (N_4275,N_4039,N_4132);
or U4276 (N_4276,N_4020,N_4182);
or U4277 (N_4277,N_4017,N_4087);
and U4278 (N_4278,N_4024,N_4133);
nand U4279 (N_4279,N_4127,N_4134);
or U4280 (N_4280,N_4057,N_4054);
xor U4281 (N_4281,N_4181,N_4010);
or U4282 (N_4282,N_4175,N_4146);
nor U4283 (N_4283,N_4041,N_4150);
xnor U4284 (N_4284,N_4167,N_4031);
nor U4285 (N_4285,N_4166,N_4048);
or U4286 (N_4286,N_4007,N_4110);
nand U4287 (N_4287,N_4101,N_4104);
xnor U4288 (N_4288,N_4119,N_4097);
xor U4289 (N_4289,N_4165,N_4100);
xor U4290 (N_4290,N_4162,N_4058);
xor U4291 (N_4291,N_4027,N_4172);
and U4292 (N_4292,N_4128,N_4093);
xor U4293 (N_4293,N_4029,N_4199);
nor U4294 (N_4294,N_4137,N_4122);
xnor U4295 (N_4295,N_4158,N_4096);
and U4296 (N_4296,N_4088,N_4124);
xnor U4297 (N_4297,N_4053,N_4116);
xor U4298 (N_4298,N_4153,N_4056);
and U4299 (N_4299,N_4194,N_4103);
nor U4300 (N_4300,N_4033,N_4088);
nor U4301 (N_4301,N_4115,N_4090);
xor U4302 (N_4302,N_4163,N_4087);
nand U4303 (N_4303,N_4162,N_4105);
nand U4304 (N_4304,N_4159,N_4154);
nand U4305 (N_4305,N_4176,N_4061);
nand U4306 (N_4306,N_4059,N_4099);
nand U4307 (N_4307,N_4179,N_4083);
xor U4308 (N_4308,N_4189,N_4096);
nor U4309 (N_4309,N_4175,N_4081);
or U4310 (N_4310,N_4089,N_4068);
or U4311 (N_4311,N_4025,N_4114);
and U4312 (N_4312,N_4094,N_4042);
nand U4313 (N_4313,N_4007,N_4160);
nand U4314 (N_4314,N_4139,N_4026);
nor U4315 (N_4315,N_4141,N_4044);
and U4316 (N_4316,N_4022,N_4182);
nand U4317 (N_4317,N_4135,N_4156);
and U4318 (N_4318,N_4141,N_4036);
and U4319 (N_4319,N_4105,N_4046);
nand U4320 (N_4320,N_4176,N_4136);
or U4321 (N_4321,N_4024,N_4054);
or U4322 (N_4322,N_4037,N_4094);
xor U4323 (N_4323,N_4078,N_4128);
xor U4324 (N_4324,N_4038,N_4095);
xnor U4325 (N_4325,N_4084,N_4185);
and U4326 (N_4326,N_4178,N_4036);
xnor U4327 (N_4327,N_4083,N_4064);
nor U4328 (N_4328,N_4166,N_4093);
and U4329 (N_4329,N_4166,N_4012);
nor U4330 (N_4330,N_4191,N_4198);
and U4331 (N_4331,N_4147,N_4188);
or U4332 (N_4332,N_4065,N_4093);
nor U4333 (N_4333,N_4085,N_4148);
and U4334 (N_4334,N_4127,N_4088);
nand U4335 (N_4335,N_4010,N_4043);
nand U4336 (N_4336,N_4042,N_4095);
nor U4337 (N_4337,N_4154,N_4140);
or U4338 (N_4338,N_4053,N_4137);
or U4339 (N_4339,N_4164,N_4031);
xor U4340 (N_4340,N_4058,N_4167);
xor U4341 (N_4341,N_4036,N_4185);
nand U4342 (N_4342,N_4181,N_4129);
and U4343 (N_4343,N_4156,N_4072);
nand U4344 (N_4344,N_4143,N_4074);
xor U4345 (N_4345,N_4087,N_4060);
and U4346 (N_4346,N_4120,N_4129);
xnor U4347 (N_4347,N_4088,N_4094);
and U4348 (N_4348,N_4011,N_4030);
nand U4349 (N_4349,N_4077,N_4133);
nor U4350 (N_4350,N_4111,N_4102);
and U4351 (N_4351,N_4139,N_4010);
and U4352 (N_4352,N_4068,N_4032);
nand U4353 (N_4353,N_4096,N_4137);
or U4354 (N_4354,N_4022,N_4092);
nor U4355 (N_4355,N_4178,N_4056);
nor U4356 (N_4356,N_4190,N_4037);
nand U4357 (N_4357,N_4131,N_4103);
xor U4358 (N_4358,N_4184,N_4056);
nand U4359 (N_4359,N_4005,N_4126);
xnor U4360 (N_4360,N_4158,N_4162);
nor U4361 (N_4361,N_4082,N_4161);
and U4362 (N_4362,N_4053,N_4199);
nand U4363 (N_4363,N_4002,N_4041);
or U4364 (N_4364,N_4053,N_4170);
nor U4365 (N_4365,N_4181,N_4127);
nand U4366 (N_4366,N_4097,N_4009);
or U4367 (N_4367,N_4027,N_4147);
or U4368 (N_4368,N_4053,N_4070);
nor U4369 (N_4369,N_4058,N_4066);
or U4370 (N_4370,N_4151,N_4045);
or U4371 (N_4371,N_4153,N_4032);
nor U4372 (N_4372,N_4157,N_4016);
nand U4373 (N_4373,N_4145,N_4199);
xor U4374 (N_4374,N_4106,N_4175);
and U4375 (N_4375,N_4129,N_4114);
nor U4376 (N_4376,N_4037,N_4187);
or U4377 (N_4377,N_4150,N_4159);
nor U4378 (N_4378,N_4077,N_4123);
or U4379 (N_4379,N_4030,N_4155);
nand U4380 (N_4380,N_4061,N_4086);
nor U4381 (N_4381,N_4066,N_4062);
xor U4382 (N_4382,N_4150,N_4104);
xor U4383 (N_4383,N_4052,N_4024);
xor U4384 (N_4384,N_4018,N_4068);
or U4385 (N_4385,N_4103,N_4164);
nor U4386 (N_4386,N_4048,N_4102);
nand U4387 (N_4387,N_4034,N_4130);
and U4388 (N_4388,N_4031,N_4106);
nor U4389 (N_4389,N_4150,N_4116);
and U4390 (N_4390,N_4153,N_4094);
and U4391 (N_4391,N_4015,N_4059);
xnor U4392 (N_4392,N_4049,N_4147);
xnor U4393 (N_4393,N_4014,N_4173);
or U4394 (N_4394,N_4195,N_4168);
and U4395 (N_4395,N_4044,N_4015);
nor U4396 (N_4396,N_4075,N_4006);
nand U4397 (N_4397,N_4007,N_4064);
nor U4398 (N_4398,N_4073,N_4103);
or U4399 (N_4399,N_4026,N_4185);
or U4400 (N_4400,N_4213,N_4235);
and U4401 (N_4401,N_4324,N_4238);
and U4402 (N_4402,N_4313,N_4248);
or U4403 (N_4403,N_4363,N_4371);
nor U4404 (N_4404,N_4201,N_4279);
xor U4405 (N_4405,N_4252,N_4267);
nand U4406 (N_4406,N_4207,N_4341);
xnor U4407 (N_4407,N_4342,N_4387);
xor U4408 (N_4408,N_4291,N_4242);
and U4409 (N_4409,N_4268,N_4228);
nand U4410 (N_4410,N_4224,N_4237);
nand U4411 (N_4411,N_4368,N_4384);
and U4412 (N_4412,N_4359,N_4318);
and U4413 (N_4413,N_4326,N_4250);
nor U4414 (N_4414,N_4397,N_4353);
nand U4415 (N_4415,N_4280,N_4394);
xor U4416 (N_4416,N_4203,N_4240);
xnor U4417 (N_4417,N_4358,N_4361);
xnor U4418 (N_4418,N_4275,N_4278);
or U4419 (N_4419,N_4297,N_4222);
nor U4420 (N_4420,N_4225,N_4316);
nor U4421 (N_4421,N_4343,N_4276);
xor U4422 (N_4422,N_4393,N_4200);
xor U4423 (N_4423,N_4372,N_4236);
or U4424 (N_4424,N_4391,N_4390);
or U4425 (N_4425,N_4241,N_4344);
nor U4426 (N_4426,N_4328,N_4334);
nand U4427 (N_4427,N_4348,N_4255);
and U4428 (N_4428,N_4367,N_4263);
or U4429 (N_4429,N_4266,N_4307);
nor U4430 (N_4430,N_4293,N_4383);
xnor U4431 (N_4431,N_4281,N_4260);
and U4432 (N_4432,N_4232,N_4253);
and U4433 (N_4433,N_4345,N_4249);
nand U4434 (N_4434,N_4336,N_4277);
and U4435 (N_4435,N_4375,N_4323);
or U4436 (N_4436,N_4381,N_4369);
or U4437 (N_4437,N_4327,N_4306);
nand U4438 (N_4438,N_4305,N_4205);
and U4439 (N_4439,N_4239,N_4354);
nor U4440 (N_4440,N_4206,N_4287);
nand U4441 (N_4441,N_4243,N_4271);
nand U4442 (N_4442,N_4370,N_4218);
and U4443 (N_4443,N_4220,N_4364);
nor U4444 (N_4444,N_4294,N_4284);
nor U4445 (N_4445,N_4265,N_4246);
xor U4446 (N_4446,N_4398,N_4319);
nor U4447 (N_4447,N_4292,N_4380);
nand U4448 (N_4448,N_4322,N_4295);
nand U4449 (N_4449,N_4216,N_4215);
or U4450 (N_4450,N_4204,N_4312);
or U4451 (N_4451,N_4258,N_4310);
nor U4452 (N_4452,N_4233,N_4352);
and U4453 (N_4453,N_4365,N_4303);
and U4454 (N_4454,N_4325,N_4257);
nor U4455 (N_4455,N_4379,N_4308);
or U4456 (N_4456,N_4320,N_4209);
xor U4457 (N_4457,N_4234,N_4332);
nor U4458 (N_4458,N_4301,N_4347);
or U4459 (N_4459,N_4360,N_4273);
and U4460 (N_4460,N_4299,N_4335);
nor U4461 (N_4461,N_4286,N_4357);
or U4462 (N_4462,N_4356,N_4210);
nor U4463 (N_4463,N_4374,N_4392);
or U4464 (N_4464,N_4270,N_4389);
xnor U4465 (N_4465,N_4282,N_4315);
and U4466 (N_4466,N_4385,N_4283);
nand U4467 (N_4467,N_4254,N_4256);
nor U4468 (N_4468,N_4288,N_4377);
nor U4469 (N_4469,N_4382,N_4355);
or U4470 (N_4470,N_4349,N_4376);
nand U4471 (N_4471,N_4211,N_4223);
or U4472 (N_4472,N_4373,N_4226);
xnor U4473 (N_4473,N_4378,N_4314);
and U4474 (N_4474,N_4366,N_4396);
nand U4475 (N_4475,N_4289,N_4330);
or U4476 (N_4476,N_4296,N_4244);
xor U4477 (N_4477,N_4350,N_4227);
nor U4478 (N_4478,N_4264,N_4338);
and U4479 (N_4479,N_4269,N_4311);
and U4480 (N_4480,N_4300,N_4229);
or U4481 (N_4481,N_4231,N_4219);
nand U4482 (N_4482,N_4386,N_4362);
nor U4483 (N_4483,N_4339,N_4214);
or U4484 (N_4484,N_4208,N_4259);
nor U4485 (N_4485,N_4321,N_4395);
or U4486 (N_4486,N_4285,N_4247);
nand U4487 (N_4487,N_4212,N_4333);
or U4488 (N_4488,N_4262,N_4298);
and U4489 (N_4489,N_4340,N_4317);
or U4490 (N_4490,N_4221,N_4245);
or U4491 (N_4491,N_4304,N_4309);
nor U4492 (N_4492,N_4331,N_4230);
and U4493 (N_4493,N_4346,N_4251);
xnor U4494 (N_4494,N_4337,N_4399);
nand U4495 (N_4495,N_4202,N_4388);
nor U4496 (N_4496,N_4351,N_4217);
nand U4497 (N_4497,N_4272,N_4290);
xnor U4498 (N_4498,N_4302,N_4329);
xnor U4499 (N_4499,N_4261,N_4274);
xor U4500 (N_4500,N_4389,N_4289);
or U4501 (N_4501,N_4361,N_4258);
xnor U4502 (N_4502,N_4391,N_4257);
or U4503 (N_4503,N_4240,N_4344);
and U4504 (N_4504,N_4204,N_4357);
nand U4505 (N_4505,N_4275,N_4203);
xnor U4506 (N_4506,N_4393,N_4360);
or U4507 (N_4507,N_4287,N_4223);
or U4508 (N_4508,N_4306,N_4382);
xnor U4509 (N_4509,N_4257,N_4360);
or U4510 (N_4510,N_4237,N_4389);
or U4511 (N_4511,N_4304,N_4378);
or U4512 (N_4512,N_4246,N_4310);
xnor U4513 (N_4513,N_4358,N_4205);
or U4514 (N_4514,N_4392,N_4212);
nand U4515 (N_4515,N_4285,N_4263);
or U4516 (N_4516,N_4349,N_4317);
or U4517 (N_4517,N_4235,N_4359);
xnor U4518 (N_4518,N_4363,N_4212);
nand U4519 (N_4519,N_4382,N_4392);
nor U4520 (N_4520,N_4269,N_4310);
nand U4521 (N_4521,N_4393,N_4380);
nand U4522 (N_4522,N_4275,N_4332);
xnor U4523 (N_4523,N_4286,N_4249);
xor U4524 (N_4524,N_4253,N_4230);
and U4525 (N_4525,N_4336,N_4239);
or U4526 (N_4526,N_4225,N_4307);
or U4527 (N_4527,N_4213,N_4270);
xor U4528 (N_4528,N_4239,N_4386);
and U4529 (N_4529,N_4357,N_4215);
or U4530 (N_4530,N_4296,N_4212);
nand U4531 (N_4531,N_4339,N_4345);
and U4532 (N_4532,N_4231,N_4333);
xor U4533 (N_4533,N_4360,N_4396);
or U4534 (N_4534,N_4238,N_4228);
nor U4535 (N_4535,N_4250,N_4397);
nor U4536 (N_4536,N_4347,N_4370);
or U4537 (N_4537,N_4229,N_4285);
and U4538 (N_4538,N_4340,N_4329);
or U4539 (N_4539,N_4299,N_4222);
or U4540 (N_4540,N_4354,N_4272);
xor U4541 (N_4541,N_4293,N_4368);
and U4542 (N_4542,N_4241,N_4392);
or U4543 (N_4543,N_4281,N_4275);
or U4544 (N_4544,N_4359,N_4372);
xor U4545 (N_4545,N_4309,N_4273);
xnor U4546 (N_4546,N_4384,N_4228);
nor U4547 (N_4547,N_4269,N_4382);
and U4548 (N_4548,N_4296,N_4232);
or U4549 (N_4549,N_4338,N_4322);
and U4550 (N_4550,N_4243,N_4276);
nand U4551 (N_4551,N_4391,N_4251);
and U4552 (N_4552,N_4238,N_4288);
xnor U4553 (N_4553,N_4368,N_4387);
and U4554 (N_4554,N_4325,N_4321);
nor U4555 (N_4555,N_4394,N_4214);
xor U4556 (N_4556,N_4241,N_4385);
and U4557 (N_4557,N_4330,N_4288);
nor U4558 (N_4558,N_4389,N_4279);
nor U4559 (N_4559,N_4217,N_4305);
or U4560 (N_4560,N_4331,N_4204);
or U4561 (N_4561,N_4376,N_4360);
nor U4562 (N_4562,N_4210,N_4348);
xor U4563 (N_4563,N_4270,N_4245);
nor U4564 (N_4564,N_4313,N_4344);
nor U4565 (N_4565,N_4362,N_4306);
or U4566 (N_4566,N_4221,N_4247);
xnor U4567 (N_4567,N_4367,N_4214);
nand U4568 (N_4568,N_4248,N_4237);
or U4569 (N_4569,N_4223,N_4338);
nor U4570 (N_4570,N_4349,N_4321);
xor U4571 (N_4571,N_4320,N_4232);
nand U4572 (N_4572,N_4394,N_4291);
xnor U4573 (N_4573,N_4372,N_4318);
or U4574 (N_4574,N_4302,N_4278);
xor U4575 (N_4575,N_4201,N_4347);
and U4576 (N_4576,N_4377,N_4296);
xor U4577 (N_4577,N_4308,N_4307);
and U4578 (N_4578,N_4218,N_4255);
or U4579 (N_4579,N_4214,N_4388);
nand U4580 (N_4580,N_4275,N_4204);
xnor U4581 (N_4581,N_4334,N_4336);
nand U4582 (N_4582,N_4382,N_4309);
or U4583 (N_4583,N_4359,N_4293);
and U4584 (N_4584,N_4204,N_4342);
or U4585 (N_4585,N_4336,N_4313);
or U4586 (N_4586,N_4271,N_4210);
xor U4587 (N_4587,N_4216,N_4272);
nor U4588 (N_4588,N_4358,N_4302);
nor U4589 (N_4589,N_4299,N_4202);
nor U4590 (N_4590,N_4390,N_4373);
xor U4591 (N_4591,N_4327,N_4385);
nor U4592 (N_4592,N_4335,N_4283);
and U4593 (N_4593,N_4393,N_4208);
nand U4594 (N_4594,N_4223,N_4359);
xnor U4595 (N_4595,N_4237,N_4291);
and U4596 (N_4596,N_4235,N_4310);
and U4597 (N_4597,N_4355,N_4313);
nand U4598 (N_4598,N_4380,N_4210);
nor U4599 (N_4599,N_4221,N_4355);
and U4600 (N_4600,N_4439,N_4494);
and U4601 (N_4601,N_4426,N_4430);
nor U4602 (N_4602,N_4500,N_4475);
and U4603 (N_4603,N_4535,N_4401);
xnor U4604 (N_4604,N_4434,N_4577);
and U4605 (N_4605,N_4530,N_4538);
and U4606 (N_4606,N_4478,N_4550);
xnor U4607 (N_4607,N_4453,N_4521);
and U4608 (N_4608,N_4507,N_4583);
or U4609 (N_4609,N_4413,N_4579);
and U4610 (N_4610,N_4597,N_4450);
xor U4611 (N_4611,N_4465,N_4573);
and U4612 (N_4612,N_4497,N_4543);
or U4613 (N_4613,N_4506,N_4463);
or U4614 (N_4614,N_4568,N_4487);
nand U4615 (N_4615,N_4437,N_4576);
nand U4616 (N_4616,N_4524,N_4540);
nor U4617 (N_4617,N_4518,N_4536);
or U4618 (N_4618,N_4508,N_4484);
nor U4619 (N_4619,N_4408,N_4404);
nand U4620 (N_4620,N_4471,N_4525);
nand U4621 (N_4621,N_4454,N_4402);
nor U4622 (N_4622,N_4489,N_4474);
and U4623 (N_4623,N_4488,N_4537);
nand U4624 (N_4624,N_4479,N_4467);
or U4625 (N_4625,N_4468,N_4517);
and U4626 (N_4626,N_4495,N_4588);
nand U4627 (N_4627,N_4476,N_4527);
and U4628 (N_4628,N_4582,N_4458);
or U4629 (N_4629,N_4455,N_4457);
nand U4630 (N_4630,N_4572,N_4586);
or U4631 (N_4631,N_4549,N_4442);
or U4632 (N_4632,N_4592,N_4539);
or U4633 (N_4633,N_4460,N_4512);
nand U4634 (N_4634,N_4425,N_4416);
nor U4635 (N_4635,N_4485,N_4526);
nand U4636 (N_4636,N_4429,N_4503);
nand U4637 (N_4637,N_4498,N_4464);
or U4638 (N_4638,N_4510,N_4505);
xor U4639 (N_4639,N_4483,N_4433);
nor U4640 (N_4640,N_4481,N_4532);
and U4641 (N_4641,N_4421,N_4417);
nor U4642 (N_4642,N_4546,N_4492);
xor U4643 (N_4643,N_4519,N_4480);
nor U4644 (N_4644,N_4559,N_4511);
nor U4645 (N_4645,N_4422,N_4569);
nand U4646 (N_4646,N_4482,N_4574);
xnor U4647 (N_4647,N_4522,N_4462);
nor U4648 (N_4648,N_4560,N_4555);
and U4649 (N_4649,N_4558,N_4581);
xnor U4650 (N_4650,N_4553,N_4420);
and U4651 (N_4651,N_4469,N_4490);
nor U4652 (N_4652,N_4590,N_4570);
nand U4653 (N_4653,N_4473,N_4591);
xor U4654 (N_4654,N_4423,N_4578);
nand U4655 (N_4655,N_4456,N_4477);
xor U4656 (N_4656,N_4584,N_4444);
or U4657 (N_4657,N_4514,N_4501);
and U4658 (N_4658,N_4571,N_4405);
or U4659 (N_4659,N_4431,N_4438);
xnor U4660 (N_4660,N_4561,N_4446);
or U4661 (N_4661,N_4427,N_4554);
nand U4662 (N_4662,N_4424,N_4580);
or U4663 (N_4663,N_4445,N_4556);
and U4664 (N_4664,N_4496,N_4403);
and U4665 (N_4665,N_4599,N_4585);
nor U4666 (N_4666,N_4428,N_4443);
or U4667 (N_4667,N_4459,N_4513);
nor U4668 (N_4668,N_4409,N_4406);
nand U4669 (N_4669,N_4436,N_4449);
or U4670 (N_4670,N_4528,N_4440);
and U4671 (N_4671,N_4541,N_4551);
nor U4672 (N_4672,N_4415,N_4520);
nor U4673 (N_4673,N_4419,N_4400);
xnor U4674 (N_4674,N_4435,N_4563);
nor U4675 (N_4675,N_4491,N_4441);
or U4676 (N_4676,N_4547,N_4410);
nor U4677 (N_4677,N_4557,N_4411);
nand U4678 (N_4678,N_4486,N_4412);
nand U4679 (N_4679,N_4504,N_4451);
nor U4680 (N_4680,N_4593,N_4565);
nand U4681 (N_4681,N_4598,N_4515);
or U4682 (N_4682,N_4564,N_4545);
nand U4683 (N_4683,N_4562,N_4502);
nand U4684 (N_4684,N_4448,N_4596);
or U4685 (N_4685,N_4447,N_4594);
xnor U4686 (N_4686,N_4589,N_4516);
or U4687 (N_4687,N_4566,N_4533);
and U4688 (N_4688,N_4542,N_4414);
nor U4689 (N_4689,N_4461,N_4548);
and U4690 (N_4690,N_4466,N_4567);
or U4691 (N_4691,N_4509,N_4534);
xor U4692 (N_4692,N_4499,N_4552);
xor U4693 (N_4693,N_4472,N_4418);
xor U4694 (N_4694,N_4407,N_4452);
nand U4695 (N_4695,N_4432,N_4587);
nor U4696 (N_4696,N_4470,N_4595);
xor U4697 (N_4697,N_4575,N_4531);
or U4698 (N_4698,N_4523,N_4544);
xnor U4699 (N_4699,N_4493,N_4529);
xnor U4700 (N_4700,N_4565,N_4596);
xor U4701 (N_4701,N_4520,N_4451);
or U4702 (N_4702,N_4588,N_4419);
nand U4703 (N_4703,N_4555,N_4490);
or U4704 (N_4704,N_4552,N_4535);
nor U4705 (N_4705,N_4559,N_4448);
nand U4706 (N_4706,N_4471,N_4421);
nor U4707 (N_4707,N_4483,N_4519);
or U4708 (N_4708,N_4558,N_4446);
and U4709 (N_4709,N_4527,N_4409);
and U4710 (N_4710,N_4582,N_4580);
and U4711 (N_4711,N_4407,N_4403);
or U4712 (N_4712,N_4403,N_4572);
or U4713 (N_4713,N_4577,N_4502);
and U4714 (N_4714,N_4473,N_4479);
nand U4715 (N_4715,N_4469,N_4582);
and U4716 (N_4716,N_4474,N_4492);
nand U4717 (N_4717,N_4409,N_4404);
xor U4718 (N_4718,N_4405,N_4503);
xnor U4719 (N_4719,N_4516,N_4408);
nor U4720 (N_4720,N_4413,N_4493);
xnor U4721 (N_4721,N_4588,N_4579);
or U4722 (N_4722,N_4522,N_4442);
or U4723 (N_4723,N_4589,N_4503);
nor U4724 (N_4724,N_4410,N_4546);
or U4725 (N_4725,N_4595,N_4439);
and U4726 (N_4726,N_4408,N_4523);
xnor U4727 (N_4727,N_4575,N_4407);
and U4728 (N_4728,N_4557,N_4489);
and U4729 (N_4729,N_4511,N_4411);
nor U4730 (N_4730,N_4520,N_4423);
nand U4731 (N_4731,N_4578,N_4433);
xnor U4732 (N_4732,N_4520,N_4538);
nor U4733 (N_4733,N_4591,N_4532);
nand U4734 (N_4734,N_4543,N_4508);
nand U4735 (N_4735,N_4580,N_4522);
or U4736 (N_4736,N_4466,N_4564);
nor U4737 (N_4737,N_4533,N_4521);
nand U4738 (N_4738,N_4467,N_4592);
and U4739 (N_4739,N_4497,N_4579);
nor U4740 (N_4740,N_4496,N_4502);
and U4741 (N_4741,N_4530,N_4535);
nand U4742 (N_4742,N_4497,N_4429);
xor U4743 (N_4743,N_4452,N_4414);
or U4744 (N_4744,N_4452,N_4408);
and U4745 (N_4745,N_4424,N_4569);
nand U4746 (N_4746,N_4433,N_4422);
and U4747 (N_4747,N_4419,N_4553);
nand U4748 (N_4748,N_4457,N_4416);
nand U4749 (N_4749,N_4428,N_4579);
nor U4750 (N_4750,N_4408,N_4580);
nor U4751 (N_4751,N_4568,N_4585);
xnor U4752 (N_4752,N_4412,N_4443);
xor U4753 (N_4753,N_4486,N_4426);
xnor U4754 (N_4754,N_4402,N_4596);
nor U4755 (N_4755,N_4435,N_4482);
or U4756 (N_4756,N_4464,N_4471);
or U4757 (N_4757,N_4454,N_4567);
and U4758 (N_4758,N_4517,N_4441);
nor U4759 (N_4759,N_4425,N_4546);
nand U4760 (N_4760,N_4509,N_4581);
xnor U4761 (N_4761,N_4486,N_4490);
or U4762 (N_4762,N_4444,N_4554);
or U4763 (N_4763,N_4568,N_4506);
xnor U4764 (N_4764,N_4532,N_4559);
and U4765 (N_4765,N_4430,N_4522);
nor U4766 (N_4766,N_4501,N_4533);
xor U4767 (N_4767,N_4586,N_4560);
nand U4768 (N_4768,N_4590,N_4529);
nor U4769 (N_4769,N_4538,N_4498);
or U4770 (N_4770,N_4544,N_4473);
xor U4771 (N_4771,N_4400,N_4593);
nor U4772 (N_4772,N_4501,N_4510);
or U4773 (N_4773,N_4530,N_4407);
nor U4774 (N_4774,N_4516,N_4444);
nor U4775 (N_4775,N_4481,N_4453);
and U4776 (N_4776,N_4577,N_4566);
and U4777 (N_4777,N_4527,N_4450);
nor U4778 (N_4778,N_4491,N_4432);
and U4779 (N_4779,N_4527,N_4540);
and U4780 (N_4780,N_4599,N_4573);
or U4781 (N_4781,N_4455,N_4495);
and U4782 (N_4782,N_4532,N_4473);
xor U4783 (N_4783,N_4543,N_4529);
nor U4784 (N_4784,N_4473,N_4474);
or U4785 (N_4785,N_4567,N_4448);
and U4786 (N_4786,N_4461,N_4425);
nand U4787 (N_4787,N_4492,N_4472);
xor U4788 (N_4788,N_4593,N_4437);
xor U4789 (N_4789,N_4595,N_4592);
nand U4790 (N_4790,N_4555,N_4461);
or U4791 (N_4791,N_4485,N_4540);
or U4792 (N_4792,N_4464,N_4486);
nand U4793 (N_4793,N_4528,N_4424);
xnor U4794 (N_4794,N_4592,N_4536);
and U4795 (N_4795,N_4414,N_4412);
or U4796 (N_4796,N_4542,N_4401);
nand U4797 (N_4797,N_4493,N_4436);
xnor U4798 (N_4798,N_4492,N_4565);
and U4799 (N_4799,N_4446,N_4580);
and U4800 (N_4800,N_4640,N_4712);
nor U4801 (N_4801,N_4611,N_4626);
nand U4802 (N_4802,N_4665,N_4787);
and U4803 (N_4803,N_4682,N_4703);
nand U4804 (N_4804,N_4649,N_4694);
and U4805 (N_4805,N_4692,N_4687);
xor U4806 (N_4806,N_4751,N_4757);
nand U4807 (N_4807,N_4653,N_4702);
nand U4808 (N_4808,N_4658,N_4614);
nor U4809 (N_4809,N_4723,N_4796);
nor U4810 (N_4810,N_4679,N_4686);
nand U4811 (N_4811,N_4747,N_4625);
or U4812 (N_4812,N_4685,N_4616);
nor U4813 (N_4813,N_4765,N_4790);
xnor U4814 (N_4814,N_4774,N_4793);
xnor U4815 (N_4815,N_4600,N_4788);
nor U4816 (N_4816,N_4607,N_4717);
nor U4817 (N_4817,N_4627,N_4630);
and U4818 (N_4818,N_4612,N_4732);
and U4819 (N_4819,N_4775,N_4759);
or U4820 (N_4820,N_4720,N_4768);
nor U4821 (N_4821,N_4719,N_4786);
or U4822 (N_4822,N_4780,N_4680);
nor U4823 (N_4823,N_4794,N_4606);
nand U4824 (N_4824,N_4672,N_4746);
xnor U4825 (N_4825,N_4709,N_4740);
nor U4826 (N_4826,N_4727,N_4769);
or U4827 (N_4827,N_4766,N_4622);
or U4828 (N_4828,N_4615,N_4754);
or U4829 (N_4829,N_4652,N_4648);
nor U4830 (N_4830,N_4738,N_4799);
nand U4831 (N_4831,N_4684,N_4735);
and U4832 (N_4832,N_4700,N_4722);
and U4833 (N_4833,N_4795,N_4742);
or U4834 (N_4834,N_4748,N_4761);
xnor U4835 (N_4835,N_4601,N_4724);
nand U4836 (N_4836,N_4666,N_4676);
nand U4837 (N_4837,N_4731,N_4755);
xnor U4838 (N_4838,N_4789,N_4613);
and U4839 (N_4839,N_4655,N_4671);
or U4840 (N_4840,N_4714,N_4739);
xnor U4841 (N_4841,N_4681,N_4741);
nor U4842 (N_4842,N_4637,N_4762);
and U4843 (N_4843,N_4688,N_4704);
and U4844 (N_4844,N_4728,N_4764);
nor U4845 (N_4845,N_4781,N_4629);
or U4846 (N_4846,N_4609,N_4784);
nand U4847 (N_4847,N_4628,N_4651);
nand U4848 (N_4848,N_4638,N_4621);
nand U4849 (N_4849,N_4699,N_4707);
xnor U4850 (N_4850,N_4696,N_4641);
nor U4851 (N_4851,N_4698,N_4752);
and U4852 (N_4852,N_4791,N_4604);
nor U4853 (N_4853,N_4753,N_4773);
xnor U4854 (N_4854,N_4770,N_4744);
nand U4855 (N_4855,N_4726,N_4677);
nand U4856 (N_4856,N_4729,N_4792);
xnor U4857 (N_4857,N_4619,N_4695);
nand U4858 (N_4858,N_4708,N_4711);
nor U4859 (N_4859,N_4624,N_4618);
nand U4860 (N_4860,N_4661,N_4697);
nand U4861 (N_4861,N_4716,N_4660);
and U4862 (N_4862,N_4771,N_4636);
nand U4863 (N_4863,N_4733,N_4634);
nor U4864 (N_4864,N_4645,N_4602);
nor U4865 (N_4865,N_4633,N_4635);
nand U4866 (N_4866,N_4617,N_4691);
nor U4867 (N_4867,N_4737,N_4797);
xnor U4868 (N_4868,N_4693,N_4767);
and U4869 (N_4869,N_4678,N_4776);
or U4870 (N_4870,N_4643,N_4659);
xnor U4871 (N_4871,N_4644,N_4646);
nor U4872 (N_4872,N_4639,N_4721);
xor U4873 (N_4873,N_4749,N_4750);
nor U4874 (N_4874,N_4760,N_4725);
and U4875 (N_4875,N_4690,N_4608);
or U4876 (N_4876,N_4675,N_4674);
nor U4877 (N_4877,N_4756,N_4654);
nand U4878 (N_4878,N_4663,N_4736);
and U4879 (N_4879,N_4785,N_4668);
and U4880 (N_4880,N_4689,N_4667);
nor U4881 (N_4881,N_4772,N_4798);
xor U4882 (N_4882,N_4713,N_4763);
xnor U4883 (N_4883,N_4743,N_4705);
xor U4884 (N_4884,N_4782,N_4718);
and U4885 (N_4885,N_4631,N_4664);
nand U4886 (N_4886,N_4662,N_4650);
or U4887 (N_4887,N_4603,N_4783);
nand U4888 (N_4888,N_4777,N_4673);
nand U4889 (N_4889,N_4758,N_4620);
or U4890 (N_4890,N_4605,N_4706);
or U4891 (N_4891,N_4730,N_4683);
nor U4892 (N_4892,N_4701,N_4623);
and U4893 (N_4893,N_4610,N_4734);
and U4894 (N_4894,N_4778,N_4656);
or U4895 (N_4895,N_4779,N_4647);
nand U4896 (N_4896,N_4642,N_4632);
nor U4897 (N_4897,N_4715,N_4657);
and U4898 (N_4898,N_4670,N_4745);
nand U4899 (N_4899,N_4710,N_4669);
and U4900 (N_4900,N_4741,N_4725);
and U4901 (N_4901,N_4653,N_4727);
or U4902 (N_4902,N_4653,N_4682);
xor U4903 (N_4903,N_4673,N_4739);
or U4904 (N_4904,N_4773,N_4776);
nor U4905 (N_4905,N_4623,N_4783);
nor U4906 (N_4906,N_4638,N_4644);
nand U4907 (N_4907,N_4737,N_4631);
and U4908 (N_4908,N_4612,N_4638);
and U4909 (N_4909,N_4783,N_4712);
or U4910 (N_4910,N_4765,N_4784);
nor U4911 (N_4911,N_4778,N_4693);
or U4912 (N_4912,N_4745,N_4722);
and U4913 (N_4913,N_4703,N_4749);
nor U4914 (N_4914,N_4672,N_4753);
xor U4915 (N_4915,N_4798,N_4776);
or U4916 (N_4916,N_4644,N_4726);
and U4917 (N_4917,N_4636,N_4764);
nor U4918 (N_4918,N_4652,N_4688);
and U4919 (N_4919,N_4703,N_4774);
nor U4920 (N_4920,N_4616,N_4744);
nor U4921 (N_4921,N_4602,N_4756);
and U4922 (N_4922,N_4686,N_4617);
xnor U4923 (N_4923,N_4725,N_4794);
nand U4924 (N_4924,N_4735,N_4719);
nand U4925 (N_4925,N_4607,N_4764);
xor U4926 (N_4926,N_4779,N_4795);
nor U4927 (N_4927,N_4660,N_4754);
or U4928 (N_4928,N_4699,N_4711);
and U4929 (N_4929,N_4659,N_4611);
xnor U4930 (N_4930,N_4711,N_4609);
or U4931 (N_4931,N_4700,N_4662);
nor U4932 (N_4932,N_4612,N_4626);
or U4933 (N_4933,N_4657,N_4698);
nand U4934 (N_4934,N_4723,N_4609);
or U4935 (N_4935,N_4622,N_4719);
or U4936 (N_4936,N_4657,N_4758);
xor U4937 (N_4937,N_4716,N_4720);
nand U4938 (N_4938,N_4724,N_4699);
nand U4939 (N_4939,N_4701,N_4683);
nand U4940 (N_4940,N_4796,N_4776);
and U4941 (N_4941,N_4635,N_4631);
and U4942 (N_4942,N_4695,N_4737);
xor U4943 (N_4943,N_4744,N_4720);
nor U4944 (N_4944,N_4737,N_4731);
and U4945 (N_4945,N_4766,N_4657);
nand U4946 (N_4946,N_4744,N_4661);
nand U4947 (N_4947,N_4694,N_4617);
nor U4948 (N_4948,N_4718,N_4770);
nor U4949 (N_4949,N_4766,N_4756);
nor U4950 (N_4950,N_4748,N_4713);
and U4951 (N_4951,N_4682,N_4734);
nand U4952 (N_4952,N_4727,N_4695);
nand U4953 (N_4953,N_4771,N_4629);
nand U4954 (N_4954,N_4659,N_4713);
xnor U4955 (N_4955,N_4634,N_4638);
xnor U4956 (N_4956,N_4793,N_4639);
and U4957 (N_4957,N_4655,N_4637);
nand U4958 (N_4958,N_4666,N_4670);
xor U4959 (N_4959,N_4784,N_4697);
nand U4960 (N_4960,N_4674,N_4670);
xnor U4961 (N_4961,N_4741,N_4654);
or U4962 (N_4962,N_4694,N_4651);
and U4963 (N_4963,N_4746,N_4753);
and U4964 (N_4964,N_4776,N_4688);
or U4965 (N_4965,N_4738,N_4725);
and U4966 (N_4966,N_4795,N_4653);
or U4967 (N_4967,N_4612,N_4796);
xnor U4968 (N_4968,N_4663,N_4638);
nand U4969 (N_4969,N_4687,N_4646);
nor U4970 (N_4970,N_4661,N_4775);
xnor U4971 (N_4971,N_4677,N_4631);
and U4972 (N_4972,N_4634,N_4796);
or U4973 (N_4973,N_4699,N_4690);
nor U4974 (N_4974,N_4653,N_4715);
and U4975 (N_4975,N_4741,N_4627);
xnor U4976 (N_4976,N_4740,N_4639);
or U4977 (N_4977,N_4662,N_4644);
or U4978 (N_4978,N_4761,N_4711);
or U4979 (N_4979,N_4681,N_4705);
nand U4980 (N_4980,N_4679,N_4602);
and U4981 (N_4981,N_4650,N_4671);
nor U4982 (N_4982,N_4630,N_4644);
nand U4983 (N_4983,N_4779,N_4685);
and U4984 (N_4984,N_4707,N_4695);
nand U4985 (N_4985,N_4666,N_4689);
nor U4986 (N_4986,N_4641,N_4747);
nor U4987 (N_4987,N_4774,N_4734);
and U4988 (N_4988,N_4664,N_4692);
nand U4989 (N_4989,N_4687,N_4688);
nand U4990 (N_4990,N_4759,N_4720);
and U4991 (N_4991,N_4772,N_4698);
xnor U4992 (N_4992,N_4713,N_4795);
nor U4993 (N_4993,N_4721,N_4619);
and U4994 (N_4994,N_4652,N_4642);
nand U4995 (N_4995,N_4660,N_4635);
xnor U4996 (N_4996,N_4749,N_4723);
and U4997 (N_4997,N_4790,N_4762);
and U4998 (N_4998,N_4637,N_4788);
nor U4999 (N_4999,N_4602,N_4662);
nor U5000 (N_5000,N_4937,N_4977);
xor U5001 (N_5001,N_4845,N_4946);
and U5002 (N_5002,N_4813,N_4951);
or U5003 (N_5003,N_4941,N_4907);
and U5004 (N_5004,N_4928,N_4875);
nor U5005 (N_5005,N_4893,N_4870);
xnor U5006 (N_5006,N_4913,N_4874);
nand U5007 (N_5007,N_4862,N_4891);
nand U5008 (N_5008,N_4814,N_4973);
nand U5009 (N_5009,N_4965,N_4803);
and U5010 (N_5010,N_4938,N_4948);
nand U5011 (N_5011,N_4877,N_4890);
and U5012 (N_5012,N_4805,N_4866);
or U5013 (N_5013,N_4978,N_4936);
xnor U5014 (N_5014,N_4921,N_4927);
nor U5015 (N_5015,N_4999,N_4915);
nor U5016 (N_5016,N_4811,N_4909);
and U5017 (N_5017,N_4993,N_4884);
or U5018 (N_5018,N_4919,N_4895);
xor U5019 (N_5019,N_4887,N_4869);
xor U5020 (N_5020,N_4853,N_4989);
and U5021 (N_5021,N_4901,N_4836);
or U5022 (N_5022,N_4850,N_4934);
nor U5023 (N_5023,N_4984,N_4806);
nor U5024 (N_5024,N_4894,N_4922);
xor U5025 (N_5025,N_4988,N_4958);
nor U5026 (N_5026,N_4840,N_4912);
or U5027 (N_5027,N_4865,N_4910);
nand U5028 (N_5028,N_4835,N_4963);
xnor U5029 (N_5029,N_4985,N_4995);
nor U5030 (N_5030,N_4983,N_4878);
nor U5031 (N_5031,N_4829,N_4810);
xnor U5032 (N_5032,N_4838,N_4943);
and U5033 (N_5033,N_4967,N_4974);
and U5034 (N_5034,N_4992,N_4807);
xnor U5035 (N_5035,N_4867,N_4952);
nand U5036 (N_5036,N_4809,N_4815);
nand U5037 (N_5037,N_4854,N_4953);
or U5038 (N_5038,N_4879,N_4966);
or U5039 (N_5039,N_4855,N_4883);
and U5040 (N_5040,N_4896,N_4846);
nor U5041 (N_5041,N_4825,N_4826);
or U5042 (N_5042,N_4960,N_4833);
nand U5043 (N_5043,N_4902,N_4804);
nor U5044 (N_5044,N_4998,N_4931);
and U5045 (N_5045,N_4820,N_4823);
xor U5046 (N_5046,N_4980,N_4860);
nor U5047 (N_5047,N_4947,N_4961);
xnor U5048 (N_5048,N_4920,N_4970);
nor U5049 (N_5049,N_4843,N_4849);
or U5050 (N_5050,N_4924,N_4905);
and U5051 (N_5051,N_4876,N_4824);
or U5052 (N_5052,N_4904,N_4819);
or U5053 (N_5053,N_4935,N_4839);
nand U5054 (N_5054,N_4817,N_4885);
xnor U5055 (N_5055,N_4997,N_4914);
xnor U5056 (N_5056,N_4945,N_4994);
or U5057 (N_5057,N_4949,N_4917);
and U5058 (N_5058,N_4933,N_4889);
and U5059 (N_5059,N_4834,N_4976);
nor U5060 (N_5060,N_4990,N_4898);
and U5061 (N_5061,N_4930,N_4880);
and U5062 (N_5062,N_4903,N_4954);
or U5063 (N_5063,N_4848,N_4856);
or U5064 (N_5064,N_4816,N_4842);
nor U5065 (N_5065,N_4906,N_4858);
or U5066 (N_5066,N_4957,N_4832);
nor U5067 (N_5067,N_4929,N_4861);
nand U5068 (N_5068,N_4981,N_4911);
or U5069 (N_5069,N_4808,N_4802);
nor U5070 (N_5070,N_4852,N_4962);
or U5071 (N_5071,N_4864,N_4987);
xor U5072 (N_5072,N_4932,N_4872);
or U5073 (N_5073,N_4897,N_4801);
or U5074 (N_5074,N_4975,N_4956);
or U5075 (N_5075,N_4955,N_4863);
nand U5076 (N_5076,N_4828,N_4982);
or U5077 (N_5077,N_4821,N_4991);
nor U5078 (N_5078,N_4837,N_4900);
nand U5079 (N_5079,N_4908,N_4859);
or U5080 (N_5080,N_4899,N_4857);
and U5081 (N_5081,N_4841,N_4959);
and U5082 (N_5082,N_4830,N_4886);
xnor U5083 (N_5083,N_4916,N_4827);
and U5084 (N_5084,N_4972,N_4888);
xnor U5085 (N_5085,N_4873,N_4996);
nand U5086 (N_5086,N_4882,N_4868);
xor U5087 (N_5087,N_4847,N_4881);
nor U5088 (N_5088,N_4926,N_4942);
or U5089 (N_5089,N_4971,N_4918);
or U5090 (N_5090,N_4818,N_4964);
and U5091 (N_5091,N_4950,N_4800);
xor U5092 (N_5092,N_4925,N_4812);
nor U5093 (N_5093,N_4940,N_4851);
nor U5094 (N_5094,N_4844,N_4968);
xnor U5095 (N_5095,N_4969,N_4979);
xnor U5096 (N_5096,N_4944,N_4892);
xnor U5097 (N_5097,N_4939,N_4986);
and U5098 (N_5098,N_4822,N_4871);
nor U5099 (N_5099,N_4923,N_4831);
nand U5100 (N_5100,N_4858,N_4859);
or U5101 (N_5101,N_4935,N_4834);
nand U5102 (N_5102,N_4873,N_4833);
nand U5103 (N_5103,N_4921,N_4973);
or U5104 (N_5104,N_4968,N_4965);
xnor U5105 (N_5105,N_4974,N_4855);
or U5106 (N_5106,N_4940,N_4902);
xor U5107 (N_5107,N_4941,N_4853);
nor U5108 (N_5108,N_4928,N_4946);
nor U5109 (N_5109,N_4881,N_4851);
and U5110 (N_5110,N_4958,N_4878);
nand U5111 (N_5111,N_4872,N_4824);
nor U5112 (N_5112,N_4922,N_4837);
nor U5113 (N_5113,N_4904,N_4882);
xnor U5114 (N_5114,N_4957,N_4996);
or U5115 (N_5115,N_4817,N_4955);
nand U5116 (N_5116,N_4941,N_4844);
nand U5117 (N_5117,N_4971,N_4944);
and U5118 (N_5118,N_4991,N_4852);
or U5119 (N_5119,N_4825,N_4995);
xor U5120 (N_5120,N_4900,N_4814);
nor U5121 (N_5121,N_4983,N_4888);
nand U5122 (N_5122,N_4865,N_4827);
nor U5123 (N_5123,N_4873,N_4945);
nor U5124 (N_5124,N_4839,N_4931);
nand U5125 (N_5125,N_4911,N_4973);
or U5126 (N_5126,N_4979,N_4843);
or U5127 (N_5127,N_4808,N_4934);
and U5128 (N_5128,N_4951,N_4935);
and U5129 (N_5129,N_4906,N_4986);
or U5130 (N_5130,N_4902,N_4860);
xor U5131 (N_5131,N_4824,N_4855);
or U5132 (N_5132,N_4867,N_4983);
nor U5133 (N_5133,N_4856,N_4892);
and U5134 (N_5134,N_4831,N_4806);
xor U5135 (N_5135,N_4965,N_4826);
and U5136 (N_5136,N_4833,N_4970);
nor U5137 (N_5137,N_4961,N_4893);
and U5138 (N_5138,N_4981,N_4929);
nand U5139 (N_5139,N_4820,N_4926);
or U5140 (N_5140,N_4978,N_4803);
and U5141 (N_5141,N_4897,N_4875);
nor U5142 (N_5142,N_4993,N_4943);
xnor U5143 (N_5143,N_4933,N_4803);
or U5144 (N_5144,N_4971,N_4896);
and U5145 (N_5145,N_4880,N_4886);
or U5146 (N_5146,N_4944,N_4848);
xor U5147 (N_5147,N_4928,N_4811);
nand U5148 (N_5148,N_4864,N_4890);
xor U5149 (N_5149,N_4998,N_4905);
xor U5150 (N_5150,N_4815,N_4936);
nand U5151 (N_5151,N_4962,N_4823);
and U5152 (N_5152,N_4920,N_4843);
or U5153 (N_5153,N_4998,N_4972);
nand U5154 (N_5154,N_4930,N_4867);
xnor U5155 (N_5155,N_4996,N_4822);
and U5156 (N_5156,N_4862,N_4818);
and U5157 (N_5157,N_4950,N_4972);
nor U5158 (N_5158,N_4954,N_4906);
or U5159 (N_5159,N_4883,N_4935);
and U5160 (N_5160,N_4853,N_4953);
nand U5161 (N_5161,N_4969,N_4940);
nor U5162 (N_5162,N_4951,N_4962);
and U5163 (N_5163,N_4912,N_4898);
and U5164 (N_5164,N_4913,N_4892);
nand U5165 (N_5165,N_4894,N_4920);
and U5166 (N_5166,N_4883,N_4957);
and U5167 (N_5167,N_4827,N_4973);
nand U5168 (N_5168,N_4990,N_4889);
and U5169 (N_5169,N_4829,N_4927);
xor U5170 (N_5170,N_4987,N_4940);
nor U5171 (N_5171,N_4974,N_4963);
xor U5172 (N_5172,N_4903,N_4969);
nand U5173 (N_5173,N_4815,N_4855);
nor U5174 (N_5174,N_4878,N_4835);
nand U5175 (N_5175,N_4932,N_4866);
xor U5176 (N_5176,N_4855,N_4825);
xor U5177 (N_5177,N_4897,N_4989);
or U5178 (N_5178,N_4856,N_4919);
xnor U5179 (N_5179,N_4892,N_4979);
or U5180 (N_5180,N_4894,N_4811);
xnor U5181 (N_5181,N_4948,N_4889);
nand U5182 (N_5182,N_4951,N_4852);
nand U5183 (N_5183,N_4888,N_4829);
xor U5184 (N_5184,N_4863,N_4928);
nor U5185 (N_5185,N_4876,N_4920);
xnor U5186 (N_5186,N_4956,N_4969);
xnor U5187 (N_5187,N_4859,N_4836);
nand U5188 (N_5188,N_4910,N_4999);
nor U5189 (N_5189,N_4857,N_4951);
nor U5190 (N_5190,N_4878,N_4991);
nand U5191 (N_5191,N_4934,N_4999);
and U5192 (N_5192,N_4870,N_4887);
nor U5193 (N_5193,N_4840,N_4867);
or U5194 (N_5194,N_4823,N_4959);
or U5195 (N_5195,N_4891,N_4910);
or U5196 (N_5196,N_4809,N_4902);
nor U5197 (N_5197,N_4902,N_4963);
nand U5198 (N_5198,N_4813,N_4843);
nor U5199 (N_5199,N_4964,N_4883);
or U5200 (N_5200,N_5095,N_5111);
or U5201 (N_5201,N_5021,N_5077);
nor U5202 (N_5202,N_5121,N_5166);
xnor U5203 (N_5203,N_5048,N_5199);
and U5204 (N_5204,N_5162,N_5159);
and U5205 (N_5205,N_5170,N_5198);
nor U5206 (N_5206,N_5144,N_5184);
or U5207 (N_5207,N_5059,N_5006);
nand U5208 (N_5208,N_5026,N_5116);
nor U5209 (N_5209,N_5132,N_5093);
nor U5210 (N_5210,N_5073,N_5051);
and U5211 (N_5211,N_5112,N_5164);
nor U5212 (N_5212,N_5137,N_5108);
nor U5213 (N_5213,N_5169,N_5083);
xnor U5214 (N_5214,N_5102,N_5045);
and U5215 (N_5215,N_5018,N_5038);
xor U5216 (N_5216,N_5053,N_5066);
xor U5217 (N_5217,N_5123,N_5193);
or U5218 (N_5218,N_5019,N_5014);
or U5219 (N_5219,N_5007,N_5020);
xor U5220 (N_5220,N_5015,N_5029);
and U5221 (N_5221,N_5003,N_5180);
nand U5222 (N_5222,N_5060,N_5145);
nand U5223 (N_5223,N_5150,N_5172);
xor U5224 (N_5224,N_5008,N_5074);
or U5225 (N_5225,N_5085,N_5161);
and U5226 (N_5226,N_5005,N_5041);
nor U5227 (N_5227,N_5151,N_5188);
nand U5228 (N_5228,N_5027,N_5192);
and U5229 (N_5229,N_5183,N_5174);
xor U5230 (N_5230,N_5129,N_5195);
xor U5231 (N_5231,N_5030,N_5067);
nand U5232 (N_5232,N_5156,N_5043);
nor U5233 (N_5233,N_5147,N_5042);
nor U5234 (N_5234,N_5013,N_5082);
nor U5235 (N_5235,N_5122,N_5040);
or U5236 (N_5236,N_5194,N_5099);
xnor U5237 (N_5237,N_5039,N_5153);
nand U5238 (N_5238,N_5107,N_5154);
nor U5239 (N_5239,N_5177,N_5143);
nand U5240 (N_5240,N_5023,N_5110);
nor U5241 (N_5241,N_5181,N_5146);
and U5242 (N_5242,N_5109,N_5179);
or U5243 (N_5243,N_5076,N_5098);
nand U5244 (N_5244,N_5057,N_5061);
and U5245 (N_5245,N_5196,N_5084);
nor U5246 (N_5246,N_5037,N_5068);
nand U5247 (N_5247,N_5106,N_5028);
and U5248 (N_5248,N_5126,N_5001);
xnor U5249 (N_5249,N_5092,N_5148);
nand U5250 (N_5250,N_5075,N_5050);
xor U5251 (N_5251,N_5114,N_5002);
or U5252 (N_5252,N_5187,N_5033);
nand U5253 (N_5253,N_5190,N_5065);
and U5254 (N_5254,N_5064,N_5191);
or U5255 (N_5255,N_5063,N_5115);
nand U5256 (N_5256,N_5127,N_5117);
and U5257 (N_5257,N_5124,N_5088);
xor U5258 (N_5258,N_5168,N_5120);
or U5259 (N_5259,N_5022,N_5157);
and U5260 (N_5260,N_5103,N_5100);
nor U5261 (N_5261,N_5087,N_5097);
xnor U5262 (N_5262,N_5130,N_5175);
nand U5263 (N_5263,N_5017,N_5049);
nand U5264 (N_5264,N_5135,N_5046);
nor U5265 (N_5265,N_5054,N_5081);
or U5266 (N_5266,N_5176,N_5080);
nor U5267 (N_5267,N_5131,N_5032);
nor U5268 (N_5268,N_5056,N_5197);
and U5269 (N_5269,N_5133,N_5178);
nor U5270 (N_5270,N_5171,N_5165);
or U5271 (N_5271,N_5118,N_5185);
nand U5272 (N_5272,N_5163,N_5072);
and U5273 (N_5273,N_5024,N_5071);
nor U5274 (N_5274,N_5094,N_5104);
or U5275 (N_5275,N_5136,N_5119);
and U5276 (N_5276,N_5089,N_5078);
and U5277 (N_5277,N_5016,N_5044);
nor U5278 (N_5278,N_5009,N_5055);
xor U5279 (N_5279,N_5025,N_5160);
nor U5280 (N_5280,N_5000,N_5105);
or U5281 (N_5281,N_5096,N_5158);
xor U5282 (N_5282,N_5142,N_5189);
nand U5283 (N_5283,N_5062,N_5034);
nand U5284 (N_5284,N_5004,N_5173);
and U5285 (N_5285,N_5069,N_5152);
nor U5286 (N_5286,N_5134,N_5011);
nand U5287 (N_5287,N_5149,N_5012);
nand U5288 (N_5288,N_5035,N_5036);
nand U5289 (N_5289,N_5113,N_5182);
or U5290 (N_5290,N_5128,N_5058);
xor U5291 (N_5291,N_5079,N_5141);
and U5292 (N_5292,N_5010,N_5125);
xor U5293 (N_5293,N_5047,N_5139);
or U5294 (N_5294,N_5091,N_5138);
nor U5295 (N_5295,N_5140,N_5155);
and U5296 (N_5296,N_5167,N_5052);
nor U5297 (N_5297,N_5031,N_5086);
nor U5298 (N_5298,N_5101,N_5090);
nand U5299 (N_5299,N_5070,N_5186);
nor U5300 (N_5300,N_5175,N_5120);
nand U5301 (N_5301,N_5145,N_5190);
nand U5302 (N_5302,N_5095,N_5109);
nor U5303 (N_5303,N_5113,N_5088);
or U5304 (N_5304,N_5151,N_5134);
nor U5305 (N_5305,N_5161,N_5113);
or U5306 (N_5306,N_5088,N_5021);
or U5307 (N_5307,N_5055,N_5185);
and U5308 (N_5308,N_5118,N_5053);
nand U5309 (N_5309,N_5146,N_5145);
xnor U5310 (N_5310,N_5028,N_5131);
or U5311 (N_5311,N_5123,N_5166);
or U5312 (N_5312,N_5140,N_5146);
nor U5313 (N_5313,N_5110,N_5009);
or U5314 (N_5314,N_5067,N_5160);
and U5315 (N_5315,N_5193,N_5132);
or U5316 (N_5316,N_5031,N_5004);
or U5317 (N_5317,N_5048,N_5017);
and U5318 (N_5318,N_5166,N_5010);
nand U5319 (N_5319,N_5041,N_5010);
nand U5320 (N_5320,N_5146,N_5001);
or U5321 (N_5321,N_5027,N_5121);
xor U5322 (N_5322,N_5108,N_5023);
and U5323 (N_5323,N_5057,N_5078);
xnor U5324 (N_5324,N_5112,N_5090);
xor U5325 (N_5325,N_5148,N_5020);
nor U5326 (N_5326,N_5026,N_5076);
or U5327 (N_5327,N_5023,N_5187);
and U5328 (N_5328,N_5151,N_5020);
nand U5329 (N_5329,N_5126,N_5105);
and U5330 (N_5330,N_5130,N_5030);
xor U5331 (N_5331,N_5052,N_5049);
or U5332 (N_5332,N_5123,N_5001);
and U5333 (N_5333,N_5036,N_5048);
and U5334 (N_5334,N_5031,N_5118);
or U5335 (N_5335,N_5039,N_5182);
nand U5336 (N_5336,N_5134,N_5159);
and U5337 (N_5337,N_5103,N_5019);
xor U5338 (N_5338,N_5138,N_5136);
nand U5339 (N_5339,N_5053,N_5135);
and U5340 (N_5340,N_5007,N_5055);
or U5341 (N_5341,N_5047,N_5109);
or U5342 (N_5342,N_5000,N_5056);
nand U5343 (N_5343,N_5067,N_5069);
xnor U5344 (N_5344,N_5127,N_5195);
or U5345 (N_5345,N_5173,N_5045);
nand U5346 (N_5346,N_5059,N_5169);
and U5347 (N_5347,N_5105,N_5199);
nand U5348 (N_5348,N_5097,N_5134);
xnor U5349 (N_5349,N_5173,N_5090);
nand U5350 (N_5350,N_5139,N_5143);
or U5351 (N_5351,N_5158,N_5084);
nor U5352 (N_5352,N_5108,N_5084);
nand U5353 (N_5353,N_5119,N_5154);
and U5354 (N_5354,N_5189,N_5072);
or U5355 (N_5355,N_5094,N_5149);
nand U5356 (N_5356,N_5171,N_5011);
xnor U5357 (N_5357,N_5012,N_5168);
xnor U5358 (N_5358,N_5128,N_5143);
nor U5359 (N_5359,N_5009,N_5019);
xnor U5360 (N_5360,N_5075,N_5045);
nand U5361 (N_5361,N_5132,N_5023);
or U5362 (N_5362,N_5022,N_5015);
nand U5363 (N_5363,N_5022,N_5094);
nor U5364 (N_5364,N_5043,N_5101);
nand U5365 (N_5365,N_5045,N_5199);
nor U5366 (N_5366,N_5166,N_5170);
xor U5367 (N_5367,N_5006,N_5184);
and U5368 (N_5368,N_5022,N_5147);
and U5369 (N_5369,N_5091,N_5108);
and U5370 (N_5370,N_5056,N_5116);
nor U5371 (N_5371,N_5094,N_5003);
and U5372 (N_5372,N_5043,N_5044);
or U5373 (N_5373,N_5058,N_5032);
nor U5374 (N_5374,N_5049,N_5072);
nor U5375 (N_5375,N_5073,N_5044);
xor U5376 (N_5376,N_5147,N_5134);
and U5377 (N_5377,N_5181,N_5177);
nor U5378 (N_5378,N_5152,N_5059);
xor U5379 (N_5379,N_5031,N_5197);
nor U5380 (N_5380,N_5009,N_5075);
nor U5381 (N_5381,N_5137,N_5000);
nor U5382 (N_5382,N_5023,N_5155);
nor U5383 (N_5383,N_5003,N_5129);
nand U5384 (N_5384,N_5016,N_5108);
nor U5385 (N_5385,N_5031,N_5063);
xor U5386 (N_5386,N_5079,N_5021);
xor U5387 (N_5387,N_5087,N_5022);
nand U5388 (N_5388,N_5156,N_5034);
or U5389 (N_5389,N_5001,N_5114);
or U5390 (N_5390,N_5145,N_5084);
or U5391 (N_5391,N_5140,N_5171);
nor U5392 (N_5392,N_5136,N_5078);
or U5393 (N_5393,N_5072,N_5123);
xnor U5394 (N_5394,N_5083,N_5186);
nand U5395 (N_5395,N_5067,N_5032);
nand U5396 (N_5396,N_5080,N_5148);
nor U5397 (N_5397,N_5090,N_5147);
nor U5398 (N_5398,N_5081,N_5102);
nor U5399 (N_5399,N_5153,N_5023);
and U5400 (N_5400,N_5368,N_5270);
and U5401 (N_5401,N_5321,N_5376);
nor U5402 (N_5402,N_5309,N_5361);
xnor U5403 (N_5403,N_5254,N_5238);
xnor U5404 (N_5404,N_5393,N_5297);
xor U5405 (N_5405,N_5200,N_5296);
nor U5406 (N_5406,N_5358,N_5252);
or U5407 (N_5407,N_5338,N_5324);
or U5408 (N_5408,N_5330,N_5326);
or U5409 (N_5409,N_5295,N_5280);
nand U5410 (N_5410,N_5255,N_5273);
nor U5411 (N_5411,N_5319,N_5300);
nor U5412 (N_5412,N_5274,N_5352);
xor U5413 (N_5413,N_5222,N_5364);
nor U5414 (N_5414,N_5267,N_5307);
and U5415 (N_5415,N_5245,N_5219);
nand U5416 (N_5416,N_5281,N_5259);
xnor U5417 (N_5417,N_5221,N_5350);
and U5418 (N_5418,N_5369,N_5397);
xnor U5419 (N_5419,N_5201,N_5204);
or U5420 (N_5420,N_5236,N_5210);
nor U5421 (N_5421,N_5353,N_5382);
and U5422 (N_5422,N_5249,N_5277);
xnor U5423 (N_5423,N_5378,N_5392);
nand U5424 (N_5424,N_5253,N_5206);
nor U5425 (N_5425,N_5208,N_5278);
xor U5426 (N_5426,N_5298,N_5264);
nand U5427 (N_5427,N_5287,N_5332);
nand U5428 (N_5428,N_5228,N_5211);
and U5429 (N_5429,N_5233,N_5363);
nor U5430 (N_5430,N_5290,N_5325);
nand U5431 (N_5431,N_5312,N_5272);
or U5432 (N_5432,N_5284,N_5289);
xnor U5433 (N_5433,N_5379,N_5327);
or U5434 (N_5434,N_5237,N_5310);
and U5435 (N_5435,N_5377,N_5302);
xor U5436 (N_5436,N_5346,N_5334);
or U5437 (N_5437,N_5225,N_5331);
or U5438 (N_5438,N_5231,N_5303);
nor U5439 (N_5439,N_5365,N_5387);
nor U5440 (N_5440,N_5360,N_5380);
nand U5441 (N_5441,N_5359,N_5243);
nor U5442 (N_5442,N_5398,N_5372);
nand U5443 (N_5443,N_5304,N_5251);
nor U5444 (N_5444,N_5329,N_5285);
and U5445 (N_5445,N_5286,N_5386);
nand U5446 (N_5446,N_5256,N_5224);
xnor U5447 (N_5447,N_5247,N_5223);
or U5448 (N_5448,N_5218,N_5362);
xnor U5449 (N_5449,N_5394,N_5235);
or U5450 (N_5450,N_5299,N_5374);
nor U5451 (N_5451,N_5239,N_5214);
xnor U5452 (N_5452,N_5265,N_5213);
nor U5453 (N_5453,N_5328,N_5306);
or U5454 (N_5454,N_5244,N_5269);
nor U5455 (N_5455,N_5395,N_5318);
nor U5456 (N_5456,N_5205,N_5260);
xor U5457 (N_5457,N_5279,N_5391);
or U5458 (N_5458,N_5314,N_5234);
nand U5459 (N_5459,N_5248,N_5226);
xnor U5460 (N_5460,N_5373,N_5323);
or U5461 (N_5461,N_5337,N_5282);
xor U5462 (N_5462,N_5355,N_5203);
xor U5463 (N_5463,N_5367,N_5202);
or U5464 (N_5464,N_5262,N_5341);
xnor U5465 (N_5465,N_5311,N_5242);
xor U5466 (N_5466,N_5292,N_5351);
and U5467 (N_5467,N_5320,N_5313);
or U5468 (N_5468,N_5383,N_5283);
or U5469 (N_5469,N_5370,N_5301);
xnor U5470 (N_5470,N_5305,N_5246);
nor U5471 (N_5471,N_5366,N_5275);
nand U5472 (N_5472,N_5227,N_5371);
nand U5473 (N_5473,N_5343,N_5385);
nand U5474 (N_5474,N_5317,N_5339);
xnor U5475 (N_5475,N_5216,N_5389);
xor U5476 (N_5476,N_5240,N_5229);
nor U5477 (N_5477,N_5207,N_5258);
and U5478 (N_5478,N_5336,N_5356);
nor U5479 (N_5479,N_5388,N_5347);
xor U5480 (N_5480,N_5340,N_5220);
xor U5481 (N_5481,N_5348,N_5230);
xor U5482 (N_5482,N_5375,N_5315);
nor U5483 (N_5483,N_5354,N_5316);
nand U5484 (N_5484,N_5266,N_5345);
or U5485 (N_5485,N_5335,N_5268);
and U5486 (N_5486,N_5232,N_5344);
nand U5487 (N_5487,N_5294,N_5276);
nand U5488 (N_5488,N_5384,N_5257);
or U5489 (N_5489,N_5250,N_5357);
and U5490 (N_5490,N_5349,N_5322);
nor U5491 (N_5491,N_5293,N_5399);
and U5492 (N_5492,N_5308,N_5390);
nand U5493 (N_5493,N_5263,N_5291);
or U5494 (N_5494,N_5241,N_5381);
or U5495 (N_5495,N_5396,N_5215);
or U5496 (N_5496,N_5271,N_5261);
nand U5497 (N_5497,N_5288,N_5342);
nor U5498 (N_5498,N_5217,N_5209);
nand U5499 (N_5499,N_5333,N_5212);
nor U5500 (N_5500,N_5216,N_5255);
or U5501 (N_5501,N_5348,N_5364);
nand U5502 (N_5502,N_5279,N_5209);
nor U5503 (N_5503,N_5314,N_5244);
nand U5504 (N_5504,N_5297,N_5380);
or U5505 (N_5505,N_5205,N_5395);
nor U5506 (N_5506,N_5266,N_5389);
xnor U5507 (N_5507,N_5245,N_5355);
and U5508 (N_5508,N_5201,N_5398);
nor U5509 (N_5509,N_5303,N_5216);
xnor U5510 (N_5510,N_5247,N_5391);
nand U5511 (N_5511,N_5355,N_5316);
and U5512 (N_5512,N_5256,N_5333);
nor U5513 (N_5513,N_5264,N_5341);
nand U5514 (N_5514,N_5239,N_5332);
nor U5515 (N_5515,N_5364,N_5238);
and U5516 (N_5516,N_5386,N_5322);
and U5517 (N_5517,N_5305,N_5236);
and U5518 (N_5518,N_5351,N_5368);
or U5519 (N_5519,N_5295,N_5282);
and U5520 (N_5520,N_5362,N_5375);
and U5521 (N_5521,N_5359,N_5319);
or U5522 (N_5522,N_5288,N_5300);
nand U5523 (N_5523,N_5239,N_5307);
nand U5524 (N_5524,N_5256,N_5259);
and U5525 (N_5525,N_5391,N_5390);
and U5526 (N_5526,N_5375,N_5345);
nor U5527 (N_5527,N_5225,N_5342);
nand U5528 (N_5528,N_5259,N_5264);
nand U5529 (N_5529,N_5345,N_5214);
nand U5530 (N_5530,N_5234,N_5321);
or U5531 (N_5531,N_5380,N_5223);
nor U5532 (N_5532,N_5252,N_5240);
nor U5533 (N_5533,N_5358,N_5394);
xor U5534 (N_5534,N_5290,N_5374);
or U5535 (N_5535,N_5369,N_5268);
or U5536 (N_5536,N_5397,N_5352);
nor U5537 (N_5537,N_5230,N_5301);
xor U5538 (N_5538,N_5394,N_5250);
and U5539 (N_5539,N_5312,N_5370);
nand U5540 (N_5540,N_5220,N_5367);
or U5541 (N_5541,N_5265,N_5234);
xnor U5542 (N_5542,N_5327,N_5227);
or U5543 (N_5543,N_5311,N_5343);
nand U5544 (N_5544,N_5324,N_5284);
and U5545 (N_5545,N_5307,N_5320);
and U5546 (N_5546,N_5262,N_5307);
nand U5547 (N_5547,N_5301,N_5240);
nor U5548 (N_5548,N_5330,N_5338);
or U5549 (N_5549,N_5383,N_5259);
xnor U5550 (N_5550,N_5312,N_5365);
xor U5551 (N_5551,N_5261,N_5209);
and U5552 (N_5552,N_5260,N_5398);
nand U5553 (N_5553,N_5298,N_5344);
xnor U5554 (N_5554,N_5312,N_5327);
xnor U5555 (N_5555,N_5271,N_5206);
or U5556 (N_5556,N_5207,N_5300);
nor U5557 (N_5557,N_5271,N_5341);
nand U5558 (N_5558,N_5317,N_5318);
xnor U5559 (N_5559,N_5382,N_5315);
xnor U5560 (N_5560,N_5387,N_5312);
or U5561 (N_5561,N_5203,N_5204);
xor U5562 (N_5562,N_5372,N_5254);
or U5563 (N_5563,N_5335,N_5299);
and U5564 (N_5564,N_5355,N_5225);
and U5565 (N_5565,N_5247,N_5336);
nor U5566 (N_5566,N_5319,N_5324);
or U5567 (N_5567,N_5372,N_5321);
xor U5568 (N_5568,N_5204,N_5356);
nor U5569 (N_5569,N_5266,N_5363);
nand U5570 (N_5570,N_5234,N_5270);
nand U5571 (N_5571,N_5330,N_5328);
or U5572 (N_5572,N_5236,N_5274);
nor U5573 (N_5573,N_5275,N_5216);
or U5574 (N_5574,N_5302,N_5317);
nand U5575 (N_5575,N_5215,N_5374);
xnor U5576 (N_5576,N_5217,N_5219);
or U5577 (N_5577,N_5216,N_5295);
or U5578 (N_5578,N_5238,N_5215);
nand U5579 (N_5579,N_5296,N_5271);
nor U5580 (N_5580,N_5210,N_5398);
or U5581 (N_5581,N_5259,N_5261);
xor U5582 (N_5582,N_5340,N_5248);
nor U5583 (N_5583,N_5246,N_5325);
nor U5584 (N_5584,N_5254,N_5276);
nand U5585 (N_5585,N_5271,N_5244);
and U5586 (N_5586,N_5293,N_5235);
or U5587 (N_5587,N_5289,N_5372);
xnor U5588 (N_5588,N_5332,N_5329);
and U5589 (N_5589,N_5272,N_5253);
xor U5590 (N_5590,N_5306,N_5213);
xor U5591 (N_5591,N_5204,N_5290);
nand U5592 (N_5592,N_5301,N_5208);
nand U5593 (N_5593,N_5310,N_5321);
nor U5594 (N_5594,N_5289,N_5259);
xor U5595 (N_5595,N_5249,N_5369);
nand U5596 (N_5596,N_5224,N_5278);
nand U5597 (N_5597,N_5340,N_5228);
xor U5598 (N_5598,N_5263,N_5219);
and U5599 (N_5599,N_5207,N_5341);
xor U5600 (N_5600,N_5445,N_5570);
nor U5601 (N_5601,N_5444,N_5536);
xor U5602 (N_5602,N_5521,N_5429);
and U5603 (N_5603,N_5526,N_5517);
or U5604 (N_5604,N_5494,N_5557);
xnor U5605 (N_5605,N_5486,N_5491);
xor U5606 (N_5606,N_5578,N_5589);
nand U5607 (N_5607,N_5558,N_5453);
xor U5608 (N_5608,N_5461,N_5477);
nor U5609 (N_5609,N_5545,N_5468);
and U5610 (N_5610,N_5503,N_5534);
nand U5611 (N_5611,N_5513,N_5406);
nand U5612 (N_5612,N_5411,N_5502);
xor U5613 (N_5613,N_5455,N_5581);
or U5614 (N_5614,N_5451,N_5405);
and U5615 (N_5615,N_5520,N_5562);
xnor U5616 (N_5616,N_5572,N_5438);
xnor U5617 (N_5617,N_5554,N_5481);
nor U5618 (N_5618,N_5447,N_5504);
and U5619 (N_5619,N_5431,N_5478);
and U5620 (N_5620,N_5579,N_5548);
nor U5621 (N_5621,N_5404,N_5592);
or U5622 (N_5622,N_5428,N_5518);
xnor U5623 (N_5623,N_5416,N_5482);
nand U5624 (N_5624,N_5496,N_5500);
nor U5625 (N_5625,N_5532,N_5471);
xor U5626 (N_5626,N_5435,N_5493);
nand U5627 (N_5627,N_5470,N_5439);
or U5628 (N_5628,N_5530,N_5559);
xor U5629 (N_5629,N_5459,N_5465);
or U5630 (N_5630,N_5522,N_5417);
and U5631 (N_5631,N_5423,N_5582);
xnor U5632 (N_5632,N_5452,N_5550);
nand U5633 (N_5633,N_5514,N_5485);
and U5634 (N_5634,N_5499,N_5539);
or U5635 (N_5635,N_5599,N_5408);
or U5636 (N_5636,N_5489,N_5402);
nand U5637 (N_5637,N_5487,N_5546);
or U5638 (N_5638,N_5426,N_5583);
and U5639 (N_5639,N_5531,N_5421);
nand U5640 (N_5640,N_5458,N_5432);
xor U5641 (N_5641,N_5565,N_5525);
xnor U5642 (N_5642,N_5454,N_5412);
nand U5643 (N_5643,N_5446,N_5456);
nor U5644 (N_5644,N_5541,N_5538);
and U5645 (N_5645,N_5568,N_5529);
nand U5646 (N_5646,N_5556,N_5480);
and U5647 (N_5647,N_5574,N_5555);
xor U5648 (N_5648,N_5575,N_5442);
and U5649 (N_5649,N_5498,N_5424);
xor U5650 (N_5650,N_5597,N_5449);
xor U5651 (N_5651,N_5472,N_5511);
and U5652 (N_5652,N_5528,N_5501);
and U5653 (N_5653,N_5587,N_5418);
nor U5654 (N_5654,N_5516,N_5507);
or U5655 (N_5655,N_5586,N_5591);
nand U5656 (N_5656,N_5523,N_5549);
nor U5657 (N_5657,N_5596,N_5422);
nor U5658 (N_5658,N_5593,N_5410);
xnor U5659 (N_5659,N_5457,N_5588);
nand U5660 (N_5660,N_5505,N_5595);
nand U5661 (N_5661,N_5508,N_5547);
xor U5662 (N_5662,N_5544,N_5497);
or U5663 (N_5663,N_5403,N_5488);
and U5664 (N_5664,N_5473,N_5483);
nand U5665 (N_5665,N_5543,N_5484);
nand U5666 (N_5666,N_5537,N_5474);
and U5667 (N_5667,N_5509,N_5479);
nand U5668 (N_5668,N_5475,N_5467);
and U5669 (N_5669,N_5492,N_5527);
and U5670 (N_5670,N_5464,N_5419);
nor U5671 (N_5671,N_5535,N_5512);
or U5672 (N_5672,N_5407,N_5466);
and U5673 (N_5673,N_5437,N_5524);
and U5674 (N_5674,N_5434,N_5564);
nor U5675 (N_5675,N_5571,N_5552);
and U5676 (N_5676,N_5413,N_5510);
xnor U5677 (N_5677,N_5409,N_5450);
nand U5678 (N_5678,N_5427,N_5580);
xor U5679 (N_5679,N_5573,N_5433);
xor U5680 (N_5680,N_5576,N_5490);
nor U5681 (N_5681,N_5569,N_5495);
nor U5682 (N_5682,N_5440,N_5430);
nor U5683 (N_5683,N_5561,N_5414);
xnor U5684 (N_5684,N_5506,N_5560);
nor U5685 (N_5685,N_5476,N_5401);
or U5686 (N_5686,N_5448,N_5567);
and U5687 (N_5687,N_5436,N_5515);
nor U5688 (N_5688,N_5463,N_5519);
nand U5689 (N_5689,N_5462,N_5563);
nand U5690 (N_5690,N_5425,N_5460);
xor U5691 (N_5691,N_5415,N_5594);
nor U5692 (N_5692,N_5598,N_5542);
and U5693 (N_5693,N_5577,N_5566);
or U5694 (N_5694,N_5551,N_5553);
or U5695 (N_5695,N_5585,N_5533);
and U5696 (N_5696,N_5584,N_5469);
or U5697 (N_5697,N_5400,N_5590);
and U5698 (N_5698,N_5443,N_5420);
nand U5699 (N_5699,N_5540,N_5441);
or U5700 (N_5700,N_5451,N_5472);
and U5701 (N_5701,N_5449,N_5550);
nor U5702 (N_5702,N_5437,N_5463);
xor U5703 (N_5703,N_5425,N_5555);
or U5704 (N_5704,N_5520,N_5557);
nor U5705 (N_5705,N_5415,N_5404);
or U5706 (N_5706,N_5478,N_5516);
and U5707 (N_5707,N_5561,N_5593);
xor U5708 (N_5708,N_5413,N_5562);
nor U5709 (N_5709,N_5548,N_5466);
and U5710 (N_5710,N_5542,N_5428);
and U5711 (N_5711,N_5416,N_5425);
nand U5712 (N_5712,N_5582,N_5593);
nand U5713 (N_5713,N_5461,N_5553);
nand U5714 (N_5714,N_5499,N_5428);
and U5715 (N_5715,N_5449,N_5544);
nand U5716 (N_5716,N_5580,N_5451);
nor U5717 (N_5717,N_5578,N_5428);
nor U5718 (N_5718,N_5563,N_5535);
and U5719 (N_5719,N_5533,N_5456);
or U5720 (N_5720,N_5574,N_5464);
and U5721 (N_5721,N_5522,N_5418);
or U5722 (N_5722,N_5401,N_5591);
or U5723 (N_5723,N_5502,N_5427);
nand U5724 (N_5724,N_5555,N_5594);
nor U5725 (N_5725,N_5553,N_5426);
or U5726 (N_5726,N_5554,N_5567);
or U5727 (N_5727,N_5546,N_5559);
nor U5728 (N_5728,N_5439,N_5475);
xor U5729 (N_5729,N_5546,N_5564);
or U5730 (N_5730,N_5431,N_5554);
and U5731 (N_5731,N_5518,N_5525);
or U5732 (N_5732,N_5578,N_5447);
nand U5733 (N_5733,N_5575,N_5425);
and U5734 (N_5734,N_5495,N_5473);
or U5735 (N_5735,N_5453,N_5565);
nor U5736 (N_5736,N_5504,N_5566);
and U5737 (N_5737,N_5557,N_5433);
and U5738 (N_5738,N_5436,N_5586);
xnor U5739 (N_5739,N_5456,N_5581);
xor U5740 (N_5740,N_5578,N_5497);
and U5741 (N_5741,N_5514,N_5421);
or U5742 (N_5742,N_5551,N_5440);
nor U5743 (N_5743,N_5554,N_5437);
nor U5744 (N_5744,N_5504,N_5441);
or U5745 (N_5745,N_5578,N_5556);
xor U5746 (N_5746,N_5477,N_5503);
and U5747 (N_5747,N_5583,N_5434);
xor U5748 (N_5748,N_5497,N_5549);
nand U5749 (N_5749,N_5597,N_5583);
nand U5750 (N_5750,N_5567,N_5565);
and U5751 (N_5751,N_5526,N_5567);
nor U5752 (N_5752,N_5419,N_5430);
xor U5753 (N_5753,N_5449,N_5572);
xnor U5754 (N_5754,N_5526,N_5557);
xor U5755 (N_5755,N_5409,N_5504);
nand U5756 (N_5756,N_5563,N_5521);
nand U5757 (N_5757,N_5530,N_5558);
or U5758 (N_5758,N_5416,N_5413);
or U5759 (N_5759,N_5468,N_5431);
nand U5760 (N_5760,N_5506,N_5488);
nor U5761 (N_5761,N_5597,N_5569);
xor U5762 (N_5762,N_5414,N_5411);
nor U5763 (N_5763,N_5592,N_5500);
and U5764 (N_5764,N_5501,N_5503);
nor U5765 (N_5765,N_5492,N_5599);
or U5766 (N_5766,N_5488,N_5518);
xnor U5767 (N_5767,N_5510,N_5486);
nor U5768 (N_5768,N_5407,N_5442);
nor U5769 (N_5769,N_5566,N_5576);
and U5770 (N_5770,N_5479,N_5520);
nor U5771 (N_5771,N_5489,N_5583);
xor U5772 (N_5772,N_5569,N_5501);
or U5773 (N_5773,N_5421,N_5577);
or U5774 (N_5774,N_5469,N_5541);
nand U5775 (N_5775,N_5533,N_5464);
nand U5776 (N_5776,N_5534,N_5459);
and U5777 (N_5777,N_5590,N_5592);
nand U5778 (N_5778,N_5493,N_5482);
or U5779 (N_5779,N_5467,N_5577);
or U5780 (N_5780,N_5523,N_5590);
nand U5781 (N_5781,N_5441,N_5506);
xnor U5782 (N_5782,N_5506,N_5562);
or U5783 (N_5783,N_5541,N_5572);
nor U5784 (N_5784,N_5588,N_5449);
and U5785 (N_5785,N_5502,N_5592);
nand U5786 (N_5786,N_5410,N_5452);
nor U5787 (N_5787,N_5433,N_5447);
nand U5788 (N_5788,N_5462,N_5416);
nor U5789 (N_5789,N_5430,N_5404);
nand U5790 (N_5790,N_5582,N_5404);
xnor U5791 (N_5791,N_5477,N_5481);
and U5792 (N_5792,N_5523,N_5468);
and U5793 (N_5793,N_5574,N_5487);
nor U5794 (N_5794,N_5429,N_5569);
nor U5795 (N_5795,N_5482,N_5429);
nor U5796 (N_5796,N_5426,N_5490);
nor U5797 (N_5797,N_5500,N_5442);
xnor U5798 (N_5798,N_5558,N_5555);
or U5799 (N_5799,N_5581,N_5541);
nor U5800 (N_5800,N_5617,N_5603);
and U5801 (N_5801,N_5699,N_5772);
or U5802 (N_5802,N_5633,N_5628);
xor U5803 (N_5803,N_5612,N_5718);
or U5804 (N_5804,N_5760,N_5719);
and U5805 (N_5805,N_5646,N_5622);
xor U5806 (N_5806,N_5717,N_5769);
xor U5807 (N_5807,N_5651,N_5744);
and U5808 (N_5808,N_5737,N_5711);
nor U5809 (N_5809,N_5792,N_5721);
nand U5810 (N_5810,N_5678,N_5654);
or U5811 (N_5811,N_5762,N_5706);
nand U5812 (N_5812,N_5667,N_5659);
or U5813 (N_5813,N_5673,N_5621);
nor U5814 (N_5814,N_5728,N_5606);
nand U5815 (N_5815,N_5668,N_5765);
xor U5816 (N_5816,N_5631,N_5784);
or U5817 (N_5817,N_5674,N_5790);
xor U5818 (N_5818,N_5695,N_5613);
xor U5819 (N_5819,N_5696,N_5641);
and U5820 (N_5820,N_5752,N_5627);
or U5821 (N_5821,N_5664,N_5618);
xor U5822 (N_5822,N_5708,N_5698);
nor U5823 (N_5823,N_5660,N_5796);
nor U5824 (N_5824,N_5670,N_5690);
or U5825 (N_5825,N_5649,N_5665);
and U5826 (N_5826,N_5643,N_5789);
xnor U5827 (N_5827,N_5632,N_5741);
and U5828 (N_5828,N_5686,N_5709);
xor U5829 (N_5829,N_5630,N_5683);
nand U5830 (N_5830,N_5733,N_5723);
and U5831 (N_5831,N_5757,N_5604);
xnor U5832 (N_5832,N_5747,N_5611);
nand U5833 (N_5833,N_5655,N_5600);
nand U5834 (N_5834,N_5773,N_5774);
xnor U5835 (N_5835,N_5701,N_5703);
nor U5836 (N_5836,N_5700,N_5602);
nor U5837 (N_5837,N_5626,N_5624);
xor U5838 (N_5838,N_5722,N_5710);
nand U5839 (N_5839,N_5745,N_5689);
and U5840 (N_5840,N_5743,N_5639);
nand U5841 (N_5841,N_5731,N_5608);
nand U5842 (N_5842,N_5691,N_5625);
nor U5843 (N_5843,N_5656,N_5637);
nand U5844 (N_5844,N_5672,N_5702);
and U5845 (N_5845,N_5730,N_5629);
or U5846 (N_5846,N_5799,N_5714);
xnor U5847 (N_5847,N_5669,N_5638);
nor U5848 (N_5848,N_5671,N_5761);
or U5849 (N_5849,N_5751,N_5783);
or U5850 (N_5850,N_5697,N_5692);
and U5851 (N_5851,N_5727,N_5739);
or U5852 (N_5852,N_5725,N_5785);
and U5853 (N_5853,N_5662,N_5687);
nand U5854 (N_5854,N_5610,N_5795);
nor U5855 (N_5855,N_5798,N_5750);
and U5856 (N_5856,N_5770,N_5647);
and U5857 (N_5857,N_5685,N_5734);
and U5858 (N_5858,N_5759,N_5793);
or U5859 (N_5859,N_5619,N_5766);
xor U5860 (N_5860,N_5688,N_5623);
nand U5861 (N_5861,N_5715,N_5712);
and U5862 (N_5862,N_5620,N_5694);
or U5863 (N_5863,N_5724,N_5726);
and U5864 (N_5864,N_5652,N_5636);
or U5865 (N_5865,N_5775,N_5729);
nand U5866 (N_5866,N_5609,N_5684);
nand U5867 (N_5867,N_5771,N_5782);
xnor U5868 (N_5868,N_5705,N_5615);
and U5869 (N_5869,N_5780,N_5680);
nor U5870 (N_5870,N_5681,N_5764);
xnor U5871 (N_5871,N_5661,N_5738);
and U5872 (N_5872,N_5776,N_5791);
or U5873 (N_5873,N_5679,N_5788);
nor U5874 (N_5874,N_5616,N_5794);
nand U5875 (N_5875,N_5736,N_5605);
xor U5876 (N_5876,N_5754,N_5735);
nor U5877 (N_5877,N_5634,N_5767);
or U5878 (N_5878,N_5644,N_5635);
or U5879 (N_5879,N_5642,N_5756);
xnor U5880 (N_5880,N_5707,N_5614);
and U5881 (N_5881,N_5716,N_5778);
nor U5882 (N_5882,N_5720,N_5653);
nand U5883 (N_5883,N_5749,N_5666);
nor U5884 (N_5884,N_5650,N_5677);
and U5885 (N_5885,N_5768,N_5779);
and U5886 (N_5886,N_5746,N_5763);
nand U5887 (N_5887,N_5607,N_5742);
or U5888 (N_5888,N_5601,N_5777);
nand U5889 (N_5889,N_5797,N_5675);
or U5890 (N_5890,N_5704,N_5781);
nor U5891 (N_5891,N_5682,N_5648);
and U5892 (N_5892,N_5740,N_5758);
or U5893 (N_5893,N_5658,N_5645);
and U5894 (N_5894,N_5748,N_5657);
nand U5895 (N_5895,N_5713,N_5753);
or U5896 (N_5896,N_5786,N_5693);
and U5897 (N_5897,N_5787,N_5640);
xor U5898 (N_5898,N_5732,N_5663);
and U5899 (N_5899,N_5755,N_5676);
or U5900 (N_5900,N_5736,N_5782);
xnor U5901 (N_5901,N_5628,N_5668);
nand U5902 (N_5902,N_5622,N_5735);
nand U5903 (N_5903,N_5787,N_5635);
or U5904 (N_5904,N_5752,N_5675);
nand U5905 (N_5905,N_5718,N_5676);
and U5906 (N_5906,N_5703,N_5793);
xor U5907 (N_5907,N_5723,N_5615);
nand U5908 (N_5908,N_5655,N_5665);
or U5909 (N_5909,N_5687,N_5600);
xor U5910 (N_5910,N_5719,N_5673);
nor U5911 (N_5911,N_5613,N_5655);
nand U5912 (N_5912,N_5787,N_5725);
nor U5913 (N_5913,N_5623,N_5771);
and U5914 (N_5914,N_5688,N_5704);
xor U5915 (N_5915,N_5734,N_5733);
nand U5916 (N_5916,N_5764,N_5714);
or U5917 (N_5917,N_5685,N_5758);
or U5918 (N_5918,N_5776,N_5637);
and U5919 (N_5919,N_5777,N_5722);
nor U5920 (N_5920,N_5639,N_5689);
nor U5921 (N_5921,N_5637,N_5715);
nor U5922 (N_5922,N_5622,N_5643);
nor U5923 (N_5923,N_5723,N_5757);
nor U5924 (N_5924,N_5783,N_5735);
nor U5925 (N_5925,N_5702,N_5657);
xnor U5926 (N_5926,N_5729,N_5601);
xor U5927 (N_5927,N_5626,N_5631);
or U5928 (N_5928,N_5786,N_5795);
nor U5929 (N_5929,N_5647,N_5745);
or U5930 (N_5930,N_5664,N_5686);
xnor U5931 (N_5931,N_5755,N_5678);
nor U5932 (N_5932,N_5703,N_5787);
or U5933 (N_5933,N_5642,N_5660);
and U5934 (N_5934,N_5648,N_5698);
or U5935 (N_5935,N_5719,N_5705);
or U5936 (N_5936,N_5755,N_5786);
xnor U5937 (N_5937,N_5683,N_5640);
or U5938 (N_5938,N_5722,N_5620);
or U5939 (N_5939,N_5742,N_5602);
nand U5940 (N_5940,N_5766,N_5667);
nand U5941 (N_5941,N_5719,N_5609);
nor U5942 (N_5942,N_5600,N_5776);
nor U5943 (N_5943,N_5615,N_5704);
nor U5944 (N_5944,N_5717,N_5601);
nor U5945 (N_5945,N_5669,N_5758);
xnor U5946 (N_5946,N_5766,N_5673);
nor U5947 (N_5947,N_5625,N_5623);
or U5948 (N_5948,N_5670,N_5752);
or U5949 (N_5949,N_5612,N_5774);
nand U5950 (N_5950,N_5659,N_5688);
nand U5951 (N_5951,N_5791,N_5715);
nand U5952 (N_5952,N_5669,N_5700);
nand U5953 (N_5953,N_5621,N_5725);
xnor U5954 (N_5954,N_5772,N_5621);
and U5955 (N_5955,N_5679,N_5627);
xnor U5956 (N_5956,N_5615,N_5646);
nand U5957 (N_5957,N_5652,N_5766);
nor U5958 (N_5958,N_5602,N_5756);
or U5959 (N_5959,N_5622,N_5798);
or U5960 (N_5960,N_5760,N_5602);
nor U5961 (N_5961,N_5757,N_5667);
xor U5962 (N_5962,N_5750,N_5616);
nand U5963 (N_5963,N_5633,N_5778);
nand U5964 (N_5964,N_5784,N_5712);
nand U5965 (N_5965,N_5622,N_5633);
and U5966 (N_5966,N_5712,N_5665);
and U5967 (N_5967,N_5636,N_5667);
or U5968 (N_5968,N_5794,N_5631);
and U5969 (N_5969,N_5650,N_5710);
xnor U5970 (N_5970,N_5668,N_5719);
xnor U5971 (N_5971,N_5600,N_5764);
or U5972 (N_5972,N_5738,N_5639);
nor U5973 (N_5973,N_5770,N_5661);
and U5974 (N_5974,N_5729,N_5694);
and U5975 (N_5975,N_5718,N_5622);
and U5976 (N_5976,N_5793,N_5700);
nor U5977 (N_5977,N_5736,N_5794);
xnor U5978 (N_5978,N_5693,N_5717);
xnor U5979 (N_5979,N_5762,N_5667);
nor U5980 (N_5980,N_5769,N_5766);
or U5981 (N_5981,N_5783,N_5707);
nor U5982 (N_5982,N_5609,N_5729);
nor U5983 (N_5983,N_5754,N_5786);
and U5984 (N_5984,N_5744,N_5660);
nor U5985 (N_5985,N_5681,N_5719);
and U5986 (N_5986,N_5703,N_5734);
nand U5987 (N_5987,N_5606,N_5704);
or U5988 (N_5988,N_5732,N_5737);
and U5989 (N_5989,N_5670,N_5663);
xor U5990 (N_5990,N_5733,N_5682);
nand U5991 (N_5991,N_5665,N_5793);
nand U5992 (N_5992,N_5604,N_5705);
nor U5993 (N_5993,N_5755,N_5631);
xor U5994 (N_5994,N_5738,N_5680);
nor U5995 (N_5995,N_5798,N_5663);
nand U5996 (N_5996,N_5660,N_5692);
or U5997 (N_5997,N_5727,N_5707);
nand U5998 (N_5998,N_5689,N_5616);
nor U5999 (N_5999,N_5633,N_5752);
and U6000 (N_6000,N_5838,N_5874);
xnor U6001 (N_6001,N_5820,N_5831);
or U6002 (N_6002,N_5960,N_5881);
nor U6003 (N_6003,N_5839,N_5912);
nor U6004 (N_6004,N_5855,N_5856);
and U6005 (N_6005,N_5919,N_5814);
or U6006 (N_6006,N_5893,N_5849);
and U6007 (N_6007,N_5827,N_5947);
xnor U6008 (N_6008,N_5823,N_5927);
nand U6009 (N_6009,N_5955,N_5869);
nand U6010 (N_6010,N_5964,N_5864);
or U6011 (N_6011,N_5997,N_5900);
xnor U6012 (N_6012,N_5819,N_5828);
nor U6013 (N_6013,N_5801,N_5981);
nand U6014 (N_6014,N_5929,N_5863);
nand U6015 (N_6015,N_5906,N_5805);
or U6016 (N_6016,N_5822,N_5809);
nand U6017 (N_6017,N_5816,N_5873);
and U6018 (N_6018,N_5815,N_5821);
or U6019 (N_6019,N_5980,N_5908);
xnor U6020 (N_6020,N_5860,N_5979);
xnor U6021 (N_6021,N_5800,N_5858);
or U6022 (N_6022,N_5969,N_5917);
and U6023 (N_6023,N_5833,N_5974);
or U6024 (N_6024,N_5852,N_5866);
nor U6025 (N_6025,N_5990,N_5968);
or U6026 (N_6026,N_5892,N_5931);
nor U6027 (N_6027,N_5899,N_5803);
and U6028 (N_6028,N_5930,N_5913);
nor U6029 (N_6029,N_5807,N_5950);
xor U6030 (N_6030,N_5896,N_5959);
and U6031 (N_6031,N_5826,N_5921);
nor U6032 (N_6032,N_5813,N_5802);
xor U6033 (N_6033,N_5998,N_5956);
xor U6034 (N_6034,N_5982,N_5905);
and U6035 (N_6035,N_5966,N_5907);
xor U6036 (N_6036,N_5859,N_5897);
or U6037 (N_6037,N_5918,N_5898);
xor U6038 (N_6038,N_5954,N_5992);
and U6039 (N_6039,N_5825,N_5817);
or U6040 (N_6040,N_5854,N_5967);
xor U6041 (N_6041,N_5901,N_5987);
nand U6042 (N_6042,N_5999,N_5888);
or U6043 (N_6043,N_5812,N_5943);
nand U6044 (N_6044,N_5984,N_5958);
xor U6045 (N_6045,N_5876,N_5951);
or U6046 (N_6046,N_5946,N_5953);
nand U6047 (N_6047,N_5887,N_5834);
or U6048 (N_6048,N_5840,N_5978);
nand U6049 (N_6049,N_5847,N_5940);
or U6050 (N_6050,N_5915,N_5845);
xor U6051 (N_6051,N_5861,N_5851);
xnor U6052 (N_6052,N_5890,N_5988);
and U6053 (N_6053,N_5832,N_5877);
xor U6054 (N_6054,N_5945,N_5884);
nor U6055 (N_6055,N_5808,N_5952);
xnor U6056 (N_6056,N_5848,N_5972);
nor U6057 (N_6057,N_5948,N_5867);
nand U6058 (N_6058,N_5975,N_5934);
nand U6059 (N_6059,N_5894,N_5875);
and U6060 (N_6060,N_5933,N_5976);
and U6061 (N_6061,N_5996,N_5830);
nand U6062 (N_6062,N_5936,N_5973);
nor U6063 (N_6063,N_5811,N_5885);
and U6064 (N_6064,N_5806,N_5920);
or U6065 (N_6065,N_5991,N_5882);
and U6066 (N_6066,N_5880,N_5895);
xnor U6067 (N_6067,N_5870,N_5911);
and U6068 (N_6068,N_5829,N_5886);
or U6069 (N_6069,N_5843,N_5824);
or U6070 (N_6070,N_5844,N_5846);
and U6071 (N_6071,N_5937,N_5970);
and U6072 (N_6072,N_5926,N_5928);
nand U6073 (N_6073,N_5957,N_5872);
nor U6074 (N_6074,N_5818,N_5914);
and U6075 (N_6075,N_5932,N_5889);
and U6076 (N_6076,N_5995,N_5902);
or U6077 (N_6077,N_5871,N_5965);
xnor U6078 (N_6078,N_5924,N_5850);
and U6079 (N_6079,N_5903,N_5842);
and U6080 (N_6080,N_5804,N_5939);
nor U6081 (N_6081,N_5922,N_5944);
nand U6082 (N_6082,N_5853,N_5986);
nand U6083 (N_6083,N_5923,N_5994);
xor U6084 (N_6084,N_5868,N_5941);
and U6085 (N_6085,N_5989,N_5862);
nor U6086 (N_6086,N_5942,N_5810);
xnor U6087 (N_6087,N_5891,N_5985);
xnor U6088 (N_6088,N_5836,N_5904);
or U6089 (N_6089,N_5878,N_5857);
and U6090 (N_6090,N_5909,N_5993);
nor U6091 (N_6091,N_5841,N_5835);
xnor U6092 (N_6092,N_5883,N_5938);
xor U6093 (N_6093,N_5910,N_5916);
and U6094 (N_6094,N_5963,N_5949);
nand U6095 (N_6095,N_5977,N_5935);
nand U6096 (N_6096,N_5962,N_5983);
xor U6097 (N_6097,N_5837,N_5925);
xnor U6098 (N_6098,N_5865,N_5961);
and U6099 (N_6099,N_5879,N_5971);
and U6100 (N_6100,N_5806,N_5895);
or U6101 (N_6101,N_5809,N_5880);
xor U6102 (N_6102,N_5971,N_5891);
and U6103 (N_6103,N_5952,N_5974);
and U6104 (N_6104,N_5960,N_5998);
nand U6105 (N_6105,N_5927,N_5879);
nand U6106 (N_6106,N_5925,N_5932);
or U6107 (N_6107,N_5866,N_5822);
or U6108 (N_6108,N_5816,N_5880);
or U6109 (N_6109,N_5802,N_5841);
nor U6110 (N_6110,N_5977,N_5822);
xor U6111 (N_6111,N_5912,N_5867);
xor U6112 (N_6112,N_5844,N_5987);
nor U6113 (N_6113,N_5945,N_5833);
nand U6114 (N_6114,N_5834,N_5922);
or U6115 (N_6115,N_5930,N_5907);
xor U6116 (N_6116,N_5907,N_5975);
nor U6117 (N_6117,N_5956,N_5903);
or U6118 (N_6118,N_5974,N_5804);
nand U6119 (N_6119,N_5924,N_5867);
and U6120 (N_6120,N_5919,N_5834);
xnor U6121 (N_6121,N_5916,N_5819);
nand U6122 (N_6122,N_5901,N_5866);
nor U6123 (N_6123,N_5950,N_5802);
xor U6124 (N_6124,N_5821,N_5972);
nand U6125 (N_6125,N_5866,N_5895);
xor U6126 (N_6126,N_5867,N_5805);
nand U6127 (N_6127,N_5889,N_5926);
nor U6128 (N_6128,N_5952,N_5876);
xnor U6129 (N_6129,N_5844,N_5807);
or U6130 (N_6130,N_5804,N_5896);
or U6131 (N_6131,N_5804,N_5887);
and U6132 (N_6132,N_5960,N_5900);
nor U6133 (N_6133,N_5910,N_5811);
or U6134 (N_6134,N_5859,N_5843);
and U6135 (N_6135,N_5810,N_5809);
or U6136 (N_6136,N_5846,N_5922);
nand U6137 (N_6137,N_5875,N_5829);
or U6138 (N_6138,N_5801,N_5941);
or U6139 (N_6139,N_5988,N_5936);
nor U6140 (N_6140,N_5803,N_5980);
nor U6141 (N_6141,N_5831,N_5818);
and U6142 (N_6142,N_5943,N_5843);
and U6143 (N_6143,N_5832,N_5947);
nor U6144 (N_6144,N_5842,N_5803);
xor U6145 (N_6145,N_5910,N_5953);
and U6146 (N_6146,N_5800,N_5883);
or U6147 (N_6147,N_5960,N_5878);
or U6148 (N_6148,N_5915,N_5925);
nand U6149 (N_6149,N_5926,N_5912);
nor U6150 (N_6150,N_5914,N_5840);
nand U6151 (N_6151,N_5883,N_5902);
nand U6152 (N_6152,N_5982,N_5932);
and U6153 (N_6153,N_5989,N_5988);
and U6154 (N_6154,N_5925,N_5909);
nand U6155 (N_6155,N_5936,N_5912);
xor U6156 (N_6156,N_5913,N_5876);
nor U6157 (N_6157,N_5845,N_5821);
xnor U6158 (N_6158,N_5869,N_5901);
and U6159 (N_6159,N_5859,N_5823);
nor U6160 (N_6160,N_5989,N_5955);
and U6161 (N_6161,N_5819,N_5858);
xor U6162 (N_6162,N_5927,N_5816);
nand U6163 (N_6163,N_5927,N_5815);
nor U6164 (N_6164,N_5811,N_5874);
nand U6165 (N_6165,N_5880,N_5995);
xor U6166 (N_6166,N_5878,N_5983);
nor U6167 (N_6167,N_5861,N_5922);
xor U6168 (N_6168,N_5836,N_5816);
nor U6169 (N_6169,N_5832,N_5810);
xnor U6170 (N_6170,N_5892,N_5994);
or U6171 (N_6171,N_5825,N_5885);
nor U6172 (N_6172,N_5956,N_5981);
xnor U6173 (N_6173,N_5952,N_5826);
nor U6174 (N_6174,N_5939,N_5850);
nand U6175 (N_6175,N_5986,N_5882);
nor U6176 (N_6176,N_5848,N_5858);
nand U6177 (N_6177,N_5905,N_5880);
and U6178 (N_6178,N_5979,N_5988);
or U6179 (N_6179,N_5963,N_5864);
or U6180 (N_6180,N_5964,N_5987);
nand U6181 (N_6181,N_5894,N_5946);
or U6182 (N_6182,N_5908,N_5976);
nand U6183 (N_6183,N_5843,N_5929);
nor U6184 (N_6184,N_5822,N_5936);
or U6185 (N_6185,N_5812,N_5894);
or U6186 (N_6186,N_5924,N_5835);
nor U6187 (N_6187,N_5854,N_5991);
xor U6188 (N_6188,N_5990,N_5974);
and U6189 (N_6189,N_5853,N_5988);
nand U6190 (N_6190,N_5979,N_5902);
xor U6191 (N_6191,N_5800,N_5965);
and U6192 (N_6192,N_5903,N_5914);
xnor U6193 (N_6193,N_5892,N_5930);
nor U6194 (N_6194,N_5999,N_5912);
nor U6195 (N_6195,N_5894,N_5831);
or U6196 (N_6196,N_5920,N_5847);
and U6197 (N_6197,N_5857,N_5899);
nand U6198 (N_6198,N_5889,N_5915);
and U6199 (N_6199,N_5921,N_5986);
nor U6200 (N_6200,N_6057,N_6029);
nand U6201 (N_6201,N_6026,N_6173);
or U6202 (N_6202,N_6030,N_6177);
nand U6203 (N_6203,N_6078,N_6009);
nand U6204 (N_6204,N_6188,N_6156);
nor U6205 (N_6205,N_6035,N_6012);
or U6206 (N_6206,N_6154,N_6043);
nand U6207 (N_6207,N_6124,N_6171);
nor U6208 (N_6208,N_6157,N_6048);
nor U6209 (N_6209,N_6070,N_6119);
and U6210 (N_6210,N_6041,N_6052);
nor U6211 (N_6211,N_6075,N_6165);
or U6212 (N_6212,N_6180,N_6102);
xnor U6213 (N_6213,N_6147,N_6169);
xnor U6214 (N_6214,N_6101,N_6187);
xnor U6215 (N_6215,N_6185,N_6120);
nor U6216 (N_6216,N_6051,N_6162);
or U6217 (N_6217,N_6056,N_6159);
or U6218 (N_6218,N_6079,N_6047);
nand U6219 (N_6219,N_6136,N_6142);
or U6220 (N_6220,N_6080,N_6045);
nor U6221 (N_6221,N_6135,N_6123);
nand U6222 (N_6222,N_6097,N_6150);
xnor U6223 (N_6223,N_6195,N_6151);
xor U6224 (N_6224,N_6103,N_6155);
nand U6225 (N_6225,N_6098,N_6131);
nand U6226 (N_6226,N_6110,N_6182);
nor U6227 (N_6227,N_6066,N_6107);
xor U6228 (N_6228,N_6065,N_6061);
or U6229 (N_6229,N_6170,N_6046);
or U6230 (N_6230,N_6090,N_6062);
and U6231 (N_6231,N_6022,N_6093);
xnor U6232 (N_6232,N_6067,N_6024);
xnor U6233 (N_6233,N_6160,N_6134);
and U6234 (N_6234,N_6161,N_6137);
or U6235 (N_6235,N_6094,N_6125);
xor U6236 (N_6236,N_6050,N_6001);
xor U6237 (N_6237,N_6194,N_6091);
and U6238 (N_6238,N_6121,N_6181);
xnor U6239 (N_6239,N_6002,N_6019);
xnor U6240 (N_6240,N_6081,N_6149);
nor U6241 (N_6241,N_6126,N_6084);
nor U6242 (N_6242,N_6192,N_6113);
nor U6243 (N_6243,N_6189,N_6072);
xor U6244 (N_6244,N_6018,N_6055);
or U6245 (N_6245,N_6143,N_6086);
nor U6246 (N_6246,N_6112,N_6031);
nor U6247 (N_6247,N_6087,N_6049);
xor U6248 (N_6248,N_6122,N_6015);
and U6249 (N_6249,N_6104,N_6039);
nor U6250 (N_6250,N_6006,N_6168);
nand U6251 (N_6251,N_6108,N_6138);
nand U6252 (N_6252,N_6083,N_6059);
xnor U6253 (N_6253,N_6077,N_6139);
or U6254 (N_6254,N_6000,N_6145);
and U6255 (N_6255,N_6127,N_6038);
nand U6256 (N_6256,N_6114,N_6141);
xnor U6257 (N_6257,N_6008,N_6088);
and U6258 (N_6258,N_6152,N_6128);
and U6259 (N_6259,N_6158,N_6199);
nand U6260 (N_6260,N_6146,N_6071);
xor U6261 (N_6261,N_6014,N_6144);
nand U6262 (N_6262,N_6186,N_6033);
nor U6263 (N_6263,N_6020,N_6054);
nor U6264 (N_6264,N_6028,N_6178);
nand U6265 (N_6265,N_6105,N_6118);
or U6266 (N_6266,N_6196,N_6004);
nand U6267 (N_6267,N_6025,N_6176);
xnor U6268 (N_6268,N_6089,N_6117);
nand U6269 (N_6269,N_6010,N_6184);
or U6270 (N_6270,N_6109,N_6191);
nand U6271 (N_6271,N_6116,N_6076);
and U6272 (N_6272,N_6044,N_6153);
or U6273 (N_6273,N_6198,N_6017);
nor U6274 (N_6274,N_6130,N_6063);
nand U6275 (N_6275,N_6034,N_6013);
or U6276 (N_6276,N_6174,N_6074);
nor U6277 (N_6277,N_6085,N_6092);
or U6278 (N_6278,N_6095,N_6197);
nor U6279 (N_6279,N_6007,N_6082);
or U6280 (N_6280,N_6140,N_6016);
xor U6281 (N_6281,N_6167,N_6129);
or U6282 (N_6282,N_6037,N_6100);
xor U6283 (N_6283,N_6106,N_6193);
or U6284 (N_6284,N_6099,N_6032);
nor U6285 (N_6285,N_6027,N_6166);
xnor U6286 (N_6286,N_6023,N_6053);
and U6287 (N_6287,N_6175,N_6069);
xor U6288 (N_6288,N_6133,N_6073);
nor U6289 (N_6289,N_6042,N_6068);
or U6290 (N_6290,N_6005,N_6164);
nand U6291 (N_6291,N_6060,N_6148);
and U6292 (N_6292,N_6003,N_6021);
nand U6293 (N_6293,N_6064,N_6183);
nor U6294 (N_6294,N_6096,N_6040);
nand U6295 (N_6295,N_6111,N_6058);
and U6296 (N_6296,N_6011,N_6179);
nor U6297 (N_6297,N_6132,N_6163);
and U6298 (N_6298,N_6190,N_6172);
nor U6299 (N_6299,N_6115,N_6036);
nand U6300 (N_6300,N_6178,N_6103);
and U6301 (N_6301,N_6114,N_6011);
nand U6302 (N_6302,N_6103,N_6140);
xnor U6303 (N_6303,N_6185,N_6050);
or U6304 (N_6304,N_6161,N_6036);
xnor U6305 (N_6305,N_6007,N_6124);
nor U6306 (N_6306,N_6153,N_6182);
nand U6307 (N_6307,N_6095,N_6011);
and U6308 (N_6308,N_6069,N_6164);
nor U6309 (N_6309,N_6037,N_6106);
nand U6310 (N_6310,N_6161,N_6075);
nor U6311 (N_6311,N_6066,N_6083);
nor U6312 (N_6312,N_6160,N_6138);
nand U6313 (N_6313,N_6030,N_6181);
xnor U6314 (N_6314,N_6104,N_6108);
xor U6315 (N_6315,N_6192,N_6142);
nor U6316 (N_6316,N_6097,N_6021);
or U6317 (N_6317,N_6077,N_6148);
and U6318 (N_6318,N_6187,N_6019);
nand U6319 (N_6319,N_6154,N_6010);
nor U6320 (N_6320,N_6162,N_6060);
xor U6321 (N_6321,N_6147,N_6141);
or U6322 (N_6322,N_6014,N_6038);
nor U6323 (N_6323,N_6061,N_6033);
or U6324 (N_6324,N_6072,N_6108);
and U6325 (N_6325,N_6003,N_6058);
nand U6326 (N_6326,N_6020,N_6171);
xnor U6327 (N_6327,N_6189,N_6127);
xnor U6328 (N_6328,N_6146,N_6042);
nand U6329 (N_6329,N_6188,N_6118);
and U6330 (N_6330,N_6128,N_6088);
nor U6331 (N_6331,N_6018,N_6195);
and U6332 (N_6332,N_6187,N_6074);
nand U6333 (N_6333,N_6086,N_6039);
nor U6334 (N_6334,N_6138,N_6176);
xor U6335 (N_6335,N_6011,N_6168);
nand U6336 (N_6336,N_6008,N_6080);
nand U6337 (N_6337,N_6115,N_6035);
xor U6338 (N_6338,N_6135,N_6051);
nor U6339 (N_6339,N_6045,N_6124);
and U6340 (N_6340,N_6007,N_6120);
nand U6341 (N_6341,N_6012,N_6013);
or U6342 (N_6342,N_6014,N_6185);
xor U6343 (N_6343,N_6056,N_6059);
or U6344 (N_6344,N_6124,N_6068);
and U6345 (N_6345,N_6128,N_6131);
nor U6346 (N_6346,N_6171,N_6045);
and U6347 (N_6347,N_6172,N_6149);
and U6348 (N_6348,N_6197,N_6007);
nand U6349 (N_6349,N_6168,N_6020);
nand U6350 (N_6350,N_6044,N_6134);
nand U6351 (N_6351,N_6109,N_6049);
or U6352 (N_6352,N_6108,N_6043);
nand U6353 (N_6353,N_6021,N_6031);
nor U6354 (N_6354,N_6168,N_6120);
nor U6355 (N_6355,N_6160,N_6081);
and U6356 (N_6356,N_6133,N_6006);
nand U6357 (N_6357,N_6015,N_6012);
xor U6358 (N_6358,N_6120,N_6110);
and U6359 (N_6359,N_6090,N_6023);
and U6360 (N_6360,N_6097,N_6027);
or U6361 (N_6361,N_6026,N_6110);
or U6362 (N_6362,N_6173,N_6134);
xnor U6363 (N_6363,N_6105,N_6171);
nand U6364 (N_6364,N_6117,N_6021);
nor U6365 (N_6365,N_6155,N_6076);
or U6366 (N_6366,N_6018,N_6179);
nor U6367 (N_6367,N_6081,N_6120);
nor U6368 (N_6368,N_6173,N_6023);
nand U6369 (N_6369,N_6135,N_6050);
nand U6370 (N_6370,N_6098,N_6130);
xor U6371 (N_6371,N_6135,N_6191);
nand U6372 (N_6372,N_6054,N_6082);
xor U6373 (N_6373,N_6080,N_6050);
xor U6374 (N_6374,N_6030,N_6067);
xnor U6375 (N_6375,N_6014,N_6005);
or U6376 (N_6376,N_6118,N_6040);
xor U6377 (N_6377,N_6091,N_6049);
nand U6378 (N_6378,N_6050,N_6196);
xor U6379 (N_6379,N_6037,N_6198);
and U6380 (N_6380,N_6038,N_6144);
or U6381 (N_6381,N_6061,N_6011);
or U6382 (N_6382,N_6079,N_6059);
or U6383 (N_6383,N_6030,N_6051);
or U6384 (N_6384,N_6148,N_6085);
or U6385 (N_6385,N_6140,N_6115);
or U6386 (N_6386,N_6157,N_6129);
nand U6387 (N_6387,N_6192,N_6029);
nand U6388 (N_6388,N_6180,N_6185);
or U6389 (N_6389,N_6152,N_6025);
nor U6390 (N_6390,N_6197,N_6028);
xor U6391 (N_6391,N_6105,N_6065);
xor U6392 (N_6392,N_6114,N_6128);
nor U6393 (N_6393,N_6157,N_6159);
or U6394 (N_6394,N_6195,N_6036);
xnor U6395 (N_6395,N_6127,N_6096);
or U6396 (N_6396,N_6124,N_6160);
nor U6397 (N_6397,N_6193,N_6025);
and U6398 (N_6398,N_6003,N_6075);
nor U6399 (N_6399,N_6037,N_6121);
and U6400 (N_6400,N_6399,N_6319);
and U6401 (N_6401,N_6263,N_6350);
nand U6402 (N_6402,N_6334,N_6243);
and U6403 (N_6403,N_6287,N_6310);
and U6404 (N_6404,N_6288,N_6228);
and U6405 (N_6405,N_6353,N_6273);
xor U6406 (N_6406,N_6214,N_6305);
or U6407 (N_6407,N_6386,N_6365);
or U6408 (N_6408,N_6380,N_6282);
nand U6409 (N_6409,N_6331,N_6314);
nand U6410 (N_6410,N_6206,N_6344);
and U6411 (N_6411,N_6240,N_6349);
nor U6412 (N_6412,N_6330,N_6359);
or U6413 (N_6413,N_6388,N_6378);
or U6414 (N_6414,N_6225,N_6213);
nand U6415 (N_6415,N_6355,N_6242);
xnor U6416 (N_6416,N_6318,N_6356);
nand U6417 (N_6417,N_6256,N_6286);
nor U6418 (N_6418,N_6204,N_6257);
or U6419 (N_6419,N_6221,N_6295);
nand U6420 (N_6420,N_6251,N_6384);
and U6421 (N_6421,N_6398,N_6338);
nor U6422 (N_6422,N_6259,N_6342);
nand U6423 (N_6423,N_6311,N_6245);
nand U6424 (N_6424,N_6304,N_6367);
and U6425 (N_6425,N_6397,N_6201);
xor U6426 (N_6426,N_6341,N_6274);
xnor U6427 (N_6427,N_6220,N_6396);
xor U6428 (N_6428,N_6382,N_6230);
xnor U6429 (N_6429,N_6200,N_6293);
nand U6430 (N_6430,N_6216,N_6373);
nand U6431 (N_6431,N_6209,N_6376);
xor U6432 (N_6432,N_6385,N_6300);
nor U6433 (N_6433,N_6390,N_6345);
and U6434 (N_6434,N_6312,N_6346);
nor U6435 (N_6435,N_6270,N_6258);
nand U6436 (N_6436,N_6358,N_6208);
nand U6437 (N_6437,N_6271,N_6381);
and U6438 (N_6438,N_6321,N_6351);
and U6439 (N_6439,N_6374,N_6361);
nand U6440 (N_6440,N_6244,N_6377);
nor U6441 (N_6441,N_6316,N_6223);
nor U6442 (N_6442,N_6227,N_6292);
nor U6443 (N_6443,N_6395,N_6336);
and U6444 (N_6444,N_6219,N_6275);
xnor U6445 (N_6445,N_6364,N_6348);
xnor U6446 (N_6446,N_6299,N_6352);
nor U6447 (N_6447,N_6301,N_6266);
nand U6448 (N_6448,N_6307,N_6335);
xnor U6449 (N_6449,N_6360,N_6264);
nand U6450 (N_6450,N_6339,N_6237);
or U6451 (N_6451,N_6327,N_6222);
nor U6452 (N_6452,N_6370,N_6366);
or U6453 (N_6453,N_6211,N_6290);
or U6454 (N_6454,N_6315,N_6302);
xnor U6455 (N_6455,N_6354,N_6248);
xnor U6456 (N_6456,N_6298,N_6332);
nand U6457 (N_6457,N_6328,N_6250);
nand U6458 (N_6458,N_6340,N_6393);
or U6459 (N_6459,N_6303,N_6323);
xor U6460 (N_6460,N_6389,N_6347);
nand U6461 (N_6461,N_6383,N_6372);
or U6462 (N_6462,N_6297,N_6379);
nand U6463 (N_6463,N_6260,N_6234);
nor U6464 (N_6464,N_6253,N_6278);
nor U6465 (N_6465,N_6255,N_6215);
xor U6466 (N_6466,N_6231,N_6369);
nand U6467 (N_6467,N_6229,N_6308);
or U6468 (N_6468,N_6313,N_6324);
nor U6469 (N_6469,N_6239,N_6212);
nand U6470 (N_6470,N_6261,N_6254);
or U6471 (N_6471,N_6357,N_6368);
xnor U6472 (N_6472,N_6247,N_6202);
and U6473 (N_6473,N_6277,N_6375);
nor U6474 (N_6474,N_6371,N_6337);
or U6475 (N_6475,N_6329,N_6363);
nand U6476 (N_6476,N_6265,N_6224);
xnor U6477 (N_6477,N_6238,N_6267);
or U6478 (N_6478,N_6235,N_6362);
and U6479 (N_6479,N_6217,N_6285);
xnor U6480 (N_6480,N_6268,N_6272);
xnor U6481 (N_6481,N_6317,N_6296);
xor U6482 (N_6482,N_6281,N_6284);
xor U6483 (N_6483,N_6262,N_6249);
or U6484 (N_6484,N_6333,N_6205);
and U6485 (N_6485,N_6322,N_6236);
xnor U6486 (N_6486,N_6252,N_6279);
nand U6487 (N_6487,N_6246,N_6241);
xnor U6488 (N_6488,N_6232,N_6291);
nand U6489 (N_6489,N_6320,N_6280);
nor U6490 (N_6490,N_6294,N_6276);
xnor U6491 (N_6491,N_6325,N_6218);
or U6492 (N_6492,N_6391,N_6210);
xnor U6493 (N_6493,N_6387,N_6269);
and U6494 (N_6494,N_6203,N_6283);
nand U6495 (N_6495,N_6309,N_6392);
nor U6496 (N_6496,N_6289,N_6226);
nor U6497 (N_6497,N_6233,N_6326);
xor U6498 (N_6498,N_6343,N_6306);
xnor U6499 (N_6499,N_6394,N_6207);
xnor U6500 (N_6500,N_6320,N_6325);
or U6501 (N_6501,N_6345,N_6381);
nor U6502 (N_6502,N_6228,N_6341);
nor U6503 (N_6503,N_6207,N_6223);
and U6504 (N_6504,N_6326,N_6339);
and U6505 (N_6505,N_6232,N_6351);
nor U6506 (N_6506,N_6304,N_6322);
nor U6507 (N_6507,N_6383,N_6279);
xnor U6508 (N_6508,N_6260,N_6253);
nor U6509 (N_6509,N_6315,N_6214);
xnor U6510 (N_6510,N_6331,N_6207);
and U6511 (N_6511,N_6371,N_6374);
nor U6512 (N_6512,N_6364,N_6217);
or U6513 (N_6513,N_6235,N_6316);
and U6514 (N_6514,N_6377,N_6203);
or U6515 (N_6515,N_6289,N_6292);
xnor U6516 (N_6516,N_6295,N_6207);
xnor U6517 (N_6517,N_6378,N_6394);
nor U6518 (N_6518,N_6206,N_6323);
and U6519 (N_6519,N_6342,N_6326);
xor U6520 (N_6520,N_6399,N_6340);
nor U6521 (N_6521,N_6338,N_6296);
and U6522 (N_6522,N_6221,N_6331);
nor U6523 (N_6523,N_6280,N_6386);
nor U6524 (N_6524,N_6338,N_6381);
nor U6525 (N_6525,N_6316,N_6380);
xnor U6526 (N_6526,N_6251,N_6398);
or U6527 (N_6527,N_6239,N_6363);
nor U6528 (N_6528,N_6238,N_6275);
nor U6529 (N_6529,N_6342,N_6210);
xnor U6530 (N_6530,N_6330,N_6335);
xnor U6531 (N_6531,N_6325,N_6265);
xnor U6532 (N_6532,N_6342,N_6257);
nand U6533 (N_6533,N_6296,N_6304);
or U6534 (N_6534,N_6218,N_6222);
nor U6535 (N_6535,N_6233,N_6377);
xnor U6536 (N_6536,N_6244,N_6259);
nand U6537 (N_6537,N_6228,N_6281);
xnor U6538 (N_6538,N_6263,N_6290);
and U6539 (N_6539,N_6203,N_6374);
nor U6540 (N_6540,N_6343,N_6369);
nor U6541 (N_6541,N_6386,N_6283);
and U6542 (N_6542,N_6397,N_6393);
nand U6543 (N_6543,N_6329,N_6301);
xnor U6544 (N_6544,N_6247,N_6336);
nor U6545 (N_6545,N_6230,N_6346);
or U6546 (N_6546,N_6268,N_6213);
xnor U6547 (N_6547,N_6333,N_6243);
and U6548 (N_6548,N_6264,N_6226);
and U6549 (N_6549,N_6347,N_6207);
nor U6550 (N_6550,N_6259,N_6203);
or U6551 (N_6551,N_6294,N_6389);
or U6552 (N_6552,N_6255,N_6296);
or U6553 (N_6553,N_6201,N_6203);
nor U6554 (N_6554,N_6284,N_6289);
xor U6555 (N_6555,N_6373,N_6298);
xnor U6556 (N_6556,N_6341,N_6269);
and U6557 (N_6557,N_6234,N_6392);
or U6558 (N_6558,N_6273,N_6275);
and U6559 (N_6559,N_6240,N_6336);
or U6560 (N_6560,N_6238,N_6247);
or U6561 (N_6561,N_6345,N_6233);
nor U6562 (N_6562,N_6370,N_6268);
or U6563 (N_6563,N_6334,N_6294);
xnor U6564 (N_6564,N_6389,N_6373);
nand U6565 (N_6565,N_6320,N_6247);
xnor U6566 (N_6566,N_6302,N_6249);
nand U6567 (N_6567,N_6308,N_6316);
xor U6568 (N_6568,N_6348,N_6392);
and U6569 (N_6569,N_6282,N_6296);
nand U6570 (N_6570,N_6346,N_6370);
xor U6571 (N_6571,N_6291,N_6246);
nor U6572 (N_6572,N_6221,N_6350);
or U6573 (N_6573,N_6308,N_6326);
nand U6574 (N_6574,N_6324,N_6296);
nor U6575 (N_6575,N_6275,N_6253);
or U6576 (N_6576,N_6319,N_6371);
nor U6577 (N_6577,N_6398,N_6271);
nand U6578 (N_6578,N_6224,N_6362);
and U6579 (N_6579,N_6211,N_6308);
xor U6580 (N_6580,N_6279,N_6205);
and U6581 (N_6581,N_6314,N_6258);
nand U6582 (N_6582,N_6319,N_6359);
nor U6583 (N_6583,N_6324,N_6342);
nand U6584 (N_6584,N_6377,N_6372);
nand U6585 (N_6585,N_6342,N_6320);
xnor U6586 (N_6586,N_6297,N_6207);
xnor U6587 (N_6587,N_6391,N_6356);
nand U6588 (N_6588,N_6226,N_6256);
nand U6589 (N_6589,N_6315,N_6326);
and U6590 (N_6590,N_6241,N_6260);
and U6591 (N_6591,N_6205,N_6374);
and U6592 (N_6592,N_6385,N_6361);
nand U6593 (N_6593,N_6215,N_6335);
or U6594 (N_6594,N_6209,N_6390);
xnor U6595 (N_6595,N_6294,N_6374);
or U6596 (N_6596,N_6319,N_6244);
nor U6597 (N_6597,N_6298,N_6235);
and U6598 (N_6598,N_6256,N_6371);
nand U6599 (N_6599,N_6375,N_6281);
xor U6600 (N_6600,N_6528,N_6438);
or U6601 (N_6601,N_6497,N_6534);
nor U6602 (N_6602,N_6410,N_6416);
nand U6603 (N_6603,N_6480,N_6421);
nor U6604 (N_6604,N_6446,N_6506);
nor U6605 (N_6605,N_6590,N_6594);
and U6606 (N_6606,N_6441,N_6427);
nor U6607 (N_6607,N_6569,N_6548);
or U6608 (N_6608,N_6495,N_6592);
or U6609 (N_6609,N_6434,N_6499);
nand U6610 (N_6610,N_6479,N_6512);
nand U6611 (N_6611,N_6537,N_6484);
or U6612 (N_6612,N_6567,N_6523);
nand U6613 (N_6613,N_6481,N_6545);
nor U6614 (N_6614,N_6544,N_6471);
nand U6615 (N_6615,N_6556,N_6496);
xnor U6616 (N_6616,N_6460,N_6500);
xor U6617 (N_6617,N_6470,N_6520);
and U6618 (N_6618,N_6587,N_6586);
and U6619 (N_6619,N_6559,N_6455);
and U6620 (N_6620,N_6541,N_6403);
and U6621 (N_6621,N_6475,N_6433);
or U6622 (N_6622,N_6498,N_6469);
and U6623 (N_6623,N_6596,N_6524);
xor U6624 (N_6624,N_6464,N_6447);
nand U6625 (N_6625,N_6593,N_6529);
or U6626 (N_6626,N_6412,N_6411);
or U6627 (N_6627,N_6458,N_6513);
xor U6628 (N_6628,N_6449,N_6597);
nand U6629 (N_6629,N_6409,N_6535);
nor U6630 (N_6630,N_6514,N_6511);
xor U6631 (N_6631,N_6502,N_6492);
nor U6632 (N_6632,N_6553,N_6473);
or U6633 (N_6633,N_6533,N_6404);
xnor U6634 (N_6634,N_6579,N_6443);
nand U6635 (N_6635,N_6482,N_6468);
nand U6636 (N_6636,N_6461,N_6422);
nor U6637 (N_6637,N_6562,N_6518);
xnor U6638 (N_6638,N_6550,N_6515);
xnor U6639 (N_6639,N_6530,N_6417);
and U6640 (N_6640,N_6531,N_6574);
nor U6641 (N_6641,N_6560,N_6572);
and U6642 (N_6642,N_6527,N_6565);
or U6643 (N_6643,N_6413,N_6580);
nor U6644 (N_6644,N_6542,N_6424);
nor U6645 (N_6645,N_6536,N_6488);
and U6646 (N_6646,N_6450,N_6486);
nand U6647 (N_6647,N_6476,N_6406);
nor U6648 (N_6648,N_6598,N_6442);
nor U6649 (N_6649,N_6564,N_6516);
nor U6650 (N_6650,N_6402,N_6576);
nand U6651 (N_6651,N_6563,N_6589);
xnor U6652 (N_6652,N_6440,N_6526);
nor U6653 (N_6653,N_6557,N_6570);
nor U6654 (N_6654,N_6477,N_6568);
nor U6655 (N_6655,N_6490,N_6507);
nand U6656 (N_6656,N_6547,N_6407);
xnor U6657 (N_6657,N_6444,N_6501);
nor U6658 (N_6658,N_6451,N_6505);
xnor U6659 (N_6659,N_6575,N_6400);
nand U6660 (N_6660,N_6466,N_6549);
or U6661 (N_6661,N_6430,N_6543);
and U6662 (N_6662,N_6573,N_6463);
or U6663 (N_6663,N_6493,N_6585);
and U6664 (N_6664,N_6510,N_6571);
xor U6665 (N_6665,N_6472,N_6418);
nand U6666 (N_6666,N_6561,N_6467);
xor U6667 (N_6667,N_6485,N_6452);
xnor U6668 (N_6668,N_6566,N_6432);
or U6669 (N_6669,N_6555,N_6423);
xor U6670 (N_6670,N_6405,N_6465);
xnor U6671 (N_6671,N_6551,N_6439);
or U6672 (N_6672,N_6436,N_6554);
xor U6673 (N_6673,N_6582,N_6532);
nor U6674 (N_6674,N_6503,N_6525);
xor U6675 (N_6675,N_6583,N_6504);
and U6676 (N_6676,N_6508,N_6429);
nor U6677 (N_6677,N_6431,N_6487);
and U6678 (N_6678,N_6415,N_6588);
nor U6679 (N_6679,N_6435,N_6595);
nor U6680 (N_6680,N_6577,N_6419);
and U6681 (N_6681,N_6578,N_6538);
nand U6682 (N_6682,N_6489,N_6509);
and U6683 (N_6683,N_6457,N_6519);
nor U6684 (N_6684,N_6420,N_6558);
xnor U6685 (N_6685,N_6474,N_6425);
xnor U6686 (N_6686,N_6540,N_6581);
and U6687 (N_6687,N_6483,N_6428);
and U6688 (N_6688,N_6426,N_6448);
nand U6689 (N_6689,N_6517,N_6591);
nor U6690 (N_6690,N_6459,N_6445);
or U6691 (N_6691,N_6437,N_6456);
nand U6692 (N_6692,N_6478,N_6552);
and U6693 (N_6693,N_6454,N_6539);
nor U6694 (N_6694,N_6408,N_6414);
nor U6695 (N_6695,N_6462,N_6453);
and U6696 (N_6696,N_6584,N_6494);
nor U6697 (N_6697,N_6599,N_6491);
nor U6698 (N_6698,N_6521,N_6401);
nand U6699 (N_6699,N_6546,N_6522);
nor U6700 (N_6700,N_6455,N_6414);
xor U6701 (N_6701,N_6438,N_6413);
xor U6702 (N_6702,N_6595,N_6529);
xor U6703 (N_6703,N_6476,N_6484);
and U6704 (N_6704,N_6485,N_6400);
nor U6705 (N_6705,N_6582,N_6466);
nand U6706 (N_6706,N_6409,N_6584);
xor U6707 (N_6707,N_6598,N_6501);
and U6708 (N_6708,N_6433,N_6412);
or U6709 (N_6709,N_6561,N_6571);
and U6710 (N_6710,N_6596,N_6547);
nor U6711 (N_6711,N_6405,N_6596);
nor U6712 (N_6712,N_6517,N_6542);
nand U6713 (N_6713,N_6577,N_6500);
and U6714 (N_6714,N_6455,N_6522);
nand U6715 (N_6715,N_6463,N_6586);
or U6716 (N_6716,N_6456,N_6508);
xnor U6717 (N_6717,N_6548,N_6592);
or U6718 (N_6718,N_6443,N_6459);
nand U6719 (N_6719,N_6544,N_6458);
nor U6720 (N_6720,N_6562,N_6564);
nand U6721 (N_6721,N_6504,N_6410);
nand U6722 (N_6722,N_6443,N_6572);
or U6723 (N_6723,N_6556,N_6451);
and U6724 (N_6724,N_6474,N_6458);
xnor U6725 (N_6725,N_6505,N_6422);
and U6726 (N_6726,N_6579,N_6486);
or U6727 (N_6727,N_6456,N_6488);
and U6728 (N_6728,N_6428,N_6554);
and U6729 (N_6729,N_6498,N_6472);
nand U6730 (N_6730,N_6444,N_6428);
xnor U6731 (N_6731,N_6413,N_6409);
xor U6732 (N_6732,N_6426,N_6444);
xnor U6733 (N_6733,N_6594,N_6465);
nor U6734 (N_6734,N_6487,N_6455);
xnor U6735 (N_6735,N_6401,N_6578);
xnor U6736 (N_6736,N_6430,N_6446);
xnor U6737 (N_6737,N_6457,N_6529);
nor U6738 (N_6738,N_6469,N_6455);
and U6739 (N_6739,N_6488,N_6415);
or U6740 (N_6740,N_6434,N_6470);
and U6741 (N_6741,N_6475,N_6412);
nor U6742 (N_6742,N_6533,N_6532);
xnor U6743 (N_6743,N_6466,N_6424);
nor U6744 (N_6744,N_6568,N_6476);
xor U6745 (N_6745,N_6583,N_6513);
xnor U6746 (N_6746,N_6569,N_6575);
nand U6747 (N_6747,N_6446,N_6537);
nand U6748 (N_6748,N_6525,N_6516);
nand U6749 (N_6749,N_6535,N_6578);
xnor U6750 (N_6750,N_6412,N_6565);
and U6751 (N_6751,N_6424,N_6496);
xor U6752 (N_6752,N_6444,N_6433);
nor U6753 (N_6753,N_6506,N_6556);
or U6754 (N_6754,N_6529,N_6446);
nand U6755 (N_6755,N_6520,N_6441);
nand U6756 (N_6756,N_6472,N_6438);
nor U6757 (N_6757,N_6422,N_6447);
and U6758 (N_6758,N_6430,N_6532);
or U6759 (N_6759,N_6446,N_6533);
nand U6760 (N_6760,N_6514,N_6469);
and U6761 (N_6761,N_6436,N_6584);
nor U6762 (N_6762,N_6445,N_6475);
xor U6763 (N_6763,N_6493,N_6579);
nor U6764 (N_6764,N_6506,N_6553);
xor U6765 (N_6765,N_6450,N_6439);
and U6766 (N_6766,N_6518,N_6452);
and U6767 (N_6767,N_6565,N_6563);
or U6768 (N_6768,N_6435,N_6500);
nor U6769 (N_6769,N_6539,N_6448);
and U6770 (N_6770,N_6548,N_6532);
and U6771 (N_6771,N_6407,N_6451);
nand U6772 (N_6772,N_6543,N_6499);
or U6773 (N_6773,N_6563,N_6504);
and U6774 (N_6774,N_6568,N_6419);
or U6775 (N_6775,N_6557,N_6580);
or U6776 (N_6776,N_6562,N_6537);
and U6777 (N_6777,N_6570,N_6588);
and U6778 (N_6778,N_6429,N_6425);
and U6779 (N_6779,N_6463,N_6530);
nand U6780 (N_6780,N_6588,N_6521);
nor U6781 (N_6781,N_6593,N_6530);
nand U6782 (N_6782,N_6532,N_6588);
and U6783 (N_6783,N_6408,N_6452);
nor U6784 (N_6784,N_6432,N_6553);
or U6785 (N_6785,N_6563,N_6468);
nor U6786 (N_6786,N_6425,N_6407);
or U6787 (N_6787,N_6574,N_6513);
or U6788 (N_6788,N_6429,N_6494);
nand U6789 (N_6789,N_6578,N_6464);
or U6790 (N_6790,N_6421,N_6565);
nor U6791 (N_6791,N_6414,N_6538);
and U6792 (N_6792,N_6513,N_6437);
and U6793 (N_6793,N_6452,N_6416);
xnor U6794 (N_6794,N_6430,N_6427);
and U6795 (N_6795,N_6542,N_6465);
and U6796 (N_6796,N_6484,N_6528);
and U6797 (N_6797,N_6465,N_6473);
or U6798 (N_6798,N_6405,N_6559);
or U6799 (N_6799,N_6587,N_6511);
or U6800 (N_6800,N_6638,N_6789);
xnor U6801 (N_6801,N_6695,N_6737);
nor U6802 (N_6802,N_6705,N_6669);
nand U6803 (N_6803,N_6693,N_6796);
xor U6804 (N_6804,N_6675,N_6655);
xnor U6805 (N_6805,N_6613,N_6702);
nor U6806 (N_6806,N_6624,N_6731);
and U6807 (N_6807,N_6630,N_6604);
nor U6808 (N_6808,N_6654,N_6696);
and U6809 (N_6809,N_6778,N_6685);
and U6810 (N_6810,N_6709,N_6661);
xnor U6811 (N_6811,N_6777,N_6622);
or U6812 (N_6812,N_6650,N_6707);
xnor U6813 (N_6813,N_6649,N_6674);
nor U6814 (N_6814,N_6615,N_6775);
and U6815 (N_6815,N_6752,N_6713);
or U6816 (N_6816,N_6714,N_6610);
and U6817 (N_6817,N_6670,N_6750);
and U6818 (N_6818,N_6697,N_6663);
nor U6819 (N_6819,N_6694,N_6761);
and U6820 (N_6820,N_6616,N_6758);
xnor U6821 (N_6821,N_6749,N_6751);
nand U6822 (N_6822,N_6739,N_6664);
nor U6823 (N_6823,N_6648,N_6641);
nor U6824 (N_6824,N_6771,N_6665);
nand U6825 (N_6825,N_6623,N_6733);
nand U6826 (N_6826,N_6619,N_6720);
xnor U6827 (N_6827,N_6755,N_6736);
nor U6828 (N_6828,N_6711,N_6620);
or U6829 (N_6829,N_6754,N_6687);
nor U6830 (N_6830,N_6688,N_6636);
nand U6831 (N_6831,N_6698,N_6717);
nor U6832 (N_6832,N_6635,N_6782);
xor U6833 (N_6833,N_6617,N_6745);
xnor U6834 (N_6834,N_6723,N_6643);
xor U6835 (N_6835,N_6657,N_6798);
nor U6836 (N_6836,N_6706,N_6639);
xor U6837 (N_6837,N_6652,N_6634);
or U6838 (N_6838,N_6601,N_6740);
nor U6839 (N_6839,N_6770,N_6708);
nand U6840 (N_6840,N_6759,N_6767);
xnor U6841 (N_6841,N_6797,N_6793);
or U6842 (N_6842,N_6779,N_6642);
or U6843 (N_6843,N_6600,N_6795);
or U6844 (N_6844,N_6757,N_6647);
nand U6845 (N_6845,N_6701,N_6774);
or U6846 (N_6846,N_6627,N_6732);
nand U6847 (N_6847,N_6728,N_6725);
and U6848 (N_6848,N_6710,N_6691);
and U6849 (N_6849,N_6676,N_6794);
nand U6850 (N_6850,N_6722,N_6718);
xnor U6851 (N_6851,N_6735,N_6662);
nor U6852 (N_6852,N_6791,N_6612);
nand U6853 (N_6853,N_6684,N_6632);
xnor U6854 (N_6854,N_6618,N_6605);
xor U6855 (N_6855,N_6776,N_6645);
or U6856 (N_6856,N_6656,N_6721);
nor U6857 (N_6857,N_6756,N_6764);
xnor U6858 (N_6858,N_6741,N_6672);
xnor U6859 (N_6859,N_6744,N_6788);
nand U6860 (N_6860,N_6727,N_6626);
nor U6861 (N_6861,N_6787,N_6773);
and U6862 (N_6862,N_6631,N_6673);
nand U6863 (N_6863,N_6699,N_6746);
nor U6864 (N_6864,N_6726,N_6785);
and U6865 (N_6865,N_6700,N_6667);
xor U6866 (N_6866,N_6609,N_6738);
xor U6867 (N_6867,N_6659,N_6747);
nor U6868 (N_6868,N_6651,N_6799);
nor U6869 (N_6869,N_6712,N_6671);
nand U6870 (N_6870,N_6792,N_6716);
or U6871 (N_6871,N_6780,N_6690);
or U6872 (N_6872,N_6781,N_6666);
nor U6873 (N_6873,N_6677,N_6633);
xnor U6874 (N_6874,N_6611,N_6682);
xor U6875 (N_6875,N_6719,N_6653);
nand U6876 (N_6876,N_6730,N_6640);
or U6877 (N_6877,N_6766,N_6603);
or U6878 (N_6878,N_6784,N_6724);
xor U6879 (N_6879,N_6762,N_6646);
xor U6880 (N_6880,N_6689,N_6790);
nor U6881 (N_6881,N_6692,N_6743);
or U6882 (N_6882,N_6742,N_6760);
and U6883 (N_6883,N_6769,N_6753);
or U6884 (N_6884,N_6763,N_6715);
and U6885 (N_6885,N_6765,N_6703);
nor U6886 (N_6886,N_6772,N_6658);
nand U6887 (N_6887,N_6606,N_6607);
nor U6888 (N_6888,N_6681,N_6614);
nand U6889 (N_6889,N_6734,N_6629);
or U6890 (N_6890,N_6786,N_6608);
nor U6891 (N_6891,N_6678,N_6686);
and U6892 (N_6892,N_6704,N_6628);
nor U6893 (N_6893,N_6680,N_6679);
nand U6894 (N_6894,N_6748,N_6637);
and U6895 (N_6895,N_6783,N_6602);
and U6896 (N_6896,N_6621,N_6729);
nor U6897 (N_6897,N_6683,N_6668);
xnor U6898 (N_6898,N_6644,N_6660);
nand U6899 (N_6899,N_6625,N_6768);
nor U6900 (N_6900,N_6697,N_6603);
nor U6901 (N_6901,N_6692,N_6718);
nor U6902 (N_6902,N_6673,N_6668);
xor U6903 (N_6903,N_6681,N_6691);
and U6904 (N_6904,N_6631,N_6610);
and U6905 (N_6905,N_6651,N_6705);
nor U6906 (N_6906,N_6745,N_6614);
nand U6907 (N_6907,N_6712,N_6689);
nor U6908 (N_6908,N_6773,N_6797);
and U6909 (N_6909,N_6722,N_6613);
nor U6910 (N_6910,N_6729,N_6643);
or U6911 (N_6911,N_6727,N_6614);
nand U6912 (N_6912,N_6639,N_6707);
xor U6913 (N_6913,N_6600,N_6604);
xor U6914 (N_6914,N_6709,N_6650);
or U6915 (N_6915,N_6647,N_6609);
nand U6916 (N_6916,N_6754,N_6625);
or U6917 (N_6917,N_6783,N_6629);
or U6918 (N_6918,N_6732,N_6769);
or U6919 (N_6919,N_6707,N_6734);
or U6920 (N_6920,N_6798,N_6689);
or U6921 (N_6921,N_6743,N_6661);
nor U6922 (N_6922,N_6628,N_6771);
and U6923 (N_6923,N_6795,N_6674);
or U6924 (N_6924,N_6722,N_6655);
and U6925 (N_6925,N_6784,N_6792);
and U6926 (N_6926,N_6621,N_6782);
nor U6927 (N_6927,N_6701,N_6749);
nor U6928 (N_6928,N_6715,N_6766);
or U6929 (N_6929,N_6760,N_6621);
xnor U6930 (N_6930,N_6617,N_6659);
or U6931 (N_6931,N_6783,N_6799);
nor U6932 (N_6932,N_6605,N_6691);
or U6933 (N_6933,N_6661,N_6613);
nor U6934 (N_6934,N_6638,N_6660);
and U6935 (N_6935,N_6744,N_6609);
and U6936 (N_6936,N_6714,N_6760);
and U6937 (N_6937,N_6728,N_6724);
xor U6938 (N_6938,N_6624,N_6748);
or U6939 (N_6939,N_6700,N_6724);
nor U6940 (N_6940,N_6707,N_6614);
xor U6941 (N_6941,N_6733,N_6704);
nor U6942 (N_6942,N_6789,N_6760);
nor U6943 (N_6943,N_6735,N_6642);
or U6944 (N_6944,N_6610,N_6782);
and U6945 (N_6945,N_6617,N_6675);
nand U6946 (N_6946,N_6728,N_6613);
and U6947 (N_6947,N_6694,N_6797);
nor U6948 (N_6948,N_6690,N_6728);
xnor U6949 (N_6949,N_6740,N_6691);
nor U6950 (N_6950,N_6746,N_6614);
or U6951 (N_6951,N_6669,N_6620);
and U6952 (N_6952,N_6652,N_6617);
nand U6953 (N_6953,N_6658,N_6773);
nor U6954 (N_6954,N_6621,N_6615);
and U6955 (N_6955,N_6623,N_6736);
and U6956 (N_6956,N_6680,N_6759);
and U6957 (N_6957,N_6715,N_6673);
or U6958 (N_6958,N_6605,N_6646);
nand U6959 (N_6959,N_6645,N_6716);
xnor U6960 (N_6960,N_6648,N_6660);
or U6961 (N_6961,N_6630,N_6734);
nand U6962 (N_6962,N_6624,N_6636);
xnor U6963 (N_6963,N_6665,N_6755);
nor U6964 (N_6964,N_6605,N_6663);
or U6965 (N_6965,N_6786,N_6687);
and U6966 (N_6966,N_6772,N_6790);
nor U6967 (N_6967,N_6646,N_6782);
xor U6968 (N_6968,N_6754,N_6770);
or U6969 (N_6969,N_6777,N_6750);
nand U6970 (N_6970,N_6772,N_6749);
nor U6971 (N_6971,N_6658,N_6720);
nor U6972 (N_6972,N_6742,N_6688);
or U6973 (N_6973,N_6736,N_6762);
and U6974 (N_6974,N_6757,N_6682);
and U6975 (N_6975,N_6646,N_6794);
nor U6976 (N_6976,N_6738,N_6623);
and U6977 (N_6977,N_6660,N_6769);
or U6978 (N_6978,N_6784,N_6664);
and U6979 (N_6979,N_6677,N_6783);
xor U6980 (N_6980,N_6690,N_6757);
nor U6981 (N_6981,N_6792,N_6621);
or U6982 (N_6982,N_6779,N_6773);
nor U6983 (N_6983,N_6606,N_6683);
nor U6984 (N_6984,N_6650,N_6793);
nor U6985 (N_6985,N_6679,N_6663);
and U6986 (N_6986,N_6740,N_6796);
nor U6987 (N_6987,N_6606,N_6649);
xor U6988 (N_6988,N_6663,N_6712);
and U6989 (N_6989,N_6636,N_6673);
nor U6990 (N_6990,N_6714,N_6697);
xnor U6991 (N_6991,N_6610,N_6732);
nor U6992 (N_6992,N_6697,N_6764);
nand U6993 (N_6993,N_6741,N_6762);
nand U6994 (N_6994,N_6614,N_6793);
and U6995 (N_6995,N_6645,N_6769);
and U6996 (N_6996,N_6635,N_6758);
or U6997 (N_6997,N_6729,N_6671);
xor U6998 (N_6998,N_6681,N_6626);
and U6999 (N_6999,N_6637,N_6656);
xnor U7000 (N_7000,N_6827,N_6875);
xor U7001 (N_7001,N_6872,N_6915);
nand U7002 (N_7002,N_6853,N_6837);
nand U7003 (N_7003,N_6836,N_6924);
nand U7004 (N_7004,N_6888,N_6809);
or U7005 (N_7005,N_6831,N_6971);
nand U7006 (N_7006,N_6974,N_6986);
nor U7007 (N_7007,N_6933,N_6873);
nand U7008 (N_7008,N_6860,N_6896);
nor U7009 (N_7009,N_6859,N_6877);
xnor U7010 (N_7010,N_6835,N_6995);
or U7011 (N_7011,N_6865,N_6893);
xor U7012 (N_7012,N_6814,N_6825);
nand U7013 (N_7013,N_6829,N_6997);
nor U7014 (N_7014,N_6891,N_6850);
or U7015 (N_7015,N_6930,N_6901);
or U7016 (N_7016,N_6921,N_6802);
and U7017 (N_7017,N_6903,N_6917);
nand U7018 (N_7018,N_6834,N_6938);
nand U7019 (N_7019,N_6838,N_6898);
or U7020 (N_7020,N_6929,N_6881);
nand U7021 (N_7021,N_6852,N_6922);
or U7022 (N_7022,N_6972,N_6812);
xor U7023 (N_7023,N_6902,N_6920);
nand U7024 (N_7024,N_6895,N_6975);
nand U7025 (N_7025,N_6887,N_6962);
and U7026 (N_7026,N_6937,N_6990);
and U7027 (N_7027,N_6886,N_6976);
or U7028 (N_7028,N_6956,N_6927);
nand U7029 (N_7029,N_6899,N_6978);
nor U7030 (N_7030,N_6925,N_6970);
nand U7031 (N_7031,N_6871,N_6818);
nand U7032 (N_7032,N_6800,N_6842);
and U7033 (N_7033,N_6806,N_6823);
nand U7034 (N_7034,N_6851,N_6841);
or U7035 (N_7035,N_6984,N_6979);
nand U7036 (N_7036,N_6821,N_6889);
nand U7037 (N_7037,N_6936,N_6856);
nand U7038 (N_7038,N_6843,N_6998);
xor U7039 (N_7039,N_6963,N_6819);
xor U7040 (N_7040,N_6828,N_6916);
xnor U7041 (N_7041,N_6897,N_6969);
nand U7042 (N_7042,N_6943,N_6992);
xnor U7043 (N_7043,N_6953,N_6878);
or U7044 (N_7044,N_6955,N_6954);
or U7045 (N_7045,N_6906,N_6876);
or U7046 (N_7046,N_6822,N_6869);
nand U7047 (N_7047,N_6805,N_6844);
nand U7048 (N_7048,N_6952,N_6833);
and U7049 (N_7049,N_6947,N_6968);
or U7050 (N_7050,N_6868,N_6914);
or U7051 (N_7051,N_6944,N_6830);
xor U7052 (N_7052,N_6857,N_6808);
xor U7053 (N_7053,N_6945,N_6950);
xor U7054 (N_7054,N_6973,N_6941);
and U7055 (N_7055,N_6863,N_6923);
or U7056 (N_7056,N_6867,N_6880);
xor U7057 (N_7057,N_6939,N_6918);
and U7058 (N_7058,N_6817,N_6824);
or U7059 (N_7059,N_6942,N_6839);
and U7060 (N_7060,N_6961,N_6988);
nand U7061 (N_7061,N_6816,N_6884);
xor U7062 (N_7062,N_6820,N_6855);
or U7063 (N_7063,N_6847,N_6928);
xor U7064 (N_7064,N_6949,N_6934);
or U7065 (N_7065,N_6815,N_6864);
nor U7066 (N_7066,N_6948,N_6967);
xor U7067 (N_7067,N_6892,N_6999);
xnor U7068 (N_7068,N_6980,N_6912);
nor U7069 (N_7069,N_6981,N_6894);
nand U7070 (N_7070,N_6882,N_6926);
and U7071 (N_7071,N_6958,N_6907);
xnor U7072 (N_7072,N_6813,N_6905);
or U7073 (N_7073,N_6803,N_6966);
nor U7074 (N_7074,N_6935,N_6885);
nand U7075 (N_7075,N_6832,N_6904);
or U7076 (N_7076,N_6861,N_6804);
nor U7077 (N_7077,N_6840,N_6879);
nor U7078 (N_7078,N_6957,N_6845);
nand U7079 (N_7079,N_6951,N_6870);
nor U7080 (N_7080,N_6807,N_6931);
and U7081 (N_7081,N_6913,N_6964);
or U7082 (N_7082,N_6874,N_6890);
and U7083 (N_7083,N_6900,N_6846);
nor U7084 (N_7084,N_6960,N_6977);
xnor U7085 (N_7085,N_6993,N_6959);
xor U7086 (N_7086,N_6996,N_6826);
xnor U7087 (N_7087,N_6932,N_6866);
or U7088 (N_7088,N_6989,N_6965);
and U7089 (N_7089,N_6983,N_6909);
nor U7090 (N_7090,N_6810,N_6848);
xnor U7091 (N_7091,N_6910,N_6940);
nor U7092 (N_7092,N_6854,N_6858);
xnor U7093 (N_7093,N_6946,N_6987);
nand U7094 (N_7094,N_6862,N_6919);
or U7095 (N_7095,N_6985,N_6908);
nor U7096 (N_7096,N_6991,N_6994);
and U7097 (N_7097,N_6883,N_6849);
or U7098 (N_7098,N_6811,N_6801);
nand U7099 (N_7099,N_6911,N_6982);
nand U7100 (N_7100,N_6944,N_6858);
and U7101 (N_7101,N_6875,N_6930);
and U7102 (N_7102,N_6980,N_6995);
nand U7103 (N_7103,N_6985,N_6860);
and U7104 (N_7104,N_6949,N_6992);
nor U7105 (N_7105,N_6917,N_6801);
nand U7106 (N_7106,N_6924,N_6831);
xnor U7107 (N_7107,N_6902,N_6911);
xor U7108 (N_7108,N_6871,N_6927);
nand U7109 (N_7109,N_6849,N_6858);
xor U7110 (N_7110,N_6978,N_6986);
nand U7111 (N_7111,N_6960,N_6985);
or U7112 (N_7112,N_6876,N_6800);
and U7113 (N_7113,N_6890,N_6974);
nand U7114 (N_7114,N_6882,N_6990);
and U7115 (N_7115,N_6863,N_6967);
xnor U7116 (N_7116,N_6977,N_6826);
and U7117 (N_7117,N_6905,N_6858);
xor U7118 (N_7118,N_6968,N_6856);
nor U7119 (N_7119,N_6815,N_6988);
nand U7120 (N_7120,N_6822,N_6868);
and U7121 (N_7121,N_6942,N_6929);
nor U7122 (N_7122,N_6924,N_6882);
xnor U7123 (N_7123,N_6855,N_6857);
or U7124 (N_7124,N_6818,N_6865);
or U7125 (N_7125,N_6878,N_6924);
and U7126 (N_7126,N_6867,N_6866);
nor U7127 (N_7127,N_6838,N_6802);
xnor U7128 (N_7128,N_6829,N_6837);
and U7129 (N_7129,N_6981,N_6895);
nand U7130 (N_7130,N_6956,N_6942);
and U7131 (N_7131,N_6864,N_6931);
nand U7132 (N_7132,N_6996,N_6984);
xnor U7133 (N_7133,N_6946,N_6836);
xor U7134 (N_7134,N_6939,N_6946);
and U7135 (N_7135,N_6901,N_6933);
or U7136 (N_7136,N_6836,N_6978);
nor U7137 (N_7137,N_6884,N_6876);
xor U7138 (N_7138,N_6813,N_6995);
nand U7139 (N_7139,N_6907,N_6868);
or U7140 (N_7140,N_6923,N_6818);
and U7141 (N_7141,N_6973,N_6889);
nand U7142 (N_7142,N_6918,N_6989);
or U7143 (N_7143,N_6910,N_6813);
xor U7144 (N_7144,N_6837,N_6970);
xor U7145 (N_7145,N_6947,N_6964);
xor U7146 (N_7146,N_6953,N_6963);
or U7147 (N_7147,N_6976,N_6937);
nand U7148 (N_7148,N_6841,N_6935);
nand U7149 (N_7149,N_6886,N_6849);
nand U7150 (N_7150,N_6822,N_6890);
xor U7151 (N_7151,N_6913,N_6837);
xor U7152 (N_7152,N_6934,N_6977);
xor U7153 (N_7153,N_6838,N_6952);
and U7154 (N_7154,N_6956,N_6941);
nand U7155 (N_7155,N_6989,N_6929);
nor U7156 (N_7156,N_6951,N_6868);
nor U7157 (N_7157,N_6962,N_6881);
xor U7158 (N_7158,N_6949,N_6873);
and U7159 (N_7159,N_6891,N_6942);
or U7160 (N_7160,N_6817,N_6906);
nand U7161 (N_7161,N_6897,N_6905);
and U7162 (N_7162,N_6994,N_6880);
nor U7163 (N_7163,N_6840,N_6970);
nor U7164 (N_7164,N_6894,N_6858);
or U7165 (N_7165,N_6897,N_6807);
nand U7166 (N_7166,N_6802,N_6988);
and U7167 (N_7167,N_6809,N_6918);
and U7168 (N_7168,N_6809,N_6865);
nor U7169 (N_7169,N_6862,N_6802);
xor U7170 (N_7170,N_6916,N_6871);
xor U7171 (N_7171,N_6861,N_6869);
xor U7172 (N_7172,N_6867,N_6821);
xor U7173 (N_7173,N_6968,N_6845);
and U7174 (N_7174,N_6917,N_6836);
or U7175 (N_7175,N_6921,N_6950);
nor U7176 (N_7176,N_6916,N_6882);
or U7177 (N_7177,N_6998,N_6947);
or U7178 (N_7178,N_6803,N_6928);
or U7179 (N_7179,N_6911,N_6907);
xor U7180 (N_7180,N_6927,N_6813);
and U7181 (N_7181,N_6844,N_6882);
nand U7182 (N_7182,N_6817,N_6822);
or U7183 (N_7183,N_6858,N_6877);
or U7184 (N_7184,N_6892,N_6906);
or U7185 (N_7185,N_6872,N_6821);
and U7186 (N_7186,N_6874,N_6812);
nand U7187 (N_7187,N_6991,N_6949);
nand U7188 (N_7188,N_6913,N_6937);
or U7189 (N_7189,N_6804,N_6882);
and U7190 (N_7190,N_6837,N_6966);
nand U7191 (N_7191,N_6830,N_6885);
and U7192 (N_7192,N_6916,N_6935);
and U7193 (N_7193,N_6958,N_6881);
nand U7194 (N_7194,N_6984,N_6869);
or U7195 (N_7195,N_6928,N_6827);
nand U7196 (N_7196,N_6926,N_6907);
and U7197 (N_7197,N_6919,N_6867);
and U7198 (N_7198,N_6950,N_6917);
nand U7199 (N_7199,N_6978,N_6871);
nor U7200 (N_7200,N_7091,N_7097);
nor U7201 (N_7201,N_7108,N_7122);
xnor U7202 (N_7202,N_7095,N_7126);
nor U7203 (N_7203,N_7060,N_7098);
and U7204 (N_7204,N_7109,N_7104);
and U7205 (N_7205,N_7088,N_7181);
and U7206 (N_7206,N_7103,N_7034);
xnor U7207 (N_7207,N_7090,N_7014);
nor U7208 (N_7208,N_7160,N_7050);
nor U7209 (N_7209,N_7128,N_7075);
xnor U7210 (N_7210,N_7172,N_7185);
nor U7211 (N_7211,N_7024,N_7120);
nand U7212 (N_7212,N_7116,N_7061);
nand U7213 (N_7213,N_7016,N_7033);
and U7214 (N_7214,N_7162,N_7038);
and U7215 (N_7215,N_7066,N_7106);
nor U7216 (N_7216,N_7112,N_7174);
nor U7217 (N_7217,N_7176,N_7115);
and U7218 (N_7218,N_7099,N_7123);
and U7219 (N_7219,N_7184,N_7030);
xor U7220 (N_7220,N_7022,N_7057);
nor U7221 (N_7221,N_7083,N_7187);
xor U7222 (N_7222,N_7025,N_7058);
nor U7223 (N_7223,N_7082,N_7002);
or U7224 (N_7224,N_7092,N_7020);
xor U7225 (N_7225,N_7144,N_7151);
nand U7226 (N_7226,N_7054,N_7149);
and U7227 (N_7227,N_7037,N_7188);
nor U7228 (N_7228,N_7093,N_7056);
xor U7229 (N_7229,N_7049,N_7031);
and U7230 (N_7230,N_7159,N_7035);
xnor U7231 (N_7231,N_7028,N_7044);
and U7232 (N_7232,N_7063,N_7130);
nand U7233 (N_7233,N_7124,N_7152);
or U7234 (N_7234,N_7113,N_7039);
or U7235 (N_7235,N_7011,N_7167);
and U7236 (N_7236,N_7125,N_7101);
xor U7237 (N_7237,N_7021,N_7196);
xor U7238 (N_7238,N_7146,N_7175);
or U7239 (N_7239,N_7043,N_7164);
or U7240 (N_7240,N_7086,N_7143);
nor U7241 (N_7241,N_7032,N_7111);
or U7242 (N_7242,N_7087,N_7163);
nand U7243 (N_7243,N_7094,N_7132);
nor U7244 (N_7244,N_7105,N_7154);
or U7245 (N_7245,N_7019,N_7141);
and U7246 (N_7246,N_7080,N_7085);
and U7247 (N_7247,N_7012,N_7138);
xnor U7248 (N_7248,N_7100,N_7195);
xor U7249 (N_7249,N_7147,N_7192);
nor U7250 (N_7250,N_7171,N_7073);
xor U7251 (N_7251,N_7003,N_7110);
nor U7252 (N_7252,N_7065,N_7046);
nor U7253 (N_7253,N_7169,N_7165);
nor U7254 (N_7254,N_7015,N_7183);
and U7255 (N_7255,N_7059,N_7077);
and U7256 (N_7256,N_7194,N_7047);
nor U7257 (N_7257,N_7179,N_7052);
and U7258 (N_7258,N_7070,N_7131);
or U7259 (N_7259,N_7153,N_7023);
nand U7260 (N_7260,N_7117,N_7155);
nor U7261 (N_7261,N_7158,N_7074);
xor U7262 (N_7262,N_7170,N_7157);
or U7263 (N_7263,N_7096,N_7089);
or U7264 (N_7264,N_7013,N_7142);
xor U7265 (N_7265,N_7026,N_7004);
xor U7266 (N_7266,N_7118,N_7027);
and U7267 (N_7267,N_7069,N_7114);
and U7268 (N_7268,N_7107,N_7051);
nor U7269 (N_7269,N_7168,N_7017);
and U7270 (N_7270,N_7199,N_7008);
xor U7271 (N_7271,N_7136,N_7177);
nor U7272 (N_7272,N_7180,N_7009);
nor U7273 (N_7273,N_7081,N_7129);
nand U7274 (N_7274,N_7048,N_7140);
xnor U7275 (N_7275,N_7000,N_7135);
and U7276 (N_7276,N_7166,N_7079);
or U7277 (N_7277,N_7150,N_7064);
or U7278 (N_7278,N_7040,N_7029);
and U7279 (N_7279,N_7053,N_7161);
nand U7280 (N_7280,N_7036,N_7055);
nand U7281 (N_7281,N_7084,N_7121);
and U7282 (N_7282,N_7178,N_7045);
nand U7283 (N_7283,N_7102,N_7197);
and U7284 (N_7284,N_7182,N_7190);
and U7285 (N_7285,N_7007,N_7134);
and U7286 (N_7286,N_7076,N_7078);
nand U7287 (N_7287,N_7018,N_7119);
xor U7288 (N_7288,N_7148,N_7041);
nand U7289 (N_7289,N_7137,N_7006);
xnor U7290 (N_7290,N_7198,N_7189);
xor U7291 (N_7291,N_7145,N_7193);
nand U7292 (N_7292,N_7139,N_7068);
nor U7293 (N_7293,N_7001,N_7186);
and U7294 (N_7294,N_7010,N_7191);
or U7295 (N_7295,N_7127,N_7062);
xnor U7296 (N_7296,N_7071,N_7005);
xnor U7297 (N_7297,N_7067,N_7173);
nor U7298 (N_7298,N_7042,N_7072);
xnor U7299 (N_7299,N_7133,N_7156);
nand U7300 (N_7300,N_7118,N_7100);
xor U7301 (N_7301,N_7084,N_7152);
or U7302 (N_7302,N_7060,N_7062);
xor U7303 (N_7303,N_7168,N_7050);
xnor U7304 (N_7304,N_7026,N_7010);
xnor U7305 (N_7305,N_7079,N_7021);
or U7306 (N_7306,N_7084,N_7043);
nor U7307 (N_7307,N_7096,N_7026);
nand U7308 (N_7308,N_7125,N_7126);
or U7309 (N_7309,N_7029,N_7088);
or U7310 (N_7310,N_7149,N_7128);
nand U7311 (N_7311,N_7175,N_7054);
xnor U7312 (N_7312,N_7038,N_7069);
xnor U7313 (N_7313,N_7004,N_7105);
nor U7314 (N_7314,N_7189,N_7003);
or U7315 (N_7315,N_7105,N_7050);
or U7316 (N_7316,N_7085,N_7155);
nand U7317 (N_7317,N_7056,N_7052);
and U7318 (N_7318,N_7117,N_7097);
nand U7319 (N_7319,N_7157,N_7188);
and U7320 (N_7320,N_7137,N_7174);
or U7321 (N_7321,N_7067,N_7151);
nor U7322 (N_7322,N_7032,N_7138);
nand U7323 (N_7323,N_7078,N_7165);
nor U7324 (N_7324,N_7168,N_7130);
nor U7325 (N_7325,N_7057,N_7088);
and U7326 (N_7326,N_7077,N_7156);
xnor U7327 (N_7327,N_7110,N_7024);
xnor U7328 (N_7328,N_7109,N_7010);
or U7329 (N_7329,N_7104,N_7123);
nand U7330 (N_7330,N_7071,N_7090);
nand U7331 (N_7331,N_7075,N_7094);
and U7332 (N_7332,N_7074,N_7005);
xnor U7333 (N_7333,N_7005,N_7114);
or U7334 (N_7334,N_7188,N_7194);
xor U7335 (N_7335,N_7175,N_7161);
nor U7336 (N_7336,N_7197,N_7146);
nor U7337 (N_7337,N_7113,N_7103);
or U7338 (N_7338,N_7094,N_7017);
or U7339 (N_7339,N_7001,N_7105);
and U7340 (N_7340,N_7170,N_7163);
nand U7341 (N_7341,N_7195,N_7012);
nand U7342 (N_7342,N_7085,N_7001);
nor U7343 (N_7343,N_7060,N_7028);
and U7344 (N_7344,N_7185,N_7093);
and U7345 (N_7345,N_7114,N_7133);
and U7346 (N_7346,N_7048,N_7060);
nand U7347 (N_7347,N_7165,N_7126);
and U7348 (N_7348,N_7002,N_7098);
xnor U7349 (N_7349,N_7175,N_7050);
nand U7350 (N_7350,N_7062,N_7131);
or U7351 (N_7351,N_7069,N_7011);
nand U7352 (N_7352,N_7118,N_7133);
and U7353 (N_7353,N_7187,N_7183);
or U7354 (N_7354,N_7128,N_7152);
xnor U7355 (N_7355,N_7136,N_7033);
nand U7356 (N_7356,N_7158,N_7082);
and U7357 (N_7357,N_7011,N_7173);
xor U7358 (N_7358,N_7087,N_7090);
or U7359 (N_7359,N_7177,N_7139);
nand U7360 (N_7360,N_7031,N_7076);
or U7361 (N_7361,N_7143,N_7192);
xnor U7362 (N_7362,N_7138,N_7011);
and U7363 (N_7363,N_7015,N_7000);
and U7364 (N_7364,N_7119,N_7006);
nor U7365 (N_7365,N_7062,N_7011);
or U7366 (N_7366,N_7174,N_7128);
xor U7367 (N_7367,N_7129,N_7011);
nor U7368 (N_7368,N_7098,N_7122);
or U7369 (N_7369,N_7091,N_7146);
nor U7370 (N_7370,N_7157,N_7186);
xor U7371 (N_7371,N_7015,N_7180);
nand U7372 (N_7372,N_7142,N_7039);
xnor U7373 (N_7373,N_7051,N_7104);
and U7374 (N_7374,N_7120,N_7134);
xnor U7375 (N_7375,N_7048,N_7152);
and U7376 (N_7376,N_7177,N_7180);
nor U7377 (N_7377,N_7195,N_7158);
nand U7378 (N_7378,N_7056,N_7133);
nand U7379 (N_7379,N_7042,N_7106);
nand U7380 (N_7380,N_7191,N_7186);
and U7381 (N_7381,N_7142,N_7005);
xnor U7382 (N_7382,N_7041,N_7161);
or U7383 (N_7383,N_7152,N_7166);
or U7384 (N_7384,N_7086,N_7176);
nor U7385 (N_7385,N_7186,N_7020);
nand U7386 (N_7386,N_7159,N_7041);
xnor U7387 (N_7387,N_7008,N_7152);
nand U7388 (N_7388,N_7147,N_7098);
nor U7389 (N_7389,N_7023,N_7149);
and U7390 (N_7390,N_7105,N_7115);
nand U7391 (N_7391,N_7017,N_7159);
nor U7392 (N_7392,N_7126,N_7119);
xnor U7393 (N_7393,N_7027,N_7040);
nand U7394 (N_7394,N_7179,N_7188);
nor U7395 (N_7395,N_7079,N_7042);
xnor U7396 (N_7396,N_7143,N_7044);
xor U7397 (N_7397,N_7155,N_7197);
xnor U7398 (N_7398,N_7189,N_7110);
nor U7399 (N_7399,N_7052,N_7198);
and U7400 (N_7400,N_7274,N_7320);
xnor U7401 (N_7401,N_7263,N_7232);
nor U7402 (N_7402,N_7265,N_7387);
xnor U7403 (N_7403,N_7377,N_7214);
nand U7404 (N_7404,N_7246,N_7375);
or U7405 (N_7405,N_7300,N_7391);
or U7406 (N_7406,N_7330,N_7213);
xor U7407 (N_7407,N_7336,N_7245);
xnor U7408 (N_7408,N_7249,N_7380);
nand U7409 (N_7409,N_7302,N_7363);
xor U7410 (N_7410,N_7399,N_7321);
or U7411 (N_7411,N_7224,N_7237);
nand U7412 (N_7412,N_7204,N_7212);
xor U7413 (N_7413,N_7386,N_7281);
and U7414 (N_7414,N_7311,N_7277);
and U7415 (N_7415,N_7240,N_7310);
and U7416 (N_7416,N_7325,N_7335);
nor U7417 (N_7417,N_7250,N_7373);
or U7418 (N_7418,N_7392,N_7307);
nand U7419 (N_7419,N_7372,N_7233);
nor U7420 (N_7420,N_7337,N_7364);
and U7421 (N_7421,N_7259,N_7266);
and U7422 (N_7422,N_7378,N_7286);
and U7423 (N_7423,N_7269,N_7275);
or U7424 (N_7424,N_7365,N_7201);
xnor U7425 (N_7425,N_7352,N_7394);
nor U7426 (N_7426,N_7206,N_7319);
or U7427 (N_7427,N_7264,N_7355);
nor U7428 (N_7428,N_7385,N_7296);
nor U7429 (N_7429,N_7228,N_7257);
or U7430 (N_7430,N_7345,N_7395);
nand U7431 (N_7431,N_7304,N_7223);
xor U7432 (N_7432,N_7348,N_7216);
nor U7433 (N_7433,N_7278,N_7203);
nor U7434 (N_7434,N_7288,N_7303);
nor U7435 (N_7435,N_7369,N_7272);
or U7436 (N_7436,N_7215,N_7258);
and U7437 (N_7437,N_7283,N_7273);
or U7438 (N_7438,N_7241,N_7368);
xor U7439 (N_7439,N_7255,N_7341);
xnor U7440 (N_7440,N_7267,N_7333);
nor U7441 (N_7441,N_7350,N_7343);
and U7442 (N_7442,N_7396,N_7353);
or U7443 (N_7443,N_7225,N_7316);
or U7444 (N_7444,N_7218,N_7211);
nand U7445 (N_7445,N_7293,N_7324);
nand U7446 (N_7446,N_7322,N_7299);
or U7447 (N_7447,N_7290,N_7226);
nor U7448 (N_7448,N_7270,N_7370);
or U7449 (N_7449,N_7313,N_7220);
or U7450 (N_7450,N_7243,N_7315);
nand U7451 (N_7451,N_7200,N_7309);
xor U7452 (N_7452,N_7292,N_7289);
nand U7453 (N_7453,N_7359,N_7217);
xnor U7454 (N_7454,N_7361,N_7235);
xor U7455 (N_7455,N_7236,N_7254);
nor U7456 (N_7456,N_7239,N_7287);
or U7457 (N_7457,N_7344,N_7398);
nor U7458 (N_7458,N_7338,N_7295);
or U7459 (N_7459,N_7230,N_7327);
or U7460 (N_7460,N_7271,N_7252);
nor U7461 (N_7461,N_7326,N_7358);
nand U7462 (N_7462,N_7347,N_7328);
xnor U7463 (N_7463,N_7314,N_7294);
or U7464 (N_7464,N_7374,N_7390);
or U7465 (N_7465,N_7312,N_7357);
or U7466 (N_7466,N_7388,N_7371);
or U7467 (N_7467,N_7356,N_7317);
and U7468 (N_7468,N_7329,N_7261);
and U7469 (N_7469,N_7279,N_7244);
and U7470 (N_7470,N_7334,N_7383);
and U7471 (N_7471,N_7382,N_7242);
nor U7472 (N_7472,N_7256,N_7339);
or U7473 (N_7473,N_7362,N_7284);
or U7474 (N_7474,N_7251,N_7367);
nor U7475 (N_7475,N_7205,N_7384);
or U7476 (N_7476,N_7210,N_7397);
xor U7477 (N_7477,N_7376,N_7209);
and U7478 (N_7478,N_7297,N_7219);
xor U7479 (N_7479,N_7360,N_7248);
xor U7480 (N_7480,N_7340,N_7238);
xor U7481 (N_7481,N_7262,N_7354);
xnor U7482 (N_7482,N_7332,N_7268);
or U7483 (N_7483,N_7282,N_7276);
xor U7484 (N_7484,N_7260,N_7305);
or U7485 (N_7485,N_7323,N_7253);
or U7486 (N_7486,N_7298,N_7342);
xnor U7487 (N_7487,N_7221,N_7285);
and U7488 (N_7488,N_7234,N_7280);
xnor U7489 (N_7489,N_7331,N_7222);
nor U7490 (N_7490,N_7381,N_7291);
or U7491 (N_7491,N_7306,N_7308);
and U7492 (N_7492,N_7247,N_7351);
and U7493 (N_7493,N_7208,N_7349);
xnor U7494 (N_7494,N_7379,N_7389);
nor U7495 (N_7495,N_7393,N_7366);
nor U7496 (N_7496,N_7227,N_7318);
xor U7497 (N_7497,N_7301,N_7346);
nand U7498 (N_7498,N_7207,N_7229);
xnor U7499 (N_7499,N_7202,N_7231);
nand U7500 (N_7500,N_7322,N_7332);
and U7501 (N_7501,N_7252,N_7300);
nor U7502 (N_7502,N_7236,N_7315);
xor U7503 (N_7503,N_7286,N_7293);
nor U7504 (N_7504,N_7288,N_7265);
nor U7505 (N_7505,N_7256,N_7315);
nor U7506 (N_7506,N_7237,N_7384);
xor U7507 (N_7507,N_7228,N_7390);
and U7508 (N_7508,N_7321,N_7290);
or U7509 (N_7509,N_7259,N_7379);
or U7510 (N_7510,N_7280,N_7347);
or U7511 (N_7511,N_7377,N_7386);
nor U7512 (N_7512,N_7248,N_7290);
or U7513 (N_7513,N_7224,N_7340);
and U7514 (N_7514,N_7283,N_7266);
xnor U7515 (N_7515,N_7215,N_7236);
and U7516 (N_7516,N_7336,N_7289);
xor U7517 (N_7517,N_7205,N_7268);
and U7518 (N_7518,N_7210,N_7227);
nor U7519 (N_7519,N_7315,N_7382);
nor U7520 (N_7520,N_7253,N_7219);
nand U7521 (N_7521,N_7236,N_7297);
nor U7522 (N_7522,N_7357,N_7346);
nand U7523 (N_7523,N_7266,N_7235);
and U7524 (N_7524,N_7367,N_7234);
nand U7525 (N_7525,N_7249,N_7279);
or U7526 (N_7526,N_7327,N_7338);
or U7527 (N_7527,N_7234,N_7324);
xnor U7528 (N_7528,N_7309,N_7330);
xnor U7529 (N_7529,N_7318,N_7201);
or U7530 (N_7530,N_7391,N_7246);
nor U7531 (N_7531,N_7294,N_7220);
nand U7532 (N_7532,N_7314,N_7352);
xor U7533 (N_7533,N_7360,N_7282);
or U7534 (N_7534,N_7200,N_7203);
nor U7535 (N_7535,N_7353,N_7358);
and U7536 (N_7536,N_7391,N_7388);
xor U7537 (N_7537,N_7218,N_7321);
nand U7538 (N_7538,N_7374,N_7335);
xor U7539 (N_7539,N_7341,N_7314);
or U7540 (N_7540,N_7209,N_7369);
and U7541 (N_7541,N_7305,N_7213);
nor U7542 (N_7542,N_7328,N_7389);
nand U7543 (N_7543,N_7276,N_7297);
nand U7544 (N_7544,N_7249,N_7319);
or U7545 (N_7545,N_7205,N_7372);
or U7546 (N_7546,N_7310,N_7331);
and U7547 (N_7547,N_7345,N_7245);
or U7548 (N_7548,N_7302,N_7200);
xor U7549 (N_7549,N_7235,N_7388);
xor U7550 (N_7550,N_7349,N_7215);
nand U7551 (N_7551,N_7324,N_7334);
or U7552 (N_7552,N_7396,N_7346);
nand U7553 (N_7553,N_7324,N_7254);
nor U7554 (N_7554,N_7364,N_7293);
nand U7555 (N_7555,N_7280,N_7323);
nand U7556 (N_7556,N_7354,N_7265);
and U7557 (N_7557,N_7382,N_7297);
and U7558 (N_7558,N_7230,N_7283);
xnor U7559 (N_7559,N_7200,N_7317);
xnor U7560 (N_7560,N_7325,N_7225);
or U7561 (N_7561,N_7204,N_7237);
or U7562 (N_7562,N_7223,N_7250);
and U7563 (N_7563,N_7317,N_7316);
nand U7564 (N_7564,N_7204,N_7230);
nand U7565 (N_7565,N_7335,N_7302);
nand U7566 (N_7566,N_7395,N_7298);
nor U7567 (N_7567,N_7264,N_7278);
nor U7568 (N_7568,N_7280,N_7228);
or U7569 (N_7569,N_7231,N_7304);
nor U7570 (N_7570,N_7284,N_7383);
nand U7571 (N_7571,N_7324,N_7233);
nand U7572 (N_7572,N_7232,N_7340);
or U7573 (N_7573,N_7397,N_7242);
and U7574 (N_7574,N_7368,N_7320);
nor U7575 (N_7575,N_7323,N_7285);
nand U7576 (N_7576,N_7200,N_7218);
and U7577 (N_7577,N_7213,N_7389);
xor U7578 (N_7578,N_7217,N_7327);
nor U7579 (N_7579,N_7386,N_7203);
nand U7580 (N_7580,N_7305,N_7323);
and U7581 (N_7581,N_7342,N_7271);
nor U7582 (N_7582,N_7278,N_7272);
or U7583 (N_7583,N_7291,N_7248);
nor U7584 (N_7584,N_7245,N_7236);
and U7585 (N_7585,N_7303,N_7339);
xnor U7586 (N_7586,N_7268,N_7386);
and U7587 (N_7587,N_7358,N_7369);
xor U7588 (N_7588,N_7320,N_7231);
or U7589 (N_7589,N_7380,N_7296);
nand U7590 (N_7590,N_7367,N_7226);
or U7591 (N_7591,N_7203,N_7356);
and U7592 (N_7592,N_7372,N_7259);
nand U7593 (N_7593,N_7354,N_7237);
nor U7594 (N_7594,N_7255,N_7232);
xor U7595 (N_7595,N_7307,N_7239);
xor U7596 (N_7596,N_7232,N_7213);
and U7597 (N_7597,N_7338,N_7306);
and U7598 (N_7598,N_7224,N_7354);
xor U7599 (N_7599,N_7305,N_7366);
nor U7600 (N_7600,N_7448,N_7410);
xnor U7601 (N_7601,N_7564,N_7403);
nand U7602 (N_7602,N_7504,N_7408);
and U7603 (N_7603,N_7434,N_7548);
xnor U7604 (N_7604,N_7498,N_7477);
nor U7605 (N_7605,N_7432,N_7509);
or U7606 (N_7606,N_7562,N_7417);
nor U7607 (N_7607,N_7453,N_7545);
nand U7608 (N_7608,N_7566,N_7522);
xnor U7609 (N_7609,N_7487,N_7428);
and U7610 (N_7610,N_7560,N_7518);
nor U7611 (N_7611,N_7430,N_7537);
nor U7612 (N_7612,N_7476,N_7494);
or U7613 (N_7613,N_7553,N_7482);
and U7614 (N_7614,N_7454,N_7473);
xor U7615 (N_7615,N_7508,N_7451);
or U7616 (N_7616,N_7593,N_7596);
and U7617 (N_7617,N_7563,N_7577);
xnor U7618 (N_7618,N_7456,N_7547);
or U7619 (N_7619,N_7471,N_7427);
nor U7620 (N_7620,N_7413,N_7507);
nor U7621 (N_7621,N_7586,N_7421);
and U7622 (N_7622,N_7503,N_7407);
nand U7623 (N_7623,N_7462,N_7524);
or U7624 (N_7624,N_7538,N_7557);
nand U7625 (N_7625,N_7543,N_7481);
nor U7626 (N_7626,N_7496,N_7419);
xnor U7627 (N_7627,N_7514,N_7485);
nand U7628 (N_7628,N_7574,N_7437);
and U7629 (N_7629,N_7597,N_7404);
nor U7630 (N_7630,N_7441,N_7549);
nor U7631 (N_7631,N_7591,N_7452);
nand U7632 (N_7632,N_7455,N_7478);
xor U7633 (N_7633,N_7429,N_7500);
or U7634 (N_7634,N_7449,N_7426);
xnor U7635 (N_7635,N_7540,N_7469);
nand U7636 (N_7636,N_7599,N_7412);
and U7637 (N_7637,N_7530,N_7536);
xor U7638 (N_7638,N_7531,N_7515);
nor U7639 (N_7639,N_7435,N_7554);
xnor U7640 (N_7640,N_7492,N_7550);
or U7641 (N_7641,N_7511,N_7439);
nor U7642 (N_7642,N_7489,N_7583);
nand U7643 (N_7643,N_7541,N_7458);
and U7644 (N_7644,N_7483,N_7443);
nand U7645 (N_7645,N_7587,N_7459);
xnor U7646 (N_7646,N_7400,N_7464);
or U7647 (N_7647,N_7474,N_7411);
or U7648 (N_7648,N_7472,N_7416);
nand U7649 (N_7649,N_7442,N_7495);
nand U7650 (N_7650,N_7488,N_7568);
or U7651 (N_7651,N_7431,N_7544);
nor U7652 (N_7652,N_7565,N_7497);
nor U7653 (N_7653,N_7516,N_7581);
xor U7654 (N_7654,N_7589,N_7571);
or U7655 (N_7655,N_7590,N_7552);
and U7656 (N_7656,N_7490,N_7491);
or U7657 (N_7657,N_7517,N_7539);
and U7658 (N_7658,N_7521,N_7493);
nor U7659 (N_7659,N_7460,N_7555);
and U7660 (N_7660,N_7512,N_7575);
nand U7661 (N_7661,N_7479,N_7450);
xnor U7662 (N_7662,N_7401,N_7466);
or U7663 (N_7663,N_7533,N_7422);
nand U7664 (N_7664,N_7440,N_7556);
and U7665 (N_7665,N_7424,N_7527);
or U7666 (N_7666,N_7570,N_7506);
and U7667 (N_7667,N_7510,N_7578);
nor U7668 (N_7668,N_7584,N_7480);
nand U7669 (N_7669,N_7519,N_7569);
xor U7670 (N_7670,N_7559,N_7461);
nor U7671 (N_7671,N_7470,N_7484);
and U7672 (N_7672,N_7501,N_7598);
xor U7673 (N_7673,N_7534,N_7582);
nand U7674 (N_7674,N_7580,N_7523);
xor U7675 (N_7675,N_7594,N_7423);
or U7676 (N_7676,N_7445,N_7468);
xnor U7677 (N_7677,N_7433,N_7588);
nor U7678 (N_7678,N_7457,N_7505);
and U7679 (N_7679,N_7595,N_7418);
and U7680 (N_7680,N_7551,N_7520);
and U7681 (N_7681,N_7513,N_7558);
nand U7682 (N_7682,N_7446,N_7532);
nor U7683 (N_7683,N_7528,N_7438);
nor U7684 (N_7684,N_7529,N_7526);
xor U7685 (N_7685,N_7502,N_7425);
xnor U7686 (N_7686,N_7415,N_7409);
and U7687 (N_7687,N_7535,N_7546);
xor U7688 (N_7688,N_7405,N_7585);
xor U7689 (N_7689,N_7592,N_7420);
xnor U7690 (N_7690,N_7567,N_7467);
nand U7691 (N_7691,N_7525,N_7573);
nor U7692 (N_7692,N_7402,N_7444);
nand U7693 (N_7693,N_7465,N_7463);
nand U7694 (N_7694,N_7436,N_7486);
nor U7695 (N_7695,N_7572,N_7561);
and U7696 (N_7696,N_7576,N_7542);
and U7697 (N_7697,N_7499,N_7579);
xnor U7698 (N_7698,N_7414,N_7447);
and U7699 (N_7699,N_7475,N_7406);
xor U7700 (N_7700,N_7474,N_7422);
nor U7701 (N_7701,N_7576,N_7454);
xor U7702 (N_7702,N_7442,N_7458);
nand U7703 (N_7703,N_7447,N_7583);
nor U7704 (N_7704,N_7425,N_7480);
and U7705 (N_7705,N_7431,N_7511);
nor U7706 (N_7706,N_7529,N_7425);
and U7707 (N_7707,N_7476,N_7527);
or U7708 (N_7708,N_7570,N_7481);
nor U7709 (N_7709,N_7404,N_7430);
or U7710 (N_7710,N_7489,N_7513);
nand U7711 (N_7711,N_7528,N_7597);
xnor U7712 (N_7712,N_7557,N_7556);
xor U7713 (N_7713,N_7570,N_7521);
nor U7714 (N_7714,N_7573,N_7584);
or U7715 (N_7715,N_7502,N_7498);
and U7716 (N_7716,N_7568,N_7517);
and U7717 (N_7717,N_7467,N_7540);
and U7718 (N_7718,N_7519,N_7497);
nor U7719 (N_7719,N_7593,N_7484);
nor U7720 (N_7720,N_7477,N_7599);
or U7721 (N_7721,N_7579,N_7593);
nand U7722 (N_7722,N_7518,N_7540);
xnor U7723 (N_7723,N_7522,N_7552);
and U7724 (N_7724,N_7585,N_7546);
nor U7725 (N_7725,N_7442,N_7467);
xor U7726 (N_7726,N_7560,N_7578);
or U7727 (N_7727,N_7538,N_7478);
and U7728 (N_7728,N_7411,N_7472);
and U7729 (N_7729,N_7460,N_7472);
xnor U7730 (N_7730,N_7461,N_7573);
or U7731 (N_7731,N_7462,N_7470);
nand U7732 (N_7732,N_7431,N_7561);
xnor U7733 (N_7733,N_7511,N_7556);
nand U7734 (N_7734,N_7494,N_7425);
nand U7735 (N_7735,N_7553,N_7569);
nand U7736 (N_7736,N_7421,N_7530);
or U7737 (N_7737,N_7582,N_7498);
and U7738 (N_7738,N_7496,N_7598);
and U7739 (N_7739,N_7559,N_7420);
xor U7740 (N_7740,N_7542,N_7498);
or U7741 (N_7741,N_7410,N_7435);
and U7742 (N_7742,N_7483,N_7493);
xnor U7743 (N_7743,N_7436,N_7550);
and U7744 (N_7744,N_7400,N_7552);
nand U7745 (N_7745,N_7405,N_7425);
or U7746 (N_7746,N_7508,N_7553);
nor U7747 (N_7747,N_7588,N_7461);
nand U7748 (N_7748,N_7435,N_7428);
nor U7749 (N_7749,N_7537,N_7478);
and U7750 (N_7750,N_7414,N_7505);
nand U7751 (N_7751,N_7538,N_7510);
nand U7752 (N_7752,N_7578,N_7511);
nand U7753 (N_7753,N_7575,N_7489);
xor U7754 (N_7754,N_7553,N_7404);
or U7755 (N_7755,N_7565,N_7450);
and U7756 (N_7756,N_7598,N_7410);
xor U7757 (N_7757,N_7412,N_7555);
nor U7758 (N_7758,N_7474,N_7466);
nor U7759 (N_7759,N_7440,N_7430);
nor U7760 (N_7760,N_7531,N_7440);
xor U7761 (N_7761,N_7427,N_7561);
nor U7762 (N_7762,N_7533,N_7425);
or U7763 (N_7763,N_7573,N_7583);
xnor U7764 (N_7764,N_7563,N_7570);
xor U7765 (N_7765,N_7427,N_7469);
nor U7766 (N_7766,N_7460,N_7593);
xnor U7767 (N_7767,N_7431,N_7539);
xnor U7768 (N_7768,N_7581,N_7588);
and U7769 (N_7769,N_7465,N_7510);
xnor U7770 (N_7770,N_7559,N_7577);
and U7771 (N_7771,N_7536,N_7537);
and U7772 (N_7772,N_7439,N_7456);
and U7773 (N_7773,N_7554,N_7516);
nor U7774 (N_7774,N_7527,N_7404);
nor U7775 (N_7775,N_7428,N_7537);
xor U7776 (N_7776,N_7405,N_7521);
nor U7777 (N_7777,N_7460,N_7500);
or U7778 (N_7778,N_7544,N_7448);
nand U7779 (N_7779,N_7534,N_7546);
xor U7780 (N_7780,N_7414,N_7493);
and U7781 (N_7781,N_7465,N_7488);
or U7782 (N_7782,N_7458,N_7592);
nand U7783 (N_7783,N_7426,N_7590);
nor U7784 (N_7784,N_7489,N_7526);
nor U7785 (N_7785,N_7567,N_7598);
and U7786 (N_7786,N_7419,N_7526);
nand U7787 (N_7787,N_7496,N_7590);
or U7788 (N_7788,N_7492,N_7437);
nand U7789 (N_7789,N_7581,N_7493);
or U7790 (N_7790,N_7504,N_7505);
nand U7791 (N_7791,N_7537,N_7517);
or U7792 (N_7792,N_7497,N_7501);
nor U7793 (N_7793,N_7430,N_7588);
xnor U7794 (N_7794,N_7462,N_7504);
nand U7795 (N_7795,N_7596,N_7404);
nand U7796 (N_7796,N_7513,N_7464);
nor U7797 (N_7797,N_7476,N_7535);
or U7798 (N_7798,N_7468,N_7477);
or U7799 (N_7799,N_7589,N_7497);
or U7800 (N_7800,N_7770,N_7735);
xor U7801 (N_7801,N_7796,N_7733);
xor U7802 (N_7802,N_7777,N_7739);
nand U7803 (N_7803,N_7757,N_7698);
nor U7804 (N_7804,N_7600,N_7743);
xnor U7805 (N_7805,N_7761,N_7660);
and U7806 (N_7806,N_7786,N_7721);
nor U7807 (N_7807,N_7621,N_7691);
nor U7808 (N_7808,N_7727,N_7681);
nor U7809 (N_7809,N_7657,N_7700);
nor U7810 (N_7810,N_7708,N_7793);
nor U7811 (N_7811,N_7688,N_7641);
and U7812 (N_7812,N_7630,N_7784);
and U7813 (N_7813,N_7622,N_7629);
nor U7814 (N_7814,N_7765,N_7731);
xor U7815 (N_7815,N_7722,N_7680);
and U7816 (N_7816,N_7764,N_7677);
and U7817 (N_7817,N_7747,N_7633);
and U7818 (N_7818,N_7610,N_7651);
or U7819 (N_7819,N_7679,N_7746);
nand U7820 (N_7820,N_7696,N_7602);
nand U7821 (N_7821,N_7617,N_7725);
and U7822 (N_7822,N_7741,N_7795);
nor U7823 (N_7823,N_7692,N_7636);
or U7824 (N_7824,N_7618,N_7789);
nor U7825 (N_7825,N_7780,N_7711);
and U7826 (N_7826,N_7763,N_7626);
or U7827 (N_7827,N_7643,N_7737);
or U7828 (N_7828,N_7669,N_7703);
nor U7829 (N_7829,N_7767,N_7707);
nor U7830 (N_7830,N_7753,N_7655);
or U7831 (N_7831,N_7799,N_7683);
nor U7832 (N_7832,N_7730,N_7705);
and U7833 (N_7833,N_7638,N_7775);
nor U7834 (N_7834,N_7615,N_7687);
xnor U7835 (N_7835,N_7738,N_7785);
nand U7836 (N_7836,N_7613,N_7774);
and U7837 (N_7837,N_7783,N_7717);
nand U7838 (N_7838,N_7697,N_7652);
xnor U7839 (N_7839,N_7625,N_7695);
xnor U7840 (N_7840,N_7750,N_7666);
xnor U7841 (N_7841,N_7720,N_7798);
nor U7842 (N_7842,N_7653,N_7693);
and U7843 (N_7843,N_7716,N_7748);
or U7844 (N_7844,N_7769,N_7637);
nor U7845 (N_7845,N_7674,N_7682);
nor U7846 (N_7846,N_7791,N_7606);
xnor U7847 (N_7847,N_7734,N_7604);
nand U7848 (N_7848,N_7646,N_7756);
or U7849 (N_7849,N_7685,N_7623);
or U7850 (N_7850,N_7671,N_7605);
nor U7851 (N_7851,N_7779,N_7794);
xor U7852 (N_7852,N_7797,N_7612);
nor U7853 (N_7853,N_7678,N_7632);
nand U7854 (N_7854,N_7776,N_7663);
xnor U7855 (N_7855,N_7662,N_7740);
xor U7856 (N_7856,N_7792,N_7694);
and U7857 (N_7857,N_7667,N_7689);
and U7858 (N_7858,N_7782,N_7611);
nand U7859 (N_7859,N_7758,N_7631);
or U7860 (N_7860,N_7749,N_7790);
nand U7861 (N_7861,N_7642,N_7648);
or U7862 (N_7862,N_7699,N_7650);
nor U7863 (N_7863,N_7787,N_7773);
xor U7864 (N_7864,N_7712,N_7742);
nor U7865 (N_7865,N_7713,N_7755);
xnor U7866 (N_7866,N_7736,N_7772);
nand U7867 (N_7867,N_7701,N_7619);
nand U7868 (N_7868,N_7668,N_7603);
or U7869 (N_7869,N_7627,N_7628);
xnor U7870 (N_7870,N_7714,N_7673);
nand U7871 (N_7871,N_7640,N_7744);
nand U7872 (N_7872,N_7715,N_7635);
nor U7873 (N_7873,N_7620,N_7684);
xor U7874 (N_7874,N_7768,N_7760);
nand U7875 (N_7875,N_7665,N_7762);
nor U7876 (N_7876,N_7658,N_7732);
nor U7877 (N_7877,N_7690,N_7607);
xnor U7878 (N_7878,N_7726,N_7723);
nor U7879 (N_7879,N_7754,N_7676);
and U7880 (N_7880,N_7778,N_7672);
nand U7881 (N_7881,N_7664,N_7766);
nor U7882 (N_7882,N_7656,N_7675);
nor U7883 (N_7883,N_7649,N_7670);
xnor U7884 (N_7884,N_7609,N_7718);
nor U7885 (N_7885,N_7644,N_7704);
nand U7886 (N_7886,N_7745,N_7654);
nor U7887 (N_7887,N_7647,N_7724);
nand U7888 (N_7888,N_7781,N_7706);
and U7889 (N_7889,N_7624,N_7709);
xor U7890 (N_7890,N_7751,N_7729);
or U7891 (N_7891,N_7661,N_7659);
or U7892 (N_7892,N_7759,N_7601);
and U7893 (N_7893,N_7634,N_7608);
nand U7894 (N_7894,N_7645,N_7616);
nor U7895 (N_7895,N_7752,N_7614);
nand U7896 (N_7896,N_7719,N_7702);
nand U7897 (N_7897,N_7728,N_7639);
nand U7898 (N_7898,N_7710,N_7788);
nor U7899 (N_7899,N_7686,N_7771);
nor U7900 (N_7900,N_7680,N_7693);
xnor U7901 (N_7901,N_7767,N_7713);
nor U7902 (N_7902,N_7735,N_7674);
nor U7903 (N_7903,N_7617,N_7630);
or U7904 (N_7904,N_7648,N_7729);
or U7905 (N_7905,N_7693,N_7736);
or U7906 (N_7906,N_7745,N_7671);
or U7907 (N_7907,N_7691,N_7756);
nor U7908 (N_7908,N_7610,N_7797);
or U7909 (N_7909,N_7719,N_7671);
nor U7910 (N_7910,N_7653,N_7636);
nand U7911 (N_7911,N_7735,N_7631);
nor U7912 (N_7912,N_7727,N_7751);
xor U7913 (N_7913,N_7669,N_7688);
nor U7914 (N_7914,N_7614,N_7611);
nand U7915 (N_7915,N_7750,N_7602);
or U7916 (N_7916,N_7693,N_7754);
nand U7917 (N_7917,N_7720,N_7754);
or U7918 (N_7918,N_7766,N_7637);
xor U7919 (N_7919,N_7705,N_7618);
and U7920 (N_7920,N_7706,N_7711);
nand U7921 (N_7921,N_7714,N_7623);
or U7922 (N_7922,N_7712,N_7676);
nor U7923 (N_7923,N_7746,N_7711);
and U7924 (N_7924,N_7708,N_7728);
nand U7925 (N_7925,N_7712,N_7620);
or U7926 (N_7926,N_7737,N_7766);
or U7927 (N_7927,N_7638,N_7781);
nor U7928 (N_7928,N_7678,N_7643);
or U7929 (N_7929,N_7684,N_7672);
or U7930 (N_7930,N_7774,N_7709);
and U7931 (N_7931,N_7697,N_7789);
nor U7932 (N_7932,N_7774,N_7766);
or U7933 (N_7933,N_7666,N_7780);
xor U7934 (N_7934,N_7680,N_7629);
nand U7935 (N_7935,N_7715,N_7634);
or U7936 (N_7936,N_7769,N_7773);
nor U7937 (N_7937,N_7784,N_7655);
and U7938 (N_7938,N_7665,N_7793);
and U7939 (N_7939,N_7756,N_7798);
nand U7940 (N_7940,N_7651,N_7630);
xnor U7941 (N_7941,N_7607,N_7723);
xor U7942 (N_7942,N_7791,N_7727);
nor U7943 (N_7943,N_7783,N_7609);
nor U7944 (N_7944,N_7785,N_7703);
or U7945 (N_7945,N_7660,N_7755);
or U7946 (N_7946,N_7711,N_7600);
nand U7947 (N_7947,N_7749,N_7799);
xnor U7948 (N_7948,N_7739,N_7700);
nand U7949 (N_7949,N_7624,N_7644);
xnor U7950 (N_7950,N_7753,N_7780);
and U7951 (N_7951,N_7735,N_7737);
or U7952 (N_7952,N_7729,N_7722);
nand U7953 (N_7953,N_7615,N_7742);
and U7954 (N_7954,N_7690,N_7681);
nand U7955 (N_7955,N_7725,N_7729);
nand U7956 (N_7956,N_7703,N_7727);
xor U7957 (N_7957,N_7729,N_7650);
nand U7958 (N_7958,N_7647,N_7671);
or U7959 (N_7959,N_7697,N_7733);
nand U7960 (N_7960,N_7609,N_7689);
and U7961 (N_7961,N_7690,N_7746);
or U7962 (N_7962,N_7753,N_7763);
nand U7963 (N_7963,N_7688,N_7779);
and U7964 (N_7964,N_7665,N_7681);
nand U7965 (N_7965,N_7621,N_7762);
and U7966 (N_7966,N_7769,N_7753);
and U7967 (N_7967,N_7662,N_7744);
or U7968 (N_7968,N_7655,N_7750);
nand U7969 (N_7969,N_7690,N_7728);
nand U7970 (N_7970,N_7677,N_7614);
xnor U7971 (N_7971,N_7611,N_7663);
or U7972 (N_7972,N_7795,N_7715);
and U7973 (N_7973,N_7744,N_7734);
nor U7974 (N_7974,N_7765,N_7727);
nor U7975 (N_7975,N_7680,N_7661);
xnor U7976 (N_7976,N_7745,N_7633);
or U7977 (N_7977,N_7715,N_7710);
xnor U7978 (N_7978,N_7632,N_7789);
or U7979 (N_7979,N_7707,N_7746);
nor U7980 (N_7980,N_7601,N_7697);
nor U7981 (N_7981,N_7658,N_7679);
nand U7982 (N_7982,N_7724,N_7613);
or U7983 (N_7983,N_7782,N_7770);
and U7984 (N_7984,N_7792,N_7671);
or U7985 (N_7985,N_7745,N_7701);
xnor U7986 (N_7986,N_7717,N_7643);
xnor U7987 (N_7987,N_7734,N_7736);
and U7988 (N_7988,N_7628,N_7797);
and U7989 (N_7989,N_7711,N_7721);
and U7990 (N_7990,N_7795,N_7725);
or U7991 (N_7991,N_7787,N_7680);
nor U7992 (N_7992,N_7782,N_7601);
nor U7993 (N_7993,N_7698,N_7668);
or U7994 (N_7994,N_7612,N_7600);
and U7995 (N_7995,N_7616,N_7769);
nand U7996 (N_7996,N_7706,N_7652);
nand U7997 (N_7997,N_7726,N_7686);
nor U7998 (N_7998,N_7762,N_7792);
and U7999 (N_7999,N_7759,N_7793);
and U8000 (N_8000,N_7861,N_7986);
or U8001 (N_8001,N_7977,N_7930);
xnor U8002 (N_8002,N_7950,N_7820);
nor U8003 (N_8003,N_7876,N_7852);
nand U8004 (N_8004,N_7998,N_7914);
nand U8005 (N_8005,N_7855,N_7902);
nand U8006 (N_8006,N_7974,N_7955);
and U8007 (N_8007,N_7886,N_7934);
or U8008 (N_8008,N_7993,N_7845);
or U8009 (N_8009,N_7846,N_7867);
xnor U8010 (N_8010,N_7979,N_7994);
or U8011 (N_8011,N_7967,N_7834);
nand U8012 (N_8012,N_7887,N_7853);
xor U8013 (N_8013,N_7984,N_7952);
nand U8014 (N_8014,N_7889,N_7919);
nand U8015 (N_8015,N_7938,N_7809);
and U8016 (N_8016,N_7838,N_7802);
nor U8017 (N_8017,N_7931,N_7971);
nor U8018 (N_8018,N_7976,N_7854);
nand U8019 (N_8019,N_7828,N_7926);
xnor U8020 (N_8020,N_7922,N_7826);
or U8021 (N_8021,N_7897,N_7801);
nand U8022 (N_8022,N_7923,N_7987);
nor U8023 (N_8023,N_7999,N_7823);
xor U8024 (N_8024,N_7858,N_7936);
xnor U8025 (N_8025,N_7829,N_7992);
and U8026 (N_8026,N_7944,N_7909);
nor U8027 (N_8027,N_7959,N_7811);
and U8028 (N_8028,N_7819,N_7804);
or U8029 (N_8029,N_7905,N_7866);
and U8030 (N_8030,N_7816,N_7806);
nor U8031 (N_8031,N_7877,N_7917);
or U8032 (N_8032,N_7895,N_7882);
xnor U8033 (N_8033,N_7808,N_7817);
xor U8034 (N_8034,N_7906,N_7958);
and U8035 (N_8035,N_7836,N_7839);
xnor U8036 (N_8036,N_7964,N_7894);
and U8037 (N_8037,N_7995,N_7966);
xnor U8038 (N_8038,N_7973,N_7830);
nor U8039 (N_8039,N_7937,N_7844);
xor U8040 (N_8040,N_7827,N_7989);
xor U8041 (N_8041,N_7975,N_7935);
or U8042 (N_8042,N_7961,N_7982);
nand U8043 (N_8043,N_7963,N_7900);
or U8044 (N_8044,N_7913,N_7821);
or U8045 (N_8045,N_7831,N_7932);
and U8046 (N_8046,N_7899,N_7878);
xnor U8047 (N_8047,N_7869,N_7837);
xnor U8048 (N_8048,N_7871,N_7945);
or U8049 (N_8049,N_7972,N_7880);
or U8050 (N_8050,N_7862,N_7856);
and U8051 (N_8051,N_7810,N_7888);
and U8052 (N_8052,N_7920,N_7847);
nand U8053 (N_8053,N_7841,N_7951);
nand U8054 (N_8054,N_7835,N_7870);
nand U8055 (N_8055,N_7881,N_7850);
nor U8056 (N_8056,N_7925,N_7884);
or U8057 (N_8057,N_7947,N_7983);
nor U8058 (N_8058,N_7814,N_7904);
xnor U8059 (N_8059,N_7903,N_7941);
or U8060 (N_8060,N_7822,N_7863);
and U8061 (N_8061,N_7840,N_7928);
nand U8062 (N_8062,N_7891,N_7875);
nor U8063 (N_8063,N_7918,N_7832);
xor U8064 (N_8064,N_7848,N_7843);
nand U8065 (N_8065,N_7818,N_7980);
nor U8066 (N_8066,N_7825,N_7910);
xor U8067 (N_8067,N_7912,N_7851);
nor U8068 (N_8068,N_7857,N_7864);
nand U8069 (N_8069,N_7872,N_7898);
nand U8070 (N_8070,N_7970,N_7924);
or U8071 (N_8071,N_7949,N_7842);
nor U8072 (N_8072,N_7978,N_7883);
nand U8073 (N_8073,N_7940,N_7956);
and U8074 (N_8074,N_7962,N_7991);
or U8075 (N_8075,N_7915,N_7907);
or U8076 (N_8076,N_7824,N_7860);
and U8077 (N_8077,N_7892,N_7946);
xnor U8078 (N_8078,N_7859,N_7868);
or U8079 (N_8079,N_7813,N_7803);
nand U8080 (N_8080,N_7873,N_7960);
or U8081 (N_8081,N_7890,N_7943);
nand U8082 (N_8082,N_7957,N_7988);
nor U8083 (N_8083,N_7885,N_7865);
nor U8084 (N_8084,N_7965,N_7879);
or U8085 (N_8085,N_7893,N_7927);
or U8086 (N_8086,N_7985,N_7815);
xor U8087 (N_8087,N_7996,N_7911);
and U8088 (N_8088,N_7916,N_7805);
nand U8089 (N_8089,N_7933,N_7921);
or U8090 (N_8090,N_7908,N_7901);
xnor U8091 (N_8091,N_7812,N_7849);
and U8092 (N_8092,N_7896,N_7874);
nand U8093 (N_8093,N_7942,N_7968);
nand U8094 (N_8094,N_7948,N_7953);
xor U8095 (N_8095,N_7997,N_7800);
nand U8096 (N_8096,N_7833,N_7981);
and U8097 (N_8097,N_7969,N_7939);
nand U8098 (N_8098,N_7929,N_7807);
xnor U8099 (N_8099,N_7954,N_7990);
nand U8100 (N_8100,N_7977,N_7868);
and U8101 (N_8101,N_7839,N_7893);
nor U8102 (N_8102,N_7844,N_7864);
or U8103 (N_8103,N_7923,N_7964);
and U8104 (N_8104,N_7882,N_7854);
and U8105 (N_8105,N_7883,N_7849);
xor U8106 (N_8106,N_7982,N_7904);
or U8107 (N_8107,N_7959,N_7831);
nor U8108 (N_8108,N_7930,N_7827);
and U8109 (N_8109,N_7927,N_7979);
or U8110 (N_8110,N_7800,N_7933);
and U8111 (N_8111,N_7848,N_7886);
and U8112 (N_8112,N_7849,N_7944);
xnor U8113 (N_8113,N_7907,N_7952);
and U8114 (N_8114,N_7931,N_7983);
xnor U8115 (N_8115,N_7891,N_7851);
and U8116 (N_8116,N_7862,N_7819);
nand U8117 (N_8117,N_7940,N_7997);
xnor U8118 (N_8118,N_7973,N_7801);
xor U8119 (N_8119,N_7958,N_7820);
and U8120 (N_8120,N_7999,N_7882);
and U8121 (N_8121,N_7933,N_7948);
nor U8122 (N_8122,N_7913,N_7804);
and U8123 (N_8123,N_7861,N_7819);
or U8124 (N_8124,N_7884,N_7995);
nor U8125 (N_8125,N_7804,N_7906);
or U8126 (N_8126,N_7821,N_7993);
nor U8127 (N_8127,N_7916,N_7951);
or U8128 (N_8128,N_7832,N_7906);
xnor U8129 (N_8129,N_7867,N_7984);
xnor U8130 (N_8130,N_7828,N_7842);
xor U8131 (N_8131,N_7906,N_7922);
nand U8132 (N_8132,N_7860,N_7828);
nor U8133 (N_8133,N_7880,N_7935);
nand U8134 (N_8134,N_7849,N_7861);
nand U8135 (N_8135,N_7923,N_7839);
xor U8136 (N_8136,N_7813,N_7972);
nor U8137 (N_8137,N_7866,N_7830);
or U8138 (N_8138,N_7891,N_7976);
nor U8139 (N_8139,N_7906,N_7893);
and U8140 (N_8140,N_7924,N_7815);
and U8141 (N_8141,N_7863,N_7935);
and U8142 (N_8142,N_7965,N_7999);
nand U8143 (N_8143,N_7843,N_7968);
or U8144 (N_8144,N_7904,N_7945);
nor U8145 (N_8145,N_7914,N_7858);
or U8146 (N_8146,N_7954,N_7817);
and U8147 (N_8147,N_7817,N_7837);
and U8148 (N_8148,N_7875,N_7896);
nor U8149 (N_8149,N_7966,N_7844);
nor U8150 (N_8150,N_7956,N_7890);
or U8151 (N_8151,N_7966,N_7814);
and U8152 (N_8152,N_7834,N_7825);
xor U8153 (N_8153,N_7873,N_7955);
xor U8154 (N_8154,N_7812,N_7986);
or U8155 (N_8155,N_7924,N_7910);
xnor U8156 (N_8156,N_7851,N_7977);
or U8157 (N_8157,N_7909,N_7953);
nand U8158 (N_8158,N_7951,N_7917);
and U8159 (N_8159,N_7922,N_7851);
nor U8160 (N_8160,N_7978,N_7933);
and U8161 (N_8161,N_7989,N_7846);
and U8162 (N_8162,N_7946,N_7871);
xnor U8163 (N_8163,N_7947,N_7951);
and U8164 (N_8164,N_7900,N_7882);
and U8165 (N_8165,N_7978,N_7998);
nor U8166 (N_8166,N_7895,N_7952);
nand U8167 (N_8167,N_7824,N_7939);
nor U8168 (N_8168,N_7905,N_7924);
nor U8169 (N_8169,N_7937,N_7982);
nand U8170 (N_8170,N_7881,N_7832);
nand U8171 (N_8171,N_7991,N_7820);
xnor U8172 (N_8172,N_7922,N_7893);
nand U8173 (N_8173,N_7877,N_7847);
or U8174 (N_8174,N_7998,N_7968);
xor U8175 (N_8175,N_7978,N_7820);
and U8176 (N_8176,N_7869,N_7814);
and U8177 (N_8177,N_7822,N_7950);
nand U8178 (N_8178,N_7822,N_7907);
nor U8179 (N_8179,N_7883,N_7965);
nor U8180 (N_8180,N_7927,N_7999);
xnor U8181 (N_8181,N_7930,N_7869);
nor U8182 (N_8182,N_7995,N_7975);
xnor U8183 (N_8183,N_7862,N_7918);
nand U8184 (N_8184,N_7842,N_7973);
nand U8185 (N_8185,N_7933,N_7980);
and U8186 (N_8186,N_7830,N_7923);
and U8187 (N_8187,N_7876,N_7802);
xnor U8188 (N_8188,N_7822,N_7946);
xnor U8189 (N_8189,N_7837,N_7936);
or U8190 (N_8190,N_7899,N_7853);
xor U8191 (N_8191,N_7902,N_7814);
nor U8192 (N_8192,N_7974,N_7908);
nor U8193 (N_8193,N_7830,N_7929);
nand U8194 (N_8194,N_7943,N_7928);
nor U8195 (N_8195,N_7991,N_7903);
xor U8196 (N_8196,N_7942,N_7865);
or U8197 (N_8197,N_7852,N_7881);
nand U8198 (N_8198,N_7901,N_7950);
nor U8199 (N_8199,N_7999,N_7957);
nand U8200 (N_8200,N_8180,N_8059);
nor U8201 (N_8201,N_8172,N_8191);
or U8202 (N_8202,N_8087,N_8041);
nand U8203 (N_8203,N_8186,N_8104);
and U8204 (N_8204,N_8011,N_8159);
nand U8205 (N_8205,N_8102,N_8066);
and U8206 (N_8206,N_8182,N_8069);
xnor U8207 (N_8207,N_8044,N_8030);
xor U8208 (N_8208,N_8153,N_8058);
or U8209 (N_8209,N_8150,N_8198);
xnor U8210 (N_8210,N_8063,N_8000);
or U8211 (N_8211,N_8192,N_8114);
xnor U8212 (N_8212,N_8196,N_8080);
xnor U8213 (N_8213,N_8048,N_8073);
nor U8214 (N_8214,N_8161,N_8072);
nor U8215 (N_8215,N_8188,N_8143);
xor U8216 (N_8216,N_8169,N_8012);
nand U8217 (N_8217,N_8117,N_8195);
or U8218 (N_8218,N_8155,N_8070);
xnor U8219 (N_8219,N_8189,N_8013);
nor U8220 (N_8220,N_8103,N_8166);
nor U8221 (N_8221,N_8164,N_8081);
nand U8222 (N_8222,N_8163,N_8038);
xnor U8223 (N_8223,N_8099,N_8168);
or U8224 (N_8224,N_8165,N_8098);
and U8225 (N_8225,N_8127,N_8090);
nand U8226 (N_8226,N_8075,N_8110);
and U8227 (N_8227,N_8015,N_8078);
nor U8228 (N_8228,N_8181,N_8167);
nor U8229 (N_8229,N_8129,N_8184);
nor U8230 (N_8230,N_8065,N_8079);
and U8231 (N_8231,N_8137,N_8146);
xor U8232 (N_8232,N_8086,N_8040);
nor U8233 (N_8233,N_8135,N_8126);
or U8234 (N_8234,N_8130,N_8091);
or U8235 (N_8235,N_8197,N_8083);
nor U8236 (N_8236,N_8039,N_8108);
and U8237 (N_8237,N_8116,N_8154);
and U8238 (N_8238,N_8122,N_8057);
nor U8239 (N_8239,N_8009,N_8095);
or U8240 (N_8240,N_8061,N_8007);
nor U8241 (N_8241,N_8094,N_8032);
nor U8242 (N_8242,N_8004,N_8084);
or U8243 (N_8243,N_8112,N_8025);
or U8244 (N_8244,N_8023,N_8014);
nand U8245 (N_8245,N_8077,N_8019);
or U8246 (N_8246,N_8131,N_8034);
or U8247 (N_8247,N_8177,N_8021);
nor U8248 (N_8248,N_8067,N_8017);
or U8249 (N_8249,N_8047,N_8042);
xnor U8250 (N_8250,N_8051,N_8187);
and U8251 (N_8251,N_8139,N_8120);
or U8252 (N_8252,N_8178,N_8128);
xnor U8253 (N_8253,N_8055,N_8107);
or U8254 (N_8254,N_8016,N_8101);
or U8255 (N_8255,N_8097,N_8046);
nand U8256 (N_8256,N_8148,N_8050);
nand U8257 (N_8257,N_8142,N_8033);
and U8258 (N_8258,N_8076,N_8132);
xor U8259 (N_8259,N_8074,N_8071);
nor U8260 (N_8260,N_8190,N_8149);
or U8261 (N_8261,N_8096,N_8160);
or U8262 (N_8262,N_8060,N_8052);
nand U8263 (N_8263,N_8141,N_8156);
xnor U8264 (N_8264,N_8006,N_8037);
nor U8265 (N_8265,N_8053,N_8133);
nand U8266 (N_8266,N_8176,N_8173);
nand U8267 (N_8267,N_8010,N_8170);
nand U8268 (N_8268,N_8064,N_8115);
nor U8269 (N_8269,N_8134,N_8027);
nor U8270 (N_8270,N_8147,N_8024);
and U8271 (N_8271,N_8183,N_8068);
and U8272 (N_8272,N_8003,N_8054);
xnor U8273 (N_8273,N_8100,N_8031);
nor U8274 (N_8274,N_8158,N_8082);
xor U8275 (N_8275,N_8056,N_8029);
xor U8276 (N_8276,N_8136,N_8185);
nor U8277 (N_8277,N_8175,N_8018);
or U8278 (N_8278,N_8085,N_8151);
xor U8279 (N_8279,N_8092,N_8026);
or U8280 (N_8280,N_8119,N_8105);
and U8281 (N_8281,N_8035,N_8028);
and U8282 (N_8282,N_8089,N_8113);
or U8283 (N_8283,N_8045,N_8174);
nor U8284 (N_8284,N_8043,N_8106);
or U8285 (N_8285,N_8020,N_8194);
or U8286 (N_8286,N_8118,N_8124);
or U8287 (N_8287,N_8062,N_8123);
xnor U8288 (N_8288,N_8121,N_8162);
or U8289 (N_8289,N_8140,N_8093);
nor U8290 (N_8290,N_8049,N_8152);
xor U8291 (N_8291,N_8088,N_8109);
xnor U8292 (N_8292,N_8022,N_8036);
nand U8293 (N_8293,N_8199,N_8145);
and U8294 (N_8294,N_8171,N_8193);
and U8295 (N_8295,N_8111,N_8157);
and U8296 (N_8296,N_8008,N_8005);
or U8297 (N_8297,N_8001,N_8138);
xnor U8298 (N_8298,N_8179,N_8125);
nor U8299 (N_8299,N_8002,N_8144);
and U8300 (N_8300,N_8062,N_8095);
xnor U8301 (N_8301,N_8173,N_8000);
or U8302 (N_8302,N_8075,N_8156);
or U8303 (N_8303,N_8153,N_8007);
xor U8304 (N_8304,N_8121,N_8172);
and U8305 (N_8305,N_8153,N_8017);
or U8306 (N_8306,N_8075,N_8024);
xnor U8307 (N_8307,N_8147,N_8123);
or U8308 (N_8308,N_8137,N_8145);
and U8309 (N_8309,N_8096,N_8168);
and U8310 (N_8310,N_8119,N_8084);
and U8311 (N_8311,N_8190,N_8046);
nand U8312 (N_8312,N_8132,N_8144);
nor U8313 (N_8313,N_8097,N_8182);
or U8314 (N_8314,N_8118,N_8099);
nand U8315 (N_8315,N_8001,N_8133);
nand U8316 (N_8316,N_8056,N_8162);
nor U8317 (N_8317,N_8082,N_8165);
nor U8318 (N_8318,N_8074,N_8016);
and U8319 (N_8319,N_8155,N_8162);
or U8320 (N_8320,N_8041,N_8008);
or U8321 (N_8321,N_8109,N_8122);
or U8322 (N_8322,N_8188,N_8023);
or U8323 (N_8323,N_8010,N_8118);
nor U8324 (N_8324,N_8066,N_8010);
nand U8325 (N_8325,N_8181,N_8099);
or U8326 (N_8326,N_8030,N_8090);
xor U8327 (N_8327,N_8145,N_8167);
nand U8328 (N_8328,N_8128,N_8175);
xor U8329 (N_8329,N_8137,N_8026);
nand U8330 (N_8330,N_8179,N_8150);
or U8331 (N_8331,N_8058,N_8079);
or U8332 (N_8332,N_8132,N_8016);
and U8333 (N_8333,N_8124,N_8175);
and U8334 (N_8334,N_8064,N_8049);
and U8335 (N_8335,N_8043,N_8014);
or U8336 (N_8336,N_8134,N_8054);
nand U8337 (N_8337,N_8161,N_8130);
and U8338 (N_8338,N_8107,N_8000);
nor U8339 (N_8339,N_8019,N_8054);
or U8340 (N_8340,N_8115,N_8173);
nand U8341 (N_8341,N_8042,N_8040);
nand U8342 (N_8342,N_8008,N_8035);
nand U8343 (N_8343,N_8060,N_8097);
and U8344 (N_8344,N_8149,N_8158);
and U8345 (N_8345,N_8147,N_8064);
nor U8346 (N_8346,N_8074,N_8061);
nand U8347 (N_8347,N_8112,N_8184);
nor U8348 (N_8348,N_8070,N_8052);
and U8349 (N_8349,N_8129,N_8105);
nand U8350 (N_8350,N_8098,N_8111);
and U8351 (N_8351,N_8005,N_8133);
or U8352 (N_8352,N_8066,N_8051);
or U8353 (N_8353,N_8141,N_8188);
nor U8354 (N_8354,N_8060,N_8001);
nand U8355 (N_8355,N_8093,N_8059);
or U8356 (N_8356,N_8143,N_8083);
or U8357 (N_8357,N_8020,N_8088);
or U8358 (N_8358,N_8101,N_8173);
nor U8359 (N_8359,N_8121,N_8065);
xnor U8360 (N_8360,N_8029,N_8045);
nand U8361 (N_8361,N_8103,N_8018);
xnor U8362 (N_8362,N_8014,N_8004);
nand U8363 (N_8363,N_8011,N_8051);
and U8364 (N_8364,N_8084,N_8153);
xnor U8365 (N_8365,N_8175,N_8103);
or U8366 (N_8366,N_8055,N_8182);
xnor U8367 (N_8367,N_8101,N_8009);
or U8368 (N_8368,N_8166,N_8145);
nand U8369 (N_8369,N_8055,N_8089);
or U8370 (N_8370,N_8066,N_8018);
xor U8371 (N_8371,N_8008,N_8056);
and U8372 (N_8372,N_8142,N_8117);
nand U8373 (N_8373,N_8086,N_8064);
or U8374 (N_8374,N_8085,N_8130);
or U8375 (N_8375,N_8033,N_8006);
xor U8376 (N_8376,N_8074,N_8060);
nor U8377 (N_8377,N_8137,N_8110);
or U8378 (N_8378,N_8004,N_8106);
xor U8379 (N_8379,N_8150,N_8025);
or U8380 (N_8380,N_8172,N_8149);
nand U8381 (N_8381,N_8139,N_8069);
or U8382 (N_8382,N_8195,N_8126);
nand U8383 (N_8383,N_8072,N_8068);
nand U8384 (N_8384,N_8071,N_8122);
and U8385 (N_8385,N_8157,N_8103);
xor U8386 (N_8386,N_8081,N_8184);
nand U8387 (N_8387,N_8045,N_8186);
nand U8388 (N_8388,N_8027,N_8111);
nand U8389 (N_8389,N_8010,N_8024);
nor U8390 (N_8390,N_8064,N_8117);
nor U8391 (N_8391,N_8055,N_8049);
nand U8392 (N_8392,N_8023,N_8055);
nor U8393 (N_8393,N_8110,N_8169);
or U8394 (N_8394,N_8176,N_8059);
xnor U8395 (N_8395,N_8103,N_8098);
nand U8396 (N_8396,N_8017,N_8035);
xnor U8397 (N_8397,N_8109,N_8060);
and U8398 (N_8398,N_8045,N_8182);
or U8399 (N_8399,N_8009,N_8012);
and U8400 (N_8400,N_8347,N_8342);
nor U8401 (N_8401,N_8297,N_8338);
nor U8402 (N_8402,N_8291,N_8350);
or U8403 (N_8403,N_8209,N_8200);
nor U8404 (N_8404,N_8252,N_8217);
nor U8405 (N_8405,N_8287,N_8399);
nand U8406 (N_8406,N_8301,N_8335);
and U8407 (N_8407,N_8339,N_8305);
nand U8408 (N_8408,N_8302,N_8355);
nand U8409 (N_8409,N_8284,N_8299);
and U8410 (N_8410,N_8282,N_8325);
xnor U8411 (N_8411,N_8249,N_8344);
or U8412 (N_8412,N_8280,N_8216);
or U8413 (N_8413,N_8296,N_8224);
nand U8414 (N_8414,N_8379,N_8393);
and U8415 (N_8415,N_8259,N_8233);
xor U8416 (N_8416,N_8245,N_8311);
xnor U8417 (N_8417,N_8211,N_8290);
nand U8418 (N_8418,N_8367,N_8227);
xnor U8419 (N_8419,N_8359,N_8271);
nand U8420 (N_8420,N_8303,N_8298);
nor U8421 (N_8421,N_8374,N_8349);
nand U8422 (N_8422,N_8219,N_8329);
xnor U8423 (N_8423,N_8395,N_8276);
nor U8424 (N_8424,N_8244,N_8377);
xor U8425 (N_8425,N_8274,N_8319);
xnor U8426 (N_8426,N_8358,N_8292);
or U8427 (N_8427,N_8340,N_8324);
nand U8428 (N_8428,N_8261,N_8215);
nand U8429 (N_8429,N_8343,N_8201);
and U8430 (N_8430,N_8314,N_8204);
nand U8431 (N_8431,N_8218,N_8354);
xor U8432 (N_8432,N_8214,N_8283);
nand U8433 (N_8433,N_8229,N_8368);
nor U8434 (N_8434,N_8238,N_8304);
or U8435 (N_8435,N_8365,N_8337);
or U8436 (N_8436,N_8231,N_8369);
xor U8437 (N_8437,N_8262,N_8246);
and U8438 (N_8438,N_8373,N_8361);
and U8439 (N_8439,N_8389,N_8388);
or U8440 (N_8440,N_8318,N_8309);
nand U8441 (N_8441,N_8264,N_8221);
nand U8442 (N_8442,N_8327,N_8241);
nor U8443 (N_8443,N_8357,N_8307);
nor U8444 (N_8444,N_8396,N_8253);
nor U8445 (N_8445,N_8308,N_8234);
nor U8446 (N_8446,N_8346,N_8352);
xor U8447 (N_8447,N_8289,N_8254);
xnor U8448 (N_8448,N_8225,N_8364);
nand U8449 (N_8449,N_8232,N_8371);
nor U8450 (N_8450,N_8378,N_8202);
nand U8451 (N_8451,N_8336,N_8334);
or U8452 (N_8452,N_8300,N_8383);
and U8453 (N_8453,N_8391,N_8382);
nand U8454 (N_8454,N_8273,N_8205);
nand U8455 (N_8455,N_8239,N_8392);
nand U8456 (N_8456,N_8356,N_8363);
xor U8457 (N_8457,N_8206,N_8295);
nor U8458 (N_8458,N_8328,N_8330);
nor U8459 (N_8459,N_8323,N_8384);
or U8460 (N_8460,N_8256,N_8317);
and U8461 (N_8461,N_8236,N_8260);
xor U8462 (N_8462,N_8288,N_8351);
xnor U8463 (N_8463,N_8257,N_8203);
nor U8464 (N_8464,N_8248,N_8370);
xor U8465 (N_8465,N_8390,N_8360);
and U8466 (N_8466,N_8397,N_8281);
or U8467 (N_8467,N_8268,N_8230);
or U8468 (N_8468,N_8277,N_8294);
or U8469 (N_8469,N_8394,N_8312);
or U8470 (N_8470,N_8348,N_8385);
or U8471 (N_8471,N_8272,N_8278);
and U8472 (N_8472,N_8228,N_8251);
xnor U8473 (N_8473,N_8285,N_8263);
and U8474 (N_8474,N_8326,N_8353);
nor U8475 (N_8475,N_8279,N_8310);
or U8476 (N_8476,N_8220,N_8398);
xor U8477 (N_8477,N_8275,N_8240);
xor U8478 (N_8478,N_8208,N_8386);
and U8479 (N_8479,N_8250,N_8286);
xnor U8480 (N_8480,N_8242,N_8381);
xor U8481 (N_8481,N_8269,N_8306);
nand U8482 (N_8482,N_8210,N_8266);
and U8483 (N_8483,N_8333,N_8222);
or U8484 (N_8484,N_8212,N_8366);
nand U8485 (N_8485,N_8362,N_8321);
and U8486 (N_8486,N_8213,N_8375);
and U8487 (N_8487,N_8315,N_8207);
nor U8488 (N_8488,N_8247,N_8258);
or U8489 (N_8489,N_8237,N_8332);
nor U8490 (N_8490,N_8322,N_8341);
nand U8491 (N_8491,N_8345,N_8267);
xnor U8492 (N_8492,N_8320,N_8316);
or U8493 (N_8493,N_8255,N_8387);
or U8494 (N_8494,N_8331,N_8293);
or U8495 (N_8495,N_8226,N_8376);
nor U8496 (N_8496,N_8265,N_8223);
xor U8497 (N_8497,N_8380,N_8243);
and U8498 (N_8498,N_8372,N_8313);
and U8499 (N_8499,N_8235,N_8270);
nand U8500 (N_8500,N_8288,N_8216);
xor U8501 (N_8501,N_8204,N_8212);
and U8502 (N_8502,N_8337,N_8222);
and U8503 (N_8503,N_8226,N_8242);
xnor U8504 (N_8504,N_8392,N_8231);
nand U8505 (N_8505,N_8349,N_8220);
or U8506 (N_8506,N_8385,N_8310);
or U8507 (N_8507,N_8295,N_8237);
or U8508 (N_8508,N_8357,N_8258);
nor U8509 (N_8509,N_8232,N_8276);
nor U8510 (N_8510,N_8302,N_8303);
nand U8511 (N_8511,N_8216,N_8309);
nand U8512 (N_8512,N_8200,N_8327);
nor U8513 (N_8513,N_8229,N_8346);
nand U8514 (N_8514,N_8253,N_8268);
or U8515 (N_8515,N_8386,N_8286);
nor U8516 (N_8516,N_8281,N_8394);
nand U8517 (N_8517,N_8391,N_8305);
and U8518 (N_8518,N_8290,N_8353);
or U8519 (N_8519,N_8307,N_8306);
and U8520 (N_8520,N_8206,N_8306);
nand U8521 (N_8521,N_8218,N_8277);
xor U8522 (N_8522,N_8313,N_8337);
nand U8523 (N_8523,N_8373,N_8313);
nand U8524 (N_8524,N_8360,N_8392);
or U8525 (N_8525,N_8360,N_8272);
xnor U8526 (N_8526,N_8353,N_8250);
nand U8527 (N_8527,N_8325,N_8264);
and U8528 (N_8528,N_8265,N_8370);
nand U8529 (N_8529,N_8266,N_8389);
nor U8530 (N_8530,N_8306,N_8389);
nand U8531 (N_8531,N_8226,N_8255);
xor U8532 (N_8532,N_8369,N_8234);
xor U8533 (N_8533,N_8244,N_8296);
xor U8534 (N_8534,N_8235,N_8328);
or U8535 (N_8535,N_8264,N_8289);
nand U8536 (N_8536,N_8304,N_8349);
and U8537 (N_8537,N_8353,N_8214);
xnor U8538 (N_8538,N_8395,N_8391);
and U8539 (N_8539,N_8218,N_8258);
and U8540 (N_8540,N_8382,N_8279);
and U8541 (N_8541,N_8327,N_8274);
or U8542 (N_8542,N_8353,N_8297);
nor U8543 (N_8543,N_8293,N_8205);
or U8544 (N_8544,N_8241,N_8224);
xor U8545 (N_8545,N_8370,N_8243);
or U8546 (N_8546,N_8330,N_8380);
nand U8547 (N_8547,N_8309,N_8334);
nand U8548 (N_8548,N_8257,N_8381);
xnor U8549 (N_8549,N_8266,N_8230);
nand U8550 (N_8550,N_8343,N_8207);
nand U8551 (N_8551,N_8385,N_8205);
and U8552 (N_8552,N_8336,N_8353);
nand U8553 (N_8553,N_8218,N_8208);
or U8554 (N_8554,N_8226,N_8340);
xnor U8555 (N_8555,N_8303,N_8202);
nand U8556 (N_8556,N_8356,N_8324);
nand U8557 (N_8557,N_8343,N_8399);
or U8558 (N_8558,N_8355,N_8223);
and U8559 (N_8559,N_8244,N_8223);
and U8560 (N_8560,N_8301,N_8381);
or U8561 (N_8561,N_8351,N_8274);
nand U8562 (N_8562,N_8283,N_8356);
or U8563 (N_8563,N_8237,N_8213);
and U8564 (N_8564,N_8215,N_8275);
and U8565 (N_8565,N_8284,N_8254);
and U8566 (N_8566,N_8299,N_8282);
nor U8567 (N_8567,N_8294,N_8220);
nand U8568 (N_8568,N_8327,N_8236);
or U8569 (N_8569,N_8316,N_8349);
and U8570 (N_8570,N_8252,N_8215);
nand U8571 (N_8571,N_8376,N_8364);
nor U8572 (N_8572,N_8322,N_8365);
nand U8573 (N_8573,N_8239,N_8216);
xor U8574 (N_8574,N_8314,N_8330);
and U8575 (N_8575,N_8240,N_8218);
nand U8576 (N_8576,N_8346,N_8383);
or U8577 (N_8577,N_8283,N_8202);
and U8578 (N_8578,N_8252,N_8293);
nor U8579 (N_8579,N_8318,N_8396);
and U8580 (N_8580,N_8286,N_8378);
nand U8581 (N_8581,N_8324,N_8248);
or U8582 (N_8582,N_8273,N_8299);
or U8583 (N_8583,N_8243,N_8392);
or U8584 (N_8584,N_8265,N_8396);
nor U8585 (N_8585,N_8223,N_8389);
or U8586 (N_8586,N_8379,N_8363);
nand U8587 (N_8587,N_8317,N_8333);
and U8588 (N_8588,N_8364,N_8371);
nor U8589 (N_8589,N_8288,N_8374);
and U8590 (N_8590,N_8338,N_8268);
and U8591 (N_8591,N_8269,N_8371);
nor U8592 (N_8592,N_8284,N_8275);
nand U8593 (N_8593,N_8313,N_8256);
xor U8594 (N_8594,N_8349,N_8268);
nand U8595 (N_8595,N_8219,N_8382);
and U8596 (N_8596,N_8318,N_8356);
or U8597 (N_8597,N_8206,N_8381);
nor U8598 (N_8598,N_8381,N_8284);
and U8599 (N_8599,N_8349,N_8357);
and U8600 (N_8600,N_8507,N_8560);
nand U8601 (N_8601,N_8553,N_8575);
or U8602 (N_8602,N_8492,N_8580);
xnor U8603 (N_8603,N_8402,N_8434);
nand U8604 (N_8604,N_8417,N_8436);
and U8605 (N_8605,N_8541,N_8564);
nor U8606 (N_8606,N_8487,N_8491);
xnor U8607 (N_8607,N_8499,N_8589);
xor U8608 (N_8608,N_8478,N_8573);
nand U8609 (N_8609,N_8486,N_8442);
or U8610 (N_8610,N_8432,N_8599);
or U8611 (N_8611,N_8456,N_8488);
or U8612 (N_8612,N_8424,N_8479);
and U8613 (N_8613,N_8538,N_8501);
and U8614 (N_8614,N_8406,N_8407);
or U8615 (N_8615,N_8531,N_8472);
and U8616 (N_8616,N_8427,N_8430);
or U8617 (N_8617,N_8482,N_8527);
and U8618 (N_8618,N_8400,N_8506);
xor U8619 (N_8619,N_8416,N_8449);
xor U8620 (N_8620,N_8550,N_8539);
and U8621 (N_8621,N_8429,N_8477);
nor U8622 (N_8622,N_8423,N_8590);
and U8623 (N_8623,N_8425,N_8464);
nand U8624 (N_8624,N_8543,N_8569);
xnor U8625 (N_8625,N_8405,N_8594);
nor U8626 (N_8626,N_8511,N_8544);
xnor U8627 (N_8627,N_8509,N_8411);
nand U8628 (N_8628,N_8444,N_8467);
xor U8629 (N_8629,N_8532,N_8495);
and U8630 (N_8630,N_8552,N_8570);
nand U8631 (N_8631,N_8502,N_8498);
and U8632 (N_8632,N_8483,N_8408);
and U8633 (N_8633,N_8582,N_8579);
xnor U8634 (N_8634,N_8525,N_8412);
nor U8635 (N_8635,N_8508,N_8535);
nor U8636 (N_8636,N_8421,N_8463);
and U8637 (N_8637,N_8583,N_8420);
and U8638 (N_8638,N_8563,N_8572);
and U8639 (N_8639,N_8439,N_8414);
nand U8640 (N_8640,N_8517,N_8476);
and U8641 (N_8641,N_8461,N_8592);
or U8642 (N_8642,N_8497,N_8526);
nor U8643 (N_8643,N_8536,N_8542);
nor U8644 (N_8644,N_8493,N_8428);
and U8645 (N_8645,N_8596,N_8410);
xor U8646 (N_8646,N_8586,N_8403);
or U8647 (N_8647,N_8513,N_8540);
nand U8648 (N_8648,N_8469,N_8473);
nand U8649 (N_8649,N_8504,N_8519);
nor U8650 (N_8650,N_8455,N_8431);
xor U8651 (N_8651,N_8593,N_8555);
or U8652 (N_8652,N_8468,N_8565);
or U8653 (N_8653,N_8462,N_8481);
and U8654 (N_8654,N_8521,N_8452);
nor U8655 (N_8655,N_8466,N_8447);
or U8656 (N_8656,N_8445,N_8401);
nand U8657 (N_8657,N_8598,N_8409);
xor U8658 (N_8658,N_8404,N_8437);
nand U8659 (N_8659,N_8528,N_8558);
nand U8660 (N_8660,N_8556,N_8480);
and U8661 (N_8661,N_8595,N_8557);
nor U8662 (N_8662,N_8474,N_8566);
or U8663 (N_8663,N_8496,N_8574);
nor U8664 (N_8664,N_8505,N_8494);
and U8665 (N_8665,N_8426,N_8551);
or U8666 (N_8666,N_8591,N_8490);
xnor U8667 (N_8667,N_8522,N_8454);
xnor U8668 (N_8668,N_8485,N_8561);
xor U8669 (N_8669,N_8446,N_8547);
nand U8670 (N_8670,N_8448,N_8576);
nor U8671 (N_8671,N_8500,N_8458);
nand U8672 (N_8672,N_8567,N_8484);
nor U8673 (N_8673,N_8453,N_8518);
and U8674 (N_8674,N_8419,N_8571);
nand U8675 (N_8675,N_8415,N_8530);
nor U8676 (N_8676,N_8581,N_8503);
xor U8677 (N_8677,N_8465,N_8435);
xor U8678 (N_8678,N_8457,N_8534);
nor U8679 (N_8679,N_8470,N_8475);
and U8680 (N_8680,N_8545,N_8597);
xor U8681 (N_8681,N_8459,N_8537);
or U8682 (N_8682,N_8584,N_8524);
nor U8683 (N_8683,N_8577,N_8440);
nor U8684 (N_8684,N_8422,N_8529);
or U8685 (N_8685,N_8516,N_8562);
nand U8686 (N_8686,N_8443,N_8441);
nand U8687 (N_8687,N_8533,N_8451);
or U8688 (N_8688,N_8568,N_8587);
xor U8689 (N_8689,N_8588,N_8418);
and U8690 (N_8690,N_8548,N_8559);
nor U8691 (N_8691,N_8512,N_8510);
xnor U8692 (N_8692,N_8450,N_8489);
and U8693 (N_8693,N_8523,N_8471);
nor U8694 (N_8694,N_8413,N_8578);
nor U8695 (N_8695,N_8585,N_8549);
and U8696 (N_8696,N_8438,N_8515);
xor U8697 (N_8697,N_8460,N_8554);
or U8698 (N_8698,N_8546,N_8433);
nand U8699 (N_8699,N_8520,N_8514);
nand U8700 (N_8700,N_8534,N_8586);
nor U8701 (N_8701,N_8489,N_8434);
nand U8702 (N_8702,N_8485,N_8451);
nor U8703 (N_8703,N_8580,N_8556);
or U8704 (N_8704,N_8582,N_8522);
nand U8705 (N_8705,N_8474,N_8598);
nand U8706 (N_8706,N_8419,N_8550);
or U8707 (N_8707,N_8488,N_8541);
nand U8708 (N_8708,N_8560,N_8446);
or U8709 (N_8709,N_8432,N_8535);
or U8710 (N_8710,N_8563,N_8506);
or U8711 (N_8711,N_8558,N_8447);
nor U8712 (N_8712,N_8401,N_8572);
nor U8713 (N_8713,N_8417,N_8504);
nor U8714 (N_8714,N_8563,N_8580);
nor U8715 (N_8715,N_8464,N_8595);
and U8716 (N_8716,N_8496,N_8410);
nand U8717 (N_8717,N_8526,N_8433);
nand U8718 (N_8718,N_8490,N_8563);
and U8719 (N_8719,N_8482,N_8461);
nand U8720 (N_8720,N_8493,N_8575);
nand U8721 (N_8721,N_8439,N_8404);
xnor U8722 (N_8722,N_8563,N_8598);
nand U8723 (N_8723,N_8486,N_8531);
xor U8724 (N_8724,N_8441,N_8415);
xor U8725 (N_8725,N_8421,N_8412);
and U8726 (N_8726,N_8473,N_8435);
xor U8727 (N_8727,N_8466,N_8415);
or U8728 (N_8728,N_8525,N_8404);
nand U8729 (N_8729,N_8408,N_8423);
and U8730 (N_8730,N_8456,N_8401);
xnor U8731 (N_8731,N_8544,N_8482);
and U8732 (N_8732,N_8442,N_8567);
and U8733 (N_8733,N_8464,N_8519);
or U8734 (N_8734,N_8576,N_8442);
and U8735 (N_8735,N_8487,N_8597);
nand U8736 (N_8736,N_8555,N_8482);
and U8737 (N_8737,N_8574,N_8565);
nor U8738 (N_8738,N_8439,N_8499);
nor U8739 (N_8739,N_8465,N_8539);
and U8740 (N_8740,N_8473,N_8521);
nand U8741 (N_8741,N_8482,N_8502);
or U8742 (N_8742,N_8511,N_8479);
nor U8743 (N_8743,N_8513,N_8496);
and U8744 (N_8744,N_8449,N_8456);
and U8745 (N_8745,N_8434,N_8414);
nand U8746 (N_8746,N_8426,N_8419);
and U8747 (N_8747,N_8526,N_8492);
nor U8748 (N_8748,N_8508,N_8487);
and U8749 (N_8749,N_8501,N_8559);
xor U8750 (N_8750,N_8414,N_8419);
or U8751 (N_8751,N_8427,N_8493);
or U8752 (N_8752,N_8428,N_8477);
nor U8753 (N_8753,N_8402,N_8474);
nand U8754 (N_8754,N_8567,N_8454);
nor U8755 (N_8755,N_8542,N_8546);
nand U8756 (N_8756,N_8472,N_8571);
and U8757 (N_8757,N_8561,N_8445);
and U8758 (N_8758,N_8537,N_8469);
nor U8759 (N_8759,N_8505,N_8531);
nand U8760 (N_8760,N_8468,N_8596);
xor U8761 (N_8761,N_8528,N_8431);
nor U8762 (N_8762,N_8567,N_8535);
xor U8763 (N_8763,N_8539,N_8584);
and U8764 (N_8764,N_8510,N_8401);
xnor U8765 (N_8765,N_8429,N_8559);
nand U8766 (N_8766,N_8411,N_8488);
and U8767 (N_8767,N_8450,N_8505);
xor U8768 (N_8768,N_8562,N_8560);
nor U8769 (N_8769,N_8466,N_8459);
and U8770 (N_8770,N_8474,N_8554);
nor U8771 (N_8771,N_8418,N_8486);
nor U8772 (N_8772,N_8526,N_8491);
and U8773 (N_8773,N_8403,N_8481);
or U8774 (N_8774,N_8474,N_8420);
xnor U8775 (N_8775,N_8465,N_8507);
nor U8776 (N_8776,N_8496,N_8419);
xnor U8777 (N_8777,N_8454,N_8459);
xnor U8778 (N_8778,N_8595,N_8547);
nand U8779 (N_8779,N_8414,N_8518);
xor U8780 (N_8780,N_8480,N_8413);
nor U8781 (N_8781,N_8455,N_8476);
or U8782 (N_8782,N_8532,N_8410);
nor U8783 (N_8783,N_8585,N_8532);
xor U8784 (N_8784,N_8455,N_8556);
xor U8785 (N_8785,N_8423,N_8511);
nor U8786 (N_8786,N_8574,N_8576);
xor U8787 (N_8787,N_8489,N_8580);
nand U8788 (N_8788,N_8458,N_8472);
nand U8789 (N_8789,N_8526,N_8586);
nand U8790 (N_8790,N_8433,N_8583);
nor U8791 (N_8791,N_8569,N_8489);
nand U8792 (N_8792,N_8567,N_8436);
nand U8793 (N_8793,N_8520,N_8598);
or U8794 (N_8794,N_8440,N_8424);
or U8795 (N_8795,N_8522,N_8456);
xor U8796 (N_8796,N_8461,N_8469);
nand U8797 (N_8797,N_8413,N_8566);
nand U8798 (N_8798,N_8576,N_8588);
nand U8799 (N_8799,N_8459,N_8489);
or U8800 (N_8800,N_8686,N_8740);
nor U8801 (N_8801,N_8624,N_8693);
nand U8802 (N_8802,N_8703,N_8723);
and U8803 (N_8803,N_8643,N_8657);
nand U8804 (N_8804,N_8653,N_8719);
and U8805 (N_8805,N_8699,N_8648);
or U8806 (N_8806,N_8731,N_8606);
nor U8807 (N_8807,N_8689,N_8766);
nor U8808 (N_8808,N_8661,N_8662);
or U8809 (N_8809,N_8732,N_8612);
nor U8810 (N_8810,N_8652,N_8639);
or U8811 (N_8811,N_8609,N_8674);
nor U8812 (N_8812,N_8678,N_8694);
xor U8813 (N_8813,N_8763,N_8664);
and U8814 (N_8814,N_8622,N_8717);
nand U8815 (N_8815,N_8666,N_8600);
and U8816 (N_8816,N_8796,N_8728);
xnor U8817 (N_8817,N_8746,N_8697);
and U8818 (N_8818,N_8619,N_8747);
or U8819 (N_8819,N_8785,N_8646);
xor U8820 (N_8820,N_8617,N_8607);
xor U8821 (N_8821,N_8601,N_8795);
nand U8822 (N_8822,N_8775,N_8668);
xnor U8823 (N_8823,N_8651,N_8791);
nand U8824 (N_8824,N_8730,N_8629);
or U8825 (N_8825,N_8616,N_8650);
or U8826 (N_8826,N_8673,N_8705);
nand U8827 (N_8827,N_8618,N_8632);
nand U8828 (N_8828,N_8783,N_8748);
nor U8829 (N_8829,N_8675,N_8782);
and U8830 (N_8830,N_8769,N_8644);
or U8831 (N_8831,N_8718,N_8663);
or U8832 (N_8832,N_8608,N_8659);
nor U8833 (N_8833,N_8628,N_8637);
or U8834 (N_8834,N_8696,N_8640);
nor U8835 (N_8835,N_8613,N_8724);
nand U8836 (N_8836,N_8721,N_8734);
or U8837 (N_8837,N_8602,N_8765);
nand U8838 (N_8838,N_8722,N_8671);
nor U8839 (N_8839,N_8756,N_8761);
nor U8840 (N_8840,N_8631,N_8647);
nor U8841 (N_8841,N_8603,N_8623);
nor U8842 (N_8842,N_8614,N_8658);
or U8843 (N_8843,N_8621,N_8700);
nand U8844 (N_8844,N_8741,N_8736);
xor U8845 (N_8845,N_8757,N_8665);
nor U8846 (N_8846,N_8780,N_8793);
nand U8847 (N_8847,N_8789,N_8704);
nand U8848 (N_8848,N_8698,N_8749);
nor U8849 (N_8849,N_8744,N_8773);
nor U8850 (N_8850,N_8672,N_8713);
and U8851 (N_8851,N_8790,N_8610);
or U8852 (N_8852,N_8690,N_8708);
or U8853 (N_8853,N_8729,N_8605);
nand U8854 (N_8854,N_8787,N_8764);
xnor U8855 (N_8855,N_8688,N_8683);
nand U8856 (N_8856,N_8611,N_8670);
nor U8857 (N_8857,N_8695,N_8778);
and U8858 (N_8858,N_8720,N_8655);
and U8859 (N_8859,N_8636,N_8738);
nor U8860 (N_8860,N_8739,N_8799);
nor U8861 (N_8861,N_8743,N_8715);
xor U8862 (N_8862,N_8711,N_8627);
nand U8863 (N_8863,N_8677,N_8776);
xor U8864 (N_8864,N_8753,N_8726);
or U8865 (N_8865,N_8633,N_8792);
nor U8866 (N_8866,N_8768,N_8667);
xor U8867 (N_8867,N_8682,N_8684);
or U8868 (N_8868,N_8681,N_8727);
or U8869 (N_8869,N_8781,N_8656);
nor U8870 (N_8870,N_8755,N_8771);
nor U8871 (N_8871,N_8679,N_8767);
nand U8872 (N_8872,N_8707,N_8716);
nand U8873 (N_8873,N_8760,N_8737);
nand U8874 (N_8874,N_8709,N_8641);
nor U8875 (N_8875,N_8714,N_8733);
nand U8876 (N_8876,N_8735,N_8798);
or U8877 (N_8877,N_8725,N_8645);
and U8878 (N_8878,N_8784,N_8615);
and U8879 (N_8879,N_8710,N_8635);
nand U8880 (N_8880,N_8754,N_8712);
nand U8881 (N_8881,N_8752,N_8680);
or U8882 (N_8882,N_8701,N_8751);
nand U8883 (N_8883,N_8706,N_8630);
nand U8884 (N_8884,N_8794,N_8742);
and U8885 (N_8885,N_8745,N_8779);
or U8886 (N_8886,N_8625,N_8620);
nand U8887 (N_8887,N_8676,N_8626);
nor U8888 (N_8888,N_8642,N_8762);
nor U8889 (N_8889,N_8634,N_8654);
nor U8890 (N_8890,N_8758,N_8788);
xnor U8891 (N_8891,N_8777,N_8691);
or U8892 (N_8892,N_8786,N_8770);
and U8893 (N_8893,N_8660,N_8750);
or U8894 (N_8894,N_8638,N_8692);
nand U8895 (N_8895,N_8759,N_8649);
and U8896 (N_8896,N_8702,N_8687);
nor U8897 (N_8897,N_8797,N_8772);
and U8898 (N_8898,N_8774,N_8685);
nor U8899 (N_8899,N_8669,N_8604);
and U8900 (N_8900,N_8714,N_8684);
or U8901 (N_8901,N_8780,N_8786);
xor U8902 (N_8902,N_8771,N_8707);
nor U8903 (N_8903,N_8730,N_8701);
nor U8904 (N_8904,N_8687,N_8759);
xnor U8905 (N_8905,N_8742,N_8625);
or U8906 (N_8906,N_8677,N_8628);
or U8907 (N_8907,N_8603,N_8695);
or U8908 (N_8908,N_8794,N_8729);
and U8909 (N_8909,N_8770,N_8654);
nand U8910 (N_8910,N_8640,N_8702);
or U8911 (N_8911,N_8766,N_8621);
xor U8912 (N_8912,N_8626,N_8640);
xnor U8913 (N_8913,N_8780,N_8617);
nand U8914 (N_8914,N_8620,N_8692);
or U8915 (N_8915,N_8796,N_8767);
nand U8916 (N_8916,N_8759,N_8707);
nand U8917 (N_8917,N_8742,N_8601);
or U8918 (N_8918,N_8683,N_8664);
xor U8919 (N_8919,N_8713,N_8780);
nor U8920 (N_8920,N_8755,N_8600);
and U8921 (N_8921,N_8750,N_8683);
nor U8922 (N_8922,N_8662,N_8669);
xor U8923 (N_8923,N_8612,N_8601);
and U8924 (N_8924,N_8794,N_8707);
nand U8925 (N_8925,N_8601,N_8643);
and U8926 (N_8926,N_8627,N_8766);
nor U8927 (N_8927,N_8676,N_8777);
and U8928 (N_8928,N_8654,N_8760);
and U8929 (N_8929,N_8635,N_8761);
and U8930 (N_8930,N_8607,N_8660);
nand U8931 (N_8931,N_8725,N_8732);
nand U8932 (N_8932,N_8710,N_8739);
and U8933 (N_8933,N_8620,N_8737);
nand U8934 (N_8934,N_8656,N_8706);
and U8935 (N_8935,N_8766,N_8732);
nor U8936 (N_8936,N_8730,N_8634);
xnor U8937 (N_8937,N_8656,N_8717);
xor U8938 (N_8938,N_8712,N_8661);
xnor U8939 (N_8939,N_8752,N_8797);
xnor U8940 (N_8940,N_8647,N_8641);
nor U8941 (N_8941,N_8671,N_8793);
xnor U8942 (N_8942,N_8681,N_8757);
or U8943 (N_8943,N_8726,N_8739);
nand U8944 (N_8944,N_8700,N_8686);
and U8945 (N_8945,N_8661,N_8719);
and U8946 (N_8946,N_8602,N_8662);
nor U8947 (N_8947,N_8797,N_8714);
or U8948 (N_8948,N_8670,N_8755);
xnor U8949 (N_8949,N_8731,N_8701);
or U8950 (N_8950,N_8615,N_8651);
nand U8951 (N_8951,N_8785,N_8771);
or U8952 (N_8952,N_8704,N_8706);
xnor U8953 (N_8953,N_8745,N_8703);
and U8954 (N_8954,N_8626,N_8712);
nor U8955 (N_8955,N_8722,N_8706);
and U8956 (N_8956,N_8713,N_8720);
and U8957 (N_8957,N_8798,N_8782);
xnor U8958 (N_8958,N_8769,N_8712);
nand U8959 (N_8959,N_8644,N_8638);
xor U8960 (N_8960,N_8649,N_8740);
and U8961 (N_8961,N_8729,N_8668);
nor U8962 (N_8962,N_8630,N_8652);
xnor U8963 (N_8963,N_8728,N_8785);
or U8964 (N_8964,N_8663,N_8668);
nand U8965 (N_8965,N_8723,N_8610);
xnor U8966 (N_8966,N_8664,N_8646);
xnor U8967 (N_8967,N_8607,N_8677);
or U8968 (N_8968,N_8622,N_8779);
or U8969 (N_8969,N_8653,N_8627);
or U8970 (N_8970,N_8766,N_8617);
or U8971 (N_8971,N_8720,N_8787);
or U8972 (N_8972,N_8782,N_8626);
and U8973 (N_8973,N_8673,N_8667);
nand U8974 (N_8974,N_8673,N_8658);
or U8975 (N_8975,N_8688,N_8758);
xnor U8976 (N_8976,N_8759,N_8673);
or U8977 (N_8977,N_8725,N_8794);
and U8978 (N_8978,N_8734,N_8789);
nor U8979 (N_8979,N_8756,N_8727);
xor U8980 (N_8980,N_8748,N_8790);
nor U8981 (N_8981,N_8728,N_8619);
or U8982 (N_8982,N_8682,N_8677);
xnor U8983 (N_8983,N_8620,N_8632);
and U8984 (N_8984,N_8736,N_8727);
nand U8985 (N_8985,N_8688,N_8608);
and U8986 (N_8986,N_8627,N_8778);
xor U8987 (N_8987,N_8732,N_8798);
nand U8988 (N_8988,N_8750,N_8686);
nand U8989 (N_8989,N_8676,N_8612);
nand U8990 (N_8990,N_8743,N_8764);
xor U8991 (N_8991,N_8742,N_8657);
and U8992 (N_8992,N_8719,N_8681);
and U8993 (N_8993,N_8749,N_8607);
xnor U8994 (N_8994,N_8745,N_8637);
or U8995 (N_8995,N_8730,N_8675);
and U8996 (N_8996,N_8610,N_8609);
or U8997 (N_8997,N_8727,N_8726);
and U8998 (N_8998,N_8679,N_8783);
nor U8999 (N_8999,N_8739,N_8778);
nand U9000 (N_9000,N_8906,N_8864);
nand U9001 (N_9001,N_8867,N_8979);
nor U9002 (N_9002,N_8839,N_8913);
xnor U9003 (N_9003,N_8896,N_8914);
nor U9004 (N_9004,N_8810,N_8882);
and U9005 (N_9005,N_8878,N_8915);
nor U9006 (N_9006,N_8980,N_8916);
nor U9007 (N_9007,N_8803,N_8822);
nor U9008 (N_9008,N_8889,N_8801);
xor U9009 (N_9009,N_8924,N_8904);
nor U9010 (N_9010,N_8826,N_8928);
xnor U9011 (N_9011,N_8912,N_8816);
nand U9012 (N_9012,N_8834,N_8974);
or U9013 (N_9013,N_8892,N_8960);
and U9014 (N_9014,N_8921,N_8901);
or U9015 (N_9015,N_8805,N_8987);
or U9016 (N_9016,N_8978,N_8966);
xnor U9017 (N_9017,N_8927,N_8871);
xnor U9018 (N_9018,N_8910,N_8903);
nor U9019 (N_9019,N_8932,N_8954);
and U9020 (N_9020,N_8837,N_8992);
xnor U9021 (N_9021,N_8929,N_8844);
xnor U9022 (N_9022,N_8829,N_8888);
nor U9023 (N_9023,N_8900,N_8847);
xnor U9024 (N_9024,N_8965,N_8948);
nor U9025 (N_9025,N_8902,N_8956);
xnor U9026 (N_9026,N_8946,N_8975);
xor U9027 (N_9027,N_8938,N_8865);
or U9028 (N_9028,N_8957,N_8973);
or U9029 (N_9029,N_8862,N_8977);
or U9030 (N_9030,N_8872,N_8989);
nand U9031 (N_9031,N_8935,N_8806);
and U9032 (N_9032,N_8962,N_8982);
nand U9033 (N_9033,N_8818,N_8999);
xnor U9034 (N_9034,N_8836,N_8814);
nor U9035 (N_9035,N_8808,N_8905);
xnor U9036 (N_9036,N_8853,N_8859);
and U9037 (N_9037,N_8942,N_8991);
nor U9038 (N_9038,N_8998,N_8953);
or U9039 (N_9039,N_8870,N_8994);
or U9040 (N_9040,N_8855,N_8841);
xor U9041 (N_9041,N_8968,N_8883);
xor U9042 (N_9042,N_8843,N_8918);
nor U9043 (N_9043,N_8894,N_8934);
nor U9044 (N_9044,N_8940,N_8925);
or U9045 (N_9045,N_8851,N_8858);
xnor U9046 (N_9046,N_8926,N_8959);
xor U9047 (N_9047,N_8874,N_8852);
nand U9048 (N_9048,N_8823,N_8885);
and U9049 (N_9049,N_8817,N_8831);
nand U9050 (N_9050,N_8950,N_8952);
and U9051 (N_9051,N_8804,N_8825);
xor U9052 (N_9052,N_8908,N_8827);
and U9053 (N_9053,N_8930,N_8949);
nand U9054 (N_9054,N_8936,N_8891);
xnor U9055 (N_9055,N_8866,N_8832);
nand U9056 (N_9056,N_8856,N_8879);
nor U9057 (N_9057,N_8923,N_8869);
xnor U9058 (N_9058,N_8984,N_8983);
nand U9059 (N_9059,N_8881,N_8838);
or U9060 (N_9060,N_8861,N_8917);
and U9061 (N_9061,N_8854,N_8812);
nor U9062 (N_9062,N_8922,N_8986);
nand U9063 (N_9063,N_8944,N_8828);
and U9064 (N_9064,N_8857,N_8990);
and U9065 (N_9065,N_8863,N_8976);
nor U9066 (N_9066,N_8860,N_8951);
xor U9067 (N_9067,N_8845,N_8988);
nor U9068 (N_9068,N_8875,N_8846);
nand U9069 (N_9069,N_8920,N_8886);
or U9070 (N_9070,N_8819,N_8947);
xnor U9071 (N_9071,N_8820,N_8969);
and U9072 (N_9072,N_8821,N_8993);
nand U9073 (N_9073,N_8995,N_8997);
xor U9074 (N_9074,N_8981,N_8911);
xor U9075 (N_9075,N_8880,N_8964);
and U9076 (N_9076,N_8945,N_8970);
nand U9077 (N_9077,N_8963,N_8849);
xnor U9078 (N_9078,N_8895,N_8876);
nand U9079 (N_9079,N_8941,N_8933);
or U9080 (N_9080,N_8815,N_8967);
nand U9081 (N_9081,N_8890,N_8877);
or U9082 (N_9082,N_8809,N_8811);
or U9083 (N_9083,N_8931,N_8873);
or U9084 (N_9084,N_8807,N_8830);
or U9085 (N_9085,N_8887,N_8840);
and U9086 (N_9086,N_8972,N_8985);
nand U9087 (N_9087,N_8943,N_8813);
xor U9088 (N_9088,N_8937,N_8833);
nand U9089 (N_9089,N_8996,N_8884);
or U9090 (N_9090,N_8955,N_8971);
xnor U9091 (N_9091,N_8898,N_8909);
nor U9092 (N_9092,N_8868,N_8802);
or U9093 (N_9093,N_8850,N_8939);
xor U9094 (N_9094,N_8824,N_8919);
or U9095 (N_9095,N_8958,N_8800);
nand U9096 (N_9096,N_8897,N_8961);
nand U9097 (N_9097,N_8848,N_8842);
or U9098 (N_9098,N_8899,N_8893);
or U9099 (N_9099,N_8907,N_8835);
and U9100 (N_9100,N_8965,N_8952);
or U9101 (N_9101,N_8949,N_8965);
and U9102 (N_9102,N_8812,N_8879);
and U9103 (N_9103,N_8838,N_8802);
and U9104 (N_9104,N_8977,N_8923);
nor U9105 (N_9105,N_8876,N_8953);
xnor U9106 (N_9106,N_8979,N_8853);
and U9107 (N_9107,N_8811,N_8951);
and U9108 (N_9108,N_8881,N_8812);
or U9109 (N_9109,N_8882,N_8912);
nor U9110 (N_9110,N_8924,N_8921);
nand U9111 (N_9111,N_8992,N_8877);
xor U9112 (N_9112,N_8961,N_8844);
and U9113 (N_9113,N_8803,N_8843);
nor U9114 (N_9114,N_8889,N_8865);
xnor U9115 (N_9115,N_8852,N_8859);
or U9116 (N_9116,N_8982,N_8993);
or U9117 (N_9117,N_8847,N_8913);
or U9118 (N_9118,N_8881,N_8970);
nand U9119 (N_9119,N_8828,N_8900);
xor U9120 (N_9120,N_8943,N_8876);
nor U9121 (N_9121,N_8802,N_8918);
or U9122 (N_9122,N_8848,N_8823);
and U9123 (N_9123,N_8947,N_8876);
xnor U9124 (N_9124,N_8814,N_8849);
and U9125 (N_9125,N_8989,N_8825);
or U9126 (N_9126,N_8993,N_8872);
nor U9127 (N_9127,N_8989,N_8920);
and U9128 (N_9128,N_8910,N_8961);
nand U9129 (N_9129,N_8819,N_8948);
nor U9130 (N_9130,N_8880,N_8851);
nor U9131 (N_9131,N_8883,N_8871);
and U9132 (N_9132,N_8929,N_8950);
nor U9133 (N_9133,N_8961,N_8950);
xnor U9134 (N_9134,N_8909,N_8911);
or U9135 (N_9135,N_8839,N_8930);
and U9136 (N_9136,N_8875,N_8952);
nand U9137 (N_9137,N_8898,N_8936);
nand U9138 (N_9138,N_8976,N_8964);
and U9139 (N_9139,N_8958,N_8995);
xnor U9140 (N_9140,N_8807,N_8838);
xor U9141 (N_9141,N_8826,N_8952);
nor U9142 (N_9142,N_8901,N_8952);
or U9143 (N_9143,N_8904,N_8981);
nor U9144 (N_9144,N_8807,N_8841);
xnor U9145 (N_9145,N_8987,N_8837);
xor U9146 (N_9146,N_8930,N_8813);
or U9147 (N_9147,N_8957,N_8909);
and U9148 (N_9148,N_8813,N_8971);
or U9149 (N_9149,N_8846,N_8992);
or U9150 (N_9150,N_8964,N_8940);
nor U9151 (N_9151,N_8948,N_8843);
xnor U9152 (N_9152,N_8950,N_8932);
nor U9153 (N_9153,N_8890,N_8863);
and U9154 (N_9154,N_8812,N_8954);
or U9155 (N_9155,N_8849,N_8962);
and U9156 (N_9156,N_8990,N_8829);
and U9157 (N_9157,N_8960,N_8961);
nor U9158 (N_9158,N_8909,N_8910);
xnor U9159 (N_9159,N_8945,N_8975);
or U9160 (N_9160,N_8953,N_8894);
nand U9161 (N_9161,N_8858,N_8812);
and U9162 (N_9162,N_8878,N_8873);
nor U9163 (N_9163,N_8891,N_8934);
nand U9164 (N_9164,N_8832,N_8840);
nor U9165 (N_9165,N_8998,N_8982);
and U9166 (N_9166,N_8949,N_8890);
or U9167 (N_9167,N_8834,N_8854);
and U9168 (N_9168,N_8943,N_8811);
nand U9169 (N_9169,N_8954,N_8916);
nor U9170 (N_9170,N_8800,N_8825);
xnor U9171 (N_9171,N_8983,N_8869);
nand U9172 (N_9172,N_8907,N_8877);
xor U9173 (N_9173,N_8930,N_8886);
xnor U9174 (N_9174,N_8893,N_8827);
nor U9175 (N_9175,N_8805,N_8999);
xnor U9176 (N_9176,N_8830,N_8867);
nor U9177 (N_9177,N_8930,N_8902);
and U9178 (N_9178,N_8816,N_8955);
nor U9179 (N_9179,N_8914,N_8888);
or U9180 (N_9180,N_8981,N_8922);
nand U9181 (N_9181,N_8845,N_8802);
nand U9182 (N_9182,N_8976,N_8866);
or U9183 (N_9183,N_8982,N_8917);
nand U9184 (N_9184,N_8840,N_8805);
nor U9185 (N_9185,N_8991,N_8948);
and U9186 (N_9186,N_8968,N_8882);
xor U9187 (N_9187,N_8906,N_8917);
nand U9188 (N_9188,N_8898,N_8837);
xor U9189 (N_9189,N_8883,N_8898);
nand U9190 (N_9190,N_8954,N_8929);
and U9191 (N_9191,N_8870,N_8896);
nor U9192 (N_9192,N_8980,N_8874);
and U9193 (N_9193,N_8922,N_8928);
xnor U9194 (N_9194,N_8823,N_8901);
and U9195 (N_9195,N_8918,N_8852);
and U9196 (N_9196,N_8984,N_8804);
xor U9197 (N_9197,N_8944,N_8964);
xor U9198 (N_9198,N_8859,N_8822);
nor U9199 (N_9199,N_8887,N_8857);
or U9200 (N_9200,N_9017,N_9185);
nor U9201 (N_9201,N_9147,N_9031);
nor U9202 (N_9202,N_9187,N_9137);
nand U9203 (N_9203,N_9067,N_9077);
nand U9204 (N_9204,N_9060,N_9135);
or U9205 (N_9205,N_9195,N_9033);
xnor U9206 (N_9206,N_9144,N_9088);
xor U9207 (N_9207,N_9120,N_9086);
and U9208 (N_9208,N_9024,N_9070);
or U9209 (N_9209,N_9157,N_9169);
nand U9210 (N_9210,N_9133,N_9174);
nand U9211 (N_9211,N_9117,N_9110);
nand U9212 (N_9212,N_9094,N_9136);
or U9213 (N_9213,N_9007,N_9038);
xnor U9214 (N_9214,N_9193,N_9107);
or U9215 (N_9215,N_9116,N_9091);
xor U9216 (N_9216,N_9182,N_9127);
nor U9217 (N_9217,N_9030,N_9064);
nand U9218 (N_9218,N_9044,N_9001);
and U9219 (N_9219,N_9037,N_9160);
nand U9220 (N_9220,N_9059,N_9139);
nand U9221 (N_9221,N_9095,N_9198);
xor U9222 (N_9222,N_9047,N_9022);
xor U9223 (N_9223,N_9162,N_9053);
and U9224 (N_9224,N_9009,N_9166);
or U9225 (N_9225,N_9036,N_9050);
and U9226 (N_9226,N_9084,N_9102);
and U9227 (N_9227,N_9002,N_9154);
nor U9228 (N_9228,N_9199,N_9076);
or U9229 (N_9229,N_9034,N_9075);
or U9230 (N_9230,N_9054,N_9003);
nand U9231 (N_9231,N_9104,N_9040);
nand U9232 (N_9232,N_9122,N_9069);
nor U9233 (N_9233,N_9015,N_9100);
nand U9234 (N_9234,N_9010,N_9073);
xor U9235 (N_9235,N_9140,N_9026);
and U9236 (N_9236,N_9066,N_9051);
nor U9237 (N_9237,N_9008,N_9131);
nor U9238 (N_9238,N_9138,N_9098);
xnor U9239 (N_9239,N_9012,N_9025);
xnor U9240 (N_9240,N_9079,N_9105);
nor U9241 (N_9241,N_9065,N_9168);
or U9242 (N_9242,N_9078,N_9042);
xor U9243 (N_9243,N_9124,N_9189);
or U9244 (N_9244,N_9179,N_9096);
nand U9245 (N_9245,N_9197,N_9048);
nor U9246 (N_9246,N_9129,N_9152);
xnor U9247 (N_9247,N_9103,N_9000);
xor U9248 (N_9248,N_9141,N_9020);
nand U9249 (N_9249,N_9004,N_9057);
nand U9250 (N_9250,N_9153,N_9043);
and U9251 (N_9251,N_9072,N_9013);
xor U9252 (N_9252,N_9019,N_9130);
or U9253 (N_9253,N_9142,N_9063);
nor U9254 (N_9254,N_9027,N_9196);
or U9255 (N_9255,N_9109,N_9183);
and U9256 (N_9256,N_9194,N_9023);
and U9257 (N_9257,N_9016,N_9118);
and U9258 (N_9258,N_9014,N_9188);
nor U9259 (N_9259,N_9167,N_9021);
or U9260 (N_9260,N_9155,N_9062);
or U9261 (N_9261,N_9032,N_9143);
nand U9262 (N_9262,N_9165,N_9145);
xnor U9263 (N_9263,N_9055,N_9006);
xor U9264 (N_9264,N_9149,N_9181);
nand U9265 (N_9265,N_9148,N_9028);
nor U9266 (N_9266,N_9058,N_9005);
xnor U9267 (N_9267,N_9082,N_9180);
xor U9268 (N_9268,N_9074,N_9011);
or U9269 (N_9269,N_9191,N_9126);
nor U9270 (N_9270,N_9128,N_9113);
xor U9271 (N_9271,N_9101,N_9045);
nor U9272 (N_9272,N_9177,N_9175);
nor U9273 (N_9273,N_9090,N_9099);
nand U9274 (N_9274,N_9186,N_9052);
nand U9275 (N_9275,N_9119,N_9184);
nor U9276 (N_9276,N_9150,N_9068);
nand U9277 (N_9277,N_9061,N_9114);
or U9278 (N_9278,N_9089,N_9159);
nand U9279 (N_9279,N_9178,N_9111);
and U9280 (N_9280,N_9161,N_9085);
or U9281 (N_9281,N_9151,N_9071);
or U9282 (N_9282,N_9163,N_9132);
and U9283 (N_9283,N_9106,N_9190);
and U9284 (N_9284,N_9172,N_9171);
or U9285 (N_9285,N_9081,N_9176);
nand U9286 (N_9286,N_9018,N_9121);
and U9287 (N_9287,N_9093,N_9115);
xor U9288 (N_9288,N_9134,N_9035);
nand U9289 (N_9289,N_9080,N_9164);
or U9290 (N_9290,N_9108,N_9146);
xor U9291 (N_9291,N_9083,N_9173);
xor U9292 (N_9292,N_9123,N_9029);
or U9293 (N_9293,N_9039,N_9056);
or U9294 (N_9294,N_9170,N_9092);
and U9295 (N_9295,N_9049,N_9192);
or U9296 (N_9296,N_9041,N_9112);
xnor U9297 (N_9297,N_9125,N_9087);
and U9298 (N_9298,N_9097,N_9156);
nand U9299 (N_9299,N_9158,N_9046);
xor U9300 (N_9300,N_9072,N_9043);
and U9301 (N_9301,N_9145,N_9146);
and U9302 (N_9302,N_9058,N_9018);
and U9303 (N_9303,N_9168,N_9117);
or U9304 (N_9304,N_9183,N_9129);
nand U9305 (N_9305,N_9018,N_9147);
or U9306 (N_9306,N_9104,N_9177);
and U9307 (N_9307,N_9001,N_9058);
and U9308 (N_9308,N_9173,N_9166);
xnor U9309 (N_9309,N_9100,N_9058);
nor U9310 (N_9310,N_9084,N_9167);
xnor U9311 (N_9311,N_9015,N_9054);
nand U9312 (N_9312,N_9174,N_9123);
nor U9313 (N_9313,N_9116,N_9162);
nor U9314 (N_9314,N_9058,N_9048);
nor U9315 (N_9315,N_9047,N_9108);
or U9316 (N_9316,N_9119,N_9097);
nand U9317 (N_9317,N_9195,N_9135);
nand U9318 (N_9318,N_9132,N_9167);
or U9319 (N_9319,N_9133,N_9144);
nor U9320 (N_9320,N_9149,N_9083);
nand U9321 (N_9321,N_9122,N_9192);
nor U9322 (N_9322,N_9086,N_9000);
xnor U9323 (N_9323,N_9078,N_9142);
and U9324 (N_9324,N_9029,N_9043);
nor U9325 (N_9325,N_9115,N_9038);
nand U9326 (N_9326,N_9023,N_9067);
and U9327 (N_9327,N_9163,N_9154);
and U9328 (N_9328,N_9015,N_9003);
or U9329 (N_9329,N_9003,N_9162);
or U9330 (N_9330,N_9059,N_9091);
nand U9331 (N_9331,N_9003,N_9063);
and U9332 (N_9332,N_9161,N_9105);
nand U9333 (N_9333,N_9024,N_9030);
and U9334 (N_9334,N_9051,N_9148);
nor U9335 (N_9335,N_9124,N_9031);
xnor U9336 (N_9336,N_9157,N_9140);
nor U9337 (N_9337,N_9096,N_9126);
xnor U9338 (N_9338,N_9019,N_9136);
nand U9339 (N_9339,N_9109,N_9020);
nor U9340 (N_9340,N_9025,N_9009);
nor U9341 (N_9341,N_9094,N_9110);
nand U9342 (N_9342,N_9056,N_9076);
nand U9343 (N_9343,N_9157,N_9039);
nor U9344 (N_9344,N_9000,N_9072);
nor U9345 (N_9345,N_9134,N_9131);
and U9346 (N_9346,N_9126,N_9041);
or U9347 (N_9347,N_9118,N_9059);
and U9348 (N_9348,N_9124,N_9092);
or U9349 (N_9349,N_9032,N_9120);
nor U9350 (N_9350,N_9199,N_9016);
nor U9351 (N_9351,N_9139,N_9158);
nor U9352 (N_9352,N_9013,N_9198);
xnor U9353 (N_9353,N_9058,N_9113);
xnor U9354 (N_9354,N_9185,N_9154);
and U9355 (N_9355,N_9054,N_9005);
or U9356 (N_9356,N_9195,N_9054);
xnor U9357 (N_9357,N_9109,N_9133);
xnor U9358 (N_9358,N_9181,N_9053);
nand U9359 (N_9359,N_9147,N_9172);
xor U9360 (N_9360,N_9135,N_9198);
nor U9361 (N_9361,N_9164,N_9054);
or U9362 (N_9362,N_9118,N_9160);
xnor U9363 (N_9363,N_9069,N_9117);
and U9364 (N_9364,N_9056,N_9130);
nand U9365 (N_9365,N_9124,N_9187);
or U9366 (N_9366,N_9109,N_9037);
nand U9367 (N_9367,N_9151,N_9183);
xnor U9368 (N_9368,N_9130,N_9142);
nor U9369 (N_9369,N_9028,N_9174);
xnor U9370 (N_9370,N_9093,N_9177);
nor U9371 (N_9371,N_9102,N_9004);
nor U9372 (N_9372,N_9003,N_9027);
xor U9373 (N_9373,N_9006,N_9124);
xor U9374 (N_9374,N_9034,N_9069);
nor U9375 (N_9375,N_9104,N_9128);
xnor U9376 (N_9376,N_9129,N_9089);
nand U9377 (N_9377,N_9143,N_9162);
nand U9378 (N_9378,N_9086,N_9179);
xnor U9379 (N_9379,N_9129,N_9063);
or U9380 (N_9380,N_9090,N_9026);
and U9381 (N_9381,N_9150,N_9011);
or U9382 (N_9382,N_9098,N_9143);
xor U9383 (N_9383,N_9139,N_9143);
and U9384 (N_9384,N_9019,N_9101);
xnor U9385 (N_9385,N_9103,N_9190);
nand U9386 (N_9386,N_9103,N_9009);
and U9387 (N_9387,N_9076,N_9136);
and U9388 (N_9388,N_9083,N_9160);
xor U9389 (N_9389,N_9184,N_9004);
and U9390 (N_9390,N_9166,N_9151);
and U9391 (N_9391,N_9066,N_9146);
xnor U9392 (N_9392,N_9035,N_9102);
nor U9393 (N_9393,N_9013,N_9189);
nand U9394 (N_9394,N_9179,N_9137);
nand U9395 (N_9395,N_9162,N_9061);
nand U9396 (N_9396,N_9025,N_9061);
and U9397 (N_9397,N_9080,N_9020);
and U9398 (N_9398,N_9022,N_9153);
or U9399 (N_9399,N_9046,N_9168);
and U9400 (N_9400,N_9325,N_9303);
nor U9401 (N_9401,N_9351,N_9269);
nand U9402 (N_9402,N_9309,N_9216);
and U9403 (N_9403,N_9297,N_9391);
nor U9404 (N_9404,N_9259,N_9247);
and U9405 (N_9405,N_9235,N_9346);
nor U9406 (N_9406,N_9249,N_9360);
or U9407 (N_9407,N_9243,N_9385);
and U9408 (N_9408,N_9217,N_9227);
nand U9409 (N_9409,N_9350,N_9337);
nor U9410 (N_9410,N_9242,N_9368);
nor U9411 (N_9411,N_9212,N_9278);
and U9412 (N_9412,N_9336,N_9327);
xnor U9413 (N_9413,N_9356,N_9328);
and U9414 (N_9414,N_9257,N_9284);
and U9415 (N_9415,N_9210,N_9205);
or U9416 (N_9416,N_9248,N_9381);
xnor U9417 (N_9417,N_9285,N_9224);
or U9418 (N_9418,N_9316,N_9355);
and U9419 (N_9419,N_9320,N_9260);
xor U9420 (N_9420,N_9252,N_9296);
or U9421 (N_9421,N_9312,N_9345);
xnor U9422 (N_9422,N_9365,N_9341);
nand U9423 (N_9423,N_9245,N_9315);
and U9424 (N_9424,N_9335,N_9322);
nand U9425 (N_9425,N_9293,N_9307);
nand U9426 (N_9426,N_9342,N_9398);
nor U9427 (N_9427,N_9330,N_9270);
and U9428 (N_9428,N_9372,N_9240);
xnor U9429 (N_9429,N_9206,N_9374);
nor U9430 (N_9430,N_9380,N_9347);
or U9431 (N_9431,N_9295,N_9213);
xor U9432 (N_9432,N_9305,N_9277);
or U9433 (N_9433,N_9340,N_9314);
or U9434 (N_9434,N_9283,N_9203);
and U9435 (N_9435,N_9384,N_9258);
and U9436 (N_9436,N_9253,N_9207);
or U9437 (N_9437,N_9282,N_9299);
nor U9438 (N_9438,N_9265,N_9236);
xor U9439 (N_9439,N_9239,N_9324);
xnor U9440 (N_9440,N_9308,N_9220);
and U9441 (N_9441,N_9382,N_9289);
nand U9442 (N_9442,N_9317,N_9311);
xor U9443 (N_9443,N_9294,N_9396);
and U9444 (N_9444,N_9228,N_9377);
xnor U9445 (N_9445,N_9202,N_9358);
nand U9446 (N_9446,N_9225,N_9389);
and U9447 (N_9447,N_9219,N_9376);
and U9448 (N_9448,N_9233,N_9390);
xnor U9449 (N_9449,N_9211,N_9275);
nand U9450 (N_9450,N_9254,N_9338);
and U9451 (N_9451,N_9201,N_9261);
nor U9452 (N_9452,N_9250,N_9367);
xor U9453 (N_9453,N_9244,N_9298);
or U9454 (N_9454,N_9238,N_9321);
xnor U9455 (N_9455,N_9369,N_9383);
and U9456 (N_9456,N_9241,N_9288);
nor U9457 (N_9457,N_9281,N_9287);
xnor U9458 (N_9458,N_9229,N_9393);
nand U9459 (N_9459,N_9373,N_9392);
nand U9460 (N_9460,N_9301,N_9348);
xor U9461 (N_9461,N_9333,N_9388);
nand U9462 (N_9462,N_9329,N_9302);
nor U9463 (N_9463,N_9349,N_9230);
or U9464 (N_9464,N_9354,N_9371);
or U9465 (N_9465,N_9352,N_9318);
xor U9466 (N_9466,N_9386,N_9370);
nand U9467 (N_9467,N_9357,N_9378);
or U9468 (N_9468,N_9223,N_9313);
xnor U9469 (N_9469,N_9221,N_9251);
and U9470 (N_9470,N_9226,N_9266);
nor U9471 (N_9471,N_9361,N_9319);
or U9472 (N_9472,N_9326,N_9300);
nand U9473 (N_9473,N_9273,N_9366);
nand U9474 (N_9474,N_9399,N_9268);
xor U9475 (N_9475,N_9274,N_9364);
or U9476 (N_9476,N_9290,N_9231);
and U9477 (N_9477,N_9363,N_9395);
or U9478 (N_9478,N_9215,N_9262);
xnor U9479 (N_9479,N_9280,N_9222);
xor U9480 (N_9480,N_9204,N_9306);
xnor U9481 (N_9481,N_9334,N_9272);
or U9482 (N_9482,N_9234,N_9267);
nor U9483 (N_9483,N_9237,N_9375);
and U9484 (N_9484,N_9359,N_9323);
or U9485 (N_9485,N_9208,N_9387);
and U9486 (N_9486,N_9394,N_9343);
xor U9487 (N_9487,N_9339,N_9246);
nor U9488 (N_9488,N_9255,N_9362);
nand U9489 (N_9489,N_9279,N_9263);
or U9490 (N_9490,N_9353,N_9397);
nand U9491 (N_9491,N_9209,N_9304);
nand U9492 (N_9492,N_9232,N_9379);
and U9493 (N_9493,N_9332,N_9292);
nand U9494 (N_9494,N_9264,N_9344);
or U9495 (N_9495,N_9331,N_9291);
xor U9496 (N_9496,N_9200,N_9218);
or U9497 (N_9497,N_9276,N_9271);
nor U9498 (N_9498,N_9310,N_9256);
nor U9499 (N_9499,N_9214,N_9286);
nor U9500 (N_9500,N_9273,N_9276);
and U9501 (N_9501,N_9306,N_9288);
or U9502 (N_9502,N_9308,N_9298);
xor U9503 (N_9503,N_9281,N_9231);
and U9504 (N_9504,N_9303,N_9234);
xnor U9505 (N_9505,N_9283,N_9311);
nand U9506 (N_9506,N_9207,N_9314);
xor U9507 (N_9507,N_9351,N_9270);
nor U9508 (N_9508,N_9329,N_9261);
nand U9509 (N_9509,N_9314,N_9277);
xor U9510 (N_9510,N_9351,N_9350);
and U9511 (N_9511,N_9385,N_9380);
nor U9512 (N_9512,N_9379,N_9289);
and U9513 (N_9513,N_9300,N_9257);
xor U9514 (N_9514,N_9215,N_9304);
and U9515 (N_9515,N_9205,N_9378);
nor U9516 (N_9516,N_9224,N_9366);
and U9517 (N_9517,N_9392,N_9381);
nand U9518 (N_9518,N_9202,N_9273);
xor U9519 (N_9519,N_9398,N_9325);
nand U9520 (N_9520,N_9379,N_9217);
nor U9521 (N_9521,N_9322,N_9247);
xor U9522 (N_9522,N_9299,N_9328);
nand U9523 (N_9523,N_9362,N_9355);
nand U9524 (N_9524,N_9331,N_9238);
nand U9525 (N_9525,N_9212,N_9311);
nand U9526 (N_9526,N_9293,N_9328);
and U9527 (N_9527,N_9384,N_9311);
and U9528 (N_9528,N_9216,N_9275);
nand U9529 (N_9529,N_9259,N_9268);
and U9530 (N_9530,N_9338,N_9320);
and U9531 (N_9531,N_9222,N_9332);
or U9532 (N_9532,N_9225,N_9200);
or U9533 (N_9533,N_9244,N_9232);
and U9534 (N_9534,N_9354,N_9258);
and U9535 (N_9535,N_9397,N_9290);
and U9536 (N_9536,N_9336,N_9333);
nand U9537 (N_9537,N_9342,N_9207);
or U9538 (N_9538,N_9320,N_9313);
and U9539 (N_9539,N_9276,N_9314);
and U9540 (N_9540,N_9393,N_9387);
and U9541 (N_9541,N_9237,N_9394);
or U9542 (N_9542,N_9304,N_9381);
and U9543 (N_9543,N_9382,N_9387);
or U9544 (N_9544,N_9303,N_9242);
nor U9545 (N_9545,N_9334,N_9352);
or U9546 (N_9546,N_9272,N_9212);
xor U9547 (N_9547,N_9296,N_9290);
nor U9548 (N_9548,N_9372,N_9378);
and U9549 (N_9549,N_9283,N_9289);
nand U9550 (N_9550,N_9328,N_9329);
or U9551 (N_9551,N_9233,N_9340);
xnor U9552 (N_9552,N_9331,N_9218);
xor U9553 (N_9553,N_9210,N_9286);
xor U9554 (N_9554,N_9253,N_9325);
xnor U9555 (N_9555,N_9288,N_9386);
or U9556 (N_9556,N_9244,N_9217);
or U9557 (N_9557,N_9211,N_9399);
nand U9558 (N_9558,N_9203,N_9321);
xor U9559 (N_9559,N_9391,N_9345);
or U9560 (N_9560,N_9306,N_9328);
nand U9561 (N_9561,N_9214,N_9339);
nand U9562 (N_9562,N_9248,N_9232);
xor U9563 (N_9563,N_9229,N_9345);
nand U9564 (N_9564,N_9296,N_9295);
nor U9565 (N_9565,N_9345,N_9205);
xnor U9566 (N_9566,N_9386,N_9286);
nand U9567 (N_9567,N_9384,N_9359);
and U9568 (N_9568,N_9261,N_9243);
nor U9569 (N_9569,N_9252,N_9267);
nand U9570 (N_9570,N_9297,N_9219);
nand U9571 (N_9571,N_9204,N_9311);
or U9572 (N_9572,N_9395,N_9340);
and U9573 (N_9573,N_9286,N_9323);
nor U9574 (N_9574,N_9258,N_9206);
nor U9575 (N_9575,N_9389,N_9257);
nand U9576 (N_9576,N_9223,N_9359);
nand U9577 (N_9577,N_9320,N_9367);
xor U9578 (N_9578,N_9297,N_9355);
and U9579 (N_9579,N_9344,N_9284);
or U9580 (N_9580,N_9312,N_9276);
and U9581 (N_9581,N_9296,N_9227);
nand U9582 (N_9582,N_9321,N_9300);
nand U9583 (N_9583,N_9278,N_9382);
nand U9584 (N_9584,N_9285,N_9280);
nand U9585 (N_9585,N_9241,N_9214);
nand U9586 (N_9586,N_9259,N_9230);
nand U9587 (N_9587,N_9339,N_9351);
and U9588 (N_9588,N_9229,N_9247);
nand U9589 (N_9589,N_9326,N_9268);
and U9590 (N_9590,N_9266,N_9303);
nor U9591 (N_9591,N_9394,N_9351);
nand U9592 (N_9592,N_9352,N_9251);
and U9593 (N_9593,N_9201,N_9244);
nor U9594 (N_9594,N_9340,N_9278);
nand U9595 (N_9595,N_9200,N_9244);
xnor U9596 (N_9596,N_9257,N_9213);
nand U9597 (N_9597,N_9227,N_9208);
nand U9598 (N_9598,N_9277,N_9316);
and U9599 (N_9599,N_9337,N_9204);
xnor U9600 (N_9600,N_9403,N_9439);
or U9601 (N_9601,N_9452,N_9474);
and U9602 (N_9602,N_9479,N_9504);
and U9603 (N_9603,N_9496,N_9543);
nand U9604 (N_9604,N_9512,N_9409);
or U9605 (N_9605,N_9402,N_9498);
nand U9606 (N_9606,N_9509,N_9541);
nor U9607 (N_9607,N_9533,N_9467);
and U9608 (N_9608,N_9511,N_9557);
nor U9609 (N_9609,N_9491,N_9429);
and U9610 (N_9610,N_9428,N_9470);
or U9611 (N_9611,N_9532,N_9586);
nand U9612 (N_9612,N_9539,N_9523);
xor U9613 (N_9613,N_9577,N_9417);
xor U9614 (N_9614,N_9550,N_9562);
nor U9615 (N_9615,N_9443,N_9423);
nor U9616 (N_9616,N_9463,N_9450);
or U9617 (N_9617,N_9489,N_9484);
nand U9618 (N_9618,N_9441,N_9535);
or U9619 (N_9619,N_9574,N_9462);
xor U9620 (N_9620,N_9405,N_9584);
nand U9621 (N_9621,N_9421,N_9570);
xnor U9622 (N_9622,N_9475,N_9506);
nor U9623 (N_9623,N_9449,N_9590);
and U9624 (N_9624,N_9499,N_9418);
nor U9625 (N_9625,N_9566,N_9519);
nor U9626 (N_9626,N_9426,N_9435);
nand U9627 (N_9627,N_9444,N_9442);
nand U9628 (N_9628,N_9582,N_9599);
xor U9629 (N_9629,N_9513,N_9478);
xnor U9630 (N_9630,N_9416,N_9553);
nor U9631 (N_9631,N_9455,N_9457);
and U9632 (N_9632,N_9583,N_9549);
or U9633 (N_9633,N_9501,N_9427);
nand U9634 (N_9634,N_9596,N_9406);
and U9635 (N_9635,N_9561,N_9530);
xnor U9636 (N_9636,N_9581,N_9521);
or U9637 (N_9637,N_9548,N_9560);
nor U9638 (N_9638,N_9554,N_9516);
nor U9639 (N_9639,N_9465,N_9414);
xnor U9640 (N_9640,N_9515,N_9424);
xor U9641 (N_9641,N_9589,N_9567);
xnor U9642 (N_9642,N_9578,N_9485);
or U9643 (N_9643,N_9555,N_9454);
nor U9644 (N_9644,N_9432,N_9447);
xnor U9645 (N_9645,N_9572,N_9565);
and U9646 (N_9646,N_9524,N_9448);
nor U9647 (N_9647,N_9453,N_9525);
xnor U9648 (N_9648,N_9587,N_9413);
xor U9649 (N_9649,N_9522,N_9547);
xor U9650 (N_9650,N_9529,N_9408);
and U9651 (N_9651,N_9461,N_9415);
and U9652 (N_9652,N_9508,N_9505);
or U9653 (N_9653,N_9526,N_9438);
and U9654 (N_9654,N_9483,N_9480);
nand U9655 (N_9655,N_9537,N_9551);
and U9656 (N_9656,N_9425,N_9588);
nand U9657 (N_9657,N_9497,N_9569);
and U9658 (N_9658,N_9410,N_9477);
nor U9659 (N_9659,N_9540,N_9528);
or U9660 (N_9660,N_9520,N_9517);
nand U9661 (N_9661,N_9445,N_9472);
nand U9662 (N_9662,N_9536,N_9404);
nor U9663 (N_9663,N_9514,N_9487);
nor U9664 (N_9664,N_9544,N_9420);
nor U9665 (N_9665,N_9564,N_9440);
or U9666 (N_9666,N_9595,N_9534);
or U9667 (N_9667,N_9401,N_9500);
and U9668 (N_9668,N_9436,N_9546);
or U9669 (N_9669,N_9431,N_9563);
nor U9670 (N_9670,N_9571,N_9486);
nor U9671 (N_9671,N_9482,N_9412);
xnor U9672 (N_9672,N_9580,N_9419);
nor U9673 (N_9673,N_9464,N_9510);
nor U9674 (N_9674,N_9579,N_9407);
nand U9675 (N_9675,N_9433,N_9495);
nor U9676 (N_9676,N_9502,N_9490);
and U9677 (N_9677,N_9503,N_9411);
nor U9678 (N_9678,N_9493,N_9527);
nor U9679 (N_9679,N_9456,N_9545);
or U9680 (N_9680,N_9481,N_9469);
xnor U9681 (N_9681,N_9400,N_9597);
xnor U9682 (N_9682,N_9437,N_9542);
nor U9683 (N_9683,N_9559,N_9507);
nor U9684 (N_9684,N_9473,N_9494);
or U9685 (N_9685,N_9518,N_9451);
xnor U9686 (N_9686,N_9459,N_9471);
nor U9687 (N_9687,N_9492,N_9531);
xnor U9688 (N_9688,N_9573,N_9598);
or U9689 (N_9689,N_9466,N_9460);
and U9690 (N_9690,N_9458,N_9594);
nand U9691 (N_9691,N_9592,N_9591);
or U9692 (N_9692,N_9552,N_9558);
nor U9693 (N_9693,N_9434,N_9576);
or U9694 (N_9694,N_9538,N_9468);
nand U9695 (N_9695,N_9568,N_9446);
nand U9696 (N_9696,N_9575,N_9593);
xnor U9697 (N_9697,N_9422,N_9585);
or U9698 (N_9698,N_9488,N_9476);
nand U9699 (N_9699,N_9430,N_9556);
or U9700 (N_9700,N_9560,N_9431);
or U9701 (N_9701,N_9440,N_9590);
and U9702 (N_9702,N_9542,N_9573);
nand U9703 (N_9703,N_9568,N_9545);
or U9704 (N_9704,N_9584,N_9570);
nor U9705 (N_9705,N_9522,N_9474);
nor U9706 (N_9706,N_9566,N_9560);
nand U9707 (N_9707,N_9509,N_9463);
and U9708 (N_9708,N_9561,N_9540);
and U9709 (N_9709,N_9402,N_9491);
nand U9710 (N_9710,N_9509,N_9599);
nor U9711 (N_9711,N_9580,N_9505);
nand U9712 (N_9712,N_9531,N_9514);
nand U9713 (N_9713,N_9564,N_9538);
nand U9714 (N_9714,N_9567,N_9486);
and U9715 (N_9715,N_9523,N_9406);
or U9716 (N_9716,N_9579,N_9483);
xor U9717 (N_9717,N_9410,N_9574);
xor U9718 (N_9718,N_9523,N_9594);
or U9719 (N_9719,N_9567,N_9598);
xor U9720 (N_9720,N_9576,N_9513);
and U9721 (N_9721,N_9565,N_9511);
xnor U9722 (N_9722,N_9467,N_9569);
xnor U9723 (N_9723,N_9414,N_9493);
and U9724 (N_9724,N_9577,N_9598);
xnor U9725 (N_9725,N_9462,N_9448);
xor U9726 (N_9726,N_9523,N_9542);
nand U9727 (N_9727,N_9413,N_9428);
or U9728 (N_9728,N_9419,N_9476);
nand U9729 (N_9729,N_9568,N_9474);
or U9730 (N_9730,N_9474,N_9489);
nand U9731 (N_9731,N_9577,N_9424);
nand U9732 (N_9732,N_9471,N_9533);
or U9733 (N_9733,N_9463,N_9569);
and U9734 (N_9734,N_9534,N_9593);
or U9735 (N_9735,N_9553,N_9436);
nor U9736 (N_9736,N_9427,N_9504);
or U9737 (N_9737,N_9520,N_9438);
nor U9738 (N_9738,N_9421,N_9457);
xor U9739 (N_9739,N_9561,N_9468);
or U9740 (N_9740,N_9481,N_9490);
and U9741 (N_9741,N_9485,N_9419);
nor U9742 (N_9742,N_9462,N_9560);
or U9743 (N_9743,N_9573,N_9510);
and U9744 (N_9744,N_9476,N_9411);
and U9745 (N_9745,N_9534,N_9568);
nand U9746 (N_9746,N_9573,N_9562);
nand U9747 (N_9747,N_9550,N_9419);
xnor U9748 (N_9748,N_9506,N_9425);
and U9749 (N_9749,N_9570,N_9542);
nor U9750 (N_9750,N_9545,N_9439);
and U9751 (N_9751,N_9577,N_9556);
xor U9752 (N_9752,N_9562,N_9591);
or U9753 (N_9753,N_9468,N_9491);
xnor U9754 (N_9754,N_9580,N_9407);
nand U9755 (N_9755,N_9406,N_9505);
nor U9756 (N_9756,N_9512,N_9549);
and U9757 (N_9757,N_9455,N_9548);
or U9758 (N_9758,N_9550,N_9494);
and U9759 (N_9759,N_9439,N_9519);
or U9760 (N_9760,N_9527,N_9472);
and U9761 (N_9761,N_9457,N_9435);
xnor U9762 (N_9762,N_9590,N_9522);
or U9763 (N_9763,N_9448,N_9472);
nor U9764 (N_9764,N_9468,N_9536);
or U9765 (N_9765,N_9576,N_9527);
or U9766 (N_9766,N_9523,N_9463);
or U9767 (N_9767,N_9447,N_9457);
or U9768 (N_9768,N_9538,N_9482);
and U9769 (N_9769,N_9526,N_9518);
nand U9770 (N_9770,N_9519,N_9403);
xor U9771 (N_9771,N_9499,N_9510);
xnor U9772 (N_9772,N_9569,N_9523);
or U9773 (N_9773,N_9500,N_9580);
nor U9774 (N_9774,N_9415,N_9474);
xnor U9775 (N_9775,N_9587,N_9557);
nand U9776 (N_9776,N_9547,N_9432);
nand U9777 (N_9777,N_9520,N_9453);
and U9778 (N_9778,N_9572,N_9471);
nor U9779 (N_9779,N_9494,N_9507);
nand U9780 (N_9780,N_9587,N_9458);
xor U9781 (N_9781,N_9425,N_9414);
nor U9782 (N_9782,N_9560,N_9559);
nand U9783 (N_9783,N_9401,N_9529);
nand U9784 (N_9784,N_9513,N_9430);
and U9785 (N_9785,N_9529,N_9426);
or U9786 (N_9786,N_9416,N_9532);
or U9787 (N_9787,N_9530,N_9461);
xnor U9788 (N_9788,N_9464,N_9552);
nor U9789 (N_9789,N_9452,N_9542);
nand U9790 (N_9790,N_9411,N_9541);
nor U9791 (N_9791,N_9535,N_9564);
xnor U9792 (N_9792,N_9460,N_9453);
xnor U9793 (N_9793,N_9501,N_9507);
nor U9794 (N_9794,N_9519,N_9443);
nor U9795 (N_9795,N_9422,N_9430);
nor U9796 (N_9796,N_9599,N_9496);
or U9797 (N_9797,N_9559,N_9575);
nand U9798 (N_9798,N_9517,N_9505);
nand U9799 (N_9799,N_9562,N_9592);
and U9800 (N_9800,N_9731,N_9717);
xor U9801 (N_9801,N_9781,N_9658);
and U9802 (N_9802,N_9651,N_9693);
or U9803 (N_9803,N_9618,N_9786);
and U9804 (N_9804,N_9615,N_9621);
xor U9805 (N_9805,N_9691,N_9637);
nor U9806 (N_9806,N_9770,N_9753);
and U9807 (N_9807,N_9733,N_9650);
or U9808 (N_9808,N_9616,N_9775);
and U9809 (N_9809,N_9631,N_9799);
nand U9810 (N_9810,N_9788,N_9738);
and U9811 (N_9811,N_9632,N_9679);
and U9812 (N_9812,N_9715,N_9719);
or U9813 (N_9813,N_9602,N_9707);
nor U9814 (N_9814,N_9692,N_9699);
or U9815 (N_9815,N_9674,N_9669);
nor U9816 (N_9816,N_9702,N_9736);
nor U9817 (N_9817,N_9667,N_9626);
or U9818 (N_9818,N_9711,N_9617);
xor U9819 (N_9819,N_9682,N_9760);
xnor U9820 (N_9820,N_9628,N_9742);
xor U9821 (N_9821,N_9722,N_9785);
xnor U9822 (N_9822,N_9782,N_9609);
nand U9823 (N_9823,N_9641,N_9622);
xor U9824 (N_9824,N_9758,N_9624);
nand U9825 (N_9825,N_9751,N_9789);
and U9826 (N_9826,N_9744,N_9735);
or U9827 (N_9827,N_9757,N_9745);
nor U9828 (N_9828,N_9734,N_9779);
xnor U9829 (N_9829,N_9625,N_9749);
or U9830 (N_9830,N_9647,N_9766);
xnor U9831 (N_9831,N_9752,N_9797);
nand U9832 (N_9832,N_9700,N_9664);
nand U9833 (N_9833,N_9683,N_9652);
nand U9834 (N_9834,N_9794,N_9644);
xnor U9835 (N_9835,N_9764,N_9776);
xnor U9836 (N_9836,N_9703,N_9605);
nor U9837 (N_9837,N_9608,N_9676);
xor U9838 (N_9838,N_9748,N_9726);
and U9839 (N_9839,N_9677,N_9623);
and U9840 (N_9840,N_9740,N_9694);
nor U9841 (N_9841,N_9607,N_9772);
nor U9842 (N_9842,N_9653,N_9680);
and U9843 (N_9843,N_9675,N_9762);
nand U9844 (N_9844,N_9633,N_9604);
or U9845 (N_9845,N_9769,N_9732);
or U9846 (N_9846,N_9755,N_9661);
and U9847 (N_9847,N_9643,N_9619);
or U9848 (N_9848,N_9787,N_9737);
nand U9849 (N_9849,N_9662,N_9646);
xor U9850 (N_9850,N_9730,N_9750);
or U9851 (N_9851,N_9690,N_9642);
xnor U9852 (N_9852,N_9796,N_9656);
nor U9853 (N_9853,N_9689,N_9771);
xnor U9854 (N_9854,N_9712,N_9721);
and U9855 (N_9855,N_9672,N_9710);
and U9856 (N_9856,N_9635,N_9739);
nand U9857 (N_9857,N_9670,N_9610);
and U9858 (N_9858,N_9640,N_9698);
and U9859 (N_9859,N_9747,N_9791);
nand U9860 (N_9860,N_9724,N_9620);
and U9861 (N_9861,N_9657,N_9774);
or U9862 (N_9862,N_9684,N_9614);
xor U9863 (N_9863,N_9767,N_9720);
or U9864 (N_9864,N_9629,N_9636);
and U9865 (N_9865,N_9665,N_9685);
xor U9866 (N_9866,N_9686,N_9798);
nand U9867 (N_9867,N_9654,N_9612);
xnor U9868 (N_9868,N_9759,N_9696);
or U9869 (N_9869,N_9663,N_9648);
nand U9870 (N_9870,N_9687,N_9761);
or U9871 (N_9871,N_9655,N_9728);
nand U9872 (N_9872,N_9613,N_9792);
and U9873 (N_9873,N_9743,N_9783);
nand U9874 (N_9874,N_9697,N_9713);
or U9875 (N_9875,N_9709,N_9630);
and U9876 (N_9876,N_9754,N_9671);
nor U9877 (N_9877,N_9688,N_9704);
or U9878 (N_9878,N_9706,N_9727);
xnor U9879 (N_9879,N_9777,N_9701);
nand U9880 (N_9880,N_9780,N_9705);
and U9881 (N_9881,N_9793,N_9600);
nand U9882 (N_9882,N_9768,N_9666);
nor U9883 (N_9883,N_9634,N_9638);
and U9884 (N_9884,N_9795,N_9659);
nand U9885 (N_9885,N_9606,N_9660);
nand U9886 (N_9886,N_9765,N_9601);
nand U9887 (N_9887,N_9763,N_9741);
or U9888 (N_9888,N_9611,N_9678);
xnor U9889 (N_9889,N_9746,N_9708);
nor U9890 (N_9890,N_9716,N_9695);
nand U9891 (N_9891,N_9627,N_9756);
nor U9892 (N_9892,N_9723,N_9645);
nand U9893 (N_9893,N_9673,N_9773);
nor U9894 (N_9894,N_9714,N_9681);
or U9895 (N_9895,N_9784,N_9603);
nand U9896 (N_9896,N_9639,N_9778);
nand U9897 (N_9897,N_9668,N_9729);
and U9898 (N_9898,N_9725,N_9649);
or U9899 (N_9899,N_9718,N_9790);
nand U9900 (N_9900,N_9785,N_9659);
or U9901 (N_9901,N_9670,N_9640);
nor U9902 (N_9902,N_9716,N_9647);
nand U9903 (N_9903,N_9738,N_9613);
xor U9904 (N_9904,N_9732,N_9630);
and U9905 (N_9905,N_9675,N_9701);
nand U9906 (N_9906,N_9765,N_9689);
nand U9907 (N_9907,N_9662,N_9751);
and U9908 (N_9908,N_9606,N_9629);
nand U9909 (N_9909,N_9730,N_9746);
or U9910 (N_9910,N_9657,N_9641);
or U9911 (N_9911,N_9684,N_9680);
nor U9912 (N_9912,N_9737,N_9740);
or U9913 (N_9913,N_9700,N_9639);
or U9914 (N_9914,N_9798,N_9680);
or U9915 (N_9915,N_9625,N_9615);
or U9916 (N_9916,N_9620,N_9672);
nor U9917 (N_9917,N_9786,N_9604);
or U9918 (N_9918,N_9735,N_9725);
and U9919 (N_9919,N_9741,N_9743);
nor U9920 (N_9920,N_9732,N_9738);
nand U9921 (N_9921,N_9745,N_9683);
nor U9922 (N_9922,N_9726,N_9693);
xor U9923 (N_9923,N_9798,N_9762);
nand U9924 (N_9924,N_9785,N_9620);
xor U9925 (N_9925,N_9678,N_9626);
xnor U9926 (N_9926,N_9663,N_9794);
nand U9927 (N_9927,N_9632,N_9691);
or U9928 (N_9928,N_9759,N_9614);
xor U9929 (N_9929,N_9725,N_9774);
nand U9930 (N_9930,N_9648,N_9769);
xnor U9931 (N_9931,N_9691,N_9720);
and U9932 (N_9932,N_9710,N_9659);
xor U9933 (N_9933,N_9633,N_9602);
and U9934 (N_9934,N_9634,N_9651);
and U9935 (N_9935,N_9719,N_9647);
nand U9936 (N_9936,N_9758,N_9652);
or U9937 (N_9937,N_9686,N_9613);
nand U9938 (N_9938,N_9676,N_9726);
xnor U9939 (N_9939,N_9707,N_9662);
nor U9940 (N_9940,N_9633,N_9724);
nor U9941 (N_9941,N_9601,N_9643);
or U9942 (N_9942,N_9625,N_9702);
xor U9943 (N_9943,N_9698,N_9603);
or U9944 (N_9944,N_9799,N_9796);
and U9945 (N_9945,N_9610,N_9739);
nand U9946 (N_9946,N_9646,N_9609);
nor U9947 (N_9947,N_9620,N_9742);
nand U9948 (N_9948,N_9623,N_9690);
nand U9949 (N_9949,N_9770,N_9744);
xnor U9950 (N_9950,N_9772,N_9674);
nand U9951 (N_9951,N_9724,N_9723);
xor U9952 (N_9952,N_9613,N_9799);
and U9953 (N_9953,N_9654,N_9653);
or U9954 (N_9954,N_9644,N_9625);
nand U9955 (N_9955,N_9610,N_9669);
nor U9956 (N_9956,N_9689,N_9672);
or U9957 (N_9957,N_9756,N_9658);
or U9958 (N_9958,N_9615,N_9750);
or U9959 (N_9959,N_9766,N_9785);
xnor U9960 (N_9960,N_9666,N_9788);
or U9961 (N_9961,N_9767,N_9654);
or U9962 (N_9962,N_9700,N_9638);
xnor U9963 (N_9963,N_9739,N_9770);
and U9964 (N_9964,N_9613,N_9781);
xnor U9965 (N_9965,N_9609,N_9776);
nand U9966 (N_9966,N_9619,N_9633);
nand U9967 (N_9967,N_9757,N_9617);
and U9968 (N_9968,N_9772,N_9636);
and U9969 (N_9969,N_9723,N_9615);
and U9970 (N_9970,N_9730,N_9743);
nand U9971 (N_9971,N_9631,N_9694);
xor U9972 (N_9972,N_9690,N_9689);
nand U9973 (N_9973,N_9773,N_9769);
or U9974 (N_9974,N_9718,N_9617);
xor U9975 (N_9975,N_9750,N_9786);
xor U9976 (N_9976,N_9606,N_9600);
nor U9977 (N_9977,N_9672,N_9687);
and U9978 (N_9978,N_9789,N_9686);
nand U9979 (N_9979,N_9653,N_9632);
or U9980 (N_9980,N_9696,N_9765);
and U9981 (N_9981,N_9659,N_9766);
and U9982 (N_9982,N_9747,N_9662);
nand U9983 (N_9983,N_9649,N_9745);
or U9984 (N_9984,N_9738,N_9662);
and U9985 (N_9985,N_9763,N_9629);
xnor U9986 (N_9986,N_9720,N_9615);
nand U9987 (N_9987,N_9696,N_9723);
nor U9988 (N_9988,N_9737,N_9765);
nand U9989 (N_9989,N_9626,N_9696);
or U9990 (N_9990,N_9784,N_9723);
xor U9991 (N_9991,N_9608,N_9619);
nand U9992 (N_9992,N_9742,N_9606);
nand U9993 (N_9993,N_9770,N_9703);
xnor U9994 (N_9994,N_9633,N_9786);
and U9995 (N_9995,N_9755,N_9758);
xor U9996 (N_9996,N_9740,N_9771);
nand U9997 (N_9997,N_9626,N_9729);
xnor U9998 (N_9998,N_9609,N_9603);
nand U9999 (N_9999,N_9650,N_9738);
nor UO_0 (O_0,N_9983,N_9973);
nor UO_1 (O_1,N_9803,N_9818);
and UO_2 (O_2,N_9958,N_9856);
xnor UO_3 (O_3,N_9890,N_9981);
and UO_4 (O_4,N_9894,N_9868);
and UO_5 (O_5,N_9881,N_9921);
or UO_6 (O_6,N_9929,N_9987);
nor UO_7 (O_7,N_9845,N_9916);
xnor UO_8 (O_8,N_9949,N_9988);
and UO_9 (O_9,N_9807,N_9804);
or UO_10 (O_10,N_9972,N_9846);
nand UO_11 (O_11,N_9909,N_9935);
xnor UO_12 (O_12,N_9933,N_9898);
xor UO_13 (O_13,N_9848,N_9998);
nand UO_14 (O_14,N_9858,N_9932);
xnor UO_15 (O_15,N_9866,N_9951);
nor UO_16 (O_16,N_9892,N_9820);
or UO_17 (O_17,N_9993,N_9838);
xnor UO_18 (O_18,N_9809,N_9940);
nand UO_19 (O_19,N_9867,N_9930);
xor UO_20 (O_20,N_9976,N_9912);
or UO_21 (O_21,N_9974,N_9851);
xor UO_22 (O_22,N_9960,N_9947);
nand UO_23 (O_23,N_9819,N_9835);
nor UO_24 (O_24,N_9842,N_9876);
xor UO_25 (O_25,N_9986,N_9982);
and UO_26 (O_26,N_9833,N_9839);
nand UO_27 (O_27,N_9887,N_9824);
and UO_28 (O_28,N_9882,N_9834);
or UO_29 (O_29,N_9891,N_9936);
xor UO_30 (O_30,N_9923,N_9830);
nor UO_31 (O_31,N_9917,N_9939);
and UO_32 (O_32,N_9897,N_9995);
nand UO_33 (O_33,N_9865,N_9875);
nand UO_34 (O_34,N_9965,N_9924);
or UO_35 (O_35,N_9963,N_9991);
or UO_36 (O_36,N_9925,N_9964);
nor UO_37 (O_37,N_9857,N_9966);
xnor UO_38 (O_38,N_9879,N_9931);
and UO_39 (O_39,N_9806,N_9802);
xnor UO_40 (O_40,N_9859,N_9905);
nor UO_41 (O_41,N_9808,N_9910);
nand UO_42 (O_42,N_9907,N_9941);
and UO_43 (O_43,N_9888,N_9978);
nand UO_44 (O_44,N_9840,N_9927);
xor UO_45 (O_45,N_9837,N_9847);
nand UO_46 (O_46,N_9979,N_9853);
and UO_47 (O_47,N_9895,N_9920);
and UO_48 (O_48,N_9985,N_9970);
xor UO_49 (O_49,N_9952,N_9919);
or UO_50 (O_50,N_9946,N_9943);
nor UO_51 (O_51,N_9823,N_9861);
or UO_52 (O_52,N_9942,N_9938);
xor UO_53 (O_53,N_9903,N_9800);
nor UO_54 (O_54,N_9953,N_9955);
or UO_55 (O_55,N_9937,N_9997);
and UO_56 (O_56,N_9954,N_9854);
nor UO_57 (O_57,N_9980,N_9827);
nand UO_58 (O_58,N_9880,N_9967);
xor UO_59 (O_59,N_9829,N_9873);
nand UO_60 (O_60,N_9814,N_9852);
nor UO_61 (O_61,N_9922,N_9812);
xnor UO_62 (O_62,N_9999,N_9908);
nand UO_63 (O_63,N_9913,N_9825);
or UO_64 (O_64,N_9815,N_9878);
nand UO_65 (O_65,N_9817,N_9844);
nand UO_66 (O_66,N_9956,N_9828);
nand UO_67 (O_67,N_9885,N_9860);
and UO_68 (O_68,N_9864,N_9926);
nand UO_69 (O_69,N_9886,N_9928);
or UO_70 (O_70,N_9869,N_9944);
nor UO_71 (O_71,N_9850,N_9957);
nor UO_72 (O_72,N_9994,N_9893);
and UO_73 (O_73,N_9961,N_9906);
nand UO_74 (O_74,N_9801,N_9901);
and UO_75 (O_75,N_9989,N_9889);
nand UO_76 (O_76,N_9900,N_9902);
nor UO_77 (O_77,N_9948,N_9877);
nor UO_78 (O_78,N_9826,N_9883);
nor UO_79 (O_79,N_9816,N_9841);
xnor UO_80 (O_80,N_9874,N_9805);
nand UO_81 (O_81,N_9813,N_9911);
nand UO_82 (O_82,N_9984,N_9884);
or UO_83 (O_83,N_9992,N_9962);
or UO_84 (O_84,N_9870,N_9996);
xor UO_85 (O_85,N_9862,N_9896);
nand UO_86 (O_86,N_9871,N_9855);
and UO_87 (O_87,N_9959,N_9918);
nor UO_88 (O_88,N_9811,N_9945);
or UO_89 (O_89,N_9904,N_9899);
xor UO_90 (O_90,N_9990,N_9977);
and UO_91 (O_91,N_9975,N_9968);
or UO_92 (O_92,N_9969,N_9832);
xor UO_93 (O_93,N_9821,N_9810);
or UO_94 (O_94,N_9934,N_9914);
nor UO_95 (O_95,N_9950,N_9849);
nand UO_96 (O_96,N_9872,N_9822);
and UO_97 (O_97,N_9843,N_9863);
and UO_98 (O_98,N_9831,N_9915);
xnor UO_99 (O_99,N_9836,N_9971);
and UO_100 (O_100,N_9816,N_9952);
nand UO_101 (O_101,N_9896,N_9969);
nand UO_102 (O_102,N_9992,N_9974);
nor UO_103 (O_103,N_9922,N_9953);
xor UO_104 (O_104,N_9808,N_9923);
xor UO_105 (O_105,N_9882,N_9924);
xor UO_106 (O_106,N_9911,N_9898);
or UO_107 (O_107,N_9914,N_9842);
and UO_108 (O_108,N_9863,N_9900);
and UO_109 (O_109,N_9984,N_9976);
and UO_110 (O_110,N_9918,N_9971);
nand UO_111 (O_111,N_9802,N_9976);
nand UO_112 (O_112,N_9921,N_9886);
or UO_113 (O_113,N_9915,N_9982);
nor UO_114 (O_114,N_9939,N_9877);
nand UO_115 (O_115,N_9838,N_9816);
or UO_116 (O_116,N_9831,N_9900);
nor UO_117 (O_117,N_9826,N_9967);
nor UO_118 (O_118,N_9893,N_9828);
nor UO_119 (O_119,N_9812,N_9969);
or UO_120 (O_120,N_9881,N_9960);
and UO_121 (O_121,N_9805,N_9922);
nand UO_122 (O_122,N_9951,N_9825);
and UO_123 (O_123,N_9950,N_9813);
nand UO_124 (O_124,N_9824,N_9901);
nor UO_125 (O_125,N_9917,N_9991);
nor UO_126 (O_126,N_9940,N_9929);
nand UO_127 (O_127,N_9881,N_9937);
nand UO_128 (O_128,N_9955,N_9885);
xor UO_129 (O_129,N_9830,N_9818);
xnor UO_130 (O_130,N_9930,N_9893);
or UO_131 (O_131,N_9917,N_9813);
nor UO_132 (O_132,N_9846,N_9975);
and UO_133 (O_133,N_9970,N_9942);
xnor UO_134 (O_134,N_9915,N_9976);
xor UO_135 (O_135,N_9854,N_9925);
or UO_136 (O_136,N_9985,N_9989);
nand UO_137 (O_137,N_9814,N_9971);
nor UO_138 (O_138,N_9936,N_9802);
or UO_139 (O_139,N_9932,N_9951);
or UO_140 (O_140,N_9809,N_9842);
or UO_141 (O_141,N_9961,N_9883);
nand UO_142 (O_142,N_9810,N_9867);
or UO_143 (O_143,N_9831,N_9824);
and UO_144 (O_144,N_9919,N_9880);
and UO_145 (O_145,N_9800,N_9955);
xnor UO_146 (O_146,N_9981,N_9937);
nor UO_147 (O_147,N_9986,N_9945);
and UO_148 (O_148,N_9886,N_9822);
or UO_149 (O_149,N_9896,N_9876);
or UO_150 (O_150,N_9885,N_9910);
and UO_151 (O_151,N_9825,N_9887);
xor UO_152 (O_152,N_9922,N_9959);
or UO_153 (O_153,N_9919,N_9971);
and UO_154 (O_154,N_9987,N_9936);
nor UO_155 (O_155,N_9967,N_9927);
xnor UO_156 (O_156,N_9804,N_9834);
nand UO_157 (O_157,N_9893,N_9865);
xor UO_158 (O_158,N_9915,N_9854);
and UO_159 (O_159,N_9988,N_9946);
and UO_160 (O_160,N_9851,N_9815);
or UO_161 (O_161,N_9979,N_9850);
nor UO_162 (O_162,N_9966,N_9914);
nor UO_163 (O_163,N_9808,N_9940);
xnor UO_164 (O_164,N_9893,N_9919);
or UO_165 (O_165,N_9981,N_9809);
and UO_166 (O_166,N_9982,N_9946);
and UO_167 (O_167,N_9814,N_9863);
nand UO_168 (O_168,N_9958,N_9996);
xnor UO_169 (O_169,N_9959,N_9998);
xor UO_170 (O_170,N_9899,N_9818);
nor UO_171 (O_171,N_9816,N_9947);
nor UO_172 (O_172,N_9991,N_9932);
nor UO_173 (O_173,N_9850,N_9965);
or UO_174 (O_174,N_9895,N_9937);
nand UO_175 (O_175,N_9867,N_9821);
xor UO_176 (O_176,N_9952,N_9832);
or UO_177 (O_177,N_9918,N_9938);
or UO_178 (O_178,N_9999,N_9936);
and UO_179 (O_179,N_9807,N_9836);
and UO_180 (O_180,N_9944,N_9912);
and UO_181 (O_181,N_9826,N_9878);
xor UO_182 (O_182,N_9887,N_9910);
and UO_183 (O_183,N_9935,N_9831);
nand UO_184 (O_184,N_9886,N_9936);
nor UO_185 (O_185,N_9852,N_9843);
and UO_186 (O_186,N_9815,N_9841);
nor UO_187 (O_187,N_9815,N_9949);
xnor UO_188 (O_188,N_9989,N_9966);
or UO_189 (O_189,N_9993,N_9986);
nand UO_190 (O_190,N_9865,N_9855);
or UO_191 (O_191,N_9999,N_9869);
or UO_192 (O_192,N_9811,N_9902);
xnor UO_193 (O_193,N_9993,N_9840);
nor UO_194 (O_194,N_9805,N_9873);
nor UO_195 (O_195,N_9843,N_9930);
nor UO_196 (O_196,N_9856,N_9894);
nand UO_197 (O_197,N_9955,N_9951);
nor UO_198 (O_198,N_9835,N_9905);
nand UO_199 (O_199,N_9912,N_9818);
nor UO_200 (O_200,N_9971,N_9808);
nor UO_201 (O_201,N_9955,N_9946);
xor UO_202 (O_202,N_9868,N_9955);
or UO_203 (O_203,N_9854,N_9881);
nor UO_204 (O_204,N_9933,N_9866);
and UO_205 (O_205,N_9915,N_9939);
or UO_206 (O_206,N_9830,N_9899);
or UO_207 (O_207,N_9962,N_9968);
and UO_208 (O_208,N_9804,N_9946);
or UO_209 (O_209,N_9947,N_9954);
xor UO_210 (O_210,N_9922,N_9813);
nand UO_211 (O_211,N_9837,N_9846);
xnor UO_212 (O_212,N_9976,N_9853);
or UO_213 (O_213,N_9921,N_9930);
and UO_214 (O_214,N_9802,N_9998);
and UO_215 (O_215,N_9823,N_9863);
nor UO_216 (O_216,N_9994,N_9864);
and UO_217 (O_217,N_9810,N_9877);
or UO_218 (O_218,N_9882,N_9966);
xnor UO_219 (O_219,N_9892,N_9913);
and UO_220 (O_220,N_9837,N_9884);
xnor UO_221 (O_221,N_9870,N_9893);
or UO_222 (O_222,N_9937,N_9955);
nor UO_223 (O_223,N_9849,N_9952);
nor UO_224 (O_224,N_9836,N_9887);
and UO_225 (O_225,N_9977,N_9916);
xnor UO_226 (O_226,N_9906,N_9803);
and UO_227 (O_227,N_9924,N_9853);
or UO_228 (O_228,N_9846,N_9923);
and UO_229 (O_229,N_9926,N_9828);
nor UO_230 (O_230,N_9920,N_9964);
xnor UO_231 (O_231,N_9836,N_9838);
xnor UO_232 (O_232,N_9894,N_9812);
and UO_233 (O_233,N_9966,N_9851);
and UO_234 (O_234,N_9969,N_9831);
nand UO_235 (O_235,N_9921,N_9975);
nand UO_236 (O_236,N_9912,N_9903);
nor UO_237 (O_237,N_9893,N_9846);
nor UO_238 (O_238,N_9850,N_9975);
nand UO_239 (O_239,N_9911,N_9844);
nor UO_240 (O_240,N_9816,N_9802);
nor UO_241 (O_241,N_9899,N_9896);
nand UO_242 (O_242,N_9915,N_9957);
or UO_243 (O_243,N_9827,N_9997);
nor UO_244 (O_244,N_9900,N_9829);
nor UO_245 (O_245,N_9832,N_9810);
and UO_246 (O_246,N_9909,N_9913);
or UO_247 (O_247,N_9872,N_9953);
and UO_248 (O_248,N_9800,N_9938);
nand UO_249 (O_249,N_9871,N_9996);
and UO_250 (O_250,N_9938,N_9813);
or UO_251 (O_251,N_9911,N_9853);
or UO_252 (O_252,N_9865,N_9832);
nand UO_253 (O_253,N_9819,N_9838);
xnor UO_254 (O_254,N_9993,N_9876);
nand UO_255 (O_255,N_9922,N_9820);
xor UO_256 (O_256,N_9807,N_9922);
or UO_257 (O_257,N_9847,N_9809);
and UO_258 (O_258,N_9814,N_9809);
xnor UO_259 (O_259,N_9819,N_9890);
and UO_260 (O_260,N_9952,N_9833);
or UO_261 (O_261,N_9963,N_9954);
xor UO_262 (O_262,N_9961,N_9867);
and UO_263 (O_263,N_9977,N_9863);
nor UO_264 (O_264,N_9924,N_9963);
xor UO_265 (O_265,N_9910,N_9975);
or UO_266 (O_266,N_9870,N_9964);
and UO_267 (O_267,N_9939,N_9874);
and UO_268 (O_268,N_9815,N_9916);
nor UO_269 (O_269,N_9848,N_9999);
and UO_270 (O_270,N_9809,N_9961);
or UO_271 (O_271,N_9963,N_9907);
nand UO_272 (O_272,N_9934,N_9805);
or UO_273 (O_273,N_9914,N_9999);
or UO_274 (O_274,N_9815,N_9933);
and UO_275 (O_275,N_9938,N_9835);
and UO_276 (O_276,N_9903,N_9923);
nor UO_277 (O_277,N_9947,N_9990);
nor UO_278 (O_278,N_9878,N_9911);
and UO_279 (O_279,N_9863,N_9869);
or UO_280 (O_280,N_9947,N_9900);
or UO_281 (O_281,N_9886,N_9830);
nand UO_282 (O_282,N_9894,N_9924);
or UO_283 (O_283,N_9847,N_9953);
xnor UO_284 (O_284,N_9999,N_9958);
or UO_285 (O_285,N_9966,N_9968);
and UO_286 (O_286,N_9838,N_9989);
nand UO_287 (O_287,N_9975,N_9885);
and UO_288 (O_288,N_9824,N_9817);
or UO_289 (O_289,N_9804,N_9896);
xnor UO_290 (O_290,N_9943,N_9884);
nand UO_291 (O_291,N_9864,N_9825);
or UO_292 (O_292,N_9887,N_9847);
nand UO_293 (O_293,N_9882,N_9954);
and UO_294 (O_294,N_9811,N_9938);
and UO_295 (O_295,N_9817,N_9948);
nor UO_296 (O_296,N_9862,N_9895);
or UO_297 (O_297,N_9832,N_9937);
xor UO_298 (O_298,N_9937,N_9943);
nand UO_299 (O_299,N_9935,N_9830);
or UO_300 (O_300,N_9999,N_9873);
xor UO_301 (O_301,N_9923,N_9912);
or UO_302 (O_302,N_9967,N_9909);
nor UO_303 (O_303,N_9860,N_9959);
and UO_304 (O_304,N_9912,N_9859);
or UO_305 (O_305,N_9939,N_9857);
or UO_306 (O_306,N_9875,N_9982);
nor UO_307 (O_307,N_9811,N_9971);
and UO_308 (O_308,N_9928,N_9822);
nand UO_309 (O_309,N_9835,N_9908);
nand UO_310 (O_310,N_9969,N_9943);
xnor UO_311 (O_311,N_9927,N_9834);
nor UO_312 (O_312,N_9957,N_9996);
nand UO_313 (O_313,N_9902,N_9860);
xnor UO_314 (O_314,N_9968,N_9835);
nand UO_315 (O_315,N_9974,N_9929);
xor UO_316 (O_316,N_9828,N_9879);
xnor UO_317 (O_317,N_9886,N_9904);
nor UO_318 (O_318,N_9813,N_9914);
or UO_319 (O_319,N_9832,N_9863);
or UO_320 (O_320,N_9839,N_9853);
and UO_321 (O_321,N_9948,N_9897);
xor UO_322 (O_322,N_9826,N_9986);
xnor UO_323 (O_323,N_9957,N_9968);
xnor UO_324 (O_324,N_9871,N_9864);
and UO_325 (O_325,N_9914,N_9824);
and UO_326 (O_326,N_9975,N_9838);
or UO_327 (O_327,N_9864,N_9989);
and UO_328 (O_328,N_9829,N_9941);
xor UO_329 (O_329,N_9990,N_9937);
and UO_330 (O_330,N_9852,N_9850);
and UO_331 (O_331,N_9936,N_9975);
nor UO_332 (O_332,N_9937,N_9872);
xor UO_333 (O_333,N_9901,N_9984);
xnor UO_334 (O_334,N_9925,N_9932);
nand UO_335 (O_335,N_9804,N_9875);
nand UO_336 (O_336,N_9908,N_9923);
and UO_337 (O_337,N_9822,N_9997);
or UO_338 (O_338,N_9840,N_9855);
nor UO_339 (O_339,N_9806,N_9902);
xor UO_340 (O_340,N_9976,N_9834);
nor UO_341 (O_341,N_9826,N_9872);
nand UO_342 (O_342,N_9896,N_9831);
nor UO_343 (O_343,N_9845,N_9859);
or UO_344 (O_344,N_9893,N_9998);
nor UO_345 (O_345,N_9899,N_9961);
nor UO_346 (O_346,N_9870,N_9828);
or UO_347 (O_347,N_9806,N_9931);
or UO_348 (O_348,N_9838,N_9991);
and UO_349 (O_349,N_9943,N_9914);
xnor UO_350 (O_350,N_9920,N_9860);
and UO_351 (O_351,N_9957,N_9994);
and UO_352 (O_352,N_9940,N_9903);
xor UO_353 (O_353,N_9927,N_9916);
xnor UO_354 (O_354,N_9808,N_9920);
xor UO_355 (O_355,N_9865,N_9971);
xnor UO_356 (O_356,N_9971,N_9824);
xor UO_357 (O_357,N_9846,N_9892);
xnor UO_358 (O_358,N_9894,N_9840);
or UO_359 (O_359,N_9981,N_9805);
or UO_360 (O_360,N_9935,N_9938);
and UO_361 (O_361,N_9973,N_9886);
or UO_362 (O_362,N_9852,N_9864);
xnor UO_363 (O_363,N_9931,N_9973);
xor UO_364 (O_364,N_9830,N_9993);
nand UO_365 (O_365,N_9920,N_9811);
or UO_366 (O_366,N_9838,N_9885);
nand UO_367 (O_367,N_9996,N_9844);
nor UO_368 (O_368,N_9819,N_9988);
nand UO_369 (O_369,N_9894,N_9861);
and UO_370 (O_370,N_9961,N_9870);
or UO_371 (O_371,N_9816,N_9982);
and UO_372 (O_372,N_9982,N_9829);
xor UO_373 (O_373,N_9880,N_9861);
and UO_374 (O_374,N_9997,N_9992);
or UO_375 (O_375,N_9892,N_9938);
or UO_376 (O_376,N_9848,N_9850);
nand UO_377 (O_377,N_9944,N_9844);
and UO_378 (O_378,N_9977,N_9972);
xnor UO_379 (O_379,N_9983,N_9815);
nand UO_380 (O_380,N_9998,N_9929);
or UO_381 (O_381,N_9872,N_9844);
nand UO_382 (O_382,N_9993,N_9952);
nand UO_383 (O_383,N_9895,N_9882);
or UO_384 (O_384,N_9905,N_9815);
or UO_385 (O_385,N_9933,N_9922);
or UO_386 (O_386,N_9963,N_9841);
or UO_387 (O_387,N_9854,N_9995);
xor UO_388 (O_388,N_9806,N_9875);
xnor UO_389 (O_389,N_9966,N_9992);
xor UO_390 (O_390,N_9893,N_9949);
xor UO_391 (O_391,N_9965,N_9804);
or UO_392 (O_392,N_9907,N_9864);
and UO_393 (O_393,N_9867,N_9831);
or UO_394 (O_394,N_9957,N_9944);
nor UO_395 (O_395,N_9807,N_9968);
xor UO_396 (O_396,N_9873,N_9855);
nor UO_397 (O_397,N_9893,N_9939);
nand UO_398 (O_398,N_9815,N_9942);
nor UO_399 (O_399,N_9813,N_9909);
and UO_400 (O_400,N_9859,N_9871);
and UO_401 (O_401,N_9886,N_9962);
and UO_402 (O_402,N_9829,N_9926);
or UO_403 (O_403,N_9949,N_9823);
or UO_404 (O_404,N_9958,N_9852);
nand UO_405 (O_405,N_9984,N_9810);
or UO_406 (O_406,N_9999,N_9820);
and UO_407 (O_407,N_9977,N_9995);
and UO_408 (O_408,N_9856,N_9919);
or UO_409 (O_409,N_9955,N_9922);
and UO_410 (O_410,N_9838,N_9861);
nand UO_411 (O_411,N_9986,N_9820);
or UO_412 (O_412,N_9840,N_9829);
nor UO_413 (O_413,N_9907,N_9967);
or UO_414 (O_414,N_9809,N_9970);
and UO_415 (O_415,N_9914,N_9951);
or UO_416 (O_416,N_9859,N_9889);
and UO_417 (O_417,N_9912,N_9918);
or UO_418 (O_418,N_9862,N_9971);
nor UO_419 (O_419,N_9948,N_9881);
xor UO_420 (O_420,N_9872,N_9885);
xor UO_421 (O_421,N_9874,N_9889);
nand UO_422 (O_422,N_9880,N_9886);
or UO_423 (O_423,N_9993,N_9818);
nor UO_424 (O_424,N_9818,N_9982);
nand UO_425 (O_425,N_9983,N_9828);
and UO_426 (O_426,N_9905,N_9959);
xnor UO_427 (O_427,N_9891,N_9914);
and UO_428 (O_428,N_9978,N_9983);
or UO_429 (O_429,N_9953,N_9981);
or UO_430 (O_430,N_9808,N_9819);
nor UO_431 (O_431,N_9936,N_9849);
or UO_432 (O_432,N_9988,N_9820);
nand UO_433 (O_433,N_9920,N_9983);
and UO_434 (O_434,N_9993,N_9965);
nor UO_435 (O_435,N_9857,N_9804);
xor UO_436 (O_436,N_9811,N_9914);
nand UO_437 (O_437,N_9847,N_9916);
xnor UO_438 (O_438,N_9950,N_9809);
nand UO_439 (O_439,N_9908,N_9910);
and UO_440 (O_440,N_9895,N_9859);
nand UO_441 (O_441,N_9972,N_9953);
and UO_442 (O_442,N_9869,N_9911);
nor UO_443 (O_443,N_9875,N_9987);
nand UO_444 (O_444,N_9868,N_9963);
or UO_445 (O_445,N_9910,N_9962);
or UO_446 (O_446,N_9840,N_9913);
xor UO_447 (O_447,N_9913,N_9823);
xor UO_448 (O_448,N_9980,N_9927);
xnor UO_449 (O_449,N_9983,N_9954);
or UO_450 (O_450,N_9951,N_9867);
nand UO_451 (O_451,N_9852,N_9938);
nand UO_452 (O_452,N_9867,N_9918);
and UO_453 (O_453,N_9839,N_9941);
nand UO_454 (O_454,N_9921,N_9899);
nor UO_455 (O_455,N_9918,N_9815);
xor UO_456 (O_456,N_9911,N_9902);
nor UO_457 (O_457,N_9838,N_9917);
nor UO_458 (O_458,N_9824,N_9990);
nand UO_459 (O_459,N_9961,N_9829);
nor UO_460 (O_460,N_9946,N_9848);
and UO_461 (O_461,N_9984,N_9939);
and UO_462 (O_462,N_9812,N_9830);
and UO_463 (O_463,N_9810,N_9895);
and UO_464 (O_464,N_9941,N_9983);
nand UO_465 (O_465,N_9964,N_9943);
and UO_466 (O_466,N_9924,N_9996);
or UO_467 (O_467,N_9893,N_9999);
nor UO_468 (O_468,N_9822,N_9863);
nor UO_469 (O_469,N_9874,N_9922);
xnor UO_470 (O_470,N_9846,N_9977);
nor UO_471 (O_471,N_9840,N_9968);
nand UO_472 (O_472,N_9944,N_9901);
nor UO_473 (O_473,N_9817,N_9892);
or UO_474 (O_474,N_9894,N_9911);
nand UO_475 (O_475,N_9907,N_9853);
nor UO_476 (O_476,N_9929,N_9970);
nor UO_477 (O_477,N_9812,N_9965);
nand UO_478 (O_478,N_9988,N_9967);
and UO_479 (O_479,N_9806,N_9935);
xnor UO_480 (O_480,N_9892,N_9907);
nand UO_481 (O_481,N_9948,N_9880);
nand UO_482 (O_482,N_9954,N_9890);
or UO_483 (O_483,N_9801,N_9963);
nand UO_484 (O_484,N_9854,N_9901);
nor UO_485 (O_485,N_9901,N_9880);
or UO_486 (O_486,N_9857,N_9955);
nand UO_487 (O_487,N_9875,N_9948);
xnor UO_488 (O_488,N_9800,N_9936);
nor UO_489 (O_489,N_9852,N_9960);
and UO_490 (O_490,N_9800,N_9912);
nand UO_491 (O_491,N_9974,N_9981);
and UO_492 (O_492,N_9834,N_9994);
nor UO_493 (O_493,N_9976,N_9993);
and UO_494 (O_494,N_9875,N_9909);
xnor UO_495 (O_495,N_9889,N_9915);
or UO_496 (O_496,N_9931,N_9943);
nor UO_497 (O_497,N_9995,N_9841);
and UO_498 (O_498,N_9997,N_9998);
nand UO_499 (O_499,N_9933,N_9830);
nand UO_500 (O_500,N_9950,N_9846);
xnor UO_501 (O_501,N_9998,N_9897);
and UO_502 (O_502,N_9810,N_9874);
xnor UO_503 (O_503,N_9981,N_9866);
nor UO_504 (O_504,N_9825,N_9982);
xor UO_505 (O_505,N_9830,N_9980);
and UO_506 (O_506,N_9921,N_9903);
and UO_507 (O_507,N_9946,N_9857);
or UO_508 (O_508,N_9996,N_9804);
nand UO_509 (O_509,N_9890,N_9885);
and UO_510 (O_510,N_9942,N_9860);
or UO_511 (O_511,N_9887,N_9976);
xor UO_512 (O_512,N_9834,N_9957);
xor UO_513 (O_513,N_9864,N_9893);
nand UO_514 (O_514,N_9851,N_9856);
and UO_515 (O_515,N_9916,N_9887);
and UO_516 (O_516,N_9949,N_9818);
nand UO_517 (O_517,N_9968,N_9852);
xor UO_518 (O_518,N_9804,N_9943);
or UO_519 (O_519,N_9975,N_9988);
or UO_520 (O_520,N_9883,N_9916);
or UO_521 (O_521,N_9998,N_9841);
xor UO_522 (O_522,N_9925,N_9852);
nand UO_523 (O_523,N_9839,N_9804);
and UO_524 (O_524,N_9828,N_9815);
or UO_525 (O_525,N_9952,N_9837);
nor UO_526 (O_526,N_9882,N_9899);
nor UO_527 (O_527,N_9819,N_9993);
and UO_528 (O_528,N_9929,N_9968);
nand UO_529 (O_529,N_9916,N_9957);
nor UO_530 (O_530,N_9929,N_9907);
xnor UO_531 (O_531,N_9816,N_9860);
nand UO_532 (O_532,N_9991,N_9802);
nor UO_533 (O_533,N_9839,N_9926);
nor UO_534 (O_534,N_9819,N_9917);
xnor UO_535 (O_535,N_9908,N_9878);
xnor UO_536 (O_536,N_9850,N_9968);
and UO_537 (O_537,N_9891,N_9803);
or UO_538 (O_538,N_9868,N_9941);
xor UO_539 (O_539,N_9961,N_9881);
or UO_540 (O_540,N_9977,N_9820);
or UO_541 (O_541,N_9892,N_9886);
nand UO_542 (O_542,N_9809,N_9821);
xnor UO_543 (O_543,N_9979,N_9975);
nand UO_544 (O_544,N_9846,N_9978);
or UO_545 (O_545,N_9816,N_9877);
nor UO_546 (O_546,N_9895,N_9994);
nor UO_547 (O_547,N_9841,N_9939);
and UO_548 (O_548,N_9945,N_9816);
nand UO_549 (O_549,N_9852,N_9984);
xor UO_550 (O_550,N_9915,N_9944);
or UO_551 (O_551,N_9880,N_9846);
and UO_552 (O_552,N_9803,N_9880);
nand UO_553 (O_553,N_9833,N_9991);
and UO_554 (O_554,N_9877,N_9805);
nand UO_555 (O_555,N_9929,N_9973);
nand UO_556 (O_556,N_9972,N_9817);
xor UO_557 (O_557,N_9811,N_9898);
or UO_558 (O_558,N_9997,N_9906);
or UO_559 (O_559,N_9805,N_9938);
xnor UO_560 (O_560,N_9824,N_9839);
and UO_561 (O_561,N_9858,N_9847);
nor UO_562 (O_562,N_9985,N_9861);
nand UO_563 (O_563,N_9820,N_9933);
xor UO_564 (O_564,N_9856,N_9885);
nor UO_565 (O_565,N_9800,N_9842);
nand UO_566 (O_566,N_9938,N_9932);
and UO_567 (O_567,N_9996,N_9893);
xor UO_568 (O_568,N_9884,N_9961);
or UO_569 (O_569,N_9833,N_9981);
xor UO_570 (O_570,N_9835,N_9838);
nor UO_571 (O_571,N_9920,N_9863);
or UO_572 (O_572,N_9825,N_9854);
and UO_573 (O_573,N_9847,N_9882);
or UO_574 (O_574,N_9842,N_9802);
nor UO_575 (O_575,N_9940,N_9892);
nand UO_576 (O_576,N_9879,N_9821);
nor UO_577 (O_577,N_9857,N_9903);
or UO_578 (O_578,N_9900,N_9852);
nand UO_579 (O_579,N_9966,N_9925);
xnor UO_580 (O_580,N_9840,N_9984);
xor UO_581 (O_581,N_9847,N_9898);
nand UO_582 (O_582,N_9920,N_9947);
nand UO_583 (O_583,N_9914,N_9817);
nand UO_584 (O_584,N_9834,N_9813);
or UO_585 (O_585,N_9994,N_9933);
nand UO_586 (O_586,N_9972,N_9979);
nor UO_587 (O_587,N_9878,N_9887);
nor UO_588 (O_588,N_9979,N_9803);
xnor UO_589 (O_589,N_9826,N_9815);
and UO_590 (O_590,N_9992,N_9955);
xnor UO_591 (O_591,N_9858,N_9881);
or UO_592 (O_592,N_9959,N_9940);
xor UO_593 (O_593,N_9923,N_9825);
nor UO_594 (O_594,N_9887,N_9989);
and UO_595 (O_595,N_9911,N_9811);
nor UO_596 (O_596,N_9853,N_9909);
nand UO_597 (O_597,N_9947,N_9898);
nor UO_598 (O_598,N_9865,N_9870);
xnor UO_599 (O_599,N_9940,N_9863);
or UO_600 (O_600,N_9815,N_9874);
or UO_601 (O_601,N_9960,N_9968);
nand UO_602 (O_602,N_9841,N_9859);
nand UO_603 (O_603,N_9821,N_9935);
nor UO_604 (O_604,N_9858,N_9958);
xor UO_605 (O_605,N_9863,N_9902);
nor UO_606 (O_606,N_9858,N_9855);
and UO_607 (O_607,N_9934,N_9921);
and UO_608 (O_608,N_9926,N_9925);
and UO_609 (O_609,N_9866,N_9844);
nor UO_610 (O_610,N_9876,N_9847);
and UO_611 (O_611,N_9907,N_9856);
nor UO_612 (O_612,N_9917,N_9999);
and UO_613 (O_613,N_9925,N_9890);
nor UO_614 (O_614,N_9981,N_9950);
and UO_615 (O_615,N_9831,N_9957);
or UO_616 (O_616,N_9838,N_9889);
nand UO_617 (O_617,N_9953,N_9837);
or UO_618 (O_618,N_9821,N_9916);
nand UO_619 (O_619,N_9894,N_9969);
nor UO_620 (O_620,N_9971,N_9921);
or UO_621 (O_621,N_9841,N_9970);
nor UO_622 (O_622,N_9911,N_9810);
nor UO_623 (O_623,N_9923,N_9863);
nand UO_624 (O_624,N_9957,N_9885);
or UO_625 (O_625,N_9851,N_9971);
xnor UO_626 (O_626,N_9998,N_9859);
xnor UO_627 (O_627,N_9908,N_9855);
or UO_628 (O_628,N_9818,N_9920);
nor UO_629 (O_629,N_9807,N_9998);
or UO_630 (O_630,N_9868,N_9832);
and UO_631 (O_631,N_9941,N_9861);
or UO_632 (O_632,N_9946,N_9891);
nor UO_633 (O_633,N_9816,N_9862);
and UO_634 (O_634,N_9839,N_9814);
and UO_635 (O_635,N_9929,N_9870);
and UO_636 (O_636,N_9964,N_9903);
and UO_637 (O_637,N_9852,N_9825);
and UO_638 (O_638,N_9936,N_9876);
or UO_639 (O_639,N_9985,N_9914);
or UO_640 (O_640,N_9910,N_9837);
nand UO_641 (O_641,N_9814,N_9941);
xnor UO_642 (O_642,N_9981,N_9877);
and UO_643 (O_643,N_9849,N_9962);
xor UO_644 (O_644,N_9936,N_9935);
or UO_645 (O_645,N_9958,N_9811);
or UO_646 (O_646,N_9935,N_9920);
or UO_647 (O_647,N_9944,N_9973);
and UO_648 (O_648,N_9802,N_9909);
nand UO_649 (O_649,N_9904,N_9964);
or UO_650 (O_650,N_9966,N_9859);
nand UO_651 (O_651,N_9814,N_9843);
nor UO_652 (O_652,N_9843,N_9881);
nor UO_653 (O_653,N_9885,N_9987);
or UO_654 (O_654,N_9920,N_9816);
nor UO_655 (O_655,N_9986,N_9814);
or UO_656 (O_656,N_9936,N_9990);
or UO_657 (O_657,N_9869,N_9970);
nor UO_658 (O_658,N_9844,N_9972);
xnor UO_659 (O_659,N_9833,N_9888);
xnor UO_660 (O_660,N_9964,N_9950);
nand UO_661 (O_661,N_9811,N_9863);
or UO_662 (O_662,N_9960,N_9964);
and UO_663 (O_663,N_9857,N_9892);
and UO_664 (O_664,N_9985,N_9811);
and UO_665 (O_665,N_9866,N_9877);
and UO_666 (O_666,N_9993,N_9964);
nor UO_667 (O_667,N_9946,N_9882);
or UO_668 (O_668,N_9990,N_9858);
and UO_669 (O_669,N_9941,N_9835);
or UO_670 (O_670,N_9851,N_9908);
and UO_671 (O_671,N_9814,N_9913);
nand UO_672 (O_672,N_9932,N_9981);
nand UO_673 (O_673,N_9995,N_9892);
nand UO_674 (O_674,N_9946,N_9870);
nand UO_675 (O_675,N_9831,N_9821);
nand UO_676 (O_676,N_9933,N_9899);
xor UO_677 (O_677,N_9862,N_9996);
nor UO_678 (O_678,N_9812,N_9961);
and UO_679 (O_679,N_9814,N_9923);
nand UO_680 (O_680,N_9813,N_9944);
nor UO_681 (O_681,N_9919,N_9958);
nand UO_682 (O_682,N_9975,N_9954);
nand UO_683 (O_683,N_9813,N_9903);
or UO_684 (O_684,N_9887,N_9874);
nand UO_685 (O_685,N_9830,N_9904);
and UO_686 (O_686,N_9841,N_9838);
or UO_687 (O_687,N_9828,N_9868);
nor UO_688 (O_688,N_9876,N_9985);
and UO_689 (O_689,N_9869,N_9888);
xor UO_690 (O_690,N_9925,N_9850);
and UO_691 (O_691,N_9929,N_9833);
or UO_692 (O_692,N_9801,N_9941);
nor UO_693 (O_693,N_9856,N_9874);
nor UO_694 (O_694,N_9881,N_9965);
nand UO_695 (O_695,N_9844,N_9842);
xnor UO_696 (O_696,N_9858,N_9910);
and UO_697 (O_697,N_9869,N_9806);
and UO_698 (O_698,N_9991,N_9939);
and UO_699 (O_699,N_9936,N_9971);
nor UO_700 (O_700,N_9948,N_9908);
and UO_701 (O_701,N_9915,N_9816);
or UO_702 (O_702,N_9887,N_9830);
nand UO_703 (O_703,N_9851,N_9898);
nand UO_704 (O_704,N_9823,N_9954);
and UO_705 (O_705,N_9850,N_9932);
or UO_706 (O_706,N_9860,N_9896);
xor UO_707 (O_707,N_9806,N_9879);
xor UO_708 (O_708,N_9897,N_9994);
nand UO_709 (O_709,N_9880,N_9951);
or UO_710 (O_710,N_9974,N_9914);
xnor UO_711 (O_711,N_9865,N_9950);
and UO_712 (O_712,N_9940,N_9827);
nand UO_713 (O_713,N_9809,N_9894);
and UO_714 (O_714,N_9857,N_9969);
nor UO_715 (O_715,N_9865,N_9964);
or UO_716 (O_716,N_9815,N_9986);
nand UO_717 (O_717,N_9905,N_9854);
nor UO_718 (O_718,N_9861,N_9862);
nor UO_719 (O_719,N_9873,N_9946);
and UO_720 (O_720,N_9823,N_9889);
or UO_721 (O_721,N_9920,N_9873);
and UO_722 (O_722,N_9892,N_9850);
and UO_723 (O_723,N_9949,N_9847);
and UO_724 (O_724,N_9820,N_9915);
and UO_725 (O_725,N_9814,N_9874);
nor UO_726 (O_726,N_9914,N_9880);
nand UO_727 (O_727,N_9932,N_9959);
nor UO_728 (O_728,N_9858,N_9967);
and UO_729 (O_729,N_9909,N_9939);
and UO_730 (O_730,N_9991,N_9979);
or UO_731 (O_731,N_9964,N_9851);
or UO_732 (O_732,N_9888,N_9853);
nand UO_733 (O_733,N_9960,N_9813);
nor UO_734 (O_734,N_9874,N_9875);
or UO_735 (O_735,N_9886,N_9945);
and UO_736 (O_736,N_9923,N_9998);
xor UO_737 (O_737,N_9929,N_9855);
and UO_738 (O_738,N_9931,N_9942);
or UO_739 (O_739,N_9862,N_9915);
nand UO_740 (O_740,N_9908,N_9877);
nand UO_741 (O_741,N_9922,N_9880);
or UO_742 (O_742,N_9912,N_9911);
and UO_743 (O_743,N_9973,N_9804);
nand UO_744 (O_744,N_9823,N_9961);
xnor UO_745 (O_745,N_9905,N_9948);
or UO_746 (O_746,N_9874,N_9932);
nor UO_747 (O_747,N_9929,N_9991);
xor UO_748 (O_748,N_9886,N_9824);
xor UO_749 (O_749,N_9984,N_9975);
nor UO_750 (O_750,N_9881,N_9856);
nand UO_751 (O_751,N_9911,N_9985);
nand UO_752 (O_752,N_9826,N_9988);
and UO_753 (O_753,N_9912,N_9863);
or UO_754 (O_754,N_9921,N_9997);
and UO_755 (O_755,N_9977,N_9960);
nor UO_756 (O_756,N_9829,N_9842);
and UO_757 (O_757,N_9949,N_9943);
nor UO_758 (O_758,N_9864,N_9854);
xor UO_759 (O_759,N_9862,N_9975);
nand UO_760 (O_760,N_9907,N_9802);
nor UO_761 (O_761,N_9878,N_9963);
nand UO_762 (O_762,N_9815,N_9802);
nand UO_763 (O_763,N_9816,N_9895);
nor UO_764 (O_764,N_9886,N_9867);
or UO_765 (O_765,N_9887,N_9895);
or UO_766 (O_766,N_9992,N_9864);
nand UO_767 (O_767,N_9943,N_9917);
or UO_768 (O_768,N_9966,N_9829);
and UO_769 (O_769,N_9916,N_9895);
xor UO_770 (O_770,N_9849,N_9896);
or UO_771 (O_771,N_9847,N_9825);
or UO_772 (O_772,N_9861,N_9943);
and UO_773 (O_773,N_9982,N_9970);
nor UO_774 (O_774,N_9950,N_9871);
or UO_775 (O_775,N_9879,N_9988);
nor UO_776 (O_776,N_9883,N_9953);
xnor UO_777 (O_777,N_9831,N_9989);
xnor UO_778 (O_778,N_9953,N_9905);
nand UO_779 (O_779,N_9889,N_9828);
nand UO_780 (O_780,N_9834,N_9946);
nor UO_781 (O_781,N_9945,N_9983);
and UO_782 (O_782,N_9886,N_9980);
and UO_783 (O_783,N_9917,N_9827);
xnor UO_784 (O_784,N_9822,N_9835);
nor UO_785 (O_785,N_9932,N_9837);
and UO_786 (O_786,N_9982,N_9882);
or UO_787 (O_787,N_9930,N_9956);
nor UO_788 (O_788,N_9890,N_9882);
nor UO_789 (O_789,N_9980,N_9981);
and UO_790 (O_790,N_9830,N_9879);
xnor UO_791 (O_791,N_9948,N_9893);
and UO_792 (O_792,N_9882,N_9986);
nor UO_793 (O_793,N_9807,N_9971);
xor UO_794 (O_794,N_9971,N_9978);
nand UO_795 (O_795,N_9956,N_9999);
or UO_796 (O_796,N_9853,N_9854);
nand UO_797 (O_797,N_9983,N_9970);
or UO_798 (O_798,N_9876,N_9884);
and UO_799 (O_799,N_9975,N_9825);
nor UO_800 (O_800,N_9911,N_9883);
nor UO_801 (O_801,N_9955,N_9952);
nor UO_802 (O_802,N_9903,N_9937);
nor UO_803 (O_803,N_9877,N_9834);
or UO_804 (O_804,N_9927,N_9943);
and UO_805 (O_805,N_9801,N_9810);
xor UO_806 (O_806,N_9918,N_9930);
nand UO_807 (O_807,N_9946,N_9801);
nand UO_808 (O_808,N_9894,N_9928);
nand UO_809 (O_809,N_9904,N_9918);
or UO_810 (O_810,N_9935,N_9891);
or UO_811 (O_811,N_9857,N_9832);
nand UO_812 (O_812,N_9826,N_9916);
and UO_813 (O_813,N_9981,N_9867);
xnor UO_814 (O_814,N_9878,N_9858);
and UO_815 (O_815,N_9811,N_9974);
nor UO_816 (O_816,N_9924,N_9843);
or UO_817 (O_817,N_9923,N_9958);
nand UO_818 (O_818,N_9944,N_9850);
and UO_819 (O_819,N_9835,N_9845);
nand UO_820 (O_820,N_9870,N_9908);
nor UO_821 (O_821,N_9876,N_9841);
xnor UO_822 (O_822,N_9982,N_9890);
or UO_823 (O_823,N_9983,N_9824);
nor UO_824 (O_824,N_9818,N_9882);
nor UO_825 (O_825,N_9987,N_9883);
or UO_826 (O_826,N_9980,N_9891);
and UO_827 (O_827,N_9956,N_9944);
xor UO_828 (O_828,N_9903,N_9947);
nor UO_829 (O_829,N_9928,N_9859);
or UO_830 (O_830,N_9809,N_9956);
xnor UO_831 (O_831,N_9907,N_9949);
or UO_832 (O_832,N_9848,N_9826);
or UO_833 (O_833,N_9899,N_9833);
and UO_834 (O_834,N_9861,N_9981);
or UO_835 (O_835,N_9940,N_9900);
xnor UO_836 (O_836,N_9920,N_9886);
or UO_837 (O_837,N_9941,N_9978);
xor UO_838 (O_838,N_9867,N_9962);
nor UO_839 (O_839,N_9995,N_9877);
and UO_840 (O_840,N_9838,N_9817);
nand UO_841 (O_841,N_9871,N_9990);
nand UO_842 (O_842,N_9919,N_9969);
or UO_843 (O_843,N_9903,N_9884);
and UO_844 (O_844,N_9826,N_9813);
nand UO_845 (O_845,N_9937,N_9954);
or UO_846 (O_846,N_9886,N_9836);
xor UO_847 (O_847,N_9820,N_9948);
or UO_848 (O_848,N_9860,N_9969);
xnor UO_849 (O_849,N_9892,N_9981);
and UO_850 (O_850,N_9849,N_9824);
nand UO_851 (O_851,N_9829,N_9950);
and UO_852 (O_852,N_9933,N_9977);
and UO_853 (O_853,N_9999,N_9915);
or UO_854 (O_854,N_9965,N_9910);
xnor UO_855 (O_855,N_9819,N_9805);
and UO_856 (O_856,N_9963,N_9936);
and UO_857 (O_857,N_9929,N_9984);
xnor UO_858 (O_858,N_9862,N_9965);
xor UO_859 (O_859,N_9841,N_9910);
and UO_860 (O_860,N_9818,N_9928);
nor UO_861 (O_861,N_9943,N_9992);
xnor UO_862 (O_862,N_9823,N_9851);
or UO_863 (O_863,N_9896,N_9889);
nor UO_864 (O_864,N_9984,N_9841);
and UO_865 (O_865,N_9835,N_9982);
and UO_866 (O_866,N_9943,N_9913);
nor UO_867 (O_867,N_9948,N_9915);
xnor UO_868 (O_868,N_9816,N_9863);
nand UO_869 (O_869,N_9956,N_9871);
nand UO_870 (O_870,N_9834,N_9979);
nand UO_871 (O_871,N_9977,N_9917);
nand UO_872 (O_872,N_9941,N_9817);
nand UO_873 (O_873,N_9970,N_9899);
nor UO_874 (O_874,N_9927,N_9824);
xor UO_875 (O_875,N_9851,N_9830);
nor UO_876 (O_876,N_9810,N_9809);
and UO_877 (O_877,N_9916,N_9881);
nand UO_878 (O_878,N_9817,N_9998);
xor UO_879 (O_879,N_9824,N_9862);
nor UO_880 (O_880,N_9895,N_9967);
xor UO_881 (O_881,N_9933,N_9924);
xor UO_882 (O_882,N_9996,N_9900);
nor UO_883 (O_883,N_9810,N_9835);
or UO_884 (O_884,N_9981,N_9994);
nand UO_885 (O_885,N_9919,N_9807);
or UO_886 (O_886,N_9941,N_9864);
nand UO_887 (O_887,N_9809,N_9882);
nor UO_888 (O_888,N_9887,N_9833);
nor UO_889 (O_889,N_9830,N_9848);
or UO_890 (O_890,N_9862,N_9841);
nor UO_891 (O_891,N_9903,N_9954);
or UO_892 (O_892,N_9946,N_9958);
xor UO_893 (O_893,N_9818,N_9877);
or UO_894 (O_894,N_9942,N_9853);
nand UO_895 (O_895,N_9983,N_9849);
nor UO_896 (O_896,N_9851,N_9840);
nor UO_897 (O_897,N_9877,N_9852);
and UO_898 (O_898,N_9956,N_9977);
nand UO_899 (O_899,N_9847,N_9893);
or UO_900 (O_900,N_9996,N_9827);
nand UO_901 (O_901,N_9803,N_9827);
nand UO_902 (O_902,N_9860,N_9821);
or UO_903 (O_903,N_9936,N_9982);
or UO_904 (O_904,N_9973,N_9976);
nand UO_905 (O_905,N_9808,N_9858);
and UO_906 (O_906,N_9993,N_9925);
and UO_907 (O_907,N_9821,N_9971);
and UO_908 (O_908,N_9807,N_9814);
nand UO_909 (O_909,N_9840,N_9820);
nand UO_910 (O_910,N_9924,N_9986);
and UO_911 (O_911,N_9916,N_9862);
and UO_912 (O_912,N_9950,N_9959);
nor UO_913 (O_913,N_9831,N_9823);
nor UO_914 (O_914,N_9839,N_9843);
nor UO_915 (O_915,N_9997,N_9971);
xor UO_916 (O_916,N_9968,N_9829);
and UO_917 (O_917,N_9936,N_9834);
and UO_918 (O_918,N_9932,N_9832);
nor UO_919 (O_919,N_9826,N_9896);
nor UO_920 (O_920,N_9858,N_9945);
nand UO_921 (O_921,N_9866,N_9983);
and UO_922 (O_922,N_9983,N_9863);
xnor UO_923 (O_923,N_9952,N_9940);
or UO_924 (O_924,N_9841,N_9882);
nor UO_925 (O_925,N_9987,N_9931);
nor UO_926 (O_926,N_9926,N_9904);
nand UO_927 (O_927,N_9945,N_9996);
nand UO_928 (O_928,N_9851,N_9818);
and UO_929 (O_929,N_9937,N_9811);
or UO_930 (O_930,N_9925,N_9943);
or UO_931 (O_931,N_9852,N_9892);
and UO_932 (O_932,N_9897,N_9904);
xor UO_933 (O_933,N_9863,N_9877);
nand UO_934 (O_934,N_9983,N_9845);
nor UO_935 (O_935,N_9830,N_9853);
xnor UO_936 (O_936,N_9823,N_9993);
or UO_937 (O_937,N_9974,N_9985);
xor UO_938 (O_938,N_9854,N_9965);
xnor UO_939 (O_939,N_9972,N_9902);
or UO_940 (O_940,N_9997,N_9967);
or UO_941 (O_941,N_9810,N_9993);
xor UO_942 (O_942,N_9913,N_9817);
nor UO_943 (O_943,N_9996,N_9840);
nand UO_944 (O_944,N_9973,N_9834);
or UO_945 (O_945,N_9961,N_9819);
nor UO_946 (O_946,N_9812,N_9852);
nand UO_947 (O_947,N_9984,N_9964);
and UO_948 (O_948,N_9982,N_9998);
and UO_949 (O_949,N_9919,N_9957);
nand UO_950 (O_950,N_9966,N_9893);
nor UO_951 (O_951,N_9890,N_9861);
nor UO_952 (O_952,N_9962,N_9977);
xnor UO_953 (O_953,N_9927,N_9962);
and UO_954 (O_954,N_9904,N_9819);
or UO_955 (O_955,N_9870,N_9930);
nand UO_956 (O_956,N_9834,N_9853);
xnor UO_957 (O_957,N_9898,N_9854);
nand UO_958 (O_958,N_9998,N_9831);
nor UO_959 (O_959,N_9963,N_9912);
or UO_960 (O_960,N_9857,N_9845);
xnor UO_961 (O_961,N_9851,N_9828);
and UO_962 (O_962,N_9812,N_9986);
nand UO_963 (O_963,N_9846,N_9979);
xnor UO_964 (O_964,N_9941,N_9980);
and UO_965 (O_965,N_9809,N_9979);
nor UO_966 (O_966,N_9990,N_9989);
and UO_967 (O_967,N_9982,N_9980);
xor UO_968 (O_968,N_9893,N_9817);
and UO_969 (O_969,N_9894,N_9900);
xnor UO_970 (O_970,N_9994,N_9927);
xnor UO_971 (O_971,N_9967,N_9970);
nor UO_972 (O_972,N_9986,N_9980);
and UO_973 (O_973,N_9814,N_9845);
xor UO_974 (O_974,N_9976,N_9810);
xor UO_975 (O_975,N_9855,N_9813);
xnor UO_976 (O_976,N_9927,N_9931);
nor UO_977 (O_977,N_9862,N_9846);
nand UO_978 (O_978,N_9917,N_9817);
nor UO_979 (O_979,N_9985,N_9884);
and UO_980 (O_980,N_9897,N_9978);
xor UO_981 (O_981,N_9952,N_9916);
nand UO_982 (O_982,N_9825,N_9967);
nor UO_983 (O_983,N_9877,N_9987);
nand UO_984 (O_984,N_9948,N_9959);
xor UO_985 (O_985,N_9934,N_9840);
and UO_986 (O_986,N_9998,N_9828);
nor UO_987 (O_987,N_9957,N_9810);
xnor UO_988 (O_988,N_9884,N_9968);
nor UO_989 (O_989,N_9815,N_9945);
or UO_990 (O_990,N_9819,N_9815);
nor UO_991 (O_991,N_9935,N_9801);
nand UO_992 (O_992,N_9837,N_9894);
nor UO_993 (O_993,N_9825,N_9989);
nor UO_994 (O_994,N_9891,N_9928);
xor UO_995 (O_995,N_9930,N_9815);
nor UO_996 (O_996,N_9807,N_9934);
and UO_997 (O_997,N_9897,N_9906);
nor UO_998 (O_998,N_9999,N_9861);
nor UO_999 (O_999,N_9877,N_9992);
nor UO_1000 (O_1000,N_9955,N_9834);
xnor UO_1001 (O_1001,N_9961,N_9836);
and UO_1002 (O_1002,N_9802,N_9984);
nor UO_1003 (O_1003,N_9841,N_9915);
or UO_1004 (O_1004,N_9967,N_9800);
nor UO_1005 (O_1005,N_9828,N_9990);
nand UO_1006 (O_1006,N_9989,N_9960);
nor UO_1007 (O_1007,N_9898,N_9812);
xor UO_1008 (O_1008,N_9895,N_9989);
nor UO_1009 (O_1009,N_9832,N_9845);
and UO_1010 (O_1010,N_9958,N_9801);
xnor UO_1011 (O_1011,N_9985,N_9891);
nor UO_1012 (O_1012,N_9950,N_9968);
or UO_1013 (O_1013,N_9800,N_9835);
nand UO_1014 (O_1014,N_9941,N_9870);
nand UO_1015 (O_1015,N_9821,N_9878);
nand UO_1016 (O_1016,N_9895,N_9836);
nor UO_1017 (O_1017,N_9998,N_9968);
nor UO_1018 (O_1018,N_9928,N_9817);
nor UO_1019 (O_1019,N_9931,N_9965);
nand UO_1020 (O_1020,N_9913,N_9966);
or UO_1021 (O_1021,N_9868,N_9949);
nor UO_1022 (O_1022,N_9929,N_9999);
nor UO_1023 (O_1023,N_9875,N_9918);
nor UO_1024 (O_1024,N_9975,N_9951);
nand UO_1025 (O_1025,N_9948,N_9815);
and UO_1026 (O_1026,N_9941,N_9977);
xor UO_1027 (O_1027,N_9970,N_9902);
nand UO_1028 (O_1028,N_9949,N_9942);
xor UO_1029 (O_1029,N_9853,N_9920);
and UO_1030 (O_1030,N_9854,N_9991);
or UO_1031 (O_1031,N_9958,N_9988);
or UO_1032 (O_1032,N_9925,N_9922);
xor UO_1033 (O_1033,N_9853,N_9963);
nand UO_1034 (O_1034,N_9993,N_9915);
and UO_1035 (O_1035,N_9927,N_9881);
xnor UO_1036 (O_1036,N_9804,N_9944);
nand UO_1037 (O_1037,N_9929,N_9975);
xnor UO_1038 (O_1038,N_9848,N_9904);
nand UO_1039 (O_1039,N_9944,N_9905);
xnor UO_1040 (O_1040,N_9866,N_9904);
xnor UO_1041 (O_1041,N_9869,N_9929);
or UO_1042 (O_1042,N_9993,N_9892);
and UO_1043 (O_1043,N_9834,N_9932);
and UO_1044 (O_1044,N_9833,N_9810);
and UO_1045 (O_1045,N_9805,N_9979);
and UO_1046 (O_1046,N_9936,N_9868);
nand UO_1047 (O_1047,N_9913,N_9891);
or UO_1048 (O_1048,N_9815,N_9830);
and UO_1049 (O_1049,N_9926,N_9874);
or UO_1050 (O_1050,N_9814,N_9877);
and UO_1051 (O_1051,N_9897,N_9960);
or UO_1052 (O_1052,N_9915,N_9985);
nor UO_1053 (O_1053,N_9884,N_9832);
and UO_1054 (O_1054,N_9919,N_9872);
nor UO_1055 (O_1055,N_9955,N_9928);
or UO_1056 (O_1056,N_9951,N_9985);
or UO_1057 (O_1057,N_9883,N_9966);
or UO_1058 (O_1058,N_9927,N_9971);
and UO_1059 (O_1059,N_9802,N_9804);
nor UO_1060 (O_1060,N_9834,N_9899);
nand UO_1061 (O_1061,N_9934,N_9953);
and UO_1062 (O_1062,N_9944,N_9810);
and UO_1063 (O_1063,N_9890,N_9888);
nor UO_1064 (O_1064,N_9808,N_9960);
nor UO_1065 (O_1065,N_9912,N_9860);
xor UO_1066 (O_1066,N_9882,N_9853);
nand UO_1067 (O_1067,N_9849,N_9953);
nand UO_1068 (O_1068,N_9886,N_9828);
and UO_1069 (O_1069,N_9958,N_9944);
or UO_1070 (O_1070,N_9970,N_9843);
nor UO_1071 (O_1071,N_9961,N_9832);
nor UO_1072 (O_1072,N_9950,N_9803);
xor UO_1073 (O_1073,N_9853,N_9860);
xnor UO_1074 (O_1074,N_9903,N_9950);
nor UO_1075 (O_1075,N_9822,N_9915);
and UO_1076 (O_1076,N_9987,N_9897);
nor UO_1077 (O_1077,N_9859,N_9883);
or UO_1078 (O_1078,N_9940,N_9916);
xnor UO_1079 (O_1079,N_9819,N_9970);
nand UO_1080 (O_1080,N_9888,N_9990);
nand UO_1081 (O_1081,N_9887,N_9867);
nand UO_1082 (O_1082,N_9815,N_9903);
and UO_1083 (O_1083,N_9890,N_9848);
nor UO_1084 (O_1084,N_9800,N_9806);
and UO_1085 (O_1085,N_9994,N_9943);
nor UO_1086 (O_1086,N_9941,N_9959);
or UO_1087 (O_1087,N_9827,N_9886);
or UO_1088 (O_1088,N_9850,N_9985);
and UO_1089 (O_1089,N_9831,N_9822);
nand UO_1090 (O_1090,N_9926,N_9909);
nand UO_1091 (O_1091,N_9878,N_9848);
xnor UO_1092 (O_1092,N_9925,N_9834);
xor UO_1093 (O_1093,N_9845,N_9972);
xor UO_1094 (O_1094,N_9970,N_9901);
nor UO_1095 (O_1095,N_9811,N_9955);
nor UO_1096 (O_1096,N_9906,N_9902);
nor UO_1097 (O_1097,N_9847,N_9804);
xnor UO_1098 (O_1098,N_9992,N_9862);
and UO_1099 (O_1099,N_9822,N_9873);
nor UO_1100 (O_1100,N_9867,N_9928);
xnor UO_1101 (O_1101,N_9821,N_9886);
or UO_1102 (O_1102,N_9897,N_9804);
and UO_1103 (O_1103,N_9933,N_9855);
and UO_1104 (O_1104,N_9948,N_9945);
nor UO_1105 (O_1105,N_9901,N_9844);
xor UO_1106 (O_1106,N_9921,N_9862);
xnor UO_1107 (O_1107,N_9867,N_9883);
nor UO_1108 (O_1108,N_9824,N_9861);
nand UO_1109 (O_1109,N_9915,N_9968);
nand UO_1110 (O_1110,N_9882,N_9977);
nand UO_1111 (O_1111,N_9821,N_9914);
or UO_1112 (O_1112,N_9863,N_9974);
xnor UO_1113 (O_1113,N_9835,N_9877);
xor UO_1114 (O_1114,N_9846,N_9809);
and UO_1115 (O_1115,N_9823,N_9981);
nand UO_1116 (O_1116,N_9862,N_9949);
or UO_1117 (O_1117,N_9985,N_9832);
or UO_1118 (O_1118,N_9825,N_9853);
or UO_1119 (O_1119,N_9831,N_9904);
nand UO_1120 (O_1120,N_9997,N_9961);
and UO_1121 (O_1121,N_9962,N_9902);
xnor UO_1122 (O_1122,N_9922,N_9896);
nand UO_1123 (O_1123,N_9847,N_9870);
nand UO_1124 (O_1124,N_9975,N_9955);
or UO_1125 (O_1125,N_9871,N_9829);
or UO_1126 (O_1126,N_9914,N_9923);
nand UO_1127 (O_1127,N_9977,N_9899);
nand UO_1128 (O_1128,N_9981,N_9984);
or UO_1129 (O_1129,N_9938,N_9901);
nor UO_1130 (O_1130,N_9964,N_9859);
or UO_1131 (O_1131,N_9989,N_9839);
and UO_1132 (O_1132,N_9947,N_9833);
xor UO_1133 (O_1133,N_9874,N_9840);
xor UO_1134 (O_1134,N_9978,N_9963);
nor UO_1135 (O_1135,N_9917,N_9981);
nor UO_1136 (O_1136,N_9898,N_9824);
and UO_1137 (O_1137,N_9971,N_9904);
nor UO_1138 (O_1138,N_9827,N_9896);
or UO_1139 (O_1139,N_9894,N_9822);
or UO_1140 (O_1140,N_9952,N_9976);
and UO_1141 (O_1141,N_9988,N_9900);
nand UO_1142 (O_1142,N_9845,N_9834);
and UO_1143 (O_1143,N_9874,N_9999);
xor UO_1144 (O_1144,N_9923,N_9865);
xnor UO_1145 (O_1145,N_9972,N_9952);
or UO_1146 (O_1146,N_9968,N_9956);
and UO_1147 (O_1147,N_9951,N_9814);
or UO_1148 (O_1148,N_9975,N_9890);
xnor UO_1149 (O_1149,N_9807,N_9839);
or UO_1150 (O_1150,N_9946,N_9899);
and UO_1151 (O_1151,N_9898,N_9801);
nand UO_1152 (O_1152,N_9846,N_9850);
or UO_1153 (O_1153,N_9963,N_9964);
and UO_1154 (O_1154,N_9914,N_9902);
and UO_1155 (O_1155,N_9808,N_9806);
xor UO_1156 (O_1156,N_9839,N_9877);
or UO_1157 (O_1157,N_9818,N_9866);
nor UO_1158 (O_1158,N_9943,N_9865);
or UO_1159 (O_1159,N_9876,N_9823);
xnor UO_1160 (O_1160,N_9841,N_9803);
and UO_1161 (O_1161,N_9909,N_9941);
or UO_1162 (O_1162,N_9895,N_9849);
or UO_1163 (O_1163,N_9955,N_9986);
nand UO_1164 (O_1164,N_9839,N_9859);
xor UO_1165 (O_1165,N_9827,N_9984);
nand UO_1166 (O_1166,N_9998,N_9822);
and UO_1167 (O_1167,N_9883,N_9976);
xor UO_1168 (O_1168,N_9930,N_9947);
or UO_1169 (O_1169,N_9984,N_9995);
nand UO_1170 (O_1170,N_9868,N_9922);
nand UO_1171 (O_1171,N_9847,N_9989);
and UO_1172 (O_1172,N_9903,N_9970);
nor UO_1173 (O_1173,N_9853,N_9930);
xnor UO_1174 (O_1174,N_9979,N_9868);
xor UO_1175 (O_1175,N_9982,N_9809);
or UO_1176 (O_1176,N_9912,N_9943);
or UO_1177 (O_1177,N_9840,N_9973);
nor UO_1178 (O_1178,N_9973,N_9803);
nor UO_1179 (O_1179,N_9927,N_9878);
nor UO_1180 (O_1180,N_9953,N_9977);
nor UO_1181 (O_1181,N_9963,N_9953);
nor UO_1182 (O_1182,N_9854,N_9940);
or UO_1183 (O_1183,N_9898,N_9918);
or UO_1184 (O_1184,N_9918,N_9800);
or UO_1185 (O_1185,N_9967,N_9822);
and UO_1186 (O_1186,N_9923,N_9853);
xnor UO_1187 (O_1187,N_9985,N_9921);
xor UO_1188 (O_1188,N_9889,N_9931);
and UO_1189 (O_1189,N_9937,N_9969);
xor UO_1190 (O_1190,N_9812,N_9819);
xnor UO_1191 (O_1191,N_9800,N_9983);
nor UO_1192 (O_1192,N_9890,N_9833);
xor UO_1193 (O_1193,N_9814,N_9908);
nor UO_1194 (O_1194,N_9931,N_9903);
nand UO_1195 (O_1195,N_9901,N_9873);
xor UO_1196 (O_1196,N_9998,N_9830);
nor UO_1197 (O_1197,N_9932,N_9927);
nor UO_1198 (O_1198,N_9974,N_9859);
nand UO_1199 (O_1199,N_9965,N_9956);
nor UO_1200 (O_1200,N_9875,N_9911);
or UO_1201 (O_1201,N_9999,N_9933);
nand UO_1202 (O_1202,N_9936,N_9809);
nand UO_1203 (O_1203,N_9908,N_9807);
xnor UO_1204 (O_1204,N_9923,N_9811);
or UO_1205 (O_1205,N_9847,N_9935);
nand UO_1206 (O_1206,N_9836,N_9851);
xnor UO_1207 (O_1207,N_9819,N_9994);
or UO_1208 (O_1208,N_9968,N_9979);
nand UO_1209 (O_1209,N_9885,N_9960);
nand UO_1210 (O_1210,N_9978,N_9891);
xor UO_1211 (O_1211,N_9959,N_9827);
nand UO_1212 (O_1212,N_9842,N_9851);
nand UO_1213 (O_1213,N_9913,N_9967);
nor UO_1214 (O_1214,N_9971,N_9938);
or UO_1215 (O_1215,N_9981,N_9829);
or UO_1216 (O_1216,N_9942,N_9933);
nand UO_1217 (O_1217,N_9975,N_9888);
nor UO_1218 (O_1218,N_9948,N_9979);
xor UO_1219 (O_1219,N_9845,N_9867);
nand UO_1220 (O_1220,N_9857,N_9930);
and UO_1221 (O_1221,N_9845,N_9914);
nor UO_1222 (O_1222,N_9879,N_9861);
nand UO_1223 (O_1223,N_9913,N_9970);
xnor UO_1224 (O_1224,N_9972,N_9992);
and UO_1225 (O_1225,N_9933,N_9804);
nand UO_1226 (O_1226,N_9940,N_9977);
nand UO_1227 (O_1227,N_9854,N_9967);
and UO_1228 (O_1228,N_9908,N_9958);
and UO_1229 (O_1229,N_9914,N_9904);
xor UO_1230 (O_1230,N_9825,N_9962);
and UO_1231 (O_1231,N_9813,N_9809);
or UO_1232 (O_1232,N_9892,N_9856);
xor UO_1233 (O_1233,N_9885,N_9803);
and UO_1234 (O_1234,N_9983,N_9997);
and UO_1235 (O_1235,N_9803,N_9849);
xor UO_1236 (O_1236,N_9883,N_9884);
or UO_1237 (O_1237,N_9986,N_9843);
nor UO_1238 (O_1238,N_9906,N_9920);
or UO_1239 (O_1239,N_9941,N_9976);
or UO_1240 (O_1240,N_9800,N_9898);
and UO_1241 (O_1241,N_9980,N_9856);
nand UO_1242 (O_1242,N_9926,N_9814);
xnor UO_1243 (O_1243,N_9875,N_9850);
and UO_1244 (O_1244,N_9813,N_9957);
and UO_1245 (O_1245,N_9876,N_9849);
and UO_1246 (O_1246,N_9865,N_9818);
xor UO_1247 (O_1247,N_9890,N_9977);
and UO_1248 (O_1248,N_9810,N_9948);
or UO_1249 (O_1249,N_9843,N_9883);
nand UO_1250 (O_1250,N_9995,N_9990);
nand UO_1251 (O_1251,N_9867,N_9820);
nor UO_1252 (O_1252,N_9844,N_9907);
xor UO_1253 (O_1253,N_9988,N_9894);
xnor UO_1254 (O_1254,N_9812,N_9823);
xor UO_1255 (O_1255,N_9856,N_9801);
and UO_1256 (O_1256,N_9904,N_9949);
nand UO_1257 (O_1257,N_9948,N_9839);
nor UO_1258 (O_1258,N_9969,N_9878);
nand UO_1259 (O_1259,N_9919,N_9914);
nor UO_1260 (O_1260,N_9806,N_9817);
or UO_1261 (O_1261,N_9896,N_9854);
nand UO_1262 (O_1262,N_9842,N_9995);
or UO_1263 (O_1263,N_9990,N_9830);
or UO_1264 (O_1264,N_9920,N_9954);
or UO_1265 (O_1265,N_9929,N_9874);
nand UO_1266 (O_1266,N_9883,N_9904);
or UO_1267 (O_1267,N_9963,N_9973);
nand UO_1268 (O_1268,N_9917,N_9898);
or UO_1269 (O_1269,N_9809,N_9833);
or UO_1270 (O_1270,N_9961,N_9941);
or UO_1271 (O_1271,N_9988,N_9839);
or UO_1272 (O_1272,N_9910,N_9875);
nor UO_1273 (O_1273,N_9910,N_9948);
xnor UO_1274 (O_1274,N_9857,N_9980);
or UO_1275 (O_1275,N_9980,N_9993);
nand UO_1276 (O_1276,N_9932,N_9804);
nand UO_1277 (O_1277,N_9951,N_9887);
xor UO_1278 (O_1278,N_9965,N_9849);
nand UO_1279 (O_1279,N_9965,N_9803);
or UO_1280 (O_1280,N_9951,N_9907);
xnor UO_1281 (O_1281,N_9852,N_9920);
nand UO_1282 (O_1282,N_9943,N_9822);
nand UO_1283 (O_1283,N_9897,N_9873);
nor UO_1284 (O_1284,N_9877,N_9836);
xnor UO_1285 (O_1285,N_9945,N_9982);
or UO_1286 (O_1286,N_9929,N_9889);
xnor UO_1287 (O_1287,N_9938,N_9990);
xor UO_1288 (O_1288,N_9879,N_9950);
or UO_1289 (O_1289,N_9869,N_9962);
and UO_1290 (O_1290,N_9990,N_9834);
or UO_1291 (O_1291,N_9812,N_9834);
and UO_1292 (O_1292,N_9991,N_9903);
xor UO_1293 (O_1293,N_9845,N_9827);
and UO_1294 (O_1294,N_9895,N_9818);
nand UO_1295 (O_1295,N_9985,N_9944);
nand UO_1296 (O_1296,N_9884,N_9979);
or UO_1297 (O_1297,N_9887,N_9999);
or UO_1298 (O_1298,N_9867,N_9975);
nand UO_1299 (O_1299,N_9831,N_9829);
and UO_1300 (O_1300,N_9846,N_9932);
or UO_1301 (O_1301,N_9914,N_9901);
nor UO_1302 (O_1302,N_9894,N_9898);
or UO_1303 (O_1303,N_9975,N_9999);
xor UO_1304 (O_1304,N_9936,N_9899);
xnor UO_1305 (O_1305,N_9869,N_9817);
or UO_1306 (O_1306,N_9821,N_9980);
and UO_1307 (O_1307,N_9994,N_9820);
nand UO_1308 (O_1308,N_9920,N_9937);
or UO_1309 (O_1309,N_9977,N_9835);
nand UO_1310 (O_1310,N_9990,N_9892);
and UO_1311 (O_1311,N_9991,N_9847);
and UO_1312 (O_1312,N_9951,N_9931);
nand UO_1313 (O_1313,N_9817,N_9946);
and UO_1314 (O_1314,N_9955,N_9835);
nor UO_1315 (O_1315,N_9930,N_9995);
nand UO_1316 (O_1316,N_9953,N_9908);
xnor UO_1317 (O_1317,N_9964,N_9893);
nor UO_1318 (O_1318,N_9846,N_9947);
xor UO_1319 (O_1319,N_9915,N_9958);
or UO_1320 (O_1320,N_9883,N_9828);
nor UO_1321 (O_1321,N_9907,N_9842);
xnor UO_1322 (O_1322,N_9971,N_9998);
xor UO_1323 (O_1323,N_9978,N_9884);
nor UO_1324 (O_1324,N_9864,N_9915);
or UO_1325 (O_1325,N_9922,N_9816);
xor UO_1326 (O_1326,N_9802,N_9801);
or UO_1327 (O_1327,N_9834,N_9833);
nand UO_1328 (O_1328,N_9995,N_9948);
nor UO_1329 (O_1329,N_9915,N_9994);
and UO_1330 (O_1330,N_9933,N_9963);
nor UO_1331 (O_1331,N_9924,N_9931);
xor UO_1332 (O_1332,N_9912,N_9802);
nor UO_1333 (O_1333,N_9826,N_9806);
xor UO_1334 (O_1334,N_9889,N_9860);
and UO_1335 (O_1335,N_9857,N_9951);
nand UO_1336 (O_1336,N_9925,N_9910);
nor UO_1337 (O_1337,N_9990,N_9882);
xor UO_1338 (O_1338,N_9877,N_9947);
nor UO_1339 (O_1339,N_9800,N_9944);
nand UO_1340 (O_1340,N_9903,N_9904);
or UO_1341 (O_1341,N_9902,N_9968);
xor UO_1342 (O_1342,N_9813,N_9941);
xor UO_1343 (O_1343,N_9967,N_9899);
nor UO_1344 (O_1344,N_9868,N_9960);
nand UO_1345 (O_1345,N_9990,N_9851);
nand UO_1346 (O_1346,N_9834,N_9965);
or UO_1347 (O_1347,N_9895,N_9899);
and UO_1348 (O_1348,N_9997,N_9858);
nor UO_1349 (O_1349,N_9886,N_9852);
and UO_1350 (O_1350,N_9974,N_9937);
or UO_1351 (O_1351,N_9918,N_9835);
xor UO_1352 (O_1352,N_9982,N_9873);
xnor UO_1353 (O_1353,N_9991,N_9882);
nand UO_1354 (O_1354,N_9825,N_9926);
or UO_1355 (O_1355,N_9965,N_9961);
and UO_1356 (O_1356,N_9877,N_9861);
nor UO_1357 (O_1357,N_9893,N_9876);
or UO_1358 (O_1358,N_9825,N_9818);
or UO_1359 (O_1359,N_9917,N_9844);
xnor UO_1360 (O_1360,N_9845,N_9903);
xnor UO_1361 (O_1361,N_9941,N_9994);
nor UO_1362 (O_1362,N_9972,N_9827);
nand UO_1363 (O_1363,N_9817,N_9820);
nand UO_1364 (O_1364,N_9959,N_9951);
nand UO_1365 (O_1365,N_9849,N_9941);
nor UO_1366 (O_1366,N_9955,N_9830);
xor UO_1367 (O_1367,N_9945,N_9882);
nand UO_1368 (O_1368,N_9931,N_9938);
or UO_1369 (O_1369,N_9978,N_9805);
nand UO_1370 (O_1370,N_9828,N_9878);
nor UO_1371 (O_1371,N_9811,N_9878);
nor UO_1372 (O_1372,N_9875,N_9801);
xnor UO_1373 (O_1373,N_9901,N_9987);
xnor UO_1374 (O_1374,N_9947,N_9820);
and UO_1375 (O_1375,N_9970,N_9994);
nor UO_1376 (O_1376,N_9903,N_9941);
and UO_1377 (O_1377,N_9893,N_9802);
xnor UO_1378 (O_1378,N_9912,N_9871);
nand UO_1379 (O_1379,N_9979,N_9826);
or UO_1380 (O_1380,N_9933,N_9905);
nand UO_1381 (O_1381,N_9955,N_9906);
nor UO_1382 (O_1382,N_9859,N_9969);
nor UO_1383 (O_1383,N_9924,N_9961);
and UO_1384 (O_1384,N_9822,N_9823);
xnor UO_1385 (O_1385,N_9807,N_9855);
nor UO_1386 (O_1386,N_9872,N_9839);
nand UO_1387 (O_1387,N_9973,N_9802);
or UO_1388 (O_1388,N_9975,N_9849);
nand UO_1389 (O_1389,N_9927,N_9867);
xor UO_1390 (O_1390,N_9913,N_9992);
nand UO_1391 (O_1391,N_9988,N_9828);
and UO_1392 (O_1392,N_9845,N_9831);
xor UO_1393 (O_1393,N_9904,N_9917);
and UO_1394 (O_1394,N_9809,N_9968);
nor UO_1395 (O_1395,N_9954,N_9930);
nor UO_1396 (O_1396,N_9982,N_9995);
or UO_1397 (O_1397,N_9808,N_9959);
xnor UO_1398 (O_1398,N_9972,N_9912);
and UO_1399 (O_1399,N_9986,N_9912);
nor UO_1400 (O_1400,N_9972,N_9961);
nand UO_1401 (O_1401,N_9867,N_9844);
nor UO_1402 (O_1402,N_9884,N_9917);
or UO_1403 (O_1403,N_9918,N_9903);
nor UO_1404 (O_1404,N_9866,N_9993);
and UO_1405 (O_1405,N_9994,N_9802);
nor UO_1406 (O_1406,N_9803,N_9896);
or UO_1407 (O_1407,N_9917,N_9846);
or UO_1408 (O_1408,N_9975,N_9880);
nor UO_1409 (O_1409,N_9800,N_9829);
xor UO_1410 (O_1410,N_9870,N_9949);
and UO_1411 (O_1411,N_9908,N_9996);
nor UO_1412 (O_1412,N_9912,N_9856);
nor UO_1413 (O_1413,N_9944,N_9909);
and UO_1414 (O_1414,N_9945,N_9848);
xor UO_1415 (O_1415,N_9812,N_9952);
nor UO_1416 (O_1416,N_9979,N_9839);
xnor UO_1417 (O_1417,N_9945,N_9863);
nand UO_1418 (O_1418,N_9873,N_9968);
nor UO_1419 (O_1419,N_9988,N_9928);
or UO_1420 (O_1420,N_9918,N_9998);
and UO_1421 (O_1421,N_9987,N_9939);
or UO_1422 (O_1422,N_9867,N_9882);
and UO_1423 (O_1423,N_9955,N_9869);
nand UO_1424 (O_1424,N_9961,N_9835);
nor UO_1425 (O_1425,N_9837,N_9830);
xnor UO_1426 (O_1426,N_9997,N_9845);
or UO_1427 (O_1427,N_9941,N_9924);
nor UO_1428 (O_1428,N_9943,N_9818);
nand UO_1429 (O_1429,N_9955,N_9935);
nand UO_1430 (O_1430,N_9853,N_9875);
or UO_1431 (O_1431,N_9853,N_9904);
and UO_1432 (O_1432,N_9972,N_9926);
xor UO_1433 (O_1433,N_9935,N_9946);
nand UO_1434 (O_1434,N_9917,N_9890);
xor UO_1435 (O_1435,N_9834,N_9890);
and UO_1436 (O_1436,N_9905,N_9823);
nand UO_1437 (O_1437,N_9926,N_9898);
or UO_1438 (O_1438,N_9909,N_9856);
xnor UO_1439 (O_1439,N_9899,N_9831);
nand UO_1440 (O_1440,N_9874,N_9872);
nor UO_1441 (O_1441,N_9939,N_9883);
xnor UO_1442 (O_1442,N_9809,N_9960);
or UO_1443 (O_1443,N_9855,N_9963);
and UO_1444 (O_1444,N_9969,N_9869);
and UO_1445 (O_1445,N_9812,N_9928);
xor UO_1446 (O_1446,N_9958,N_9945);
xor UO_1447 (O_1447,N_9922,N_9814);
nand UO_1448 (O_1448,N_9998,N_9896);
xnor UO_1449 (O_1449,N_9871,N_9836);
xnor UO_1450 (O_1450,N_9820,N_9987);
xnor UO_1451 (O_1451,N_9891,N_9917);
nand UO_1452 (O_1452,N_9879,N_9854);
nor UO_1453 (O_1453,N_9937,N_9907);
and UO_1454 (O_1454,N_9856,N_9953);
nor UO_1455 (O_1455,N_9939,N_9947);
nand UO_1456 (O_1456,N_9943,N_9814);
and UO_1457 (O_1457,N_9930,N_9855);
and UO_1458 (O_1458,N_9825,N_9812);
nand UO_1459 (O_1459,N_9839,N_9836);
nor UO_1460 (O_1460,N_9824,N_9951);
nor UO_1461 (O_1461,N_9977,N_9873);
nand UO_1462 (O_1462,N_9879,N_9896);
nand UO_1463 (O_1463,N_9830,N_9821);
nand UO_1464 (O_1464,N_9918,N_9810);
nand UO_1465 (O_1465,N_9912,N_9854);
nor UO_1466 (O_1466,N_9817,N_9989);
and UO_1467 (O_1467,N_9989,N_9865);
nor UO_1468 (O_1468,N_9867,N_9878);
or UO_1469 (O_1469,N_9997,N_9928);
or UO_1470 (O_1470,N_9828,N_9941);
xnor UO_1471 (O_1471,N_9806,N_9816);
or UO_1472 (O_1472,N_9954,N_9858);
xor UO_1473 (O_1473,N_9802,N_9856);
nand UO_1474 (O_1474,N_9855,N_9902);
nor UO_1475 (O_1475,N_9896,N_9900);
nor UO_1476 (O_1476,N_9836,N_9981);
nand UO_1477 (O_1477,N_9934,N_9937);
nor UO_1478 (O_1478,N_9818,N_9879);
xnor UO_1479 (O_1479,N_9899,N_9990);
xor UO_1480 (O_1480,N_9851,N_9998);
xnor UO_1481 (O_1481,N_9894,N_9889);
xnor UO_1482 (O_1482,N_9886,N_9925);
xor UO_1483 (O_1483,N_9999,N_9899);
xor UO_1484 (O_1484,N_9962,N_9916);
xnor UO_1485 (O_1485,N_9933,N_9927);
nor UO_1486 (O_1486,N_9877,N_9926);
nor UO_1487 (O_1487,N_9933,N_9894);
or UO_1488 (O_1488,N_9903,N_9958);
nand UO_1489 (O_1489,N_9871,N_9877);
xor UO_1490 (O_1490,N_9924,N_9923);
or UO_1491 (O_1491,N_9807,N_9876);
or UO_1492 (O_1492,N_9992,N_9944);
xor UO_1493 (O_1493,N_9987,N_9839);
nand UO_1494 (O_1494,N_9870,N_9920);
xor UO_1495 (O_1495,N_9920,N_9881);
and UO_1496 (O_1496,N_9821,N_9862);
nor UO_1497 (O_1497,N_9991,N_9951);
and UO_1498 (O_1498,N_9811,N_9918);
xor UO_1499 (O_1499,N_9819,N_9996);
endmodule