module basic_1000_10000_1500_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_927,In_516);
nor U1 (N_1,In_104,In_586);
and U2 (N_2,In_783,In_771);
xnor U3 (N_3,In_979,In_671);
xor U4 (N_4,In_686,In_898);
xor U5 (N_5,In_740,In_751);
nand U6 (N_6,In_39,In_450);
or U7 (N_7,In_305,In_553);
xor U8 (N_8,In_398,In_931);
xor U9 (N_9,In_344,In_907);
nand U10 (N_10,In_571,In_619);
xor U11 (N_11,In_690,In_590);
or U12 (N_12,In_567,In_718);
or U13 (N_13,In_174,In_465);
nor U14 (N_14,In_6,In_521);
xor U15 (N_15,In_573,In_112);
or U16 (N_16,In_741,In_318);
or U17 (N_17,In_90,In_727);
or U18 (N_18,In_446,In_152);
and U19 (N_19,In_724,In_426);
nor U20 (N_20,In_44,In_642);
or U21 (N_21,In_796,In_443);
nor U22 (N_22,In_591,In_944);
xor U23 (N_23,In_986,In_476);
and U24 (N_24,In_494,In_468);
nand U25 (N_25,In_933,In_752);
nand U26 (N_26,In_525,In_714);
nor U27 (N_27,In_60,In_940);
and U28 (N_28,In_142,In_925);
nand U29 (N_29,In_851,In_462);
xor U30 (N_30,In_330,In_206);
and U31 (N_31,In_618,In_456);
nor U32 (N_32,In_71,In_599);
nand U33 (N_33,In_916,In_273);
nand U34 (N_34,In_262,In_773);
nor U35 (N_35,In_864,In_762);
xor U36 (N_36,In_80,In_185);
and U37 (N_37,In_164,In_277);
and U38 (N_38,In_95,In_540);
nor U39 (N_39,In_939,In_326);
and U40 (N_40,In_255,In_761);
nand U41 (N_41,In_113,In_982);
nand U42 (N_42,In_106,In_375);
nand U43 (N_43,In_186,In_632);
and U44 (N_44,In_269,In_792);
nand U45 (N_45,In_872,In_109);
and U46 (N_46,In_656,In_423);
nor U47 (N_47,In_86,In_329);
and U48 (N_48,In_876,In_767);
xnor U49 (N_49,In_454,In_806);
and U50 (N_50,In_484,In_341);
nand U51 (N_51,In_922,In_148);
nand U52 (N_52,In_665,In_801);
nand U53 (N_53,In_854,In_968);
or U54 (N_54,In_886,In_144);
xnor U55 (N_55,In_75,In_808);
xor U56 (N_56,In_988,In_256);
nand U57 (N_57,In_627,In_202);
xnor U58 (N_58,In_23,In_178);
xnor U59 (N_59,In_477,In_531);
xnor U60 (N_60,In_452,In_649);
and U61 (N_61,In_629,In_388);
xor U62 (N_62,In_409,In_950);
xor U63 (N_63,In_893,In_296);
xor U64 (N_64,In_879,In_820);
or U65 (N_65,In_897,In_810);
nor U66 (N_66,In_858,In_600);
xor U67 (N_67,In_617,In_63);
and U68 (N_68,In_948,In_194);
and U69 (N_69,In_622,In_680);
or U70 (N_70,In_809,In_62);
nor U71 (N_71,In_190,In_403);
and U72 (N_72,In_140,In_957);
nand U73 (N_73,In_570,In_10);
xnor U74 (N_74,In_254,In_669);
or U75 (N_75,In_830,In_17);
or U76 (N_76,In_216,In_662);
or U77 (N_77,In_928,In_706);
and U78 (N_78,In_974,In_753);
nor U79 (N_79,In_710,In_882);
xnor U80 (N_80,In_955,In_374);
xor U81 (N_81,In_735,In_471);
nor U82 (N_82,In_803,In_719);
and U83 (N_83,In_3,In_565);
or U84 (N_84,In_538,In_582);
xor U85 (N_85,In_906,In_239);
xor U86 (N_86,In_187,In_523);
or U87 (N_87,In_343,In_778);
or U88 (N_88,In_924,In_844);
xnor U89 (N_89,In_739,In_514);
nor U90 (N_90,In_597,In_744);
and U91 (N_91,In_831,In_956);
nor U92 (N_92,In_77,In_559);
and U93 (N_93,In_840,In_660);
and U94 (N_94,In_711,In_377);
or U95 (N_95,In_807,In_989);
xor U96 (N_96,In_880,In_506);
nand U97 (N_97,In_73,In_580);
xor U98 (N_98,In_247,In_742);
and U99 (N_99,In_659,In_288);
or U100 (N_100,In_438,In_261);
and U101 (N_101,In_522,In_654);
nand U102 (N_102,In_302,In_308);
and U103 (N_103,In_589,In_683);
or U104 (N_104,In_346,In_736);
or U105 (N_105,In_102,In_648);
and U106 (N_106,In_25,In_132);
or U107 (N_107,In_675,In_640);
nand U108 (N_108,In_472,In_413);
or U109 (N_109,In_392,In_391);
nor U110 (N_110,In_238,In_157);
nand U111 (N_111,In_895,In_250);
nand U112 (N_112,In_757,In_942);
or U113 (N_113,In_123,In_337);
and U114 (N_114,In_168,In_101);
or U115 (N_115,In_869,In_917);
and U116 (N_116,In_53,In_292);
nand U117 (N_117,In_972,In_685);
nand U118 (N_118,In_356,In_415);
nand U119 (N_119,In_585,In_821);
nand U120 (N_120,In_878,In_765);
or U121 (N_121,In_394,In_676);
nor U122 (N_122,In_130,In_84);
xnor U123 (N_123,In_702,In_899);
and U124 (N_124,In_362,In_966);
or U125 (N_125,In_832,In_816);
xnor U126 (N_126,In_520,In_606);
nand U127 (N_127,In_442,In_644);
or U128 (N_128,In_376,In_78);
xor U129 (N_129,In_625,In_327);
or U130 (N_130,In_64,In_647);
or U131 (N_131,In_38,In_533);
or U132 (N_132,In_379,In_843);
xor U133 (N_133,In_7,In_993);
nand U134 (N_134,In_331,In_387);
and U135 (N_135,In_593,In_2);
nor U136 (N_136,In_746,In_252);
or U137 (N_137,In_910,In_873);
nor U138 (N_138,In_902,In_290);
or U139 (N_139,In_709,In_99);
nand U140 (N_140,In_126,In_729);
or U141 (N_141,In_207,In_431);
nand U142 (N_142,In_501,In_371);
xnor U143 (N_143,In_713,In_965);
and U144 (N_144,In_354,In_732);
or U145 (N_145,In_58,In_776);
nor U146 (N_146,In_389,In_889);
nand U147 (N_147,In_511,In_240);
nor U148 (N_148,In_425,In_340);
or U149 (N_149,In_135,In_698);
and U150 (N_150,In_29,In_615);
xor U151 (N_151,In_963,In_51);
and U152 (N_152,In_310,In_264);
and U153 (N_153,In_473,In_951);
xnor U154 (N_154,In_169,In_518);
and U155 (N_155,In_900,In_118);
and U156 (N_156,In_74,In_634);
xnor U157 (N_157,In_34,In_201);
and U158 (N_158,In_233,In_797);
xnor U159 (N_159,In_549,In_891);
xor U160 (N_160,In_550,In_195);
and U161 (N_161,In_8,In_564);
and U162 (N_162,In_969,In_381);
or U163 (N_163,In_855,In_496);
or U164 (N_164,In_373,In_937);
nand U165 (N_165,In_351,In_603);
or U166 (N_166,In_115,In_877);
nand U167 (N_167,In_556,In_466);
or U168 (N_168,In_401,In_664);
nand U169 (N_169,In_631,In_971);
xor U170 (N_170,In_213,In_592);
and U171 (N_171,In_445,In_774);
nor U172 (N_172,In_227,In_892);
or U173 (N_173,In_777,In_52);
nand U174 (N_174,In_246,In_694);
and U175 (N_175,In_205,In_661);
and U176 (N_176,In_562,In_530);
xor U177 (N_177,In_587,In_15);
or U178 (N_178,In_267,In_336);
nor U179 (N_179,In_18,In_812);
nor U180 (N_180,In_791,In_846);
or U181 (N_181,In_865,In_265);
xnor U182 (N_182,In_172,In_919);
nand U183 (N_183,In_167,In_474);
xor U184 (N_184,In_111,In_650);
nor U185 (N_185,In_242,In_87);
or U186 (N_186,In_498,In_114);
xnor U187 (N_187,In_323,In_842);
or U188 (N_188,In_226,In_316);
and U189 (N_189,In_847,In_49);
and U190 (N_190,In_594,In_555);
nand U191 (N_191,In_574,In_845);
and U192 (N_192,In_867,In_70);
nor U193 (N_193,In_779,In_723);
and U194 (N_194,In_527,In_197);
or U195 (N_195,In_82,In_756);
xnor U196 (N_196,In_420,In_992);
nand U197 (N_197,In_962,In_361);
or U198 (N_198,In_674,In_700);
nor U199 (N_199,In_704,In_835);
nand U200 (N_200,In_321,In_65);
and U201 (N_201,In_360,In_176);
nor U202 (N_202,In_27,N_169);
or U203 (N_203,In_314,In_994);
and U204 (N_204,In_677,N_180);
nor U205 (N_205,N_136,N_3);
xor U206 (N_206,In_657,In_639);
nand U207 (N_207,In_16,In_519);
nand U208 (N_208,In_46,In_291);
nor U209 (N_209,In_949,In_224);
or U210 (N_210,N_143,In_165);
or U211 (N_211,In_509,In_253);
or U212 (N_212,In_98,In_544);
nor U213 (N_213,In_163,In_563);
nand U214 (N_214,In_754,N_195);
or U215 (N_215,In_93,N_119);
or U216 (N_216,In_769,In_188);
nand U217 (N_217,N_58,In_838);
xnor U218 (N_218,In_766,In_747);
xor U219 (N_219,In_486,N_186);
xor U220 (N_220,In_107,In_935);
and U221 (N_221,In_566,In_503);
or U222 (N_222,In_282,In_119);
nor U223 (N_223,In_287,In_930);
or U224 (N_224,In_100,In_324);
or U225 (N_225,In_738,In_673);
nor U226 (N_226,In_30,In_705);
and U227 (N_227,In_623,In_491);
and U228 (N_228,N_124,In_802);
nor U229 (N_229,In_526,In_546);
nor U230 (N_230,In_568,In_991);
and U231 (N_231,In_954,In_120);
xor U232 (N_232,N_17,In_457);
or U233 (N_233,In_572,In_689);
and U234 (N_234,In_651,In_870);
or U235 (N_235,In_733,In_973);
xnor U236 (N_236,N_116,In_607);
or U237 (N_237,In_231,In_787);
nor U238 (N_238,In_663,In_493);
nor U239 (N_239,In_192,In_785);
nand U240 (N_240,N_57,N_167);
or U241 (N_241,In_784,In_887);
or U242 (N_242,In_162,In_536);
nand U243 (N_243,In_976,In_449);
or U244 (N_244,In_145,In_96);
and U245 (N_245,In_596,In_978);
xor U246 (N_246,In_608,In_492);
or U247 (N_247,In_883,N_53);
or U248 (N_248,N_45,In_155);
or U249 (N_249,N_170,In_487);
nor U250 (N_250,In_652,In_913);
xnor U251 (N_251,In_911,In_958);
nor U252 (N_252,N_90,In_0);
and U253 (N_253,N_86,In_304);
xor U254 (N_254,In_577,N_22);
and U255 (N_255,In_551,In_137);
nor U256 (N_256,In_655,In_624);
nor U257 (N_257,In_278,In_745);
nand U258 (N_258,In_97,In_868);
and U259 (N_259,In_85,In_860);
nor U260 (N_260,In_626,In_103);
nand U261 (N_261,In_799,In_293);
nand U262 (N_262,In_69,In_357);
or U263 (N_263,In_110,In_271);
nor U264 (N_264,In_959,In_576);
nand U265 (N_265,N_72,In_241);
and U266 (N_266,In_981,In_453);
and U267 (N_267,In_859,In_862);
xnor U268 (N_268,N_41,N_85);
nand U269 (N_269,In_975,In_154);
and U270 (N_270,In_461,In_579);
nor U271 (N_271,N_112,In_179);
nor U272 (N_272,In_703,In_434);
and U273 (N_273,In_419,N_153);
and U274 (N_274,In_805,N_160);
and U275 (N_275,N_12,In_339);
xor U276 (N_276,In_517,N_26);
nand U277 (N_277,In_279,In_441);
or U278 (N_278,In_363,In_717);
or U279 (N_279,In_478,In_204);
and U280 (N_280,In_888,In_485);
nor U281 (N_281,In_149,N_62);
nand U282 (N_282,In_189,N_61);
and U283 (N_283,In_504,N_139);
nand U284 (N_284,In_153,N_49);
nand U285 (N_285,In_249,In_901);
or U286 (N_286,In_621,In_598);
and U287 (N_287,In_309,In_696);
and U288 (N_288,In_217,In_970);
nand U289 (N_289,In_708,N_89);
nor U290 (N_290,N_175,N_199);
and U291 (N_291,In_138,In_370);
and U292 (N_292,In_12,In_483);
or U293 (N_293,In_372,In_946);
xor U294 (N_294,In_228,N_113);
and U295 (N_295,N_105,In_482);
and U296 (N_296,In_405,In_795);
nand U297 (N_297,In_307,N_37);
or U298 (N_298,In_894,In_347);
or U299 (N_299,In_236,In_141);
nand U300 (N_300,N_88,N_0);
nand U301 (N_301,N_64,In_156);
nor U302 (N_302,N_68,In_404);
and U303 (N_303,In_637,In_824);
xor U304 (N_304,In_804,In_932);
xor U305 (N_305,N_184,In_116);
and U306 (N_306,N_43,In_407);
or U307 (N_307,In_800,In_43);
xnor U308 (N_308,In_682,In_512);
or U309 (N_309,In_915,In_850);
or U310 (N_310,In_643,In_281);
nand U311 (N_311,In_697,N_23);
nand U312 (N_312,In_251,In_358);
nor U313 (N_313,In_578,In_715);
xnor U314 (N_314,In_181,N_187);
xor U315 (N_315,In_76,In_211);
and U316 (N_316,In_418,In_725);
nor U317 (N_317,In_45,In_635);
xnor U318 (N_318,In_208,N_135);
or U319 (N_319,In_408,N_122);
xnor U320 (N_320,N_133,N_120);
xnor U321 (N_321,In_908,N_35);
and U322 (N_322,N_188,In_871);
or U323 (N_323,In_166,In_881);
nand U324 (N_324,N_141,In_410);
or U325 (N_325,In_257,N_87);
nand U326 (N_326,In_244,In_945);
nand U327 (N_327,N_157,N_185);
nand U328 (N_328,In_569,In_641);
and U329 (N_329,In_819,N_163);
or U330 (N_330,In_272,In_366);
nand U331 (N_331,In_128,In_400);
nand U332 (N_332,In_737,N_193);
xnor U333 (N_333,In_385,In_311);
nor U334 (N_334,In_633,In_40);
or U335 (N_335,In_961,In_319);
and U336 (N_336,In_37,In_583);
or U337 (N_337,In_333,In_667);
xor U338 (N_338,N_178,In_416);
and U339 (N_339,In_368,In_488);
and U340 (N_340,In_601,In_59);
nand U341 (N_341,In_929,In_548);
or U342 (N_342,In_209,In_460);
nand U343 (N_343,In_658,In_313);
nor U344 (N_344,In_758,In_620);
nand U345 (N_345,N_155,In_720);
or U346 (N_346,N_125,In_79);
nand U347 (N_347,N_106,In_604);
xor U348 (N_348,In_191,N_118);
and U349 (N_349,In_61,N_137);
xnor U350 (N_350,N_50,In_378);
nand U351 (N_351,N_31,In_535);
and U352 (N_352,In_768,N_161);
nand U353 (N_353,In_849,In_263);
and U354 (N_354,In_837,In_595);
or U355 (N_355,N_93,In_276);
nor U356 (N_356,In_874,In_818);
nor U357 (N_357,In_382,In_225);
nand U358 (N_358,In_616,In_193);
nor U359 (N_359,In_575,In_513);
nand U360 (N_360,N_171,In_380);
xor U361 (N_361,In_730,In_383);
nand U362 (N_362,In_50,In_646);
xor U363 (N_363,N_39,N_32);
or U364 (N_364,In_853,N_168);
xor U365 (N_365,In_275,In_489);
nor U366 (N_366,N_9,N_140);
and U367 (N_367,In_749,N_151);
xnor U368 (N_368,In_350,In_124);
or U369 (N_369,In_429,In_731);
nand U370 (N_370,In_299,In_605);
or U371 (N_371,In_322,In_500);
nor U372 (N_372,N_10,In_560);
xor U373 (N_373,In_35,N_38);
nor U374 (N_374,In_508,In_428);
nand U375 (N_375,In_875,In_760);
nand U376 (N_376,In_136,In_335);
or U377 (N_377,N_129,In_537);
nand U378 (N_378,In_543,N_28);
and U379 (N_379,In_48,In_220);
xor U380 (N_380,N_63,In_545);
or U381 (N_381,In_440,In_121);
or U382 (N_382,N_145,In_306);
nand U383 (N_383,In_841,N_29);
and U384 (N_384,In_237,In_836);
and U385 (N_385,N_131,In_490);
nor U386 (N_386,In_848,In_67);
xor U387 (N_387,In_127,In_811);
xor U388 (N_388,In_348,N_4);
or U389 (N_389,N_148,In_414);
nor U390 (N_390,In_558,N_71);
nor U391 (N_391,In_763,In_105);
or U392 (N_392,In_89,N_198);
nand U393 (N_393,In_399,In_588);
nor U394 (N_394,In_701,In_817);
and U395 (N_395,N_20,N_14);
or U396 (N_396,N_162,In_934);
or U397 (N_397,In_11,In_829);
xnor U398 (N_398,In_469,In_14);
nand U399 (N_399,In_266,In_55);
or U400 (N_400,In_611,In_180);
and U401 (N_401,N_210,In_171);
xor U402 (N_402,In_947,In_967);
nor U403 (N_403,N_245,In_557);
xor U404 (N_404,In_941,N_204);
nand U405 (N_405,In_258,N_268);
xor U406 (N_406,In_628,In_36);
nand U407 (N_407,N_275,In_147);
and U408 (N_408,N_381,In_903);
nor U409 (N_409,In_210,N_292);
and U410 (N_410,N_375,In_561);
nor U411 (N_411,N_36,In_699);
nand U412 (N_412,In_57,In_502);
xnor U413 (N_413,N_44,In_143);
or U414 (N_414,In_386,In_539);
xnor U415 (N_415,N_386,In_444);
or U416 (N_416,In_134,In_32);
or U417 (N_417,In_54,N_363);
or U418 (N_418,N_310,In_983);
or U419 (N_419,In_91,In_759);
or U420 (N_420,N_285,N_261);
xnor U421 (N_421,In_479,In_295);
or U422 (N_422,N_102,In_781);
xor U423 (N_423,In_235,In_430);
and U424 (N_424,In_325,In_613);
and U425 (N_425,In_367,In_447);
nor U426 (N_426,N_304,N_279);
nand U427 (N_427,In_748,In_232);
xor U428 (N_428,In_997,In_198);
or U429 (N_429,N_230,N_321);
and U430 (N_430,In_609,N_387);
and U431 (N_431,N_114,In_668);
nand U432 (N_432,In_712,N_257);
nor U433 (N_433,In_707,In_355);
nor U434 (N_434,N_266,N_130);
xor U435 (N_435,In_170,N_60);
xor U436 (N_436,N_296,N_225);
or U437 (N_437,N_344,In_780);
nand U438 (N_438,N_108,In_734);
or U439 (N_439,In_995,In_480);
or U440 (N_440,In_670,N_297);
nor U441 (N_441,N_356,N_206);
nand U442 (N_442,N_132,N_336);
and U443 (N_443,In_393,N_391);
nand U444 (N_444,In_693,In_775);
and U445 (N_445,N_150,In_390);
nor U446 (N_446,N_330,N_121);
or U447 (N_447,In_638,N_329);
xnor U448 (N_448,In_301,In_117);
and U449 (N_449,N_367,N_281);
nor U450 (N_450,N_227,In_790);
or U451 (N_451,In_412,In_83);
and U452 (N_452,N_115,N_360);
nand U453 (N_453,In_369,In_183);
and U454 (N_454,In_56,In_980);
and U455 (N_455,N_191,N_5);
and U456 (N_456,In_532,In_984);
nor U457 (N_457,N_27,In_822);
xnor U458 (N_458,In_270,N_364);
or U459 (N_459,In_219,N_397);
or U460 (N_460,N_318,In_199);
nand U461 (N_461,N_394,In_19);
and U462 (N_462,In_653,N_197);
nand U463 (N_463,N_107,N_368);
xor U464 (N_464,In_436,N_214);
nor U465 (N_465,N_189,N_181);
or U466 (N_466,In_688,N_383);
nor U467 (N_467,N_276,N_104);
nor U468 (N_468,N_332,In_495);
and U469 (N_469,N_253,N_79);
nor U470 (N_470,N_389,In_547);
and U471 (N_471,In_459,N_399);
nand U472 (N_472,N_333,In_402);
or U473 (N_473,In_636,In_728);
nor U474 (N_474,N_277,In_541);
and U475 (N_475,N_235,N_248);
and U476 (N_476,In_964,N_220);
and U477 (N_477,N_390,In_451);
nand U478 (N_478,N_208,In_827);
nor U479 (N_479,In_68,In_534);
nor U480 (N_480,In_150,N_215);
or U481 (N_481,In_212,In_33);
xor U482 (N_482,In_320,N_305);
nor U483 (N_483,In_139,In_72);
or U484 (N_484,In_248,N_357);
xor U485 (N_485,In_798,N_325);
nor U486 (N_486,N_270,In_826);
or U487 (N_487,N_369,N_34);
or U488 (N_488,N_341,N_19);
xor U489 (N_489,N_73,N_237);
nand U490 (N_490,In_926,In_602);
xnor U491 (N_491,N_324,In_66);
or U492 (N_492,N_289,N_40);
nor U493 (N_493,N_94,In_554);
xnor U494 (N_494,In_612,N_379);
nor U495 (N_495,In_524,N_252);
xnor U496 (N_496,In_510,N_372);
or U497 (N_497,In_125,N_349);
nor U498 (N_498,In_904,N_350);
nand U499 (N_499,N_144,In_131);
nor U500 (N_500,In_814,In_182);
nand U501 (N_501,In_88,N_174);
or U502 (N_502,N_345,N_373);
nand U503 (N_503,In_681,In_552);
nand U504 (N_504,N_316,In_221);
and U505 (N_505,In_828,In_716);
nor U506 (N_506,N_59,In_200);
and U507 (N_507,In_890,In_481);
or U508 (N_508,N_219,N_211);
xor U509 (N_509,N_142,N_398);
or U510 (N_510,N_339,N_343);
nor U511 (N_511,N_322,N_30);
nor U512 (N_512,N_250,N_282);
xnor U513 (N_513,In_458,In_259);
nand U514 (N_514,N_286,N_205);
nand U515 (N_515,N_393,N_66);
nor U516 (N_516,In_315,N_384);
and U517 (N_517,In_294,N_177);
xor U518 (N_518,N_103,In_943);
nor U519 (N_519,N_111,In_173);
xnor U520 (N_520,N_16,In_21);
xnor U521 (N_521,In_297,In_866);
or U522 (N_522,In_755,N_154);
xor U523 (N_523,In_24,N_238);
or U524 (N_524,In_692,N_242);
xnor U525 (N_525,N_239,In_678);
or U526 (N_526,N_272,In_122);
or U527 (N_527,N_91,N_265);
and U528 (N_528,N_280,In_750);
and U529 (N_529,N_300,In_280);
xor U530 (N_530,N_337,N_11);
nor U531 (N_531,In_825,N_224);
xor U532 (N_532,In_345,N_6);
or U533 (N_533,In_788,In_448);
and U534 (N_534,N_320,In_396);
xor U535 (N_535,In_856,N_351);
or U536 (N_536,In_542,N_361);
xnor U537 (N_537,In_289,In_218);
or U538 (N_538,N_84,In_857);
or U539 (N_539,In_4,N_366);
nand U540 (N_540,N_251,In_645);
or U541 (N_541,N_75,In_245);
and U542 (N_542,In_914,N_346);
xnor U543 (N_543,N_236,In_839);
and U544 (N_544,In_334,N_274);
xnor U545 (N_545,N_200,In_433);
and U546 (N_546,In_905,N_98);
or U547 (N_547,In_146,N_331);
nand U548 (N_548,In_987,N_221);
xor U549 (N_549,N_326,N_247);
or U550 (N_550,N_212,In_721);
xor U551 (N_551,N_48,In_177);
or U552 (N_552,In_317,In_223);
or U553 (N_553,N_149,N_376);
and U554 (N_554,N_291,N_258);
and U555 (N_555,In_852,In_312);
and U556 (N_556,N_70,N_317);
xnor U557 (N_557,N_288,N_342);
and U558 (N_558,N_352,In_960);
and U559 (N_559,In_229,N_335);
xor U560 (N_560,In_13,In_672);
nor U561 (N_561,In_151,In_20);
or U562 (N_562,In_41,N_158);
nand U563 (N_563,N_2,N_232);
nor U564 (N_564,In_772,N_359);
nor U565 (N_565,N_159,In_794);
xor U566 (N_566,In_953,In_395);
or U567 (N_567,In_497,In_160);
nand U568 (N_568,N_298,N_82);
nand U569 (N_569,N_92,In_359);
xnor U570 (N_570,N_314,N_126);
or U571 (N_571,N_234,N_301);
and U572 (N_572,N_52,N_217);
and U573 (N_573,In_424,N_99);
xnor U574 (N_574,In_985,In_764);
nand U575 (N_575,In_529,N_382);
or U576 (N_576,In_863,In_349);
nand U577 (N_577,N_110,In_284);
xnor U578 (N_578,N_269,N_340);
and U579 (N_579,N_354,N_392);
or U580 (N_580,N_147,N_311);
nand U581 (N_581,N_284,N_378);
or U582 (N_582,N_213,In_92);
xnor U583 (N_583,N_134,N_176);
xor U584 (N_584,In_793,In_365);
and U585 (N_585,N_55,In_432);
xnor U586 (N_586,In_230,In_435);
xor U587 (N_587,N_319,In_463);
nor U588 (N_588,N_18,N_377);
xor U589 (N_589,In_42,N_260);
nand U590 (N_590,N_202,In_786);
nor U591 (N_591,In_397,N_183);
or U592 (N_592,In_499,N_179);
xnor U593 (N_593,N_80,In_614);
xnor U594 (N_594,In_215,N_388);
nand U595 (N_595,N_228,N_255);
xor U596 (N_596,In_417,In_214);
nand U597 (N_597,N_209,In_920);
nor U598 (N_598,N_81,N_15);
or U599 (N_599,N_334,N_309);
or U600 (N_600,In_789,N_567);
nor U601 (N_601,N_65,N_444);
or U602 (N_602,N_430,N_509);
xor U603 (N_603,In_384,N_484);
and U604 (N_604,N_489,N_487);
nor U605 (N_605,N_582,In_952);
or U606 (N_606,N_313,N_417);
nor U607 (N_607,In_161,N_42);
xnor U608 (N_608,N_194,N_540);
nand U609 (N_609,N_517,N_164);
nor U610 (N_610,N_433,In_918);
or U611 (N_611,N_464,N_299);
xnor U612 (N_612,N_467,N_485);
nand U613 (N_613,N_222,N_401);
or U614 (N_614,N_515,N_374);
xor U615 (N_615,N_207,N_422);
and U616 (N_616,N_457,N_428);
nor U617 (N_617,In_439,N_506);
nor U618 (N_618,N_592,N_264);
xnor U619 (N_619,In_998,N_462);
nor U620 (N_620,In_921,In_938);
or U621 (N_621,In_515,In_833);
or U622 (N_622,In_427,N_499);
nand U623 (N_623,N_568,N_166);
or U624 (N_624,N_495,N_165);
xor U625 (N_625,N_408,N_138);
xnor U626 (N_626,N_271,N_460);
and U627 (N_627,In_823,N_295);
xor U628 (N_628,N_461,In_158);
or U629 (N_629,N_290,N_480);
or U630 (N_630,N_283,N_564);
or U631 (N_631,In_437,N_293);
nand U632 (N_632,N_543,In_222);
and U633 (N_633,N_454,N_231);
xnor U634 (N_634,N_596,N_481);
xnor U635 (N_635,N_501,N_524);
nor U636 (N_636,In_129,N_76);
or U637 (N_637,N_246,N_51);
nor U638 (N_638,N_598,N_463);
nand U639 (N_639,N_404,N_557);
nor U640 (N_640,N_445,N_554);
nand U641 (N_641,N_533,N_565);
xor U642 (N_642,N_553,In_990);
nand U643 (N_643,N_312,N_503);
nor U644 (N_644,N_24,N_262);
and U645 (N_645,In_422,N_423);
or U646 (N_646,In_303,N_256);
nand U647 (N_647,N_323,N_406);
nor U648 (N_648,N_450,N_405);
and U649 (N_649,N_385,In_528);
nor U650 (N_650,N_581,In_353);
nand U651 (N_651,N_196,N_496);
xor U652 (N_652,N_407,In_684);
or U653 (N_653,N_465,N_522);
or U654 (N_654,N_69,N_441);
or U655 (N_655,N_528,N_584);
xnor U656 (N_656,N_371,In_996);
or U657 (N_657,In_909,N_590);
or U658 (N_658,In_81,In_159);
or U659 (N_659,N_512,N_365);
xnor U660 (N_660,In_912,N_419);
nand U661 (N_661,In_342,In_695);
nor U662 (N_662,N_446,N_491);
nor U663 (N_663,N_67,N_527);
or U664 (N_664,N_513,In_726);
nor U665 (N_665,N_532,N_100);
nand U666 (N_666,N_152,In_834);
xor U667 (N_667,N_451,N_396);
or U668 (N_668,N_558,In_505);
nor U669 (N_669,N_477,In_722);
nor U670 (N_670,N_498,N_74);
xor U671 (N_671,N_420,N_249);
nor U672 (N_672,N_573,N_229);
and U673 (N_673,N_595,N_358);
xor U674 (N_674,N_287,In_813);
xor U675 (N_675,N_478,N_443);
and U676 (N_676,N_504,N_431);
or U677 (N_677,In_999,In_9);
or U678 (N_678,In_5,N_347);
or U679 (N_679,N_555,N_545);
nor U680 (N_680,N_46,N_471);
nand U681 (N_681,N_439,N_482);
nor U682 (N_682,N_294,N_117);
xor U683 (N_683,N_559,N_33);
xnor U684 (N_684,N_437,N_534);
xor U685 (N_685,N_556,In_507);
or U686 (N_686,In_133,In_352);
nor U687 (N_687,In_610,N_473);
nor U688 (N_688,N_505,In_260);
nor U689 (N_689,N_580,N_440);
or U690 (N_690,N_327,N_458);
or U691 (N_691,N_529,N_490);
nor U692 (N_692,N_583,N_54);
nor U693 (N_693,N_432,N_267);
nand U694 (N_694,N_442,In_770);
xor U695 (N_695,N_526,N_427);
xor U696 (N_696,In_923,In_22);
xnor U697 (N_697,N_146,In_581);
and U698 (N_698,N_78,N_599);
xor U699 (N_699,N_475,N_438);
xor U700 (N_700,N_552,N_476);
xor U701 (N_701,N_576,In_464);
nor U702 (N_702,N_338,N_127);
nand U703 (N_703,N_412,N_560);
nand U704 (N_704,N_566,N_469);
xnor U705 (N_705,N_410,N_572);
or U706 (N_706,N_508,N_192);
xor U707 (N_707,N_418,N_578);
and U708 (N_708,N_25,N_8);
and U709 (N_709,N_518,N_273);
and U710 (N_710,N_426,In_470);
nand U711 (N_711,N_470,N_353);
nor U712 (N_712,N_13,N_561);
nor U713 (N_713,N_546,N_453);
or U714 (N_714,N_83,N_307);
nand U715 (N_715,N_424,N_570);
nor U716 (N_716,In_285,N_537);
and U717 (N_717,N_216,N_486);
xnor U718 (N_718,In_1,In_274);
xnor U719 (N_719,In_743,N_571);
nand U720 (N_720,N_551,N_594);
or U721 (N_721,N_173,N_243);
xor U722 (N_722,N_411,N_579);
and U723 (N_723,In_26,N_452);
or U724 (N_724,N_519,N_577);
and U725 (N_725,In_47,N_409);
xnor U726 (N_726,N_574,N_308);
xor U727 (N_727,N_400,N_541);
nor U728 (N_728,N_539,N_362);
and U729 (N_729,N_494,In_467);
xor U730 (N_730,N_587,N_259);
or U731 (N_731,N_414,N_535);
nand U732 (N_732,N_456,In_421);
xnor U733 (N_733,N_586,In_687);
nand U734 (N_734,N_593,N_355);
or U735 (N_735,N_492,In_175);
nor U736 (N_736,N_123,N_514);
nand U737 (N_737,N_497,In_584);
nor U738 (N_738,N_223,N_455);
xor U739 (N_739,N_483,N_575);
and U740 (N_740,N_525,N_523);
nand U741 (N_741,In_243,N_536);
and U742 (N_742,N_370,N_95);
xnor U743 (N_743,N_436,In_286);
nand U744 (N_744,In_184,N_302);
xnor U745 (N_745,N_328,N_507);
and U746 (N_746,N_97,N_591);
nand U747 (N_747,N_395,N_226);
nand U748 (N_748,In_338,In_691);
xor U749 (N_749,N_562,N_550);
or U750 (N_750,N_172,N_500);
xor U751 (N_751,N_348,N_402);
nor U752 (N_752,N_7,N_474);
xnor U753 (N_753,N_241,In_475);
or U754 (N_754,In_936,N_109);
xnor U755 (N_755,N_96,N_569);
nor U756 (N_756,N_429,In_630);
xnor U757 (N_757,In_283,N_240);
and U758 (N_758,N_597,N_233);
nand U759 (N_759,N_201,N_547);
or U760 (N_760,In_28,N_520);
or U761 (N_761,N_538,N_413);
or U762 (N_762,In_782,N_77);
nand U763 (N_763,In_815,N_435);
xor U764 (N_764,N_306,N_278);
nand U765 (N_765,In_896,N_263);
nor U766 (N_766,In_885,N_421);
xor U767 (N_767,In_679,N_425);
xnor U768 (N_768,N_511,N_101);
xnor U769 (N_769,In_861,In_298);
nor U770 (N_770,N_47,In_666);
or U771 (N_771,N_190,N_493);
nand U772 (N_772,N_472,N_563);
nor U773 (N_773,N_218,In_234);
or U774 (N_774,N_203,N_588);
nand U775 (N_775,N_521,N_531);
nor U776 (N_776,In_328,N_488);
and U777 (N_777,In_300,N_468);
and U778 (N_778,N_434,N_1);
nor U779 (N_779,In_364,N_447);
xor U780 (N_780,N_449,N_182);
nor U781 (N_781,N_315,N_303);
xor U782 (N_782,N_585,In_196);
or U783 (N_783,N_544,N_502);
nor U784 (N_784,N_530,N_416);
and U785 (N_785,N_466,N_21);
or U786 (N_786,In_977,N_254);
nand U787 (N_787,N_56,In_332);
or U788 (N_788,In_31,N_415);
nor U789 (N_789,N_156,N_549);
and U790 (N_790,N_244,N_459);
nor U791 (N_791,N_542,N_548);
or U792 (N_792,N_516,N_128);
and U793 (N_793,In_455,In_108);
and U794 (N_794,In_884,In_411);
nor U795 (N_795,In_94,In_268);
or U796 (N_796,N_510,N_403);
nand U797 (N_797,N_589,In_406);
nor U798 (N_798,N_479,N_448);
or U799 (N_799,In_203,N_380);
nor U800 (N_800,N_640,N_735);
nor U801 (N_801,N_742,N_621);
nor U802 (N_802,N_762,N_789);
xor U803 (N_803,N_715,N_603);
nand U804 (N_804,N_708,N_688);
nor U805 (N_805,N_639,N_738);
nor U806 (N_806,N_689,N_709);
nand U807 (N_807,N_772,N_630);
and U808 (N_808,N_756,N_788);
and U809 (N_809,N_623,N_669);
nor U810 (N_810,N_635,N_707);
or U811 (N_811,N_729,N_695);
and U812 (N_812,N_720,N_607);
or U813 (N_813,N_684,N_677);
xor U814 (N_814,N_636,N_693);
or U815 (N_815,N_612,N_725);
xnor U816 (N_816,N_653,N_629);
nand U817 (N_817,N_681,N_671);
xor U818 (N_818,N_701,N_786);
xor U819 (N_819,N_631,N_744);
and U820 (N_820,N_615,N_652);
and U821 (N_821,N_647,N_705);
and U822 (N_822,N_773,N_604);
nor U823 (N_823,N_672,N_664);
nor U824 (N_824,N_643,N_673);
nor U825 (N_825,N_782,N_609);
nor U826 (N_826,N_732,N_627);
and U827 (N_827,N_678,N_722);
or U828 (N_828,N_764,N_601);
xor U829 (N_829,N_700,N_702);
and U830 (N_830,N_711,N_641);
nor U831 (N_831,N_608,N_675);
xor U832 (N_832,N_775,N_765);
nor U833 (N_833,N_686,N_622);
or U834 (N_834,N_763,N_799);
nor U835 (N_835,N_710,N_787);
nand U836 (N_836,N_713,N_645);
nor U837 (N_837,N_637,N_613);
and U838 (N_838,N_600,N_611);
nand U839 (N_839,N_747,N_741);
nand U840 (N_840,N_749,N_646);
or U841 (N_841,N_644,N_634);
or U842 (N_842,N_650,N_661);
xor U843 (N_843,N_724,N_794);
xnor U844 (N_844,N_687,N_795);
or U845 (N_845,N_758,N_654);
xnor U846 (N_846,N_751,N_679);
xnor U847 (N_847,N_798,N_614);
or U848 (N_848,N_760,N_655);
and U849 (N_849,N_676,N_670);
nor U850 (N_850,N_698,N_781);
and U851 (N_851,N_696,N_649);
nor U852 (N_852,N_659,N_752);
nand U853 (N_853,N_754,N_726);
nor U854 (N_854,N_626,N_727);
and U855 (N_855,N_750,N_737);
or U856 (N_856,N_616,N_721);
nand U857 (N_857,N_777,N_784);
nor U858 (N_858,N_716,N_605);
nor U859 (N_859,N_680,N_719);
xnor U860 (N_860,N_642,N_620);
xnor U861 (N_861,N_663,N_667);
nand U862 (N_862,N_731,N_779);
or U863 (N_863,N_674,N_769);
nand U864 (N_864,N_692,N_718);
nand U865 (N_865,N_704,N_699);
and U866 (N_866,N_743,N_797);
and U867 (N_867,N_791,N_624);
xnor U868 (N_868,N_761,N_657);
xor U869 (N_869,N_619,N_768);
nand U870 (N_870,N_618,N_771);
nor U871 (N_871,N_723,N_628);
xnor U872 (N_872,N_660,N_753);
nand U873 (N_873,N_691,N_685);
nand U874 (N_874,N_717,N_730);
nor U875 (N_875,N_739,N_682);
nand U876 (N_876,N_666,N_774);
or U877 (N_877,N_759,N_662);
or U878 (N_878,N_755,N_712);
or U879 (N_879,N_778,N_656);
or U880 (N_880,N_740,N_703);
nor U881 (N_881,N_648,N_748);
nor U882 (N_882,N_697,N_736);
xor U883 (N_883,N_632,N_638);
and U884 (N_884,N_767,N_746);
nor U885 (N_885,N_683,N_706);
and U886 (N_886,N_668,N_796);
nor U887 (N_887,N_658,N_745);
xnor U888 (N_888,N_633,N_792);
xor U889 (N_889,N_766,N_651);
or U890 (N_890,N_728,N_606);
xor U891 (N_891,N_780,N_610);
or U892 (N_892,N_757,N_625);
and U893 (N_893,N_617,N_690);
nor U894 (N_894,N_783,N_793);
and U895 (N_895,N_776,N_734);
or U896 (N_896,N_714,N_770);
or U897 (N_897,N_665,N_733);
or U898 (N_898,N_694,N_785);
nor U899 (N_899,N_602,N_790);
or U900 (N_900,N_766,N_676);
or U901 (N_901,N_761,N_731);
xnor U902 (N_902,N_756,N_768);
xor U903 (N_903,N_664,N_728);
nor U904 (N_904,N_677,N_607);
xnor U905 (N_905,N_694,N_620);
xnor U906 (N_906,N_679,N_736);
nor U907 (N_907,N_765,N_799);
xor U908 (N_908,N_682,N_643);
nor U909 (N_909,N_686,N_621);
or U910 (N_910,N_652,N_618);
xor U911 (N_911,N_604,N_737);
nor U912 (N_912,N_676,N_689);
and U913 (N_913,N_775,N_715);
and U914 (N_914,N_672,N_680);
nor U915 (N_915,N_689,N_751);
or U916 (N_916,N_690,N_747);
xor U917 (N_917,N_773,N_742);
and U918 (N_918,N_782,N_722);
xor U919 (N_919,N_683,N_676);
nand U920 (N_920,N_768,N_765);
and U921 (N_921,N_717,N_735);
and U922 (N_922,N_671,N_692);
and U923 (N_923,N_714,N_697);
nand U924 (N_924,N_653,N_767);
and U925 (N_925,N_642,N_680);
nand U926 (N_926,N_628,N_780);
nor U927 (N_927,N_720,N_647);
and U928 (N_928,N_700,N_753);
nor U929 (N_929,N_656,N_781);
nor U930 (N_930,N_637,N_649);
and U931 (N_931,N_695,N_605);
or U932 (N_932,N_612,N_781);
or U933 (N_933,N_607,N_622);
or U934 (N_934,N_713,N_629);
or U935 (N_935,N_789,N_698);
nand U936 (N_936,N_698,N_759);
and U937 (N_937,N_775,N_778);
nor U938 (N_938,N_751,N_617);
nor U939 (N_939,N_724,N_766);
nor U940 (N_940,N_707,N_607);
nand U941 (N_941,N_626,N_657);
nand U942 (N_942,N_693,N_726);
nand U943 (N_943,N_752,N_747);
nor U944 (N_944,N_626,N_606);
xor U945 (N_945,N_732,N_784);
or U946 (N_946,N_618,N_766);
xnor U947 (N_947,N_789,N_671);
or U948 (N_948,N_627,N_770);
and U949 (N_949,N_779,N_686);
and U950 (N_950,N_602,N_619);
xnor U951 (N_951,N_621,N_756);
nor U952 (N_952,N_665,N_638);
nand U953 (N_953,N_697,N_636);
and U954 (N_954,N_754,N_617);
nor U955 (N_955,N_620,N_677);
xnor U956 (N_956,N_668,N_603);
and U957 (N_957,N_687,N_657);
nor U958 (N_958,N_668,N_604);
and U959 (N_959,N_738,N_768);
xor U960 (N_960,N_625,N_663);
and U961 (N_961,N_694,N_615);
nor U962 (N_962,N_603,N_616);
and U963 (N_963,N_627,N_667);
nand U964 (N_964,N_652,N_701);
and U965 (N_965,N_647,N_773);
and U966 (N_966,N_753,N_621);
or U967 (N_967,N_642,N_755);
and U968 (N_968,N_799,N_650);
and U969 (N_969,N_727,N_600);
nand U970 (N_970,N_607,N_632);
xnor U971 (N_971,N_728,N_662);
nor U972 (N_972,N_790,N_735);
or U973 (N_973,N_792,N_771);
xor U974 (N_974,N_690,N_771);
or U975 (N_975,N_763,N_735);
xnor U976 (N_976,N_704,N_767);
nand U977 (N_977,N_673,N_702);
or U978 (N_978,N_689,N_777);
or U979 (N_979,N_611,N_637);
nor U980 (N_980,N_623,N_693);
and U981 (N_981,N_646,N_674);
or U982 (N_982,N_616,N_690);
xor U983 (N_983,N_783,N_635);
nand U984 (N_984,N_787,N_619);
or U985 (N_985,N_609,N_620);
nand U986 (N_986,N_670,N_651);
nand U987 (N_987,N_754,N_737);
xor U988 (N_988,N_617,N_667);
nor U989 (N_989,N_726,N_781);
nand U990 (N_990,N_756,N_778);
and U991 (N_991,N_696,N_629);
or U992 (N_992,N_636,N_725);
nand U993 (N_993,N_730,N_684);
and U994 (N_994,N_743,N_772);
xor U995 (N_995,N_646,N_630);
xnor U996 (N_996,N_733,N_636);
nor U997 (N_997,N_659,N_672);
nand U998 (N_998,N_694,N_633);
nand U999 (N_999,N_769,N_646);
nor U1000 (N_1000,N_975,N_982);
or U1001 (N_1001,N_961,N_916);
nor U1002 (N_1002,N_991,N_819);
nor U1003 (N_1003,N_840,N_863);
and U1004 (N_1004,N_940,N_918);
or U1005 (N_1005,N_892,N_854);
or U1006 (N_1006,N_905,N_915);
nand U1007 (N_1007,N_953,N_837);
nor U1008 (N_1008,N_936,N_999);
and U1009 (N_1009,N_812,N_862);
nor U1010 (N_1010,N_979,N_985);
xor U1011 (N_1011,N_954,N_907);
or U1012 (N_1012,N_908,N_852);
and U1013 (N_1013,N_869,N_900);
xnor U1014 (N_1014,N_951,N_996);
nor U1015 (N_1015,N_993,N_899);
xnor U1016 (N_1016,N_844,N_963);
or U1017 (N_1017,N_937,N_807);
nand U1018 (N_1018,N_945,N_893);
xor U1019 (N_1019,N_864,N_952);
xor U1020 (N_1020,N_926,N_972);
nor U1021 (N_1021,N_947,N_986);
or U1022 (N_1022,N_824,N_828);
nand U1023 (N_1023,N_883,N_948);
and U1024 (N_1024,N_888,N_811);
nor U1025 (N_1025,N_998,N_830);
xnor U1026 (N_1026,N_970,N_962);
nand U1027 (N_1027,N_849,N_873);
xor U1028 (N_1028,N_988,N_942);
nand U1029 (N_1029,N_813,N_827);
xor U1030 (N_1030,N_805,N_867);
and U1031 (N_1031,N_987,N_842);
or U1032 (N_1032,N_941,N_974);
nor U1033 (N_1033,N_959,N_990);
and U1034 (N_1034,N_898,N_885);
nor U1035 (N_1035,N_914,N_816);
or U1036 (N_1036,N_834,N_902);
xor U1037 (N_1037,N_847,N_976);
or U1038 (N_1038,N_801,N_901);
nand U1039 (N_1039,N_833,N_946);
or U1040 (N_1040,N_804,N_971);
and U1041 (N_1041,N_957,N_871);
or U1042 (N_1042,N_821,N_823);
nand U1043 (N_1043,N_835,N_968);
xnor U1044 (N_1044,N_956,N_890);
nor U1045 (N_1045,N_853,N_876);
xor U1046 (N_1046,N_960,N_910);
and U1047 (N_1047,N_992,N_882);
and U1048 (N_1048,N_904,N_989);
nand U1049 (N_1049,N_906,N_860);
or U1050 (N_1050,N_930,N_995);
nor U1051 (N_1051,N_843,N_955);
and U1052 (N_1052,N_870,N_866);
or U1053 (N_1053,N_950,N_938);
xnor U1054 (N_1054,N_881,N_848);
nand U1055 (N_1055,N_856,N_829);
xnor U1056 (N_1056,N_809,N_994);
nand U1057 (N_1057,N_943,N_822);
xnor U1058 (N_1058,N_980,N_978);
or U1059 (N_1059,N_949,N_879);
xnor U1060 (N_1060,N_832,N_920);
and U1061 (N_1061,N_855,N_912);
xnor U1062 (N_1062,N_984,N_923);
nand U1063 (N_1063,N_927,N_934);
nor U1064 (N_1064,N_818,N_838);
or U1065 (N_1065,N_969,N_831);
and U1066 (N_1066,N_880,N_977);
or U1067 (N_1067,N_958,N_868);
or U1068 (N_1068,N_846,N_889);
nand U1069 (N_1069,N_932,N_894);
and U1070 (N_1070,N_886,N_913);
xor U1071 (N_1071,N_933,N_967);
and U1072 (N_1072,N_983,N_817);
or U1073 (N_1073,N_814,N_925);
nand U1074 (N_1074,N_878,N_825);
nor U1075 (N_1075,N_973,N_851);
xnor U1076 (N_1076,N_891,N_808);
nand U1077 (N_1077,N_931,N_929);
nor U1078 (N_1078,N_865,N_858);
or U1079 (N_1079,N_820,N_841);
nand U1080 (N_1080,N_826,N_895);
xnor U1081 (N_1081,N_810,N_935);
xnor U1082 (N_1082,N_921,N_965);
and U1083 (N_1083,N_877,N_981);
xnor U1084 (N_1084,N_845,N_997);
nor U1085 (N_1085,N_806,N_861);
xor U1086 (N_1086,N_966,N_839);
nand U1087 (N_1087,N_815,N_802);
nor U1088 (N_1088,N_872,N_850);
nand U1089 (N_1089,N_884,N_896);
nor U1090 (N_1090,N_875,N_897);
or U1091 (N_1091,N_909,N_919);
and U1092 (N_1092,N_939,N_887);
nor U1093 (N_1093,N_857,N_944);
and U1094 (N_1094,N_924,N_800);
nor U1095 (N_1095,N_803,N_917);
nand U1096 (N_1096,N_964,N_922);
nor U1097 (N_1097,N_836,N_874);
and U1098 (N_1098,N_911,N_928);
and U1099 (N_1099,N_903,N_859);
or U1100 (N_1100,N_860,N_949);
xnor U1101 (N_1101,N_876,N_825);
xor U1102 (N_1102,N_972,N_867);
nor U1103 (N_1103,N_903,N_845);
nand U1104 (N_1104,N_975,N_927);
and U1105 (N_1105,N_828,N_904);
xnor U1106 (N_1106,N_893,N_927);
or U1107 (N_1107,N_950,N_956);
nor U1108 (N_1108,N_980,N_890);
nor U1109 (N_1109,N_891,N_875);
and U1110 (N_1110,N_999,N_838);
xor U1111 (N_1111,N_903,N_945);
xor U1112 (N_1112,N_943,N_899);
or U1113 (N_1113,N_906,N_921);
xnor U1114 (N_1114,N_998,N_984);
xnor U1115 (N_1115,N_929,N_841);
xnor U1116 (N_1116,N_983,N_953);
or U1117 (N_1117,N_941,N_971);
nand U1118 (N_1118,N_983,N_841);
xor U1119 (N_1119,N_807,N_942);
and U1120 (N_1120,N_962,N_833);
and U1121 (N_1121,N_888,N_832);
and U1122 (N_1122,N_894,N_923);
nor U1123 (N_1123,N_822,N_992);
or U1124 (N_1124,N_939,N_870);
and U1125 (N_1125,N_996,N_891);
or U1126 (N_1126,N_910,N_876);
nand U1127 (N_1127,N_977,N_847);
and U1128 (N_1128,N_957,N_890);
nand U1129 (N_1129,N_951,N_953);
nor U1130 (N_1130,N_828,N_801);
and U1131 (N_1131,N_896,N_977);
nand U1132 (N_1132,N_915,N_959);
and U1133 (N_1133,N_832,N_860);
xnor U1134 (N_1134,N_802,N_901);
or U1135 (N_1135,N_912,N_986);
nor U1136 (N_1136,N_805,N_954);
nand U1137 (N_1137,N_945,N_932);
nor U1138 (N_1138,N_992,N_825);
nor U1139 (N_1139,N_843,N_831);
xnor U1140 (N_1140,N_999,N_803);
and U1141 (N_1141,N_819,N_866);
nand U1142 (N_1142,N_968,N_814);
nor U1143 (N_1143,N_952,N_860);
nand U1144 (N_1144,N_843,N_880);
nor U1145 (N_1145,N_919,N_994);
nand U1146 (N_1146,N_955,N_876);
or U1147 (N_1147,N_909,N_921);
or U1148 (N_1148,N_854,N_974);
or U1149 (N_1149,N_869,N_821);
nor U1150 (N_1150,N_886,N_989);
or U1151 (N_1151,N_917,N_807);
and U1152 (N_1152,N_942,N_992);
and U1153 (N_1153,N_985,N_986);
nand U1154 (N_1154,N_853,N_904);
nor U1155 (N_1155,N_989,N_970);
xnor U1156 (N_1156,N_971,N_877);
xnor U1157 (N_1157,N_872,N_947);
and U1158 (N_1158,N_964,N_981);
nand U1159 (N_1159,N_864,N_893);
or U1160 (N_1160,N_862,N_965);
or U1161 (N_1161,N_877,N_954);
nor U1162 (N_1162,N_823,N_804);
xor U1163 (N_1163,N_993,N_946);
or U1164 (N_1164,N_899,N_810);
and U1165 (N_1165,N_963,N_805);
xor U1166 (N_1166,N_944,N_970);
xor U1167 (N_1167,N_914,N_801);
and U1168 (N_1168,N_999,N_840);
nand U1169 (N_1169,N_975,N_881);
xor U1170 (N_1170,N_969,N_977);
or U1171 (N_1171,N_897,N_911);
nand U1172 (N_1172,N_805,N_893);
or U1173 (N_1173,N_922,N_833);
nor U1174 (N_1174,N_808,N_855);
nand U1175 (N_1175,N_867,N_903);
nand U1176 (N_1176,N_934,N_908);
nor U1177 (N_1177,N_925,N_807);
and U1178 (N_1178,N_866,N_825);
xnor U1179 (N_1179,N_889,N_813);
nand U1180 (N_1180,N_945,N_889);
nor U1181 (N_1181,N_928,N_804);
nand U1182 (N_1182,N_862,N_895);
or U1183 (N_1183,N_829,N_928);
or U1184 (N_1184,N_827,N_927);
or U1185 (N_1185,N_818,N_922);
and U1186 (N_1186,N_926,N_928);
or U1187 (N_1187,N_885,N_847);
or U1188 (N_1188,N_833,N_851);
or U1189 (N_1189,N_814,N_919);
and U1190 (N_1190,N_813,N_839);
nor U1191 (N_1191,N_951,N_982);
and U1192 (N_1192,N_856,N_816);
xnor U1193 (N_1193,N_863,N_888);
or U1194 (N_1194,N_867,N_885);
and U1195 (N_1195,N_898,N_936);
and U1196 (N_1196,N_934,N_909);
xnor U1197 (N_1197,N_917,N_862);
xnor U1198 (N_1198,N_961,N_842);
or U1199 (N_1199,N_979,N_800);
xor U1200 (N_1200,N_1161,N_1173);
nand U1201 (N_1201,N_1093,N_1110);
nor U1202 (N_1202,N_1164,N_1169);
and U1203 (N_1203,N_1143,N_1134);
or U1204 (N_1204,N_1028,N_1045);
or U1205 (N_1205,N_1010,N_1176);
or U1206 (N_1206,N_1195,N_1021);
nand U1207 (N_1207,N_1139,N_1054);
xor U1208 (N_1208,N_1071,N_1165);
or U1209 (N_1209,N_1097,N_1152);
or U1210 (N_1210,N_1146,N_1072);
or U1211 (N_1211,N_1124,N_1175);
xor U1212 (N_1212,N_1055,N_1184);
or U1213 (N_1213,N_1131,N_1109);
nor U1214 (N_1214,N_1101,N_1114);
or U1215 (N_1215,N_1000,N_1057);
or U1216 (N_1216,N_1138,N_1056);
nor U1217 (N_1217,N_1081,N_1122);
nand U1218 (N_1218,N_1074,N_1193);
nand U1219 (N_1219,N_1182,N_1127);
and U1220 (N_1220,N_1002,N_1064);
and U1221 (N_1221,N_1188,N_1151);
xor U1222 (N_1222,N_1020,N_1062);
nor U1223 (N_1223,N_1177,N_1060);
or U1224 (N_1224,N_1157,N_1179);
nor U1225 (N_1225,N_1191,N_1168);
nor U1226 (N_1226,N_1065,N_1026);
and U1227 (N_1227,N_1186,N_1133);
nor U1228 (N_1228,N_1194,N_1059);
nor U1229 (N_1229,N_1012,N_1132);
nand U1230 (N_1230,N_1166,N_1106);
nand U1231 (N_1231,N_1199,N_1008);
nand U1232 (N_1232,N_1135,N_1047);
and U1233 (N_1233,N_1043,N_1086);
nand U1234 (N_1234,N_1128,N_1033);
nand U1235 (N_1235,N_1156,N_1118);
xnor U1236 (N_1236,N_1113,N_1196);
or U1237 (N_1237,N_1084,N_1100);
and U1238 (N_1238,N_1070,N_1050);
and U1239 (N_1239,N_1170,N_1107);
nor U1240 (N_1240,N_1015,N_1142);
and U1241 (N_1241,N_1190,N_1096);
xnor U1242 (N_1242,N_1068,N_1119);
nor U1243 (N_1243,N_1123,N_1125);
xor U1244 (N_1244,N_1046,N_1116);
nor U1245 (N_1245,N_1187,N_1129);
xor U1246 (N_1246,N_1058,N_1159);
nand U1247 (N_1247,N_1094,N_1042);
xor U1248 (N_1248,N_1183,N_1019);
nor U1249 (N_1249,N_1089,N_1063);
or U1250 (N_1250,N_1076,N_1174);
or U1251 (N_1251,N_1117,N_1039);
nand U1252 (N_1252,N_1080,N_1115);
or U1253 (N_1253,N_1163,N_1083);
nor U1254 (N_1254,N_1085,N_1037);
xor U1255 (N_1255,N_1016,N_1120);
and U1256 (N_1256,N_1171,N_1067);
or U1257 (N_1257,N_1181,N_1024);
nand U1258 (N_1258,N_1051,N_1189);
xor U1259 (N_1259,N_1052,N_1004);
nor U1260 (N_1260,N_1147,N_1022);
or U1261 (N_1261,N_1144,N_1029);
and U1262 (N_1262,N_1141,N_1077);
and U1263 (N_1263,N_1030,N_1198);
and U1264 (N_1264,N_1155,N_1178);
nand U1265 (N_1265,N_1025,N_1040);
nand U1266 (N_1266,N_1053,N_1108);
xnor U1267 (N_1267,N_1034,N_1145);
xnor U1268 (N_1268,N_1136,N_1087);
xor U1269 (N_1269,N_1009,N_1090);
or U1270 (N_1270,N_1073,N_1036);
nor U1271 (N_1271,N_1023,N_1075);
nor U1272 (N_1272,N_1111,N_1121);
or U1273 (N_1273,N_1149,N_1148);
xor U1274 (N_1274,N_1103,N_1017);
xor U1275 (N_1275,N_1003,N_1098);
or U1276 (N_1276,N_1061,N_1192);
xnor U1277 (N_1277,N_1035,N_1088);
nor U1278 (N_1278,N_1153,N_1049);
xor U1279 (N_1279,N_1041,N_1048);
or U1280 (N_1280,N_1112,N_1167);
or U1281 (N_1281,N_1069,N_1092);
nor U1282 (N_1282,N_1018,N_1006);
xor U1283 (N_1283,N_1197,N_1140);
xnor U1284 (N_1284,N_1079,N_1102);
or U1285 (N_1285,N_1160,N_1185);
xor U1286 (N_1286,N_1011,N_1078);
nand U1287 (N_1287,N_1044,N_1162);
and U1288 (N_1288,N_1014,N_1154);
and U1289 (N_1289,N_1104,N_1099);
or U1290 (N_1290,N_1091,N_1013);
and U1291 (N_1291,N_1005,N_1032);
xnor U1292 (N_1292,N_1137,N_1038);
and U1293 (N_1293,N_1126,N_1105);
nor U1294 (N_1294,N_1158,N_1180);
xnor U1295 (N_1295,N_1031,N_1172);
xor U1296 (N_1296,N_1027,N_1066);
nand U1297 (N_1297,N_1001,N_1095);
nand U1298 (N_1298,N_1007,N_1082);
xor U1299 (N_1299,N_1130,N_1150);
nand U1300 (N_1300,N_1152,N_1158);
nor U1301 (N_1301,N_1022,N_1120);
or U1302 (N_1302,N_1073,N_1147);
nor U1303 (N_1303,N_1000,N_1133);
nor U1304 (N_1304,N_1131,N_1159);
xor U1305 (N_1305,N_1153,N_1168);
nand U1306 (N_1306,N_1021,N_1177);
and U1307 (N_1307,N_1034,N_1160);
and U1308 (N_1308,N_1172,N_1156);
nand U1309 (N_1309,N_1152,N_1054);
nand U1310 (N_1310,N_1078,N_1030);
and U1311 (N_1311,N_1176,N_1161);
xor U1312 (N_1312,N_1040,N_1001);
and U1313 (N_1313,N_1079,N_1016);
and U1314 (N_1314,N_1192,N_1086);
xnor U1315 (N_1315,N_1114,N_1142);
xor U1316 (N_1316,N_1078,N_1044);
nor U1317 (N_1317,N_1000,N_1140);
and U1318 (N_1318,N_1076,N_1179);
nand U1319 (N_1319,N_1192,N_1003);
xor U1320 (N_1320,N_1070,N_1061);
and U1321 (N_1321,N_1103,N_1042);
xor U1322 (N_1322,N_1001,N_1053);
nand U1323 (N_1323,N_1072,N_1145);
nand U1324 (N_1324,N_1174,N_1015);
or U1325 (N_1325,N_1125,N_1033);
nand U1326 (N_1326,N_1092,N_1062);
nand U1327 (N_1327,N_1000,N_1135);
nand U1328 (N_1328,N_1088,N_1179);
xnor U1329 (N_1329,N_1149,N_1032);
nor U1330 (N_1330,N_1165,N_1139);
nand U1331 (N_1331,N_1075,N_1186);
or U1332 (N_1332,N_1037,N_1030);
nand U1333 (N_1333,N_1019,N_1188);
xnor U1334 (N_1334,N_1046,N_1160);
and U1335 (N_1335,N_1109,N_1067);
or U1336 (N_1336,N_1063,N_1164);
nand U1337 (N_1337,N_1052,N_1023);
or U1338 (N_1338,N_1005,N_1076);
and U1339 (N_1339,N_1175,N_1015);
xnor U1340 (N_1340,N_1094,N_1164);
and U1341 (N_1341,N_1106,N_1049);
and U1342 (N_1342,N_1061,N_1183);
nor U1343 (N_1343,N_1056,N_1163);
nand U1344 (N_1344,N_1144,N_1070);
or U1345 (N_1345,N_1110,N_1039);
and U1346 (N_1346,N_1005,N_1077);
nor U1347 (N_1347,N_1007,N_1145);
and U1348 (N_1348,N_1116,N_1122);
nor U1349 (N_1349,N_1000,N_1099);
xor U1350 (N_1350,N_1071,N_1008);
nand U1351 (N_1351,N_1078,N_1175);
or U1352 (N_1352,N_1048,N_1171);
nand U1353 (N_1353,N_1032,N_1043);
xor U1354 (N_1354,N_1077,N_1173);
or U1355 (N_1355,N_1150,N_1176);
xnor U1356 (N_1356,N_1188,N_1001);
xnor U1357 (N_1357,N_1116,N_1099);
nand U1358 (N_1358,N_1063,N_1068);
or U1359 (N_1359,N_1068,N_1185);
or U1360 (N_1360,N_1088,N_1121);
nand U1361 (N_1361,N_1120,N_1150);
nor U1362 (N_1362,N_1139,N_1123);
and U1363 (N_1363,N_1159,N_1187);
xnor U1364 (N_1364,N_1004,N_1151);
xor U1365 (N_1365,N_1155,N_1104);
nor U1366 (N_1366,N_1131,N_1154);
or U1367 (N_1367,N_1103,N_1138);
xnor U1368 (N_1368,N_1111,N_1053);
nand U1369 (N_1369,N_1192,N_1006);
and U1370 (N_1370,N_1117,N_1065);
nor U1371 (N_1371,N_1146,N_1076);
and U1372 (N_1372,N_1045,N_1057);
xnor U1373 (N_1373,N_1113,N_1012);
nand U1374 (N_1374,N_1106,N_1036);
nand U1375 (N_1375,N_1149,N_1169);
and U1376 (N_1376,N_1004,N_1074);
and U1377 (N_1377,N_1077,N_1133);
or U1378 (N_1378,N_1096,N_1199);
and U1379 (N_1379,N_1114,N_1128);
nand U1380 (N_1380,N_1126,N_1062);
xor U1381 (N_1381,N_1060,N_1151);
xnor U1382 (N_1382,N_1018,N_1110);
or U1383 (N_1383,N_1180,N_1163);
nor U1384 (N_1384,N_1056,N_1015);
xnor U1385 (N_1385,N_1043,N_1187);
and U1386 (N_1386,N_1084,N_1156);
or U1387 (N_1387,N_1092,N_1010);
nor U1388 (N_1388,N_1171,N_1013);
and U1389 (N_1389,N_1115,N_1048);
nand U1390 (N_1390,N_1055,N_1109);
xnor U1391 (N_1391,N_1176,N_1121);
nor U1392 (N_1392,N_1002,N_1115);
or U1393 (N_1393,N_1155,N_1185);
nand U1394 (N_1394,N_1044,N_1163);
xnor U1395 (N_1395,N_1153,N_1073);
nor U1396 (N_1396,N_1103,N_1149);
and U1397 (N_1397,N_1121,N_1022);
xor U1398 (N_1398,N_1152,N_1165);
xnor U1399 (N_1399,N_1187,N_1009);
xnor U1400 (N_1400,N_1323,N_1210);
xor U1401 (N_1401,N_1265,N_1297);
or U1402 (N_1402,N_1306,N_1280);
nor U1403 (N_1403,N_1230,N_1277);
or U1404 (N_1404,N_1202,N_1328);
and U1405 (N_1405,N_1367,N_1307);
and U1406 (N_1406,N_1236,N_1361);
nand U1407 (N_1407,N_1331,N_1244);
xor U1408 (N_1408,N_1300,N_1369);
xor U1409 (N_1409,N_1313,N_1376);
nand U1410 (N_1410,N_1336,N_1251);
nor U1411 (N_1411,N_1312,N_1345);
nand U1412 (N_1412,N_1375,N_1200);
nor U1413 (N_1413,N_1247,N_1326);
xor U1414 (N_1414,N_1386,N_1397);
and U1415 (N_1415,N_1310,N_1393);
nor U1416 (N_1416,N_1366,N_1344);
nand U1417 (N_1417,N_1253,N_1235);
xor U1418 (N_1418,N_1260,N_1221);
nor U1419 (N_1419,N_1392,N_1281);
xnor U1420 (N_1420,N_1296,N_1285);
nor U1421 (N_1421,N_1261,N_1232);
xnor U1422 (N_1422,N_1324,N_1275);
nand U1423 (N_1423,N_1282,N_1292);
or U1424 (N_1424,N_1231,N_1321);
and U1425 (N_1425,N_1320,N_1342);
or U1426 (N_1426,N_1363,N_1316);
xnor U1427 (N_1427,N_1303,N_1272);
and U1428 (N_1428,N_1274,N_1377);
xor U1429 (N_1429,N_1388,N_1325);
nand U1430 (N_1430,N_1359,N_1206);
and U1431 (N_1431,N_1238,N_1372);
xor U1432 (N_1432,N_1276,N_1295);
nor U1433 (N_1433,N_1314,N_1399);
nor U1434 (N_1434,N_1243,N_1264);
nor U1435 (N_1435,N_1252,N_1207);
xor U1436 (N_1436,N_1353,N_1224);
nor U1437 (N_1437,N_1246,N_1315);
or U1438 (N_1438,N_1364,N_1337);
and U1439 (N_1439,N_1268,N_1319);
xnor U1440 (N_1440,N_1370,N_1245);
and U1441 (N_1441,N_1254,N_1341);
or U1442 (N_1442,N_1209,N_1287);
xnor U1443 (N_1443,N_1360,N_1343);
or U1444 (N_1444,N_1284,N_1346);
and U1445 (N_1445,N_1380,N_1215);
nand U1446 (N_1446,N_1212,N_1213);
nor U1447 (N_1447,N_1394,N_1239);
xor U1448 (N_1448,N_1271,N_1349);
and U1449 (N_1449,N_1299,N_1368);
and U1450 (N_1450,N_1354,N_1290);
and U1451 (N_1451,N_1233,N_1226);
xnor U1452 (N_1452,N_1242,N_1347);
or U1453 (N_1453,N_1257,N_1217);
and U1454 (N_1454,N_1240,N_1220);
or U1455 (N_1455,N_1269,N_1355);
or U1456 (N_1456,N_1241,N_1203);
or U1457 (N_1457,N_1216,N_1278);
and U1458 (N_1458,N_1309,N_1229);
nor U1459 (N_1459,N_1334,N_1234);
or U1460 (N_1460,N_1317,N_1373);
and U1461 (N_1461,N_1270,N_1329);
xnor U1462 (N_1462,N_1298,N_1279);
nand U1463 (N_1463,N_1291,N_1225);
xor U1464 (N_1464,N_1294,N_1338);
or U1465 (N_1465,N_1382,N_1389);
or U1466 (N_1466,N_1396,N_1339);
and U1467 (N_1467,N_1381,N_1356);
nand U1468 (N_1468,N_1350,N_1387);
and U1469 (N_1469,N_1286,N_1384);
and U1470 (N_1470,N_1333,N_1378);
or U1471 (N_1471,N_1273,N_1222);
nor U1472 (N_1472,N_1374,N_1223);
nand U1473 (N_1473,N_1214,N_1258);
or U1474 (N_1474,N_1228,N_1357);
and U1475 (N_1475,N_1391,N_1289);
nor U1476 (N_1476,N_1249,N_1390);
nand U1477 (N_1477,N_1358,N_1255);
xor U1478 (N_1478,N_1340,N_1259);
or U1479 (N_1479,N_1301,N_1395);
nand U1480 (N_1480,N_1352,N_1379);
xnor U1481 (N_1481,N_1311,N_1348);
nand U1482 (N_1482,N_1205,N_1219);
nand U1483 (N_1483,N_1266,N_1383);
and U1484 (N_1484,N_1211,N_1305);
and U1485 (N_1485,N_1304,N_1371);
and U1486 (N_1486,N_1385,N_1365);
or U1487 (N_1487,N_1283,N_1256);
nand U1488 (N_1488,N_1293,N_1288);
nor U1489 (N_1489,N_1267,N_1237);
xnor U1490 (N_1490,N_1204,N_1330);
and U1491 (N_1491,N_1218,N_1250);
nor U1492 (N_1492,N_1308,N_1362);
nor U1493 (N_1493,N_1351,N_1322);
xnor U1494 (N_1494,N_1335,N_1302);
and U1495 (N_1495,N_1263,N_1248);
nand U1496 (N_1496,N_1208,N_1201);
xor U1497 (N_1497,N_1227,N_1398);
xnor U1498 (N_1498,N_1262,N_1318);
nor U1499 (N_1499,N_1327,N_1332);
nand U1500 (N_1500,N_1200,N_1221);
or U1501 (N_1501,N_1352,N_1279);
xor U1502 (N_1502,N_1258,N_1338);
xnor U1503 (N_1503,N_1224,N_1297);
xor U1504 (N_1504,N_1203,N_1238);
and U1505 (N_1505,N_1396,N_1202);
or U1506 (N_1506,N_1378,N_1260);
nor U1507 (N_1507,N_1265,N_1324);
xnor U1508 (N_1508,N_1399,N_1337);
xor U1509 (N_1509,N_1388,N_1211);
or U1510 (N_1510,N_1321,N_1235);
and U1511 (N_1511,N_1206,N_1239);
nand U1512 (N_1512,N_1380,N_1214);
xor U1513 (N_1513,N_1326,N_1248);
and U1514 (N_1514,N_1362,N_1304);
nor U1515 (N_1515,N_1245,N_1243);
nor U1516 (N_1516,N_1372,N_1377);
or U1517 (N_1517,N_1367,N_1351);
nor U1518 (N_1518,N_1398,N_1207);
nand U1519 (N_1519,N_1394,N_1271);
or U1520 (N_1520,N_1397,N_1329);
and U1521 (N_1521,N_1216,N_1309);
or U1522 (N_1522,N_1317,N_1261);
nor U1523 (N_1523,N_1335,N_1218);
xor U1524 (N_1524,N_1371,N_1219);
and U1525 (N_1525,N_1224,N_1279);
or U1526 (N_1526,N_1279,N_1332);
nor U1527 (N_1527,N_1387,N_1264);
nor U1528 (N_1528,N_1292,N_1204);
nor U1529 (N_1529,N_1353,N_1371);
xnor U1530 (N_1530,N_1382,N_1260);
xor U1531 (N_1531,N_1309,N_1379);
and U1532 (N_1532,N_1334,N_1261);
or U1533 (N_1533,N_1239,N_1256);
and U1534 (N_1534,N_1263,N_1316);
nand U1535 (N_1535,N_1243,N_1399);
and U1536 (N_1536,N_1332,N_1322);
and U1537 (N_1537,N_1243,N_1375);
nor U1538 (N_1538,N_1354,N_1243);
and U1539 (N_1539,N_1235,N_1272);
xnor U1540 (N_1540,N_1355,N_1244);
nand U1541 (N_1541,N_1383,N_1215);
nand U1542 (N_1542,N_1269,N_1399);
nand U1543 (N_1543,N_1378,N_1266);
and U1544 (N_1544,N_1212,N_1243);
nand U1545 (N_1545,N_1316,N_1222);
nand U1546 (N_1546,N_1225,N_1304);
and U1547 (N_1547,N_1375,N_1392);
xor U1548 (N_1548,N_1266,N_1208);
nand U1549 (N_1549,N_1240,N_1221);
xor U1550 (N_1550,N_1395,N_1278);
or U1551 (N_1551,N_1385,N_1222);
nor U1552 (N_1552,N_1307,N_1240);
nor U1553 (N_1553,N_1245,N_1213);
and U1554 (N_1554,N_1324,N_1348);
nor U1555 (N_1555,N_1259,N_1230);
or U1556 (N_1556,N_1201,N_1350);
xor U1557 (N_1557,N_1383,N_1298);
nand U1558 (N_1558,N_1342,N_1263);
xor U1559 (N_1559,N_1253,N_1393);
or U1560 (N_1560,N_1309,N_1382);
and U1561 (N_1561,N_1296,N_1306);
or U1562 (N_1562,N_1294,N_1391);
nand U1563 (N_1563,N_1378,N_1304);
nor U1564 (N_1564,N_1213,N_1271);
xnor U1565 (N_1565,N_1219,N_1330);
nor U1566 (N_1566,N_1327,N_1241);
and U1567 (N_1567,N_1207,N_1282);
xor U1568 (N_1568,N_1238,N_1366);
nor U1569 (N_1569,N_1212,N_1394);
nand U1570 (N_1570,N_1376,N_1250);
nor U1571 (N_1571,N_1373,N_1379);
and U1572 (N_1572,N_1311,N_1217);
and U1573 (N_1573,N_1347,N_1225);
and U1574 (N_1574,N_1327,N_1220);
nor U1575 (N_1575,N_1205,N_1242);
nor U1576 (N_1576,N_1353,N_1251);
nand U1577 (N_1577,N_1316,N_1375);
nand U1578 (N_1578,N_1251,N_1367);
and U1579 (N_1579,N_1302,N_1276);
and U1580 (N_1580,N_1390,N_1283);
xnor U1581 (N_1581,N_1367,N_1208);
xor U1582 (N_1582,N_1239,N_1371);
nand U1583 (N_1583,N_1208,N_1388);
xnor U1584 (N_1584,N_1271,N_1372);
nand U1585 (N_1585,N_1201,N_1386);
nand U1586 (N_1586,N_1266,N_1236);
nand U1587 (N_1587,N_1243,N_1270);
or U1588 (N_1588,N_1364,N_1349);
nand U1589 (N_1589,N_1373,N_1339);
nor U1590 (N_1590,N_1297,N_1217);
nand U1591 (N_1591,N_1347,N_1332);
and U1592 (N_1592,N_1299,N_1311);
or U1593 (N_1593,N_1373,N_1283);
or U1594 (N_1594,N_1354,N_1361);
or U1595 (N_1595,N_1257,N_1348);
or U1596 (N_1596,N_1250,N_1382);
and U1597 (N_1597,N_1342,N_1201);
xor U1598 (N_1598,N_1350,N_1279);
nor U1599 (N_1599,N_1222,N_1302);
nand U1600 (N_1600,N_1423,N_1558);
xnor U1601 (N_1601,N_1527,N_1468);
and U1602 (N_1602,N_1418,N_1460);
or U1603 (N_1603,N_1471,N_1454);
nand U1604 (N_1604,N_1456,N_1432);
or U1605 (N_1605,N_1495,N_1469);
and U1606 (N_1606,N_1565,N_1400);
or U1607 (N_1607,N_1451,N_1444);
nor U1608 (N_1608,N_1455,N_1516);
xnor U1609 (N_1609,N_1493,N_1443);
nand U1610 (N_1610,N_1467,N_1539);
or U1611 (N_1611,N_1434,N_1429);
xnor U1612 (N_1612,N_1478,N_1419);
nand U1613 (N_1613,N_1492,N_1591);
or U1614 (N_1614,N_1531,N_1563);
and U1615 (N_1615,N_1413,N_1596);
nor U1616 (N_1616,N_1550,N_1557);
xor U1617 (N_1617,N_1409,N_1485);
nand U1618 (N_1618,N_1502,N_1564);
nand U1619 (N_1619,N_1504,N_1554);
nand U1620 (N_1620,N_1496,N_1580);
and U1621 (N_1621,N_1599,N_1431);
xor U1622 (N_1622,N_1545,N_1405);
xnor U1623 (N_1623,N_1517,N_1543);
and U1624 (N_1624,N_1421,N_1500);
xor U1625 (N_1625,N_1537,N_1403);
or U1626 (N_1626,N_1466,N_1404);
or U1627 (N_1627,N_1586,N_1506);
and U1628 (N_1628,N_1523,N_1453);
and U1629 (N_1629,N_1452,N_1530);
or U1630 (N_1630,N_1512,N_1576);
or U1631 (N_1631,N_1570,N_1511);
or U1632 (N_1632,N_1417,N_1437);
and U1633 (N_1633,N_1542,N_1435);
and U1634 (N_1634,N_1473,N_1498);
or U1635 (N_1635,N_1551,N_1470);
nor U1636 (N_1636,N_1572,N_1441);
or U1637 (N_1637,N_1491,N_1535);
nand U1638 (N_1638,N_1401,N_1503);
xor U1639 (N_1639,N_1406,N_1497);
nand U1640 (N_1640,N_1465,N_1509);
nand U1641 (N_1641,N_1578,N_1448);
and U1642 (N_1642,N_1488,N_1449);
or U1643 (N_1643,N_1522,N_1479);
nand U1644 (N_1644,N_1507,N_1583);
nor U1645 (N_1645,N_1582,N_1556);
nor U1646 (N_1646,N_1597,N_1529);
nor U1647 (N_1647,N_1445,N_1414);
or U1648 (N_1648,N_1490,N_1568);
xor U1649 (N_1649,N_1501,N_1459);
nor U1650 (N_1650,N_1415,N_1426);
nor U1651 (N_1651,N_1487,N_1528);
nand U1652 (N_1652,N_1581,N_1584);
and U1653 (N_1653,N_1446,N_1571);
or U1654 (N_1654,N_1588,N_1475);
and U1655 (N_1655,N_1519,N_1520);
and U1656 (N_1656,N_1515,N_1579);
nor U1657 (N_1657,N_1433,N_1561);
and U1658 (N_1658,N_1447,N_1411);
nand U1659 (N_1659,N_1463,N_1440);
xor U1660 (N_1660,N_1424,N_1518);
nand U1661 (N_1661,N_1547,N_1590);
xnor U1662 (N_1662,N_1457,N_1482);
and U1663 (N_1663,N_1593,N_1461);
nand U1664 (N_1664,N_1562,N_1589);
and U1665 (N_1665,N_1489,N_1499);
and U1666 (N_1666,N_1428,N_1476);
and U1667 (N_1667,N_1477,N_1508);
or U1668 (N_1668,N_1514,N_1534);
nor U1669 (N_1669,N_1464,N_1458);
nand U1670 (N_1670,N_1513,N_1587);
or U1671 (N_1671,N_1430,N_1480);
xnor U1672 (N_1672,N_1462,N_1532);
xor U1673 (N_1673,N_1544,N_1574);
and U1674 (N_1674,N_1472,N_1510);
nor U1675 (N_1675,N_1573,N_1598);
nand U1676 (N_1676,N_1402,N_1553);
nor U1677 (N_1677,N_1484,N_1575);
xor U1678 (N_1678,N_1422,N_1536);
nor U1679 (N_1679,N_1486,N_1416);
nand U1680 (N_1680,N_1420,N_1566);
or U1681 (N_1681,N_1538,N_1552);
nor U1682 (N_1682,N_1567,N_1541);
nand U1683 (N_1683,N_1577,N_1540);
and U1684 (N_1684,N_1410,N_1585);
nor U1685 (N_1685,N_1436,N_1427);
and U1686 (N_1686,N_1483,N_1425);
nand U1687 (N_1687,N_1442,N_1524);
and U1688 (N_1688,N_1569,N_1412);
xnor U1689 (N_1689,N_1546,N_1521);
nor U1690 (N_1690,N_1548,N_1474);
or U1691 (N_1691,N_1439,N_1525);
or U1692 (N_1692,N_1481,N_1560);
xor U1693 (N_1693,N_1594,N_1494);
or U1694 (N_1694,N_1505,N_1592);
nor U1695 (N_1695,N_1526,N_1407);
xnor U1696 (N_1696,N_1438,N_1549);
or U1697 (N_1697,N_1533,N_1450);
xor U1698 (N_1698,N_1555,N_1559);
or U1699 (N_1699,N_1595,N_1408);
and U1700 (N_1700,N_1518,N_1466);
nand U1701 (N_1701,N_1566,N_1431);
or U1702 (N_1702,N_1597,N_1527);
xor U1703 (N_1703,N_1545,N_1540);
nand U1704 (N_1704,N_1458,N_1444);
nor U1705 (N_1705,N_1473,N_1548);
or U1706 (N_1706,N_1479,N_1553);
xor U1707 (N_1707,N_1547,N_1476);
nor U1708 (N_1708,N_1457,N_1554);
or U1709 (N_1709,N_1570,N_1523);
and U1710 (N_1710,N_1562,N_1499);
xnor U1711 (N_1711,N_1505,N_1411);
or U1712 (N_1712,N_1406,N_1403);
xor U1713 (N_1713,N_1561,N_1464);
nor U1714 (N_1714,N_1531,N_1400);
xor U1715 (N_1715,N_1580,N_1561);
nor U1716 (N_1716,N_1474,N_1585);
nor U1717 (N_1717,N_1553,N_1571);
or U1718 (N_1718,N_1402,N_1567);
nand U1719 (N_1719,N_1468,N_1441);
xor U1720 (N_1720,N_1406,N_1433);
and U1721 (N_1721,N_1586,N_1417);
nor U1722 (N_1722,N_1473,N_1488);
or U1723 (N_1723,N_1557,N_1459);
and U1724 (N_1724,N_1406,N_1501);
nor U1725 (N_1725,N_1441,N_1475);
xor U1726 (N_1726,N_1432,N_1429);
nor U1727 (N_1727,N_1532,N_1476);
nand U1728 (N_1728,N_1423,N_1512);
and U1729 (N_1729,N_1473,N_1587);
nand U1730 (N_1730,N_1508,N_1461);
xor U1731 (N_1731,N_1562,N_1559);
xor U1732 (N_1732,N_1539,N_1483);
and U1733 (N_1733,N_1475,N_1538);
and U1734 (N_1734,N_1545,N_1444);
xor U1735 (N_1735,N_1415,N_1473);
or U1736 (N_1736,N_1409,N_1405);
and U1737 (N_1737,N_1512,N_1503);
nor U1738 (N_1738,N_1547,N_1475);
and U1739 (N_1739,N_1526,N_1531);
or U1740 (N_1740,N_1525,N_1425);
nand U1741 (N_1741,N_1529,N_1451);
or U1742 (N_1742,N_1499,N_1449);
nor U1743 (N_1743,N_1488,N_1565);
or U1744 (N_1744,N_1594,N_1493);
and U1745 (N_1745,N_1575,N_1586);
xor U1746 (N_1746,N_1449,N_1458);
xor U1747 (N_1747,N_1529,N_1420);
nand U1748 (N_1748,N_1565,N_1427);
nand U1749 (N_1749,N_1418,N_1511);
nor U1750 (N_1750,N_1554,N_1434);
xor U1751 (N_1751,N_1514,N_1556);
xnor U1752 (N_1752,N_1539,N_1597);
xnor U1753 (N_1753,N_1472,N_1430);
nand U1754 (N_1754,N_1599,N_1480);
xnor U1755 (N_1755,N_1526,N_1516);
nor U1756 (N_1756,N_1463,N_1423);
nor U1757 (N_1757,N_1455,N_1567);
nand U1758 (N_1758,N_1521,N_1554);
nor U1759 (N_1759,N_1415,N_1577);
or U1760 (N_1760,N_1583,N_1400);
xnor U1761 (N_1761,N_1419,N_1539);
xnor U1762 (N_1762,N_1459,N_1507);
nand U1763 (N_1763,N_1405,N_1410);
xnor U1764 (N_1764,N_1478,N_1523);
or U1765 (N_1765,N_1560,N_1461);
nor U1766 (N_1766,N_1592,N_1567);
nand U1767 (N_1767,N_1447,N_1500);
nor U1768 (N_1768,N_1477,N_1570);
nor U1769 (N_1769,N_1469,N_1530);
nor U1770 (N_1770,N_1590,N_1521);
and U1771 (N_1771,N_1428,N_1590);
nor U1772 (N_1772,N_1549,N_1545);
or U1773 (N_1773,N_1460,N_1424);
nand U1774 (N_1774,N_1577,N_1517);
nand U1775 (N_1775,N_1497,N_1544);
xor U1776 (N_1776,N_1447,N_1477);
and U1777 (N_1777,N_1424,N_1489);
xnor U1778 (N_1778,N_1455,N_1595);
and U1779 (N_1779,N_1460,N_1432);
and U1780 (N_1780,N_1448,N_1517);
and U1781 (N_1781,N_1566,N_1450);
nand U1782 (N_1782,N_1491,N_1404);
nand U1783 (N_1783,N_1580,N_1576);
or U1784 (N_1784,N_1510,N_1537);
and U1785 (N_1785,N_1409,N_1511);
nor U1786 (N_1786,N_1443,N_1465);
xnor U1787 (N_1787,N_1588,N_1476);
xnor U1788 (N_1788,N_1424,N_1498);
xnor U1789 (N_1789,N_1569,N_1490);
or U1790 (N_1790,N_1531,N_1463);
or U1791 (N_1791,N_1437,N_1553);
nand U1792 (N_1792,N_1596,N_1499);
and U1793 (N_1793,N_1541,N_1523);
nor U1794 (N_1794,N_1465,N_1468);
nor U1795 (N_1795,N_1569,N_1561);
xnor U1796 (N_1796,N_1489,N_1403);
or U1797 (N_1797,N_1491,N_1556);
or U1798 (N_1798,N_1427,N_1407);
nand U1799 (N_1799,N_1470,N_1460);
or U1800 (N_1800,N_1648,N_1656);
or U1801 (N_1801,N_1735,N_1659);
nand U1802 (N_1802,N_1715,N_1708);
nor U1803 (N_1803,N_1742,N_1621);
and U1804 (N_1804,N_1691,N_1617);
nand U1805 (N_1805,N_1745,N_1679);
and U1806 (N_1806,N_1615,N_1701);
nand U1807 (N_1807,N_1794,N_1752);
or U1808 (N_1808,N_1685,N_1601);
xnor U1809 (N_1809,N_1793,N_1729);
nand U1810 (N_1810,N_1636,N_1781);
and U1811 (N_1811,N_1790,N_1632);
nand U1812 (N_1812,N_1756,N_1605);
nand U1813 (N_1813,N_1643,N_1670);
or U1814 (N_1814,N_1719,N_1754);
nand U1815 (N_1815,N_1792,N_1624);
nor U1816 (N_1816,N_1777,N_1630);
nand U1817 (N_1817,N_1619,N_1799);
xor U1818 (N_1818,N_1710,N_1649);
and U1819 (N_1819,N_1626,N_1640);
and U1820 (N_1820,N_1780,N_1749);
xnor U1821 (N_1821,N_1655,N_1700);
xor U1822 (N_1822,N_1722,N_1771);
xor U1823 (N_1823,N_1690,N_1646);
xor U1824 (N_1824,N_1681,N_1712);
xor U1825 (N_1825,N_1741,N_1772);
and U1826 (N_1826,N_1608,N_1653);
nand U1827 (N_1827,N_1694,N_1686);
and U1828 (N_1828,N_1634,N_1695);
xor U1829 (N_1829,N_1744,N_1689);
nand U1830 (N_1830,N_1737,N_1674);
or U1831 (N_1831,N_1618,N_1609);
nor U1832 (N_1832,N_1673,N_1676);
nor U1833 (N_1833,N_1782,N_1714);
nor U1834 (N_1834,N_1740,N_1769);
nand U1835 (N_1835,N_1651,N_1760);
or U1836 (N_1836,N_1731,N_1684);
or U1837 (N_1837,N_1774,N_1638);
or U1838 (N_1838,N_1660,N_1797);
nor U1839 (N_1839,N_1658,N_1633);
and U1840 (N_1840,N_1704,N_1620);
xnor U1841 (N_1841,N_1709,N_1600);
nand U1842 (N_1842,N_1604,N_1637);
and U1843 (N_1843,N_1642,N_1688);
nor U1844 (N_1844,N_1785,N_1678);
nor U1845 (N_1845,N_1762,N_1711);
nand U1846 (N_1846,N_1661,N_1697);
nand U1847 (N_1847,N_1664,N_1786);
nand U1848 (N_1848,N_1706,N_1759);
nand U1849 (N_1849,N_1767,N_1627);
nor U1850 (N_1850,N_1666,N_1779);
nor U1851 (N_1851,N_1692,N_1625);
and U1852 (N_1852,N_1764,N_1611);
xor U1853 (N_1853,N_1758,N_1721);
nand U1854 (N_1854,N_1727,N_1789);
nor U1855 (N_1855,N_1736,N_1716);
or U1856 (N_1856,N_1641,N_1650);
nand U1857 (N_1857,N_1602,N_1662);
xor U1858 (N_1858,N_1761,N_1613);
xnor U1859 (N_1859,N_1622,N_1603);
and U1860 (N_1860,N_1672,N_1763);
or U1861 (N_1861,N_1788,N_1607);
nand U1862 (N_1862,N_1610,N_1726);
and U1863 (N_1863,N_1628,N_1734);
and U1864 (N_1864,N_1765,N_1753);
xnor U1865 (N_1865,N_1644,N_1614);
nor U1866 (N_1866,N_1796,N_1787);
nor U1867 (N_1867,N_1705,N_1730);
nand U1868 (N_1868,N_1669,N_1748);
xor U1869 (N_1869,N_1612,N_1687);
nor U1870 (N_1870,N_1616,N_1738);
nand U1871 (N_1871,N_1629,N_1783);
nand U1872 (N_1872,N_1720,N_1723);
or U1873 (N_1873,N_1703,N_1635);
and U1874 (N_1874,N_1791,N_1718);
or U1875 (N_1875,N_1770,N_1747);
xor U1876 (N_1876,N_1683,N_1675);
xor U1877 (N_1877,N_1652,N_1657);
xnor U1878 (N_1878,N_1784,N_1778);
or U1879 (N_1879,N_1647,N_1775);
nor U1880 (N_1880,N_1671,N_1768);
xor U1881 (N_1881,N_1663,N_1698);
or U1882 (N_1882,N_1746,N_1631);
xor U1883 (N_1883,N_1739,N_1733);
nor U1884 (N_1884,N_1798,N_1713);
or U1885 (N_1885,N_1665,N_1766);
and U1886 (N_1886,N_1728,N_1693);
or U1887 (N_1887,N_1639,N_1795);
and U1888 (N_1888,N_1743,N_1702);
nor U1889 (N_1889,N_1750,N_1773);
or U1890 (N_1890,N_1667,N_1677);
nand U1891 (N_1891,N_1696,N_1725);
and U1892 (N_1892,N_1654,N_1732);
nand U1893 (N_1893,N_1668,N_1645);
nand U1894 (N_1894,N_1751,N_1757);
nand U1895 (N_1895,N_1680,N_1776);
or U1896 (N_1896,N_1717,N_1682);
nor U1897 (N_1897,N_1606,N_1724);
xor U1898 (N_1898,N_1755,N_1623);
nand U1899 (N_1899,N_1707,N_1699);
and U1900 (N_1900,N_1744,N_1784);
nor U1901 (N_1901,N_1711,N_1688);
xor U1902 (N_1902,N_1745,N_1640);
xnor U1903 (N_1903,N_1701,N_1608);
nor U1904 (N_1904,N_1710,N_1672);
nand U1905 (N_1905,N_1645,N_1684);
nand U1906 (N_1906,N_1607,N_1695);
and U1907 (N_1907,N_1623,N_1796);
xnor U1908 (N_1908,N_1736,N_1766);
or U1909 (N_1909,N_1797,N_1629);
xor U1910 (N_1910,N_1631,N_1790);
and U1911 (N_1911,N_1725,N_1663);
nand U1912 (N_1912,N_1652,N_1766);
and U1913 (N_1913,N_1669,N_1623);
xnor U1914 (N_1914,N_1738,N_1663);
xor U1915 (N_1915,N_1732,N_1648);
and U1916 (N_1916,N_1790,N_1718);
xnor U1917 (N_1917,N_1696,N_1729);
nor U1918 (N_1918,N_1762,N_1639);
nand U1919 (N_1919,N_1681,N_1769);
nand U1920 (N_1920,N_1788,N_1616);
xnor U1921 (N_1921,N_1692,N_1752);
or U1922 (N_1922,N_1619,N_1744);
nor U1923 (N_1923,N_1719,N_1610);
nor U1924 (N_1924,N_1770,N_1677);
nand U1925 (N_1925,N_1649,N_1705);
xor U1926 (N_1926,N_1733,N_1763);
nand U1927 (N_1927,N_1660,N_1708);
or U1928 (N_1928,N_1600,N_1693);
xor U1929 (N_1929,N_1736,N_1675);
and U1930 (N_1930,N_1744,N_1723);
or U1931 (N_1931,N_1643,N_1615);
nand U1932 (N_1932,N_1659,N_1761);
nand U1933 (N_1933,N_1751,N_1706);
xnor U1934 (N_1934,N_1639,N_1797);
nor U1935 (N_1935,N_1661,N_1731);
nand U1936 (N_1936,N_1719,N_1691);
and U1937 (N_1937,N_1715,N_1625);
nor U1938 (N_1938,N_1672,N_1623);
or U1939 (N_1939,N_1678,N_1783);
and U1940 (N_1940,N_1745,N_1781);
xor U1941 (N_1941,N_1764,N_1792);
xor U1942 (N_1942,N_1687,N_1674);
or U1943 (N_1943,N_1793,N_1664);
nand U1944 (N_1944,N_1626,N_1729);
nor U1945 (N_1945,N_1623,N_1795);
or U1946 (N_1946,N_1691,N_1726);
nand U1947 (N_1947,N_1790,N_1698);
xnor U1948 (N_1948,N_1765,N_1634);
nand U1949 (N_1949,N_1764,N_1706);
nand U1950 (N_1950,N_1778,N_1709);
nor U1951 (N_1951,N_1658,N_1730);
xnor U1952 (N_1952,N_1752,N_1761);
or U1953 (N_1953,N_1664,N_1609);
nand U1954 (N_1954,N_1667,N_1724);
and U1955 (N_1955,N_1685,N_1633);
xor U1956 (N_1956,N_1660,N_1793);
or U1957 (N_1957,N_1753,N_1770);
nand U1958 (N_1958,N_1757,N_1647);
xor U1959 (N_1959,N_1746,N_1643);
nand U1960 (N_1960,N_1754,N_1675);
or U1961 (N_1961,N_1769,N_1788);
nand U1962 (N_1962,N_1645,N_1695);
xnor U1963 (N_1963,N_1623,N_1621);
nor U1964 (N_1964,N_1625,N_1777);
nor U1965 (N_1965,N_1698,N_1608);
or U1966 (N_1966,N_1633,N_1686);
nand U1967 (N_1967,N_1607,N_1755);
xnor U1968 (N_1968,N_1682,N_1635);
nor U1969 (N_1969,N_1701,N_1607);
nor U1970 (N_1970,N_1678,N_1662);
nand U1971 (N_1971,N_1622,N_1625);
and U1972 (N_1972,N_1780,N_1628);
and U1973 (N_1973,N_1633,N_1694);
xor U1974 (N_1974,N_1677,N_1710);
nand U1975 (N_1975,N_1639,N_1798);
or U1976 (N_1976,N_1716,N_1776);
xnor U1977 (N_1977,N_1638,N_1753);
xor U1978 (N_1978,N_1656,N_1618);
and U1979 (N_1979,N_1708,N_1781);
nand U1980 (N_1980,N_1617,N_1660);
xor U1981 (N_1981,N_1729,N_1615);
nor U1982 (N_1982,N_1639,N_1679);
nand U1983 (N_1983,N_1705,N_1625);
and U1984 (N_1984,N_1712,N_1723);
xor U1985 (N_1985,N_1733,N_1645);
nand U1986 (N_1986,N_1704,N_1747);
or U1987 (N_1987,N_1666,N_1729);
nand U1988 (N_1988,N_1727,N_1685);
and U1989 (N_1989,N_1642,N_1696);
nor U1990 (N_1990,N_1603,N_1629);
and U1991 (N_1991,N_1686,N_1755);
and U1992 (N_1992,N_1687,N_1754);
xnor U1993 (N_1993,N_1744,N_1720);
or U1994 (N_1994,N_1726,N_1678);
xnor U1995 (N_1995,N_1681,N_1640);
nand U1996 (N_1996,N_1722,N_1648);
nor U1997 (N_1997,N_1751,N_1698);
or U1998 (N_1998,N_1736,N_1720);
nand U1999 (N_1999,N_1784,N_1651);
xnor U2000 (N_2000,N_1912,N_1973);
nand U2001 (N_2001,N_1806,N_1940);
or U2002 (N_2002,N_1913,N_1856);
nor U2003 (N_2003,N_1843,N_1994);
and U2004 (N_2004,N_1801,N_1953);
or U2005 (N_2005,N_1834,N_1984);
or U2006 (N_2006,N_1860,N_1833);
nor U2007 (N_2007,N_1919,N_1935);
and U2008 (N_2008,N_1904,N_1849);
xnor U2009 (N_2009,N_1944,N_1946);
nor U2010 (N_2010,N_1976,N_1829);
or U2011 (N_2011,N_1985,N_1866);
and U2012 (N_2012,N_1952,N_1903);
or U2013 (N_2013,N_1881,N_1871);
nand U2014 (N_2014,N_1998,N_1805);
xnor U2015 (N_2015,N_1966,N_1960);
nor U2016 (N_2016,N_1852,N_1876);
or U2017 (N_2017,N_1879,N_1921);
nand U2018 (N_2018,N_1995,N_1978);
or U2019 (N_2019,N_1991,N_1915);
nand U2020 (N_2020,N_1885,N_1990);
xor U2021 (N_2021,N_1957,N_1857);
xor U2022 (N_2022,N_1877,N_1883);
xnor U2023 (N_2023,N_1875,N_1955);
and U2024 (N_2024,N_1932,N_1943);
and U2025 (N_2025,N_1910,N_1949);
or U2026 (N_2026,N_1977,N_1812);
or U2027 (N_2027,N_1850,N_1959);
xor U2028 (N_2028,N_1926,N_1958);
xor U2029 (N_2029,N_1815,N_1880);
nor U2030 (N_2030,N_1804,N_1870);
and U2031 (N_2031,N_1865,N_1917);
and U2032 (N_2032,N_1841,N_1964);
and U2033 (N_2033,N_1937,N_1899);
or U2034 (N_2034,N_1811,N_1873);
and U2035 (N_2035,N_1909,N_1988);
xnor U2036 (N_2036,N_1824,N_1851);
and U2037 (N_2037,N_1947,N_1882);
or U2038 (N_2038,N_1918,N_1891);
and U2039 (N_2039,N_1982,N_1950);
nor U2040 (N_2040,N_1836,N_1983);
or U2041 (N_2041,N_1837,N_1816);
nand U2042 (N_2042,N_1832,N_1965);
or U2043 (N_2043,N_1864,N_1987);
xor U2044 (N_2044,N_1825,N_1925);
xor U2045 (N_2045,N_1842,N_1808);
nor U2046 (N_2046,N_1892,N_1826);
and U2047 (N_2047,N_1906,N_1800);
nor U2048 (N_2048,N_1817,N_1928);
or U2049 (N_2049,N_1869,N_1890);
xor U2050 (N_2050,N_1969,N_1989);
or U2051 (N_2051,N_1907,N_1945);
or U2052 (N_2052,N_1996,N_1810);
nor U2053 (N_2053,N_1974,N_1874);
or U2054 (N_2054,N_1867,N_1938);
and U2055 (N_2055,N_1993,N_1920);
xor U2056 (N_2056,N_1911,N_1897);
nor U2057 (N_2057,N_1819,N_1894);
xor U2058 (N_2058,N_1986,N_1927);
nor U2059 (N_2059,N_1835,N_1901);
xnor U2060 (N_2060,N_1847,N_1902);
and U2061 (N_2061,N_1948,N_1809);
or U2062 (N_2062,N_1884,N_1954);
nand U2063 (N_2063,N_1863,N_1916);
xnor U2064 (N_2064,N_1936,N_1827);
nand U2065 (N_2065,N_1886,N_1862);
xnor U2066 (N_2066,N_1981,N_1830);
nor U2067 (N_2067,N_1962,N_1814);
and U2068 (N_2068,N_1839,N_1853);
nand U2069 (N_2069,N_1818,N_1888);
xor U2070 (N_2070,N_1859,N_1951);
or U2071 (N_2071,N_1845,N_1905);
xnor U2072 (N_2072,N_1896,N_1861);
and U2073 (N_2073,N_1968,N_1908);
or U2074 (N_2074,N_1846,N_1887);
nand U2075 (N_2075,N_1999,N_1971);
nor U2076 (N_2076,N_1929,N_1807);
or U2077 (N_2077,N_1813,N_1914);
nand U2078 (N_2078,N_1980,N_1840);
or U2079 (N_2079,N_1820,N_1934);
nor U2080 (N_2080,N_1838,N_1992);
nor U2081 (N_2081,N_1970,N_1931);
or U2082 (N_2082,N_1997,N_1848);
or U2083 (N_2083,N_1923,N_1831);
nand U2084 (N_2084,N_1803,N_1941);
or U2085 (N_2085,N_1963,N_1872);
xnor U2086 (N_2086,N_1922,N_1844);
or U2087 (N_2087,N_1979,N_1967);
xor U2088 (N_2088,N_1975,N_1972);
xnor U2089 (N_2089,N_1878,N_1821);
xnor U2090 (N_2090,N_1855,N_1823);
nor U2091 (N_2091,N_1933,N_1900);
or U2092 (N_2092,N_1898,N_1858);
nand U2093 (N_2093,N_1854,N_1924);
xor U2094 (N_2094,N_1942,N_1961);
or U2095 (N_2095,N_1939,N_1828);
nand U2096 (N_2096,N_1889,N_1893);
or U2097 (N_2097,N_1868,N_1895);
nand U2098 (N_2098,N_1930,N_1822);
xnor U2099 (N_2099,N_1956,N_1802);
or U2100 (N_2100,N_1846,N_1842);
nor U2101 (N_2101,N_1983,N_1838);
and U2102 (N_2102,N_1922,N_1959);
or U2103 (N_2103,N_1831,N_1843);
xnor U2104 (N_2104,N_1842,N_1816);
or U2105 (N_2105,N_1890,N_1803);
and U2106 (N_2106,N_1919,N_1838);
nand U2107 (N_2107,N_1853,N_1815);
xnor U2108 (N_2108,N_1948,N_1868);
or U2109 (N_2109,N_1856,N_1990);
nor U2110 (N_2110,N_1821,N_1936);
nand U2111 (N_2111,N_1877,N_1906);
and U2112 (N_2112,N_1839,N_1854);
nor U2113 (N_2113,N_1949,N_1851);
and U2114 (N_2114,N_1953,N_1887);
and U2115 (N_2115,N_1839,N_1947);
xor U2116 (N_2116,N_1949,N_1857);
or U2117 (N_2117,N_1901,N_1930);
nor U2118 (N_2118,N_1836,N_1961);
nor U2119 (N_2119,N_1860,N_1889);
nand U2120 (N_2120,N_1943,N_1994);
or U2121 (N_2121,N_1805,N_1809);
nor U2122 (N_2122,N_1890,N_1905);
nand U2123 (N_2123,N_1821,N_1861);
xnor U2124 (N_2124,N_1869,N_1938);
nor U2125 (N_2125,N_1994,N_1912);
nand U2126 (N_2126,N_1826,N_1948);
nor U2127 (N_2127,N_1941,N_1914);
or U2128 (N_2128,N_1816,N_1922);
xor U2129 (N_2129,N_1897,N_1979);
and U2130 (N_2130,N_1807,N_1882);
xnor U2131 (N_2131,N_1836,N_1859);
xor U2132 (N_2132,N_1840,N_1941);
xor U2133 (N_2133,N_1961,N_1878);
and U2134 (N_2134,N_1806,N_1921);
nor U2135 (N_2135,N_1872,N_1876);
and U2136 (N_2136,N_1989,N_1926);
xnor U2137 (N_2137,N_1890,N_1836);
xnor U2138 (N_2138,N_1919,N_1890);
nand U2139 (N_2139,N_1883,N_1829);
xor U2140 (N_2140,N_1985,N_1897);
nand U2141 (N_2141,N_1819,N_1871);
nand U2142 (N_2142,N_1846,N_1814);
nand U2143 (N_2143,N_1845,N_1958);
and U2144 (N_2144,N_1892,N_1843);
nand U2145 (N_2145,N_1841,N_1961);
xnor U2146 (N_2146,N_1826,N_1875);
xnor U2147 (N_2147,N_1807,N_1968);
nor U2148 (N_2148,N_1898,N_1986);
xnor U2149 (N_2149,N_1986,N_1952);
nor U2150 (N_2150,N_1965,N_1889);
xnor U2151 (N_2151,N_1981,N_1956);
or U2152 (N_2152,N_1824,N_1874);
or U2153 (N_2153,N_1819,N_1993);
xnor U2154 (N_2154,N_1854,N_1953);
xor U2155 (N_2155,N_1933,N_1941);
nand U2156 (N_2156,N_1949,N_1909);
xor U2157 (N_2157,N_1863,N_1890);
nor U2158 (N_2158,N_1988,N_1839);
or U2159 (N_2159,N_1842,N_1864);
and U2160 (N_2160,N_1949,N_1993);
xor U2161 (N_2161,N_1853,N_1879);
or U2162 (N_2162,N_1986,N_1843);
nor U2163 (N_2163,N_1926,N_1842);
or U2164 (N_2164,N_1965,N_1839);
and U2165 (N_2165,N_1944,N_1896);
nand U2166 (N_2166,N_1896,N_1855);
or U2167 (N_2167,N_1890,N_1962);
or U2168 (N_2168,N_1881,N_1970);
xnor U2169 (N_2169,N_1978,N_1967);
nor U2170 (N_2170,N_1815,N_1984);
or U2171 (N_2171,N_1904,N_1856);
and U2172 (N_2172,N_1916,N_1968);
xnor U2173 (N_2173,N_1868,N_1801);
nand U2174 (N_2174,N_1889,N_1958);
or U2175 (N_2175,N_1905,N_1919);
nand U2176 (N_2176,N_1874,N_1892);
nor U2177 (N_2177,N_1994,N_1944);
nand U2178 (N_2178,N_1945,N_1829);
xnor U2179 (N_2179,N_1901,N_1989);
and U2180 (N_2180,N_1868,N_1961);
and U2181 (N_2181,N_1880,N_1916);
xor U2182 (N_2182,N_1907,N_1985);
nand U2183 (N_2183,N_1897,N_1863);
nor U2184 (N_2184,N_1837,N_1843);
xor U2185 (N_2185,N_1885,N_1899);
nor U2186 (N_2186,N_1876,N_1998);
nor U2187 (N_2187,N_1892,N_1905);
nor U2188 (N_2188,N_1974,N_1800);
nand U2189 (N_2189,N_1894,N_1970);
nor U2190 (N_2190,N_1851,N_1843);
or U2191 (N_2191,N_1879,N_1831);
and U2192 (N_2192,N_1839,N_1811);
xnor U2193 (N_2193,N_1881,N_1910);
xor U2194 (N_2194,N_1822,N_1841);
nor U2195 (N_2195,N_1971,N_1845);
or U2196 (N_2196,N_1960,N_1940);
nand U2197 (N_2197,N_1997,N_1807);
or U2198 (N_2198,N_1998,N_1884);
nand U2199 (N_2199,N_1995,N_1935);
nor U2200 (N_2200,N_2016,N_2026);
nand U2201 (N_2201,N_2030,N_2053);
or U2202 (N_2202,N_2051,N_2127);
nand U2203 (N_2203,N_2007,N_2038);
or U2204 (N_2204,N_2090,N_2072);
nor U2205 (N_2205,N_2186,N_2155);
nor U2206 (N_2206,N_2075,N_2121);
nand U2207 (N_2207,N_2058,N_2138);
xor U2208 (N_2208,N_2180,N_2045);
nor U2209 (N_2209,N_2039,N_2130);
nor U2210 (N_2210,N_2035,N_2021);
nand U2211 (N_2211,N_2061,N_2123);
and U2212 (N_2212,N_2184,N_2082);
nor U2213 (N_2213,N_2119,N_2011);
nand U2214 (N_2214,N_2197,N_2163);
nand U2215 (N_2215,N_2086,N_2176);
nor U2216 (N_2216,N_2098,N_2084);
nand U2217 (N_2217,N_2027,N_2073);
or U2218 (N_2218,N_2151,N_2063);
nand U2219 (N_2219,N_2042,N_2081);
nor U2220 (N_2220,N_2020,N_2187);
and U2221 (N_2221,N_2141,N_2158);
nand U2222 (N_2222,N_2052,N_2004);
xnor U2223 (N_2223,N_2171,N_2164);
xor U2224 (N_2224,N_2024,N_2146);
nor U2225 (N_2225,N_2162,N_2143);
xnor U2226 (N_2226,N_2170,N_2196);
or U2227 (N_2227,N_2067,N_2116);
nor U2228 (N_2228,N_2077,N_2111);
nand U2229 (N_2229,N_2142,N_2165);
and U2230 (N_2230,N_2156,N_2074);
and U2231 (N_2231,N_2140,N_2161);
nand U2232 (N_2232,N_2008,N_2115);
or U2233 (N_2233,N_2055,N_2131);
or U2234 (N_2234,N_2124,N_2150);
nand U2235 (N_2235,N_2069,N_2071);
or U2236 (N_2236,N_2190,N_2023);
xor U2237 (N_2237,N_2166,N_2134);
xor U2238 (N_2238,N_2113,N_2152);
nand U2239 (N_2239,N_2110,N_2087);
nor U2240 (N_2240,N_2083,N_2109);
or U2241 (N_2241,N_2065,N_2188);
and U2242 (N_2242,N_2010,N_2006);
or U2243 (N_2243,N_2128,N_2037);
nor U2244 (N_2244,N_2080,N_2070);
nand U2245 (N_2245,N_2117,N_2018);
xor U2246 (N_2246,N_2047,N_2104);
xor U2247 (N_2247,N_2017,N_2044);
xor U2248 (N_2248,N_2107,N_2198);
and U2249 (N_2249,N_2172,N_2102);
xor U2250 (N_2250,N_2085,N_2112);
or U2251 (N_2251,N_2133,N_2033);
or U2252 (N_2252,N_2003,N_2101);
and U2253 (N_2253,N_2097,N_2029);
and U2254 (N_2254,N_2168,N_2174);
nand U2255 (N_2255,N_2091,N_2132);
nor U2256 (N_2256,N_2159,N_2129);
xor U2257 (N_2257,N_2108,N_2013);
nor U2258 (N_2258,N_2002,N_2157);
and U2259 (N_2259,N_2088,N_2145);
xnor U2260 (N_2260,N_2177,N_2034);
nand U2261 (N_2261,N_2175,N_2185);
and U2262 (N_2262,N_2022,N_2000);
nor U2263 (N_2263,N_2079,N_2094);
nand U2264 (N_2264,N_2005,N_2036);
xor U2265 (N_2265,N_2032,N_2193);
nor U2266 (N_2266,N_2153,N_2122);
nand U2267 (N_2267,N_2089,N_2114);
or U2268 (N_2268,N_2050,N_2173);
xor U2269 (N_2269,N_2059,N_2169);
or U2270 (N_2270,N_2056,N_2057);
nor U2271 (N_2271,N_2031,N_2178);
nand U2272 (N_2272,N_2120,N_2103);
or U2273 (N_2273,N_2105,N_2012);
nand U2274 (N_2274,N_2106,N_2040);
nand U2275 (N_2275,N_2066,N_2095);
nand U2276 (N_2276,N_2136,N_2078);
nand U2277 (N_2277,N_2096,N_2100);
xnor U2278 (N_2278,N_2014,N_2194);
nor U2279 (N_2279,N_2167,N_2179);
nor U2280 (N_2280,N_2025,N_2048);
or U2281 (N_2281,N_2093,N_2118);
nor U2282 (N_2282,N_2092,N_2064);
nand U2283 (N_2283,N_2147,N_2126);
nor U2284 (N_2284,N_2135,N_2144);
nor U2285 (N_2285,N_2076,N_2099);
and U2286 (N_2286,N_2148,N_2195);
nand U2287 (N_2287,N_2192,N_2199);
or U2288 (N_2288,N_2183,N_2181);
or U2289 (N_2289,N_2046,N_2062);
nand U2290 (N_2290,N_2054,N_2154);
or U2291 (N_2291,N_2125,N_2068);
nor U2292 (N_2292,N_2060,N_2149);
xor U2293 (N_2293,N_2182,N_2041);
nor U2294 (N_2294,N_2049,N_2015);
or U2295 (N_2295,N_2043,N_2139);
xnor U2296 (N_2296,N_2009,N_2191);
or U2297 (N_2297,N_2028,N_2137);
and U2298 (N_2298,N_2189,N_2019);
nor U2299 (N_2299,N_2001,N_2160);
xor U2300 (N_2300,N_2125,N_2051);
nor U2301 (N_2301,N_2148,N_2162);
xnor U2302 (N_2302,N_2134,N_2104);
or U2303 (N_2303,N_2116,N_2090);
nand U2304 (N_2304,N_2133,N_2024);
nand U2305 (N_2305,N_2059,N_2083);
nor U2306 (N_2306,N_2169,N_2063);
or U2307 (N_2307,N_2095,N_2092);
nand U2308 (N_2308,N_2161,N_2194);
nor U2309 (N_2309,N_2090,N_2118);
xnor U2310 (N_2310,N_2006,N_2166);
and U2311 (N_2311,N_2156,N_2127);
xor U2312 (N_2312,N_2133,N_2181);
and U2313 (N_2313,N_2138,N_2108);
xor U2314 (N_2314,N_2136,N_2162);
or U2315 (N_2315,N_2134,N_2047);
xor U2316 (N_2316,N_2080,N_2038);
and U2317 (N_2317,N_2026,N_2054);
or U2318 (N_2318,N_2121,N_2085);
nor U2319 (N_2319,N_2097,N_2039);
xnor U2320 (N_2320,N_2199,N_2069);
nand U2321 (N_2321,N_2015,N_2192);
or U2322 (N_2322,N_2166,N_2144);
or U2323 (N_2323,N_2155,N_2041);
and U2324 (N_2324,N_2024,N_2084);
nor U2325 (N_2325,N_2131,N_2043);
and U2326 (N_2326,N_2070,N_2029);
xnor U2327 (N_2327,N_2040,N_2099);
nor U2328 (N_2328,N_2118,N_2184);
xor U2329 (N_2329,N_2176,N_2182);
xor U2330 (N_2330,N_2031,N_2087);
nand U2331 (N_2331,N_2176,N_2000);
xor U2332 (N_2332,N_2012,N_2075);
nand U2333 (N_2333,N_2025,N_2152);
xor U2334 (N_2334,N_2110,N_2077);
xor U2335 (N_2335,N_2062,N_2155);
nand U2336 (N_2336,N_2044,N_2199);
xor U2337 (N_2337,N_2103,N_2076);
nand U2338 (N_2338,N_2063,N_2181);
and U2339 (N_2339,N_2161,N_2040);
xnor U2340 (N_2340,N_2124,N_2120);
and U2341 (N_2341,N_2056,N_2035);
nor U2342 (N_2342,N_2155,N_2013);
xnor U2343 (N_2343,N_2133,N_2064);
or U2344 (N_2344,N_2173,N_2096);
xnor U2345 (N_2345,N_2024,N_2088);
nand U2346 (N_2346,N_2060,N_2089);
nor U2347 (N_2347,N_2110,N_2185);
and U2348 (N_2348,N_2185,N_2133);
and U2349 (N_2349,N_2108,N_2186);
or U2350 (N_2350,N_2198,N_2084);
nand U2351 (N_2351,N_2001,N_2011);
or U2352 (N_2352,N_2082,N_2039);
and U2353 (N_2353,N_2192,N_2148);
nor U2354 (N_2354,N_2127,N_2114);
nor U2355 (N_2355,N_2135,N_2117);
nand U2356 (N_2356,N_2089,N_2138);
nand U2357 (N_2357,N_2150,N_2093);
xor U2358 (N_2358,N_2074,N_2110);
xor U2359 (N_2359,N_2013,N_2117);
nand U2360 (N_2360,N_2120,N_2119);
nand U2361 (N_2361,N_2152,N_2109);
nand U2362 (N_2362,N_2033,N_2127);
nor U2363 (N_2363,N_2073,N_2147);
nor U2364 (N_2364,N_2127,N_2190);
xor U2365 (N_2365,N_2075,N_2092);
or U2366 (N_2366,N_2165,N_2061);
nand U2367 (N_2367,N_2173,N_2071);
nand U2368 (N_2368,N_2176,N_2096);
xor U2369 (N_2369,N_2048,N_2111);
or U2370 (N_2370,N_2119,N_2020);
or U2371 (N_2371,N_2136,N_2130);
or U2372 (N_2372,N_2110,N_2199);
and U2373 (N_2373,N_2072,N_2199);
nand U2374 (N_2374,N_2174,N_2105);
nand U2375 (N_2375,N_2163,N_2042);
and U2376 (N_2376,N_2156,N_2080);
or U2377 (N_2377,N_2179,N_2198);
or U2378 (N_2378,N_2094,N_2089);
and U2379 (N_2379,N_2091,N_2061);
nand U2380 (N_2380,N_2129,N_2026);
or U2381 (N_2381,N_2046,N_2182);
and U2382 (N_2382,N_2073,N_2177);
nor U2383 (N_2383,N_2041,N_2023);
or U2384 (N_2384,N_2109,N_2147);
xor U2385 (N_2385,N_2167,N_2005);
xor U2386 (N_2386,N_2032,N_2033);
xor U2387 (N_2387,N_2045,N_2077);
xnor U2388 (N_2388,N_2135,N_2037);
and U2389 (N_2389,N_2178,N_2155);
nor U2390 (N_2390,N_2106,N_2006);
nor U2391 (N_2391,N_2130,N_2197);
nand U2392 (N_2392,N_2049,N_2121);
or U2393 (N_2393,N_2080,N_2096);
or U2394 (N_2394,N_2107,N_2019);
nand U2395 (N_2395,N_2109,N_2117);
or U2396 (N_2396,N_2076,N_2051);
nand U2397 (N_2397,N_2169,N_2123);
and U2398 (N_2398,N_2135,N_2181);
and U2399 (N_2399,N_2161,N_2007);
xor U2400 (N_2400,N_2286,N_2297);
nand U2401 (N_2401,N_2321,N_2384);
xnor U2402 (N_2402,N_2343,N_2211);
nor U2403 (N_2403,N_2280,N_2247);
xor U2404 (N_2404,N_2223,N_2373);
and U2405 (N_2405,N_2396,N_2354);
and U2406 (N_2406,N_2302,N_2331);
xnor U2407 (N_2407,N_2242,N_2225);
and U2408 (N_2408,N_2371,N_2393);
nand U2409 (N_2409,N_2271,N_2217);
and U2410 (N_2410,N_2287,N_2291);
nand U2411 (N_2411,N_2324,N_2257);
or U2412 (N_2412,N_2281,N_2227);
nand U2413 (N_2413,N_2215,N_2203);
nand U2414 (N_2414,N_2251,N_2221);
or U2415 (N_2415,N_2216,N_2289);
or U2416 (N_2416,N_2311,N_2261);
nor U2417 (N_2417,N_2220,N_2278);
or U2418 (N_2418,N_2334,N_2201);
nand U2419 (N_2419,N_2268,N_2323);
nor U2420 (N_2420,N_2341,N_2369);
nor U2421 (N_2421,N_2350,N_2347);
nor U2422 (N_2422,N_2330,N_2310);
and U2423 (N_2423,N_2243,N_2249);
nor U2424 (N_2424,N_2307,N_2274);
and U2425 (N_2425,N_2372,N_2344);
nor U2426 (N_2426,N_2277,N_2245);
nand U2427 (N_2427,N_2325,N_2218);
nand U2428 (N_2428,N_2362,N_2391);
nor U2429 (N_2429,N_2356,N_2288);
nand U2430 (N_2430,N_2241,N_2337);
or U2431 (N_2431,N_2386,N_2283);
xor U2432 (N_2432,N_2340,N_2208);
xnor U2433 (N_2433,N_2328,N_2359);
or U2434 (N_2434,N_2219,N_2226);
or U2435 (N_2435,N_2352,N_2316);
nor U2436 (N_2436,N_2317,N_2366);
nor U2437 (N_2437,N_2205,N_2230);
nor U2438 (N_2438,N_2282,N_2301);
xnor U2439 (N_2439,N_2200,N_2336);
nand U2440 (N_2440,N_2264,N_2304);
xor U2441 (N_2441,N_2231,N_2236);
or U2442 (N_2442,N_2240,N_2381);
xnor U2443 (N_2443,N_2228,N_2349);
and U2444 (N_2444,N_2364,N_2379);
or U2445 (N_2445,N_2399,N_2265);
or U2446 (N_2446,N_2390,N_2314);
or U2447 (N_2447,N_2296,N_2375);
or U2448 (N_2448,N_2284,N_2276);
xnor U2449 (N_2449,N_2235,N_2210);
nand U2450 (N_2450,N_2244,N_2374);
xor U2451 (N_2451,N_2239,N_2367);
nand U2452 (N_2452,N_2232,N_2285);
or U2453 (N_2453,N_2252,N_2273);
and U2454 (N_2454,N_2295,N_2353);
and U2455 (N_2455,N_2256,N_2275);
xor U2456 (N_2456,N_2229,N_2319);
xnor U2457 (N_2457,N_2299,N_2348);
xnor U2458 (N_2458,N_2212,N_2397);
and U2459 (N_2459,N_2389,N_2394);
nor U2460 (N_2460,N_2392,N_2315);
nand U2461 (N_2461,N_2300,N_2260);
nor U2462 (N_2462,N_2398,N_2254);
and U2463 (N_2463,N_2320,N_2233);
nand U2464 (N_2464,N_2370,N_2270);
or U2465 (N_2465,N_2395,N_2322);
or U2466 (N_2466,N_2207,N_2209);
or U2467 (N_2467,N_2238,N_2365);
nor U2468 (N_2468,N_2380,N_2318);
and U2469 (N_2469,N_2266,N_2292);
nor U2470 (N_2470,N_2262,N_2355);
xnor U2471 (N_2471,N_2358,N_2255);
or U2472 (N_2472,N_2339,N_2338);
xor U2473 (N_2473,N_2313,N_2378);
and U2474 (N_2474,N_2383,N_2222);
nand U2475 (N_2475,N_2346,N_2294);
nor U2476 (N_2476,N_2250,N_2345);
nand U2477 (N_2477,N_2388,N_2259);
nor U2478 (N_2478,N_2224,N_2368);
or U2479 (N_2479,N_2308,N_2312);
xnor U2480 (N_2480,N_2204,N_2214);
or U2481 (N_2481,N_2306,N_2290);
nand U2482 (N_2482,N_2327,N_2309);
and U2483 (N_2483,N_2361,N_2206);
xor U2484 (N_2484,N_2298,N_2234);
nor U2485 (N_2485,N_2246,N_2279);
nor U2486 (N_2486,N_2382,N_2360);
nor U2487 (N_2487,N_2351,N_2332);
nand U2488 (N_2488,N_2329,N_2272);
and U2489 (N_2489,N_2213,N_2326);
nand U2490 (N_2490,N_2335,N_2202);
xnor U2491 (N_2491,N_2385,N_2387);
and U2492 (N_2492,N_2269,N_2267);
or U2493 (N_2493,N_2357,N_2333);
and U2494 (N_2494,N_2305,N_2376);
nand U2495 (N_2495,N_2303,N_2248);
or U2496 (N_2496,N_2253,N_2293);
or U2497 (N_2497,N_2237,N_2377);
nor U2498 (N_2498,N_2258,N_2263);
or U2499 (N_2499,N_2363,N_2342);
nand U2500 (N_2500,N_2288,N_2236);
nand U2501 (N_2501,N_2326,N_2338);
nor U2502 (N_2502,N_2275,N_2361);
and U2503 (N_2503,N_2341,N_2334);
nor U2504 (N_2504,N_2252,N_2227);
xor U2505 (N_2505,N_2332,N_2205);
nor U2506 (N_2506,N_2292,N_2249);
nor U2507 (N_2507,N_2205,N_2350);
nand U2508 (N_2508,N_2368,N_2354);
nand U2509 (N_2509,N_2232,N_2319);
and U2510 (N_2510,N_2322,N_2257);
nor U2511 (N_2511,N_2399,N_2224);
or U2512 (N_2512,N_2245,N_2396);
nor U2513 (N_2513,N_2270,N_2390);
nand U2514 (N_2514,N_2362,N_2284);
nor U2515 (N_2515,N_2394,N_2238);
xnor U2516 (N_2516,N_2241,N_2375);
or U2517 (N_2517,N_2282,N_2298);
or U2518 (N_2518,N_2325,N_2347);
nor U2519 (N_2519,N_2220,N_2274);
nor U2520 (N_2520,N_2345,N_2204);
and U2521 (N_2521,N_2359,N_2332);
xor U2522 (N_2522,N_2256,N_2302);
and U2523 (N_2523,N_2209,N_2317);
or U2524 (N_2524,N_2232,N_2247);
or U2525 (N_2525,N_2202,N_2287);
and U2526 (N_2526,N_2317,N_2314);
nor U2527 (N_2527,N_2293,N_2376);
nand U2528 (N_2528,N_2268,N_2251);
and U2529 (N_2529,N_2385,N_2254);
or U2530 (N_2530,N_2200,N_2319);
xor U2531 (N_2531,N_2296,N_2339);
nand U2532 (N_2532,N_2228,N_2360);
nand U2533 (N_2533,N_2243,N_2366);
and U2534 (N_2534,N_2340,N_2359);
nand U2535 (N_2535,N_2266,N_2313);
and U2536 (N_2536,N_2365,N_2245);
or U2537 (N_2537,N_2334,N_2342);
nand U2538 (N_2538,N_2234,N_2208);
xnor U2539 (N_2539,N_2319,N_2256);
nor U2540 (N_2540,N_2348,N_2342);
and U2541 (N_2541,N_2230,N_2286);
nor U2542 (N_2542,N_2283,N_2245);
nor U2543 (N_2543,N_2222,N_2343);
nand U2544 (N_2544,N_2281,N_2373);
nand U2545 (N_2545,N_2372,N_2387);
nand U2546 (N_2546,N_2345,N_2377);
nor U2547 (N_2547,N_2305,N_2222);
and U2548 (N_2548,N_2264,N_2216);
xor U2549 (N_2549,N_2231,N_2369);
nor U2550 (N_2550,N_2252,N_2266);
and U2551 (N_2551,N_2271,N_2327);
or U2552 (N_2552,N_2356,N_2314);
nand U2553 (N_2553,N_2337,N_2216);
xnor U2554 (N_2554,N_2262,N_2316);
nand U2555 (N_2555,N_2354,N_2349);
and U2556 (N_2556,N_2260,N_2254);
or U2557 (N_2557,N_2312,N_2380);
or U2558 (N_2558,N_2255,N_2361);
nor U2559 (N_2559,N_2338,N_2303);
nor U2560 (N_2560,N_2346,N_2339);
nor U2561 (N_2561,N_2299,N_2388);
and U2562 (N_2562,N_2319,N_2209);
and U2563 (N_2563,N_2385,N_2216);
nor U2564 (N_2564,N_2283,N_2335);
nor U2565 (N_2565,N_2220,N_2275);
or U2566 (N_2566,N_2317,N_2287);
and U2567 (N_2567,N_2302,N_2338);
xor U2568 (N_2568,N_2216,N_2366);
nand U2569 (N_2569,N_2284,N_2397);
or U2570 (N_2570,N_2312,N_2399);
xor U2571 (N_2571,N_2281,N_2394);
nor U2572 (N_2572,N_2249,N_2379);
nor U2573 (N_2573,N_2395,N_2276);
xnor U2574 (N_2574,N_2282,N_2209);
xnor U2575 (N_2575,N_2376,N_2390);
nand U2576 (N_2576,N_2242,N_2316);
or U2577 (N_2577,N_2280,N_2376);
and U2578 (N_2578,N_2284,N_2373);
or U2579 (N_2579,N_2284,N_2314);
nand U2580 (N_2580,N_2284,N_2280);
or U2581 (N_2581,N_2360,N_2293);
nand U2582 (N_2582,N_2227,N_2218);
xnor U2583 (N_2583,N_2306,N_2295);
nand U2584 (N_2584,N_2262,N_2229);
nor U2585 (N_2585,N_2238,N_2368);
nor U2586 (N_2586,N_2277,N_2201);
xnor U2587 (N_2587,N_2395,N_2354);
and U2588 (N_2588,N_2229,N_2286);
nor U2589 (N_2589,N_2297,N_2296);
or U2590 (N_2590,N_2263,N_2391);
nand U2591 (N_2591,N_2306,N_2207);
nor U2592 (N_2592,N_2396,N_2303);
nand U2593 (N_2593,N_2368,N_2276);
xor U2594 (N_2594,N_2367,N_2279);
or U2595 (N_2595,N_2274,N_2246);
xor U2596 (N_2596,N_2332,N_2221);
or U2597 (N_2597,N_2237,N_2244);
xnor U2598 (N_2598,N_2204,N_2296);
nor U2599 (N_2599,N_2238,N_2219);
and U2600 (N_2600,N_2599,N_2428);
and U2601 (N_2601,N_2552,N_2475);
and U2602 (N_2602,N_2460,N_2593);
nand U2603 (N_2603,N_2544,N_2568);
xnor U2604 (N_2604,N_2554,N_2512);
nand U2605 (N_2605,N_2490,N_2556);
or U2606 (N_2606,N_2441,N_2470);
nor U2607 (N_2607,N_2455,N_2506);
or U2608 (N_2608,N_2476,N_2551);
or U2609 (N_2609,N_2561,N_2513);
nor U2610 (N_2610,N_2469,N_2411);
or U2611 (N_2611,N_2497,N_2493);
xor U2612 (N_2612,N_2539,N_2445);
and U2613 (N_2613,N_2545,N_2586);
and U2614 (N_2614,N_2520,N_2591);
or U2615 (N_2615,N_2427,N_2403);
or U2616 (N_2616,N_2590,N_2430);
xnor U2617 (N_2617,N_2564,N_2525);
nand U2618 (N_2618,N_2450,N_2436);
or U2619 (N_2619,N_2589,N_2404);
xor U2620 (N_2620,N_2482,N_2594);
xor U2621 (N_2621,N_2408,N_2565);
or U2622 (N_2622,N_2504,N_2446);
xnor U2623 (N_2623,N_2531,N_2402);
nor U2624 (N_2624,N_2465,N_2548);
nor U2625 (N_2625,N_2521,N_2412);
xor U2626 (N_2626,N_2543,N_2420);
xnor U2627 (N_2627,N_2517,N_2515);
or U2628 (N_2628,N_2487,N_2529);
and U2629 (N_2629,N_2588,N_2443);
nor U2630 (N_2630,N_2474,N_2547);
and U2631 (N_2631,N_2424,N_2486);
nand U2632 (N_2632,N_2527,N_2570);
nand U2633 (N_2633,N_2581,N_2549);
nand U2634 (N_2634,N_2562,N_2558);
and U2635 (N_2635,N_2598,N_2526);
nand U2636 (N_2636,N_2406,N_2414);
xnor U2637 (N_2637,N_2555,N_2505);
and U2638 (N_2638,N_2431,N_2473);
nand U2639 (N_2639,N_2439,N_2563);
nand U2640 (N_2640,N_2532,N_2458);
xnor U2641 (N_2641,N_2472,N_2560);
and U2642 (N_2642,N_2464,N_2478);
nor U2643 (N_2643,N_2550,N_2495);
or U2644 (N_2644,N_2422,N_2444);
and U2645 (N_2645,N_2442,N_2535);
or U2646 (N_2646,N_2440,N_2519);
or U2647 (N_2647,N_2530,N_2524);
xor U2648 (N_2648,N_2425,N_2438);
and U2649 (N_2649,N_2540,N_2534);
nor U2650 (N_2650,N_2468,N_2454);
nand U2651 (N_2651,N_2480,N_2522);
and U2652 (N_2652,N_2583,N_2511);
xor U2653 (N_2653,N_2418,N_2503);
nand U2654 (N_2654,N_2485,N_2566);
xor U2655 (N_2655,N_2456,N_2567);
or U2656 (N_2656,N_2433,N_2541);
nor U2657 (N_2657,N_2409,N_2553);
nand U2658 (N_2658,N_2523,N_2516);
or U2659 (N_2659,N_2575,N_2569);
nor U2660 (N_2660,N_2508,N_2514);
or U2661 (N_2661,N_2577,N_2538);
nand U2662 (N_2662,N_2559,N_2415);
xor U2663 (N_2663,N_2423,N_2489);
and U2664 (N_2664,N_2499,N_2466);
or U2665 (N_2665,N_2576,N_2587);
xnor U2666 (N_2666,N_2434,N_2571);
nor U2667 (N_2667,N_2447,N_2417);
and U2668 (N_2668,N_2405,N_2467);
nand U2669 (N_2669,N_2582,N_2481);
xnor U2670 (N_2670,N_2435,N_2410);
nand U2671 (N_2671,N_2462,N_2483);
nand U2672 (N_2672,N_2449,N_2537);
nand U2673 (N_2673,N_2510,N_2400);
xnor U2674 (N_2674,N_2471,N_2580);
nand U2675 (N_2675,N_2574,N_2597);
xor U2676 (N_2676,N_2484,N_2419);
nor U2677 (N_2677,N_2596,N_2572);
nor U2678 (N_2678,N_2461,N_2492);
or U2679 (N_2679,N_2584,N_2500);
or U2680 (N_2680,N_2498,N_2528);
xnor U2681 (N_2681,N_2502,N_2477);
or U2682 (N_2682,N_2421,N_2437);
or U2683 (N_2683,N_2557,N_2491);
and U2684 (N_2684,N_2451,N_2453);
and U2685 (N_2685,N_2536,N_2429);
nor U2686 (N_2686,N_2585,N_2579);
and U2687 (N_2687,N_2494,N_2542);
or U2688 (N_2688,N_2573,N_2413);
xor U2689 (N_2689,N_2459,N_2401);
and U2690 (N_2690,N_2592,N_2457);
nand U2691 (N_2691,N_2479,N_2496);
nand U2692 (N_2692,N_2509,N_2407);
xor U2693 (N_2693,N_2578,N_2432);
nand U2694 (N_2694,N_2501,N_2463);
nor U2695 (N_2695,N_2448,N_2533);
nand U2696 (N_2696,N_2518,N_2595);
xor U2697 (N_2697,N_2452,N_2546);
nand U2698 (N_2698,N_2416,N_2488);
nand U2699 (N_2699,N_2426,N_2507);
nand U2700 (N_2700,N_2485,N_2464);
nand U2701 (N_2701,N_2402,N_2429);
nand U2702 (N_2702,N_2480,N_2594);
and U2703 (N_2703,N_2549,N_2501);
nor U2704 (N_2704,N_2455,N_2444);
nand U2705 (N_2705,N_2585,N_2505);
or U2706 (N_2706,N_2550,N_2513);
nor U2707 (N_2707,N_2424,N_2592);
or U2708 (N_2708,N_2558,N_2411);
and U2709 (N_2709,N_2444,N_2441);
and U2710 (N_2710,N_2550,N_2430);
or U2711 (N_2711,N_2405,N_2403);
or U2712 (N_2712,N_2449,N_2581);
nand U2713 (N_2713,N_2586,N_2479);
or U2714 (N_2714,N_2433,N_2556);
or U2715 (N_2715,N_2484,N_2464);
and U2716 (N_2716,N_2413,N_2408);
and U2717 (N_2717,N_2575,N_2443);
or U2718 (N_2718,N_2416,N_2417);
nand U2719 (N_2719,N_2415,N_2489);
xnor U2720 (N_2720,N_2439,N_2465);
and U2721 (N_2721,N_2587,N_2434);
xor U2722 (N_2722,N_2530,N_2523);
and U2723 (N_2723,N_2476,N_2524);
and U2724 (N_2724,N_2433,N_2569);
or U2725 (N_2725,N_2569,N_2462);
and U2726 (N_2726,N_2540,N_2477);
nor U2727 (N_2727,N_2596,N_2599);
nand U2728 (N_2728,N_2476,N_2508);
xnor U2729 (N_2729,N_2504,N_2494);
nand U2730 (N_2730,N_2455,N_2417);
nand U2731 (N_2731,N_2511,N_2559);
xnor U2732 (N_2732,N_2504,N_2428);
nand U2733 (N_2733,N_2422,N_2449);
nor U2734 (N_2734,N_2456,N_2575);
nor U2735 (N_2735,N_2513,N_2452);
nor U2736 (N_2736,N_2431,N_2524);
and U2737 (N_2737,N_2427,N_2540);
nand U2738 (N_2738,N_2549,N_2418);
or U2739 (N_2739,N_2534,N_2542);
and U2740 (N_2740,N_2469,N_2458);
or U2741 (N_2741,N_2412,N_2413);
nand U2742 (N_2742,N_2532,N_2418);
or U2743 (N_2743,N_2577,N_2491);
nand U2744 (N_2744,N_2482,N_2502);
nor U2745 (N_2745,N_2557,N_2534);
nor U2746 (N_2746,N_2551,N_2588);
and U2747 (N_2747,N_2541,N_2532);
and U2748 (N_2748,N_2499,N_2566);
xor U2749 (N_2749,N_2551,N_2409);
nor U2750 (N_2750,N_2534,N_2520);
and U2751 (N_2751,N_2461,N_2597);
and U2752 (N_2752,N_2585,N_2475);
nand U2753 (N_2753,N_2500,N_2521);
or U2754 (N_2754,N_2557,N_2598);
and U2755 (N_2755,N_2482,N_2561);
nor U2756 (N_2756,N_2480,N_2443);
nor U2757 (N_2757,N_2465,N_2423);
nor U2758 (N_2758,N_2569,N_2531);
and U2759 (N_2759,N_2571,N_2517);
nor U2760 (N_2760,N_2410,N_2540);
nor U2761 (N_2761,N_2524,N_2517);
nor U2762 (N_2762,N_2556,N_2447);
and U2763 (N_2763,N_2425,N_2420);
nand U2764 (N_2764,N_2469,N_2596);
and U2765 (N_2765,N_2565,N_2560);
nor U2766 (N_2766,N_2509,N_2461);
or U2767 (N_2767,N_2558,N_2502);
nor U2768 (N_2768,N_2517,N_2500);
and U2769 (N_2769,N_2410,N_2525);
xor U2770 (N_2770,N_2408,N_2443);
nand U2771 (N_2771,N_2560,N_2493);
nand U2772 (N_2772,N_2527,N_2563);
nor U2773 (N_2773,N_2496,N_2485);
nor U2774 (N_2774,N_2537,N_2570);
or U2775 (N_2775,N_2529,N_2450);
nand U2776 (N_2776,N_2512,N_2429);
and U2777 (N_2777,N_2550,N_2510);
or U2778 (N_2778,N_2430,N_2463);
nand U2779 (N_2779,N_2511,N_2478);
and U2780 (N_2780,N_2401,N_2490);
nor U2781 (N_2781,N_2451,N_2537);
nand U2782 (N_2782,N_2517,N_2529);
xor U2783 (N_2783,N_2486,N_2464);
and U2784 (N_2784,N_2485,N_2411);
or U2785 (N_2785,N_2521,N_2481);
nor U2786 (N_2786,N_2481,N_2441);
or U2787 (N_2787,N_2590,N_2480);
xor U2788 (N_2788,N_2533,N_2532);
nand U2789 (N_2789,N_2432,N_2558);
or U2790 (N_2790,N_2528,N_2577);
and U2791 (N_2791,N_2463,N_2459);
or U2792 (N_2792,N_2452,N_2563);
xor U2793 (N_2793,N_2551,N_2545);
nor U2794 (N_2794,N_2537,N_2522);
xor U2795 (N_2795,N_2402,N_2516);
and U2796 (N_2796,N_2544,N_2494);
xor U2797 (N_2797,N_2515,N_2590);
xor U2798 (N_2798,N_2541,N_2463);
xnor U2799 (N_2799,N_2447,N_2502);
or U2800 (N_2800,N_2702,N_2746);
and U2801 (N_2801,N_2730,N_2708);
xnor U2802 (N_2802,N_2786,N_2707);
nand U2803 (N_2803,N_2682,N_2763);
xnor U2804 (N_2804,N_2605,N_2637);
and U2805 (N_2805,N_2737,N_2698);
xor U2806 (N_2806,N_2632,N_2614);
and U2807 (N_2807,N_2661,N_2743);
or U2808 (N_2808,N_2624,N_2695);
or U2809 (N_2809,N_2745,N_2700);
xor U2810 (N_2810,N_2710,N_2795);
nand U2811 (N_2811,N_2738,N_2753);
or U2812 (N_2812,N_2717,N_2623);
nor U2813 (N_2813,N_2780,N_2785);
xnor U2814 (N_2814,N_2756,N_2607);
and U2815 (N_2815,N_2754,N_2645);
or U2816 (N_2816,N_2705,N_2676);
or U2817 (N_2817,N_2663,N_2787);
xor U2818 (N_2818,N_2751,N_2742);
nor U2819 (N_2819,N_2651,N_2616);
nor U2820 (N_2820,N_2619,N_2770);
nor U2821 (N_2821,N_2715,N_2739);
and U2822 (N_2822,N_2627,N_2653);
nor U2823 (N_2823,N_2668,N_2779);
nor U2824 (N_2824,N_2631,N_2658);
nor U2825 (N_2825,N_2797,N_2720);
or U2826 (N_2826,N_2621,N_2610);
xnor U2827 (N_2827,N_2686,N_2703);
xnor U2828 (N_2828,N_2636,N_2733);
xnor U2829 (N_2829,N_2692,N_2602);
nor U2830 (N_2830,N_2618,N_2666);
nor U2831 (N_2831,N_2638,N_2647);
nand U2832 (N_2832,N_2600,N_2799);
or U2833 (N_2833,N_2630,N_2781);
xnor U2834 (N_2834,N_2687,N_2603);
and U2835 (N_2835,N_2758,N_2628);
xor U2836 (N_2836,N_2766,N_2713);
xor U2837 (N_2837,N_2723,N_2747);
nand U2838 (N_2838,N_2671,N_2721);
and U2839 (N_2839,N_2657,N_2792);
and U2840 (N_2840,N_2622,N_2772);
or U2841 (N_2841,N_2641,N_2725);
nand U2842 (N_2842,N_2634,N_2771);
or U2843 (N_2843,N_2709,N_2752);
xor U2844 (N_2844,N_2642,N_2776);
xor U2845 (N_2845,N_2654,N_2777);
or U2846 (N_2846,N_2635,N_2625);
nor U2847 (N_2847,N_2768,N_2727);
and U2848 (N_2848,N_2615,N_2793);
nand U2849 (N_2849,N_2646,N_2722);
or U2850 (N_2850,N_2644,N_2685);
and U2851 (N_2851,N_2704,N_2764);
or U2852 (N_2852,N_2794,N_2660);
nor U2853 (N_2853,N_2699,N_2665);
or U2854 (N_2854,N_2719,N_2664);
nor U2855 (N_2855,N_2788,N_2667);
nor U2856 (N_2856,N_2778,N_2690);
and U2857 (N_2857,N_2681,N_2640);
nor U2858 (N_2858,N_2675,N_2656);
xor U2859 (N_2859,N_2726,N_2711);
nand U2860 (N_2860,N_2798,N_2683);
nor U2861 (N_2861,N_2673,N_2782);
or U2862 (N_2862,N_2694,N_2652);
and U2863 (N_2863,N_2716,N_2796);
or U2864 (N_2864,N_2735,N_2612);
nand U2865 (N_2865,N_2769,N_2740);
or U2866 (N_2866,N_2744,N_2718);
nand U2867 (N_2867,N_2649,N_2749);
or U2868 (N_2868,N_2790,N_2655);
and U2869 (N_2869,N_2608,N_2791);
or U2870 (N_2870,N_2601,N_2750);
and U2871 (N_2871,N_2773,N_2762);
nand U2872 (N_2872,N_2693,N_2755);
or U2873 (N_2873,N_2669,N_2670);
xor U2874 (N_2874,N_2789,N_2650);
or U2875 (N_2875,N_2604,N_2748);
or U2876 (N_2876,N_2757,N_2678);
nor U2877 (N_2877,N_2774,N_2629);
and U2878 (N_2878,N_2677,N_2741);
nand U2879 (N_2879,N_2761,N_2767);
nor U2880 (N_2880,N_2728,N_2659);
xor U2881 (N_2881,N_2611,N_2759);
xor U2882 (N_2882,N_2760,N_2706);
nor U2883 (N_2883,N_2783,N_2696);
or U2884 (N_2884,N_2684,N_2674);
or U2885 (N_2885,N_2732,N_2714);
xor U2886 (N_2886,N_2620,N_2688);
xor U2887 (N_2887,N_2689,N_2672);
nor U2888 (N_2888,N_2648,N_2784);
nand U2889 (N_2889,N_2662,N_2712);
and U2890 (N_2890,N_2617,N_2613);
nand U2891 (N_2891,N_2729,N_2639);
nor U2892 (N_2892,N_2609,N_2680);
nand U2893 (N_2893,N_2765,N_2643);
xnor U2894 (N_2894,N_2736,N_2633);
nand U2895 (N_2895,N_2679,N_2691);
or U2896 (N_2896,N_2734,N_2626);
nand U2897 (N_2897,N_2606,N_2731);
and U2898 (N_2898,N_2697,N_2701);
nor U2899 (N_2899,N_2724,N_2775);
nor U2900 (N_2900,N_2644,N_2739);
nor U2901 (N_2901,N_2722,N_2719);
nor U2902 (N_2902,N_2677,N_2736);
xnor U2903 (N_2903,N_2640,N_2669);
nand U2904 (N_2904,N_2787,N_2714);
nor U2905 (N_2905,N_2683,N_2749);
and U2906 (N_2906,N_2673,N_2747);
xor U2907 (N_2907,N_2733,N_2658);
xor U2908 (N_2908,N_2719,N_2612);
nor U2909 (N_2909,N_2645,N_2637);
or U2910 (N_2910,N_2752,N_2605);
xnor U2911 (N_2911,N_2711,N_2626);
xnor U2912 (N_2912,N_2661,N_2613);
and U2913 (N_2913,N_2765,N_2637);
nand U2914 (N_2914,N_2636,N_2783);
or U2915 (N_2915,N_2690,N_2619);
nor U2916 (N_2916,N_2747,N_2645);
nand U2917 (N_2917,N_2609,N_2704);
xnor U2918 (N_2918,N_2645,N_2685);
nand U2919 (N_2919,N_2626,N_2735);
nor U2920 (N_2920,N_2611,N_2657);
nor U2921 (N_2921,N_2651,N_2650);
nand U2922 (N_2922,N_2768,N_2684);
and U2923 (N_2923,N_2650,N_2733);
xnor U2924 (N_2924,N_2782,N_2702);
nor U2925 (N_2925,N_2698,N_2656);
nand U2926 (N_2926,N_2697,N_2668);
and U2927 (N_2927,N_2658,N_2708);
nor U2928 (N_2928,N_2654,N_2776);
nor U2929 (N_2929,N_2674,N_2756);
and U2930 (N_2930,N_2602,N_2694);
xor U2931 (N_2931,N_2738,N_2611);
nand U2932 (N_2932,N_2726,N_2729);
and U2933 (N_2933,N_2662,N_2728);
xor U2934 (N_2934,N_2731,N_2796);
nor U2935 (N_2935,N_2650,N_2760);
nor U2936 (N_2936,N_2697,N_2635);
xnor U2937 (N_2937,N_2645,N_2646);
xnor U2938 (N_2938,N_2710,N_2786);
nor U2939 (N_2939,N_2626,N_2738);
and U2940 (N_2940,N_2754,N_2761);
nand U2941 (N_2941,N_2601,N_2727);
nand U2942 (N_2942,N_2731,N_2664);
and U2943 (N_2943,N_2790,N_2672);
nand U2944 (N_2944,N_2730,N_2738);
and U2945 (N_2945,N_2658,N_2721);
xor U2946 (N_2946,N_2774,N_2676);
nand U2947 (N_2947,N_2704,N_2767);
and U2948 (N_2948,N_2740,N_2749);
nand U2949 (N_2949,N_2742,N_2646);
or U2950 (N_2950,N_2754,N_2771);
nand U2951 (N_2951,N_2772,N_2711);
or U2952 (N_2952,N_2686,N_2721);
xor U2953 (N_2953,N_2739,N_2646);
or U2954 (N_2954,N_2611,N_2729);
nor U2955 (N_2955,N_2691,N_2662);
nor U2956 (N_2956,N_2634,N_2651);
and U2957 (N_2957,N_2629,N_2780);
or U2958 (N_2958,N_2722,N_2670);
or U2959 (N_2959,N_2701,N_2641);
xor U2960 (N_2960,N_2606,N_2755);
nand U2961 (N_2961,N_2649,N_2729);
or U2962 (N_2962,N_2664,N_2626);
xor U2963 (N_2963,N_2666,N_2732);
nor U2964 (N_2964,N_2670,N_2638);
nand U2965 (N_2965,N_2639,N_2735);
nor U2966 (N_2966,N_2702,N_2769);
nand U2967 (N_2967,N_2758,N_2684);
or U2968 (N_2968,N_2612,N_2642);
and U2969 (N_2969,N_2702,N_2759);
xor U2970 (N_2970,N_2751,N_2646);
nor U2971 (N_2971,N_2651,N_2657);
or U2972 (N_2972,N_2736,N_2756);
nand U2973 (N_2973,N_2639,N_2676);
nor U2974 (N_2974,N_2785,N_2662);
and U2975 (N_2975,N_2631,N_2789);
and U2976 (N_2976,N_2750,N_2656);
nor U2977 (N_2977,N_2630,N_2754);
nor U2978 (N_2978,N_2665,N_2730);
nand U2979 (N_2979,N_2736,N_2770);
or U2980 (N_2980,N_2635,N_2783);
nand U2981 (N_2981,N_2795,N_2648);
xor U2982 (N_2982,N_2684,N_2618);
xnor U2983 (N_2983,N_2754,N_2799);
and U2984 (N_2984,N_2773,N_2754);
xnor U2985 (N_2985,N_2704,N_2712);
nor U2986 (N_2986,N_2652,N_2756);
or U2987 (N_2987,N_2682,N_2795);
xnor U2988 (N_2988,N_2700,N_2704);
and U2989 (N_2989,N_2718,N_2770);
or U2990 (N_2990,N_2762,N_2638);
nor U2991 (N_2991,N_2782,N_2722);
nand U2992 (N_2992,N_2627,N_2639);
nor U2993 (N_2993,N_2760,N_2673);
xor U2994 (N_2994,N_2766,N_2608);
and U2995 (N_2995,N_2766,N_2748);
or U2996 (N_2996,N_2660,N_2698);
nand U2997 (N_2997,N_2667,N_2790);
or U2998 (N_2998,N_2789,N_2728);
xor U2999 (N_2999,N_2742,N_2700);
or U3000 (N_3000,N_2930,N_2814);
and U3001 (N_3001,N_2804,N_2836);
and U3002 (N_3002,N_2897,N_2988);
and U3003 (N_3003,N_2900,N_2828);
nand U3004 (N_3004,N_2990,N_2980);
and U3005 (N_3005,N_2856,N_2840);
nor U3006 (N_3006,N_2855,N_2895);
nand U3007 (N_3007,N_2934,N_2971);
nor U3008 (N_3008,N_2904,N_2819);
nand U3009 (N_3009,N_2929,N_2834);
xnor U3010 (N_3010,N_2801,N_2974);
xnor U3011 (N_3011,N_2953,N_2908);
or U3012 (N_3012,N_2941,N_2898);
nand U3013 (N_3013,N_2920,N_2818);
or U3014 (N_3014,N_2885,N_2862);
xnor U3015 (N_3015,N_2910,N_2865);
nor U3016 (N_3016,N_2997,N_2917);
nand U3017 (N_3017,N_2803,N_2926);
nor U3018 (N_3018,N_2939,N_2868);
nor U3019 (N_3019,N_2924,N_2972);
nand U3020 (N_3020,N_2809,N_2861);
nor U3021 (N_3021,N_2876,N_2902);
and U3022 (N_3022,N_2956,N_2932);
nand U3023 (N_3023,N_2874,N_2817);
and U3024 (N_3024,N_2979,N_2882);
or U3025 (N_3025,N_2950,N_2849);
nor U3026 (N_3026,N_2806,N_2984);
and U3027 (N_3027,N_2987,N_2867);
xor U3028 (N_3028,N_2852,N_2948);
xnor U3029 (N_3029,N_2824,N_2883);
nor U3030 (N_3030,N_2909,N_2927);
and U3031 (N_3031,N_2802,N_2976);
or U3032 (N_3032,N_2966,N_2843);
and U3033 (N_3033,N_2944,N_2866);
and U3034 (N_3034,N_2813,N_2918);
and U3035 (N_3035,N_2854,N_2845);
nor U3036 (N_3036,N_2848,N_2998);
nor U3037 (N_3037,N_2815,N_2901);
or U3038 (N_3038,N_2969,N_2820);
nor U3039 (N_3039,N_2911,N_2928);
and U3040 (N_3040,N_2915,N_2823);
xor U3041 (N_3041,N_2933,N_2850);
xnor U3042 (N_3042,N_2916,N_2838);
nor U3043 (N_3043,N_2958,N_2835);
nand U3044 (N_3044,N_2912,N_2903);
nand U3045 (N_3045,N_2955,N_2986);
xnor U3046 (N_3046,N_2875,N_2921);
or U3047 (N_3047,N_2860,N_2957);
nand U3048 (N_3048,N_2978,N_2935);
xor U3049 (N_3049,N_2800,N_2888);
xnor U3050 (N_3050,N_2894,N_2946);
nand U3051 (N_3051,N_2816,N_2870);
and U3052 (N_3052,N_2880,N_2983);
or U3053 (N_3053,N_2973,N_2994);
and U3054 (N_3054,N_2832,N_2942);
and U3055 (N_3055,N_2938,N_2877);
and U3056 (N_3056,N_2991,N_2847);
xnor U3057 (N_3057,N_2830,N_2826);
xor U3058 (N_3058,N_2853,N_2831);
xor U3059 (N_3059,N_2959,N_2945);
xnor U3060 (N_3060,N_2937,N_2881);
nor U3061 (N_3061,N_2869,N_2822);
nand U3062 (N_3062,N_2837,N_2851);
xnor U3063 (N_3063,N_2951,N_2812);
or U3064 (N_3064,N_2841,N_2947);
or U3065 (N_3065,N_2906,N_2872);
xor U3066 (N_3066,N_2879,N_2954);
and U3067 (N_3067,N_2949,N_2977);
nand U3068 (N_3068,N_2846,N_2981);
nor U3069 (N_3069,N_2863,N_2962);
nor U3070 (N_3070,N_2985,N_2923);
nor U3071 (N_3071,N_2996,N_2825);
nor U3072 (N_3072,N_2913,N_2891);
or U3073 (N_3073,N_2961,N_2952);
xor U3074 (N_3074,N_2992,N_2960);
nor U3075 (N_3075,N_2931,N_2964);
or U3076 (N_3076,N_2968,N_2975);
nand U3077 (N_3077,N_2967,N_2886);
nand U3078 (N_3078,N_2873,N_2982);
or U3079 (N_3079,N_2811,N_2892);
xor U3080 (N_3080,N_2833,N_2807);
nor U3081 (N_3081,N_2993,N_2859);
or U3082 (N_3082,N_2936,N_2890);
nor U3083 (N_3083,N_2995,N_2899);
or U3084 (N_3084,N_2827,N_2871);
and U3085 (N_3085,N_2810,N_2857);
xor U3086 (N_3086,N_2842,N_2905);
xor U3087 (N_3087,N_2887,N_2858);
or U3088 (N_3088,N_2963,N_2922);
nor U3089 (N_3089,N_2878,N_2925);
xnor U3090 (N_3090,N_2829,N_2805);
xnor U3091 (N_3091,N_2965,N_2884);
and U3092 (N_3092,N_2999,N_2970);
xnor U3093 (N_3093,N_2896,N_2940);
or U3094 (N_3094,N_2821,N_2844);
xor U3095 (N_3095,N_2989,N_2919);
xor U3096 (N_3096,N_2943,N_2914);
or U3097 (N_3097,N_2864,N_2893);
and U3098 (N_3098,N_2889,N_2907);
nor U3099 (N_3099,N_2839,N_2808);
nor U3100 (N_3100,N_2907,N_2952);
or U3101 (N_3101,N_2823,N_2913);
or U3102 (N_3102,N_2991,N_2948);
nor U3103 (N_3103,N_2881,N_2996);
or U3104 (N_3104,N_2901,N_2930);
or U3105 (N_3105,N_2862,N_2865);
or U3106 (N_3106,N_2835,N_2840);
or U3107 (N_3107,N_2976,N_2954);
nor U3108 (N_3108,N_2903,N_2823);
xor U3109 (N_3109,N_2873,N_2839);
or U3110 (N_3110,N_2880,N_2827);
nand U3111 (N_3111,N_2811,N_2874);
and U3112 (N_3112,N_2885,N_2817);
nor U3113 (N_3113,N_2969,N_2942);
and U3114 (N_3114,N_2811,N_2946);
nand U3115 (N_3115,N_2906,N_2881);
or U3116 (N_3116,N_2911,N_2984);
xnor U3117 (N_3117,N_2980,N_2947);
xnor U3118 (N_3118,N_2988,N_2942);
nand U3119 (N_3119,N_2959,N_2974);
xor U3120 (N_3120,N_2949,N_2971);
nand U3121 (N_3121,N_2922,N_2995);
nor U3122 (N_3122,N_2973,N_2917);
nor U3123 (N_3123,N_2949,N_2829);
or U3124 (N_3124,N_2993,N_2848);
or U3125 (N_3125,N_2824,N_2927);
nand U3126 (N_3126,N_2872,N_2963);
and U3127 (N_3127,N_2838,N_2994);
xor U3128 (N_3128,N_2835,N_2970);
and U3129 (N_3129,N_2905,N_2935);
nand U3130 (N_3130,N_2970,N_2951);
xnor U3131 (N_3131,N_2856,N_2921);
nor U3132 (N_3132,N_2822,N_2880);
or U3133 (N_3133,N_2923,N_2880);
or U3134 (N_3134,N_2984,N_2936);
and U3135 (N_3135,N_2918,N_2942);
nand U3136 (N_3136,N_2888,N_2875);
nand U3137 (N_3137,N_2901,N_2805);
or U3138 (N_3138,N_2892,N_2838);
nor U3139 (N_3139,N_2956,N_2906);
or U3140 (N_3140,N_2921,N_2944);
and U3141 (N_3141,N_2920,N_2944);
or U3142 (N_3142,N_2925,N_2801);
or U3143 (N_3143,N_2960,N_2860);
nor U3144 (N_3144,N_2833,N_2800);
and U3145 (N_3145,N_2987,N_2922);
nand U3146 (N_3146,N_2851,N_2958);
nor U3147 (N_3147,N_2805,N_2953);
xnor U3148 (N_3148,N_2861,N_2984);
and U3149 (N_3149,N_2958,N_2933);
nor U3150 (N_3150,N_2905,N_2999);
and U3151 (N_3151,N_2897,N_2972);
nor U3152 (N_3152,N_2909,N_2900);
or U3153 (N_3153,N_2900,N_2988);
or U3154 (N_3154,N_2876,N_2964);
nand U3155 (N_3155,N_2930,N_2899);
xnor U3156 (N_3156,N_2967,N_2870);
or U3157 (N_3157,N_2922,N_2929);
and U3158 (N_3158,N_2913,N_2979);
nand U3159 (N_3159,N_2867,N_2863);
nor U3160 (N_3160,N_2873,N_2901);
or U3161 (N_3161,N_2894,N_2989);
nand U3162 (N_3162,N_2838,N_2873);
or U3163 (N_3163,N_2809,N_2937);
or U3164 (N_3164,N_2881,N_2894);
nor U3165 (N_3165,N_2923,N_2852);
or U3166 (N_3166,N_2948,N_2862);
and U3167 (N_3167,N_2823,N_2898);
or U3168 (N_3168,N_2821,N_2840);
and U3169 (N_3169,N_2964,N_2973);
and U3170 (N_3170,N_2940,N_2906);
nand U3171 (N_3171,N_2961,N_2906);
and U3172 (N_3172,N_2962,N_2810);
nand U3173 (N_3173,N_2896,N_2860);
nor U3174 (N_3174,N_2994,N_2872);
or U3175 (N_3175,N_2931,N_2870);
and U3176 (N_3176,N_2936,N_2840);
nand U3177 (N_3177,N_2825,N_2883);
xor U3178 (N_3178,N_2813,N_2845);
xor U3179 (N_3179,N_2922,N_2818);
or U3180 (N_3180,N_2887,N_2802);
or U3181 (N_3181,N_2984,N_2823);
nor U3182 (N_3182,N_2812,N_2824);
nand U3183 (N_3183,N_2828,N_2801);
xnor U3184 (N_3184,N_2848,N_2844);
nand U3185 (N_3185,N_2839,N_2835);
xnor U3186 (N_3186,N_2876,N_2909);
nor U3187 (N_3187,N_2836,N_2854);
and U3188 (N_3188,N_2937,N_2815);
nand U3189 (N_3189,N_2807,N_2828);
xnor U3190 (N_3190,N_2976,N_2883);
xor U3191 (N_3191,N_2935,N_2847);
and U3192 (N_3192,N_2809,N_2900);
xnor U3193 (N_3193,N_2907,N_2881);
and U3194 (N_3194,N_2825,N_2988);
nand U3195 (N_3195,N_2977,N_2849);
nor U3196 (N_3196,N_2890,N_2904);
nor U3197 (N_3197,N_2871,N_2894);
and U3198 (N_3198,N_2813,N_2968);
and U3199 (N_3199,N_2898,N_2817);
xnor U3200 (N_3200,N_3156,N_3182);
nor U3201 (N_3201,N_3036,N_3013);
xnor U3202 (N_3202,N_3078,N_3059);
xor U3203 (N_3203,N_3108,N_3189);
xor U3204 (N_3204,N_3174,N_3141);
nor U3205 (N_3205,N_3090,N_3019);
nor U3206 (N_3206,N_3129,N_3155);
and U3207 (N_3207,N_3198,N_3065);
nand U3208 (N_3208,N_3143,N_3011);
xnor U3209 (N_3209,N_3096,N_3180);
nor U3210 (N_3210,N_3058,N_3023);
nand U3211 (N_3211,N_3002,N_3161);
and U3212 (N_3212,N_3068,N_3124);
and U3213 (N_3213,N_3111,N_3004);
nor U3214 (N_3214,N_3031,N_3063);
xor U3215 (N_3215,N_3089,N_3020);
nand U3216 (N_3216,N_3103,N_3092);
nor U3217 (N_3217,N_3107,N_3098);
xor U3218 (N_3218,N_3018,N_3024);
nand U3219 (N_3219,N_3120,N_3010);
or U3220 (N_3220,N_3052,N_3177);
or U3221 (N_3221,N_3115,N_3191);
xnor U3222 (N_3222,N_3147,N_3076);
xnor U3223 (N_3223,N_3151,N_3194);
xnor U3224 (N_3224,N_3122,N_3051);
nor U3225 (N_3225,N_3038,N_3171);
xnor U3226 (N_3226,N_3088,N_3094);
nor U3227 (N_3227,N_3037,N_3150);
or U3228 (N_3228,N_3164,N_3184);
nor U3229 (N_3229,N_3170,N_3101);
and U3230 (N_3230,N_3160,N_3095);
and U3231 (N_3231,N_3033,N_3116);
nand U3232 (N_3232,N_3022,N_3032);
and U3233 (N_3233,N_3025,N_3006);
or U3234 (N_3234,N_3030,N_3181);
xnor U3235 (N_3235,N_3162,N_3043);
xor U3236 (N_3236,N_3159,N_3126);
nand U3237 (N_3237,N_3087,N_3130);
nand U3238 (N_3238,N_3127,N_3080);
nor U3239 (N_3239,N_3121,N_3119);
nor U3240 (N_3240,N_3142,N_3028);
nand U3241 (N_3241,N_3081,N_3075);
or U3242 (N_3242,N_3153,N_3082);
nand U3243 (N_3243,N_3035,N_3166);
xnor U3244 (N_3244,N_3050,N_3085);
nor U3245 (N_3245,N_3134,N_3154);
xor U3246 (N_3246,N_3079,N_3099);
and U3247 (N_3247,N_3117,N_3000);
nor U3248 (N_3248,N_3179,N_3072);
nor U3249 (N_3249,N_3172,N_3001);
and U3250 (N_3250,N_3186,N_3026);
nand U3251 (N_3251,N_3086,N_3062);
and U3252 (N_3252,N_3047,N_3040);
and U3253 (N_3253,N_3183,N_3145);
nand U3254 (N_3254,N_3027,N_3015);
and U3255 (N_3255,N_3137,N_3128);
nor U3256 (N_3256,N_3014,N_3021);
nor U3257 (N_3257,N_3056,N_3138);
and U3258 (N_3258,N_3048,N_3069);
xnor U3259 (N_3259,N_3034,N_3070);
nor U3260 (N_3260,N_3054,N_3167);
or U3261 (N_3261,N_3199,N_3046);
nand U3262 (N_3262,N_3060,N_3123);
nor U3263 (N_3263,N_3148,N_3144);
or U3264 (N_3264,N_3178,N_3003);
nor U3265 (N_3265,N_3196,N_3193);
nor U3266 (N_3266,N_3114,N_3192);
nand U3267 (N_3267,N_3039,N_3017);
and U3268 (N_3268,N_3016,N_3008);
nand U3269 (N_3269,N_3113,N_3173);
or U3270 (N_3270,N_3175,N_3149);
nand U3271 (N_3271,N_3045,N_3100);
nor U3272 (N_3272,N_3135,N_3074);
or U3273 (N_3273,N_3110,N_3139);
or U3274 (N_3274,N_3152,N_3146);
and U3275 (N_3275,N_3168,N_3157);
and U3276 (N_3276,N_3187,N_3163);
xnor U3277 (N_3277,N_3071,N_3109);
nand U3278 (N_3278,N_3073,N_3140);
xor U3279 (N_3279,N_3102,N_3125);
and U3280 (N_3280,N_3097,N_3197);
or U3281 (N_3281,N_3136,N_3112);
xnor U3282 (N_3282,N_3169,N_3055);
nor U3283 (N_3283,N_3133,N_3093);
xnor U3284 (N_3284,N_3195,N_3105);
nand U3285 (N_3285,N_3057,N_3053);
nand U3286 (N_3286,N_3165,N_3083);
and U3287 (N_3287,N_3061,N_3044);
nor U3288 (N_3288,N_3188,N_3176);
nand U3289 (N_3289,N_3066,N_3005);
and U3290 (N_3290,N_3009,N_3012);
and U3291 (N_3291,N_3077,N_3084);
xnor U3292 (N_3292,N_3067,N_3190);
nor U3293 (N_3293,N_3091,N_3118);
nand U3294 (N_3294,N_3029,N_3132);
or U3295 (N_3295,N_3185,N_3106);
nand U3296 (N_3296,N_3131,N_3041);
and U3297 (N_3297,N_3064,N_3104);
nor U3298 (N_3298,N_3042,N_3049);
nand U3299 (N_3299,N_3007,N_3158);
nand U3300 (N_3300,N_3016,N_3170);
xor U3301 (N_3301,N_3134,N_3099);
and U3302 (N_3302,N_3016,N_3006);
xnor U3303 (N_3303,N_3063,N_3181);
or U3304 (N_3304,N_3036,N_3056);
nand U3305 (N_3305,N_3190,N_3071);
xor U3306 (N_3306,N_3080,N_3110);
nor U3307 (N_3307,N_3144,N_3170);
and U3308 (N_3308,N_3098,N_3057);
or U3309 (N_3309,N_3052,N_3050);
and U3310 (N_3310,N_3005,N_3197);
nor U3311 (N_3311,N_3138,N_3049);
and U3312 (N_3312,N_3164,N_3148);
or U3313 (N_3313,N_3138,N_3039);
or U3314 (N_3314,N_3132,N_3104);
xor U3315 (N_3315,N_3061,N_3013);
or U3316 (N_3316,N_3171,N_3183);
and U3317 (N_3317,N_3142,N_3143);
nand U3318 (N_3318,N_3022,N_3044);
nand U3319 (N_3319,N_3051,N_3147);
nor U3320 (N_3320,N_3139,N_3071);
and U3321 (N_3321,N_3099,N_3155);
or U3322 (N_3322,N_3005,N_3010);
nor U3323 (N_3323,N_3041,N_3185);
nand U3324 (N_3324,N_3081,N_3018);
nand U3325 (N_3325,N_3132,N_3141);
xnor U3326 (N_3326,N_3145,N_3185);
xor U3327 (N_3327,N_3128,N_3092);
or U3328 (N_3328,N_3027,N_3199);
xor U3329 (N_3329,N_3067,N_3124);
nand U3330 (N_3330,N_3121,N_3196);
and U3331 (N_3331,N_3071,N_3111);
nor U3332 (N_3332,N_3078,N_3188);
xor U3333 (N_3333,N_3072,N_3125);
nand U3334 (N_3334,N_3185,N_3053);
xor U3335 (N_3335,N_3090,N_3145);
nand U3336 (N_3336,N_3061,N_3134);
or U3337 (N_3337,N_3029,N_3184);
xnor U3338 (N_3338,N_3071,N_3122);
and U3339 (N_3339,N_3062,N_3194);
xnor U3340 (N_3340,N_3038,N_3072);
or U3341 (N_3341,N_3177,N_3060);
nand U3342 (N_3342,N_3175,N_3081);
or U3343 (N_3343,N_3049,N_3118);
xor U3344 (N_3344,N_3081,N_3128);
xnor U3345 (N_3345,N_3022,N_3087);
or U3346 (N_3346,N_3002,N_3042);
nand U3347 (N_3347,N_3030,N_3155);
and U3348 (N_3348,N_3094,N_3055);
nand U3349 (N_3349,N_3134,N_3072);
and U3350 (N_3350,N_3042,N_3138);
nor U3351 (N_3351,N_3011,N_3131);
nor U3352 (N_3352,N_3177,N_3006);
and U3353 (N_3353,N_3141,N_3013);
nor U3354 (N_3354,N_3141,N_3053);
nand U3355 (N_3355,N_3087,N_3000);
or U3356 (N_3356,N_3074,N_3078);
or U3357 (N_3357,N_3109,N_3031);
and U3358 (N_3358,N_3158,N_3153);
or U3359 (N_3359,N_3089,N_3048);
xnor U3360 (N_3360,N_3004,N_3169);
or U3361 (N_3361,N_3008,N_3166);
nor U3362 (N_3362,N_3063,N_3173);
xor U3363 (N_3363,N_3184,N_3150);
xor U3364 (N_3364,N_3144,N_3057);
xor U3365 (N_3365,N_3092,N_3154);
or U3366 (N_3366,N_3055,N_3172);
and U3367 (N_3367,N_3174,N_3033);
xnor U3368 (N_3368,N_3042,N_3070);
xor U3369 (N_3369,N_3130,N_3077);
and U3370 (N_3370,N_3197,N_3178);
xnor U3371 (N_3371,N_3024,N_3180);
xnor U3372 (N_3372,N_3056,N_3049);
or U3373 (N_3373,N_3059,N_3021);
nor U3374 (N_3374,N_3111,N_3137);
nand U3375 (N_3375,N_3052,N_3060);
or U3376 (N_3376,N_3142,N_3169);
or U3377 (N_3377,N_3158,N_3004);
xnor U3378 (N_3378,N_3150,N_3154);
nand U3379 (N_3379,N_3005,N_3185);
or U3380 (N_3380,N_3182,N_3035);
xor U3381 (N_3381,N_3162,N_3051);
and U3382 (N_3382,N_3170,N_3093);
nor U3383 (N_3383,N_3004,N_3082);
xnor U3384 (N_3384,N_3037,N_3160);
nand U3385 (N_3385,N_3046,N_3111);
nand U3386 (N_3386,N_3080,N_3165);
xnor U3387 (N_3387,N_3111,N_3053);
xor U3388 (N_3388,N_3058,N_3108);
nor U3389 (N_3389,N_3086,N_3130);
nand U3390 (N_3390,N_3035,N_3189);
nand U3391 (N_3391,N_3126,N_3064);
nand U3392 (N_3392,N_3152,N_3113);
xnor U3393 (N_3393,N_3163,N_3189);
and U3394 (N_3394,N_3052,N_3020);
or U3395 (N_3395,N_3164,N_3142);
and U3396 (N_3396,N_3145,N_3122);
nor U3397 (N_3397,N_3132,N_3090);
or U3398 (N_3398,N_3136,N_3061);
nand U3399 (N_3399,N_3026,N_3151);
nand U3400 (N_3400,N_3372,N_3244);
or U3401 (N_3401,N_3376,N_3206);
nor U3402 (N_3402,N_3219,N_3290);
nand U3403 (N_3403,N_3297,N_3200);
or U3404 (N_3404,N_3288,N_3271);
xor U3405 (N_3405,N_3229,N_3242);
xor U3406 (N_3406,N_3260,N_3396);
nand U3407 (N_3407,N_3309,N_3385);
xor U3408 (N_3408,N_3388,N_3319);
and U3409 (N_3409,N_3258,N_3276);
and U3410 (N_3410,N_3380,N_3212);
and U3411 (N_3411,N_3291,N_3217);
nand U3412 (N_3412,N_3213,N_3381);
xor U3413 (N_3413,N_3216,N_3337);
nand U3414 (N_3414,N_3354,N_3361);
xor U3415 (N_3415,N_3312,N_3253);
and U3416 (N_3416,N_3329,N_3320);
nor U3417 (N_3417,N_3239,N_3268);
or U3418 (N_3418,N_3371,N_3339);
or U3419 (N_3419,N_3259,N_3221);
xnor U3420 (N_3420,N_3318,N_3278);
xor U3421 (N_3421,N_3334,N_3275);
nor U3422 (N_3422,N_3323,N_3251);
nor U3423 (N_3423,N_3296,N_3340);
nand U3424 (N_3424,N_3250,N_3370);
and U3425 (N_3425,N_3220,N_3395);
nand U3426 (N_3426,N_3285,N_3365);
nand U3427 (N_3427,N_3204,N_3351);
and U3428 (N_3428,N_3358,N_3224);
and U3429 (N_3429,N_3336,N_3349);
or U3430 (N_3430,N_3305,N_3232);
nor U3431 (N_3431,N_3369,N_3310);
and U3432 (N_3432,N_3227,N_3246);
and U3433 (N_3433,N_3324,N_3367);
nand U3434 (N_3434,N_3211,N_3243);
and U3435 (N_3435,N_3269,N_3287);
nand U3436 (N_3436,N_3386,N_3325);
or U3437 (N_3437,N_3399,N_3373);
and U3438 (N_3438,N_3267,N_3279);
nor U3439 (N_3439,N_3207,N_3289);
xnor U3440 (N_3440,N_3222,N_3214);
nor U3441 (N_3441,N_3352,N_3378);
xnor U3442 (N_3442,N_3231,N_3353);
nand U3443 (N_3443,N_3233,N_3355);
nand U3444 (N_3444,N_3256,N_3299);
or U3445 (N_3445,N_3298,N_3238);
or U3446 (N_3446,N_3248,N_3374);
xnor U3447 (N_3447,N_3247,N_3317);
and U3448 (N_3448,N_3368,N_3341);
nor U3449 (N_3449,N_3311,N_3280);
nand U3450 (N_3450,N_3350,N_3328);
nor U3451 (N_3451,N_3326,N_3223);
xnor U3452 (N_3452,N_3230,N_3215);
nand U3453 (N_3453,N_3241,N_3286);
or U3454 (N_3454,N_3252,N_3272);
or U3455 (N_3455,N_3363,N_3281);
xor U3456 (N_3456,N_3240,N_3270);
or U3457 (N_3457,N_3307,N_3282);
nand U3458 (N_3458,N_3321,N_3342);
or U3459 (N_3459,N_3273,N_3393);
and U3460 (N_3460,N_3234,N_3218);
xnor U3461 (N_3461,N_3346,N_3284);
xnor U3462 (N_3462,N_3316,N_3201);
nand U3463 (N_3463,N_3263,N_3283);
xnor U3464 (N_3464,N_3375,N_3356);
or U3465 (N_3465,N_3394,N_3387);
and U3466 (N_3466,N_3235,N_3266);
and U3467 (N_3467,N_3357,N_3254);
nand U3468 (N_3468,N_3315,N_3236);
and U3469 (N_3469,N_3277,N_3333);
and U3470 (N_3470,N_3257,N_3262);
xor U3471 (N_3471,N_3382,N_3265);
or U3472 (N_3472,N_3314,N_3377);
nor U3473 (N_3473,N_3237,N_3332);
and U3474 (N_3474,N_3303,N_3274);
nand U3475 (N_3475,N_3292,N_3392);
and U3476 (N_3476,N_3383,N_3360);
nor U3477 (N_3477,N_3245,N_3344);
and U3478 (N_3478,N_3379,N_3210);
and U3479 (N_3479,N_3327,N_3389);
nor U3480 (N_3480,N_3362,N_3293);
nor U3481 (N_3481,N_3304,N_3331);
and U3482 (N_3482,N_3330,N_3335);
xor U3483 (N_3483,N_3343,N_3295);
xnor U3484 (N_3484,N_3306,N_3294);
nand U3485 (N_3485,N_3398,N_3359);
xor U3486 (N_3486,N_3384,N_3225);
and U3487 (N_3487,N_3300,N_3366);
or U3488 (N_3488,N_3208,N_3228);
nand U3489 (N_3489,N_3364,N_3203);
and U3490 (N_3490,N_3249,N_3390);
nand U3491 (N_3491,N_3313,N_3348);
and U3492 (N_3492,N_3226,N_3255);
nand U3493 (N_3493,N_3347,N_3205);
xnor U3494 (N_3494,N_3202,N_3264);
nor U3495 (N_3495,N_3322,N_3397);
nand U3496 (N_3496,N_3261,N_3338);
or U3497 (N_3497,N_3308,N_3209);
xor U3498 (N_3498,N_3391,N_3345);
nor U3499 (N_3499,N_3302,N_3301);
nor U3500 (N_3500,N_3311,N_3208);
and U3501 (N_3501,N_3214,N_3288);
and U3502 (N_3502,N_3382,N_3290);
and U3503 (N_3503,N_3327,N_3333);
xnor U3504 (N_3504,N_3253,N_3348);
xor U3505 (N_3505,N_3280,N_3286);
nand U3506 (N_3506,N_3302,N_3278);
or U3507 (N_3507,N_3262,N_3361);
or U3508 (N_3508,N_3399,N_3344);
xor U3509 (N_3509,N_3202,N_3351);
nor U3510 (N_3510,N_3375,N_3395);
or U3511 (N_3511,N_3218,N_3306);
nand U3512 (N_3512,N_3288,N_3326);
and U3513 (N_3513,N_3217,N_3278);
and U3514 (N_3514,N_3236,N_3219);
xor U3515 (N_3515,N_3221,N_3243);
nor U3516 (N_3516,N_3331,N_3276);
xor U3517 (N_3517,N_3380,N_3227);
nor U3518 (N_3518,N_3249,N_3200);
and U3519 (N_3519,N_3325,N_3361);
nor U3520 (N_3520,N_3264,N_3208);
xnor U3521 (N_3521,N_3390,N_3317);
nand U3522 (N_3522,N_3275,N_3230);
or U3523 (N_3523,N_3291,N_3386);
or U3524 (N_3524,N_3353,N_3387);
or U3525 (N_3525,N_3364,N_3283);
and U3526 (N_3526,N_3297,N_3353);
nor U3527 (N_3527,N_3393,N_3309);
or U3528 (N_3528,N_3286,N_3311);
or U3529 (N_3529,N_3298,N_3297);
xor U3530 (N_3530,N_3276,N_3348);
nor U3531 (N_3531,N_3258,N_3215);
xor U3532 (N_3532,N_3383,N_3256);
and U3533 (N_3533,N_3268,N_3301);
and U3534 (N_3534,N_3241,N_3319);
nand U3535 (N_3535,N_3293,N_3281);
or U3536 (N_3536,N_3248,N_3272);
xnor U3537 (N_3537,N_3388,N_3380);
nand U3538 (N_3538,N_3307,N_3235);
and U3539 (N_3539,N_3290,N_3309);
and U3540 (N_3540,N_3260,N_3267);
or U3541 (N_3541,N_3273,N_3345);
xor U3542 (N_3542,N_3276,N_3233);
or U3543 (N_3543,N_3217,N_3227);
and U3544 (N_3544,N_3399,N_3330);
or U3545 (N_3545,N_3290,N_3317);
and U3546 (N_3546,N_3206,N_3346);
or U3547 (N_3547,N_3350,N_3351);
nand U3548 (N_3548,N_3323,N_3386);
xnor U3549 (N_3549,N_3308,N_3379);
nand U3550 (N_3550,N_3322,N_3373);
and U3551 (N_3551,N_3384,N_3243);
and U3552 (N_3552,N_3301,N_3295);
or U3553 (N_3553,N_3271,N_3328);
nor U3554 (N_3554,N_3335,N_3286);
nor U3555 (N_3555,N_3313,N_3269);
or U3556 (N_3556,N_3254,N_3349);
nor U3557 (N_3557,N_3302,N_3359);
and U3558 (N_3558,N_3332,N_3356);
xor U3559 (N_3559,N_3245,N_3297);
nor U3560 (N_3560,N_3230,N_3204);
and U3561 (N_3561,N_3241,N_3269);
nand U3562 (N_3562,N_3369,N_3200);
nand U3563 (N_3563,N_3399,N_3294);
or U3564 (N_3564,N_3326,N_3305);
and U3565 (N_3565,N_3234,N_3273);
or U3566 (N_3566,N_3274,N_3280);
nor U3567 (N_3567,N_3383,N_3313);
xor U3568 (N_3568,N_3392,N_3373);
nand U3569 (N_3569,N_3337,N_3218);
nor U3570 (N_3570,N_3245,N_3280);
nand U3571 (N_3571,N_3380,N_3394);
nand U3572 (N_3572,N_3248,N_3315);
or U3573 (N_3573,N_3268,N_3261);
or U3574 (N_3574,N_3373,N_3311);
nor U3575 (N_3575,N_3373,N_3210);
and U3576 (N_3576,N_3245,N_3391);
nor U3577 (N_3577,N_3352,N_3232);
or U3578 (N_3578,N_3310,N_3283);
nor U3579 (N_3579,N_3398,N_3352);
and U3580 (N_3580,N_3252,N_3328);
nor U3581 (N_3581,N_3220,N_3244);
and U3582 (N_3582,N_3330,N_3253);
and U3583 (N_3583,N_3327,N_3381);
nand U3584 (N_3584,N_3245,N_3266);
nand U3585 (N_3585,N_3393,N_3265);
nand U3586 (N_3586,N_3213,N_3361);
nor U3587 (N_3587,N_3267,N_3207);
nand U3588 (N_3588,N_3348,N_3237);
xor U3589 (N_3589,N_3371,N_3252);
nand U3590 (N_3590,N_3253,N_3247);
nand U3591 (N_3591,N_3266,N_3258);
or U3592 (N_3592,N_3363,N_3235);
and U3593 (N_3593,N_3354,N_3207);
nor U3594 (N_3594,N_3287,N_3395);
or U3595 (N_3595,N_3261,N_3310);
nor U3596 (N_3596,N_3307,N_3327);
xor U3597 (N_3597,N_3295,N_3390);
and U3598 (N_3598,N_3283,N_3387);
and U3599 (N_3599,N_3384,N_3230);
xnor U3600 (N_3600,N_3545,N_3405);
or U3601 (N_3601,N_3417,N_3404);
nor U3602 (N_3602,N_3485,N_3549);
nand U3603 (N_3603,N_3423,N_3563);
or U3604 (N_3604,N_3578,N_3587);
nor U3605 (N_3605,N_3512,N_3418);
nand U3606 (N_3606,N_3480,N_3593);
or U3607 (N_3607,N_3531,N_3498);
or U3608 (N_3608,N_3516,N_3449);
nor U3609 (N_3609,N_3580,N_3497);
nor U3610 (N_3610,N_3412,N_3536);
nor U3611 (N_3611,N_3478,N_3453);
xor U3612 (N_3612,N_3503,N_3567);
xor U3613 (N_3613,N_3594,N_3413);
and U3614 (N_3614,N_3486,N_3442);
and U3615 (N_3615,N_3586,N_3592);
and U3616 (N_3616,N_3505,N_3466);
nor U3617 (N_3617,N_3517,N_3556);
and U3618 (N_3618,N_3583,N_3523);
nand U3619 (N_3619,N_3427,N_3542);
xor U3620 (N_3620,N_3425,N_3566);
or U3621 (N_3621,N_3464,N_3455);
or U3622 (N_3622,N_3491,N_3483);
or U3623 (N_3623,N_3471,N_3515);
or U3624 (N_3624,N_3598,N_3557);
nor U3625 (N_3625,N_3450,N_3513);
nor U3626 (N_3626,N_3481,N_3408);
nor U3627 (N_3627,N_3579,N_3514);
and U3628 (N_3628,N_3562,N_3508);
or U3629 (N_3629,N_3543,N_3554);
nor U3630 (N_3630,N_3452,N_3465);
nor U3631 (N_3631,N_3477,N_3470);
xnor U3632 (N_3632,N_3475,N_3506);
or U3633 (N_3633,N_3597,N_3538);
or U3634 (N_3634,N_3570,N_3469);
or U3635 (N_3635,N_3502,N_3422);
or U3636 (N_3636,N_3415,N_3457);
or U3637 (N_3637,N_3495,N_3473);
xor U3638 (N_3638,N_3432,N_3552);
xnor U3639 (N_3639,N_3537,N_3489);
nor U3640 (N_3640,N_3401,N_3458);
and U3641 (N_3641,N_3454,N_3595);
or U3642 (N_3642,N_3484,N_3421);
or U3643 (N_3643,N_3496,N_3407);
or U3644 (N_3644,N_3448,N_3520);
nor U3645 (N_3645,N_3510,N_3400);
nor U3646 (N_3646,N_3574,N_3546);
or U3647 (N_3647,N_3482,N_3555);
nand U3648 (N_3648,N_3560,N_3461);
nand U3649 (N_3649,N_3456,N_3569);
nand U3650 (N_3650,N_3532,N_3559);
nand U3651 (N_3651,N_3582,N_3527);
nor U3652 (N_3652,N_3476,N_3534);
nor U3653 (N_3653,N_3500,N_3444);
or U3654 (N_3654,N_3447,N_3540);
nor U3655 (N_3655,N_3460,N_3521);
xor U3656 (N_3656,N_3535,N_3433);
or U3657 (N_3657,N_3487,N_3430);
nor U3658 (N_3658,N_3522,N_3507);
nand U3659 (N_3659,N_3509,N_3591);
and U3660 (N_3660,N_3564,N_3596);
and U3661 (N_3661,N_3424,N_3519);
xor U3662 (N_3662,N_3494,N_3434);
nand U3663 (N_3663,N_3436,N_3524);
nand U3664 (N_3664,N_3446,N_3588);
nor U3665 (N_3665,N_3467,N_3565);
xnor U3666 (N_3666,N_3548,N_3416);
or U3667 (N_3667,N_3439,N_3402);
nand U3668 (N_3668,N_3550,N_3581);
xnor U3669 (N_3669,N_3419,N_3590);
nand U3670 (N_3670,N_3530,N_3437);
nand U3671 (N_3671,N_3406,N_3428);
nand U3672 (N_3672,N_3493,N_3529);
and U3673 (N_3673,N_3445,N_3585);
xor U3674 (N_3674,N_3575,N_3572);
or U3675 (N_3675,N_3504,N_3438);
and U3676 (N_3676,N_3490,N_3440);
nor U3677 (N_3677,N_3553,N_3468);
nor U3678 (N_3678,N_3589,N_3492);
and U3679 (N_3679,N_3435,N_3429);
xnor U3680 (N_3680,N_3431,N_3474);
or U3681 (N_3681,N_3568,N_3414);
nor U3682 (N_3682,N_3526,N_3451);
nand U3683 (N_3683,N_3463,N_3561);
nand U3684 (N_3684,N_3472,N_3441);
xnor U3685 (N_3685,N_3459,N_3544);
xnor U3686 (N_3686,N_3584,N_3499);
and U3687 (N_3687,N_3533,N_3511);
and U3688 (N_3688,N_3571,N_3539);
nor U3689 (N_3689,N_3410,N_3599);
or U3690 (N_3690,N_3479,N_3551);
nand U3691 (N_3691,N_3577,N_3518);
or U3692 (N_3692,N_3576,N_3443);
xnor U3693 (N_3693,N_3573,N_3525);
nand U3694 (N_3694,N_3411,N_3528);
and U3695 (N_3695,N_3462,N_3558);
xnor U3696 (N_3696,N_3409,N_3403);
or U3697 (N_3697,N_3501,N_3541);
or U3698 (N_3698,N_3426,N_3420);
nor U3699 (N_3699,N_3547,N_3488);
xor U3700 (N_3700,N_3440,N_3473);
nand U3701 (N_3701,N_3472,N_3574);
nand U3702 (N_3702,N_3459,N_3539);
or U3703 (N_3703,N_3581,N_3433);
and U3704 (N_3704,N_3424,N_3440);
nor U3705 (N_3705,N_3547,N_3574);
or U3706 (N_3706,N_3484,N_3518);
nor U3707 (N_3707,N_3586,N_3405);
xnor U3708 (N_3708,N_3492,N_3531);
or U3709 (N_3709,N_3546,N_3488);
and U3710 (N_3710,N_3582,N_3420);
and U3711 (N_3711,N_3585,N_3598);
and U3712 (N_3712,N_3544,N_3505);
and U3713 (N_3713,N_3504,N_3511);
and U3714 (N_3714,N_3589,N_3524);
nand U3715 (N_3715,N_3460,N_3491);
nor U3716 (N_3716,N_3557,N_3532);
xnor U3717 (N_3717,N_3516,N_3470);
nor U3718 (N_3718,N_3597,N_3580);
or U3719 (N_3719,N_3581,N_3597);
nand U3720 (N_3720,N_3491,N_3552);
nand U3721 (N_3721,N_3466,N_3433);
nor U3722 (N_3722,N_3409,N_3404);
xor U3723 (N_3723,N_3567,N_3526);
and U3724 (N_3724,N_3547,N_3483);
or U3725 (N_3725,N_3581,N_3405);
xnor U3726 (N_3726,N_3571,N_3562);
xor U3727 (N_3727,N_3533,N_3571);
xnor U3728 (N_3728,N_3402,N_3430);
or U3729 (N_3729,N_3587,N_3495);
nor U3730 (N_3730,N_3511,N_3578);
xnor U3731 (N_3731,N_3497,N_3599);
xnor U3732 (N_3732,N_3465,N_3460);
nor U3733 (N_3733,N_3462,N_3406);
or U3734 (N_3734,N_3535,N_3482);
nand U3735 (N_3735,N_3558,N_3592);
nor U3736 (N_3736,N_3416,N_3428);
nor U3737 (N_3737,N_3575,N_3497);
or U3738 (N_3738,N_3596,N_3490);
xnor U3739 (N_3739,N_3547,N_3451);
nor U3740 (N_3740,N_3461,N_3533);
xnor U3741 (N_3741,N_3543,N_3540);
nor U3742 (N_3742,N_3558,N_3532);
nor U3743 (N_3743,N_3526,N_3571);
xnor U3744 (N_3744,N_3430,N_3489);
nor U3745 (N_3745,N_3544,N_3575);
xnor U3746 (N_3746,N_3503,N_3406);
or U3747 (N_3747,N_3582,N_3442);
nand U3748 (N_3748,N_3539,N_3496);
nor U3749 (N_3749,N_3559,N_3482);
or U3750 (N_3750,N_3457,N_3475);
xor U3751 (N_3751,N_3463,N_3442);
or U3752 (N_3752,N_3548,N_3493);
and U3753 (N_3753,N_3504,N_3456);
or U3754 (N_3754,N_3551,N_3506);
and U3755 (N_3755,N_3530,N_3500);
and U3756 (N_3756,N_3567,N_3420);
nor U3757 (N_3757,N_3455,N_3461);
nor U3758 (N_3758,N_3417,N_3454);
xnor U3759 (N_3759,N_3506,N_3441);
xnor U3760 (N_3760,N_3599,N_3577);
nand U3761 (N_3761,N_3578,N_3499);
xor U3762 (N_3762,N_3454,N_3458);
or U3763 (N_3763,N_3586,N_3477);
nor U3764 (N_3764,N_3563,N_3564);
nor U3765 (N_3765,N_3455,N_3457);
nor U3766 (N_3766,N_3497,N_3436);
nor U3767 (N_3767,N_3479,N_3468);
xor U3768 (N_3768,N_3574,N_3414);
nand U3769 (N_3769,N_3584,N_3444);
xnor U3770 (N_3770,N_3456,N_3453);
xor U3771 (N_3771,N_3542,N_3488);
and U3772 (N_3772,N_3416,N_3475);
xor U3773 (N_3773,N_3518,N_3439);
or U3774 (N_3774,N_3403,N_3584);
or U3775 (N_3775,N_3404,N_3420);
nor U3776 (N_3776,N_3565,N_3459);
xnor U3777 (N_3777,N_3570,N_3531);
nand U3778 (N_3778,N_3406,N_3533);
xnor U3779 (N_3779,N_3471,N_3407);
or U3780 (N_3780,N_3500,N_3546);
or U3781 (N_3781,N_3435,N_3567);
or U3782 (N_3782,N_3552,N_3480);
nor U3783 (N_3783,N_3461,N_3586);
nand U3784 (N_3784,N_3426,N_3409);
xnor U3785 (N_3785,N_3594,N_3426);
nor U3786 (N_3786,N_3557,N_3519);
and U3787 (N_3787,N_3594,N_3488);
and U3788 (N_3788,N_3446,N_3547);
or U3789 (N_3789,N_3466,N_3554);
xor U3790 (N_3790,N_3497,N_3587);
nor U3791 (N_3791,N_3453,N_3477);
or U3792 (N_3792,N_3537,N_3405);
nand U3793 (N_3793,N_3429,N_3458);
and U3794 (N_3794,N_3473,N_3461);
xor U3795 (N_3795,N_3513,N_3519);
and U3796 (N_3796,N_3405,N_3505);
or U3797 (N_3797,N_3460,N_3446);
xor U3798 (N_3798,N_3445,N_3449);
nand U3799 (N_3799,N_3535,N_3562);
or U3800 (N_3800,N_3626,N_3791);
nand U3801 (N_3801,N_3761,N_3618);
nand U3802 (N_3802,N_3723,N_3682);
and U3803 (N_3803,N_3779,N_3754);
and U3804 (N_3804,N_3632,N_3649);
or U3805 (N_3805,N_3681,N_3660);
nor U3806 (N_3806,N_3733,N_3620);
nor U3807 (N_3807,N_3750,N_3781);
nor U3808 (N_3808,N_3794,N_3748);
or U3809 (N_3809,N_3651,N_3668);
or U3810 (N_3810,N_3696,N_3767);
xor U3811 (N_3811,N_3621,N_3743);
xnor U3812 (N_3812,N_3629,N_3677);
xnor U3813 (N_3813,N_3770,N_3640);
nor U3814 (N_3814,N_3695,N_3790);
xnor U3815 (N_3815,N_3675,N_3687);
or U3816 (N_3816,N_3663,N_3730);
nor U3817 (N_3817,N_3707,N_3753);
and U3818 (N_3818,N_3751,N_3669);
and U3819 (N_3819,N_3613,N_3670);
xnor U3820 (N_3820,N_3732,N_3785);
nor U3821 (N_3821,N_3659,N_3686);
and U3822 (N_3822,N_3740,N_3777);
xnor U3823 (N_3823,N_3728,N_3658);
xnor U3824 (N_3824,N_3611,N_3724);
xor U3825 (N_3825,N_3721,N_3617);
and U3826 (N_3826,N_3711,N_3671);
nor U3827 (N_3827,N_3657,N_3600);
nand U3828 (N_3828,N_3757,N_3624);
nor U3829 (N_3829,N_3709,N_3776);
xnor U3830 (N_3830,N_3644,N_3713);
xor U3831 (N_3831,N_3765,N_3688);
and U3832 (N_3832,N_3666,N_3604);
nand U3833 (N_3833,N_3633,N_3737);
or U3834 (N_3834,N_3698,N_3716);
nor U3835 (N_3835,N_3678,N_3714);
and U3836 (N_3836,N_3648,N_3741);
or U3837 (N_3837,N_3672,N_3742);
xor U3838 (N_3838,N_3771,N_3784);
nand U3839 (N_3839,N_3758,N_3631);
or U3840 (N_3840,N_3639,N_3614);
nand U3841 (N_3841,N_3705,N_3609);
and U3842 (N_3842,N_3645,N_3769);
xnor U3843 (N_3843,N_3685,N_3755);
nor U3844 (N_3844,N_3684,N_3792);
and U3845 (N_3845,N_3789,N_3607);
or U3846 (N_3846,N_3637,N_3622);
and U3847 (N_3847,N_3653,N_3702);
or U3848 (N_3848,N_3704,N_3766);
and U3849 (N_3849,N_3768,N_3634);
and U3850 (N_3850,N_3662,N_3756);
nor U3851 (N_3851,N_3787,N_3606);
xor U3852 (N_3852,N_3774,N_3615);
nor U3853 (N_3853,N_3654,N_3734);
nand U3854 (N_3854,N_3693,N_3652);
and U3855 (N_3855,N_3661,N_3778);
and U3856 (N_3856,N_3788,N_3628);
and U3857 (N_3857,N_3601,N_3674);
and U3858 (N_3858,N_3673,N_3627);
nor U3859 (N_3859,N_3676,N_3783);
nor U3860 (N_3860,N_3638,N_3616);
or U3861 (N_3861,N_3797,N_3694);
nand U3862 (N_3862,N_3646,N_3643);
nand U3863 (N_3863,N_3736,N_3665);
or U3864 (N_3864,N_3725,N_3719);
nor U3865 (N_3865,N_3796,N_3680);
or U3866 (N_3866,N_3772,N_3717);
nor U3867 (N_3867,N_3602,N_3689);
nor U3868 (N_3868,N_3720,N_3799);
nand U3869 (N_3869,N_3735,N_3739);
and U3870 (N_3870,N_3744,N_3712);
and U3871 (N_3871,N_3726,N_3738);
or U3872 (N_3872,N_3610,N_3773);
nor U3873 (N_3873,N_3780,N_3745);
and U3874 (N_3874,N_3752,N_3715);
or U3875 (N_3875,N_3706,N_3786);
nor U3876 (N_3876,N_3650,N_3729);
or U3877 (N_3877,N_3703,N_3641);
or U3878 (N_3878,N_3605,N_3718);
and U3879 (N_3879,N_3731,N_3608);
xnor U3880 (N_3880,N_3763,N_3795);
or U3881 (N_3881,N_3722,N_3775);
nand U3882 (N_3882,N_3667,N_3699);
nor U3883 (N_3883,N_3762,N_3746);
or U3884 (N_3884,N_3625,N_3690);
nor U3885 (N_3885,N_3691,N_3727);
nor U3886 (N_3886,N_3679,N_3697);
nand U3887 (N_3887,N_3636,N_3710);
nand U3888 (N_3888,N_3683,N_3623);
and U3889 (N_3889,N_3647,N_3619);
nand U3890 (N_3890,N_3798,N_3612);
nor U3891 (N_3891,N_3635,N_3747);
and U3892 (N_3892,N_3759,N_3782);
and U3893 (N_3893,N_3664,N_3630);
or U3894 (N_3894,N_3760,N_3700);
or U3895 (N_3895,N_3642,N_3708);
nand U3896 (N_3896,N_3655,N_3701);
nor U3897 (N_3897,N_3692,N_3793);
nand U3898 (N_3898,N_3603,N_3764);
or U3899 (N_3899,N_3749,N_3656);
or U3900 (N_3900,N_3768,N_3644);
nor U3901 (N_3901,N_3746,N_3742);
and U3902 (N_3902,N_3692,N_3736);
nor U3903 (N_3903,N_3789,N_3780);
nand U3904 (N_3904,N_3652,N_3642);
nor U3905 (N_3905,N_3773,N_3727);
or U3906 (N_3906,N_3621,N_3619);
or U3907 (N_3907,N_3766,N_3792);
or U3908 (N_3908,N_3630,N_3724);
xor U3909 (N_3909,N_3738,N_3788);
and U3910 (N_3910,N_3600,N_3746);
and U3911 (N_3911,N_3767,N_3625);
nor U3912 (N_3912,N_3733,N_3674);
nor U3913 (N_3913,N_3734,N_3698);
nor U3914 (N_3914,N_3787,N_3639);
and U3915 (N_3915,N_3652,N_3623);
nand U3916 (N_3916,N_3628,N_3786);
nor U3917 (N_3917,N_3618,N_3790);
and U3918 (N_3918,N_3615,N_3607);
and U3919 (N_3919,N_3610,N_3626);
nand U3920 (N_3920,N_3790,N_3699);
or U3921 (N_3921,N_3713,N_3732);
nand U3922 (N_3922,N_3682,N_3654);
or U3923 (N_3923,N_3762,N_3709);
xnor U3924 (N_3924,N_3770,N_3745);
nand U3925 (N_3925,N_3671,N_3693);
and U3926 (N_3926,N_3660,N_3785);
nand U3927 (N_3927,N_3713,N_3617);
or U3928 (N_3928,N_3762,N_3683);
or U3929 (N_3929,N_3603,N_3691);
and U3930 (N_3930,N_3787,N_3712);
nand U3931 (N_3931,N_3787,N_3630);
and U3932 (N_3932,N_3798,N_3791);
xnor U3933 (N_3933,N_3607,N_3791);
nand U3934 (N_3934,N_3624,N_3616);
nor U3935 (N_3935,N_3770,N_3606);
and U3936 (N_3936,N_3732,N_3639);
and U3937 (N_3937,N_3662,N_3629);
xnor U3938 (N_3938,N_3608,N_3733);
nor U3939 (N_3939,N_3706,N_3655);
xnor U3940 (N_3940,N_3735,N_3681);
and U3941 (N_3941,N_3645,N_3636);
xor U3942 (N_3942,N_3662,N_3762);
xor U3943 (N_3943,N_3671,N_3718);
or U3944 (N_3944,N_3615,N_3701);
or U3945 (N_3945,N_3769,N_3615);
nand U3946 (N_3946,N_3705,N_3749);
nor U3947 (N_3947,N_3606,N_3605);
and U3948 (N_3948,N_3735,N_3683);
xnor U3949 (N_3949,N_3771,N_3692);
xnor U3950 (N_3950,N_3643,N_3776);
xnor U3951 (N_3951,N_3786,N_3775);
and U3952 (N_3952,N_3663,N_3685);
or U3953 (N_3953,N_3689,N_3745);
nand U3954 (N_3954,N_3775,N_3616);
or U3955 (N_3955,N_3746,N_3633);
nor U3956 (N_3956,N_3678,N_3780);
or U3957 (N_3957,N_3606,N_3630);
xor U3958 (N_3958,N_3657,N_3662);
and U3959 (N_3959,N_3707,N_3756);
xor U3960 (N_3960,N_3677,N_3676);
xnor U3961 (N_3961,N_3675,N_3752);
or U3962 (N_3962,N_3636,N_3772);
and U3963 (N_3963,N_3703,N_3732);
and U3964 (N_3964,N_3695,N_3674);
and U3965 (N_3965,N_3775,N_3789);
nor U3966 (N_3966,N_3725,N_3702);
or U3967 (N_3967,N_3688,N_3707);
nor U3968 (N_3968,N_3795,N_3746);
or U3969 (N_3969,N_3665,N_3637);
nor U3970 (N_3970,N_3658,N_3737);
nor U3971 (N_3971,N_3761,N_3620);
nand U3972 (N_3972,N_3702,N_3797);
xor U3973 (N_3973,N_3700,N_3711);
nand U3974 (N_3974,N_3667,N_3663);
and U3975 (N_3975,N_3750,N_3714);
nor U3976 (N_3976,N_3696,N_3643);
xnor U3977 (N_3977,N_3795,N_3718);
nand U3978 (N_3978,N_3648,N_3785);
nand U3979 (N_3979,N_3768,N_3602);
or U3980 (N_3980,N_3767,N_3769);
nand U3981 (N_3981,N_3636,N_3655);
nor U3982 (N_3982,N_3737,N_3743);
and U3983 (N_3983,N_3784,N_3672);
xor U3984 (N_3984,N_3693,N_3724);
nand U3985 (N_3985,N_3628,N_3785);
and U3986 (N_3986,N_3654,N_3628);
and U3987 (N_3987,N_3644,N_3682);
nor U3988 (N_3988,N_3673,N_3632);
xor U3989 (N_3989,N_3654,N_3659);
or U3990 (N_3990,N_3708,N_3656);
or U3991 (N_3991,N_3619,N_3689);
nor U3992 (N_3992,N_3747,N_3724);
nand U3993 (N_3993,N_3794,N_3734);
or U3994 (N_3994,N_3779,N_3677);
nand U3995 (N_3995,N_3758,N_3778);
xor U3996 (N_3996,N_3675,N_3712);
nor U3997 (N_3997,N_3720,N_3614);
and U3998 (N_3998,N_3662,N_3717);
and U3999 (N_3999,N_3744,N_3655);
and U4000 (N_4000,N_3838,N_3867);
nor U4001 (N_4001,N_3994,N_3857);
xnor U4002 (N_4002,N_3810,N_3985);
xnor U4003 (N_4003,N_3832,N_3960);
xnor U4004 (N_4004,N_3885,N_3828);
and U4005 (N_4005,N_3860,N_3854);
or U4006 (N_4006,N_3874,N_3822);
nor U4007 (N_4007,N_3817,N_3925);
or U4008 (N_4008,N_3927,N_3870);
or U4009 (N_4009,N_3891,N_3981);
or U4010 (N_4010,N_3820,N_3932);
and U4011 (N_4011,N_3955,N_3949);
or U4012 (N_4012,N_3951,N_3993);
or U4013 (N_4013,N_3824,N_3956);
nor U4014 (N_4014,N_3992,N_3914);
nor U4015 (N_4015,N_3851,N_3945);
and U4016 (N_4016,N_3829,N_3868);
xnor U4017 (N_4017,N_3903,N_3908);
xnor U4018 (N_4018,N_3998,N_3937);
nand U4019 (N_4019,N_3827,N_3971);
xnor U4020 (N_4020,N_3977,N_3912);
nor U4021 (N_4021,N_3896,N_3946);
and U4022 (N_4022,N_3865,N_3926);
nor U4023 (N_4023,N_3941,N_3880);
and U4024 (N_4024,N_3808,N_3899);
nand U4025 (N_4025,N_3906,N_3879);
nor U4026 (N_4026,N_3889,N_3848);
xnor U4027 (N_4027,N_3934,N_3833);
or U4028 (N_4028,N_3920,N_3904);
xnor U4029 (N_4029,N_3964,N_3815);
and U4030 (N_4030,N_3866,N_3967);
and U4031 (N_4031,N_3959,N_3845);
nor U4032 (N_4032,N_3890,N_3961);
xor U4033 (N_4033,N_3907,N_3846);
or U4034 (N_4034,N_3929,N_3893);
nor U4035 (N_4035,N_3864,N_3913);
xor U4036 (N_4036,N_3826,N_3861);
nand U4037 (N_4037,N_3917,N_3969);
and U4038 (N_4038,N_3915,N_3999);
and U4039 (N_4039,N_3919,N_3805);
xnor U4040 (N_4040,N_3898,N_3947);
or U4041 (N_4041,N_3989,N_3843);
and U4042 (N_4042,N_3834,N_3821);
nor U4043 (N_4043,N_3886,N_3931);
or U4044 (N_4044,N_3948,N_3982);
xor U4045 (N_4045,N_3935,N_3952);
nand U4046 (N_4046,N_3863,N_3922);
or U4047 (N_4047,N_3975,N_3943);
or U4048 (N_4048,N_3856,N_3997);
nor U4049 (N_4049,N_3847,N_3958);
nor U4050 (N_4050,N_3849,N_3963);
and U4051 (N_4051,N_3850,N_3840);
xnor U4052 (N_4052,N_3962,N_3816);
nand U4053 (N_4053,N_3819,N_3910);
xnor U4054 (N_4054,N_3804,N_3823);
xnor U4055 (N_4055,N_3965,N_3825);
nand U4056 (N_4056,N_3916,N_3811);
nor U4057 (N_4057,N_3901,N_3921);
xnor U4058 (N_4058,N_3887,N_3897);
nor U4059 (N_4059,N_3980,N_3803);
nand U4060 (N_4060,N_3974,N_3942);
and U4061 (N_4061,N_3875,N_3938);
xnor U4062 (N_4062,N_3983,N_3814);
nand U4063 (N_4063,N_3950,N_3930);
xor U4064 (N_4064,N_3968,N_3895);
xnor U4065 (N_4065,N_3883,N_3924);
xor U4066 (N_4066,N_3806,N_3873);
and U4067 (N_4067,N_3972,N_3877);
nor U4068 (N_4068,N_3995,N_3988);
nor U4069 (N_4069,N_3839,N_3918);
nor U4070 (N_4070,N_3812,N_3978);
and U4071 (N_4071,N_3872,N_3830);
and U4072 (N_4072,N_3836,N_3973);
and U4073 (N_4073,N_3888,N_3855);
xor U4074 (N_4074,N_3841,N_3801);
nand U4075 (N_4075,N_3986,N_3996);
nor U4076 (N_4076,N_3953,N_3987);
nand U4077 (N_4077,N_3944,N_3807);
or U4078 (N_4078,N_3842,N_3818);
xnor U4079 (N_4079,N_3882,N_3979);
and U4080 (N_4080,N_3869,N_3976);
and U4081 (N_4081,N_3902,N_3923);
nand U4082 (N_4082,N_3957,N_3862);
nand U4083 (N_4083,N_3911,N_3892);
nand U4084 (N_4084,N_3970,N_3966);
nor U4085 (N_4085,N_3991,N_3858);
xor U4086 (N_4086,N_3894,N_3852);
nor U4087 (N_4087,N_3831,N_3876);
nor U4088 (N_4088,N_3909,N_3940);
nor U4089 (N_4089,N_3853,N_3954);
nand U4090 (N_4090,N_3933,N_3900);
and U4091 (N_4091,N_3939,N_3928);
and U4092 (N_4092,N_3878,N_3881);
and U4093 (N_4093,N_3859,N_3905);
xnor U4094 (N_4094,N_3800,N_3936);
nor U4095 (N_4095,N_3809,N_3813);
nand U4096 (N_4096,N_3871,N_3884);
xor U4097 (N_4097,N_3802,N_3837);
nand U4098 (N_4098,N_3835,N_3990);
xor U4099 (N_4099,N_3844,N_3984);
and U4100 (N_4100,N_3874,N_3980);
nor U4101 (N_4101,N_3815,N_3923);
xor U4102 (N_4102,N_3836,N_3940);
or U4103 (N_4103,N_3858,N_3897);
nor U4104 (N_4104,N_3824,N_3859);
nand U4105 (N_4105,N_3958,N_3810);
nand U4106 (N_4106,N_3944,N_3952);
nor U4107 (N_4107,N_3904,N_3983);
nand U4108 (N_4108,N_3957,N_3892);
nor U4109 (N_4109,N_3854,N_3889);
xor U4110 (N_4110,N_3878,N_3984);
and U4111 (N_4111,N_3870,N_3965);
nand U4112 (N_4112,N_3861,N_3911);
and U4113 (N_4113,N_3870,N_3864);
xnor U4114 (N_4114,N_3868,N_3878);
and U4115 (N_4115,N_3991,N_3888);
or U4116 (N_4116,N_3857,N_3821);
nand U4117 (N_4117,N_3876,N_3951);
nor U4118 (N_4118,N_3907,N_3893);
nand U4119 (N_4119,N_3883,N_3935);
and U4120 (N_4120,N_3918,N_3826);
nor U4121 (N_4121,N_3801,N_3833);
xnor U4122 (N_4122,N_3810,N_3868);
and U4123 (N_4123,N_3989,N_3849);
nor U4124 (N_4124,N_3827,N_3964);
nand U4125 (N_4125,N_3829,N_3865);
nand U4126 (N_4126,N_3856,N_3893);
xor U4127 (N_4127,N_3853,N_3977);
xnor U4128 (N_4128,N_3919,N_3836);
nand U4129 (N_4129,N_3981,N_3949);
nor U4130 (N_4130,N_3985,N_3881);
xor U4131 (N_4131,N_3896,N_3957);
or U4132 (N_4132,N_3953,N_3940);
nand U4133 (N_4133,N_3824,N_3862);
or U4134 (N_4134,N_3997,N_3927);
and U4135 (N_4135,N_3802,N_3990);
nor U4136 (N_4136,N_3821,N_3848);
and U4137 (N_4137,N_3980,N_3832);
xnor U4138 (N_4138,N_3900,N_3881);
and U4139 (N_4139,N_3843,N_3835);
nor U4140 (N_4140,N_3861,N_3851);
or U4141 (N_4141,N_3914,N_3804);
or U4142 (N_4142,N_3933,N_3981);
and U4143 (N_4143,N_3936,N_3889);
nand U4144 (N_4144,N_3868,N_3834);
or U4145 (N_4145,N_3847,N_3857);
xor U4146 (N_4146,N_3932,N_3892);
nor U4147 (N_4147,N_3964,N_3844);
and U4148 (N_4148,N_3812,N_3842);
nand U4149 (N_4149,N_3995,N_3817);
nand U4150 (N_4150,N_3833,N_3992);
and U4151 (N_4151,N_3905,N_3805);
and U4152 (N_4152,N_3930,N_3887);
xnor U4153 (N_4153,N_3845,N_3971);
or U4154 (N_4154,N_3877,N_3916);
nor U4155 (N_4155,N_3916,N_3860);
xnor U4156 (N_4156,N_3885,N_3962);
nor U4157 (N_4157,N_3995,N_3933);
nor U4158 (N_4158,N_3871,N_3840);
and U4159 (N_4159,N_3912,N_3807);
nor U4160 (N_4160,N_3909,N_3999);
or U4161 (N_4161,N_3888,N_3914);
or U4162 (N_4162,N_3889,N_3964);
nand U4163 (N_4163,N_3849,N_3871);
nand U4164 (N_4164,N_3827,N_3984);
nand U4165 (N_4165,N_3842,N_3836);
nand U4166 (N_4166,N_3989,N_3983);
xor U4167 (N_4167,N_3876,N_3802);
nor U4168 (N_4168,N_3981,N_3877);
xnor U4169 (N_4169,N_3854,N_3989);
or U4170 (N_4170,N_3921,N_3900);
nand U4171 (N_4171,N_3814,N_3987);
nand U4172 (N_4172,N_3827,N_3802);
nand U4173 (N_4173,N_3957,N_3979);
or U4174 (N_4174,N_3939,N_3835);
and U4175 (N_4175,N_3860,N_3892);
nand U4176 (N_4176,N_3973,N_3817);
or U4177 (N_4177,N_3910,N_3839);
xnor U4178 (N_4178,N_3931,N_3881);
nor U4179 (N_4179,N_3907,N_3820);
and U4180 (N_4180,N_3962,N_3936);
xnor U4181 (N_4181,N_3841,N_3989);
or U4182 (N_4182,N_3914,N_3882);
xor U4183 (N_4183,N_3852,N_3878);
nand U4184 (N_4184,N_3921,N_3962);
or U4185 (N_4185,N_3979,N_3836);
xor U4186 (N_4186,N_3853,N_3867);
nand U4187 (N_4187,N_3848,N_3988);
and U4188 (N_4188,N_3832,N_3867);
nand U4189 (N_4189,N_3859,N_3891);
and U4190 (N_4190,N_3880,N_3869);
and U4191 (N_4191,N_3888,N_3919);
nand U4192 (N_4192,N_3873,N_3836);
nand U4193 (N_4193,N_3872,N_3818);
nand U4194 (N_4194,N_3800,N_3964);
nor U4195 (N_4195,N_3855,N_3978);
nor U4196 (N_4196,N_3933,N_3918);
and U4197 (N_4197,N_3802,N_3902);
and U4198 (N_4198,N_3818,N_3852);
or U4199 (N_4199,N_3987,N_3960);
and U4200 (N_4200,N_4106,N_4198);
xor U4201 (N_4201,N_4001,N_4055);
nand U4202 (N_4202,N_4023,N_4130);
xnor U4203 (N_4203,N_4170,N_4167);
nor U4204 (N_4204,N_4082,N_4156);
or U4205 (N_4205,N_4073,N_4092);
xor U4206 (N_4206,N_4123,N_4184);
nor U4207 (N_4207,N_4072,N_4191);
or U4208 (N_4208,N_4060,N_4128);
nor U4209 (N_4209,N_4042,N_4044);
or U4210 (N_4210,N_4062,N_4158);
and U4211 (N_4211,N_4013,N_4047);
nand U4212 (N_4212,N_4122,N_4175);
or U4213 (N_4213,N_4083,N_4153);
nor U4214 (N_4214,N_4144,N_4081);
xnor U4215 (N_4215,N_4117,N_4077);
and U4216 (N_4216,N_4032,N_4193);
and U4217 (N_4217,N_4068,N_4096);
nand U4218 (N_4218,N_4059,N_4053);
or U4219 (N_4219,N_4026,N_4134);
xor U4220 (N_4220,N_4008,N_4034);
or U4221 (N_4221,N_4003,N_4131);
nor U4222 (N_4222,N_4155,N_4129);
and U4223 (N_4223,N_4126,N_4196);
or U4224 (N_4224,N_4190,N_4145);
nand U4225 (N_4225,N_4186,N_4015);
nand U4226 (N_4226,N_4125,N_4133);
nor U4227 (N_4227,N_4182,N_4192);
nand U4228 (N_4228,N_4140,N_4039);
or U4229 (N_4229,N_4118,N_4009);
nand U4230 (N_4230,N_4031,N_4159);
nor U4231 (N_4231,N_4037,N_4102);
or U4232 (N_4232,N_4172,N_4074);
nand U4233 (N_4233,N_4025,N_4116);
and U4234 (N_4234,N_4048,N_4107);
and U4235 (N_4235,N_4054,N_4137);
nor U4236 (N_4236,N_4188,N_4132);
xor U4237 (N_4237,N_4104,N_4151);
or U4238 (N_4238,N_4024,N_4120);
and U4239 (N_4239,N_4088,N_4010);
or U4240 (N_4240,N_4051,N_4098);
nand U4241 (N_4241,N_4127,N_4165);
nand U4242 (N_4242,N_4089,N_4057);
and U4243 (N_4243,N_4181,N_4091);
xor U4244 (N_4244,N_4064,N_4056);
and U4245 (N_4245,N_4052,N_4078);
xor U4246 (N_4246,N_4021,N_4194);
nand U4247 (N_4247,N_4119,N_4149);
or U4248 (N_4248,N_4079,N_4017);
nand U4249 (N_4249,N_4020,N_4076);
and U4250 (N_4250,N_4006,N_4195);
and U4251 (N_4251,N_4121,N_4012);
xnor U4252 (N_4252,N_4178,N_4046);
or U4253 (N_4253,N_4136,N_4018);
and U4254 (N_4254,N_4166,N_4148);
xnor U4255 (N_4255,N_4093,N_4146);
nor U4256 (N_4256,N_4169,N_4085);
or U4257 (N_4257,N_4071,N_4110);
or U4258 (N_4258,N_4069,N_4027);
xor U4259 (N_4259,N_4142,N_4029);
nand U4260 (N_4260,N_4111,N_4004);
and U4261 (N_4261,N_4011,N_4080);
nor U4262 (N_4262,N_4038,N_4138);
xor U4263 (N_4263,N_4177,N_4014);
xnor U4264 (N_4264,N_4199,N_4143);
and U4265 (N_4265,N_4152,N_4176);
and U4266 (N_4266,N_4019,N_4114);
or U4267 (N_4267,N_4000,N_4028);
and U4268 (N_4268,N_4050,N_4139);
xor U4269 (N_4269,N_4007,N_4183);
nand U4270 (N_4270,N_4150,N_4108);
or U4271 (N_4271,N_4036,N_4063);
xor U4272 (N_4272,N_4171,N_4066);
and U4273 (N_4273,N_4084,N_4109);
nand U4274 (N_4274,N_4100,N_4163);
nor U4275 (N_4275,N_4095,N_4090);
and U4276 (N_4276,N_4067,N_4035);
and U4277 (N_4277,N_4180,N_4162);
or U4278 (N_4278,N_4157,N_4168);
nor U4279 (N_4279,N_4002,N_4030);
nor U4280 (N_4280,N_4070,N_4005);
nor U4281 (N_4281,N_4179,N_4141);
xnor U4282 (N_4282,N_4147,N_4103);
and U4283 (N_4283,N_4112,N_4185);
or U4284 (N_4284,N_4061,N_4154);
nand U4285 (N_4285,N_4016,N_4187);
nand U4286 (N_4286,N_4173,N_4160);
and U4287 (N_4287,N_4101,N_4043);
or U4288 (N_4288,N_4124,N_4058);
nand U4289 (N_4289,N_4086,N_4045);
nand U4290 (N_4290,N_4135,N_4041);
xnor U4291 (N_4291,N_4065,N_4099);
or U4292 (N_4292,N_4105,N_4113);
xnor U4293 (N_4293,N_4189,N_4097);
nand U4294 (N_4294,N_4087,N_4022);
and U4295 (N_4295,N_4033,N_4174);
xnor U4296 (N_4296,N_4094,N_4161);
or U4297 (N_4297,N_4040,N_4164);
xor U4298 (N_4298,N_4049,N_4075);
xor U4299 (N_4299,N_4197,N_4115);
nand U4300 (N_4300,N_4085,N_4009);
nor U4301 (N_4301,N_4148,N_4162);
nor U4302 (N_4302,N_4182,N_4089);
and U4303 (N_4303,N_4026,N_4130);
xor U4304 (N_4304,N_4175,N_4114);
xor U4305 (N_4305,N_4038,N_4177);
and U4306 (N_4306,N_4006,N_4194);
or U4307 (N_4307,N_4166,N_4137);
or U4308 (N_4308,N_4069,N_4036);
nand U4309 (N_4309,N_4190,N_4088);
and U4310 (N_4310,N_4146,N_4124);
nor U4311 (N_4311,N_4173,N_4072);
nand U4312 (N_4312,N_4085,N_4000);
or U4313 (N_4313,N_4180,N_4157);
nor U4314 (N_4314,N_4071,N_4044);
nand U4315 (N_4315,N_4078,N_4189);
or U4316 (N_4316,N_4036,N_4060);
or U4317 (N_4317,N_4015,N_4086);
and U4318 (N_4318,N_4061,N_4051);
and U4319 (N_4319,N_4128,N_4011);
and U4320 (N_4320,N_4141,N_4010);
xor U4321 (N_4321,N_4009,N_4171);
and U4322 (N_4322,N_4169,N_4015);
and U4323 (N_4323,N_4197,N_4108);
nor U4324 (N_4324,N_4088,N_4108);
or U4325 (N_4325,N_4168,N_4059);
nor U4326 (N_4326,N_4165,N_4034);
nand U4327 (N_4327,N_4170,N_4161);
xnor U4328 (N_4328,N_4031,N_4104);
and U4329 (N_4329,N_4076,N_4008);
nand U4330 (N_4330,N_4143,N_4061);
nand U4331 (N_4331,N_4086,N_4143);
nor U4332 (N_4332,N_4180,N_4113);
or U4333 (N_4333,N_4061,N_4036);
xnor U4334 (N_4334,N_4171,N_4051);
nand U4335 (N_4335,N_4053,N_4078);
or U4336 (N_4336,N_4035,N_4119);
nand U4337 (N_4337,N_4076,N_4060);
or U4338 (N_4338,N_4055,N_4186);
or U4339 (N_4339,N_4084,N_4096);
or U4340 (N_4340,N_4149,N_4024);
and U4341 (N_4341,N_4105,N_4085);
or U4342 (N_4342,N_4137,N_4138);
and U4343 (N_4343,N_4186,N_4178);
nand U4344 (N_4344,N_4173,N_4086);
xnor U4345 (N_4345,N_4127,N_4092);
and U4346 (N_4346,N_4051,N_4000);
nand U4347 (N_4347,N_4048,N_4178);
nand U4348 (N_4348,N_4179,N_4070);
nor U4349 (N_4349,N_4123,N_4178);
or U4350 (N_4350,N_4172,N_4044);
xnor U4351 (N_4351,N_4043,N_4089);
and U4352 (N_4352,N_4100,N_4197);
xor U4353 (N_4353,N_4167,N_4135);
nand U4354 (N_4354,N_4005,N_4129);
and U4355 (N_4355,N_4194,N_4144);
and U4356 (N_4356,N_4023,N_4175);
or U4357 (N_4357,N_4024,N_4106);
and U4358 (N_4358,N_4008,N_4103);
and U4359 (N_4359,N_4168,N_4018);
nor U4360 (N_4360,N_4088,N_4030);
nor U4361 (N_4361,N_4191,N_4004);
or U4362 (N_4362,N_4147,N_4077);
nor U4363 (N_4363,N_4003,N_4018);
nor U4364 (N_4364,N_4042,N_4195);
and U4365 (N_4365,N_4035,N_4013);
nor U4366 (N_4366,N_4024,N_4008);
or U4367 (N_4367,N_4186,N_4151);
and U4368 (N_4368,N_4026,N_4058);
and U4369 (N_4369,N_4055,N_4144);
nand U4370 (N_4370,N_4003,N_4096);
or U4371 (N_4371,N_4071,N_4169);
and U4372 (N_4372,N_4079,N_4144);
xor U4373 (N_4373,N_4126,N_4102);
nor U4374 (N_4374,N_4106,N_4020);
nor U4375 (N_4375,N_4117,N_4157);
xnor U4376 (N_4376,N_4032,N_4092);
nor U4377 (N_4377,N_4183,N_4108);
and U4378 (N_4378,N_4051,N_4112);
nor U4379 (N_4379,N_4072,N_4076);
nor U4380 (N_4380,N_4037,N_4023);
xnor U4381 (N_4381,N_4035,N_4189);
nor U4382 (N_4382,N_4108,N_4035);
or U4383 (N_4383,N_4003,N_4195);
nor U4384 (N_4384,N_4072,N_4160);
and U4385 (N_4385,N_4081,N_4007);
nor U4386 (N_4386,N_4150,N_4008);
nor U4387 (N_4387,N_4064,N_4135);
xor U4388 (N_4388,N_4080,N_4111);
nor U4389 (N_4389,N_4130,N_4151);
or U4390 (N_4390,N_4133,N_4157);
xnor U4391 (N_4391,N_4075,N_4101);
or U4392 (N_4392,N_4183,N_4051);
and U4393 (N_4393,N_4045,N_4048);
nand U4394 (N_4394,N_4114,N_4021);
or U4395 (N_4395,N_4074,N_4083);
xor U4396 (N_4396,N_4086,N_4185);
or U4397 (N_4397,N_4115,N_4122);
or U4398 (N_4398,N_4048,N_4119);
and U4399 (N_4399,N_4032,N_4096);
nand U4400 (N_4400,N_4341,N_4309);
nand U4401 (N_4401,N_4293,N_4388);
xnor U4402 (N_4402,N_4396,N_4366);
xor U4403 (N_4403,N_4263,N_4246);
nand U4404 (N_4404,N_4382,N_4365);
and U4405 (N_4405,N_4235,N_4218);
or U4406 (N_4406,N_4286,N_4206);
and U4407 (N_4407,N_4267,N_4299);
nand U4408 (N_4408,N_4323,N_4390);
or U4409 (N_4409,N_4214,N_4321);
or U4410 (N_4410,N_4345,N_4250);
nand U4411 (N_4411,N_4335,N_4387);
nand U4412 (N_4412,N_4330,N_4240);
or U4413 (N_4413,N_4236,N_4278);
nand U4414 (N_4414,N_4255,N_4301);
xor U4415 (N_4415,N_4319,N_4205);
or U4416 (N_4416,N_4303,N_4350);
and U4417 (N_4417,N_4326,N_4312);
and U4418 (N_4418,N_4351,N_4363);
nand U4419 (N_4419,N_4295,N_4360);
or U4420 (N_4420,N_4339,N_4216);
nand U4421 (N_4421,N_4227,N_4313);
xor U4422 (N_4422,N_4222,N_4308);
xor U4423 (N_4423,N_4234,N_4220);
nand U4424 (N_4424,N_4362,N_4364);
and U4425 (N_4425,N_4392,N_4356);
nand U4426 (N_4426,N_4386,N_4252);
nand U4427 (N_4427,N_4297,N_4268);
and U4428 (N_4428,N_4219,N_4348);
or U4429 (N_4429,N_4274,N_4296);
or U4430 (N_4430,N_4361,N_4324);
xor U4431 (N_4431,N_4398,N_4343);
nand U4432 (N_4432,N_4352,N_4336);
nor U4433 (N_4433,N_4359,N_4254);
or U4434 (N_4434,N_4358,N_4311);
and U4435 (N_4435,N_4317,N_4210);
or U4436 (N_4436,N_4258,N_4389);
xor U4437 (N_4437,N_4229,N_4273);
xnor U4438 (N_4438,N_4318,N_4344);
nand U4439 (N_4439,N_4300,N_4269);
nor U4440 (N_4440,N_4393,N_4338);
or U4441 (N_4441,N_4237,N_4249);
xor U4442 (N_4442,N_4231,N_4283);
or U4443 (N_4443,N_4251,N_4287);
or U4444 (N_4444,N_4367,N_4353);
or U4445 (N_4445,N_4337,N_4349);
nand U4446 (N_4446,N_4232,N_4381);
nor U4447 (N_4447,N_4298,N_4376);
or U4448 (N_4448,N_4280,N_4354);
nand U4449 (N_4449,N_4207,N_4332);
xor U4450 (N_4450,N_4355,N_4257);
or U4451 (N_4451,N_4265,N_4346);
nor U4452 (N_4452,N_4290,N_4200);
nor U4453 (N_4453,N_4377,N_4256);
and U4454 (N_4454,N_4285,N_4310);
nand U4455 (N_4455,N_4371,N_4275);
and U4456 (N_4456,N_4325,N_4281);
or U4457 (N_4457,N_4347,N_4380);
nand U4458 (N_4458,N_4209,N_4375);
nor U4459 (N_4459,N_4245,N_4378);
nor U4460 (N_4460,N_4368,N_4394);
nor U4461 (N_4461,N_4284,N_4230);
or U4462 (N_4462,N_4391,N_4253);
xnor U4463 (N_4463,N_4333,N_4276);
nor U4464 (N_4464,N_4395,N_4316);
or U4465 (N_4465,N_4288,N_4292);
or U4466 (N_4466,N_4320,N_4329);
or U4467 (N_4467,N_4202,N_4397);
nand U4468 (N_4468,N_4305,N_4277);
nand U4469 (N_4469,N_4370,N_4244);
xor U4470 (N_4470,N_4331,N_4294);
and U4471 (N_4471,N_4233,N_4279);
nor U4472 (N_4472,N_4282,N_4208);
or U4473 (N_4473,N_4306,N_4289);
or U4474 (N_4474,N_4259,N_4357);
and U4475 (N_4475,N_4322,N_4248);
or U4476 (N_4476,N_4262,N_4201);
xor U4477 (N_4477,N_4374,N_4241);
nand U4478 (N_4478,N_4307,N_4247);
nand U4479 (N_4479,N_4261,N_4224);
and U4480 (N_4480,N_4264,N_4228);
and U4481 (N_4481,N_4243,N_4223);
nand U4482 (N_4482,N_4373,N_4383);
nand U4483 (N_4483,N_4242,N_4213);
nor U4484 (N_4484,N_4204,N_4304);
or U4485 (N_4485,N_4369,N_4226);
xor U4486 (N_4486,N_4342,N_4239);
or U4487 (N_4487,N_4379,N_4225);
or U4488 (N_4488,N_4334,N_4212);
nand U4489 (N_4489,N_4399,N_4328);
xor U4490 (N_4490,N_4266,N_4327);
nand U4491 (N_4491,N_4211,N_4314);
or U4492 (N_4492,N_4203,N_4271);
and U4493 (N_4493,N_4291,N_4302);
and U4494 (N_4494,N_4217,N_4340);
or U4495 (N_4495,N_4221,N_4272);
nor U4496 (N_4496,N_4385,N_4238);
nor U4497 (N_4497,N_4260,N_4215);
or U4498 (N_4498,N_4315,N_4384);
or U4499 (N_4499,N_4270,N_4372);
nand U4500 (N_4500,N_4200,N_4204);
xnor U4501 (N_4501,N_4358,N_4246);
nand U4502 (N_4502,N_4230,N_4252);
and U4503 (N_4503,N_4381,N_4289);
nand U4504 (N_4504,N_4340,N_4365);
xnor U4505 (N_4505,N_4311,N_4333);
nor U4506 (N_4506,N_4342,N_4297);
nand U4507 (N_4507,N_4279,N_4340);
xnor U4508 (N_4508,N_4214,N_4208);
or U4509 (N_4509,N_4397,N_4389);
xor U4510 (N_4510,N_4247,N_4303);
or U4511 (N_4511,N_4249,N_4385);
and U4512 (N_4512,N_4299,N_4293);
xor U4513 (N_4513,N_4290,N_4248);
and U4514 (N_4514,N_4360,N_4351);
nor U4515 (N_4515,N_4329,N_4308);
or U4516 (N_4516,N_4291,N_4260);
xor U4517 (N_4517,N_4387,N_4303);
xnor U4518 (N_4518,N_4239,N_4221);
xor U4519 (N_4519,N_4373,N_4235);
and U4520 (N_4520,N_4376,N_4237);
or U4521 (N_4521,N_4282,N_4223);
xor U4522 (N_4522,N_4394,N_4302);
or U4523 (N_4523,N_4381,N_4370);
and U4524 (N_4524,N_4241,N_4319);
nor U4525 (N_4525,N_4349,N_4386);
xnor U4526 (N_4526,N_4206,N_4248);
nand U4527 (N_4527,N_4384,N_4212);
or U4528 (N_4528,N_4250,N_4305);
or U4529 (N_4529,N_4275,N_4258);
and U4530 (N_4530,N_4382,N_4290);
xor U4531 (N_4531,N_4302,N_4290);
or U4532 (N_4532,N_4235,N_4376);
nand U4533 (N_4533,N_4241,N_4372);
nand U4534 (N_4534,N_4212,N_4362);
nor U4535 (N_4535,N_4238,N_4211);
nand U4536 (N_4536,N_4332,N_4210);
nand U4537 (N_4537,N_4324,N_4350);
or U4538 (N_4538,N_4319,N_4264);
nor U4539 (N_4539,N_4332,N_4318);
or U4540 (N_4540,N_4253,N_4236);
and U4541 (N_4541,N_4246,N_4353);
nor U4542 (N_4542,N_4213,N_4362);
nor U4543 (N_4543,N_4388,N_4224);
or U4544 (N_4544,N_4340,N_4335);
nor U4545 (N_4545,N_4225,N_4390);
xor U4546 (N_4546,N_4306,N_4318);
nand U4547 (N_4547,N_4297,N_4301);
and U4548 (N_4548,N_4312,N_4364);
nor U4549 (N_4549,N_4354,N_4285);
and U4550 (N_4550,N_4227,N_4390);
and U4551 (N_4551,N_4394,N_4356);
nor U4552 (N_4552,N_4250,N_4244);
nand U4553 (N_4553,N_4315,N_4251);
nor U4554 (N_4554,N_4367,N_4287);
nor U4555 (N_4555,N_4326,N_4251);
nor U4556 (N_4556,N_4220,N_4250);
nor U4557 (N_4557,N_4337,N_4282);
nand U4558 (N_4558,N_4249,N_4339);
or U4559 (N_4559,N_4255,N_4294);
nand U4560 (N_4560,N_4247,N_4294);
nor U4561 (N_4561,N_4271,N_4368);
nand U4562 (N_4562,N_4342,N_4358);
xnor U4563 (N_4563,N_4378,N_4351);
or U4564 (N_4564,N_4382,N_4275);
nand U4565 (N_4565,N_4346,N_4254);
xnor U4566 (N_4566,N_4269,N_4345);
nand U4567 (N_4567,N_4295,N_4331);
xnor U4568 (N_4568,N_4294,N_4364);
nand U4569 (N_4569,N_4227,N_4266);
xnor U4570 (N_4570,N_4242,N_4332);
nand U4571 (N_4571,N_4357,N_4356);
nand U4572 (N_4572,N_4288,N_4340);
nand U4573 (N_4573,N_4383,N_4233);
nand U4574 (N_4574,N_4333,N_4231);
xor U4575 (N_4575,N_4223,N_4391);
and U4576 (N_4576,N_4303,N_4354);
nor U4577 (N_4577,N_4344,N_4261);
nor U4578 (N_4578,N_4303,N_4365);
nand U4579 (N_4579,N_4243,N_4273);
xor U4580 (N_4580,N_4279,N_4296);
nand U4581 (N_4581,N_4317,N_4376);
nand U4582 (N_4582,N_4280,N_4370);
nand U4583 (N_4583,N_4282,N_4303);
nand U4584 (N_4584,N_4305,N_4244);
and U4585 (N_4585,N_4328,N_4376);
nor U4586 (N_4586,N_4344,N_4396);
nor U4587 (N_4587,N_4204,N_4332);
and U4588 (N_4588,N_4240,N_4263);
nor U4589 (N_4589,N_4359,N_4309);
nand U4590 (N_4590,N_4251,N_4314);
nor U4591 (N_4591,N_4274,N_4397);
or U4592 (N_4592,N_4339,N_4360);
nand U4593 (N_4593,N_4351,N_4342);
nand U4594 (N_4594,N_4371,N_4310);
nor U4595 (N_4595,N_4320,N_4301);
and U4596 (N_4596,N_4357,N_4277);
or U4597 (N_4597,N_4322,N_4256);
xor U4598 (N_4598,N_4304,N_4276);
xnor U4599 (N_4599,N_4283,N_4396);
xor U4600 (N_4600,N_4571,N_4595);
nand U4601 (N_4601,N_4401,N_4457);
and U4602 (N_4602,N_4444,N_4469);
nand U4603 (N_4603,N_4577,N_4442);
nand U4604 (N_4604,N_4417,N_4539);
or U4605 (N_4605,N_4541,N_4565);
xnor U4606 (N_4606,N_4415,N_4581);
xnor U4607 (N_4607,N_4440,N_4512);
nand U4608 (N_4608,N_4479,N_4515);
or U4609 (N_4609,N_4447,N_4426);
nor U4610 (N_4610,N_4566,N_4455);
and U4611 (N_4611,N_4547,N_4575);
nand U4612 (N_4612,N_4453,N_4433);
nand U4613 (N_4613,N_4436,N_4582);
or U4614 (N_4614,N_4569,N_4475);
and U4615 (N_4615,N_4431,N_4592);
xor U4616 (N_4616,N_4496,N_4471);
xnor U4617 (N_4617,N_4410,N_4574);
nor U4618 (N_4618,N_4518,N_4553);
nand U4619 (N_4619,N_4540,N_4528);
nor U4620 (N_4620,N_4580,N_4494);
or U4621 (N_4621,N_4524,N_4591);
xnor U4622 (N_4622,N_4480,N_4400);
or U4623 (N_4623,N_4481,N_4472);
xnor U4624 (N_4624,N_4502,N_4517);
or U4625 (N_4625,N_4503,N_4414);
and U4626 (N_4626,N_4483,N_4576);
and U4627 (N_4627,N_4506,N_4519);
or U4628 (N_4628,N_4461,N_4434);
and U4629 (N_4629,N_4551,N_4543);
and U4630 (N_4630,N_4509,N_4572);
or U4631 (N_4631,N_4555,N_4559);
nand U4632 (N_4632,N_4594,N_4439);
and U4633 (N_4633,N_4467,N_4548);
nand U4634 (N_4634,N_4498,N_4516);
nor U4635 (N_4635,N_4521,N_4550);
nor U4636 (N_4636,N_4549,N_4441);
or U4637 (N_4637,N_4588,N_4449);
or U4638 (N_4638,N_4527,N_4557);
nand U4639 (N_4639,N_4424,N_4456);
xor U4640 (N_4640,N_4466,N_4584);
xor U4641 (N_4641,N_4529,N_4493);
nor U4642 (N_4642,N_4437,N_4465);
nor U4643 (N_4643,N_4507,N_4482);
or U4644 (N_4644,N_4554,N_4593);
xor U4645 (N_4645,N_4463,N_4586);
and U4646 (N_4646,N_4508,N_4407);
and U4647 (N_4647,N_4597,N_4545);
nand U4648 (N_4648,N_4428,N_4589);
nor U4649 (N_4649,N_4448,N_4564);
nor U4650 (N_4650,N_4435,N_4462);
nor U4651 (N_4651,N_4531,N_4489);
nand U4652 (N_4652,N_4510,N_4533);
or U4653 (N_4653,N_4487,N_4599);
nor U4654 (N_4654,N_4544,N_4451);
or U4655 (N_4655,N_4413,N_4470);
nor U4656 (N_4656,N_4477,N_4443);
and U4657 (N_4657,N_4523,N_4425);
nor U4658 (N_4658,N_4535,N_4596);
xnor U4659 (N_4659,N_4537,N_4526);
xnor U4660 (N_4660,N_4427,N_4485);
nor U4661 (N_4661,N_4474,N_4567);
xnor U4662 (N_4662,N_4430,N_4459);
and U4663 (N_4663,N_4402,N_4450);
xnor U4664 (N_4664,N_4546,N_4416);
nor U4665 (N_4665,N_4538,N_4499);
nand U4666 (N_4666,N_4558,N_4573);
or U4667 (N_4667,N_4570,N_4583);
nor U4668 (N_4668,N_4411,N_4495);
xnor U4669 (N_4669,N_4492,N_4542);
nand U4670 (N_4670,N_4412,N_4408);
and U4671 (N_4671,N_4590,N_4490);
xor U4672 (N_4672,N_4561,N_4585);
nor U4673 (N_4673,N_4464,N_4404);
xor U4674 (N_4674,N_4418,N_4598);
nor U4675 (N_4675,N_4514,N_4587);
or U4676 (N_4676,N_4468,N_4432);
nand U4677 (N_4677,N_4504,N_4520);
and U4678 (N_4678,N_4473,N_4491);
nand U4679 (N_4679,N_4488,N_4478);
nand U4680 (N_4680,N_4568,N_4458);
xor U4681 (N_4681,N_4438,N_4405);
nand U4682 (N_4682,N_4534,N_4445);
nor U4683 (N_4683,N_4560,N_4452);
xnor U4684 (N_4684,N_4476,N_4552);
nor U4685 (N_4685,N_4532,N_4446);
or U4686 (N_4686,N_4536,N_4563);
and U4687 (N_4687,N_4505,N_4484);
or U4688 (N_4688,N_4522,N_4513);
or U4689 (N_4689,N_4530,N_4501);
nor U4690 (N_4690,N_4406,N_4511);
nor U4691 (N_4691,N_4422,N_4578);
nand U4692 (N_4692,N_4421,N_4429);
xor U4693 (N_4693,N_4419,N_4579);
xnor U4694 (N_4694,N_4500,N_4403);
nand U4695 (N_4695,N_4556,N_4497);
xnor U4696 (N_4696,N_4486,N_4454);
nor U4697 (N_4697,N_4525,N_4423);
nor U4698 (N_4698,N_4562,N_4460);
or U4699 (N_4699,N_4420,N_4409);
xor U4700 (N_4700,N_4420,N_4521);
nand U4701 (N_4701,N_4420,N_4588);
xnor U4702 (N_4702,N_4520,N_4460);
and U4703 (N_4703,N_4435,N_4571);
and U4704 (N_4704,N_4582,N_4557);
or U4705 (N_4705,N_4564,N_4402);
nand U4706 (N_4706,N_4446,N_4586);
and U4707 (N_4707,N_4509,N_4577);
and U4708 (N_4708,N_4541,N_4570);
and U4709 (N_4709,N_4534,N_4504);
or U4710 (N_4710,N_4517,N_4518);
nand U4711 (N_4711,N_4457,N_4592);
or U4712 (N_4712,N_4586,N_4478);
and U4713 (N_4713,N_4454,N_4583);
and U4714 (N_4714,N_4441,N_4543);
nor U4715 (N_4715,N_4435,N_4599);
nor U4716 (N_4716,N_4512,N_4561);
or U4717 (N_4717,N_4478,N_4573);
nor U4718 (N_4718,N_4599,N_4467);
nor U4719 (N_4719,N_4504,N_4543);
nor U4720 (N_4720,N_4441,N_4464);
or U4721 (N_4721,N_4507,N_4540);
xor U4722 (N_4722,N_4415,N_4528);
or U4723 (N_4723,N_4574,N_4564);
or U4724 (N_4724,N_4453,N_4449);
xor U4725 (N_4725,N_4521,N_4405);
nor U4726 (N_4726,N_4444,N_4513);
xnor U4727 (N_4727,N_4437,N_4467);
nor U4728 (N_4728,N_4562,N_4510);
nand U4729 (N_4729,N_4438,N_4543);
xor U4730 (N_4730,N_4436,N_4422);
and U4731 (N_4731,N_4536,N_4534);
or U4732 (N_4732,N_4594,N_4558);
or U4733 (N_4733,N_4426,N_4566);
nand U4734 (N_4734,N_4413,N_4596);
nand U4735 (N_4735,N_4560,N_4427);
nor U4736 (N_4736,N_4405,N_4539);
or U4737 (N_4737,N_4517,N_4432);
xor U4738 (N_4738,N_4457,N_4513);
nor U4739 (N_4739,N_4536,N_4585);
and U4740 (N_4740,N_4456,N_4420);
nor U4741 (N_4741,N_4462,N_4512);
or U4742 (N_4742,N_4591,N_4519);
nand U4743 (N_4743,N_4501,N_4489);
or U4744 (N_4744,N_4446,N_4431);
nand U4745 (N_4745,N_4488,N_4501);
and U4746 (N_4746,N_4525,N_4589);
nor U4747 (N_4747,N_4559,N_4592);
nand U4748 (N_4748,N_4578,N_4598);
xnor U4749 (N_4749,N_4528,N_4440);
xnor U4750 (N_4750,N_4482,N_4595);
nand U4751 (N_4751,N_4553,N_4434);
or U4752 (N_4752,N_4533,N_4444);
nor U4753 (N_4753,N_4535,N_4489);
xor U4754 (N_4754,N_4500,N_4591);
or U4755 (N_4755,N_4533,N_4592);
nand U4756 (N_4756,N_4415,N_4547);
xnor U4757 (N_4757,N_4479,N_4431);
nor U4758 (N_4758,N_4497,N_4447);
and U4759 (N_4759,N_4436,N_4481);
and U4760 (N_4760,N_4428,N_4571);
or U4761 (N_4761,N_4448,N_4540);
and U4762 (N_4762,N_4505,N_4582);
xnor U4763 (N_4763,N_4478,N_4464);
xnor U4764 (N_4764,N_4594,N_4426);
nand U4765 (N_4765,N_4510,N_4429);
nand U4766 (N_4766,N_4597,N_4427);
xnor U4767 (N_4767,N_4499,N_4513);
or U4768 (N_4768,N_4494,N_4577);
nor U4769 (N_4769,N_4491,N_4490);
nor U4770 (N_4770,N_4521,N_4597);
xnor U4771 (N_4771,N_4487,N_4409);
nor U4772 (N_4772,N_4501,N_4441);
xnor U4773 (N_4773,N_4501,N_4484);
xnor U4774 (N_4774,N_4426,N_4572);
nand U4775 (N_4775,N_4464,N_4466);
nor U4776 (N_4776,N_4569,N_4524);
nor U4777 (N_4777,N_4427,N_4496);
nor U4778 (N_4778,N_4438,N_4490);
nor U4779 (N_4779,N_4481,N_4533);
nor U4780 (N_4780,N_4442,N_4476);
nor U4781 (N_4781,N_4531,N_4572);
nand U4782 (N_4782,N_4425,N_4567);
and U4783 (N_4783,N_4403,N_4438);
nand U4784 (N_4784,N_4546,N_4401);
or U4785 (N_4785,N_4528,N_4565);
or U4786 (N_4786,N_4505,N_4455);
xnor U4787 (N_4787,N_4530,N_4595);
or U4788 (N_4788,N_4459,N_4528);
or U4789 (N_4789,N_4510,N_4532);
or U4790 (N_4790,N_4433,N_4543);
nand U4791 (N_4791,N_4415,N_4459);
xor U4792 (N_4792,N_4568,N_4424);
nor U4793 (N_4793,N_4540,N_4549);
xor U4794 (N_4794,N_4485,N_4522);
and U4795 (N_4795,N_4423,N_4557);
or U4796 (N_4796,N_4504,N_4583);
and U4797 (N_4797,N_4453,N_4564);
and U4798 (N_4798,N_4469,N_4421);
or U4799 (N_4799,N_4433,N_4405);
or U4800 (N_4800,N_4653,N_4697);
xor U4801 (N_4801,N_4768,N_4666);
nand U4802 (N_4802,N_4709,N_4628);
or U4803 (N_4803,N_4613,N_4725);
nor U4804 (N_4804,N_4771,N_4609);
xnor U4805 (N_4805,N_4680,N_4606);
nand U4806 (N_4806,N_4649,N_4700);
or U4807 (N_4807,N_4636,N_4671);
xor U4808 (N_4808,N_4728,N_4756);
or U4809 (N_4809,N_4748,N_4717);
nand U4810 (N_4810,N_4757,N_4678);
nor U4811 (N_4811,N_4611,N_4705);
or U4812 (N_4812,N_4670,N_4618);
xnor U4813 (N_4813,N_4690,N_4601);
nor U4814 (N_4814,N_4719,N_4754);
or U4815 (N_4815,N_4752,N_4746);
nor U4816 (N_4816,N_4655,N_4600);
nand U4817 (N_4817,N_4731,N_4646);
xor U4818 (N_4818,N_4763,N_4774);
or U4819 (N_4819,N_4724,N_4647);
or U4820 (N_4820,N_4762,N_4707);
nor U4821 (N_4821,N_4755,N_4723);
or U4822 (N_4822,N_4704,N_4753);
nor U4823 (N_4823,N_4749,N_4665);
nor U4824 (N_4824,N_4750,N_4651);
nand U4825 (N_4825,N_4619,N_4638);
nor U4826 (N_4826,N_4621,N_4727);
xnor U4827 (N_4827,N_4694,N_4760);
or U4828 (N_4828,N_4738,N_4782);
nand U4829 (N_4829,N_4699,N_4730);
xnor U4830 (N_4830,N_4688,N_4726);
xor U4831 (N_4831,N_4658,N_4789);
nor U4832 (N_4832,N_4720,N_4681);
or U4833 (N_4833,N_4634,N_4716);
or U4834 (N_4834,N_4603,N_4793);
nor U4835 (N_4835,N_4626,N_4759);
or U4836 (N_4836,N_4764,N_4721);
nor U4837 (N_4837,N_4663,N_4652);
nand U4838 (N_4838,N_4775,N_4718);
and U4839 (N_4839,N_4711,N_4790);
and U4840 (N_4840,N_4604,N_4769);
and U4841 (N_4841,N_4676,N_4677);
xor U4842 (N_4842,N_4695,N_4796);
xnor U4843 (N_4843,N_4777,N_4708);
or U4844 (N_4844,N_4672,N_4605);
nor U4845 (N_4845,N_4622,N_4650);
nor U4846 (N_4846,N_4644,N_4693);
and U4847 (N_4847,N_4686,N_4641);
nor U4848 (N_4848,N_4740,N_4743);
nand U4849 (N_4849,N_4770,N_4675);
nand U4850 (N_4850,N_4722,N_4703);
nor U4851 (N_4851,N_4627,N_4661);
or U4852 (N_4852,N_4691,N_4631);
and U4853 (N_4853,N_4625,N_4736);
nand U4854 (N_4854,N_4714,N_4766);
xor U4855 (N_4855,N_4667,N_4778);
or U4856 (N_4856,N_4662,N_4660);
or U4857 (N_4857,N_4642,N_4787);
and U4858 (N_4858,N_4732,N_4773);
xor U4859 (N_4859,N_4610,N_4794);
or U4860 (N_4860,N_4780,N_4602);
and U4861 (N_4861,N_4702,N_4698);
nor U4862 (N_4862,N_4633,N_4639);
nor U4863 (N_4863,N_4735,N_4706);
nor U4864 (N_4864,N_4684,N_4623);
nor U4865 (N_4865,N_4786,N_4645);
and U4866 (N_4866,N_4729,N_4744);
xor U4867 (N_4867,N_4765,N_4772);
nor U4868 (N_4868,N_4664,N_4657);
xnor U4869 (N_4869,N_4669,N_4791);
nor U4870 (N_4870,N_4692,N_4781);
nor U4871 (N_4871,N_4632,N_4734);
and U4872 (N_4872,N_4799,N_4624);
and U4873 (N_4873,N_4614,N_4620);
xnor U4874 (N_4874,N_4612,N_4715);
xnor U4875 (N_4875,N_4654,N_4685);
or U4876 (N_4876,N_4784,N_4798);
nor U4877 (N_4877,N_4785,N_4795);
nor U4878 (N_4878,N_4733,N_4629);
or U4879 (N_4879,N_4643,N_4761);
xnor U4880 (N_4880,N_4751,N_4674);
and U4881 (N_4881,N_4689,N_4608);
xnor U4882 (N_4882,N_4696,N_4712);
nand U4883 (N_4883,N_4741,N_4668);
nand U4884 (N_4884,N_4616,N_4747);
nand U4885 (N_4885,N_4745,N_4648);
nor U4886 (N_4886,N_4713,N_4687);
nand U4887 (N_4887,N_4797,N_4792);
or U4888 (N_4888,N_4656,N_4779);
xnor U4889 (N_4889,N_4701,N_4788);
xnor U4890 (N_4890,N_4607,N_4739);
xnor U4891 (N_4891,N_4682,N_4767);
or U4892 (N_4892,N_4758,N_4659);
and U4893 (N_4893,N_4673,N_4635);
xor U4894 (N_4894,N_4710,N_4637);
and U4895 (N_4895,N_4776,N_4783);
nand U4896 (N_4896,N_4617,N_4640);
and U4897 (N_4897,N_4615,N_4683);
nor U4898 (N_4898,N_4630,N_4737);
nor U4899 (N_4899,N_4742,N_4679);
or U4900 (N_4900,N_4630,N_4794);
nand U4901 (N_4901,N_4658,N_4716);
or U4902 (N_4902,N_4696,N_4749);
and U4903 (N_4903,N_4691,N_4698);
nand U4904 (N_4904,N_4700,N_4609);
or U4905 (N_4905,N_4772,N_4730);
and U4906 (N_4906,N_4710,N_4626);
xnor U4907 (N_4907,N_4720,N_4769);
nand U4908 (N_4908,N_4642,N_4718);
nor U4909 (N_4909,N_4703,N_4610);
nand U4910 (N_4910,N_4601,N_4747);
or U4911 (N_4911,N_4621,N_4761);
nor U4912 (N_4912,N_4713,N_4646);
nor U4913 (N_4913,N_4715,N_4734);
or U4914 (N_4914,N_4612,N_4783);
nor U4915 (N_4915,N_4717,N_4622);
or U4916 (N_4916,N_4727,N_4742);
xnor U4917 (N_4917,N_4791,N_4691);
xnor U4918 (N_4918,N_4680,N_4638);
nand U4919 (N_4919,N_4651,N_4640);
nor U4920 (N_4920,N_4629,N_4600);
nand U4921 (N_4921,N_4733,N_4644);
xnor U4922 (N_4922,N_4701,N_4625);
nand U4923 (N_4923,N_4760,N_4749);
and U4924 (N_4924,N_4701,N_4790);
nand U4925 (N_4925,N_4762,N_4667);
nand U4926 (N_4926,N_4636,N_4691);
or U4927 (N_4927,N_4774,N_4736);
nor U4928 (N_4928,N_4603,N_4616);
nand U4929 (N_4929,N_4740,N_4645);
xor U4930 (N_4930,N_4715,N_4732);
nand U4931 (N_4931,N_4643,N_4716);
nand U4932 (N_4932,N_4609,N_4778);
nor U4933 (N_4933,N_4679,N_4726);
or U4934 (N_4934,N_4639,N_4621);
and U4935 (N_4935,N_4624,N_4706);
nand U4936 (N_4936,N_4630,N_4663);
nor U4937 (N_4937,N_4641,N_4647);
and U4938 (N_4938,N_4701,N_4638);
nor U4939 (N_4939,N_4703,N_4783);
nand U4940 (N_4940,N_4621,N_4687);
nor U4941 (N_4941,N_4604,N_4666);
nand U4942 (N_4942,N_4619,N_4604);
nand U4943 (N_4943,N_4706,N_4795);
nor U4944 (N_4944,N_4778,N_4676);
nand U4945 (N_4945,N_4692,N_4616);
xnor U4946 (N_4946,N_4795,N_4733);
and U4947 (N_4947,N_4754,N_4679);
nand U4948 (N_4948,N_4633,N_4624);
or U4949 (N_4949,N_4792,N_4776);
or U4950 (N_4950,N_4720,N_4678);
xnor U4951 (N_4951,N_4619,N_4600);
nor U4952 (N_4952,N_4769,N_4704);
xor U4953 (N_4953,N_4627,N_4782);
and U4954 (N_4954,N_4661,N_4795);
nand U4955 (N_4955,N_4724,N_4730);
or U4956 (N_4956,N_4721,N_4677);
xor U4957 (N_4957,N_4764,N_4796);
and U4958 (N_4958,N_4748,N_4767);
or U4959 (N_4959,N_4789,N_4777);
nand U4960 (N_4960,N_4652,N_4670);
nor U4961 (N_4961,N_4741,N_4779);
and U4962 (N_4962,N_4770,N_4633);
nor U4963 (N_4963,N_4772,N_4762);
nor U4964 (N_4964,N_4723,N_4663);
and U4965 (N_4965,N_4608,N_4658);
nor U4966 (N_4966,N_4740,N_4785);
nand U4967 (N_4967,N_4616,N_4625);
nand U4968 (N_4968,N_4787,N_4685);
nand U4969 (N_4969,N_4607,N_4783);
or U4970 (N_4970,N_4685,N_4783);
xor U4971 (N_4971,N_4750,N_4688);
xnor U4972 (N_4972,N_4629,N_4649);
or U4973 (N_4973,N_4615,N_4768);
and U4974 (N_4974,N_4759,N_4667);
nor U4975 (N_4975,N_4601,N_4661);
nand U4976 (N_4976,N_4716,N_4785);
nor U4977 (N_4977,N_4670,N_4691);
and U4978 (N_4978,N_4693,N_4652);
xor U4979 (N_4979,N_4656,N_4622);
nor U4980 (N_4980,N_4783,N_4792);
or U4981 (N_4981,N_4684,N_4651);
nand U4982 (N_4982,N_4783,N_4794);
xor U4983 (N_4983,N_4723,N_4641);
xnor U4984 (N_4984,N_4725,N_4719);
or U4985 (N_4985,N_4730,N_4773);
nand U4986 (N_4986,N_4744,N_4683);
nand U4987 (N_4987,N_4778,N_4756);
or U4988 (N_4988,N_4685,N_4756);
nor U4989 (N_4989,N_4679,N_4715);
xor U4990 (N_4990,N_4772,N_4725);
and U4991 (N_4991,N_4605,N_4697);
or U4992 (N_4992,N_4799,N_4671);
nor U4993 (N_4993,N_4630,N_4651);
and U4994 (N_4994,N_4648,N_4670);
xor U4995 (N_4995,N_4786,N_4784);
or U4996 (N_4996,N_4773,N_4650);
xnor U4997 (N_4997,N_4643,N_4764);
or U4998 (N_4998,N_4782,N_4699);
xor U4999 (N_4999,N_4722,N_4751);
nand U5000 (N_5000,N_4973,N_4976);
nor U5001 (N_5001,N_4813,N_4902);
nand U5002 (N_5002,N_4962,N_4847);
xnor U5003 (N_5003,N_4836,N_4920);
or U5004 (N_5004,N_4959,N_4971);
nand U5005 (N_5005,N_4824,N_4979);
and U5006 (N_5006,N_4879,N_4963);
and U5007 (N_5007,N_4818,N_4896);
xnor U5008 (N_5008,N_4881,N_4840);
or U5009 (N_5009,N_4849,N_4834);
and U5010 (N_5010,N_4980,N_4974);
and U5011 (N_5011,N_4841,N_4821);
or U5012 (N_5012,N_4995,N_4858);
nand U5013 (N_5013,N_4871,N_4884);
nor U5014 (N_5014,N_4823,N_4877);
nor U5015 (N_5015,N_4904,N_4956);
and U5016 (N_5016,N_4855,N_4942);
nor U5017 (N_5017,N_4872,N_4955);
nand U5018 (N_5018,N_4989,N_4977);
xnor U5019 (N_5019,N_4965,N_4897);
nand U5020 (N_5020,N_4819,N_4814);
or U5021 (N_5021,N_4915,N_4999);
and U5022 (N_5022,N_4891,N_4831);
xor U5023 (N_5023,N_4909,N_4903);
nand U5024 (N_5024,N_4870,N_4857);
xor U5025 (N_5025,N_4945,N_4865);
or U5026 (N_5026,N_4894,N_4827);
or U5027 (N_5027,N_4961,N_4862);
nor U5028 (N_5028,N_4820,N_4993);
nor U5029 (N_5029,N_4816,N_4987);
and U5030 (N_5030,N_4856,N_4806);
nand U5031 (N_5031,N_4975,N_4889);
xnor U5032 (N_5032,N_4907,N_4917);
nand U5033 (N_5033,N_4922,N_4859);
or U5034 (N_5034,N_4940,N_4938);
nor U5035 (N_5035,N_4941,N_4804);
xnor U5036 (N_5036,N_4828,N_4800);
xor U5037 (N_5037,N_4805,N_4851);
and U5038 (N_5038,N_4960,N_4867);
nand U5039 (N_5039,N_4924,N_4803);
and U5040 (N_5040,N_4936,N_4983);
xnor U5041 (N_5041,N_4815,N_4978);
or U5042 (N_5042,N_4913,N_4817);
or U5043 (N_5043,N_4811,N_4900);
and U5044 (N_5044,N_4927,N_4893);
nand U5045 (N_5045,N_4886,N_4967);
and U5046 (N_5046,N_4997,N_4845);
nor U5047 (N_5047,N_4990,N_4829);
xor U5048 (N_5048,N_4966,N_4944);
nor U5049 (N_5049,N_4848,N_4808);
and U5050 (N_5050,N_4876,N_4918);
nor U5051 (N_5051,N_4985,N_4998);
nor U5052 (N_5052,N_4935,N_4899);
or U5053 (N_5053,N_4933,N_4996);
nand U5054 (N_5054,N_4910,N_4954);
nand U5055 (N_5055,N_4957,N_4992);
nor U5056 (N_5056,N_4929,N_4892);
nor U5057 (N_5057,N_4868,N_4890);
nor U5058 (N_5058,N_4968,N_4825);
nand U5059 (N_5059,N_4835,N_4947);
and U5060 (N_5060,N_4873,N_4964);
and U5061 (N_5061,N_4949,N_4844);
and U5062 (N_5062,N_4842,N_4852);
xor U5063 (N_5063,N_4953,N_4875);
nor U5064 (N_5064,N_4991,N_4943);
nor U5065 (N_5065,N_4928,N_4994);
nand U5066 (N_5066,N_4958,N_4853);
xnor U5067 (N_5067,N_4926,N_4812);
xnor U5068 (N_5068,N_4946,N_4986);
xor U5069 (N_5069,N_4981,N_4860);
nand U5070 (N_5070,N_4911,N_4908);
and U5071 (N_5071,N_4802,N_4984);
and U5072 (N_5072,N_4937,N_4901);
or U5073 (N_5073,N_4822,N_4846);
or U5074 (N_5074,N_4912,N_4861);
or U5075 (N_5075,N_4864,N_4914);
xor U5076 (N_5076,N_4898,N_4838);
nor U5077 (N_5077,N_4930,N_4801);
or U5078 (N_5078,N_4969,N_4916);
xor U5079 (N_5079,N_4837,N_4931);
nand U5080 (N_5080,N_4970,N_4887);
xnor U5081 (N_5081,N_4830,N_4939);
and U5082 (N_5082,N_4906,N_4882);
nand U5083 (N_5083,N_4863,N_4826);
nand U5084 (N_5084,N_4866,N_4885);
nand U5085 (N_5085,N_4932,N_4988);
nand U5086 (N_5086,N_4832,N_4948);
xnor U5087 (N_5087,N_4921,N_4895);
xnor U5088 (N_5088,N_4839,N_4809);
nand U5089 (N_5089,N_4888,N_4833);
and U5090 (N_5090,N_4843,N_4854);
nand U5091 (N_5091,N_4923,N_4880);
xor U5092 (N_5092,N_4950,N_4934);
nand U5093 (N_5093,N_4807,N_4850);
nor U5094 (N_5094,N_4810,N_4951);
nor U5095 (N_5095,N_4874,N_4972);
and U5096 (N_5096,N_4905,N_4869);
or U5097 (N_5097,N_4952,N_4982);
or U5098 (N_5098,N_4925,N_4883);
nand U5099 (N_5099,N_4878,N_4919);
xnor U5100 (N_5100,N_4847,N_4849);
nand U5101 (N_5101,N_4887,N_4873);
and U5102 (N_5102,N_4822,N_4860);
or U5103 (N_5103,N_4839,N_4949);
or U5104 (N_5104,N_4892,N_4849);
xnor U5105 (N_5105,N_4964,N_4872);
nand U5106 (N_5106,N_4843,N_4867);
and U5107 (N_5107,N_4851,N_4802);
and U5108 (N_5108,N_4903,N_4955);
xor U5109 (N_5109,N_4827,N_4981);
xnor U5110 (N_5110,N_4980,N_4840);
xor U5111 (N_5111,N_4863,N_4952);
nor U5112 (N_5112,N_4939,N_4887);
and U5113 (N_5113,N_4903,N_4889);
or U5114 (N_5114,N_4920,N_4915);
nand U5115 (N_5115,N_4879,N_4896);
and U5116 (N_5116,N_4984,N_4844);
xnor U5117 (N_5117,N_4983,N_4829);
nand U5118 (N_5118,N_4901,N_4858);
and U5119 (N_5119,N_4912,N_4914);
or U5120 (N_5120,N_4931,N_4908);
xor U5121 (N_5121,N_4883,N_4800);
and U5122 (N_5122,N_4908,N_4980);
xor U5123 (N_5123,N_4906,N_4915);
xnor U5124 (N_5124,N_4824,N_4987);
nand U5125 (N_5125,N_4910,N_4996);
nor U5126 (N_5126,N_4830,N_4805);
and U5127 (N_5127,N_4904,N_4941);
xor U5128 (N_5128,N_4829,N_4997);
xor U5129 (N_5129,N_4842,N_4870);
and U5130 (N_5130,N_4923,N_4887);
or U5131 (N_5131,N_4914,N_4855);
xor U5132 (N_5132,N_4846,N_4843);
and U5133 (N_5133,N_4932,N_4826);
nand U5134 (N_5134,N_4958,N_4886);
nand U5135 (N_5135,N_4961,N_4955);
nand U5136 (N_5136,N_4968,N_4809);
xnor U5137 (N_5137,N_4889,N_4932);
nand U5138 (N_5138,N_4995,N_4951);
and U5139 (N_5139,N_4974,N_4869);
nand U5140 (N_5140,N_4914,N_4821);
xor U5141 (N_5141,N_4997,N_4805);
or U5142 (N_5142,N_4885,N_4954);
and U5143 (N_5143,N_4978,N_4887);
or U5144 (N_5144,N_4935,N_4957);
nor U5145 (N_5145,N_4821,N_4974);
nand U5146 (N_5146,N_4860,N_4973);
xor U5147 (N_5147,N_4920,N_4949);
and U5148 (N_5148,N_4870,N_4935);
nor U5149 (N_5149,N_4958,N_4861);
nand U5150 (N_5150,N_4939,N_4972);
nor U5151 (N_5151,N_4815,N_4868);
nand U5152 (N_5152,N_4927,N_4957);
xor U5153 (N_5153,N_4971,N_4976);
nor U5154 (N_5154,N_4971,N_4887);
nand U5155 (N_5155,N_4948,N_4853);
nand U5156 (N_5156,N_4929,N_4989);
nand U5157 (N_5157,N_4998,N_4951);
nand U5158 (N_5158,N_4995,N_4831);
nand U5159 (N_5159,N_4905,N_4817);
xnor U5160 (N_5160,N_4958,N_4906);
or U5161 (N_5161,N_4908,N_4960);
nand U5162 (N_5162,N_4807,N_4844);
xor U5163 (N_5163,N_4862,N_4811);
or U5164 (N_5164,N_4849,N_4871);
nand U5165 (N_5165,N_4892,N_4824);
and U5166 (N_5166,N_4878,N_4946);
or U5167 (N_5167,N_4929,N_4946);
nand U5168 (N_5168,N_4863,N_4815);
or U5169 (N_5169,N_4845,N_4981);
nor U5170 (N_5170,N_4927,N_4926);
nor U5171 (N_5171,N_4833,N_4876);
and U5172 (N_5172,N_4923,N_4998);
and U5173 (N_5173,N_4943,N_4930);
and U5174 (N_5174,N_4965,N_4819);
and U5175 (N_5175,N_4869,N_4835);
and U5176 (N_5176,N_4857,N_4829);
nand U5177 (N_5177,N_4937,N_4833);
nor U5178 (N_5178,N_4993,N_4946);
xnor U5179 (N_5179,N_4983,N_4808);
xor U5180 (N_5180,N_4926,N_4800);
nor U5181 (N_5181,N_4957,N_4824);
or U5182 (N_5182,N_4899,N_4894);
or U5183 (N_5183,N_4885,N_4845);
and U5184 (N_5184,N_4859,N_4814);
or U5185 (N_5185,N_4844,N_4920);
or U5186 (N_5186,N_4839,N_4934);
nand U5187 (N_5187,N_4895,N_4934);
nand U5188 (N_5188,N_4958,N_4810);
nor U5189 (N_5189,N_4850,N_4839);
nand U5190 (N_5190,N_4855,N_4935);
xor U5191 (N_5191,N_4854,N_4995);
xor U5192 (N_5192,N_4911,N_4947);
xor U5193 (N_5193,N_4934,N_4818);
nand U5194 (N_5194,N_4864,N_4894);
nor U5195 (N_5195,N_4982,N_4840);
xor U5196 (N_5196,N_4885,N_4817);
or U5197 (N_5197,N_4892,N_4853);
nand U5198 (N_5198,N_4893,N_4881);
and U5199 (N_5199,N_4857,N_4947);
or U5200 (N_5200,N_5156,N_5159);
nor U5201 (N_5201,N_5026,N_5035);
and U5202 (N_5202,N_5121,N_5050);
and U5203 (N_5203,N_5010,N_5029);
nand U5204 (N_5204,N_5087,N_5163);
xnor U5205 (N_5205,N_5179,N_5124);
nand U5206 (N_5206,N_5167,N_5103);
or U5207 (N_5207,N_5090,N_5018);
or U5208 (N_5208,N_5119,N_5042);
and U5209 (N_5209,N_5081,N_5068);
nand U5210 (N_5210,N_5014,N_5092);
and U5211 (N_5211,N_5065,N_5181);
nor U5212 (N_5212,N_5182,N_5079);
xor U5213 (N_5213,N_5019,N_5194);
nand U5214 (N_5214,N_5172,N_5047);
and U5215 (N_5215,N_5170,N_5171);
xor U5216 (N_5216,N_5017,N_5021);
nand U5217 (N_5217,N_5034,N_5045);
nor U5218 (N_5218,N_5073,N_5143);
xor U5219 (N_5219,N_5011,N_5084);
nand U5220 (N_5220,N_5039,N_5174);
and U5221 (N_5221,N_5036,N_5110);
xor U5222 (N_5222,N_5098,N_5193);
nand U5223 (N_5223,N_5129,N_5180);
nand U5224 (N_5224,N_5144,N_5027);
nor U5225 (N_5225,N_5096,N_5072);
nor U5226 (N_5226,N_5152,N_5107);
nor U5227 (N_5227,N_5185,N_5162);
nand U5228 (N_5228,N_5062,N_5085);
or U5229 (N_5229,N_5191,N_5127);
xnor U5230 (N_5230,N_5038,N_5115);
nor U5231 (N_5231,N_5074,N_5055);
and U5232 (N_5232,N_5016,N_5151);
or U5233 (N_5233,N_5120,N_5089);
or U5234 (N_5234,N_5177,N_5132);
or U5235 (N_5235,N_5139,N_5175);
and U5236 (N_5236,N_5161,N_5125);
xor U5237 (N_5237,N_5105,N_5028);
and U5238 (N_5238,N_5112,N_5168);
nand U5239 (N_5239,N_5199,N_5091);
nor U5240 (N_5240,N_5135,N_5069);
and U5241 (N_5241,N_5109,N_5048);
nor U5242 (N_5242,N_5195,N_5012);
and U5243 (N_5243,N_5086,N_5066);
nand U5244 (N_5244,N_5082,N_5005);
nor U5245 (N_5245,N_5056,N_5196);
nand U5246 (N_5246,N_5043,N_5190);
xor U5247 (N_5247,N_5064,N_5130);
or U5248 (N_5248,N_5013,N_5114);
and U5249 (N_5249,N_5070,N_5116);
nand U5250 (N_5250,N_5024,N_5118);
or U5251 (N_5251,N_5025,N_5032);
nand U5252 (N_5252,N_5002,N_5146);
or U5253 (N_5253,N_5145,N_5040);
nor U5254 (N_5254,N_5007,N_5009);
or U5255 (N_5255,N_5192,N_5051);
and U5256 (N_5256,N_5001,N_5111);
xnor U5257 (N_5257,N_5128,N_5154);
or U5258 (N_5258,N_5052,N_5142);
and U5259 (N_5259,N_5178,N_5150);
xor U5260 (N_5260,N_5183,N_5008);
and U5261 (N_5261,N_5100,N_5094);
xnor U5262 (N_5262,N_5067,N_5148);
xnor U5263 (N_5263,N_5102,N_5157);
and U5264 (N_5264,N_5101,N_5134);
or U5265 (N_5265,N_5058,N_5198);
nor U5266 (N_5266,N_5164,N_5189);
or U5267 (N_5267,N_5020,N_5137);
nor U5268 (N_5268,N_5080,N_5133);
xor U5269 (N_5269,N_5037,N_5097);
nor U5270 (N_5270,N_5057,N_5166);
nor U5271 (N_5271,N_5054,N_5141);
xor U5272 (N_5272,N_5044,N_5188);
nand U5273 (N_5273,N_5131,N_5030);
nand U5274 (N_5274,N_5078,N_5031);
xnor U5275 (N_5275,N_5140,N_5046);
nand U5276 (N_5276,N_5108,N_5004);
nand U5277 (N_5277,N_5076,N_5184);
and U5278 (N_5278,N_5136,N_5155);
and U5279 (N_5279,N_5153,N_5158);
and U5280 (N_5280,N_5117,N_5022);
nand U5281 (N_5281,N_5049,N_5053);
xor U5282 (N_5282,N_5197,N_5061);
and U5283 (N_5283,N_5165,N_5095);
and U5284 (N_5284,N_5160,N_5083);
nor U5285 (N_5285,N_5104,N_5138);
or U5286 (N_5286,N_5186,N_5176);
nand U5287 (N_5287,N_5169,N_5077);
xor U5288 (N_5288,N_5113,N_5122);
nand U5289 (N_5289,N_5075,N_5063);
nor U5290 (N_5290,N_5000,N_5123);
xor U5291 (N_5291,N_5060,N_5147);
xor U5292 (N_5292,N_5023,N_5071);
nor U5293 (N_5293,N_5033,N_5106);
and U5294 (N_5294,N_5099,N_5059);
nand U5295 (N_5295,N_5015,N_5173);
or U5296 (N_5296,N_5126,N_5088);
nor U5297 (N_5297,N_5149,N_5041);
nand U5298 (N_5298,N_5003,N_5093);
and U5299 (N_5299,N_5187,N_5006);
and U5300 (N_5300,N_5199,N_5046);
and U5301 (N_5301,N_5195,N_5193);
nand U5302 (N_5302,N_5185,N_5116);
and U5303 (N_5303,N_5076,N_5070);
nand U5304 (N_5304,N_5062,N_5090);
nor U5305 (N_5305,N_5132,N_5141);
and U5306 (N_5306,N_5028,N_5101);
nor U5307 (N_5307,N_5140,N_5108);
xnor U5308 (N_5308,N_5063,N_5154);
and U5309 (N_5309,N_5103,N_5184);
xnor U5310 (N_5310,N_5092,N_5125);
or U5311 (N_5311,N_5007,N_5053);
and U5312 (N_5312,N_5141,N_5194);
nand U5313 (N_5313,N_5140,N_5159);
or U5314 (N_5314,N_5085,N_5195);
or U5315 (N_5315,N_5075,N_5177);
nand U5316 (N_5316,N_5101,N_5183);
nand U5317 (N_5317,N_5123,N_5185);
and U5318 (N_5318,N_5094,N_5193);
nand U5319 (N_5319,N_5065,N_5026);
nand U5320 (N_5320,N_5166,N_5033);
xor U5321 (N_5321,N_5021,N_5035);
xor U5322 (N_5322,N_5171,N_5000);
or U5323 (N_5323,N_5076,N_5008);
or U5324 (N_5324,N_5182,N_5109);
or U5325 (N_5325,N_5087,N_5056);
nor U5326 (N_5326,N_5091,N_5007);
nand U5327 (N_5327,N_5108,N_5117);
xnor U5328 (N_5328,N_5096,N_5051);
or U5329 (N_5329,N_5041,N_5063);
or U5330 (N_5330,N_5007,N_5033);
nor U5331 (N_5331,N_5106,N_5124);
or U5332 (N_5332,N_5128,N_5169);
nor U5333 (N_5333,N_5111,N_5010);
xor U5334 (N_5334,N_5199,N_5158);
nand U5335 (N_5335,N_5070,N_5063);
xor U5336 (N_5336,N_5198,N_5136);
nor U5337 (N_5337,N_5028,N_5115);
nor U5338 (N_5338,N_5031,N_5036);
or U5339 (N_5339,N_5195,N_5096);
and U5340 (N_5340,N_5080,N_5079);
nor U5341 (N_5341,N_5054,N_5113);
and U5342 (N_5342,N_5142,N_5033);
and U5343 (N_5343,N_5054,N_5088);
or U5344 (N_5344,N_5171,N_5092);
xnor U5345 (N_5345,N_5134,N_5095);
nor U5346 (N_5346,N_5049,N_5020);
and U5347 (N_5347,N_5175,N_5164);
or U5348 (N_5348,N_5187,N_5022);
nor U5349 (N_5349,N_5182,N_5126);
and U5350 (N_5350,N_5038,N_5195);
nand U5351 (N_5351,N_5163,N_5050);
xor U5352 (N_5352,N_5103,N_5112);
nor U5353 (N_5353,N_5099,N_5108);
nor U5354 (N_5354,N_5134,N_5107);
nor U5355 (N_5355,N_5155,N_5028);
nand U5356 (N_5356,N_5176,N_5174);
xnor U5357 (N_5357,N_5050,N_5194);
xnor U5358 (N_5358,N_5103,N_5095);
or U5359 (N_5359,N_5122,N_5049);
or U5360 (N_5360,N_5124,N_5032);
xnor U5361 (N_5361,N_5098,N_5046);
nand U5362 (N_5362,N_5194,N_5100);
nand U5363 (N_5363,N_5144,N_5043);
nor U5364 (N_5364,N_5168,N_5152);
nor U5365 (N_5365,N_5106,N_5034);
or U5366 (N_5366,N_5140,N_5133);
and U5367 (N_5367,N_5029,N_5161);
nor U5368 (N_5368,N_5056,N_5079);
or U5369 (N_5369,N_5155,N_5187);
xnor U5370 (N_5370,N_5063,N_5011);
xor U5371 (N_5371,N_5118,N_5027);
nand U5372 (N_5372,N_5076,N_5139);
nand U5373 (N_5373,N_5137,N_5078);
nand U5374 (N_5374,N_5018,N_5023);
or U5375 (N_5375,N_5114,N_5089);
nand U5376 (N_5376,N_5155,N_5077);
nand U5377 (N_5377,N_5192,N_5098);
nand U5378 (N_5378,N_5196,N_5197);
or U5379 (N_5379,N_5032,N_5031);
nand U5380 (N_5380,N_5176,N_5091);
or U5381 (N_5381,N_5134,N_5074);
nor U5382 (N_5382,N_5070,N_5192);
xnor U5383 (N_5383,N_5184,N_5063);
or U5384 (N_5384,N_5107,N_5062);
nand U5385 (N_5385,N_5109,N_5194);
or U5386 (N_5386,N_5083,N_5092);
xor U5387 (N_5387,N_5142,N_5133);
nor U5388 (N_5388,N_5077,N_5094);
nor U5389 (N_5389,N_5013,N_5072);
nor U5390 (N_5390,N_5061,N_5120);
xnor U5391 (N_5391,N_5180,N_5026);
nand U5392 (N_5392,N_5171,N_5161);
and U5393 (N_5393,N_5155,N_5007);
xor U5394 (N_5394,N_5185,N_5053);
and U5395 (N_5395,N_5128,N_5174);
and U5396 (N_5396,N_5181,N_5099);
and U5397 (N_5397,N_5074,N_5136);
nand U5398 (N_5398,N_5031,N_5055);
nor U5399 (N_5399,N_5084,N_5059);
and U5400 (N_5400,N_5278,N_5311);
nand U5401 (N_5401,N_5378,N_5265);
or U5402 (N_5402,N_5395,N_5248);
nand U5403 (N_5403,N_5244,N_5290);
nor U5404 (N_5404,N_5221,N_5299);
nor U5405 (N_5405,N_5200,N_5391);
and U5406 (N_5406,N_5230,N_5225);
and U5407 (N_5407,N_5243,N_5317);
xnor U5408 (N_5408,N_5306,N_5328);
xor U5409 (N_5409,N_5284,N_5319);
or U5410 (N_5410,N_5301,N_5274);
and U5411 (N_5411,N_5213,N_5307);
and U5412 (N_5412,N_5294,N_5336);
nor U5413 (N_5413,N_5340,N_5305);
and U5414 (N_5414,N_5330,N_5285);
nand U5415 (N_5415,N_5335,N_5296);
nand U5416 (N_5416,N_5329,N_5254);
or U5417 (N_5417,N_5323,N_5333);
and U5418 (N_5418,N_5316,N_5308);
or U5419 (N_5419,N_5262,N_5269);
or U5420 (N_5420,N_5348,N_5232);
nor U5421 (N_5421,N_5390,N_5292);
and U5422 (N_5422,N_5233,N_5372);
nor U5423 (N_5423,N_5327,N_5315);
and U5424 (N_5424,N_5347,N_5281);
xnor U5425 (N_5425,N_5320,N_5326);
nor U5426 (N_5426,N_5396,N_5277);
and U5427 (N_5427,N_5272,N_5208);
xnor U5428 (N_5428,N_5246,N_5321);
nand U5429 (N_5429,N_5352,N_5354);
nand U5430 (N_5430,N_5385,N_5288);
nor U5431 (N_5431,N_5291,N_5268);
nand U5432 (N_5432,N_5392,N_5236);
xnor U5433 (N_5433,N_5356,N_5267);
nand U5434 (N_5434,N_5374,N_5367);
or U5435 (N_5435,N_5271,N_5252);
xor U5436 (N_5436,N_5393,N_5295);
nor U5437 (N_5437,N_5217,N_5371);
nor U5438 (N_5438,N_5261,N_5234);
or U5439 (N_5439,N_5364,N_5344);
nor U5440 (N_5440,N_5249,N_5359);
and U5441 (N_5441,N_5388,N_5245);
nand U5442 (N_5442,N_5280,N_5331);
and U5443 (N_5443,N_5239,N_5383);
xnor U5444 (N_5444,N_5216,N_5273);
and U5445 (N_5445,N_5286,N_5343);
and U5446 (N_5446,N_5210,N_5287);
nor U5447 (N_5447,N_5357,N_5253);
nor U5448 (N_5448,N_5386,N_5341);
xor U5449 (N_5449,N_5302,N_5309);
xor U5450 (N_5450,N_5209,N_5384);
nand U5451 (N_5451,N_5237,N_5358);
or U5452 (N_5452,N_5322,N_5223);
xor U5453 (N_5453,N_5238,N_5227);
xor U5454 (N_5454,N_5334,N_5289);
nor U5455 (N_5455,N_5264,N_5338);
and U5456 (N_5456,N_5382,N_5314);
and U5457 (N_5457,N_5211,N_5279);
and U5458 (N_5458,N_5380,N_5270);
xnor U5459 (N_5459,N_5318,N_5398);
xnor U5460 (N_5460,N_5298,N_5250);
nand U5461 (N_5461,N_5205,N_5263);
xnor U5462 (N_5462,N_5282,N_5214);
xnor U5463 (N_5463,N_5399,N_5207);
nand U5464 (N_5464,N_5342,N_5370);
nand U5465 (N_5465,N_5215,N_5375);
xor U5466 (N_5466,N_5293,N_5355);
or U5467 (N_5467,N_5349,N_5247);
and U5468 (N_5468,N_5297,N_5346);
or U5469 (N_5469,N_5257,N_5310);
nor U5470 (N_5470,N_5381,N_5276);
and U5471 (N_5471,N_5377,N_5373);
nor U5472 (N_5472,N_5397,N_5332);
or U5473 (N_5473,N_5219,N_5231);
xnor U5474 (N_5474,N_5212,N_5304);
and U5475 (N_5475,N_5255,N_5260);
nand U5476 (N_5476,N_5361,N_5353);
nor U5477 (N_5477,N_5206,N_5222);
nor U5478 (N_5478,N_5379,N_5368);
nand U5479 (N_5479,N_5394,N_5365);
and U5480 (N_5480,N_5362,N_5345);
or U5481 (N_5481,N_5240,N_5337);
nand U5482 (N_5482,N_5303,N_5203);
nand U5483 (N_5483,N_5259,N_5324);
nor U5484 (N_5484,N_5275,N_5283);
nor U5485 (N_5485,N_5325,N_5226);
nand U5486 (N_5486,N_5300,N_5313);
or U5487 (N_5487,N_5224,N_5266);
or U5488 (N_5488,N_5229,N_5376);
xor U5489 (N_5489,N_5369,N_5350);
and U5490 (N_5490,N_5312,N_5251);
xor U5491 (N_5491,N_5360,N_5387);
xnor U5492 (N_5492,N_5351,N_5202);
or U5493 (N_5493,N_5220,N_5339);
and U5494 (N_5494,N_5242,N_5389);
and U5495 (N_5495,N_5241,N_5256);
or U5496 (N_5496,N_5201,N_5218);
and U5497 (N_5497,N_5366,N_5363);
and U5498 (N_5498,N_5235,N_5204);
or U5499 (N_5499,N_5258,N_5228);
or U5500 (N_5500,N_5290,N_5282);
nor U5501 (N_5501,N_5326,N_5259);
and U5502 (N_5502,N_5262,N_5319);
xor U5503 (N_5503,N_5312,N_5362);
xnor U5504 (N_5504,N_5341,N_5297);
nor U5505 (N_5505,N_5366,N_5330);
and U5506 (N_5506,N_5200,N_5303);
or U5507 (N_5507,N_5384,N_5227);
xnor U5508 (N_5508,N_5259,N_5303);
nor U5509 (N_5509,N_5224,N_5260);
and U5510 (N_5510,N_5366,N_5365);
and U5511 (N_5511,N_5229,N_5282);
nand U5512 (N_5512,N_5356,N_5293);
and U5513 (N_5513,N_5252,N_5202);
nand U5514 (N_5514,N_5277,N_5322);
or U5515 (N_5515,N_5241,N_5230);
nand U5516 (N_5516,N_5381,N_5350);
nor U5517 (N_5517,N_5270,N_5225);
nor U5518 (N_5518,N_5280,N_5391);
nand U5519 (N_5519,N_5333,N_5220);
and U5520 (N_5520,N_5317,N_5301);
xnor U5521 (N_5521,N_5330,N_5214);
xor U5522 (N_5522,N_5231,N_5310);
and U5523 (N_5523,N_5257,N_5216);
nand U5524 (N_5524,N_5259,N_5390);
or U5525 (N_5525,N_5252,N_5211);
xor U5526 (N_5526,N_5235,N_5245);
xor U5527 (N_5527,N_5217,N_5242);
xor U5528 (N_5528,N_5390,N_5341);
xnor U5529 (N_5529,N_5214,N_5363);
or U5530 (N_5530,N_5268,N_5305);
or U5531 (N_5531,N_5315,N_5316);
or U5532 (N_5532,N_5228,N_5324);
and U5533 (N_5533,N_5219,N_5241);
or U5534 (N_5534,N_5308,N_5298);
nor U5535 (N_5535,N_5334,N_5304);
nor U5536 (N_5536,N_5310,N_5283);
and U5537 (N_5537,N_5362,N_5352);
nand U5538 (N_5538,N_5367,N_5383);
and U5539 (N_5539,N_5224,N_5324);
or U5540 (N_5540,N_5258,N_5213);
xnor U5541 (N_5541,N_5332,N_5231);
nand U5542 (N_5542,N_5345,N_5249);
xnor U5543 (N_5543,N_5248,N_5388);
and U5544 (N_5544,N_5306,N_5286);
and U5545 (N_5545,N_5306,N_5283);
or U5546 (N_5546,N_5360,N_5319);
or U5547 (N_5547,N_5290,N_5287);
nor U5548 (N_5548,N_5242,N_5210);
and U5549 (N_5549,N_5364,N_5375);
or U5550 (N_5550,N_5353,N_5309);
xnor U5551 (N_5551,N_5289,N_5236);
or U5552 (N_5552,N_5290,N_5360);
nor U5553 (N_5553,N_5376,N_5285);
nand U5554 (N_5554,N_5300,N_5223);
xnor U5555 (N_5555,N_5266,N_5371);
nor U5556 (N_5556,N_5295,N_5325);
nand U5557 (N_5557,N_5345,N_5208);
or U5558 (N_5558,N_5352,N_5232);
and U5559 (N_5559,N_5248,N_5268);
and U5560 (N_5560,N_5347,N_5300);
xor U5561 (N_5561,N_5249,N_5382);
or U5562 (N_5562,N_5225,N_5291);
or U5563 (N_5563,N_5320,N_5374);
nor U5564 (N_5564,N_5304,N_5341);
and U5565 (N_5565,N_5357,N_5384);
and U5566 (N_5566,N_5269,N_5305);
and U5567 (N_5567,N_5318,N_5228);
nand U5568 (N_5568,N_5362,N_5276);
nand U5569 (N_5569,N_5326,N_5335);
nand U5570 (N_5570,N_5267,N_5260);
or U5571 (N_5571,N_5257,N_5344);
and U5572 (N_5572,N_5250,N_5345);
and U5573 (N_5573,N_5348,N_5268);
xor U5574 (N_5574,N_5210,N_5224);
or U5575 (N_5575,N_5205,N_5399);
xor U5576 (N_5576,N_5350,N_5297);
nand U5577 (N_5577,N_5261,N_5394);
or U5578 (N_5578,N_5310,N_5208);
or U5579 (N_5579,N_5280,N_5381);
nor U5580 (N_5580,N_5234,N_5368);
xnor U5581 (N_5581,N_5387,N_5344);
xor U5582 (N_5582,N_5269,N_5304);
nor U5583 (N_5583,N_5372,N_5218);
nor U5584 (N_5584,N_5307,N_5211);
xnor U5585 (N_5585,N_5272,N_5397);
or U5586 (N_5586,N_5363,N_5208);
xor U5587 (N_5587,N_5368,N_5236);
xnor U5588 (N_5588,N_5354,N_5263);
nand U5589 (N_5589,N_5329,N_5311);
and U5590 (N_5590,N_5231,N_5243);
xor U5591 (N_5591,N_5347,N_5255);
and U5592 (N_5592,N_5363,N_5267);
or U5593 (N_5593,N_5362,N_5231);
and U5594 (N_5594,N_5331,N_5390);
or U5595 (N_5595,N_5307,N_5357);
nor U5596 (N_5596,N_5281,N_5374);
or U5597 (N_5597,N_5324,N_5342);
or U5598 (N_5598,N_5383,N_5238);
xor U5599 (N_5599,N_5252,N_5317);
nor U5600 (N_5600,N_5525,N_5537);
and U5601 (N_5601,N_5572,N_5538);
and U5602 (N_5602,N_5509,N_5407);
and U5603 (N_5603,N_5520,N_5585);
nor U5604 (N_5604,N_5469,N_5547);
and U5605 (N_5605,N_5405,N_5511);
nor U5606 (N_5606,N_5458,N_5505);
nor U5607 (N_5607,N_5557,N_5527);
nor U5608 (N_5608,N_5597,N_5488);
nand U5609 (N_5609,N_5522,N_5559);
nor U5610 (N_5610,N_5516,N_5549);
or U5611 (N_5611,N_5579,N_5513);
nor U5612 (N_5612,N_5453,N_5420);
or U5613 (N_5613,N_5497,N_5440);
or U5614 (N_5614,N_5482,N_5580);
xnor U5615 (N_5615,N_5462,N_5571);
or U5616 (N_5616,N_5536,N_5587);
or U5617 (N_5617,N_5493,N_5445);
nor U5618 (N_5618,N_5530,N_5539);
or U5619 (N_5619,N_5401,N_5568);
and U5620 (N_5620,N_5491,N_5551);
xnor U5621 (N_5621,N_5564,N_5582);
xnor U5622 (N_5622,N_5577,N_5442);
xor U5623 (N_5623,N_5499,N_5455);
nor U5624 (N_5624,N_5415,N_5583);
or U5625 (N_5625,N_5463,N_5428);
or U5626 (N_5626,N_5502,N_5535);
nand U5627 (N_5627,N_5555,N_5431);
and U5628 (N_5628,N_5457,N_5473);
xnor U5629 (N_5629,N_5487,N_5529);
xor U5630 (N_5630,N_5599,N_5427);
or U5631 (N_5631,N_5452,N_5596);
and U5632 (N_5632,N_5561,N_5588);
nand U5633 (N_5633,N_5432,N_5546);
and U5634 (N_5634,N_5436,N_5531);
nor U5635 (N_5635,N_5425,N_5517);
and U5636 (N_5636,N_5408,N_5454);
xnor U5637 (N_5637,N_5423,N_5501);
xor U5638 (N_5638,N_5434,N_5451);
xor U5639 (N_5639,N_5567,N_5576);
and U5640 (N_5640,N_5406,N_5475);
nand U5641 (N_5641,N_5515,N_5532);
xnor U5642 (N_5642,N_5592,N_5574);
nor U5643 (N_5643,N_5562,N_5595);
nand U5644 (N_5644,N_5543,N_5590);
nand U5645 (N_5645,N_5569,N_5550);
xor U5646 (N_5646,N_5429,N_5483);
or U5647 (N_5647,N_5554,N_5495);
nor U5648 (N_5648,N_5476,N_5477);
nor U5649 (N_5649,N_5500,N_5447);
nor U5650 (N_5650,N_5533,N_5479);
and U5651 (N_5651,N_5553,N_5410);
nand U5652 (N_5652,N_5417,N_5506);
nor U5653 (N_5653,N_5426,N_5402);
nor U5654 (N_5654,N_5421,N_5466);
and U5655 (N_5655,N_5548,N_5518);
nor U5656 (N_5656,N_5578,N_5474);
and U5657 (N_5657,N_5558,N_5514);
or U5658 (N_5658,N_5540,N_5492);
and U5659 (N_5659,N_5461,N_5504);
xor U5660 (N_5660,N_5521,N_5486);
and U5661 (N_5661,N_5416,N_5419);
nand U5662 (N_5662,N_5494,N_5409);
xnor U5663 (N_5663,N_5480,N_5435);
and U5664 (N_5664,N_5570,N_5565);
or U5665 (N_5665,N_5484,N_5575);
xor U5666 (N_5666,N_5534,N_5446);
xnor U5667 (N_5667,N_5441,N_5544);
nor U5668 (N_5668,N_5508,N_5526);
xor U5669 (N_5669,N_5418,N_5528);
and U5670 (N_5670,N_5470,N_5519);
nor U5671 (N_5671,N_5591,N_5560);
and U5672 (N_5672,N_5507,N_5566);
or U5673 (N_5673,N_5456,N_5545);
nor U5674 (N_5674,N_5598,N_5437);
and U5675 (N_5675,N_5496,N_5552);
nor U5676 (N_5676,N_5510,N_5478);
xnor U5677 (N_5677,N_5584,N_5589);
xor U5678 (N_5678,N_5443,N_5424);
or U5679 (N_5679,N_5503,N_5464);
and U5680 (N_5680,N_5444,N_5400);
nand U5681 (N_5681,N_5524,N_5413);
and U5682 (N_5682,N_5485,N_5563);
or U5683 (N_5683,N_5422,N_5448);
and U5684 (N_5684,N_5586,N_5512);
xor U5685 (N_5685,N_5593,N_5472);
or U5686 (N_5686,N_5541,N_5460);
or U5687 (N_5687,N_5481,N_5542);
nand U5688 (N_5688,N_5414,N_5412);
nor U5689 (N_5689,N_5411,N_5556);
nor U5690 (N_5690,N_5489,N_5449);
or U5691 (N_5691,N_5450,N_5573);
nand U5692 (N_5692,N_5430,N_5468);
and U5693 (N_5693,N_5459,N_5498);
nand U5694 (N_5694,N_5433,N_5439);
xor U5695 (N_5695,N_5465,N_5581);
or U5696 (N_5696,N_5594,N_5403);
or U5697 (N_5697,N_5490,N_5438);
and U5698 (N_5698,N_5404,N_5467);
xor U5699 (N_5699,N_5471,N_5523);
and U5700 (N_5700,N_5499,N_5472);
nor U5701 (N_5701,N_5418,N_5431);
or U5702 (N_5702,N_5536,N_5501);
nor U5703 (N_5703,N_5522,N_5568);
xor U5704 (N_5704,N_5515,N_5446);
or U5705 (N_5705,N_5464,N_5525);
and U5706 (N_5706,N_5585,N_5546);
nor U5707 (N_5707,N_5502,N_5446);
and U5708 (N_5708,N_5444,N_5573);
nand U5709 (N_5709,N_5495,N_5586);
or U5710 (N_5710,N_5561,N_5495);
xor U5711 (N_5711,N_5549,N_5412);
and U5712 (N_5712,N_5402,N_5596);
and U5713 (N_5713,N_5469,N_5483);
or U5714 (N_5714,N_5420,N_5427);
or U5715 (N_5715,N_5531,N_5490);
nor U5716 (N_5716,N_5543,N_5514);
nand U5717 (N_5717,N_5412,N_5542);
or U5718 (N_5718,N_5450,N_5467);
or U5719 (N_5719,N_5538,N_5445);
nor U5720 (N_5720,N_5598,N_5587);
and U5721 (N_5721,N_5517,N_5541);
xnor U5722 (N_5722,N_5441,N_5522);
nand U5723 (N_5723,N_5453,N_5480);
nand U5724 (N_5724,N_5548,N_5551);
xnor U5725 (N_5725,N_5584,N_5437);
nand U5726 (N_5726,N_5405,N_5512);
xor U5727 (N_5727,N_5505,N_5592);
nand U5728 (N_5728,N_5541,N_5454);
xnor U5729 (N_5729,N_5552,N_5443);
and U5730 (N_5730,N_5439,N_5577);
nor U5731 (N_5731,N_5449,N_5589);
nand U5732 (N_5732,N_5485,N_5568);
or U5733 (N_5733,N_5468,N_5475);
nor U5734 (N_5734,N_5527,N_5525);
xor U5735 (N_5735,N_5499,N_5427);
xnor U5736 (N_5736,N_5412,N_5570);
and U5737 (N_5737,N_5445,N_5570);
or U5738 (N_5738,N_5404,N_5457);
and U5739 (N_5739,N_5401,N_5558);
and U5740 (N_5740,N_5590,N_5421);
nand U5741 (N_5741,N_5590,N_5497);
and U5742 (N_5742,N_5407,N_5519);
or U5743 (N_5743,N_5470,N_5558);
nand U5744 (N_5744,N_5539,N_5512);
and U5745 (N_5745,N_5580,N_5408);
nand U5746 (N_5746,N_5449,N_5402);
or U5747 (N_5747,N_5489,N_5429);
nor U5748 (N_5748,N_5539,N_5481);
or U5749 (N_5749,N_5513,N_5554);
nand U5750 (N_5750,N_5550,N_5531);
or U5751 (N_5751,N_5596,N_5474);
and U5752 (N_5752,N_5510,N_5472);
nand U5753 (N_5753,N_5424,N_5434);
nor U5754 (N_5754,N_5451,N_5509);
or U5755 (N_5755,N_5412,N_5474);
nand U5756 (N_5756,N_5581,N_5570);
xnor U5757 (N_5757,N_5531,N_5455);
xor U5758 (N_5758,N_5433,N_5455);
nand U5759 (N_5759,N_5506,N_5567);
or U5760 (N_5760,N_5472,N_5571);
xor U5761 (N_5761,N_5518,N_5436);
xnor U5762 (N_5762,N_5413,N_5487);
nand U5763 (N_5763,N_5476,N_5581);
nand U5764 (N_5764,N_5581,N_5530);
or U5765 (N_5765,N_5482,N_5503);
xnor U5766 (N_5766,N_5547,N_5468);
and U5767 (N_5767,N_5401,N_5490);
or U5768 (N_5768,N_5571,N_5579);
or U5769 (N_5769,N_5445,N_5532);
or U5770 (N_5770,N_5520,N_5408);
and U5771 (N_5771,N_5508,N_5468);
xnor U5772 (N_5772,N_5490,N_5585);
nand U5773 (N_5773,N_5541,N_5425);
nand U5774 (N_5774,N_5452,N_5568);
nand U5775 (N_5775,N_5453,N_5582);
and U5776 (N_5776,N_5438,N_5479);
nor U5777 (N_5777,N_5401,N_5592);
nor U5778 (N_5778,N_5427,N_5482);
and U5779 (N_5779,N_5549,N_5430);
or U5780 (N_5780,N_5536,N_5510);
nor U5781 (N_5781,N_5462,N_5543);
xnor U5782 (N_5782,N_5404,N_5518);
nor U5783 (N_5783,N_5536,N_5406);
nor U5784 (N_5784,N_5574,N_5416);
and U5785 (N_5785,N_5534,N_5417);
nor U5786 (N_5786,N_5539,N_5533);
nor U5787 (N_5787,N_5520,N_5575);
xnor U5788 (N_5788,N_5451,N_5475);
xnor U5789 (N_5789,N_5491,N_5472);
and U5790 (N_5790,N_5576,N_5409);
nor U5791 (N_5791,N_5472,N_5446);
nor U5792 (N_5792,N_5573,N_5454);
xor U5793 (N_5793,N_5560,N_5598);
xnor U5794 (N_5794,N_5571,N_5413);
nor U5795 (N_5795,N_5541,N_5405);
xor U5796 (N_5796,N_5400,N_5475);
nor U5797 (N_5797,N_5495,N_5510);
nor U5798 (N_5798,N_5540,N_5471);
and U5799 (N_5799,N_5594,N_5569);
nor U5800 (N_5800,N_5665,N_5618);
xnor U5801 (N_5801,N_5641,N_5722);
nor U5802 (N_5802,N_5706,N_5727);
nor U5803 (N_5803,N_5602,N_5749);
nand U5804 (N_5804,N_5607,N_5707);
and U5805 (N_5805,N_5685,N_5745);
xor U5806 (N_5806,N_5776,N_5697);
and U5807 (N_5807,N_5659,N_5767);
or U5808 (N_5808,N_5628,N_5717);
nand U5809 (N_5809,N_5627,N_5703);
nor U5810 (N_5810,N_5636,N_5721);
nand U5811 (N_5811,N_5712,N_5638);
xor U5812 (N_5812,N_5662,N_5605);
xnor U5813 (N_5813,N_5741,N_5770);
or U5814 (N_5814,N_5698,N_5666);
xor U5815 (N_5815,N_5624,N_5787);
nand U5816 (N_5816,N_5780,N_5623);
or U5817 (N_5817,N_5789,N_5732);
and U5818 (N_5818,N_5630,N_5629);
and U5819 (N_5819,N_5664,N_5743);
or U5820 (N_5820,N_5614,N_5740);
xnor U5821 (N_5821,N_5700,N_5634);
and U5822 (N_5822,N_5615,N_5736);
xnor U5823 (N_5823,N_5635,N_5731);
or U5824 (N_5824,N_5796,N_5788);
nand U5825 (N_5825,N_5699,N_5794);
nor U5826 (N_5826,N_5739,N_5651);
xnor U5827 (N_5827,N_5750,N_5642);
nand U5828 (N_5828,N_5755,N_5723);
nand U5829 (N_5829,N_5715,N_5693);
nand U5830 (N_5830,N_5619,N_5751);
nand U5831 (N_5831,N_5729,N_5649);
xor U5832 (N_5832,N_5674,N_5654);
nor U5833 (N_5833,N_5771,N_5719);
or U5834 (N_5834,N_5669,N_5673);
nor U5835 (N_5835,N_5668,N_5686);
nor U5836 (N_5836,N_5606,N_5670);
xor U5837 (N_5837,N_5769,N_5784);
xor U5838 (N_5838,N_5678,N_5768);
xor U5839 (N_5839,N_5748,N_5675);
or U5840 (N_5840,N_5701,N_5653);
xnor U5841 (N_5841,N_5765,N_5695);
and U5842 (N_5842,N_5646,N_5734);
or U5843 (N_5843,N_5785,N_5786);
or U5844 (N_5844,N_5783,N_5632);
xor U5845 (N_5845,N_5792,N_5756);
and U5846 (N_5846,N_5718,N_5775);
or U5847 (N_5847,N_5696,N_5603);
xor U5848 (N_5848,N_5793,N_5708);
nand U5849 (N_5849,N_5766,N_5680);
or U5850 (N_5850,N_5730,N_5795);
nor U5851 (N_5851,N_5791,N_5705);
nand U5852 (N_5852,N_5689,N_5681);
xor U5853 (N_5853,N_5798,N_5613);
and U5854 (N_5854,N_5759,N_5645);
or U5855 (N_5855,N_5742,N_5747);
nor U5856 (N_5856,N_5762,N_5643);
nor U5857 (N_5857,N_5640,N_5657);
xor U5858 (N_5858,N_5625,N_5671);
or U5859 (N_5859,N_5774,N_5692);
or U5860 (N_5860,N_5648,N_5622);
and U5861 (N_5861,N_5644,N_5763);
or U5862 (N_5862,N_5620,N_5611);
and U5863 (N_5863,N_5710,N_5626);
xor U5864 (N_5864,N_5728,N_5639);
and U5865 (N_5865,N_5631,N_5672);
and U5866 (N_5866,N_5650,N_5682);
nand U5867 (N_5867,N_5612,N_5746);
and U5868 (N_5868,N_5601,N_5690);
xnor U5869 (N_5869,N_5781,N_5752);
or U5870 (N_5870,N_5655,N_5663);
nand U5871 (N_5871,N_5687,N_5683);
or U5872 (N_5872,N_5617,N_5637);
or U5873 (N_5873,N_5677,N_5737);
and U5874 (N_5874,N_5757,N_5726);
and U5875 (N_5875,N_5704,N_5621);
nand U5876 (N_5876,N_5661,N_5797);
xnor U5877 (N_5877,N_5660,N_5724);
nand U5878 (N_5878,N_5760,N_5609);
nand U5879 (N_5879,N_5633,N_5773);
or U5880 (N_5880,N_5790,N_5600);
and U5881 (N_5881,N_5684,N_5725);
or U5882 (N_5882,N_5711,N_5610);
or U5883 (N_5883,N_5778,N_5604);
nand U5884 (N_5884,N_5744,N_5753);
xnor U5885 (N_5885,N_5738,N_5616);
or U5886 (N_5886,N_5716,N_5691);
or U5887 (N_5887,N_5799,N_5702);
or U5888 (N_5888,N_5782,N_5652);
or U5889 (N_5889,N_5714,N_5772);
xnor U5890 (N_5890,N_5764,N_5720);
nand U5891 (N_5891,N_5779,N_5713);
nor U5892 (N_5892,N_5709,N_5667);
or U5893 (N_5893,N_5658,N_5735);
and U5894 (N_5894,N_5733,N_5694);
or U5895 (N_5895,N_5761,N_5777);
nor U5896 (N_5896,N_5608,N_5754);
xor U5897 (N_5897,N_5688,N_5679);
and U5898 (N_5898,N_5656,N_5676);
nor U5899 (N_5899,N_5758,N_5647);
or U5900 (N_5900,N_5708,N_5737);
xnor U5901 (N_5901,N_5610,N_5797);
xnor U5902 (N_5902,N_5762,N_5777);
nand U5903 (N_5903,N_5690,N_5641);
and U5904 (N_5904,N_5770,N_5638);
nor U5905 (N_5905,N_5643,N_5612);
nor U5906 (N_5906,N_5775,N_5659);
nor U5907 (N_5907,N_5618,N_5779);
xor U5908 (N_5908,N_5750,N_5716);
nand U5909 (N_5909,N_5655,N_5621);
nor U5910 (N_5910,N_5608,N_5784);
nand U5911 (N_5911,N_5749,N_5775);
xor U5912 (N_5912,N_5691,N_5711);
or U5913 (N_5913,N_5650,N_5713);
xor U5914 (N_5914,N_5713,N_5662);
nand U5915 (N_5915,N_5740,N_5748);
xor U5916 (N_5916,N_5709,N_5768);
or U5917 (N_5917,N_5618,N_5764);
nand U5918 (N_5918,N_5773,N_5759);
xor U5919 (N_5919,N_5651,N_5634);
nand U5920 (N_5920,N_5667,N_5762);
nand U5921 (N_5921,N_5602,N_5677);
xnor U5922 (N_5922,N_5619,N_5798);
xnor U5923 (N_5923,N_5726,N_5739);
xnor U5924 (N_5924,N_5640,N_5690);
nand U5925 (N_5925,N_5651,N_5679);
nor U5926 (N_5926,N_5680,N_5720);
and U5927 (N_5927,N_5791,N_5722);
nand U5928 (N_5928,N_5730,N_5708);
xnor U5929 (N_5929,N_5732,N_5705);
and U5930 (N_5930,N_5749,N_5727);
or U5931 (N_5931,N_5611,N_5735);
nor U5932 (N_5932,N_5631,N_5696);
nand U5933 (N_5933,N_5606,N_5613);
xor U5934 (N_5934,N_5630,N_5723);
xnor U5935 (N_5935,N_5660,N_5761);
and U5936 (N_5936,N_5736,N_5781);
or U5937 (N_5937,N_5736,N_5737);
nor U5938 (N_5938,N_5748,N_5712);
nand U5939 (N_5939,N_5771,N_5779);
nor U5940 (N_5940,N_5799,N_5785);
xnor U5941 (N_5941,N_5623,N_5613);
or U5942 (N_5942,N_5610,N_5684);
xnor U5943 (N_5943,N_5720,N_5622);
or U5944 (N_5944,N_5710,N_5701);
xnor U5945 (N_5945,N_5656,N_5612);
xor U5946 (N_5946,N_5688,N_5617);
xnor U5947 (N_5947,N_5602,N_5606);
nor U5948 (N_5948,N_5716,N_5740);
nand U5949 (N_5949,N_5762,N_5670);
nand U5950 (N_5950,N_5620,N_5601);
xnor U5951 (N_5951,N_5744,N_5764);
or U5952 (N_5952,N_5684,N_5740);
nor U5953 (N_5953,N_5641,N_5654);
nand U5954 (N_5954,N_5793,N_5749);
and U5955 (N_5955,N_5773,N_5700);
or U5956 (N_5956,N_5736,N_5787);
or U5957 (N_5957,N_5637,N_5642);
and U5958 (N_5958,N_5775,N_5642);
xor U5959 (N_5959,N_5602,N_5796);
nor U5960 (N_5960,N_5664,N_5744);
nor U5961 (N_5961,N_5676,N_5637);
nand U5962 (N_5962,N_5757,N_5673);
nor U5963 (N_5963,N_5733,N_5782);
nor U5964 (N_5964,N_5670,N_5677);
or U5965 (N_5965,N_5650,N_5633);
and U5966 (N_5966,N_5725,N_5698);
nor U5967 (N_5967,N_5757,N_5689);
or U5968 (N_5968,N_5723,N_5760);
or U5969 (N_5969,N_5686,N_5697);
nand U5970 (N_5970,N_5797,N_5603);
nand U5971 (N_5971,N_5714,N_5777);
and U5972 (N_5972,N_5701,N_5753);
nand U5973 (N_5973,N_5643,N_5632);
and U5974 (N_5974,N_5771,N_5715);
or U5975 (N_5975,N_5670,N_5728);
nand U5976 (N_5976,N_5679,N_5672);
nor U5977 (N_5977,N_5696,N_5670);
and U5978 (N_5978,N_5745,N_5774);
or U5979 (N_5979,N_5778,N_5795);
xnor U5980 (N_5980,N_5733,N_5637);
xnor U5981 (N_5981,N_5611,N_5694);
nor U5982 (N_5982,N_5645,N_5621);
nand U5983 (N_5983,N_5612,N_5715);
and U5984 (N_5984,N_5684,N_5653);
nor U5985 (N_5985,N_5648,N_5647);
or U5986 (N_5986,N_5716,N_5720);
nor U5987 (N_5987,N_5705,N_5707);
xor U5988 (N_5988,N_5652,N_5710);
xnor U5989 (N_5989,N_5740,N_5746);
or U5990 (N_5990,N_5710,N_5607);
and U5991 (N_5991,N_5769,N_5655);
xnor U5992 (N_5992,N_5680,N_5731);
and U5993 (N_5993,N_5689,N_5772);
xnor U5994 (N_5994,N_5615,N_5773);
nor U5995 (N_5995,N_5730,N_5661);
xnor U5996 (N_5996,N_5796,N_5607);
nor U5997 (N_5997,N_5729,N_5685);
xor U5998 (N_5998,N_5656,N_5708);
nand U5999 (N_5999,N_5745,N_5647);
nor U6000 (N_6000,N_5910,N_5982);
or U6001 (N_6001,N_5839,N_5845);
nand U6002 (N_6002,N_5899,N_5961);
or U6003 (N_6003,N_5846,N_5983);
xnor U6004 (N_6004,N_5953,N_5804);
nor U6005 (N_6005,N_5944,N_5822);
nand U6006 (N_6006,N_5969,N_5968);
and U6007 (N_6007,N_5924,N_5902);
nor U6008 (N_6008,N_5891,N_5909);
and U6009 (N_6009,N_5841,N_5932);
and U6010 (N_6010,N_5927,N_5896);
and U6011 (N_6011,N_5866,N_5959);
nor U6012 (N_6012,N_5869,N_5936);
xor U6013 (N_6013,N_5859,N_5990);
nor U6014 (N_6014,N_5939,N_5883);
nand U6015 (N_6015,N_5905,N_5963);
nor U6016 (N_6016,N_5817,N_5865);
nand U6017 (N_6017,N_5997,N_5907);
xor U6018 (N_6018,N_5950,N_5964);
and U6019 (N_6019,N_5832,N_5831);
or U6020 (N_6020,N_5986,N_5917);
and U6021 (N_6021,N_5818,N_5823);
nor U6022 (N_6022,N_5914,N_5943);
xnor U6023 (N_6023,N_5854,N_5908);
and U6024 (N_6024,N_5806,N_5807);
xnor U6025 (N_6025,N_5826,N_5858);
nand U6026 (N_6026,N_5893,N_5989);
or U6027 (N_6027,N_5918,N_5894);
nand U6028 (N_6028,N_5829,N_5887);
nor U6029 (N_6029,N_5980,N_5864);
or U6030 (N_6030,N_5835,N_5849);
nand U6031 (N_6031,N_5809,N_5985);
xor U6032 (N_6032,N_5926,N_5922);
and U6033 (N_6033,N_5940,N_5840);
or U6034 (N_6034,N_5844,N_5971);
or U6035 (N_6035,N_5906,N_5856);
xor U6036 (N_6036,N_5888,N_5930);
and U6037 (N_6037,N_5923,N_5945);
xnor U6038 (N_6038,N_5904,N_5988);
xnor U6039 (N_6039,N_5855,N_5947);
and U6040 (N_6040,N_5946,N_5848);
nor U6041 (N_6041,N_5890,N_5975);
xnor U6042 (N_6042,N_5973,N_5895);
nor U6043 (N_6043,N_5929,N_5955);
and U6044 (N_6044,N_5937,N_5995);
or U6045 (N_6045,N_5814,N_5802);
nor U6046 (N_6046,N_5819,N_5903);
xor U6047 (N_6047,N_5898,N_5965);
xor U6048 (N_6048,N_5877,N_5957);
or U6049 (N_6049,N_5879,N_5885);
nor U6050 (N_6050,N_5816,N_5941);
nand U6051 (N_6051,N_5842,N_5827);
xnor U6052 (N_6052,N_5825,N_5970);
xnor U6053 (N_6053,N_5960,N_5886);
nand U6054 (N_6054,N_5884,N_5935);
or U6055 (N_6055,N_5913,N_5892);
nand U6056 (N_6056,N_5801,N_5824);
xor U6057 (N_6057,N_5833,N_5836);
nor U6058 (N_6058,N_5921,N_5808);
or U6059 (N_6059,N_5919,N_5984);
xor U6060 (N_6060,N_5838,N_5862);
and U6061 (N_6061,N_5981,N_5911);
and U6062 (N_6062,N_5948,N_5897);
nor U6063 (N_6063,N_5872,N_5870);
or U6064 (N_6064,N_5912,N_5942);
and U6065 (N_6065,N_5812,N_5954);
nor U6066 (N_6066,N_5811,N_5852);
nor U6067 (N_6067,N_5999,N_5815);
nand U6068 (N_6068,N_5876,N_5925);
or U6069 (N_6069,N_5998,N_5837);
or U6070 (N_6070,N_5851,N_5979);
and U6071 (N_6071,N_5933,N_5882);
or U6072 (N_6072,N_5900,N_5991);
xnor U6073 (N_6073,N_5915,N_5949);
nor U6074 (N_6074,N_5976,N_5920);
or U6075 (N_6075,N_5861,N_5987);
xor U6076 (N_6076,N_5934,N_5850);
or U6077 (N_6077,N_5938,N_5805);
and U6078 (N_6078,N_5810,N_5871);
nor U6079 (N_6079,N_5928,N_5868);
nand U6080 (N_6080,N_5974,N_5873);
nor U6081 (N_6081,N_5951,N_5875);
xnor U6082 (N_6082,N_5843,N_5931);
xor U6083 (N_6083,N_5901,N_5853);
xnor U6084 (N_6084,N_5800,N_5972);
xnor U6085 (N_6085,N_5803,N_5958);
nand U6086 (N_6086,N_5828,N_5830);
nand U6087 (N_6087,N_5857,N_5874);
nor U6088 (N_6088,N_5977,N_5978);
nor U6089 (N_6089,N_5889,N_5863);
nand U6090 (N_6090,N_5962,N_5821);
xnor U6091 (N_6091,N_5993,N_5952);
nor U6092 (N_6092,N_5916,N_5860);
xnor U6093 (N_6093,N_5878,N_5994);
nor U6094 (N_6094,N_5966,N_5834);
nor U6095 (N_6095,N_5813,N_5847);
nand U6096 (N_6096,N_5880,N_5992);
xor U6097 (N_6097,N_5820,N_5996);
nor U6098 (N_6098,N_5881,N_5967);
and U6099 (N_6099,N_5867,N_5956);
xor U6100 (N_6100,N_5924,N_5928);
nor U6101 (N_6101,N_5919,N_5873);
and U6102 (N_6102,N_5910,N_5992);
or U6103 (N_6103,N_5859,N_5995);
xnor U6104 (N_6104,N_5981,N_5893);
xnor U6105 (N_6105,N_5942,N_5974);
and U6106 (N_6106,N_5847,N_5956);
and U6107 (N_6107,N_5867,N_5810);
xnor U6108 (N_6108,N_5995,N_5820);
xor U6109 (N_6109,N_5862,N_5905);
or U6110 (N_6110,N_5929,N_5846);
xnor U6111 (N_6111,N_5982,N_5953);
nand U6112 (N_6112,N_5898,N_5877);
xnor U6113 (N_6113,N_5828,N_5898);
xnor U6114 (N_6114,N_5870,N_5808);
and U6115 (N_6115,N_5971,N_5960);
or U6116 (N_6116,N_5999,N_5821);
and U6117 (N_6117,N_5931,N_5848);
nand U6118 (N_6118,N_5943,N_5827);
nand U6119 (N_6119,N_5963,N_5844);
nand U6120 (N_6120,N_5959,N_5998);
nor U6121 (N_6121,N_5906,N_5899);
nor U6122 (N_6122,N_5835,N_5983);
xor U6123 (N_6123,N_5846,N_5976);
nand U6124 (N_6124,N_5872,N_5990);
nor U6125 (N_6125,N_5896,N_5925);
or U6126 (N_6126,N_5954,N_5801);
nand U6127 (N_6127,N_5900,N_5948);
nor U6128 (N_6128,N_5972,N_5810);
nor U6129 (N_6129,N_5953,N_5889);
and U6130 (N_6130,N_5800,N_5946);
xor U6131 (N_6131,N_5980,N_5939);
and U6132 (N_6132,N_5834,N_5976);
or U6133 (N_6133,N_5890,N_5969);
nand U6134 (N_6134,N_5839,N_5997);
nor U6135 (N_6135,N_5834,N_5913);
and U6136 (N_6136,N_5847,N_5900);
xor U6137 (N_6137,N_5839,N_5849);
nor U6138 (N_6138,N_5994,N_5918);
and U6139 (N_6139,N_5957,N_5838);
xor U6140 (N_6140,N_5908,N_5832);
or U6141 (N_6141,N_5824,N_5896);
nor U6142 (N_6142,N_5857,N_5910);
or U6143 (N_6143,N_5911,N_5978);
or U6144 (N_6144,N_5931,N_5896);
nand U6145 (N_6145,N_5906,N_5959);
nand U6146 (N_6146,N_5891,N_5835);
or U6147 (N_6147,N_5909,N_5899);
nor U6148 (N_6148,N_5924,N_5931);
xnor U6149 (N_6149,N_5800,N_5892);
and U6150 (N_6150,N_5884,N_5850);
nand U6151 (N_6151,N_5893,N_5975);
nor U6152 (N_6152,N_5901,N_5997);
nor U6153 (N_6153,N_5846,N_5916);
nor U6154 (N_6154,N_5917,N_5823);
nand U6155 (N_6155,N_5998,N_5896);
or U6156 (N_6156,N_5944,N_5847);
or U6157 (N_6157,N_5821,N_5862);
nor U6158 (N_6158,N_5940,N_5886);
or U6159 (N_6159,N_5957,N_5923);
or U6160 (N_6160,N_5913,N_5947);
nor U6161 (N_6161,N_5998,N_5973);
xor U6162 (N_6162,N_5929,N_5996);
nor U6163 (N_6163,N_5944,N_5851);
and U6164 (N_6164,N_5920,N_5977);
xor U6165 (N_6165,N_5967,N_5812);
nand U6166 (N_6166,N_5831,N_5934);
nand U6167 (N_6167,N_5829,N_5833);
and U6168 (N_6168,N_5843,N_5832);
or U6169 (N_6169,N_5815,N_5811);
or U6170 (N_6170,N_5850,N_5945);
and U6171 (N_6171,N_5840,N_5876);
and U6172 (N_6172,N_5980,N_5931);
nor U6173 (N_6173,N_5968,N_5932);
xnor U6174 (N_6174,N_5861,N_5824);
xnor U6175 (N_6175,N_5938,N_5976);
or U6176 (N_6176,N_5929,N_5979);
nor U6177 (N_6177,N_5936,N_5960);
or U6178 (N_6178,N_5839,N_5889);
nor U6179 (N_6179,N_5930,N_5886);
xnor U6180 (N_6180,N_5831,N_5996);
nand U6181 (N_6181,N_5867,N_5866);
or U6182 (N_6182,N_5847,N_5855);
and U6183 (N_6183,N_5903,N_5918);
and U6184 (N_6184,N_5877,N_5814);
and U6185 (N_6185,N_5801,N_5887);
and U6186 (N_6186,N_5891,N_5953);
nand U6187 (N_6187,N_5907,N_5995);
or U6188 (N_6188,N_5892,N_5802);
nand U6189 (N_6189,N_5928,N_5876);
and U6190 (N_6190,N_5919,N_5922);
xnor U6191 (N_6191,N_5838,N_5852);
nand U6192 (N_6192,N_5898,N_5887);
and U6193 (N_6193,N_5886,N_5961);
xor U6194 (N_6194,N_5959,N_5928);
and U6195 (N_6195,N_5897,N_5820);
nand U6196 (N_6196,N_5835,N_5805);
and U6197 (N_6197,N_5918,N_5875);
nand U6198 (N_6198,N_5984,N_5831);
xor U6199 (N_6199,N_5805,N_5909);
or U6200 (N_6200,N_6060,N_6156);
and U6201 (N_6201,N_6036,N_6034);
or U6202 (N_6202,N_6185,N_6016);
xnor U6203 (N_6203,N_6132,N_6173);
nor U6204 (N_6204,N_6138,N_6179);
and U6205 (N_6205,N_6196,N_6168);
xor U6206 (N_6206,N_6116,N_6198);
and U6207 (N_6207,N_6142,N_6133);
nand U6208 (N_6208,N_6178,N_6035);
nand U6209 (N_6209,N_6046,N_6105);
nand U6210 (N_6210,N_6021,N_6024);
nand U6211 (N_6211,N_6090,N_6051);
and U6212 (N_6212,N_6123,N_6127);
nor U6213 (N_6213,N_6159,N_6114);
xnor U6214 (N_6214,N_6120,N_6059);
or U6215 (N_6215,N_6033,N_6048);
xor U6216 (N_6216,N_6172,N_6010);
and U6217 (N_6217,N_6062,N_6137);
nor U6218 (N_6218,N_6118,N_6134);
nand U6219 (N_6219,N_6095,N_6027);
xor U6220 (N_6220,N_6191,N_6102);
or U6221 (N_6221,N_6056,N_6079);
nand U6222 (N_6222,N_6001,N_6160);
and U6223 (N_6223,N_6157,N_6042);
or U6224 (N_6224,N_6111,N_6082);
xor U6225 (N_6225,N_6012,N_6065);
and U6226 (N_6226,N_6002,N_6125);
nand U6227 (N_6227,N_6041,N_6075);
nand U6228 (N_6228,N_6195,N_6014);
xor U6229 (N_6229,N_6091,N_6040);
or U6230 (N_6230,N_6175,N_6136);
and U6231 (N_6231,N_6007,N_6163);
and U6232 (N_6232,N_6152,N_6167);
or U6233 (N_6233,N_6084,N_6081);
or U6234 (N_6234,N_6140,N_6004);
and U6235 (N_6235,N_6199,N_6028);
nor U6236 (N_6236,N_6061,N_6052);
xor U6237 (N_6237,N_6192,N_6100);
nor U6238 (N_6238,N_6078,N_6176);
nand U6239 (N_6239,N_6110,N_6113);
nor U6240 (N_6240,N_6135,N_6130);
nand U6241 (N_6241,N_6047,N_6031);
nor U6242 (N_6242,N_6023,N_6005);
nand U6243 (N_6243,N_6018,N_6072);
xnor U6244 (N_6244,N_6112,N_6000);
nor U6245 (N_6245,N_6089,N_6043);
and U6246 (N_6246,N_6182,N_6129);
nand U6247 (N_6247,N_6143,N_6187);
or U6248 (N_6248,N_6154,N_6166);
nor U6249 (N_6249,N_6099,N_6026);
or U6250 (N_6250,N_6038,N_6170);
xor U6251 (N_6251,N_6063,N_6119);
nand U6252 (N_6252,N_6126,N_6069);
xnor U6253 (N_6253,N_6106,N_6077);
and U6254 (N_6254,N_6109,N_6039);
xor U6255 (N_6255,N_6020,N_6149);
or U6256 (N_6256,N_6074,N_6019);
and U6257 (N_6257,N_6071,N_6197);
or U6258 (N_6258,N_6108,N_6164);
nor U6259 (N_6259,N_6150,N_6011);
and U6260 (N_6260,N_6013,N_6015);
and U6261 (N_6261,N_6189,N_6055);
nand U6262 (N_6262,N_6147,N_6003);
or U6263 (N_6263,N_6128,N_6068);
xnor U6264 (N_6264,N_6045,N_6158);
and U6265 (N_6265,N_6083,N_6139);
xor U6266 (N_6266,N_6066,N_6022);
nand U6267 (N_6267,N_6092,N_6169);
and U6268 (N_6268,N_6155,N_6183);
or U6269 (N_6269,N_6144,N_6181);
nor U6270 (N_6270,N_6073,N_6008);
xnor U6271 (N_6271,N_6148,N_6193);
nand U6272 (N_6272,N_6053,N_6097);
nor U6273 (N_6273,N_6094,N_6190);
xor U6274 (N_6274,N_6054,N_6104);
nor U6275 (N_6275,N_6177,N_6121);
or U6276 (N_6276,N_6064,N_6080);
or U6277 (N_6277,N_6194,N_6115);
nand U6278 (N_6278,N_6171,N_6124);
nand U6279 (N_6279,N_6025,N_6188);
and U6280 (N_6280,N_6146,N_6153);
xnor U6281 (N_6281,N_6009,N_6086);
nor U6282 (N_6282,N_6180,N_6057);
and U6283 (N_6283,N_6174,N_6162);
nand U6284 (N_6284,N_6098,N_6165);
and U6285 (N_6285,N_6070,N_6049);
nand U6286 (N_6286,N_6067,N_6141);
xor U6287 (N_6287,N_6006,N_6186);
and U6288 (N_6288,N_6117,N_6037);
or U6289 (N_6289,N_6151,N_6161);
xnor U6290 (N_6290,N_6087,N_6096);
xor U6291 (N_6291,N_6044,N_6058);
or U6292 (N_6292,N_6145,N_6076);
nand U6293 (N_6293,N_6030,N_6122);
nand U6294 (N_6294,N_6088,N_6050);
xnor U6295 (N_6295,N_6184,N_6085);
nor U6296 (N_6296,N_6131,N_6107);
or U6297 (N_6297,N_6029,N_6032);
xnor U6298 (N_6298,N_6017,N_6103);
and U6299 (N_6299,N_6101,N_6093);
xnor U6300 (N_6300,N_6017,N_6074);
xnor U6301 (N_6301,N_6164,N_6115);
nor U6302 (N_6302,N_6199,N_6093);
nand U6303 (N_6303,N_6060,N_6029);
and U6304 (N_6304,N_6158,N_6181);
nor U6305 (N_6305,N_6061,N_6137);
nand U6306 (N_6306,N_6055,N_6154);
xnor U6307 (N_6307,N_6031,N_6100);
nor U6308 (N_6308,N_6157,N_6129);
and U6309 (N_6309,N_6169,N_6140);
or U6310 (N_6310,N_6161,N_6138);
nand U6311 (N_6311,N_6147,N_6016);
nand U6312 (N_6312,N_6036,N_6142);
or U6313 (N_6313,N_6043,N_6077);
nor U6314 (N_6314,N_6088,N_6033);
and U6315 (N_6315,N_6198,N_6089);
and U6316 (N_6316,N_6130,N_6005);
nand U6317 (N_6317,N_6184,N_6168);
xnor U6318 (N_6318,N_6015,N_6114);
or U6319 (N_6319,N_6023,N_6049);
and U6320 (N_6320,N_6181,N_6091);
nand U6321 (N_6321,N_6147,N_6130);
xnor U6322 (N_6322,N_6102,N_6056);
or U6323 (N_6323,N_6063,N_6044);
xor U6324 (N_6324,N_6031,N_6187);
xor U6325 (N_6325,N_6155,N_6091);
nand U6326 (N_6326,N_6133,N_6030);
or U6327 (N_6327,N_6056,N_6067);
and U6328 (N_6328,N_6018,N_6107);
nand U6329 (N_6329,N_6170,N_6172);
and U6330 (N_6330,N_6131,N_6173);
nand U6331 (N_6331,N_6136,N_6086);
xor U6332 (N_6332,N_6049,N_6193);
and U6333 (N_6333,N_6158,N_6109);
and U6334 (N_6334,N_6152,N_6033);
and U6335 (N_6335,N_6094,N_6161);
xnor U6336 (N_6336,N_6165,N_6190);
or U6337 (N_6337,N_6163,N_6144);
and U6338 (N_6338,N_6166,N_6086);
or U6339 (N_6339,N_6138,N_6199);
xnor U6340 (N_6340,N_6181,N_6183);
nand U6341 (N_6341,N_6191,N_6014);
nand U6342 (N_6342,N_6091,N_6179);
nand U6343 (N_6343,N_6134,N_6011);
xnor U6344 (N_6344,N_6119,N_6072);
nor U6345 (N_6345,N_6075,N_6183);
and U6346 (N_6346,N_6087,N_6149);
and U6347 (N_6347,N_6190,N_6111);
nor U6348 (N_6348,N_6063,N_6064);
or U6349 (N_6349,N_6146,N_6195);
xor U6350 (N_6350,N_6134,N_6184);
xnor U6351 (N_6351,N_6113,N_6049);
nor U6352 (N_6352,N_6131,N_6158);
nor U6353 (N_6353,N_6169,N_6079);
xor U6354 (N_6354,N_6034,N_6138);
xnor U6355 (N_6355,N_6034,N_6008);
nand U6356 (N_6356,N_6031,N_6044);
xor U6357 (N_6357,N_6182,N_6176);
xor U6358 (N_6358,N_6147,N_6142);
nand U6359 (N_6359,N_6019,N_6197);
nor U6360 (N_6360,N_6126,N_6112);
or U6361 (N_6361,N_6012,N_6020);
nor U6362 (N_6362,N_6013,N_6166);
xnor U6363 (N_6363,N_6144,N_6085);
and U6364 (N_6364,N_6125,N_6199);
nand U6365 (N_6365,N_6086,N_6004);
nor U6366 (N_6366,N_6169,N_6149);
or U6367 (N_6367,N_6174,N_6081);
or U6368 (N_6368,N_6198,N_6189);
nand U6369 (N_6369,N_6155,N_6134);
and U6370 (N_6370,N_6130,N_6017);
xor U6371 (N_6371,N_6167,N_6140);
nand U6372 (N_6372,N_6183,N_6050);
and U6373 (N_6373,N_6146,N_6033);
xnor U6374 (N_6374,N_6175,N_6110);
and U6375 (N_6375,N_6019,N_6091);
and U6376 (N_6376,N_6148,N_6087);
nand U6377 (N_6377,N_6056,N_6130);
xor U6378 (N_6378,N_6005,N_6079);
or U6379 (N_6379,N_6005,N_6195);
and U6380 (N_6380,N_6183,N_6032);
or U6381 (N_6381,N_6135,N_6052);
xor U6382 (N_6382,N_6121,N_6157);
and U6383 (N_6383,N_6063,N_6127);
nor U6384 (N_6384,N_6125,N_6101);
nand U6385 (N_6385,N_6194,N_6018);
nor U6386 (N_6386,N_6173,N_6110);
or U6387 (N_6387,N_6070,N_6018);
and U6388 (N_6388,N_6173,N_6032);
or U6389 (N_6389,N_6143,N_6191);
and U6390 (N_6390,N_6096,N_6153);
nand U6391 (N_6391,N_6160,N_6035);
nor U6392 (N_6392,N_6032,N_6080);
or U6393 (N_6393,N_6182,N_6071);
or U6394 (N_6394,N_6181,N_6134);
nor U6395 (N_6395,N_6052,N_6162);
nor U6396 (N_6396,N_6166,N_6162);
nand U6397 (N_6397,N_6002,N_6014);
and U6398 (N_6398,N_6022,N_6058);
nor U6399 (N_6399,N_6026,N_6153);
nor U6400 (N_6400,N_6231,N_6341);
and U6401 (N_6401,N_6297,N_6315);
xor U6402 (N_6402,N_6261,N_6336);
or U6403 (N_6403,N_6201,N_6397);
or U6404 (N_6404,N_6301,N_6391);
or U6405 (N_6405,N_6304,N_6228);
nor U6406 (N_6406,N_6330,N_6312);
xnor U6407 (N_6407,N_6242,N_6212);
nor U6408 (N_6408,N_6272,N_6357);
nand U6409 (N_6409,N_6363,N_6374);
xor U6410 (N_6410,N_6396,N_6246);
or U6411 (N_6411,N_6383,N_6210);
nand U6412 (N_6412,N_6290,N_6288);
and U6413 (N_6413,N_6305,N_6337);
xnor U6414 (N_6414,N_6342,N_6329);
and U6415 (N_6415,N_6227,N_6292);
or U6416 (N_6416,N_6253,N_6308);
and U6417 (N_6417,N_6259,N_6276);
and U6418 (N_6418,N_6247,N_6327);
and U6419 (N_6419,N_6318,N_6240);
nor U6420 (N_6420,N_6207,N_6347);
or U6421 (N_6421,N_6249,N_6239);
or U6422 (N_6422,N_6300,N_6204);
and U6423 (N_6423,N_6281,N_6332);
nor U6424 (N_6424,N_6203,N_6394);
or U6425 (N_6425,N_6248,N_6202);
nor U6426 (N_6426,N_6268,N_6226);
or U6427 (N_6427,N_6235,N_6265);
xor U6428 (N_6428,N_6271,N_6358);
or U6429 (N_6429,N_6244,N_6386);
nor U6430 (N_6430,N_6263,N_6262);
nand U6431 (N_6431,N_6215,N_6379);
xor U6432 (N_6432,N_6243,N_6388);
nor U6433 (N_6433,N_6291,N_6254);
xor U6434 (N_6434,N_6325,N_6369);
or U6435 (N_6435,N_6322,N_6283);
nor U6436 (N_6436,N_6303,N_6209);
and U6437 (N_6437,N_6314,N_6216);
and U6438 (N_6438,N_6373,N_6324);
and U6439 (N_6439,N_6277,N_6296);
xor U6440 (N_6440,N_6372,N_6392);
or U6441 (N_6441,N_6298,N_6229);
nor U6442 (N_6442,N_6217,N_6377);
nor U6443 (N_6443,N_6398,N_6345);
nand U6444 (N_6444,N_6355,N_6360);
or U6445 (N_6445,N_6295,N_6343);
and U6446 (N_6446,N_6359,N_6311);
xnor U6447 (N_6447,N_6278,N_6376);
nand U6448 (N_6448,N_6211,N_6393);
nand U6449 (N_6449,N_6351,N_6387);
and U6450 (N_6450,N_6293,N_6350);
or U6451 (N_6451,N_6331,N_6274);
xnor U6452 (N_6452,N_6238,N_6284);
nor U6453 (N_6453,N_6258,N_6326);
nand U6454 (N_6454,N_6237,N_6310);
nor U6455 (N_6455,N_6333,N_6371);
and U6456 (N_6456,N_6319,N_6214);
nor U6457 (N_6457,N_6241,N_6251);
or U6458 (N_6458,N_6356,N_6285);
nor U6459 (N_6459,N_6221,N_6368);
nor U6460 (N_6460,N_6399,N_6380);
and U6461 (N_6461,N_6313,N_6213);
nand U6462 (N_6462,N_6354,N_6346);
xnor U6463 (N_6463,N_6250,N_6282);
nand U6464 (N_6464,N_6234,N_6316);
xor U6465 (N_6465,N_6302,N_6299);
xnor U6466 (N_6466,N_6306,N_6279);
nand U6467 (N_6467,N_6362,N_6287);
nor U6468 (N_6468,N_6381,N_6390);
xor U6469 (N_6469,N_6321,N_6352);
and U6470 (N_6470,N_6267,N_6382);
nor U6471 (N_6471,N_6220,N_6206);
nand U6472 (N_6472,N_6219,N_6275);
nor U6473 (N_6473,N_6208,N_6270);
nor U6474 (N_6474,N_6349,N_6232);
or U6475 (N_6475,N_6286,N_6338);
and U6476 (N_6476,N_6395,N_6236);
nand U6477 (N_6477,N_6289,N_6364);
and U6478 (N_6478,N_6266,N_6320);
nor U6479 (N_6479,N_6273,N_6309);
nor U6480 (N_6480,N_6384,N_6200);
xor U6481 (N_6481,N_6367,N_6245);
and U6482 (N_6482,N_6340,N_6385);
or U6483 (N_6483,N_6222,N_6205);
and U6484 (N_6484,N_6264,N_6323);
and U6485 (N_6485,N_6224,N_6328);
nor U6486 (N_6486,N_6218,N_6344);
xor U6487 (N_6487,N_6233,N_6280);
and U6488 (N_6488,N_6255,N_6256);
or U6489 (N_6489,N_6294,N_6260);
or U6490 (N_6490,N_6334,N_6252);
or U6491 (N_6491,N_6370,N_6348);
nand U6492 (N_6492,N_6257,N_6375);
nor U6493 (N_6493,N_6335,N_6389);
or U6494 (N_6494,N_6230,N_6361);
or U6495 (N_6495,N_6365,N_6223);
nor U6496 (N_6496,N_6225,N_6339);
nor U6497 (N_6497,N_6269,N_6366);
and U6498 (N_6498,N_6317,N_6307);
or U6499 (N_6499,N_6378,N_6353);
and U6500 (N_6500,N_6271,N_6395);
and U6501 (N_6501,N_6365,N_6210);
and U6502 (N_6502,N_6225,N_6283);
nand U6503 (N_6503,N_6286,N_6368);
or U6504 (N_6504,N_6209,N_6349);
or U6505 (N_6505,N_6225,N_6229);
nor U6506 (N_6506,N_6379,N_6372);
nor U6507 (N_6507,N_6262,N_6317);
and U6508 (N_6508,N_6309,N_6256);
xnor U6509 (N_6509,N_6271,N_6223);
nand U6510 (N_6510,N_6268,N_6276);
nor U6511 (N_6511,N_6272,N_6207);
nand U6512 (N_6512,N_6209,N_6214);
and U6513 (N_6513,N_6357,N_6353);
nand U6514 (N_6514,N_6236,N_6277);
or U6515 (N_6515,N_6351,N_6286);
or U6516 (N_6516,N_6318,N_6259);
or U6517 (N_6517,N_6317,N_6234);
or U6518 (N_6518,N_6238,N_6246);
and U6519 (N_6519,N_6221,N_6323);
xor U6520 (N_6520,N_6354,N_6353);
nor U6521 (N_6521,N_6220,N_6386);
or U6522 (N_6522,N_6250,N_6213);
and U6523 (N_6523,N_6221,N_6336);
nand U6524 (N_6524,N_6355,N_6265);
nor U6525 (N_6525,N_6224,N_6386);
nand U6526 (N_6526,N_6281,N_6265);
xnor U6527 (N_6527,N_6236,N_6350);
and U6528 (N_6528,N_6223,N_6334);
nor U6529 (N_6529,N_6320,N_6309);
or U6530 (N_6530,N_6299,N_6317);
nand U6531 (N_6531,N_6246,N_6341);
xor U6532 (N_6532,N_6306,N_6233);
xnor U6533 (N_6533,N_6332,N_6262);
and U6534 (N_6534,N_6234,N_6219);
nor U6535 (N_6535,N_6242,N_6376);
and U6536 (N_6536,N_6320,N_6285);
xnor U6537 (N_6537,N_6242,N_6311);
nand U6538 (N_6538,N_6216,N_6231);
nor U6539 (N_6539,N_6234,N_6367);
and U6540 (N_6540,N_6213,N_6200);
nor U6541 (N_6541,N_6204,N_6343);
or U6542 (N_6542,N_6250,N_6296);
xor U6543 (N_6543,N_6318,N_6330);
or U6544 (N_6544,N_6285,N_6323);
and U6545 (N_6545,N_6333,N_6389);
nor U6546 (N_6546,N_6222,N_6208);
or U6547 (N_6547,N_6324,N_6218);
or U6548 (N_6548,N_6211,N_6392);
nor U6549 (N_6549,N_6364,N_6234);
xor U6550 (N_6550,N_6322,N_6300);
nor U6551 (N_6551,N_6221,N_6365);
or U6552 (N_6552,N_6318,N_6256);
nor U6553 (N_6553,N_6312,N_6319);
nor U6554 (N_6554,N_6293,N_6294);
nor U6555 (N_6555,N_6326,N_6276);
xor U6556 (N_6556,N_6200,N_6371);
nand U6557 (N_6557,N_6263,N_6353);
and U6558 (N_6558,N_6314,N_6301);
xor U6559 (N_6559,N_6368,N_6365);
or U6560 (N_6560,N_6237,N_6231);
nand U6561 (N_6561,N_6290,N_6200);
or U6562 (N_6562,N_6376,N_6298);
nand U6563 (N_6563,N_6349,N_6206);
and U6564 (N_6564,N_6213,N_6383);
xnor U6565 (N_6565,N_6227,N_6378);
nor U6566 (N_6566,N_6387,N_6230);
or U6567 (N_6567,N_6235,N_6279);
and U6568 (N_6568,N_6370,N_6225);
nand U6569 (N_6569,N_6321,N_6379);
nor U6570 (N_6570,N_6225,N_6234);
nand U6571 (N_6571,N_6257,N_6224);
or U6572 (N_6572,N_6256,N_6322);
and U6573 (N_6573,N_6351,N_6281);
xnor U6574 (N_6574,N_6305,N_6297);
or U6575 (N_6575,N_6304,N_6217);
and U6576 (N_6576,N_6280,N_6358);
and U6577 (N_6577,N_6375,N_6283);
nor U6578 (N_6578,N_6302,N_6390);
or U6579 (N_6579,N_6216,N_6278);
or U6580 (N_6580,N_6285,N_6223);
nor U6581 (N_6581,N_6357,N_6281);
nand U6582 (N_6582,N_6377,N_6373);
xor U6583 (N_6583,N_6302,N_6367);
or U6584 (N_6584,N_6357,N_6238);
xnor U6585 (N_6585,N_6244,N_6373);
xor U6586 (N_6586,N_6314,N_6307);
and U6587 (N_6587,N_6339,N_6384);
or U6588 (N_6588,N_6264,N_6321);
nor U6589 (N_6589,N_6339,N_6266);
nor U6590 (N_6590,N_6392,N_6342);
nand U6591 (N_6591,N_6389,N_6238);
nand U6592 (N_6592,N_6281,N_6254);
nand U6593 (N_6593,N_6216,N_6364);
nor U6594 (N_6594,N_6313,N_6224);
nand U6595 (N_6595,N_6306,N_6226);
or U6596 (N_6596,N_6316,N_6378);
nand U6597 (N_6597,N_6230,N_6289);
nand U6598 (N_6598,N_6380,N_6259);
or U6599 (N_6599,N_6336,N_6354);
or U6600 (N_6600,N_6445,N_6480);
or U6601 (N_6601,N_6591,N_6554);
nor U6602 (N_6602,N_6473,N_6497);
or U6603 (N_6603,N_6440,N_6495);
and U6604 (N_6604,N_6403,N_6546);
nor U6605 (N_6605,N_6413,N_6446);
nand U6606 (N_6606,N_6417,N_6562);
nor U6607 (N_6607,N_6581,N_6430);
nand U6608 (N_6608,N_6574,N_6448);
and U6609 (N_6609,N_6513,N_6578);
and U6610 (N_6610,N_6537,N_6443);
xor U6611 (N_6611,N_6585,N_6593);
nand U6612 (N_6612,N_6561,N_6421);
xor U6613 (N_6613,N_6577,N_6565);
or U6614 (N_6614,N_6540,N_6521);
xnor U6615 (N_6615,N_6427,N_6538);
nand U6616 (N_6616,N_6486,N_6525);
xnor U6617 (N_6617,N_6447,N_6425);
or U6618 (N_6618,N_6559,N_6594);
nand U6619 (N_6619,N_6514,N_6586);
or U6620 (N_6620,N_6457,N_6583);
nor U6621 (N_6621,N_6478,N_6428);
nand U6622 (N_6622,N_6483,N_6579);
and U6623 (N_6623,N_6512,N_6547);
nand U6624 (N_6624,N_6558,N_6508);
nand U6625 (N_6625,N_6541,N_6534);
nor U6626 (N_6626,N_6568,N_6501);
nor U6627 (N_6627,N_6460,N_6432);
and U6628 (N_6628,N_6436,N_6529);
and U6629 (N_6629,N_6477,N_6535);
xor U6630 (N_6630,N_6418,N_6438);
or U6631 (N_6631,N_6596,N_6557);
nor U6632 (N_6632,N_6416,N_6400);
nor U6633 (N_6633,N_6548,N_6465);
or U6634 (N_6634,N_6450,N_6429);
and U6635 (N_6635,N_6412,N_6479);
and U6636 (N_6636,N_6588,N_6544);
xnor U6637 (N_6637,N_6598,N_6408);
or U6638 (N_6638,N_6556,N_6406);
xor U6639 (N_6639,N_6464,N_6407);
nand U6640 (N_6640,N_6563,N_6506);
or U6641 (N_6641,N_6491,N_6461);
and U6642 (N_6642,N_6481,N_6519);
xnor U6643 (N_6643,N_6552,N_6505);
nand U6644 (N_6644,N_6597,N_6433);
and U6645 (N_6645,N_6507,N_6553);
nand U6646 (N_6646,N_6459,N_6455);
xnor U6647 (N_6647,N_6405,N_6437);
nor U6648 (N_6648,N_6402,N_6410);
and U6649 (N_6649,N_6543,N_6462);
and U6650 (N_6650,N_6571,N_6422);
nand U6651 (N_6651,N_6442,N_6489);
and U6652 (N_6652,N_6549,N_6490);
or U6653 (N_6653,N_6415,N_6502);
and U6654 (N_6654,N_6569,N_6470);
xor U6655 (N_6655,N_6466,N_6409);
nor U6656 (N_6656,N_6527,N_6524);
and U6657 (N_6657,N_6496,N_6589);
xnor U6658 (N_6658,N_6522,N_6471);
xor U6659 (N_6659,N_6456,N_6426);
nor U6660 (N_6660,N_6551,N_6492);
nand U6661 (N_6661,N_6511,N_6494);
or U6662 (N_6662,N_6587,N_6475);
and U6663 (N_6663,N_6444,N_6449);
and U6664 (N_6664,N_6482,N_6555);
nor U6665 (N_6665,N_6420,N_6528);
nand U6666 (N_6666,N_6504,N_6404);
nand U6667 (N_6667,N_6510,N_6573);
xnor U6668 (N_6668,N_6564,N_6570);
xor U6669 (N_6669,N_6531,N_6542);
and U6670 (N_6670,N_6434,N_6414);
and U6671 (N_6671,N_6498,N_6560);
nor U6672 (N_6672,N_6485,N_6423);
or U6673 (N_6673,N_6545,N_6493);
xor U6674 (N_6674,N_6592,N_6539);
and U6675 (N_6675,N_6441,N_6575);
or U6676 (N_6676,N_6530,N_6572);
nor U6677 (N_6677,N_6424,N_6520);
or U6678 (N_6678,N_6463,N_6467);
nor U6679 (N_6679,N_6476,N_6435);
nor U6680 (N_6680,N_6595,N_6472);
and U6681 (N_6681,N_6468,N_6536);
xor U6682 (N_6682,N_6517,N_6453);
or U6683 (N_6683,N_6439,N_6431);
and U6684 (N_6684,N_6458,N_6500);
nand U6685 (N_6685,N_6401,N_6452);
and U6686 (N_6686,N_6532,N_6584);
xnor U6687 (N_6687,N_6533,N_6516);
or U6688 (N_6688,N_6582,N_6419);
or U6689 (N_6689,N_6469,N_6515);
and U6690 (N_6690,N_6474,N_6509);
nand U6691 (N_6691,N_6599,N_6590);
and U6692 (N_6692,N_6576,N_6566);
nor U6693 (N_6693,N_6518,N_6484);
or U6694 (N_6694,N_6523,N_6580);
or U6695 (N_6695,N_6411,N_6488);
nor U6696 (N_6696,N_6451,N_6499);
xnor U6697 (N_6697,N_6567,N_6503);
and U6698 (N_6698,N_6550,N_6454);
and U6699 (N_6699,N_6487,N_6526);
or U6700 (N_6700,N_6548,N_6472);
and U6701 (N_6701,N_6478,N_6539);
xnor U6702 (N_6702,N_6556,N_6571);
nand U6703 (N_6703,N_6509,N_6405);
or U6704 (N_6704,N_6530,N_6552);
nand U6705 (N_6705,N_6551,N_6447);
or U6706 (N_6706,N_6473,N_6427);
xor U6707 (N_6707,N_6508,N_6518);
nor U6708 (N_6708,N_6551,N_6472);
nand U6709 (N_6709,N_6460,N_6549);
or U6710 (N_6710,N_6411,N_6410);
xor U6711 (N_6711,N_6429,N_6545);
or U6712 (N_6712,N_6568,N_6404);
xnor U6713 (N_6713,N_6419,N_6501);
nand U6714 (N_6714,N_6527,N_6441);
nor U6715 (N_6715,N_6461,N_6523);
nand U6716 (N_6716,N_6562,N_6483);
nand U6717 (N_6717,N_6514,N_6402);
or U6718 (N_6718,N_6433,N_6572);
or U6719 (N_6719,N_6593,N_6423);
nor U6720 (N_6720,N_6515,N_6414);
nor U6721 (N_6721,N_6493,N_6445);
xor U6722 (N_6722,N_6506,N_6415);
or U6723 (N_6723,N_6414,N_6444);
and U6724 (N_6724,N_6525,N_6540);
xor U6725 (N_6725,N_6580,N_6525);
and U6726 (N_6726,N_6523,N_6519);
and U6727 (N_6727,N_6490,N_6585);
or U6728 (N_6728,N_6508,N_6438);
xor U6729 (N_6729,N_6438,N_6404);
xor U6730 (N_6730,N_6455,N_6563);
or U6731 (N_6731,N_6555,N_6574);
nand U6732 (N_6732,N_6535,N_6501);
nor U6733 (N_6733,N_6457,N_6469);
nand U6734 (N_6734,N_6471,N_6463);
xnor U6735 (N_6735,N_6506,N_6586);
or U6736 (N_6736,N_6575,N_6577);
nor U6737 (N_6737,N_6516,N_6574);
or U6738 (N_6738,N_6408,N_6546);
and U6739 (N_6739,N_6483,N_6471);
or U6740 (N_6740,N_6583,N_6544);
or U6741 (N_6741,N_6555,N_6450);
nand U6742 (N_6742,N_6466,N_6571);
and U6743 (N_6743,N_6521,N_6470);
nor U6744 (N_6744,N_6497,N_6536);
xnor U6745 (N_6745,N_6532,N_6451);
or U6746 (N_6746,N_6407,N_6480);
xor U6747 (N_6747,N_6448,N_6427);
and U6748 (N_6748,N_6552,N_6446);
or U6749 (N_6749,N_6453,N_6555);
and U6750 (N_6750,N_6571,N_6518);
or U6751 (N_6751,N_6516,N_6548);
or U6752 (N_6752,N_6534,N_6473);
nand U6753 (N_6753,N_6474,N_6493);
nand U6754 (N_6754,N_6564,N_6417);
or U6755 (N_6755,N_6504,N_6525);
and U6756 (N_6756,N_6403,N_6597);
nor U6757 (N_6757,N_6423,N_6461);
nand U6758 (N_6758,N_6516,N_6535);
nand U6759 (N_6759,N_6498,N_6458);
nand U6760 (N_6760,N_6484,N_6435);
and U6761 (N_6761,N_6553,N_6456);
nand U6762 (N_6762,N_6445,N_6401);
nand U6763 (N_6763,N_6414,N_6405);
nand U6764 (N_6764,N_6540,N_6532);
nor U6765 (N_6765,N_6530,N_6448);
xnor U6766 (N_6766,N_6469,N_6528);
or U6767 (N_6767,N_6488,N_6413);
nand U6768 (N_6768,N_6587,N_6507);
xnor U6769 (N_6769,N_6436,N_6589);
nor U6770 (N_6770,N_6524,N_6419);
xor U6771 (N_6771,N_6447,N_6418);
nor U6772 (N_6772,N_6444,N_6466);
or U6773 (N_6773,N_6543,N_6499);
or U6774 (N_6774,N_6483,N_6427);
or U6775 (N_6775,N_6548,N_6416);
and U6776 (N_6776,N_6507,N_6584);
and U6777 (N_6777,N_6564,N_6452);
nand U6778 (N_6778,N_6479,N_6579);
nor U6779 (N_6779,N_6472,N_6414);
nand U6780 (N_6780,N_6428,N_6410);
xnor U6781 (N_6781,N_6416,N_6519);
or U6782 (N_6782,N_6402,N_6481);
nor U6783 (N_6783,N_6552,N_6448);
or U6784 (N_6784,N_6500,N_6556);
and U6785 (N_6785,N_6409,N_6565);
nor U6786 (N_6786,N_6401,N_6521);
nor U6787 (N_6787,N_6405,N_6468);
xor U6788 (N_6788,N_6484,N_6433);
or U6789 (N_6789,N_6493,N_6587);
xnor U6790 (N_6790,N_6545,N_6414);
nor U6791 (N_6791,N_6592,N_6519);
nor U6792 (N_6792,N_6408,N_6494);
xor U6793 (N_6793,N_6503,N_6507);
and U6794 (N_6794,N_6575,N_6460);
nand U6795 (N_6795,N_6443,N_6534);
or U6796 (N_6796,N_6471,N_6523);
nor U6797 (N_6797,N_6417,N_6532);
nand U6798 (N_6798,N_6555,N_6498);
nand U6799 (N_6799,N_6446,N_6530);
or U6800 (N_6800,N_6797,N_6715);
xor U6801 (N_6801,N_6682,N_6697);
nand U6802 (N_6802,N_6648,N_6745);
nand U6803 (N_6803,N_6725,N_6664);
and U6804 (N_6804,N_6646,N_6754);
nand U6805 (N_6805,N_6683,N_6778);
or U6806 (N_6806,N_6724,N_6676);
nor U6807 (N_6807,N_6623,N_6631);
or U6808 (N_6808,N_6638,N_6726);
nand U6809 (N_6809,N_6708,N_6776);
nand U6810 (N_6810,N_6767,N_6758);
xor U6811 (N_6811,N_6639,N_6600);
nand U6812 (N_6812,N_6735,N_6762);
xnor U6813 (N_6813,N_6627,N_6771);
nand U6814 (N_6814,N_6605,N_6662);
nor U6815 (N_6815,N_6670,N_6783);
or U6816 (N_6816,N_6789,N_6606);
nor U6817 (N_6817,N_6685,N_6748);
or U6818 (N_6818,N_6667,N_6669);
xnor U6819 (N_6819,N_6739,N_6652);
xnor U6820 (N_6820,N_6668,N_6782);
nor U6821 (N_6821,N_6659,N_6624);
nand U6822 (N_6822,N_6722,N_6677);
or U6823 (N_6823,N_6728,N_6717);
xor U6824 (N_6824,N_6770,N_6755);
or U6825 (N_6825,N_6614,N_6740);
nand U6826 (N_6826,N_6780,N_6727);
nand U6827 (N_6827,N_6759,N_6633);
xor U6828 (N_6828,N_6637,N_6622);
or U6829 (N_6829,N_6634,N_6651);
and U6830 (N_6830,N_6751,N_6732);
and U6831 (N_6831,N_6793,N_6753);
nand U6832 (N_6832,N_6635,N_6684);
nor U6833 (N_6833,N_6699,N_6680);
or U6834 (N_6834,N_6613,N_6774);
or U6835 (N_6835,N_6612,N_6742);
and U6836 (N_6836,N_6773,N_6690);
nor U6837 (N_6837,N_6629,N_6616);
and U6838 (N_6838,N_6709,N_6747);
and U6839 (N_6839,N_6731,N_6628);
nor U6840 (N_6840,N_6647,N_6666);
and U6841 (N_6841,N_6791,N_6686);
nand U6842 (N_6842,N_6607,N_6632);
nor U6843 (N_6843,N_6763,N_6746);
or U6844 (N_6844,N_6723,N_6781);
and U6845 (N_6845,N_6772,N_6665);
nor U6846 (N_6846,N_6744,N_6719);
nor U6847 (N_6847,N_6649,N_6660);
nand U6848 (N_6848,N_6604,N_6714);
xnor U6849 (N_6849,N_6757,N_6673);
and U6850 (N_6850,N_6626,N_6784);
or U6851 (N_6851,N_6752,N_6603);
or U6852 (N_6852,N_6703,N_6701);
nand U6853 (N_6853,N_6679,N_6795);
nor U6854 (N_6854,N_6650,N_6602);
xnor U6855 (N_6855,N_6702,N_6687);
and U6856 (N_6856,N_6707,N_6678);
and U6857 (N_6857,N_6619,N_6796);
nor U6858 (N_6858,N_6644,N_6672);
nand U6859 (N_6859,N_6716,N_6601);
nand U6860 (N_6860,N_6658,N_6645);
xor U6861 (N_6861,N_6705,N_6734);
and U6862 (N_6862,N_6769,N_6653);
nor U6863 (N_6863,N_6711,N_6766);
or U6864 (N_6864,N_6741,N_6698);
xor U6865 (N_6865,N_6640,N_6790);
nand U6866 (N_6866,N_6736,N_6794);
nor U6867 (N_6867,N_6663,N_6636);
or U6868 (N_6868,N_6610,N_6733);
or U6869 (N_6869,N_6694,N_6661);
and U6870 (N_6870,N_6787,N_6765);
xor U6871 (N_6871,N_6729,N_6712);
nor U6872 (N_6872,N_6691,N_6655);
xnor U6873 (N_6873,N_6799,N_6798);
xnor U6874 (N_6874,N_6617,N_6764);
xnor U6875 (N_6875,N_6775,N_6630);
or U6876 (N_6876,N_6611,N_6761);
xnor U6877 (N_6877,N_6720,N_6768);
nor U6878 (N_6878,N_6608,N_6738);
and U6879 (N_6879,N_6641,N_6643);
nor U6880 (N_6880,N_6693,N_6760);
and U6881 (N_6881,N_6788,N_6625);
nor U6882 (N_6882,N_6743,N_6786);
nor U6883 (N_6883,N_6671,N_6721);
or U6884 (N_6884,N_6730,N_6615);
xor U6885 (N_6885,N_6710,N_6696);
or U6886 (N_6886,N_6656,N_6737);
nand U6887 (N_6887,N_6777,N_6695);
or U6888 (N_6888,N_6785,N_6700);
or U6889 (N_6889,N_6618,N_6642);
and U6890 (N_6890,N_6750,N_6713);
nand U6891 (N_6891,N_6675,N_6756);
nor U6892 (N_6892,N_6792,N_6620);
or U6893 (N_6893,N_6749,N_6609);
nor U6894 (N_6894,N_6654,N_6681);
nand U6895 (N_6895,N_6706,N_6689);
or U6896 (N_6896,N_6718,N_6779);
or U6897 (N_6897,N_6674,N_6688);
and U6898 (N_6898,N_6657,N_6704);
xor U6899 (N_6899,N_6621,N_6692);
nand U6900 (N_6900,N_6630,N_6601);
and U6901 (N_6901,N_6717,N_6650);
or U6902 (N_6902,N_6674,N_6615);
xor U6903 (N_6903,N_6687,N_6686);
xor U6904 (N_6904,N_6714,N_6784);
xnor U6905 (N_6905,N_6736,N_6656);
nand U6906 (N_6906,N_6665,N_6660);
nand U6907 (N_6907,N_6684,N_6686);
or U6908 (N_6908,N_6737,N_6633);
xnor U6909 (N_6909,N_6786,N_6667);
nand U6910 (N_6910,N_6797,N_6654);
or U6911 (N_6911,N_6660,N_6676);
or U6912 (N_6912,N_6649,N_6696);
nand U6913 (N_6913,N_6776,N_6642);
nand U6914 (N_6914,N_6750,N_6732);
or U6915 (N_6915,N_6797,N_6635);
xor U6916 (N_6916,N_6601,N_6771);
nor U6917 (N_6917,N_6643,N_6626);
and U6918 (N_6918,N_6725,N_6674);
and U6919 (N_6919,N_6684,N_6657);
nor U6920 (N_6920,N_6775,N_6636);
and U6921 (N_6921,N_6628,N_6780);
xor U6922 (N_6922,N_6740,N_6721);
and U6923 (N_6923,N_6669,N_6721);
and U6924 (N_6924,N_6684,N_6601);
and U6925 (N_6925,N_6712,N_6751);
xor U6926 (N_6926,N_6661,N_6651);
nand U6927 (N_6927,N_6749,N_6669);
nand U6928 (N_6928,N_6709,N_6687);
nor U6929 (N_6929,N_6783,N_6773);
xnor U6930 (N_6930,N_6657,N_6702);
nor U6931 (N_6931,N_6667,N_6731);
nand U6932 (N_6932,N_6741,N_6738);
xnor U6933 (N_6933,N_6699,N_6657);
or U6934 (N_6934,N_6760,N_6671);
xnor U6935 (N_6935,N_6688,N_6785);
xnor U6936 (N_6936,N_6758,N_6648);
xnor U6937 (N_6937,N_6703,N_6636);
and U6938 (N_6938,N_6683,N_6773);
xnor U6939 (N_6939,N_6641,N_6790);
and U6940 (N_6940,N_6733,N_6669);
and U6941 (N_6941,N_6735,N_6668);
xor U6942 (N_6942,N_6747,N_6688);
xor U6943 (N_6943,N_6603,N_6714);
and U6944 (N_6944,N_6651,N_6656);
xor U6945 (N_6945,N_6737,N_6634);
nor U6946 (N_6946,N_6739,N_6767);
and U6947 (N_6947,N_6634,N_6790);
nor U6948 (N_6948,N_6637,N_6740);
or U6949 (N_6949,N_6695,N_6706);
and U6950 (N_6950,N_6625,N_6708);
or U6951 (N_6951,N_6780,N_6668);
nor U6952 (N_6952,N_6636,N_6789);
or U6953 (N_6953,N_6790,N_6700);
or U6954 (N_6954,N_6701,N_6716);
nand U6955 (N_6955,N_6747,N_6783);
nor U6956 (N_6956,N_6677,N_6634);
or U6957 (N_6957,N_6604,N_6772);
nor U6958 (N_6958,N_6624,N_6792);
nand U6959 (N_6959,N_6653,N_6605);
nor U6960 (N_6960,N_6762,N_6682);
nor U6961 (N_6961,N_6650,N_6743);
nor U6962 (N_6962,N_6711,N_6657);
nor U6963 (N_6963,N_6757,N_6747);
nor U6964 (N_6964,N_6720,N_6654);
or U6965 (N_6965,N_6692,N_6743);
and U6966 (N_6966,N_6625,N_6705);
nand U6967 (N_6967,N_6741,N_6685);
nand U6968 (N_6968,N_6674,N_6768);
xnor U6969 (N_6969,N_6655,N_6722);
nor U6970 (N_6970,N_6632,N_6774);
nor U6971 (N_6971,N_6773,N_6747);
xor U6972 (N_6972,N_6724,N_6654);
and U6973 (N_6973,N_6764,N_6783);
xor U6974 (N_6974,N_6703,N_6735);
nand U6975 (N_6975,N_6634,N_6600);
nand U6976 (N_6976,N_6760,N_6710);
or U6977 (N_6977,N_6718,N_6746);
and U6978 (N_6978,N_6682,N_6719);
nor U6979 (N_6979,N_6695,N_6717);
nand U6980 (N_6980,N_6618,N_6689);
xor U6981 (N_6981,N_6614,N_6759);
nor U6982 (N_6982,N_6779,N_6639);
nand U6983 (N_6983,N_6799,N_6783);
nand U6984 (N_6984,N_6658,N_6737);
or U6985 (N_6985,N_6664,N_6742);
nand U6986 (N_6986,N_6675,N_6634);
and U6987 (N_6987,N_6762,N_6772);
nor U6988 (N_6988,N_6676,N_6694);
and U6989 (N_6989,N_6769,N_6784);
nand U6990 (N_6990,N_6731,N_6792);
nor U6991 (N_6991,N_6614,N_6604);
and U6992 (N_6992,N_6666,N_6731);
or U6993 (N_6993,N_6694,N_6727);
xnor U6994 (N_6994,N_6669,N_6790);
and U6995 (N_6995,N_6737,N_6716);
and U6996 (N_6996,N_6787,N_6747);
xnor U6997 (N_6997,N_6788,N_6694);
xor U6998 (N_6998,N_6695,N_6758);
and U6999 (N_6999,N_6711,N_6790);
xnor U7000 (N_7000,N_6985,N_6839);
or U7001 (N_7001,N_6992,N_6855);
or U7002 (N_7002,N_6853,N_6967);
xor U7003 (N_7003,N_6826,N_6838);
nor U7004 (N_7004,N_6902,N_6983);
nand U7005 (N_7005,N_6963,N_6968);
nor U7006 (N_7006,N_6820,N_6828);
xnor U7007 (N_7007,N_6837,N_6805);
nor U7008 (N_7008,N_6958,N_6980);
nor U7009 (N_7009,N_6941,N_6823);
and U7010 (N_7010,N_6906,N_6933);
and U7011 (N_7011,N_6897,N_6912);
or U7012 (N_7012,N_6971,N_6830);
or U7013 (N_7013,N_6871,N_6896);
nand U7014 (N_7014,N_6850,N_6928);
or U7015 (N_7015,N_6852,N_6993);
and U7016 (N_7016,N_6973,N_6869);
nor U7017 (N_7017,N_6816,N_6931);
or U7018 (N_7018,N_6865,N_6870);
xnor U7019 (N_7019,N_6821,N_6894);
xnor U7020 (N_7020,N_6951,N_6898);
and U7021 (N_7021,N_6950,N_6920);
or U7022 (N_7022,N_6803,N_6909);
and U7023 (N_7023,N_6978,N_6910);
nor U7024 (N_7024,N_6945,N_6974);
xor U7025 (N_7025,N_6943,N_6988);
nand U7026 (N_7026,N_6825,N_6995);
and U7027 (N_7027,N_6848,N_6884);
nand U7028 (N_7028,N_6877,N_6957);
nor U7029 (N_7029,N_6913,N_6812);
nand U7030 (N_7030,N_6858,N_6955);
xnor U7031 (N_7031,N_6999,N_6804);
nor U7032 (N_7032,N_6881,N_6873);
nand U7033 (N_7033,N_6972,N_6827);
and U7034 (N_7034,N_6814,N_6960);
xor U7035 (N_7035,N_6859,N_6867);
nand U7036 (N_7036,N_6854,N_6815);
and U7037 (N_7037,N_6806,N_6887);
xnor U7038 (N_7038,N_6885,N_6856);
nand U7039 (N_7039,N_6818,N_6914);
or U7040 (N_7040,N_6901,N_6948);
nand U7041 (N_7041,N_6890,N_6861);
nor U7042 (N_7042,N_6840,N_6969);
xnor U7043 (N_7043,N_6918,N_6886);
nand U7044 (N_7044,N_6893,N_6936);
nor U7045 (N_7045,N_6811,N_6998);
nor U7046 (N_7046,N_6961,N_6868);
nand U7047 (N_7047,N_6834,N_6964);
or U7048 (N_7048,N_6975,N_6833);
xnor U7049 (N_7049,N_6925,N_6824);
nor U7050 (N_7050,N_6846,N_6956);
nor U7051 (N_7051,N_6832,N_6882);
nand U7052 (N_7052,N_6862,N_6892);
nor U7053 (N_7053,N_6940,N_6900);
xnor U7054 (N_7054,N_6908,N_6875);
and U7055 (N_7055,N_6949,N_6891);
and U7056 (N_7056,N_6845,N_6970);
nor U7057 (N_7057,N_6919,N_6847);
nand U7058 (N_7058,N_6903,N_6986);
and U7059 (N_7059,N_6874,N_6997);
xor U7060 (N_7060,N_6981,N_6899);
nor U7061 (N_7061,N_6879,N_6926);
nor U7062 (N_7062,N_6810,N_6917);
and U7063 (N_7063,N_6801,N_6813);
xnor U7064 (N_7064,N_6939,N_6905);
nor U7065 (N_7065,N_6921,N_6924);
or U7066 (N_7066,N_6984,N_6937);
nand U7067 (N_7067,N_6935,N_6907);
xor U7068 (N_7068,N_6916,N_6883);
nor U7069 (N_7069,N_6944,N_6994);
nor U7070 (N_7070,N_6831,N_6932);
and U7071 (N_7071,N_6895,N_6965);
nand U7072 (N_7072,N_6991,N_6987);
nand U7073 (N_7073,N_6982,N_6817);
nand U7074 (N_7074,N_6849,N_6923);
xnor U7075 (N_7075,N_6990,N_6915);
or U7076 (N_7076,N_6947,N_6819);
nor U7077 (N_7077,N_6876,N_6977);
and U7078 (N_7078,N_6864,N_6942);
nand U7079 (N_7079,N_6996,N_6880);
or U7080 (N_7080,N_6946,N_6857);
or U7081 (N_7081,N_6952,N_6872);
nand U7082 (N_7082,N_6904,N_6843);
and U7083 (N_7083,N_6842,N_6976);
or U7084 (N_7084,N_6927,N_6959);
or U7085 (N_7085,N_6929,N_6922);
nor U7086 (N_7086,N_6930,N_6866);
and U7087 (N_7087,N_6809,N_6800);
nor U7088 (N_7088,N_6953,N_6829);
nor U7089 (N_7089,N_6989,N_6822);
nor U7090 (N_7090,N_6863,N_6934);
nor U7091 (N_7091,N_6979,N_6808);
nand U7092 (N_7092,N_6889,N_6844);
xor U7093 (N_7093,N_6802,N_6966);
and U7094 (N_7094,N_6851,N_6938);
and U7095 (N_7095,N_6878,N_6962);
nand U7096 (N_7096,N_6835,N_6860);
nand U7097 (N_7097,N_6807,N_6888);
and U7098 (N_7098,N_6841,N_6911);
xor U7099 (N_7099,N_6954,N_6836);
nand U7100 (N_7100,N_6876,N_6832);
and U7101 (N_7101,N_6869,N_6960);
and U7102 (N_7102,N_6882,N_6944);
nand U7103 (N_7103,N_6843,N_6971);
nor U7104 (N_7104,N_6854,N_6893);
nand U7105 (N_7105,N_6944,N_6853);
and U7106 (N_7106,N_6935,N_6983);
xor U7107 (N_7107,N_6988,N_6903);
or U7108 (N_7108,N_6804,N_6924);
nor U7109 (N_7109,N_6841,N_6965);
nand U7110 (N_7110,N_6951,N_6927);
and U7111 (N_7111,N_6821,N_6936);
nor U7112 (N_7112,N_6991,N_6818);
nor U7113 (N_7113,N_6985,N_6875);
nor U7114 (N_7114,N_6830,N_6889);
xnor U7115 (N_7115,N_6966,N_6948);
nand U7116 (N_7116,N_6848,N_6856);
xnor U7117 (N_7117,N_6920,N_6954);
nor U7118 (N_7118,N_6869,N_6828);
nor U7119 (N_7119,N_6955,N_6800);
nor U7120 (N_7120,N_6955,N_6975);
xnor U7121 (N_7121,N_6970,N_6860);
or U7122 (N_7122,N_6991,N_6928);
xor U7123 (N_7123,N_6972,N_6872);
or U7124 (N_7124,N_6922,N_6847);
nor U7125 (N_7125,N_6978,N_6874);
nor U7126 (N_7126,N_6977,N_6834);
nor U7127 (N_7127,N_6847,N_6881);
xnor U7128 (N_7128,N_6977,N_6978);
nor U7129 (N_7129,N_6809,N_6877);
xor U7130 (N_7130,N_6953,N_6818);
and U7131 (N_7131,N_6960,N_6889);
and U7132 (N_7132,N_6954,N_6945);
nor U7133 (N_7133,N_6850,N_6950);
xor U7134 (N_7134,N_6806,N_6996);
nand U7135 (N_7135,N_6811,N_6901);
xor U7136 (N_7136,N_6946,N_6854);
or U7137 (N_7137,N_6872,N_6953);
nor U7138 (N_7138,N_6972,N_6849);
nand U7139 (N_7139,N_6881,N_6861);
and U7140 (N_7140,N_6857,N_6853);
xnor U7141 (N_7141,N_6883,N_6992);
xor U7142 (N_7142,N_6931,N_6986);
nand U7143 (N_7143,N_6893,N_6989);
or U7144 (N_7144,N_6935,N_6829);
nor U7145 (N_7145,N_6908,N_6825);
nand U7146 (N_7146,N_6852,N_6903);
nand U7147 (N_7147,N_6814,N_6991);
nand U7148 (N_7148,N_6928,N_6894);
xnor U7149 (N_7149,N_6829,N_6965);
and U7150 (N_7150,N_6986,N_6907);
and U7151 (N_7151,N_6911,N_6902);
xnor U7152 (N_7152,N_6922,N_6899);
nand U7153 (N_7153,N_6978,N_6834);
and U7154 (N_7154,N_6958,N_6857);
nor U7155 (N_7155,N_6891,N_6800);
and U7156 (N_7156,N_6931,N_6972);
nand U7157 (N_7157,N_6884,N_6983);
xor U7158 (N_7158,N_6865,N_6984);
nand U7159 (N_7159,N_6869,N_6892);
and U7160 (N_7160,N_6872,N_6986);
nand U7161 (N_7161,N_6859,N_6996);
and U7162 (N_7162,N_6996,N_6804);
nor U7163 (N_7163,N_6903,N_6893);
nor U7164 (N_7164,N_6978,N_6963);
xnor U7165 (N_7165,N_6818,N_6945);
xor U7166 (N_7166,N_6862,N_6986);
and U7167 (N_7167,N_6840,N_6876);
nand U7168 (N_7168,N_6804,N_6808);
xor U7169 (N_7169,N_6972,N_6927);
and U7170 (N_7170,N_6867,N_6991);
or U7171 (N_7171,N_6902,N_6816);
nand U7172 (N_7172,N_6870,N_6999);
nor U7173 (N_7173,N_6868,N_6827);
xnor U7174 (N_7174,N_6922,N_6952);
and U7175 (N_7175,N_6817,N_6845);
and U7176 (N_7176,N_6969,N_6937);
nand U7177 (N_7177,N_6890,N_6896);
and U7178 (N_7178,N_6853,N_6836);
xor U7179 (N_7179,N_6905,N_6884);
nand U7180 (N_7180,N_6949,N_6810);
nor U7181 (N_7181,N_6898,N_6966);
xnor U7182 (N_7182,N_6966,N_6883);
nand U7183 (N_7183,N_6983,N_6835);
nor U7184 (N_7184,N_6990,N_6881);
or U7185 (N_7185,N_6893,N_6803);
nor U7186 (N_7186,N_6925,N_6866);
or U7187 (N_7187,N_6879,N_6844);
and U7188 (N_7188,N_6996,N_6803);
and U7189 (N_7189,N_6870,N_6914);
and U7190 (N_7190,N_6806,N_6848);
and U7191 (N_7191,N_6966,N_6882);
and U7192 (N_7192,N_6817,N_6814);
nor U7193 (N_7193,N_6969,N_6923);
and U7194 (N_7194,N_6870,N_6900);
nor U7195 (N_7195,N_6951,N_6804);
and U7196 (N_7196,N_6840,N_6899);
or U7197 (N_7197,N_6808,N_6921);
or U7198 (N_7198,N_6920,N_6862);
and U7199 (N_7199,N_6894,N_6807);
and U7200 (N_7200,N_7001,N_7024);
xnor U7201 (N_7201,N_7078,N_7195);
xor U7202 (N_7202,N_7002,N_7067);
xnor U7203 (N_7203,N_7039,N_7079);
nand U7204 (N_7204,N_7167,N_7106);
and U7205 (N_7205,N_7189,N_7083);
nand U7206 (N_7206,N_7111,N_7118);
nand U7207 (N_7207,N_7093,N_7066);
nand U7208 (N_7208,N_7133,N_7197);
nand U7209 (N_7209,N_7035,N_7100);
or U7210 (N_7210,N_7187,N_7003);
and U7211 (N_7211,N_7082,N_7037);
xor U7212 (N_7212,N_7096,N_7006);
or U7213 (N_7213,N_7041,N_7159);
and U7214 (N_7214,N_7053,N_7177);
nor U7215 (N_7215,N_7031,N_7130);
nand U7216 (N_7216,N_7050,N_7112);
nand U7217 (N_7217,N_7184,N_7058);
nor U7218 (N_7218,N_7152,N_7073);
nor U7219 (N_7219,N_7188,N_7153);
nor U7220 (N_7220,N_7116,N_7007);
and U7221 (N_7221,N_7014,N_7183);
and U7222 (N_7222,N_7095,N_7028);
or U7223 (N_7223,N_7127,N_7179);
xor U7224 (N_7224,N_7036,N_7155);
nor U7225 (N_7225,N_7180,N_7142);
nand U7226 (N_7226,N_7048,N_7134);
or U7227 (N_7227,N_7145,N_7047);
nor U7228 (N_7228,N_7056,N_7062);
nor U7229 (N_7229,N_7172,N_7015);
or U7230 (N_7230,N_7054,N_7123);
xnor U7231 (N_7231,N_7136,N_7161);
or U7232 (N_7232,N_7021,N_7104);
and U7233 (N_7233,N_7072,N_7023);
nor U7234 (N_7234,N_7141,N_7119);
or U7235 (N_7235,N_7005,N_7191);
and U7236 (N_7236,N_7122,N_7102);
nand U7237 (N_7237,N_7089,N_7160);
nor U7238 (N_7238,N_7055,N_7107);
nor U7239 (N_7239,N_7128,N_7109);
nor U7240 (N_7240,N_7193,N_7090);
or U7241 (N_7241,N_7069,N_7174);
nand U7242 (N_7242,N_7144,N_7080);
nand U7243 (N_7243,N_7076,N_7008);
nand U7244 (N_7244,N_7020,N_7018);
xnor U7245 (N_7245,N_7052,N_7022);
nor U7246 (N_7246,N_7040,N_7097);
or U7247 (N_7247,N_7171,N_7060);
and U7248 (N_7248,N_7046,N_7051);
and U7249 (N_7249,N_7017,N_7173);
nor U7250 (N_7250,N_7148,N_7010);
or U7251 (N_7251,N_7091,N_7032);
and U7252 (N_7252,N_7086,N_7027);
or U7253 (N_7253,N_7074,N_7131);
xor U7254 (N_7254,N_7084,N_7168);
and U7255 (N_7255,N_7016,N_7140);
nor U7256 (N_7256,N_7113,N_7175);
and U7257 (N_7257,N_7170,N_7138);
or U7258 (N_7258,N_7164,N_7192);
and U7259 (N_7259,N_7059,N_7038);
xor U7260 (N_7260,N_7110,N_7042);
nand U7261 (N_7261,N_7114,N_7099);
nand U7262 (N_7262,N_7129,N_7157);
or U7263 (N_7263,N_7045,N_7156);
nor U7264 (N_7264,N_7019,N_7065);
xor U7265 (N_7265,N_7194,N_7057);
nor U7266 (N_7266,N_7166,N_7199);
xor U7267 (N_7267,N_7196,N_7165);
nor U7268 (N_7268,N_7154,N_7009);
and U7269 (N_7269,N_7124,N_7012);
xor U7270 (N_7270,N_7176,N_7061);
nand U7271 (N_7271,N_7101,N_7013);
nand U7272 (N_7272,N_7182,N_7185);
and U7273 (N_7273,N_7139,N_7070);
nor U7274 (N_7274,N_7120,N_7181);
and U7275 (N_7275,N_7143,N_7063);
or U7276 (N_7276,N_7087,N_7092);
xnor U7277 (N_7277,N_7158,N_7103);
nor U7278 (N_7278,N_7098,N_7094);
nand U7279 (N_7279,N_7146,N_7132);
nand U7280 (N_7280,N_7043,N_7137);
nor U7281 (N_7281,N_7044,N_7034);
nor U7282 (N_7282,N_7162,N_7026);
and U7283 (N_7283,N_7033,N_7108);
and U7284 (N_7284,N_7169,N_7105);
or U7285 (N_7285,N_7049,N_7075);
and U7286 (N_7286,N_7004,N_7088);
or U7287 (N_7287,N_7186,N_7163);
nand U7288 (N_7288,N_7121,N_7077);
nor U7289 (N_7289,N_7125,N_7064);
and U7290 (N_7290,N_7081,N_7149);
nor U7291 (N_7291,N_7000,N_7071);
or U7292 (N_7292,N_7190,N_7178);
or U7293 (N_7293,N_7025,N_7135);
nand U7294 (N_7294,N_7068,N_7085);
nor U7295 (N_7295,N_7147,N_7126);
nand U7296 (N_7296,N_7115,N_7011);
and U7297 (N_7297,N_7151,N_7030);
or U7298 (N_7298,N_7198,N_7029);
or U7299 (N_7299,N_7117,N_7150);
and U7300 (N_7300,N_7113,N_7100);
nor U7301 (N_7301,N_7061,N_7084);
or U7302 (N_7302,N_7118,N_7077);
or U7303 (N_7303,N_7070,N_7101);
nor U7304 (N_7304,N_7159,N_7107);
and U7305 (N_7305,N_7161,N_7085);
and U7306 (N_7306,N_7061,N_7161);
nand U7307 (N_7307,N_7193,N_7176);
or U7308 (N_7308,N_7001,N_7180);
nor U7309 (N_7309,N_7121,N_7067);
and U7310 (N_7310,N_7192,N_7089);
nand U7311 (N_7311,N_7107,N_7076);
or U7312 (N_7312,N_7155,N_7025);
xnor U7313 (N_7313,N_7189,N_7023);
xnor U7314 (N_7314,N_7178,N_7129);
nor U7315 (N_7315,N_7097,N_7100);
xnor U7316 (N_7316,N_7061,N_7175);
or U7317 (N_7317,N_7036,N_7135);
or U7318 (N_7318,N_7042,N_7004);
nor U7319 (N_7319,N_7020,N_7098);
xnor U7320 (N_7320,N_7021,N_7030);
nor U7321 (N_7321,N_7114,N_7102);
nand U7322 (N_7322,N_7096,N_7055);
or U7323 (N_7323,N_7091,N_7040);
xor U7324 (N_7324,N_7147,N_7114);
nor U7325 (N_7325,N_7100,N_7062);
nand U7326 (N_7326,N_7164,N_7187);
xnor U7327 (N_7327,N_7116,N_7142);
nand U7328 (N_7328,N_7188,N_7033);
nand U7329 (N_7329,N_7046,N_7057);
nand U7330 (N_7330,N_7077,N_7060);
nor U7331 (N_7331,N_7087,N_7031);
xnor U7332 (N_7332,N_7054,N_7149);
and U7333 (N_7333,N_7032,N_7082);
or U7334 (N_7334,N_7100,N_7044);
xnor U7335 (N_7335,N_7164,N_7160);
and U7336 (N_7336,N_7145,N_7151);
nand U7337 (N_7337,N_7060,N_7199);
nand U7338 (N_7338,N_7172,N_7100);
or U7339 (N_7339,N_7187,N_7098);
nor U7340 (N_7340,N_7124,N_7153);
and U7341 (N_7341,N_7018,N_7121);
xnor U7342 (N_7342,N_7114,N_7003);
xor U7343 (N_7343,N_7093,N_7159);
and U7344 (N_7344,N_7009,N_7182);
nor U7345 (N_7345,N_7085,N_7032);
xor U7346 (N_7346,N_7000,N_7075);
and U7347 (N_7347,N_7012,N_7003);
xor U7348 (N_7348,N_7032,N_7138);
or U7349 (N_7349,N_7184,N_7092);
xnor U7350 (N_7350,N_7021,N_7132);
xor U7351 (N_7351,N_7111,N_7139);
xnor U7352 (N_7352,N_7174,N_7050);
and U7353 (N_7353,N_7075,N_7031);
nand U7354 (N_7354,N_7165,N_7193);
xnor U7355 (N_7355,N_7098,N_7181);
or U7356 (N_7356,N_7019,N_7022);
nor U7357 (N_7357,N_7081,N_7080);
nand U7358 (N_7358,N_7052,N_7095);
nand U7359 (N_7359,N_7148,N_7054);
nor U7360 (N_7360,N_7176,N_7144);
nor U7361 (N_7361,N_7108,N_7162);
xor U7362 (N_7362,N_7149,N_7005);
or U7363 (N_7363,N_7010,N_7144);
nand U7364 (N_7364,N_7091,N_7105);
nor U7365 (N_7365,N_7136,N_7087);
and U7366 (N_7366,N_7081,N_7045);
xnor U7367 (N_7367,N_7061,N_7128);
and U7368 (N_7368,N_7158,N_7145);
nor U7369 (N_7369,N_7025,N_7080);
nor U7370 (N_7370,N_7180,N_7058);
and U7371 (N_7371,N_7047,N_7171);
or U7372 (N_7372,N_7109,N_7032);
nand U7373 (N_7373,N_7044,N_7054);
nor U7374 (N_7374,N_7020,N_7008);
or U7375 (N_7375,N_7078,N_7100);
nor U7376 (N_7376,N_7175,N_7130);
and U7377 (N_7377,N_7077,N_7116);
nand U7378 (N_7378,N_7086,N_7054);
or U7379 (N_7379,N_7065,N_7161);
xor U7380 (N_7380,N_7126,N_7030);
nand U7381 (N_7381,N_7009,N_7140);
nand U7382 (N_7382,N_7024,N_7143);
nand U7383 (N_7383,N_7009,N_7113);
and U7384 (N_7384,N_7030,N_7159);
nand U7385 (N_7385,N_7196,N_7132);
nor U7386 (N_7386,N_7047,N_7050);
or U7387 (N_7387,N_7061,N_7115);
xnor U7388 (N_7388,N_7172,N_7193);
nor U7389 (N_7389,N_7026,N_7167);
nand U7390 (N_7390,N_7198,N_7127);
and U7391 (N_7391,N_7046,N_7184);
and U7392 (N_7392,N_7180,N_7197);
xnor U7393 (N_7393,N_7031,N_7166);
and U7394 (N_7394,N_7054,N_7059);
or U7395 (N_7395,N_7038,N_7139);
xnor U7396 (N_7396,N_7052,N_7126);
and U7397 (N_7397,N_7177,N_7171);
nand U7398 (N_7398,N_7184,N_7130);
xor U7399 (N_7399,N_7033,N_7026);
xor U7400 (N_7400,N_7243,N_7300);
xor U7401 (N_7401,N_7214,N_7384);
nor U7402 (N_7402,N_7237,N_7268);
or U7403 (N_7403,N_7219,N_7335);
nand U7404 (N_7404,N_7336,N_7211);
or U7405 (N_7405,N_7210,N_7275);
or U7406 (N_7406,N_7235,N_7390);
nand U7407 (N_7407,N_7303,N_7256);
and U7408 (N_7408,N_7247,N_7231);
or U7409 (N_7409,N_7249,N_7254);
or U7410 (N_7410,N_7397,N_7362);
xnor U7411 (N_7411,N_7216,N_7332);
xor U7412 (N_7412,N_7307,N_7244);
and U7413 (N_7413,N_7264,N_7358);
or U7414 (N_7414,N_7238,N_7343);
xor U7415 (N_7415,N_7273,N_7392);
nand U7416 (N_7416,N_7215,N_7274);
xor U7417 (N_7417,N_7355,N_7338);
or U7418 (N_7418,N_7224,N_7360);
xnor U7419 (N_7419,N_7262,N_7333);
or U7420 (N_7420,N_7290,N_7346);
nor U7421 (N_7421,N_7311,N_7318);
and U7422 (N_7422,N_7341,N_7283);
or U7423 (N_7423,N_7316,N_7351);
or U7424 (N_7424,N_7205,N_7320);
nand U7425 (N_7425,N_7385,N_7323);
and U7426 (N_7426,N_7242,N_7306);
xnor U7427 (N_7427,N_7310,N_7302);
xnor U7428 (N_7428,N_7329,N_7291);
nand U7429 (N_7429,N_7348,N_7387);
nor U7430 (N_7430,N_7255,N_7299);
xnor U7431 (N_7431,N_7276,N_7269);
xnor U7432 (N_7432,N_7296,N_7218);
or U7433 (N_7433,N_7202,N_7361);
or U7434 (N_7434,N_7277,N_7271);
and U7435 (N_7435,N_7378,N_7293);
nor U7436 (N_7436,N_7380,N_7305);
nand U7437 (N_7437,N_7353,N_7394);
xnor U7438 (N_7438,N_7337,N_7388);
nand U7439 (N_7439,N_7373,N_7261);
or U7440 (N_7440,N_7280,N_7233);
or U7441 (N_7441,N_7201,N_7294);
xnor U7442 (N_7442,N_7288,N_7344);
nor U7443 (N_7443,N_7399,N_7395);
xnor U7444 (N_7444,N_7327,N_7374);
nand U7445 (N_7445,N_7315,N_7354);
nor U7446 (N_7446,N_7286,N_7213);
and U7447 (N_7447,N_7364,N_7228);
xor U7448 (N_7448,N_7350,N_7356);
xor U7449 (N_7449,N_7357,N_7270);
xnor U7450 (N_7450,N_7321,N_7207);
nor U7451 (N_7451,N_7345,N_7248);
nand U7452 (N_7452,N_7314,N_7295);
nor U7453 (N_7453,N_7232,N_7381);
nand U7454 (N_7454,N_7279,N_7375);
nand U7455 (N_7455,N_7372,N_7209);
nor U7456 (N_7456,N_7206,N_7366);
and U7457 (N_7457,N_7227,N_7204);
nand U7458 (N_7458,N_7221,N_7250);
nor U7459 (N_7459,N_7347,N_7339);
xnor U7460 (N_7460,N_7257,N_7222);
and U7461 (N_7461,N_7359,N_7379);
xor U7462 (N_7462,N_7229,N_7342);
nand U7463 (N_7463,N_7317,N_7251);
and U7464 (N_7464,N_7308,N_7284);
xor U7465 (N_7465,N_7259,N_7328);
xor U7466 (N_7466,N_7234,N_7241);
xor U7467 (N_7467,N_7282,N_7309);
nor U7468 (N_7468,N_7278,N_7340);
nor U7469 (N_7469,N_7368,N_7253);
or U7470 (N_7470,N_7263,N_7292);
nand U7471 (N_7471,N_7217,N_7312);
nor U7472 (N_7472,N_7246,N_7304);
or U7473 (N_7473,N_7230,N_7225);
and U7474 (N_7474,N_7200,N_7363);
nand U7475 (N_7475,N_7391,N_7301);
nand U7476 (N_7476,N_7377,N_7371);
nor U7477 (N_7477,N_7240,N_7331);
and U7478 (N_7478,N_7349,N_7365);
xor U7479 (N_7479,N_7245,N_7326);
or U7480 (N_7480,N_7386,N_7239);
nand U7481 (N_7481,N_7298,N_7252);
or U7482 (N_7482,N_7226,N_7212);
nor U7483 (N_7483,N_7367,N_7370);
and U7484 (N_7484,N_7398,N_7383);
nor U7485 (N_7485,N_7260,N_7334);
or U7486 (N_7486,N_7297,N_7382);
or U7487 (N_7487,N_7287,N_7267);
and U7488 (N_7488,N_7208,N_7223);
or U7489 (N_7489,N_7396,N_7285);
nor U7490 (N_7490,N_7324,N_7313);
nand U7491 (N_7491,N_7319,N_7330);
or U7492 (N_7492,N_7236,N_7322);
xor U7493 (N_7493,N_7220,N_7272);
and U7494 (N_7494,N_7266,N_7393);
and U7495 (N_7495,N_7389,N_7352);
xor U7496 (N_7496,N_7325,N_7281);
xor U7497 (N_7497,N_7289,N_7376);
or U7498 (N_7498,N_7265,N_7258);
xnor U7499 (N_7499,N_7369,N_7203);
and U7500 (N_7500,N_7358,N_7346);
or U7501 (N_7501,N_7210,N_7228);
nand U7502 (N_7502,N_7246,N_7253);
nand U7503 (N_7503,N_7378,N_7261);
nand U7504 (N_7504,N_7237,N_7340);
nand U7505 (N_7505,N_7248,N_7336);
nand U7506 (N_7506,N_7358,N_7301);
xor U7507 (N_7507,N_7221,N_7280);
or U7508 (N_7508,N_7340,N_7351);
or U7509 (N_7509,N_7279,N_7205);
xnor U7510 (N_7510,N_7396,N_7235);
nand U7511 (N_7511,N_7264,N_7282);
nor U7512 (N_7512,N_7310,N_7206);
or U7513 (N_7513,N_7298,N_7347);
and U7514 (N_7514,N_7317,N_7337);
nand U7515 (N_7515,N_7204,N_7286);
xor U7516 (N_7516,N_7263,N_7329);
xor U7517 (N_7517,N_7322,N_7217);
xor U7518 (N_7518,N_7269,N_7327);
nand U7519 (N_7519,N_7224,N_7251);
and U7520 (N_7520,N_7308,N_7346);
nor U7521 (N_7521,N_7308,N_7297);
nand U7522 (N_7522,N_7315,N_7259);
and U7523 (N_7523,N_7225,N_7201);
nor U7524 (N_7524,N_7214,N_7294);
xor U7525 (N_7525,N_7388,N_7307);
nor U7526 (N_7526,N_7295,N_7364);
xnor U7527 (N_7527,N_7211,N_7397);
nor U7528 (N_7528,N_7380,N_7222);
or U7529 (N_7529,N_7331,N_7243);
nand U7530 (N_7530,N_7200,N_7279);
xnor U7531 (N_7531,N_7274,N_7334);
nor U7532 (N_7532,N_7219,N_7286);
or U7533 (N_7533,N_7317,N_7306);
xnor U7534 (N_7534,N_7206,N_7372);
nor U7535 (N_7535,N_7354,N_7202);
nor U7536 (N_7536,N_7218,N_7316);
nor U7537 (N_7537,N_7249,N_7341);
xor U7538 (N_7538,N_7379,N_7314);
nor U7539 (N_7539,N_7340,N_7376);
nand U7540 (N_7540,N_7212,N_7275);
nand U7541 (N_7541,N_7208,N_7322);
nor U7542 (N_7542,N_7264,N_7351);
nand U7543 (N_7543,N_7239,N_7361);
and U7544 (N_7544,N_7284,N_7365);
and U7545 (N_7545,N_7309,N_7344);
and U7546 (N_7546,N_7264,N_7288);
nand U7547 (N_7547,N_7311,N_7230);
or U7548 (N_7548,N_7321,N_7384);
xnor U7549 (N_7549,N_7367,N_7227);
or U7550 (N_7550,N_7254,N_7270);
and U7551 (N_7551,N_7210,N_7376);
nand U7552 (N_7552,N_7348,N_7322);
and U7553 (N_7553,N_7312,N_7282);
nand U7554 (N_7554,N_7245,N_7369);
nand U7555 (N_7555,N_7225,N_7369);
or U7556 (N_7556,N_7271,N_7261);
xnor U7557 (N_7557,N_7271,N_7349);
nor U7558 (N_7558,N_7395,N_7321);
nor U7559 (N_7559,N_7241,N_7360);
and U7560 (N_7560,N_7248,N_7363);
nand U7561 (N_7561,N_7226,N_7202);
nand U7562 (N_7562,N_7294,N_7337);
and U7563 (N_7563,N_7224,N_7274);
xnor U7564 (N_7564,N_7268,N_7316);
nor U7565 (N_7565,N_7390,N_7249);
and U7566 (N_7566,N_7215,N_7279);
xnor U7567 (N_7567,N_7366,N_7225);
nor U7568 (N_7568,N_7236,N_7244);
nand U7569 (N_7569,N_7355,N_7361);
or U7570 (N_7570,N_7201,N_7208);
xnor U7571 (N_7571,N_7281,N_7330);
nor U7572 (N_7572,N_7381,N_7216);
xor U7573 (N_7573,N_7253,N_7309);
nor U7574 (N_7574,N_7298,N_7291);
and U7575 (N_7575,N_7211,N_7213);
or U7576 (N_7576,N_7354,N_7259);
nor U7577 (N_7577,N_7336,N_7390);
xor U7578 (N_7578,N_7379,N_7241);
or U7579 (N_7579,N_7302,N_7307);
nor U7580 (N_7580,N_7363,N_7278);
nor U7581 (N_7581,N_7228,N_7257);
nand U7582 (N_7582,N_7354,N_7226);
nor U7583 (N_7583,N_7374,N_7261);
and U7584 (N_7584,N_7253,N_7270);
nor U7585 (N_7585,N_7379,N_7254);
or U7586 (N_7586,N_7295,N_7221);
xor U7587 (N_7587,N_7303,N_7311);
xnor U7588 (N_7588,N_7314,N_7275);
nor U7589 (N_7589,N_7204,N_7256);
and U7590 (N_7590,N_7214,N_7351);
nor U7591 (N_7591,N_7394,N_7354);
nand U7592 (N_7592,N_7312,N_7229);
and U7593 (N_7593,N_7210,N_7248);
or U7594 (N_7594,N_7235,N_7387);
nand U7595 (N_7595,N_7361,N_7382);
and U7596 (N_7596,N_7302,N_7261);
xor U7597 (N_7597,N_7294,N_7393);
nand U7598 (N_7598,N_7210,N_7254);
nand U7599 (N_7599,N_7286,N_7340);
nand U7600 (N_7600,N_7424,N_7450);
nor U7601 (N_7601,N_7407,N_7533);
and U7602 (N_7602,N_7472,N_7421);
nor U7603 (N_7603,N_7556,N_7491);
xnor U7604 (N_7604,N_7546,N_7591);
nor U7605 (N_7605,N_7587,N_7578);
or U7606 (N_7606,N_7436,N_7518);
or U7607 (N_7607,N_7457,N_7559);
xor U7608 (N_7608,N_7554,N_7530);
xnor U7609 (N_7609,N_7400,N_7401);
nand U7610 (N_7610,N_7418,N_7557);
xnor U7611 (N_7611,N_7566,N_7583);
nand U7612 (N_7612,N_7465,N_7456);
and U7613 (N_7613,N_7506,N_7464);
nand U7614 (N_7614,N_7505,N_7597);
nor U7615 (N_7615,N_7434,N_7453);
nor U7616 (N_7616,N_7598,N_7416);
nand U7617 (N_7617,N_7480,N_7510);
nor U7618 (N_7618,N_7543,N_7599);
xor U7619 (N_7619,N_7443,N_7479);
xor U7620 (N_7620,N_7575,N_7516);
or U7621 (N_7621,N_7414,N_7590);
nor U7622 (N_7622,N_7417,N_7425);
and U7623 (N_7623,N_7439,N_7489);
and U7624 (N_7624,N_7511,N_7487);
nand U7625 (N_7625,N_7573,N_7508);
or U7626 (N_7626,N_7405,N_7455);
nand U7627 (N_7627,N_7492,N_7521);
nor U7628 (N_7628,N_7515,N_7523);
and U7629 (N_7629,N_7474,N_7551);
nor U7630 (N_7630,N_7589,N_7576);
or U7631 (N_7631,N_7481,N_7477);
xor U7632 (N_7632,N_7545,N_7519);
nand U7633 (N_7633,N_7475,N_7503);
xnor U7634 (N_7634,N_7524,N_7529);
or U7635 (N_7635,N_7577,N_7442);
xor U7636 (N_7636,N_7486,N_7494);
xor U7637 (N_7637,N_7541,N_7446);
nor U7638 (N_7638,N_7447,N_7413);
and U7639 (N_7639,N_7570,N_7544);
nand U7640 (N_7640,N_7565,N_7520);
xor U7641 (N_7641,N_7476,N_7579);
nand U7642 (N_7642,N_7538,N_7540);
and U7643 (N_7643,N_7504,N_7430);
and U7644 (N_7644,N_7493,N_7558);
and U7645 (N_7645,N_7572,N_7444);
xnor U7646 (N_7646,N_7502,N_7466);
nor U7647 (N_7647,N_7470,N_7488);
and U7648 (N_7648,N_7406,N_7592);
and U7649 (N_7649,N_7468,N_7451);
nor U7650 (N_7650,N_7426,N_7564);
nor U7651 (N_7651,N_7408,N_7484);
xor U7652 (N_7652,N_7452,N_7458);
nand U7653 (N_7653,N_7526,N_7478);
xor U7654 (N_7654,N_7482,N_7500);
nor U7655 (N_7655,N_7422,N_7582);
xnor U7656 (N_7656,N_7548,N_7563);
nand U7657 (N_7657,N_7496,N_7420);
nand U7658 (N_7658,N_7527,N_7509);
xor U7659 (N_7659,N_7550,N_7586);
or U7660 (N_7660,N_7460,N_7445);
or U7661 (N_7661,N_7483,N_7534);
nor U7662 (N_7662,N_7459,N_7435);
nor U7663 (N_7663,N_7471,N_7410);
and U7664 (N_7664,N_7448,N_7469);
nand U7665 (N_7665,N_7549,N_7402);
nor U7666 (N_7666,N_7580,N_7507);
nor U7667 (N_7667,N_7498,N_7404);
or U7668 (N_7668,N_7585,N_7522);
and U7669 (N_7669,N_7594,N_7454);
or U7670 (N_7670,N_7553,N_7428);
xor U7671 (N_7671,N_7595,N_7539);
or U7672 (N_7672,N_7432,N_7412);
xnor U7673 (N_7673,N_7461,N_7429);
xor U7674 (N_7674,N_7449,N_7490);
or U7675 (N_7675,N_7513,N_7552);
and U7676 (N_7676,N_7581,N_7467);
or U7677 (N_7677,N_7473,N_7441);
or U7678 (N_7678,N_7562,N_7512);
nand U7679 (N_7679,N_7588,N_7532);
nand U7680 (N_7680,N_7537,N_7463);
and U7681 (N_7681,N_7497,N_7517);
or U7682 (N_7682,N_7568,N_7561);
and U7683 (N_7683,N_7499,N_7462);
and U7684 (N_7684,N_7584,N_7571);
nor U7685 (N_7685,N_7409,N_7531);
nor U7686 (N_7686,N_7593,N_7431);
and U7687 (N_7687,N_7433,N_7536);
xor U7688 (N_7688,N_7485,N_7542);
and U7689 (N_7689,N_7437,N_7440);
nor U7690 (N_7690,N_7501,N_7415);
nor U7691 (N_7691,N_7495,N_7569);
and U7692 (N_7692,N_7528,N_7403);
and U7693 (N_7693,N_7411,N_7427);
xnor U7694 (N_7694,N_7535,N_7419);
and U7695 (N_7695,N_7525,N_7438);
nor U7696 (N_7696,N_7567,N_7555);
or U7697 (N_7697,N_7423,N_7574);
and U7698 (N_7698,N_7560,N_7596);
nand U7699 (N_7699,N_7547,N_7514);
and U7700 (N_7700,N_7510,N_7522);
nand U7701 (N_7701,N_7443,N_7532);
or U7702 (N_7702,N_7503,N_7494);
or U7703 (N_7703,N_7537,N_7528);
nand U7704 (N_7704,N_7545,N_7439);
and U7705 (N_7705,N_7469,N_7416);
nor U7706 (N_7706,N_7566,N_7560);
or U7707 (N_7707,N_7428,N_7517);
or U7708 (N_7708,N_7493,N_7454);
nor U7709 (N_7709,N_7458,N_7480);
or U7710 (N_7710,N_7577,N_7419);
nor U7711 (N_7711,N_7507,N_7530);
nand U7712 (N_7712,N_7545,N_7465);
xor U7713 (N_7713,N_7458,N_7424);
nand U7714 (N_7714,N_7536,N_7574);
or U7715 (N_7715,N_7511,N_7537);
or U7716 (N_7716,N_7423,N_7447);
nor U7717 (N_7717,N_7558,N_7560);
xnor U7718 (N_7718,N_7434,N_7420);
nor U7719 (N_7719,N_7591,N_7405);
xor U7720 (N_7720,N_7485,N_7511);
nand U7721 (N_7721,N_7525,N_7460);
and U7722 (N_7722,N_7421,N_7490);
xor U7723 (N_7723,N_7581,N_7527);
nand U7724 (N_7724,N_7594,N_7514);
nor U7725 (N_7725,N_7490,N_7545);
nor U7726 (N_7726,N_7514,N_7596);
nand U7727 (N_7727,N_7580,N_7499);
and U7728 (N_7728,N_7538,N_7499);
or U7729 (N_7729,N_7542,N_7506);
nand U7730 (N_7730,N_7462,N_7596);
xnor U7731 (N_7731,N_7532,N_7516);
nor U7732 (N_7732,N_7493,N_7540);
nor U7733 (N_7733,N_7487,N_7496);
nand U7734 (N_7734,N_7494,N_7591);
or U7735 (N_7735,N_7475,N_7505);
nor U7736 (N_7736,N_7560,N_7595);
nand U7737 (N_7737,N_7559,N_7413);
nand U7738 (N_7738,N_7445,N_7567);
xor U7739 (N_7739,N_7528,N_7569);
nand U7740 (N_7740,N_7565,N_7525);
xnor U7741 (N_7741,N_7489,N_7449);
xor U7742 (N_7742,N_7507,N_7587);
nor U7743 (N_7743,N_7530,N_7504);
xnor U7744 (N_7744,N_7471,N_7445);
or U7745 (N_7745,N_7444,N_7533);
or U7746 (N_7746,N_7444,N_7496);
and U7747 (N_7747,N_7410,N_7546);
xnor U7748 (N_7748,N_7492,N_7443);
nor U7749 (N_7749,N_7467,N_7528);
and U7750 (N_7750,N_7476,N_7454);
xor U7751 (N_7751,N_7437,N_7413);
and U7752 (N_7752,N_7568,N_7424);
and U7753 (N_7753,N_7507,N_7440);
and U7754 (N_7754,N_7551,N_7409);
xor U7755 (N_7755,N_7410,N_7541);
nand U7756 (N_7756,N_7523,N_7521);
xor U7757 (N_7757,N_7502,N_7405);
nor U7758 (N_7758,N_7428,N_7429);
xnor U7759 (N_7759,N_7539,N_7432);
nand U7760 (N_7760,N_7469,N_7543);
nor U7761 (N_7761,N_7436,N_7574);
nand U7762 (N_7762,N_7446,N_7521);
and U7763 (N_7763,N_7577,N_7523);
nor U7764 (N_7764,N_7486,N_7559);
xor U7765 (N_7765,N_7563,N_7440);
xnor U7766 (N_7766,N_7428,N_7439);
nand U7767 (N_7767,N_7406,N_7441);
nand U7768 (N_7768,N_7509,N_7474);
or U7769 (N_7769,N_7539,N_7463);
xor U7770 (N_7770,N_7537,N_7434);
or U7771 (N_7771,N_7547,N_7402);
nor U7772 (N_7772,N_7464,N_7493);
nand U7773 (N_7773,N_7516,N_7413);
nor U7774 (N_7774,N_7585,N_7485);
nor U7775 (N_7775,N_7534,N_7566);
and U7776 (N_7776,N_7402,N_7532);
xor U7777 (N_7777,N_7483,N_7422);
or U7778 (N_7778,N_7557,N_7408);
nand U7779 (N_7779,N_7405,N_7529);
xor U7780 (N_7780,N_7440,N_7431);
nand U7781 (N_7781,N_7513,N_7459);
or U7782 (N_7782,N_7407,N_7563);
xnor U7783 (N_7783,N_7543,N_7418);
or U7784 (N_7784,N_7559,N_7541);
xor U7785 (N_7785,N_7544,N_7572);
or U7786 (N_7786,N_7571,N_7567);
xnor U7787 (N_7787,N_7560,N_7562);
xor U7788 (N_7788,N_7531,N_7532);
nand U7789 (N_7789,N_7504,N_7461);
or U7790 (N_7790,N_7412,N_7480);
xnor U7791 (N_7791,N_7488,N_7424);
nor U7792 (N_7792,N_7463,N_7461);
or U7793 (N_7793,N_7448,N_7516);
nand U7794 (N_7794,N_7448,N_7533);
nand U7795 (N_7795,N_7468,N_7569);
nor U7796 (N_7796,N_7545,N_7449);
and U7797 (N_7797,N_7417,N_7538);
or U7798 (N_7798,N_7464,N_7482);
nand U7799 (N_7799,N_7525,N_7597);
xnor U7800 (N_7800,N_7651,N_7628);
nand U7801 (N_7801,N_7629,N_7699);
xnor U7802 (N_7802,N_7691,N_7676);
nor U7803 (N_7803,N_7659,N_7734);
nor U7804 (N_7804,N_7793,N_7665);
or U7805 (N_7805,N_7606,N_7754);
or U7806 (N_7806,N_7695,N_7761);
nand U7807 (N_7807,N_7635,N_7716);
or U7808 (N_7808,N_7710,N_7786);
nor U7809 (N_7809,N_7681,N_7634);
xnor U7810 (N_7810,N_7742,N_7767);
nand U7811 (N_7811,N_7747,N_7748);
xnor U7812 (N_7812,N_7608,N_7631);
and U7813 (N_7813,N_7668,N_7610);
and U7814 (N_7814,N_7779,N_7797);
and U7815 (N_7815,N_7655,N_7702);
nand U7816 (N_7816,N_7660,N_7787);
nand U7817 (N_7817,N_7618,N_7639);
nand U7818 (N_7818,N_7724,N_7707);
nand U7819 (N_7819,N_7620,N_7649);
nor U7820 (N_7820,N_7648,N_7619);
nor U7821 (N_7821,N_7617,N_7791);
nor U7822 (N_7822,N_7693,N_7607);
xor U7823 (N_7823,N_7621,N_7763);
and U7824 (N_7824,N_7600,N_7687);
and U7825 (N_7825,N_7638,N_7614);
or U7826 (N_7826,N_7750,N_7769);
or U7827 (N_7827,N_7682,N_7753);
nor U7828 (N_7828,N_7664,N_7616);
and U7829 (N_7829,N_7774,N_7775);
nand U7830 (N_7830,N_7715,N_7626);
and U7831 (N_7831,N_7746,N_7794);
nand U7832 (N_7832,N_7719,N_7743);
or U7833 (N_7833,N_7661,N_7640);
nand U7834 (N_7834,N_7749,N_7788);
xnor U7835 (N_7835,N_7680,N_7784);
nand U7836 (N_7836,N_7611,N_7694);
nand U7837 (N_7837,N_7689,N_7677);
xor U7838 (N_7838,N_7632,N_7641);
and U7839 (N_7839,N_7789,N_7704);
or U7840 (N_7840,N_7765,N_7729);
and U7841 (N_7841,N_7674,N_7673);
nor U7842 (N_7842,N_7698,N_7782);
and U7843 (N_7843,N_7780,N_7727);
and U7844 (N_7844,N_7685,N_7633);
or U7845 (N_7845,N_7623,N_7609);
nand U7846 (N_7846,N_7714,N_7785);
and U7847 (N_7847,N_7656,N_7757);
nor U7848 (N_7848,N_7678,N_7650);
nor U7849 (N_7849,N_7652,N_7658);
or U7850 (N_7850,N_7790,N_7679);
xnor U7851 (N_7851,N_7718,N_7795);
xnor U7852 (N_7852,N_7603,N_7799);
nand U7853 (N_7853,N_7684,N_7736);
and U7854 (N_7854,N_7643,N_7770);
and U7855 (N_7855,N_7604,N_7733);
xor U7856 (N_7856,N_7613,N_7756);
and U7857 (N_7857,N_7692,N_7771);
nand U7858 (N_7858,N_7722,N_7705);
or U7859 (N_7859,N_7735,N_7624);
xnor U7860 (N_7860,N_7697,N_7706);
nand U7861 (N_7861,N_7745,N_7711);
nand U7862 (N_7862,N_7713,N_7657);
and U7863 (N_7863,N_7708,N_7764);
nor U7864 (N_7864,N_7671,N_7778);
xor U7865 (N_7865,N_7783,N_7726);
or U7866 (N_7866,N_7667,N_7696);
nand U7867 (N_7867,N_7712,N_7637);
nand U7868 (N_7868,N_7690,N_7653);
nand U7869 (N_7869,N_7602,N_7777);
nand U7870 (N_7870,N_7738,N_7737);
xnor U7871 (N_7871,N_7762,N_7636);
or U7872 (N_7872,N_7728,N_7796);
xor U7873 (N_7873,N_7672,N_7701);
nand U7874 (N_7874,N_7720,N_7776);
and U7875 (N_7875,N_7670,N_7751);
xnor U7876 (N_7876,N_7675,N_7612);
xor U7877 (N_7877,N_7615,N_7723);
and U7878 (N_7878,N_7683,N_7625);
nor U7879 (N_7879,N_7654,N_7798);
and U7880 (N_7880,N_7700,N_7663);
and U7881 (N_7881,N_7741,N_7646);
nor U7882 (N_7882,N_7666,N_7739);
and U7883 (N_7883,N_7755,N_7645);
nand U7884 (N_7884,N_7766,N_7744);
xor U7885 (N_7885,N_7647,N_7644);
nor U7886 (N_7886,N_7717,N_7703);
nor U7887 (N_7887,N_7630,N_7725);
nand U7888 (N_7888,N_7622,N_7601);
xnor U7889 (N_7889,N_7709,N_7721);
or U7890 (N_7890,N_7730,N_7792);
and U7891 (N_7891,N_7740,N_7773);
and U7892 (N_7892,N_7760,N_7662);
or U7893 (N_7893,N_7752,N_7759);
xor U7894 (N_7894,N_7605,N_7686);
nor U7895 (N_7895,N_7732,N_7768);
or U7896 (N_7896,N_7731,N_7772);
xor U7897 (N_7897,N_7688,N_7642);
nor U7898 (N_7898,N_7669,N_7781);
xnor U7899 (N_7899,N_7758,N_7627);
and U7900 (N_7900,N_7628,N_7749);
or U7901 (N_7901,N_7610,N_7666);
and U7902 (N_7902,N_7782,N_7613);
nor U7903 (N_7903,N_7763,N_7684);
xor U7904 (N_7904,N_7634,N_7642);
and U7905 (N_7905,N_7601,N_7671);
or U7906 (N_7906,N_7638,N_7741);
and U7907 (N_7907,N_7776,N_7621);
and U7908 (N_7908,N_7775,N_7696);
nor U7909 (N_7909,N_7781,N_7714);
nor U7910 (N_7910,N_7616,N_7677);
or U7911 (N_7911,N_7639,N_7798);
nor U7912 (N_7912,N_7664,N_7663);
xor U7913 (N_7913,N_7795,N_7711);
nor U7914 (N_7914,N_7751,N_7659);
or U7915 (N_7915,N_7700,N_7713);
xnor U7916 (N_7916,N_7656,N_7729);
and U7917 (N_7917,N_7674,N_7786);
or U7918 (N_7918,N_7687,N_7739);
or U7919 (N_7919,N_7630,N_7654);
nor U7920 (N_7920,N_7715,N_7789);
nand U7921 (N_7921,N_7723,N_7702);
nor U7922 (N_7922,N_7702,N_7706);
or U7923 (N_7923,N_7609,N_7790);
xnor U7924 (N_7924,N_7670,N_7715);
nor U7925 (N_7925,N_7666,N_7698);
nor U7926 (N_7926,N_7787,N_7798);
or U7927 (N_7927,N_7670,N_7764);
nor U7928 (N_7928,N_7650,N_7647);
xor U7929 (N_7929,N_7644,N_7751);
nand U7930 (N_7930,N_7742,N_7713);
nand U7931 (N_7931,N_7660,N_7618);
or U7932 (N_7932,N_7779,N_7761);
and U7933 (N_7933,N_7618,N_7727);
or U7934 (N_7934,N_7693,N_7761);
nand U7935 (N_7935,N_7657,N_7747);
nand U7936 (N_7936,N_7758,N_7628);
nand U7937 (N_7937,N_7673,N_7660);
nor U7938 (N_7938,N_7685,N_7605);
nand U7939 (N_7939,N_7652,N_7649);
nand U7940 (N_7940,N_7624,N_7680);
and U7941 (N_7941,N_7714,N_7713);
nand U7942 (N_7942,N_7716,N_7678);
nor U7943 (N_7943,N_7609,N_7712);
nor U7944 (N_7944,N_7675,N_7741);
xor U7945 (N_7945,N_7650,N_7602);
and U7946 (N_7946,N_7763,N_7667);
xor U7947 (N_7947,N_7740,N_7793);
nor U7948 (N_7948,N_7767,N_7666);
or U7949 (N_7949,N_7795,N_7631);
and U7950 (N_7950,N_7679,N_7612);
xnor U7951 (N_7951,N_7640,N_7606);
nand U7952 (N_7952,N_7655,N_7786);
or U7953 (N_7953,N_7648,N_7753);
and U7954 (N_7954,N_7786,N_7606);
xor U7955 (N_7955,N_7723,N_7634);
or U7956 (N_7956,N_7754,N_7740);
nor U7957 (N_7957,N_7613,N_7788);
nand U7958 (N_7958,N_7726,N_7685);
and U7959 (N_7959,N_7677,N_7727);
xnor U7960 (N_7960,N_7727,N_7659);
xnor U7961 (N_7961,N_7755,N_7658);
xor U7962 (N_7962,N_7796,N_7642);
or U7963 (N_7963,N_7689,N_7699);
or U7964 (N_7964,N_7602,N_7775);
and U7965 (N_7965,N_7777,N_7652);
nor U7966 (N_7966,N_7755,N_7656);
nor U7967 (N_7967,N_7660,N_7735);
xor U7968 (N_7968,N_7791,N_7771);
or U7969 (N_7969,N_7751,N_7648);
or U7970 (N_7970,N_7652,N_7686);
and U7971 (N_7971,N_7715,N_7777);
xnor U7972 (N_7972,N_7689,N_7759);
nor U7973 (N_7973,N_7764,N_7689);
nand U7974 (N_7974,N_7751,N_7797);
xor U7975 (N_7975,N_7770,N_7711);
nand U7976 (N_7976,N_7665,N_7620);
and U7977 (N_7977,N_7704,N_7780);
or U7978 (N_7978,N_7783,N_7612);
xor U7979 (N_7979,N_7607,N_7789);
xnor U7980 (N_7980,N_7642,N_7784);
xor U7981 (N_7981,N_7708,N_7660);
and U7982 (N_7982,N_7696,N_7706);
nand U7983 (N_7983,N_7745,N_7605);
and U7984 (N_7984,N_7778,N_7676);
or U7985 (N_7985,N_7605,N_7698);
nor U7986 (N_7986,N_7734,N_7664);
xor U7987 (N_7987,N_7782,N_7700);
xor U7988 (N_7988,N_7763,N_7776);
xor U7989 (N_7989,N_7783,N_7747);
and U7990 (N_7990,N_7741,N_7778);
nand U7991 (N_7991,N_7713,N_7724);
xnor U7992 (N_7992,N_7608,N_7772);
nor U7993 (N_7993,N_7640,N_7674);
and U7994 (N_7994,N_7788,N_7626);
nor U7995 (N_7995,N_7665,N_7710);
or U7996 (N_7996,N_7603,N_7713);
xor U7997 (N_7997,N_7691,N_7755);
nand U7998 (N_7998,N_7711,N_7659);
or U7999 (N_7999,N_7624,N_7798);
nand U8000 (N_8000,N_7860,N_7898);
or U8001 (N_8001,N_7980,N_7970);
xor U8002 (N_8002,N_7938,N_7988);
and U8003 (N_8003,N_7825,N_7866);
nor U8004 (N_8004,N_7909,N_7837);
and U8005 (N_8005,N_7829,N_7808);
nor U8006 (N_8006,N_7900,N_7977);
and U8007 (N_8007,N_7806,N_7946);
and U8008 (N_8008,N_7884,N_7819);
or U8009 (N_8009,N_7902,N_7992);
xnor U8010 (N_8010,N_7816,N_7960);
nand U8011 (N_8011,N_7892,N_7936);
and U8012 (N_8012,N_7879,N_7836);
nor U8013 (N_8013,N_7944,N_7858);
and U8014 (N_8014,N_7962,N_7958);
or U8015 (N_8015,N_7863,N_7887);
nand U8016 (N_8016,N_7993,N_7840);
or U8017 (N_8017,N_7928,N_7817);
nor U8018 (N_8018,N_7953,N_7971);
xor U8019 (N_8019,N_7846,N_7803);
xor U8020 (N_8020,N_7951,N_7838);
xor U8021 (N_8021,N_7824,N_7812);
xor U8022 (N_8022,N_7982,N_7845);
nor U8023 (N_8023,N_7901,N_7850);
and U8024 (N_8024,N_7875,N_7952);
and U8025 (N_8025,N_7888,N_7893);
xnor U8026 (N_8026,N_7922,N_7811);
xnor U8027 (N_8027,N_7800,N_7929);
nand U8028 (N_8028,N_7979,N_7990);
or U8029 (N_8029,N_7826,N_7853);
nand U8030 (N_8030,N_7986,N_7915);
or U8031 (N_8031,N_7882,N_7809);
and U8032 (N_8032,N_7984,N_7847);
and U8033 (N_8033,N_7823,N_7949);
xor U8034 (N_8034,N_7950,N_7868);
xor U8035 (N_8035,N_7849,N_7939);
nand U8036 (N_8036,N_7947,N_7923);
nor U8037 (N_8037,N_7839,N_7930);
nor U8038 (N_8038,N_7996,N_7967);
nand U8039 (N_8039,N_7942,N_7885);
or U8040 (N_8040,N_7999,N_7802);
or U8041 (N_8041,N_7896,N_7918);
or U8042 (N_8042,N_7961,N_7869);
and U8043 (N_8043,N_7865,N_7818);
or U8044 (N_8044,N_7924,N_7919);
or U8045 (N_8045,N_7920,N_7855);
or U8046 (N_8046,N_7877,N_7981);
nor U8047 (N_8047,N_7859,N_7976);
nand U8048 (N_8048,N_7948,N_7903);
xnor U8049 (N_8049,N_7910,N_7821);
nand U8050 (N_8050,N_7932,N_7810);
or U8051 (N_8051,N_7881,N_7842);
xnor U8052 (N_8052,N_7973,N_7978);
and U8053 (N_8053,N_7956,N_7974);
nor U8054 (N_8054,N_7911,N_7983);
nor U8055 (N_8055,N_7876,N_7874);
nor U8056 (N_8056,N_7880,N_7916);
nand U8057 (N_8057,N_7886,N_7943);
or U8058 (N_8058,N_7895,N_7987);
and U8059 (N_8059,N_7832,N_7995);
nand U8060 (N_8060,N_7890,N_7854);
nor U8061 (N_8061,N_7989,N_7841);
or U8062 (N_8062,N_7934,N_7872);
or U8063 (N_8063,N_7985,N_7921);
or U8064 (N_8064,N_7965,N_7937);
or U8065 (N_8065,N_7926,N_7856);
or U8066 (N_8066,N_7870,N_7975);
nor U8067 (N_8067,N_7864,N_7807);
nor U8068 (N_8068,N_7899,N_7964);
xnor U8069 (N_8069,N_7871,N_7966);
nor U8070 (N_8070,N_7827,N_7933);
nor U8071 (N_8071,N_7907,N_7941);
and U8072 (N_8072,N_7830,N_7843);
xnor U8073 (N_8073,N_7867,N_7955);
nor U8074 (N_8074,N_7908,N_7891);
or U8075 (N_8075,N_7894,N_7844);
nor U8076 (N_8076,N_7805,N_7997);
nor U8077 (N_8077,N_7904,N_7857);
and U8078 (N_8078,N_7889,N_7852);
nor U8079 (N_8079,N_7862,N_7834);
nor U8080 (N_8080,N_7972,N_7814);
nor U8081 (N_8081,N_7851,N_7905);
nand U8082 (N_8082,N_7912,N_7940);
and U8083 (N_8083,N_7927,N_7991);
or U8084 (N_8084,N_7813,N_7968);
and U8085 (N_8085,N_7848,N_7820);
or U8086 (N_8086,N_7931,N_7917);
nor U8087 (N_8087,N_7801,N_7994);
and U8088 (N_8088,N_7913,N_7897);
nor U8089 (N_8089,N_7833,N_7861);
nor U8090 (N_8090,N_7954,N_7959);
and U8091 (N_8091,N_7878,N_7963);
and U8092 (N_8092,N_7831,N_7914);
or U8093 (N_8093,N_7969,N_7935);
nor U8094 (N_8094,N_7957,N_7822);
nor U8095 (N_8095,N_7804,N_7873);
xor U8096 (N_8096,N_7906,N_7945);
nor U8097 (N_8097,N_7835,N_7883);
nand U8098 (N_8098,N_7925,N_7828);
xnor U8099 (N_8099,N_7998,N_7815);
or U8100 (N_8100,N_7966,N_7919);
nor U8101 (N_8101,N_7848,N_7950);
nor U8102 (N_8102,N_7862,N_7886);
xnor U8103 (N_8103,N_7829,N_7831);
or U8104 (N_8104,N_7969,N_7954);
or U8105 (N_8105,N_7853,N_7986);
nor U8106 (N_8106,N_7863,N_7804);
or U8107 (N_8107,N_7902,N_7980);
or U8108 (N_8108,N_7919,N_7898);
and U8109 (N_8109,N_7877,N_7832);
nor U8110 (N_8110,N_7963,N_7881);
nand U8111 (N_8111,N_7916,N_7971);
and U8112 (N_8112,N_7880,N_7818);
and U8113 (N_8113,N_7953,N_7876);
or U8114 (N_8114,N_7924,N_7816);
xor U8115 (N_8115,N_7833,N_7912);
xnor U8116 (N_8116,N_7843,N_7882);
xor U8117 (N_8117,N_7803,N_7850);
or U8118 (N_8118,N_7972,N_7847);
and U8119 (N_8119,N_7811,N_7812);
or U8120 (N_8120,N_7901,N_7810);
xnor U8121 (N_8121,N_7985,N_7849);
xnor U8122 (N_8122,N_7932,N_7888);
or U8123 (N_8123,N_7993,N_7889);
and U8124 (N_8124,N_7866,N_7818);
nand U8125 (N_8125,N_7858,N_7849);
and U8126 (N_8126,N_7930,N_7910);
and U8127 (N_8127,N_7868,N_7928);
nand U8128 (N_8128,N_7844,N_7831);
or U8129 (N_8129,N_7941,N_7843);
xor U8130 (N_8130,N_7985,N_7868);
and U8131 (N_8131,N_7915,N_7987);
nor U8132 (N_8132,N_7997,N_7828);
and U8133 (N_8133,N_7874,N_7823);
or U8134 (N_8134,N_7840,N_7934);
nand U8135 (N_8135,N_7986,N_7814);
and U8136 (N_8136,N_7805,N_7962);
or U8137 (N_8137,N_7971,N_7940);
nor U8138 (N_8138,N_7819,N_7860);
or U8139 (N_8139,N_7885,N_7814);
nand U8140 (N_8140,N_7912,N_7904);
and U8141 (N_8141,N_7821,N_7917);
nand U8142 (N_8142,N_7919,N_7930);
or U8143 (N_8143,N_7866,N_7885);
or U8144 (N_8144,N_7813,N_7956);
or U8145 (N_8145,N_7818,N_7910);
nand U8146 (N_8146,N_7968,N_7999);
nand U8147 (N_8147,N_7962,N_7860);
nor U8148 (N_8148,N_7871,N_7896);
and U8149 (N_8149,N_7902,N_7874);
nand U8150 (N_8150,N_7902,N_7852);
nor U8151 (N_8151,N_7878,N_7887);
or U8152 (N_8152,N_7948,N_7826);
xor U8153 (N_8153,N_7824,N_7813);
or U8154 (N_8154,N_7938,N_7819);
and U8155 (N_8155,N_7862,N_7804);
nand U8156 (N_8156,N_7866,N_7838);
or U8157 (N_8157,N_7856,N_7950);
nand U8158 (N_8158,N_7844,N_7974);
or U8159 (N_8159,N_7872,N_7949);
or U8160 (N_8160,N_7903,N_7853);
nor U8161 (N_8161,N_7906,N_7848);
or U8162 (N_8162,N_7943,N_7809);
or U8163 (N_8163,N_7948,N_7842);
nand U8164 (N_8164,N_7989,N_7927);
nor U8165 (N_8165,N_7832,N_7923);
nor U8166 (N_8166,N_7822,N_7978);
nand U8167 (N_8167,N_7808,N_7873);
nand U8168 (N_8168,N_7935,N_7868);
and U8169 (N_8169,N_7800,N_7984);
xor U8170 (N_8170,N_7999,N_7915);
nand U8171 (N_8171,N_7891,N_7875);
nand U8172 (N_8172,N_7807,N_7835);
or U8173 (N_8173,N_7968,N_7833);
nand U8174 (N_8174,N_7979,N_7951);
or U8175 (N_8175,N_7944,N_7844);
xor U8176 (N_8176,N_7824,N_7818);
or U8177 (N_8177,N_7881,N_7891);
xnor U8178 (N_8178,N_7992,N_7883);
and U8179 (N_8179,N_7970,N_7883);
nor U8180 (N_8180,N_7963,N_7807);
and U8181 (N_8181,N_7903,N_7969);
or U8182 (N_8182,N_7825,N_7967);
and U8183 (N_8183,N_7809,N_7956);
or U8184 (N_8184,N_7945,N_7805);
or U8185 (N_8185,N_7819,N_7972);
and U8186 (N_8186,N_7976,N_7844);
and U8187 (N_8187,N_7930,N_7987);
or U8188 (N_8188,N_7917,N_7912);
xor U8189 (N_8189,N_7952,N_7971);
and U8190 (N_8190,N_7897,N_7867);
or U8191 (N_8191,N_7973,N_7860);
nand U8192 (N_8192,N_7917,N_7829);
xor U8193 (N_8193,N_7910,N_7847);
nor U8194 (N_8194,N_7979,N_7823);
or U8195 (N_8195,N_7945,N_7968);
or U8196 (N_8196,N_7915,N_7962);
xor U8197 (N_8197,N_7991,N_7829);
nor U8198 (N_8198,N_7930,N_7807);
or U8199 (N_8199,N_7910,N_7895);
or U8200 (N_8200,N_8026,N_8021);
xor U8201 (N_8201,N_8054,N_8086);
nand U8202 (N_8202,N_8074,N_8092);
nand U8203 (N_8203,N_8186,N_8046);
nand U8204 (N_8204,N_8047,N_8088);
nand U8205 (N_8205,N_8159,N_8121);
or U8206 (N_8206,N_8187,N_8083);
xnor U8207 (N_8207,N_8194,N_8037);
or U8208 (N_8208,N_8188,N_8031);
or U8209 (N_8209,N_8107,N_8003);
and U8210 (N_8210,N_8012,N_8087);
or U8211 (N_8211,N_8033,N_8096);
or U8212 (N_8212,N_8028,N_8075);
and U8213 (N_8213,N_8052,N_8103);
and U8214 (N_8214,N_8178,N_8111);
nor U8215 (N_8215,N_8167,N_8191);
nand U8216 (N_8216,N_8017,N_8179);
nand U8217 (N_8217,N_8155,N_8039);
and U8218 (N_8218,N_8129,N_8142);
nand U8219 (N_8219,N_8098,N_8141);
xnor U8220 (N_8220,N_8101,N_8170);
and U8221 (N_8221,N_8057,N_8114);
nand U8222 (N_8222,N_8135,N_8036);
xor U8223 (N_8223,N_8120,N_8064);
and U8224 (N_8224,N_8171,N_8070);
nor U8225 (N_8225,N_8174,N_8190);
and U8226 (N_8226,N_8065,N_8062);
and U8227 (N_8227,N_8177,N_8115);
nand U8228 (N_8228,N_8136,N_8061);
or U8229 (N_8229,N_8079,N_8069);
or U8230 (N_8230,N_8049,N_8175);
xor U8231 (N_8231,N_8143,N_8117);
xor U8232 (N_8232,N_8192,N_8160);
nor U8233 (N_8233,N_8063,N_8197);
and U8234 (N_8234,N_8108,N_8076);
nor U8235 (N_8235,N_8011,N_8055);
xor U8236 (N_8236,N_8004,N_8019);
or U8237 (N_8237,N_8007,N_8199);
or U8238 (N_8238,N_8176,N_8168);
xnor U8239 (N_8239,N_8072,N_8181);
nand U8240 (N_8240,N_8027,N_8035);
nand U8241 (N_8241,N_8193,N_8093);
nand U8242 (N_8242,N_8109,N_8158);
nor U8243 (N_8243,N_8034,N_8102);
nand U8244 (N_8244,N_8150,N_8131);
and U8245 (N_8245,N_8058,N_8038);
nand U8246 (N_8246,N_8060,N_8173);
and U8247 (N_8247,N_8022,N_8042);
and U8248 (N_8248,N_8156,N_8154);
and U8249 (N_8249,N_8094,N_8073);
nor U8250 (N_8250,N_8014,N_8163);
nor U8251 (N_8251,N_8009,N_8169);
nand U8252 (N_8252,N_8095,N_8104);
or U8253 (N_8253,N_8123,N_8008);
nand U8254 (N_8254,N_8133,N_8182);
nor U8255 (N_8255,N_8091,N_8016);
and U8256 (N_8256,N_8110,N_8081);
nand U8257 (N_8257,N_8068,N_8005);
nand U8258 (N_8258,N_8162,N_8151);
xnor U8259 (N_8259,N_8090,N_8097);
nand U8260 (N_8260,N_8024,N_8041);
or U8261 (N_8261,N_8124,N_8010);
xor U8262 (N_8262,N_8020,N_8001);
nand U8263 (N_8263,N_8180,N_8040);
xor U8264 (N_8264,N_8195,N_8185);
nor U8265 (N_8265,N_8126,N_8149);
nor U8266 (N_8266,N_8085,N_8018);
or U8267 (N_8267,N_8122,N_8144);
nor U8268 (N_8268,N_8147,N_8077);
xor U8269 (N_8269,N_8183,N_8113);
or U8270 (N_8270,N_8189,N_8153);
and U8271 (N_8271,N_8116,N_8099);
nand U8272 (N_8272,N_8148,N_8006);
or U8273 (N_8273,N_8196,N_8157);
nand U8274 (N_8274,N_8172,N_8050);
nand U8275 (N_8275,N_8165,N_8139);
nand U8276 (N_8276,N_8032,N_8128);
nand U8277 (N_8277,N_8130,N_8137);
xnor U8278 (N_8278,N_8084,N_8045);
xor U8279 (N_8279,N_8080,N_8112);
nor U8280 (N_8280,N_8198,N_8056);
nand U8281 (N_8281,N_8127,N_8089);
nor U8282 (N_8282,N_8043,N_8082);
and U8283 (N_8283,N_8138,N_8132);
and U8284 (N_8284,N_8152,N_8119);
nand U8285 (N_8285,N_8023,N_8053);
or U8286 (N_8286,N_8067,N_8161);
nor U8287 (N_8287,N_8166,N_8134);
and U8288 (N_8288,N_8100,N_8071);
xnor U8289 (N_8289,N_8015,N_8140);
nand U8290 (N_8290,N_8184,N_8106);
nor U8291 (N_8291,N_8000,N_8078);
and U8292 (N_8292,N_8145,N_8048);
or U8293 (N_8293,N_8002,N_8029);
and U8294 (N_8294,N_8118,N_8013);
and U8295 (N_8295,N_8051,N_8105);
xnor U8296 (N_8296,N_8059,N_8044);
or U8297 (N_8297,N_8066,N_8025);
nor U8298 (N_8298,N_8146,N_8030);
or U8299 (N_8299,N_8125,N_8164);
or U8300 (N_8300,N_8192,N_8184);
and U8301 (N_8301,N_8155,N_8150);
and U8302 (N_8302,N_8099,N_8095);
nand U8303 (N_8303,N_8072,N_8081);
or U8304 (N_8304,N_8125,N_8155);
nor U8305 (N_8305,N_8046,N_8112);
xnor U8306 (N_8306,N_8161,N_8077);
or U8307 (N_8307,N_8147,N_8020);
nand U8308 (N_8308,N_8007,N_8072);
or U8309 (N_8309,N_8010,N_8182);
nor U8310 (N_8310,N_8056,N_8032);
nand U8311 (N_8311,N_8148,N_8004);
xor U8312 (N_8312,N_8013,N_8181);
and U8313 (N_8313,N_8085,N_8185);
xnor U8314 (N_8314,N_8109,N_8199);
nand U8315 (N_8315,N_8126,N_8084);
nand U8316 (N_8316,N_8051,N_8056);
xor U8317 (N_8317,N_8163,N_8173);
xnor U8318 (N_8318,N_8114,N_8084);
and U8319 (N_8319,N_8042,N_8066);
or U8320 (N_8320,N_8157,N_8030);
and U8321 (N_8321,N_8035,N_8160);
or U8322 (N_8322,N_8088,N_8034);
nand U8323 (N_8323,N_8038,N_8042);
xnor U8324 (N_8324,N_8053,N_8154);
xor U8325 (N_8325,N_8135,N_8003);
xnor U8326 (N_8326,N_8037,N_8140);
xnor U8327 (N_8327,N_8153,N_8080);
nor U8328 (N_8328,N_8006,N_8020);
or U8329 (N_8329,N_8154,N_8057);
xor U8330 (N_8330,N_8077,N_8198);
or U8331 (N_8331,N_8069,N_8044);
or U8332 (N_8332,N_8181,N_8048);
nand U8333 (N_8333,N_8032,N_8193);
or U8334 (N_8334,N_8122,N_8148);
nor U8335 (N_8335,N_8178,N_8134);
nor U8336 (N_8336,N_8139,N_8125);
or U8337 (N_8337,N_8184,N_8096);
nor U8338 (N_8338,N_8044,N_8194);
or U8339 (N_8339,N_8045,N_8102);
and U8340 (N_8340,N_8035,N_8114);
or U8341 (N_8341,N_8008,N_8137);
and U8342 (N_8342,N_8085,N_8166);
xnor U8343 (N_8343,N_8030,N_8046);
nor U8344 (N_8344,N_8121,N_8176);
or U8345 (N_8345,N_8167,N_8062);
nand U8346 (N_8346,N_8025,N_8113);
or U8347 (N_8347,N_8125,N_8176);
or U8348 (N_8348,N_8180,N_8144);
nand U8349 (N_8349,N_8093,N_8087);
nand U8350 (N_8350,N_8048,N_8075);
or U8351 (N_8351,N_8027,N_8150);
or U8352 (N_8352,N_8113,N_8067);
or U8353 (N_8353,N_8082,N_8136);
nor U8354 (N_8354,N_8088,N_8194);
nor U8355 (N_8355,N_8071,N_8169);
nand U8356 (N_8356,N_8159,N_8006);
and U8357 (N_8357,N_8118,N_8057);
or U8358 (N_8358,N_8135,N_8173);
or U8359 (N_8359,N_8081,N_8008);
nand U8360 (N_8360,N_8117,N_8116);
nand U8361 (N_8361,N_8199,N_8108);
xnor U8362 (N_8362,N_8183,N_8096);
nand U8363 (N_8363,N_8054,N_8172);
or U8364 (N_8364,N_8119,N_8104);
or U8365 (N_8365,N_8164,N_8195);
or U8366 (N_8366,N_8069,N_8059);
nor U8367 (N_8367,N_8073,N_8178);
and U8368 (N_8368,N_8095,N_8045);
and U8369 (N_8369,N_8167,N_8134);
and U8370 (N_8370,N_8127,N_8071);
nand U8371 (N_8371,N_8056,N_8035);
and U8372 (N_8372,N_8148,N_8187);
nor U8373 (N_8373,N_8134,N_8016);
nand U8374 (N_8374,N_8086,N_8034);
xor U8375 (N_8375,N_8034,N_8011);
nor U8376 (N_8376,N_8053,N_8123);
xor U8377 (N_8377,N_8155,N_8082);
nand U8378 (N_8378,N_8151,N_8189);
nor U8379 (N_8379,N_8108,N_8084);
nor U8380 (N_8380,N_8113,N_8081);
nand U8381 (N_8381,N_8198,N_8064);
and U8382 (N_8382,N_8030,N_8133);
nor U8383 (N_8383,N_8129,N_8128);
xor U8384 (N_8384,N_8176,N_8095);
or U8385 (N_8385,N_8025,N_8068);
and U8386 (N_8386,N_8090,N_8082);
and U8387 (N_8387,N_8182,N_8083);
nand U8388 (N_8388,N_8056,N_8057);
or U8389 (N_8389,N_8043,N_8040);
nor U8390 (N_8390,N_8182,N_8159);
and U8391 (N_8391,N_8192,N_8011);
and U8392 (N_8392,N_8197,N_8096);
xnor U8393 (N_8393,N_8097,N_8011);
xnor U8394 (N_8394,N_8184,N_8019);
nor U8395 (N_8395,N_8012,N_8180);
or U8396 (N_8396,N_8171,N_8154);
nand U8397 (N_8397,N_8054,N_8019);
xnor U8398 (N_8398,N_8038,N_8141);
xnor U8399 (N_8399,N_8176,N_8186);
or U8400 (N_8400,N_8283,N_8391);
xor U8401 (N_8401,N_8294,N_8336);
and U8402 (N_8402,N_8360,N_8318);
or U8403 (N_8403,N_8220,N_8348);
nor U8404 (N_8404,N_8202,N_8344);
nor U8405 (N_8405,N_8252,N_8253);
or U8406 (N_8406,N_8244,N_8365);
xor U8407 (N_8407,N_8240,N_8298);
or U8408 (N_8408,N_8397,N_8367);
nand U8409 (N_8409,N_8339,N_8284);
nand U8410 (N_8410,N_8349,N_8297);
and U8411 (N_8411,N_8395,N_8357);
or U8412 (N_8412,N_8239,N_8387);
and U8413 (N_8413,N_8275,N_8375);
nor U8414 (N_8414,N_8225,N_8354);
or U8415 (N_8415,N_8388,N_8302);
xor U8416 (N_8416,N_8351,N_8209);
nand U8417 (N_8417,N_8271,N_8290);
xnor U8418 (N_8418,N_8361,N_8301);
nand U8419 (N_8419,N_8203,N_8260);
nor U8420 (N_8420,N_8346,N_8330);
xor U8421 (N_8421,N_8303,N_8214);
or U8422 (N_8422,N_8317,N_8287);
nor U8423 (N_8423,N_8266,N_8381);
or U8424 (N_8424,N_8245,N_8257);
nor U8425 (N_8425,N_8255,N_8394);
and U8426 (N_8426,N_8216,N_8272);
and U8427 (N_8427,N_8286,N_8385);
xor U8428 (N_8428,N_8293,N_8332);
or U8429 (N_8429,N_8396,N_8378);
xor U8430 (N_8430,N_8370,N_8208);
nor U8431 (N_8431,N_8325,N_8250);
and U8432 (N_8432,N_8377,N_8236);
or U8433 (N_8433,N_8259,N_8247);
and U8434 (N_8434,N_8308,N_8235);
nor U8435 (N_8435,N_8398,N_8364);
nand U8436 (N_8436,N_8368,N_8315);
nand U8437 (N_8437,N_8393,N_8281);
xor U8438 (N_8438,N_8341,N_8241);
or U8439 (N_8439,N_8224,N_8373);
and U8440 (N_8440,N_8264,N_8249);
nor U8441 (N_8441,N_8372,N_8307);
xor U8442 (N_8442,N_8270,N_8321);
nand U8443 (N_8443,N_8333,N_8324);
or U8444 (N_8444,N_8269,N_8399);
and U8445 (N_8445,N_8223,N_8320);
nand U8446 (N_8446,N_8386,N_8359);
nor U8447 (N_8447,N_8292,N_8384);
nand U8448 (N_8448,N_8237,N_8215);
and U8449 (N_8449,N_8379,N_8347);
or U8450 (N_8450,N_8211,N_8299);
or U8451 (N_8451,N_8256,N_8355);
xor U8452 (N_8452,N_8219,N_8280);
and U8453 (N_8453,N_8276,N_8366);
or U8454 (N_8454,N_8311,N_8242);
xor U8455 (N_8455,N_8234,N_8331);
xnor U8456 (N_8456,N_8218,N_8227);
xor U8457 (N_8457,N_8226,N_8343);
nor U8458 (N_8458,N_8291,N_8322);
and U8459 (N_8459,N_8289,N_8374);
nor U8460 (N_8460,N_8238,N_8251);
and U8461 (N_8461,N_8267,N_8210);
nor U8462 (N_8462,N_8345,N_8353);
and U8463 (N_8463,N_8313,N_8314);
nor U8464 (N_8464,N_8248,N_8312);
or U8465 (N_8465,N_8338,N_8230);
or U8466 (N_8466,N_8229,N_8340);
nand U8467 (N_8467,N_8207,N_8356);
and U8468 (N_8468,N_8296,N_8228);
or U8469 (N_8469,N_8304,N_8380);
xor U8470 (N_8470,N_8389,N_8323);
xnor U8471 (N_8471,N_8383,N_8274);
or U8472 (N_8472,N_8212,N_8316);
or U8473 (N_8473,N_8376,N_8201);
nand U8474 (N_8474,N_8200,N_8295);
nor U8475 (N_8475,N_8262,N_8288);
nor U8476 (N_8476,N_8371,N_8273);
xnor U8477 (N_8477,N_8246,N_8278);
nand U8478 (N_8478,N_8282,N_8350);
nand U8479 (N_8479,N_8369,N_8306);
and U8480 (N_8480,N_8390,N_8285);
nor U8481 (N_8481,N_8243,N_8335);
and U8482 (N_8482,N_8254,N_8337);
xor U8483 (N_8483,N_8352,N_8232);
or U8484 (N_8484,N_8217,N_8319);
nand U8485 (N_8485,N_8309,N_8326);
and U8486 (N_8486,N_8382,N_8358);
and U8487 (N_8487,N_8204,N_8342);
nand U8488 (N_8488,N_8213,N_8327);
or U8489 (N_8489,N_8300,N_8205);
nor U8490 (N_8490,N_8261,N_8277);
nor U8491 (N_8491,N_8392,N_8233);
xnor U8492 (N_8492,N_8310,N_8279);
nand U8493 (N_8493,N_8362,N_8329);
xor U8494 (N_8494,N_8231,N_8363);
nor U8495 (N_8495,N_8334,N_8222);
and U8496 (N_8496,N_8206,N_8263);
and U8497 (N_8497,N_8258,N_8305);
nand U8498 (N_8498,N_8221,N_8265);
nand U8499 (N_8499,N_8328,N_8268);
xnor U8500 (N_8500,N_8210,N_8341);
xnor U8501 (N_8501,N_8218,N_8317);
xor U8502 (N_8502,N_8374,N_8360);
nand U8503 (N_8503,N_8359,N_8247);
nor U8504 (N_8504,N_8300,N_8244);
nor U8505 (N_8505,N_8210,N_8360);
nor U8506 (N_8506,N_8357,N_8217);
or U8507 (N_8507,N_8314,N_8324);
nand U8508 (N_8508,N_8296,N_8305);
nor U8509 (N_8509,N_8371,N_8358);
nor U8510 (N_8510,N_8245,N_8309);
xnor U8511 (N_8511,N_8367,N_8259);
nand U8512 (N_8512,N_8231,N_8287);
or U8513 (N_8513,N_8236,N_8207);
nand U8514 (N_8514,N_8203,N_8393);
nor U8515 (N_8515,N_8355,N_8344);
nor U8516 (N_8516,N_8325,N_8318);
nand U8517 (N_8517,N_8334,N_8312);
and U8518 (N_8518,N_8360,N_8232);
nand U8519 (N_8519,N_8245,N_8261);
xor U8520 (N_8520,N_8239,N_8283);
xnor U8521 (N_8521,N_8274,N_8354);
nor U8522 (N_8522,N_8317,N_8323);
and U8523 (N_8523,N_8322,N_8323);
nor U8524 (N_8524,N_8387,N_8341);
xor U8525 (N_8525,N_8202,N_8327);
and U8526 (N_8526,N_8320,N_8256);
nand U8527 (N_8527,N_8325,N_8320);
nand U8528 (N_8528,N_8255,N_8317);
nand U8529 (N_8529,N_8224,N_8266);
nor U8530 (N_8530,N_8251,N_8293);
nand U8531 (N_8531,N_8315,N_8327);
or U8532 (N_8532,N_8329,N_8213);
and U8533 (N_8533,N_8212,N_8262);
nor U8534 (N_8534,N_8278,N_8320);
nand U8535 (N_8535,N_8254,N_8394);
and U8536 (N_8536,N_8234,N_8386);
nor U8537 (N_8537,N_8253,N_8390);
or U8538 (N_8538,N_8362,N_8331);
nor U8539 (N_8539,N_8330,N_8323);
and U8540 (N_8540,N_8279,N_8221);
nor U8541 (N_8541,N_8319,N_8266);
or U8542 (N_8542,N_8202,N_8383);
xor U8543 (N_8543,N_8311,N_8344);
xor U8544 (N_8544,N_8330,N_8240);
and U8545 (N_8545,N_8262,N_8360);
or U8546 (N_8546,N_8387,N_8395);
xor U8547 (N_8547,N_8296,N_8307);
and U8548 (N_8548,N_8239,N_8264);
xnor U8549 (N_8549,N_8215,N_8297);
nand U8550 (N_8550,N_8212,N_8249);
and U8551 (N_8551,N_8379,N_8387);
or U8552 (N_8552,N_8388,N_8308);
or U8553 (N_8553,N_8244,N_8249);
and U8554 (N_8554,N_8231,N_8393);
xor U8555 (N_8555,N_8322,N_8370);
and U8556 (N_8556,N_8248,N_8370);
xor U8557 (N_8557,N_8340,N_8303);
or U8558 (N_8558,N_8398,N_8360);
xnor U8559 (N_8559,N_8210,N_8276);
nand U8560 (N_8560,N_8244,N_8266);
or U8561 (N_8561,N_8370,N_8244);
xnor U8562 (N_8562,N_8340,N_8356);
and U8563 (N_8563,N_8208,N_8223);
nand U8564 (N_8564,N_8395,N_8350);
and U8565 (N_8565,N_8356,N_8380);
nor U8566 (N_8566,N_8283,N_8355);
and U8567 (N_8567,N_8274,N_8336);
nor U8568 (N_8568,N_8238,N_8264);
and U8569 (N_8569,N_8282,N_8233);
nor U8570 (N_8570,N_8251,N_8291);
and U8571 (N_8571,N_8361,N_8321);
and U8572 (N_8572,N_8321,N_8248);
nor U8573 (N_8573,N_8388,N_8342);
nor U8574 (N_8574,N_8253,N_8398);
nand U8575 (N_8575,N_8246,N_8341);
xor U8576 (N_8576,N_8305,N_8320);
or U8577 (N_8577,N_8212,N_8294);
nand U8578 (N_8578,N_8216,N_8269);
nand U8579 (N_8579,N_8275,N_8391);
nand U8580 (N_8580,N_8387,N_8265);
or U8581 (N_8581,N_8385,N_8301);
nor U8582 (N_8582,N_8306,N_8351);
nor U8583 (N_8583,N_8288,N_8253);
xor U8584 (N_8584,N_8209,N_8279);
nor U8585 (N_8585,N_8316,N_8387);
nand U8586 (N_8586,N_8370,N_8319);
nand U8587 (N_8587,N_8226,N_8316);
or U8588 (N_8588,N_8265,N_8222);
nand U8589 (N_8589,N_8382,N_8292);
and U8590 (N_8590,N_8254,N_8369);
and U8591 (N_8591,N_8229,N_8391);
nor U8592 (N_8592,N_8243,N_8311);
nor U8593 (N_8593,N_8240,N_8234);
nor U8594 (N_8594,N_8396,N_8217);
nand U8595 (N_8595,N_8223,N_8294);
and U8596 (N_8596,N_8210,N_8385);
nand U8597 (N_8597,N_8365,N_8342);
xor U8598 (N_8598,N_8304,N_8276);
nand U8599 (N_8599,N_8273,N_8325);
and U8600 (N_8600,N_8565,N_8562);
xor U8601 (N_8601,N_8426,N_8530);
xnor U8602 (N_8602,N_8524,N_8519);
nand U8603 (N_8603,N_8420,N_8534);
or U8604 (N_8604,N_8590,N_8513);
and U8605 (N_8605,N_8526,N_8425);
nand U8606 (N_8606,N_8536,N_8592);
xor U8607 (N_8607,N_8517,N_8484);
xnor U8608 (N_8608,N_8483,N_8544);
xnor U8609 (N_8609,N_8458,N_8591);
or U8610 (N_8610,N_8545,N_8515);
nor U8611 (N_8611,N_8474,N_8404);
or U8612 (N_8612,N_8480,N_8585);
nor U8613 (N_8613,N_8435,N_8464);
xnor U8614 (N_8614,N_8581,N_8569);
nand U8615 (N_8615,N_8532,N_8593);
nand U8616 (N_8616,N_8462,N_8559);
xnor U8617 (N_8617,N_8577,N_8598);
xnor U8618 (N_8618,N_8537,N_8401);
or U8619 (N_8619,N_8413,N_8495);
xor U8620 (N_8620,N_8440,N_8518);
or U8621 (N_8621,N_8410,N_8557);
or U8622 (N_8622,N_8475,N_8502);
nand U8623 (N_8623,N_8538,N_8564);
xnor U8624 (N_8624,N_8571,N_8457);
nand U8625 (N_8625,N_8533,N_8402);
or U8626 (N_8626,N_8477,N_8575);
nor U8627 (N_8627,N_8546,N_8578);
or U8628 (N_8628,N_8540,N_8451);
and U8629 (N_8629,N_8535,N_8408);
and U8630 (N_8630,N_8409,N_8560);
and U8631 (N_8631,N_8550,N_8478);
nand U8632 (N_8632,N_8563,N_8449);
or U8633 (N_8633,N_8572,N_8547);
xor U8634 (N_8634,N_8417,N_8493);
xor U8635 (N_8635,N_8423,N_8487);
or U8636 (N_8636,N_8439,N_8596);
xnor U8637 (N_8637,N_8594,N_8430);
nor U8638 (N_8638,N_8573,N_8414);
and U8639 (N_8639,N_8433,N_8541);
nand U8640 (N_8640,N_8488,N_8442);
nand U8641 (N_8641,N_8511,N_8567);
nand U8642 (N_8642,N_8586,N_8421);
nor U8643 (N_8643,N_8485,N_8482);
nand U8644 (N_8644,N_8496,N_8516);
nor U8645 (N_8645,N_8525,N_8498);
nand U8646 (N_8646,N_8422,N_8509);
nand U8647 (N_8647,N_8529,N_8510);
nand U8648 (N_8648,N_8463,N_8549);
nand U8649 (N_8649,N_8428,N_8494);
xnor U8650 (N_8650,N_8489,N_8467);
nor U8651 (N_8651,N_8522,N_8437);
or U8652 (N_8652,N_8406,N_8456);
xnor U8653 (N_8653,N_8471,N_8500);
xor U8654 (N_8654,N_8561,N_8461);
nor U8655 (N_8655,N_8470,N_8579);
nor U8656 (N_8656,N_8432,N_8528);
nand U8657 (N_8657,N_8450,N_8583);
and U8658 (N_8658,N_8403,N_8452);
nand U8659 (N_8659,N_8584,N_8445);
and U8660 (N_8660,N_8427,N_8527);
or U8661 (N_8661,N_8405,N_8446);
or U8662 (N_8662,N_8444,N_8523);
nor U8663 (N_8663,N_8595,N_8438);
or U8664 (N_8664,N_8459,N_8501);
or U8665 (N_8665,N_8580,N_8554);
and U8666 (N_8666,N_8507,N_8447);
xnor U8667 (N_8667,N_8424,N_8481);
xor U8668 (N_8668,N_8492,N_8506);
xor U8669 (N_8669,N_8531,N_8556);
nor U8670 (N_8670,N_8448,N_8505);
or U8671 (N_8671,N_8419,N_8543);
or U8672 (N_8672,N_8552,N_8434);
and U8673 (N_8673,N_8508,N_8521);
or U8674 (N_8674,N_8411,N_8412);
and U8675 (N_8675,N_8443,N_8465);
nor U8676 (N_8676,N_8454,N_8520);
and U8677 (N_8677,N_8418,N_8441);
nor U8678 (N_8678,N_8551,N_8407);
nor U8679 (N_8679,N_8460,N_8479);
xnor U8680 (N_8680,N_8476,N_8574);
nand U8681 (N_8681,N_8473,N_8555);
or U8682 (N_8682,N_8504,N_8548);
and U8683 (N_8683,N_8587,N_8415);
nor U8684 (N_8684,N_8503,N_8453);
xnor U8685 (N_8685,N_8466,N_8553);
or U8686 (N_8686,N_8582,N_8542);
or U8687 (N_8687,N_8416,N_8455);
xnor U8688 (N_8688,N_8499,N_8576);
and U8689 (N_8689,N_8469,N_8468);
and U8690 (N_8690,N_8539,N_8568);
and U8691 (N_8691,N_8588,N_8599);
nor U8692 (N_8692,N_8429,N_8512);
and U8693 (N_8693,N_8566,N_8472);
or U8694 (N_8694,N_8597,N_8558);
nor U8695 (N_8695,N_8491,N_8431);
nor U8696 (N_8696,N_8490,N_8570);
and U8697 (N_8697,N_8486,N_8589);
xnor U8698 (N_8698,N_8497,N_8436);
and U8699 (N_8699,N_8514,N_8400);
nor U8700 (N_8700,N_8402,N_8452);
xor U8701 (N_8701,N_8478,N_8599);
nor U8702 (N_8702,N_8408,N_8590);
or U8703 (N_8703,N_8574,N_8585);
or U8704 (N_8704,N_8468,N_8478);
or U8705 (N_8705,N_8556,N_8455);
nand U8706 (N_8706,N_8501,N_8497);
or U8707 (N_8707,N_8447,N_8525);
nor U8708 (N_8708,N_8448,N_8521);
nand U8709 (N_8709,N_8509,N_8419);
and U8710 (N_8710,N_8551,N_8513);
nor U8711 (N_8711,N_8462,N_8446);
xor U8712 (N_8712,N_8435,N_8520);
or U8713 (N_8713,N_8544,N_8498);
nor U8714 (N_8714,N_8481,N_8585);
and U8715 (N_8715,N_8405,N_8497);
and U8716 (N_8716,N_8407,N_8463);
and U8717 (N_8717,N_8483,N_8457);
and U8718 (N_8718,N_8446,N_8493);
or U8719 (N_8719,N_8538,N_8473);
and U8720 (N_8720,N_8530,N_8431);
nor U8721 (N_8721,N_8573,N_8546);
and U8722 (N_8722,N_8566,N_8557);
xnor U8723 (N_8723,N_8578,N_8459);
nor U8724 (N_8724,N_8457,N_8536);
and U8725 (N_8725,N_8483,N_8404);
nor U8726 (N_8726,N_8438,N_8486);
or U8727 (N_8727,N_8404,N_8413);
nand U8728 (N_8728,N_8480,N_8598);
or U8729 (N_8729,N_8413,N_8571);
xor U8730 (N_8730,N_8468,N_8484);
and U8731 (N_8731,N_8503,N_8454);
nor U8732 (N_8732,N_8421,N_8544);
xor U8733 (N_8733,N_8481,N_8522);
nor U8734 (N_8734,N_8555,N_8483);
or U8735 (N_8735,N_8405,N_8489);
nand U8736 (N_8736,N_8411,N_8450);
nand U8737 (N_8737,N_8578,N_8536);
xor U8738 (N_8738,N_8595,N_8434);
xnor U8739 (N_8739,N_8463,N_8595);
nor U8740 (N_8740,N_8505,N_8485);
nand U8741 (N_8741,N_8583,N_8420);
nor U8742 (N_8742,N_8456,N_8424);
or U8743 (N_8743,N_8474,N_8580);
nor U8744 (N_8744,N_8479,N_8438);
xnor U8745 (N_8745,N_8540,N_8489);
nor U8746 (N_8746,N_8499,N_8595);
nand U8747 (N_8747,N_8522,N_8465);
nor U8748 (N_8748,N_8565,N_8460);
nand U8749 (N_8749,N_8541,N_8427);
xnor U8750 (N_8750,N_8595,N_8559);
or U8751 (N_8751,N_8505,N_8501);
nand U8752 (N_8752,N_8546,N_8569);
nor U8753 (N_8753,N_8599,N_8576);
or U8754 (N_8754,N_8466,N_8497);
and U8755 (N_8755,N_8530,N_8526);
nand U8756 (N_8756,N_8589,N_8425);
and U8757 (N_8757,N_8460,N_8509);
and U8758 (N_8758,N_8581,N_8411);
nor U8759 (N_8759,N_8508,N_8409);
xnor U8760 (N_8760,N_8480,N_8447);
nor U8761 (N_8761,N_8502,N_8512);
xor U8762 (N_8762,N_8537,N_8430);
xnor U8763 (N_8763,N_8507,N_8437);
and U8764 (N_8764,N_8479,N_8587);
and U8765 (N_8765,N_8490,N_8576);
and U8766 (N_8766,N_8588,N_8547);
or U8767 (N_8767,N_8433,N_8501);
xnor U8768 (N_8768,N_8402,N_8445);
or U8769 (N_8769,N_8587,N_8550);
and U8770 (N_8770,N_8453,N_8522);
xnor U8771 (N_8771,N_8515,N_8438);
xnor U8772 (N_8772,N_8464,N_8409);
nand U8773 (N_8773,N_8522,N_8461);
or U8774 (N_8774,N_8534,N_8595);
xnor U8775 (N_8775,N_8534,N_8417);
nor U8776 (N_8776,N_8436,N_8468);
xor U8777 (N_8777,N_8408,N_8591);
and U8778 (N_8778,N_8425,N_8583);
or U8779 (N_8779,N_8565,N_8571);
and U8780 (N_8780,N_8483,N_8510);
or U8781 (N_8781,N_8470,N_8437);
xnor U8782 (N_8782,N_8519,N_8525);
or U8783 (N_8783,N_8545,N_8496);
xor U8784 (N_8784,N_8496,N_8595);
nand U8785 (N_8785,N_8566,N_8465);
nand U8786 (N_8786,N_8598,N_8481);
nor U8787 (N_8787,N_8513,N_8489);
nand U8788 (N_8788,N_8532,N_8404);
or U8789 (N_8789,N_8569,N_8543);
nand U8790 (N_8790,N_8420,N_8568);
nand U8791 (N_8791,N_8582,N_8478);
or U8792 (N_8792,N_8413,N_8465);
nor U8793 (N_8793,N_8461,N_8504);
or U8794 (N_8794,N_8469,N_8418);
or U8795 (N_8795,N_8558,N_8468);
nor U8796 (N_8796,N_8588,N_8573);
and U8797 (N_8797,N_8504,N_8410);
xor U8798 (N_8798,N_8598,N_8548);
and U8799 (N_8799,N_8456,N_8439);
xor U8800 (N_8800,N_8757,N_8660);
or U8801 (N_8801,N_8651,N_8730);
nor U8802 (N_8802,N_8618,N_8695);
nor U8803 (N_8803,N_8728,N_8710);
xnor U8804 (N_8804,N_8763,N_8793);
and U8805 (N_8805,N_8671,N_8631);
nor U8806 (N_8806,N_8739,N_8636);
xor U8807 (N_8807,N_8766,N_8609);
nor U8808 (N_8808,N_8760,N_8605);
nand U8809 (N_8809,N_8770,N_8784);
or U8810 (N_8810,N_8691,N_8679);
and U8811 (N_8811,N_8738,N_8753);
nand U8812 (N_8812,N_8792,N_8602);
xnor U8813 (N_8813,N_8683,N_8657);
xor U8814 (N_8814,N_8771,N_8720);
nor U8815 (N_8815,N_8702,N_8717);
nand U8816 (N_8816,N_8659,N_8632);
xor U8817 (N_8817,N_8669,N_8685);
nand U8818 (N_8818,N_8666,N_8707);
or U8819 (N_8819,N_8667,N_8721);
and U8820 (N_8820,N_8773,N_8662);
xor U8821 (N_8821,N_8733,N_8604);
xnor U8822 (N_8822,N_8655,N_8790);
xor U8823 (N_8823,N_8718,N_8644);
nor U8824 (N_8824,N_8670,N_8622);
nand U8825 (N_8825,N_8626,N_8700);
and U8826 (N_8826,N_8789,N_8656);
nor U8827 (N_8827,N_8729,N_8603);
or U8828 (N_8828,N_8608,N_8616);
xnor U8829 (N_8829,N_8752,N_8712);
nand U8830 (N_8830,N_8780,N_8779);
and U8831 (N_8831,N_8617,N_8647);
or U8832 (N_8832,N_8676,N_8740);
nor U8833 (N_8833,N_8797,N_8787);
nor U8834 (N_8834,N_8765,N_8736);
nor U8835 (N_8835,N_8758,N_8648);
nor U8836 (N_8836,N_8678,N_8762);
and U8837 (N_8837,N_8689,N_8737);
and U8838 (N_8838,N_8697,N_8751);
or U8839 (N_8839,N_8782,N_8675);
xnor U8840 (N_8840,N_8630,N_8688);
xor U8841 (N_8841,N_8791,N_8615);
and U8842 (N_8842,N_8600,N_8637);
or U8843 (N_8843,N_8634,N_8607);
nor U8844 (N_8844,N_8638,N_8681);
or U8845 (N_8845,N_8749,N_8725);
and U8846 (N_8846,N_8682,N_8744);
and U8847 (N_8847,N_8723,N_8799);
or U8848 (N_8848,N_8743,N_8783);
and U8849 (N_8849,N_8654,N_8620);
or U8850 (N_8850,N_8614,N_8680);
nor U8851 (N_8851,N_8703,N_8708);
nand U8852 (N_8852,N_8696,N_8724);
or U8853 (N_8853,N_8714,N_8750);
or U8854 (N_8854,N_8642,N_8687);
nor U8855 (N_8855,N_8694,N_8668);
and U8856 (N_8856,N_8719,N_8623);
or U8857 (N_8857,N_8774,N_8767);
nor U8858 (N_8858,N_8650,N_8633);
nand U8859 (N_8859,N_8619,N_8745);
and U8860 (N_8860,N_8741,N_8768);
or U8861 (N_8861,N_8798,N_8726);
xnor U8862 (N_8862,N_8735,N_8628);
or U8863 (N_8863,N_8713,N_8775);
or U8864 (N_8864,N_8621,N_8716);
and U8865 (N_8865,N_8673,N_8652);
xor U8866 (N_8866,N_8706,N_8665);
xor U8867 (N_8867,N_8627,N_8701);
and U8868 (N_8868,N_8734,N_8722);
xor U8869 (N_8869,N_8759,N_8663);
or U8870 (N_8870,N_8778,N_8794);
and U8871 (N_8871,N_8612,N_8640);
xor U8872 (N_8872,N_8742,N_8788);
nor U8873 (N_8873,N_8769,N_8732);
or U8874 (N_8874,N_8606,N_8764);
and U8875 (N_8875,N_8777,N_8613);
nand U8876 (N_8876,N_8645,N_8727);
or U8877 (N_8877,N_8776,N_8693);
xor U8878 (N_8878,N_8698,N_8692);
nor U8879 (N_8879,N_8674,N_8658);
xor U8880 (N_8880,N_8709,N_8625);
nand U8881 (N_8881,N_8684,N_8699);
nor U8882 (N_8882,N_8796,N_8690);
and U8883 (N_8883,N_8661,N_8672);
or U8884 (N_8884,N_8747,N_8649);
and U8885 (N_8885,N_8629,N_8610);
nand U8886 (N_8886,N_8686,N_8731);
nor U8887 (N_8887,N_8711,N_8705);
and U8888 (N_8888,N_8748,N_8755);
nor U8889 (N_8889,N_8639,N_8677);
and U8890 (N_8890,N_8795,N_8624);
or U8891 (N_8891,N_8646,N_8746);
nand U8892 (N_8892,N_8715,N_8786);
and U8893 (N_8893,N_8653,N_8761);
xor U8894 (N_8894,N_8785,N_8611);
or U8895 (N_8895,N_8641,N_8643);
nand U8896 (N_8896,N_8635,N_8754);
or U8897 (N_8897,N_8601,N_8756);
or U8898 (N_8898,N_8704,N_8781);
nand U8899 (N_8899,N_8772,N_8664);
nand U8900 (N_8900,N_8709,N_8613);
or U8901 (N_8901,N_8649,N_8792);
nor U8902 (N_8902,N_8672,N_8689);
and U8903 (N_8903,N_8757,N_8782);
and U8904 (N_8904,N_8752,N_8669);
nand U8905 (N_8905,N_8764,N_8761);
and U8906 (N_8906,N_8682,N_8629);
and U8907 (N_8907,N_8682,N_8699);
xor U8908 (N_8908,N_8668,N_8764);
nor U8909 (N_8909,N_8601,N_8620);
nand U8910 (N_8910,N_8620,N_8628);
and U8911 (N_8911,N_8600,N_8733);
nand U8912 (N_8912,N_8655,N_8623);
xor U8913 (N_8913,N_8768,N_8646);
xor U8914 (N_8914,N_8763,N_8791);
nor U8915 (N_8915,N_8625,N_8786);
or U8916 (N_8916,N_8726,N_8619);
nand U8917 (N_8917,N_8639,N_8745);
xor U8918 (N_8918,N_8651,N_8704);
xor U8919 (N_8919,N_8769,N_8624);
and U8920 (N_8920,N_8719,N_8754);
and U8921 (N_8921,N_8617,N_8798);
nand U8922 (N_8922,N_8740,N_8600);
or U8923 (N_8923,N_8794,N_8671);
and U8924 (N_8924,N_8781,N_8755);
and U8925 (N_8925,N_8652,N_8629);
nand U8926 (N_8926,N_8784,N_8733);
and U8927 (N_8927,N_8693,N_8716);
and U8928 (N_8928,N_8657,N_8634);
xor U8929 (N_8929,N_8680,N_8795);
nor U8930 (N_8930,N_8657,N_8776);
and U8931 (N_8931,N_8757,N_8719);
nor U8932 (N_8932,N_8647,N_8646);
xnor U8933 (N_8933,N_8787,N_8733);
xor U8934 (N_8934,N_8665,N_8712);
nor U8935 (N_8935,N_8686,N_8609);
or U8936 (N_8936,N_8722,N_8612);
nor U8937 (N_8937,N_8672,N_8680);
nand U8938 (N_8938,N_8605,N_8737);
and U8939 (N_8939,N_8688,N_8644);
or U8940 (N_8940,N_8728,N_8646);
nor U8941 (N_8941,N_8617,N_8779);
xnor U8942 (N_8942,N_8630,N_8752);
or U8943 (N_8943,N_8607,N_8754);
nor U8944 (N_8944,N_8672,N_8615);
nand U8945 (N_8945,N_8696,N_8616);
or U8946 (N_8946,N_8634,N_8674);
or U8947 (N_8947,N_8730,N_8700);
and U8948 (N_8948,N_8706,N_8629);
nor U8949 (N_8949,N_8757,N_8762);
nor U8950 (N_8950,N_8638,N_8720);
and U8951 (N_8951,N_8785,N_8767);
nand U8952 (N_8952,N_8615,N_8610);
nand U8953 (N_8953,N_8627,N_8665);
and U8954 (N_8954,N_8698,N_8686);
nand U8955 (N_8955,N_8689,N_8721);
nor U8956 (N_8956,N_8613,N_8736);
and U8957 (N_8957,N_8766,N_8789);
nor U8958 (N_8958,N_8786,N_8791);
nor U8959 (N_8959,N_8635,N_8663);
xnor U8960 (N_8960,N_8730,N_8721);
nand U8961 (N_8961,N_8602,N_8722);
xnor U8962 (N_8962,N_8663,N_8614);
xor U8963 (N_8963,N_8744,N_8728);
xnor U8964 (N_8964,N_8796,N_8667);
or U8965 (N_8965,N_8702,N_8670);
nand U8966 (N_8966,N_8708,N_8615);
and U8967 (N_8967,N_8724,N_8777);
and U8968 (N_8968,N_8699,N_8733);
nor U8969 (N_8969,N_8781,N_8716);
or U8970 (N_8970,N_8626,N_8676);
or U8971 (N_8971,N_8726,N_8794);
or U8972 (N_8972,N_8666,N_8725);
nand U8973 (N_8973,N_8761,N_8630);
and U8974 (N_8974,N_8766,N_8622);
nand U8975 (N_8975,N_8675,N_8634);
or U8976 (N_8976,N_8612,N_8719);
and U8977 (N_8977,N_8669,N_8639);
nand U8978 (N_8978,N_8758,N_8605);
nand U8979 (N_8979,N_8712,N_8677);
xor U8980 (N_8980,N_8748,N_8739);
nor U8981 (N_8981,N_8701,N_8674);
xor U8982 (N_8982,N_8602,N_8747);
nand U8983 (N_8983,N_8627,N_8636);
xnor U8984 (N_8984,N_8762,N_8708);
or U8985 (N_8985,N_8700,N_8758);
nand U8986 (N_8986,N_8646,N_8716);
xnor U8987 (N_8987,N_8723,N_8606);
and U8988 (N_8988,N_8764,N_8662);
nor U8989 (N_8989,N_8641,N_8792);
and U8990 (N_8990,N_8724,N_8705);
and U8991 (N_8991,N_8726,N_8623);
nand U8992 (N_8992,N_8735,N_8632);
xnor U8993 (N_8993,N_8714,N_8760);
nor U8994 (N_8994,N_8617,N_8744);
nand U8995 (N_8995,N_8634,N_8755);
xor U8996 (N_8996,N_8646,N_8616);
and U8997 (N_8997,N_8690,N_8789);
xor U8998 (N_8998,N_8689,N_8692);
or U8999 (N_8999,N_8695,N_8640);
or U9000 (N_9000,N_8898,N_8892);
nor U9001 (N_9001,N_8843,N_8986);
and U9002 (N_9002,N_8854,N_8861);
and U9003 (N_9003,N_8912,N_8981);
or U9004 (N_9004,N_8872,N_8888);
and U9005 (N_9005,N_8869,N_8859);
and U9006 (N_9006,N_8936,N_8988);
nor U9007 (N_9007,N_8978,N_8865);
or U9008 (N_9008,N_8969,N_8958);
nor U9009 (N_9009,N_8954,N_8808);
or U9010 (N_9010,N_8935,N_8873);
nand U9011 (N_9011,N_8910,N_8991);
or U9012 (N_9012,N_8966,N_8868);
xnor U9013 (N_9013,N_8922,N_8864);
or U9014 (N_9014,N_8887,N_8820);
or U9015 (N_9015,N_8812,N_8879);
nor U9016 (N_9016,N_8827,N_8909);
or U9017 (N_9017,N_8943,N_8976);
nand U9018 (N_9018,N_8870,N_8832);
and U9019 (N_9019,N_8916,N_8955);
xor U9020 (N_9020,N_8924,N_8894);
xnor U9021 (N_9021,N_8996,N_8886);
or U9022 (N_9022,N_8972,N_8825);
or U9023 (N_9023,N_8877,N_8884);
nor U9024 (N_9024,N_8850,N_8855);
nand U9025 (N_9025,N_8907,N_8973);
and U9026 (N_9026,N_8993,N_8921);
or U9027 (N_9027,N_8878,N_8807);
or U9028 (N_9028,N_8919,N_8891);
or U9029 (N_9029,N_8800,N_8893);
and U9030 (N_9030,N_8944,N_8862);
and U9031 (N_9031,N_8956,N_8951);
nor U9032 (N_9032,N_8881,N_8974);
nand U9033 (N_9033,N_8945,N_8942);
xor U9034 (N_9034,N_8918,N_8901);
or U9035 (N_9035,N_8815,N_8964);
nor U9036 (N_9036,N_8933,N_8947);
xnor U9037 (N_9037,N_8831,N_8897);
nand U9038 (N_9038,N_8851,N_8937);
nand U9039 (N_9039,N_8880,N_8914);
nand U9040 (N_9040,N_8906,N_8997);
xnor U9041 (N_9041,N_8813,N_8876);
and U9042 (N_9042,N_8806,N_8983);
nand U9043 (N_9043,N_8835,N_8801);
nand U9044 (N_9044,N_8828,N_8804);
nand U9045 (N_9045,N_8809,N_8938);
nand U9046 (N_9046,N_8890,N_8840);
or U9047 (N_9047,N_8814,N_8928);
or U9048 (N_9048,N_8932,N_8911);
and U9049 (N_9049,N_8853,N_8823);
or U9050 (N_9050,N_8989,N_8905);
xor U9051 (N_9051,N_8948,N_8883);
nand U9052 (N_9052,N_8805,N_8963);
and U9053 (N_9053,N_8839,N_8882);
and U9054 (N_9054,N_8957,N_8803);
or U9055 (N_9055,N_8939,N_8908);
or U9056 (N_9056,N_8959,N_8841);
xnor U9057 (N_9057,N_8925,N_8930);
nor U9058 (N_9058,N_8857,N_8979);
nor U9059 (N_9059,N_8816,N_8889);
xnor U9060 (N_9060,N_8999,N_8817);
xor U9061 (N_9061,N_8995,N_8849);
or U9062 (N_9062,N_8977,N_8950);
and U9063 (N_9063,N_8940,N_8949);
and U9064 (N_9064,N_8846,N_8915);
nand U9065 (N_9065,N_8975,N_8852);
and U9066 (N_9066,N_8941,N_8867);
and U9067 (N_9067,N_8837,N_8818);
or U9068 (N_9068,N_8962,N_8871);
and U9069 (N_9069,N_8833,N_8965);
or U9070 (N_9070,N_8967,N_8926);
nand U9071 (N_9071,N_8844,N_8931);
nand U9072 (N_9072,N_8848,N_8987);
xor U9073 (N_9073,N_8992,N_8953);
and U9074 (N_9074,N_8834,N_8970);
xnor U9075 (N_9075,N_8971,N_8904);
or U9076 (N_9076,N_8811,N_8845);
or U9077 (N_9077,N_8990,N_8824);
nand U9078 (N_9078,N_8860,N_8899);
nor U9079 (N_9079,N_8920,N_8842);
xnor U9080 (N_9080,N_8980,N_8896);
xor U9081 (N_9081,N_8994,N_8985);
xor U9082 (N_9082,N_8895,N_8952);
or U9083 (N_9083,N_8902,N_8838);
and U9084 (N_9084,N_8830,N_8802);
and U9085 (N_9085,N_8829,N_8961);
xor U9086 (N_9086,N_8847,N_8913);
or U9087 (N_9087,N_8984,N_8875);
nor U9088 (N_9088,N_8968,N_8810);
nand U9089 (N_9089,N_8822,N_8903);
nor U9090 (N_9090,N_8998,N_8982);
or U9091 (N_9091,N_8934,N_8923);
and U9092 (N_9092,N_8863,N_8917);
xnor U9093 (N_9093,N_8836,N_8826);
nand U9094 (N_9094,N_8900,N_8821);
nor U9095 (N_9095,N_8960,N_8856);
or U9096 (N_9096,N_8927,N_8885);
nand U9097 (N_9097,N_8866,N_8929);
nand U9098 (N_9098,N_8946,N_8819);
or U9099 (N_9099,N_8858,N_8874);
xor U9100 (N_9100,N_8885,N_8806);
and U9101 (N_9101,N_8966,N_8851);
xor U9102 (N_9102,N_8983,N_8889);
and U9103 (N_9103,N_8921,N_8994);
xor U9104 (N_9104,N_8830,N_8833);
xnor U9105 (N_9105,N_8941,N_8804);
nand U9106 (N_9106,N_8906,N_8811);
nand U9107 (N_9107,N_8971,N_8909);
or U9108 (N_9108,N_8813,N_8892);
nand U9109 (N_9109,N_8911,N_8869);
or U9110 (N_9110,N_8855,N_8880);
xnor U9111 (N_9111,N_8946,N_8963);
xnor U9112 (N_9112,N_8861,N_8845);
nor U9113 (N_9113,N_8822,N_8930);
and U9114 (N_9114,N_8836,N_8810);
xnor U9115 (N_9115,N_8818,N_8971);
nand U9116 (N_9116,N_8877,N_8891);
or U9117 (N_9117,N_8940,N_8817);
or U9118 (N_9118,N_8800,N_8910);
nor U9119 (N_9119,N_8816,N_8992);
and U9120 (N_9120,N_8929,N_8920);
and U9121 (N_9121,N_8945,N_8896);
nand U9122 (N_9122,N_8878,N_8914);
or U9123 (N_9123,N_8812,N_8970);
nor U9124 (N_9124,N_8914,N_8823);
and U9125 (N_9125,N_8867,N_8830);
or U9126 (N_9126,N_8845,N_8937);
xnor U9127 (N_9127,N_8886,N_8990);
and U9128 (N_9128,N_8853,N_8827);
nor U9129 (N_9129,N_8857,N_8830);
nor U9130 (N_9130,N_8824,N_8847);
xor U9131 (N_9131,N_8879,N_8857);
and U9132 (N_9132,N_8800,N_8834);
nand U9133 (N_9133,N_8949,N_8982);
and U9134 (N_9134,N_8805,N_8887);
nor U9135 (N_9135,N_8995,N_8865);
xnor U9136 (N_9136,N_8946,N_8845);
and U9137 (N_9137,N_8973,N_8998);
nor U9138 (N_9138,N_8909,N_8899);
or U9139 (N_9139,N_8921,N_8801);
xor U9140 (N_9140,N_8989,N_8859);
and U9141 (N_9141,N_8919,N_8845);
nor U9142 (N_9142,N_8851,N_8847);
nand U9143 (N_9143,N_8885,N_8883);
nor U9144 (N_9144,N_8800,N_8802);
and U9145 (N_9145,N_8818,N_8862);
and U9146 (N_9146,N_8818,N_8858);
and U9147 (N_9147,N_8872,N_8802);
xnor U9148 (N_9148,N_8955,N_8890);
nand U9149 (N_9149,N_8808,N_8977);
or U9150 (N_9150,N_8803,N_8909);
nand U9151 (N_9151,N_8857,N_8898);
nand U9152 (N_9152,N_8859,N_8825);
xnor U9153 (N_9153,N_8852,N_8823);
or U9154 (N_9154,N_8831,N_8972);
nor U9155 (N_9155,N_8892,N_8877);
nand U9156 (N_9156,N_8860,N_8862);
nor U9157 (N_9157,N_8996,N_8889);
nor U9158 (N_9158,N_8973,N_8908);
and U9159 (N_9159,N_8835,N_8938);
nor U9160 (N_9160,N_8864,N_8990);
and U9161 (N_9161,N_8835,N_8941);
xor U9162 (N_9162,N_8857,N_8934);
nand U9163 (N_9163,N_8851,N_8982);
xnor U9164 (N_9164,N_8960,N_8865);
nand U9165 (N_9165,N_8990,N_8939);
nor U9166 (N_9166,N_8865,N_8956);
or U9167 (N_9167,N_8800,N_8830);
and U9168 (N_9168,N_8806,N_8834);
nor U9169 (N_9169,N_8896,N_8857);
xnor U9170 (N_9170,N_8986,N_8901);
or U9171 (N_9171,N_8920,N_8904);
or U9172 (N_9172,N_8938,N_8948);
or U9173 (N_9173,N_8988,N_8825);
nand U9174 (N_9174,N_8937,N_8972);
nor U9175 (N_9175,N_8839,N_8803);
nand U9176 (N_9176,N_8801,N_8934);
xor U9177 (N_9177,N_8919,N_8992);
or U9178 (N_9178,N_8821,N_8956);
nor U9179 (N_9179,N_8833,N_8853);
nor U9180 (N_9180,N_8821,N_8823);
xor U9181 (N_9181,N_8808,N_8998);
nand U9182 (N_9182,N_8983,N_8816);
or U9183 (N_9183,N_8824,N_8854);
nor U9184 (N_9184,N_8944,N_8957);
nand U9185 (N_9185,N_8899,N_8813);
nor U9186 (N_9186,N_8963,N_8856);
and U9187 (N_9187,N_8933,N_8856);
or U9188 (N_9188,N_8950,N_8899);
nand U9189 (N_9189,N_8947,N_8938);
nor U9190 (N_9190,N_8983,N_8873);
and U9191 (N_9191,N_8877,N_8829);
xnor U9192 (N_9192,N_8915,N_8989);
nor U9193 (N_9193,N_8869,N_8947);
xor U9194 (N_9194,N_8962,N_8998);
nand U9195 (N_9195,N_8971,N_8959);
and U9196 (N_9196,N_8854,N_8922);
nor U9197 (N_9197,N_8918,N_8907);
and U9198 (N_9198,N_8951,N_8972);
nor U9199 (N_9199,N_8944,N_8962);
xor U9200 (N_9200,N_9192,N_9036);
nor U9201 (N_9201,N_9015,N_9139);
and U9202 (N_9202,N_9122,N_9153);
nand U9203 (N_9203,N_9029,N_9049);
nand U9204 (N_9204,N_9003,N_9148);
and U9205 (N_9205,N_9088,N_9109);
and U9206 (N_9206,N_9188,N_9190);
nor U9207 (N_9207,N_9103,N_9063);
or U9208 (N_9208,N_9017,N_9030);
xor U9209 (N_9209,N_9054,N_9039);
or U9210 (N_9210,N_9105,N_9066);
or U9211 (N_9211,N_9115,N_9126);
or U9212 (N_9212,N_9038,N_9171);
or U9213 (N_9213,N_9018,N_9113);
or U9214 (N_9214,N_9092,N_9133);
nor U9215 (N_9215,N_9140,N_9072);
nor U9216 (N_9216,N_9043,N_9175);
and U9217 (N_9217,N_9014,N_9123);
or U9218 (N_9218,N_9021,N_9080);
xnor U9219 (N_9219,N_9197,N_9187);
or U9220 (N_9220,N_9004,N_9112);
nand U9221 (N_9221,N_9095,N_9068);
xor U9222 (N_9222,N_9114,N_9193);
nor U9223 (N_9223,N_9041,N_9138);
and U9224 (N_9224,N_9044,N_9056);
xnor U9225 (N_9225,N_9013,N_9087);
nor U9226 (N_9226,N_9045,N_9019);
and U9227 (N_9227,N_9048,N_9195);
and U9228 (N_9228,N_9006,N_9034);
nand U9229 (N_9229,N_9132,N_9178);
nor U9230 (N_9230,N_9141,N_9129);
nand U9231 (N_9231,N_9011,N_9137);
nand U9232 (N_9232,N_9067,N_9009);
or U9233 (N_9233,N_9104,N_9128);
and U9234 (N_9234,N_9145,N_9010);
or U9235 (N_9235,N_9191,N_9162);
nor U9236 (N_9236,N_9119,N_9108);
xor U9237 (N_9237,N_9199,N_9196);
and U9238 (N_9238,N_9179,N_9173);
xor U9239 (N_9239,N_9079,N_9055);
xnor U9240 (N_9240,N_9099,N_9110);
or U9241 (N_9241,N_9177,N_9157);
or U9242 (N_9242,N_9125,N_9118);
and U9243 (N_9243,N_9016,N_9028);
or U9244 (N_9244,N_9012,N_9127);
nor U9245 (N_9245,N_9078,N_9089);
xnor U9246 (N_9246,N_9024,N_9098);
xor U9247 (N_9247,N_9147,N_9025);
and U9248 (N_9248,N_9052,N_9007);
and U9249 (N_9249,N_9154,N_9184);
xor U9250 (N_9250,N_9176,N_9073);
nand U9251 (N_9251,N_9047,N_9168);
nor U9252 (N_9252,N_9163,N_9060);
or U9253 (N_9253,N_9155,N_9093);
nor U9254 (N_9254,N_9158,N_9000);
nor U9255 (N_9255,N_9146,N_9090);
nand U9256 (N_9256,N_9094,N_9117);
nand U9257 (N_9257,N_9035,N_9111);
nand U9258 (N_9258,N_9031,N_9160);
and U9259 (N_9259,N_9074,N_9005);
nor U9260 (N_9260,N_9001,N_9165);
nor U9261 (N_9261,N_9070,N_9050);
nor U9262 (N_9262,N_9164,N_9037);
or U9263 (N_9263,N_9076,N_9120);
xor U9264 (N_9264,N_9069,N_9149);
nand U9265 (N_9265,N_9102,N_9057);
xor U9266 (N_9266,N_9027,N_9002);
or U9267 (N_9267,N_9042,N_9169);
and U9268 (N_9268,N_9033,N_9058);
nand U9269 (N_9269,N_9046,N_9062);
and U9270 (N_9270,N_9084,N_9064);
and U9271 (N_9271,N_9151,N_9135);
nand U9272 (N_9272,N_9100,N_9083);
xnor U9273 (N_9273,N_9065,N_9101);
nand U9274 (N_9274,N_9194,N_9061);
and U9275 (N_9275,N_9124,N_9131);
xor U9276 (N_9276,N_9059,N_9023);
or U9277 (N_9277,N_9040,N_9121);
nand U9278 (N_9278,N_9020,N_9134);
or U9279 (N_9279,N_9075,N_9142);
or U9280 (N_9280,N_9174,N_9032);
nand U9281 (N_9281,N_9051,N_9150);
nor U9282 (N_9282,N_9186,N_9143);
and U9283 (N_9283,N_9152,N_9096);
xor U9284 (N_9284,N_9077,N_9185);
nor U9285 (N_9285,N_9159,N_9091);
or U9286 (N_9286,N_9116,N_9161);
nand U9287 (N_9287,N_9167,N_9097);
or U9288 (N_9288,N_9086,N_9085);
and U9289 (N_9289,N_9181,N_9081);
nand U9290 (N_9290,N_9022,N_9198);
or U9291 (N_9291,N_9107,N_9189);
nand U9292 (N_9292,N_9183,N_9170);
nand U9293 (N_9293,N_9053,N_9082);
xnor U9294 (N_9294,N_9130,N_9172);
or U9295 (N_9295,N_9106,N_9156);
nand U9296 (N_9296,N_9136,N_9026);
xnor U9297 (N_9297,N_9180,N_9182);
nand U9298 (N_9298,N_9008,N_9166);
and U9299 (N_9299,N_9071,N_9144);
xnor U9300 (N_9300,N_9054,N_9001);
xnor U9301 (N_9301,N_9195,N_9140);
xnor U9302 (N_9302,N_9069,N_9077);
nand U9303 (N_9303,N_9182,N_9026);
or U9304 (N_9304,N_9036,N_9127);
xnor U9305 (N_9305,N_9036,N_9113);
or U9306 (N_9306,N_9055,N_9177);
or U9307 (N_9307,N_9183,N_9149);
nor U9308 (N_9308,N_9170,N_9199);
xor U9309 (N_9309,N_9163,N_9051);
nor U9310 (N_9310,N_9113,N_9112);
xnor U9311 (N_9311,N_9132,N_9160);
and U9312 (N_9312,N_9127,N_9076);
xor U9313 (N_9313,N_9071,N_9122);
nor U9314 (N_9314,N_9190,N_9101);
or U9315 (N_9315,N_9176,N_9187);
xnor U9316 (N_9316,N_9065,N_9193);
nor U9317 (N_9317,N_9172,N_9192);
nor U9318 (N_9318,N_9075,N_9058);
and U9319 (N_9319,N_9182,N_9039);
nor U9320 (N_9320,N_9016,N_9124);
nand U9321 (N_9321,N_9034,N_9111);
xnor U9322 (N_9322,N_9061,N_9153);
and U9323 (N_9323,N_9148,N_9121);
and U9324 (N_9324,N_9082,N_9103);
or U9325 (N_9325,N_9194,N_9134);
or U9326 (N_9326,N_9106,N_9088);
and U9327 (N_9327,N_9101,N_9163);
or U9328 (N_9328,N_9019,N_9158);
and U9329 (N_9329,N_9091,N_9152);
and U9330 (N_9330,N_9053,N_9042);
nand U9331 (N_9331,N_9156,N_9048);
nand U9332 (N_9332,N_9090,N_9114);
nor U9333 (N_9333,N_9197,N_9160);
and U9334 (N_9334,N_9137,N_9058);
or U9335 (N_9335,N_9158,N_9029);
or U9336 (N_9336,N_9189,N_9038);
nand U9337 (N_9337,N_9189,N_9146);
xor U9338 (N_9338,N_9129,N_9082);
and U9339 (N_9339,N_9034,N_9066);
nor U9340 (N_9340,N_9023,N_9097);
or U9341 (N_9341,N_9075,N_9046);
and U9342 (N_9342,N_9026,N_9096);
nand U9343 (N_9343,N_9193,N_9121);
nand U9344 (N_9344,N_9033,N_9086);
nor U9345 (N_9345,N_9140,N_9054);
xor U9346 (N_9346,N_9113,N_9060);
and U9347 (N_9347,N_9147,N_9173);
or U9348 (N_9348,N_9165,N_9023);
and U9349 (N_9349,N_9033,N_9002);
xnor U9350 (N_9350,N_9180,N_9131);
or U9351 (N_9351,N_9174,N_9066);
or U9352 (N_9352,N_9147,N_9040);
or U9353 (N_9353,N_9147,N_9132);
nor U9354 (N_9354,N_9020,N_9101);
and U9355 (N_9355,N_9043,N_9069);
or U9356 (N_9356,N_9077,N_9071);
nand U9357 (N_9357,N_9176,N_9042);
and U9358 (N_9358,N_9019,N_9128);
or U9359 (N_9359,N_9028,N_9145);
or U9360 (N_9360,N_9013,N_9006);
and U9361 (N_9361,N_9108,N_9127);
nor U9362 (N_9362,N_9000,N_9194);
xnor U9363 (N_9363,N_9053,N_9116);
and U9364 (N_9364,N_9153,N_9020);
xnor U9365 (N_9365,N_9021,N_9173);
and U9366 (N_9366,N_9070,N_9008);
xor U9367 (N_9367,N_9000,N_9045);
or U9368 (N_9368,N_9086,N_9186);
xor U9369 (N_9369,N_9020,N_9177);
or U9370 (N_9370,N_9144,N_9069);
xnor U9371 (N_9371,N_9061,N_9056);
xnor U9372 (N_9372,N_9101,N_9096);
xnor U9373 (N_9373,N_9051,N_9077);
or U9374 (N_9374,N_9170,N_9061);
or U9375 (N_9375,N_9027,N_9010);
nor U9376 (N_9376,N_9024,N_9034);
or U9377 (N_9377,N_9025,N_9031);
and U9378 (N_9378,N_9185,N_9052);
nor U9379 (N_9379,N_9114,N_9086);
or U9380 (N_9380,N_9174,N_9026);
xor U9381 (N_9381,N_9025,N_9132);
and U9382 (N_9382,N_9061,N_9122);
nor U9383 (N_9383,N_9190,N_9110);
or U9384 (N_9384,N_9035,N_9157);
xor U9385 (N_9385,N_9098,N_9064);
and U9386 (N_9386,N_9028,N_9012);
nor U9387 (N_9387,N_9124,N_9133);
nor U9388 (N_9388,N_9084,N_9016);
nand U9389 (N_9389,N_9161,N_9125);
xnor U9390 (N_9390,N_9029,N_9000);
and U9391 (N_9391,N_9137,N_9014);
xor U9392 (N_9392,N_9025,N_9087);
and U9393 (N_9393,N_9000,N_9155);
and U9394 (N_9394,N_9103,N_9182);
nor U9395 (N_9395,N_9197,N_9077);
nand U9396 (N_9396,N_9079,N_9039);
xor U9397 (N_9397,N_9112,N_9138);
xor U9398 (N_9398,N_9101,N_9004);
nand U9399 (N_9399,N_9007,N_9140);
xor U9400 (N_9400,N_9291,N_9315);
or U9401 (N_9401,N_9320,N_9245);
and U9402 (N_9402,N_9243,N_9346);
nor U9403 (N_9403,N_9336,N_9331);
or U9404 (N_9404,N_9378,N_9298);
and U9405 (N_9405,N_9307,N_9257);
xnor U9406 (N_9406,N_9224,N_9314);
nand U9407 (N_9407,N_9312,N_9348);
or U9408 (N_9408,N_9205,N_9204);
nand U9409 (N_9409,N_9286,N_9393);
nor U9410 (N_9410,N_9284,N_9367);
nor U9411 (N_9411,N_9354,N_9337);
xor U9412 (N_9412,N_9203,N_9231);
and U9413 (N_9413,N_9392,N_9221);
or U9414 (N_9414,N_9325,N_9214);
or U9415 (N_9415,N_9271,N_9283);
nor U9416 (N_9416,N_9328,N_9310);
or U9417 (N_9417,N_9368,N_9247);
nor U9418 (N_9418,N_9351,N_9326);
and U9419 (N_9419,N_9287,N_9381);
and U9420 (N_9420,N_9294,N_9342);
nand U9421 (N_9421,N_9263,N_9226);
xnor U9422 (N_9422,N_9251,N_9281);
xnor U9423 (N_9423,N_9345,N_9202);
or U9424 (N_9424,N_9222,N_9282);
xor U9425 (N_9425,N_9277,N_9249);
or U9426 (N_9426,N_9279,N_9292);
or U9427 (N_9427,N_9219,N_9208);
nor U9428 (N_9428,N_9356,N_9352);
nor U9429 (N_9429,N_9382,N_9275);
or U9430 (N_9430,N_9323,N_9327);
nand U9431 (N_9431,N_9297,N_9280);
and U9432 (N_9432,N_9340,N_9268);
or U9433 (N_9433,N_9376,N_9335);
nand U9434 (N_9434,N_9359,N_9293);
or U9435 (N_9435,N_9217,N_9240);
nor U9436 (N_9436,N_9261,N_9313);
nor U9437 (N_9437,N_9252,N_9383);
nor U9438 (N_9438,N_9216,N_9225);
nand U9439 (N_9439,N_9397,N_9250);
xor U9440 (N_9440,N_9303,N_9248);
and U9441 (N_9441,N_9301,N_9375);
nand U9442 (N_9442,N_9230,N_9329);
or U9443 (N_9443,N_9264,N_9322);
xnor U9444 (N_9444,N_9209,N_9344);
or U9445 (N_9445,N_9387,N_9339);
nor U9446 (N_9446,N_9333,N_9255);
xor U9447 (N_9447,N_9259,N_9318);
nand U9448 (N_9448,N_9385,N_9396);
nor U9449 (N_9449,N_9373,N_9377);
or U9450 (N_9450,N_9372,N_9229);
or U9451 (N_9451,N_9364,N_9207);
nand U9452 (N_9452,N_9347,N_9390);
and U9453 (N_9453,N_9234,N_9309);
xnor U9454 (N_9454,N_9253,N_9305);
nor U9455 (N_9455,N_9285,N_9210);
or U9456 (N_9456,N_9311,N_9350);
nor U9457 (N_9457,N_9357,N_9227);
or U9458 (N_9458,N_9272,N_9276);
nand U9459 (N_9459,N_9353,N_9299);
or U9460 (N_9460,N_9338,N_9295);
and U9461 (N_9461,N_9366,N_9256);
nor U9462 (N_9462,N_9233,N_9395);
nand U9463 (N_9463,N_9241,N_9278);
and U9464 (N_9464,N_9270,N_9391);
xnor U9465 (N_9465,N_9206,N_9317);
and U9466 (N_9466,N_9370,N_9324);
nor U9467 (N_9467,N_9386,N_9237);
nor U9468 (N_9468,N_9365,N_9330);
and U9469 (N_9469,N_9265,N_9288);
xor U9470 (N_9470,N_9296,N_9399);
xnor U9471 (N_9471,N_9398,N_9319);
xnor U9472 (N_9472,N_9316,N_9369);
nor U9473 (N_9473,N_9246,N_9300);
nor U9474 (N_9474,N_9238,N_9262);
nand U9475 (N_9475,N_9242,N_9258);
or U9476 (N_9476,N_9200,N_9306);
or U9477 (N_9477,N_9360,N_9349);
xor U9478 (N_9478,N_9380,N_9212);
nand U9479 (N_9479,N_9361,N_9304);
or U9480 (N_9480,N_9239,N_9235);
xnor U9481 (N_9481,N_9362,N_9228);
or U9482 (N_9482,N_9355,N_9374);
nand U9483 (N_9483,N_9358,N_9371);
xor U9484 (N_9484,N_9273,N_9289);
nand U9485 (N_9485,N_9223,N_9388);
xnor U9486 (N_9486,N_9220,N_9384);
nand U9487 (N_9487,N_9201,N_9363);
nor U9488 (N_9488,N_9236,N_9308);
nor U9489 (N_9489,N_9394,N_9343);
nor U9490 (N_9490,N_9266,N_9334);
or U9491 (N_9491,N_9290,N_9260);
nand U9492 (N_9492,N_9321,N_9341);
nor U9493 (N_9493,N_9244,N_9215);
xor U9494 (N_9494,N_9213,N_9267);
nor U9495 (N_9495,N_9211,N_9274);
and U9496 (N_9496,N_9379,N_9269);
xnor U9497 (N_9497,N_9232,N_9389);
and U9498 (N_9498,N_9332,N_9302);
nand U9499 (N_9499,N_9218,N_9254);
nand U9500 (N_9500,N_9342,N_9327);
and U9501 (N_9501,N_9211,N_9371);
or U9502 (N_9502,N_9240,N_9270);
nor U9503 (N_9503,N_9215,N_9373);
nand U9504 (N_9504,N_9344,N_9320);
or U9505 (N_9505,N_9288,N_9377);
and U9506 (N_9506,N_9372,N_9274);
or U9507 (N_9507,N_9292,N_9249);
xor U9508 (N_9508,N_9371,N_9308);
nor U9509 (N_9509,N_9375,N_9205);
and U9510 (N_9510,N_9248,N_9294);
or U9511 (N_9511,N_9345,N_9239);
nor U9512 (N_9512,N_9318,N_9326);
nand U9513 (N_9513,N_9306,N_9295);
and U9514 (N_9514,N_9374,N_9202);
nor U9515 (N_9515,N_9378,N_9377);
or U9516 (N_9516,N_9211,N_9276);
or U9517 (N_9517,N_9383,N_9211);
or U9518 (N_9518,N_9241,N_9237);
and U9519 (N_9519,N_9287,N_9397);
or U9520 (N_9520,N_9270,N_9392);
and U9521 (N_9521,N_9333,N_9383);
nand U9522 (N_9522,N_9292,N_9208);
xor U9523 (N_9523,N_9324,N_9249);
nor U9524 (N_9524,N_9216,N_9351);
and U9525 (N_9525,N_9364,N_9226);
or U9526 (N_9526,N_9336,N_9202);
nand U9527 (N_9527,N_9252,N_9351);
nand U9528 (N_9528,N_9312,N_9343);
nand U9529 (N_9529,N_9220,N_9355);
nor U9530 (N_9530,N_9395,N_9271);
nor U9531 (N_9531,N_9217,N_9280);
nand U9532 (N_9532,N_9396,N_9339);
and U9533 (N_9533,N_9296,N_9349);
xor U9534 (N_9534,N_9234,N_9382);
or U9535 (N_9535,N_9211,N_9234);
and U9536 (N_9536,N_9373,N_9260);
and U9537 (N_9537,N_9300,N_9238);
or U9538 (N_9538,N_9289,N_9296);
xnor U9539 (N_9539,N_9273,N_9363);
nand U9540 (N_9540,N_9337,N_9343);
xnor U9541 (N_9541,N_9386,N_9231);
nor U9542 (N_9542,N_9334,N_9362);
xnor U9543 (N_9543,N_9298,N_9327);
and U9544 (N_9544,N_9375,N_9244);
or U9545 (N_9545,N_9264,N_9341);
nor U9546 (N_9546,N_9343,N_9331);
nand U9547 (N_9547,N_9221,N_9314);
nand U9548 (N_9548,N_9327,N_9228);
or U9549 (N_9549,N_9351,N_9390);
xnor U9550 (N_9550,N_9276,N_9249);
and U9551 (N_9551,N_9370,N_9332);
nor U9552 (N_9552,N_9326,N_9244);
nand U9553 (N_9553,N_9218,N_9245);
xor U9554 (N_9554,N_9232,N_9384);
nand U9555 (N_9555,N_9216,N_9281);
xor U9556 (N_9556,N_9370,N_9204);
nor U9557 (N_9557,N_9310,N_9230);
and U9558 (N_9558,N_9236,N_9298);
nor U9559 (N_9559,N_9273,N_9298);
xnor U9560 (N_9560,N_9349,N_9269);
xor U9561 (N_9561,N_9247,N_9385);
xor U9562 (N_9562,N_9288,N_9362);
nand U9563 (N_9563,N_9305,N_9378);
nand U9564 (N_9564,N_9278,N_9315);
nor U9565 (N_9565,N_9373,N_9285);
and U9566 (N_9566,N_9393,N_9321);
and U9567 (N_9567,N_9223,N_9205);
xnor U9568 (N_9568,N_9263,N_9314);
nor U9569 (N_9569,N_9217,N_9224);
and U9570 (N_9570,N_9253,N_9359);
and U9571 (N_9571,N_9269,N_9251);
nand U9572 (N_9572,N_9262,N_9229);
nand U9573 (N_9573,N_9264,N_9340);
nor U9574 (N_9574,N_9384,N_9355);
xnor U9575 (N_9575,N_9298,N_9395);
and U9576 (N_9576,N_9295,N_9398);
or U9577 (N_9577,N_9371,N_9396);
and U9578 (N_9578,N_9292,N_9379);
nand U9579 (N_9579,N_9313,N_9394);
xnor U9580 (N_9580,N_9313,N_9334);
and U9581 (N_9581,N_9358,N_9384);
or U9582 (N_9582,N_9319,N_9220);
nor U9583 (N_9583,N_9343,N_9305);
and U9584 (N_9584,N_9375,N_9337);
nand U9585 (N_9585,N_9237,N_9321);
or U9586 (N_9586,N_9334,N_9298);
nand U9587 (N_9587,N_9245,N_9247);
and U9588 (N_9588,N_9350,N_9339);
and U9589 (N_9589,N_9331,N_9373);
and U9590 (N_9590,N_9303,N_9318);
and U9591 (N_9591,N_9329,N_9304);
nand U9592 (N_9592,N_9273,N_9200);
nor U9593 (N_9593,N_9257,N_9239);
xnor U9594 (N_9594,N_9345,N_9368);
or U9595 (N_9595,N_9368,N_9207);
nor U9596 (N_9596,N_9210,N_9283);
xor U9597 (N_9597,N_9219,N_9255);
xnor U9598 (N_9598,N_9345,N_9233);
nor U9599 (N_9599,N_9295,N_9299);
nor U9600 (N_9600,N_9457,N_9475);
nand U9601 (N_9601,N_9551,N_9554);
or U9602 (N_9602,N_9435,N_9413);
xnor U9603 (N_9603,N_9584,N_9522);
and U9604 (N_9604,N_9410,N_9478);
nor U9605 (N_9605,N_9582,N_9425);
xor U9606 (N_9606,N_9568,N_9552);
and U9607 (N_9607,N_9585,N_9456);
and U9608 (N_9608,N_9524,N_9485);
and U9609 (N_9609,N_9559,N_9437);
nand U9610 (N_9610,N_9495,N_9556);
xor U9611 (N_9611,N_9521,N_9569);
nor U9612 (N_9612,N_9581,N_9484);
or U9613 (N_9613,N_9507,N_9498);
nor U9614 (N_9614,N_9586,N_9451);
nor U9615 (N_9615,N_9492,N_9563);
or U9616 (N_9616,N_9543,N_9516);
nand U9617 (N_9617,N_9580,N_9481);
and U9618 (N_9618,N_9578,N_9421);
nand U9619 (N_9619,N_9547,N_9414);
or U9620 (N_9620,N_9434,N_9509);
and U9621 (N_9621,N_9549,N_9426);
xor U9622 (N_9622,N_9428,N_9496);
and U9623 (N_9623,N_9400,N_9419);
or U9624 (N_9624,N_9598,N_9473);
nor U9625 (N_9625,N_9486,N_9430);
nor U9626 (N_9626,N_9594,N_9560);
nor U9627 (N_9627,N_9442,N_9561);
xor U9628 (N_9628,N_9511,N_9577);
nor U9629 (N_9629,N_9592,N_9520);
or U9630 (N_9630,N_9534,N_9401);
nor U9631 (N_9631,N_9490,N_9468);
nand U9632 (N_9632,N_9503,N_9440);
or U9633 (N_9633,N_9494,N_9469);
or U9634 (N_9634,N_9436,N_9542);
xor U9635 (N_9635,N_9593,N_9525);
and U9636 (N_9636,N_9429,N_9504);
nor U9637 (N_9637,N_9596,N_9589);
and U9638 (N_9638,N_9449,N_9512);
or U9639 (N_9639,N_9579,N_9446);
nand U9640 (N_9640,N_9573,N_9567);
xor U9641 (N_9641,N_9443,N_9477);
or U9642 (N_9642,N_9572,N_9450);
nor U9643 (N_9643,N_9583,N_9487);
nor U9644 (N_9644,N_9558,N_9408);
nor U9645 (N_9645,N_9523,N_9452);
nand U9646 (N_9646,N_9555,N_9590);
nand U9647 (N_9647,N_9424,N_9566);
or U9648 (N_9648,N_9447,N_9538);
nand U9649 (N_9649,N_9467,N_9576);
and U9650 (N_9650,N_9459,N_9497);
nand U9651 (N_9651,N_9412,N_9541);
xnor U9652 (N_9652,N_9407,N_9518);
nand U9653 (N_9653,N_9420,N_9545);
or U9654 (N_9654,N_9553,N_9570);
nor U9655 (N_9655,N_9409,N_9448);
nor U9656 (N_9656,N_9532,N_9445);
or U9657 (N_9657,N_9453,N_9533);
nand U9658 (N_9658,N_9539,N_9438);
and U9659 (N_9659,N_9432,N_9535);
nor U9660 (N_9660,N_9544,N_9406);
and U9661 (N_9661,N_9489,N_9422);
nor U9662 (N_9662,N_9471,N_9427);
nor U9663 (N_9663,N_9500,N_9527);
nand U9664 (N_9664,N_9595,N_9415);
or U9665 (N_9665,N_9506,N_9565);
nand U9666 (N_9666,N_9441,N_9465);
xnor U9667 (N_9667,N_9405,N_9529);
and U9668 (N_9668,N_9530,N_9466);
xnor U9669 (N_9669,N_9433,N_9528);
nand U9670 (N_9670,N_9536,N_9423);
nand U9671 (N_9671,N_9562,N_9548);
xor U9672 (N_9672,N_9479,N_9411);
and U9673 (N_9673,N_9482,N_9502);
or U9674 (N_9674,N_9472,N_9460);
or U9675 (N_9675,N_9513,N_9404);
nor U9676 (N_9676,N_9455,N_9458);
nor U9677 (N_9677,N_9588,N_9597);
or U9678 (N_9678,N_9474,N_9515);
and U9679 (N_9679,N_9461,N_9462);
or U9680 (N_9680,N_9463,N_9416);
or U9681 (N_9681,N_9564,N_9499);
and U9682 (N_9682,N_9508,N_9480);
nand U9683 (N_9683,N_9537,N_9403);
nand U9684 (N_9684,N_9571,N_9575);
nand U9685 (N_9685,N_9476,N_9402);
nand U9686 (N_9686,N_9483,N_9439);
nand U9687 (N_9687,N_9493,N_9519);
xor U9688 (N_9688,N_9454,N_9491);
or U9689 (N_9689,N_9587,N_9488);
nor U9690 (N_9690,N_9599,N_9444);
nor U9691 (N_9691,N_9550,N_9417);
nand U9692 (N_9692,N_9531,N_9557);
nor U9693 (N_9693,N_9546,N_9501);
nor U9694 (N_9694,N_9505,N_9464);
xor U9695 (N_9695,N_9510,N_9591);
xor U9696 (N_9696,N_9470,N_9540);
nand U9697 (N_9697,N_9431,N_9514);
xnor U9698 (N_9698,N_9526,N_9418);
nand U9699 (N_9699,N_9574,N_9517);
nor U9700 (N_9700,N_9591,N_9516);
nand U9701 (N_9701,N_9429,N_9500);
or U9702 (N_9702,N_9427,N_9494);
nor U9703 (N_9703,N_9448,N_9539);
nor U9704 (N_9704,N_9401,N_9494);
nand U9705 (N_9705,N_9436,N_9559);
xor U9706 (N_9706,N_9528,N_9465);
and U9707 (N_9707,N_9553,N_9426);
nand U9708 (N_9708,N_9521,N_9562);
or U9709 (N_9709,N_9560,N_9555);
xnor U9710 (N_9710,N_9585,N_9449);
xor U9711 (N_9711,N_9511,N_9456);
or U9712 (N_9712,N_9508,N_9529);
nor U9713 (N_9713,N_9472,N_9438);
nor U9714 (N_9714,N_9536,N_9576);
nand U9715 (N_9715,N_9429,N_9562);
or U9716 (N_9716,N_9520,N_9545);
nor U9717 (N_9717,N_9420,N_9587);
xor U9718 (N_9718,N_9545,N_9406);
nor U9719 (N_9719,N_9427,N_9450);
or U9720 (N_9720,N_9414,N_9420);
nand U9721 (N_9721,N_9562,N_9434);
nand U9722 (N_9722,N_9569,N_9550);
and U9723 (N_9723,N_9591,N_9452);
nand U9724 (N_9724,N_9565,N_9550);
and U9725 (N_9725,N_9567,N_9437);
nor U9726 (N_9726,N_9580,N_9484);
or U9727 (N_9727,N_9576,N_9514);
nor U9728 (N_9728,N_9562,N_9540);
nor U9729 (N_9729,N_9447,N_9499);
and U9730 (N_9730,N_9459,N_9435);
xor U9731 (N_9731,N_9420,N_9425);
nand U9732 (N_9732,N_9432,N_9515);
nor U9733 (N_9733,N_9421,N_9597);
and U9734 (N_9734,N_9580,N_9450);
and U9735 (N_9735,N_9559,N_9446);
nand U9736 (N_9736,N_9481,N_9487);
xor U9737 (N_9737,N_9540,N_9558);
nor U9738 (N_9738,N_9521,N_9417);
or U9739 (N_9739,N_9512,N_9535);
nor U9740 (N_9740,N_9414,N_9470);
nand U9741 (N_9741,N_9439,N_9475);
or U9742 (N_9742,N_9556,N_9488);
nand U9743 (N_9743,N_9529,N_9441);
or U9744 (N_9744,N_9413,N_9547);
xnor U9745 (N_9745,N_9476,N_9529);
nor U9746 (N_9746,N_9406,N_9531);
nand U9747 (N_9747,N_9483,N_9482);
or U9748 (N_9748,N_9480,N_9446);
nand U9749 (N_9749,N_9521,N_9506);
nand U9750 (N_9750,N_9401,N_9573);
nor U9751 (N_9751,N_9514,N_9445);
xnor U9752 (N_9752,N_9513,N_9422);
and U9753 (N_9753,N_9406,N_9569);
or U9754 (N_9754,N_9494,N_9503);
nor U9755 (N_9755,N_9563,N_9528);
nand U9756 (N_9756,N_9567,N_9551);
xnor U9757 (N_9757,N_9510,N_9468);
and U9758 (N_9758,N_9566,N_9538);
and U9759 (N_9759,N_9598,N_9515);
nand U9760 (N_9760,N_9587,N_9483);
nand U9761 (N_9761,N_9484,N_9477);
nand U9762 (N_9762,N_9482,N_9471);
and U9763 (N_9763,N_9461,N_9465);
xor U9764 (N_9764,N_9574,N_9590);
nor U9765 (N_9765,N_9530,N_9566);
and U9766 (N_9766,N_9536,N_9421);
nor U9767 (N_9767,N_9575,N_9591);
and U9768 (N_9768,N_9549,N_9458);
or U9769 (N_9769,N_9517,N_9576);
or U9770 (N_9770,N_9441,N_9412);
nand U9771 (N_9771,N_9445,N_9428);
or U9772 (N_9772,N_9544,N_9536);
or U9773 (N_9773,N_9413,N_9582);
and U9774 (N_9774,N_9555,N_9557);
nand U9775 (N_9775,N_9568,N_9583);
nand U9776 (N_9776,N_9530,N_9559);
and U9777 (N_9777,N_9545,N_9462);
nor U9778 (N_9778,N_9439,N_9570);
xnor U9779 (N_9779,N_9556,N_9499);
and U9780 (N_9780,N_9507,N_9531);
or U9781 (N_9781,N_9552,N_9456);
xor U9782 (N_9782,N_9590,N_9588);
nor U9783 (N_9783,N_9533,N_9442);
or U9784 (N_9784,N_9412,N_9559);
or U9785 (N_9785,N_9575,N_9463);
or U9786 (N_9786,N_9508,N_9598);
or U9787 (N_9787,N_9464,N_9483);
nor U9788 (N_9788,N_9440,N_9557);
or U9789 (N_9789,N_9562,N_9519);
nand U9790 (N_9790,N_9400,N_9459);
or U9791 (N_9791,N_9466,N_9423);
nand U9792 (N_9792,N_9507,N_9597);
nand U9793 (N_9793,N_9445,N_9451);
and U9794 (N_9794,N_9452,N_9551);
nand U9795 (N_9795,N_9596,N_9400);
nand U9796 (N_9796,N_9563,N_9529);
or U9797 (N_9797,N_9562,N_9589);
nor U9798 (N_9798,N_9589,N_9587);
nor U9799 (N_9799,N_9468,N_9593);
nand U9800 (N_9800,N_9676,N_9724);
nor U9801 (N_9801,N_9601,N_9710);
and U9802 (N_9802,N_9618,N_9786);
and U9803 (N_9803,N_9721,N_9625);
nor U9804 (N_9804,N_9739,N_9667);
nor U9805 (N_9805,N_9619,N_9797);
nand U9806 (N_9806,N_9778,N_9622);
or U9807 (N_9807,N_9736,N_9730);
or U9808 (N_9808,N_9678,N_9604);
nand U9809 (N_9809,N_9712,N_9783);
and U9810 (N_9810,N_9767,N_9615);
xnor U9811 (N_9811,N_9654,N_9706);
or U9812 (N_9812,N_9629,N_9715);
and U9813 (N_9813,N_9745,N_9791);
nand U9814 (N_9814,N_9661,N_9703);
xnor U9815 (N_9815,N_9610,N_9764);
or U9816 (N_9816,N_9699,N_9662);
and U9817 (N_9817,N_9691,N_9673);
xnor U9818 (N_9818,N_9748,N_9686);
xnor U9819 (N_9819,N_9746,N_9643);
and U9820 (N_9820,N_9663,N_9749);
nand U9821 (N_9821,N_9747,N_9689);
nor U9822 (N_9822,N_9755,N_9688);
and U9823 (N_9823,N_9696,N_9626);
or U9824 (N_9824,N_9693,N_9718);
nand U9825 (N_9825,N_9633,N_9717);
xor U9826 (N_9826,N_9731,N_9640);
and U9827 (N_9827,N_9639,N_9621);
nor U9828 (N_9828,N_9762,N_9743);
nand U9829 (N_9829,N_9741,N_9641);
or U9830 (N_9830,N_9628,N_9729);
nand U9831 (N_9831,N_9790,N_9714);
nor U9832 (N_9832,N_9716,N_9702);
and U9833 (N_9833,N_9675,N_9700);
and U9834 (N_9834,N_9726,N_9649);
nand U9835 (N_9835,N_9612,N_9770);
nor U9836 (N_9836,N_9658,N_9734);
or U9837 (N_9837,N_9723,N_9757);
or U9838 (N_9838,N_9728,N_9793);
and U9839 (N_9839,N_9759,N_9634);
or U9840 (N_9840,N_9738,N_9682);
nor U9841 (N_9841,N_9630,N_9735);
or U9842 (N_9842,N_9613,N_9646);
nor U9843 (N_9843,N_9653,N_9701);
nor U9844 (N_9844,N_9668,N_9644);
or U9845 (N_9845,N_9680,N_9695);
xor U9846 (N_9846,N_9677,N_9685);
nand U9847 (N_9847,N_9608,N_9664);
xnor U9848 (N_9848,N_9611,N_9674);
nor U9849 (N_9849,N_9697,N_9733);
nand U9850 (N_9850,N_9623,N_9707);
and U9851 (N_9851,N_9636,N_9788);
nand U9852 (N_9852,N_9624,N_9627);
nand U9853 (N_9853,N_9792,N_9616);
and U9854 (N_9854,N_9765,N_9799);
nand U9855 (N_9855,N_9603,N_9719);
and U9856 (N_9856,N_9698,N_9672);
and U9857 (N_9857,N_9725,N_9766);
xnor U9858 (N_9858,N_9752,N_9768);
or U9859 (N_9859,N_9774,N_9796);
nor U9860 (N_9860,N_9781,N_9687);
nand U9861 (N_9861,N_9750,N_9681);
xnor U9862 (N_9862,N_9775,N_9751);
xnor U9863 (N_9863,N_9671,N_9660);
xor U9864 (N_9864,N_9753,N_9650);
and U9865 (N_9865,N_9690,N_9784);
xor U9866 (N_9866,N_9787,N_9694);
nand U9867 (N_9867,N_9760,N_9679);
or U9868 (N_9868,N_9683,N_9756);
or U9869 (N_9869,N_9656,N_9722);
and U9870 (N_9870,N_9794,N_9665);
nor U9871 (N_9871,N_9727,N_9772);
or U9872 (N_9872,N_9705,N_9684);
xnor U9873 (N_9873,N_9773,N_9637);
nand U9874 (N_9874,N_9744,N_9614);
nor U9875 (N_9875,N_9645,N_9789);
nand U9876 (N_9876,N_9754,N_9607);
nand U9877 (N_9877,N_9651,N_9779);
and U9878 (N_9878,N_9620,N_9666);
nor U9879 (N_9879,N_9708,N_9777);
or U9880 (N_9880,N_9670,N_9655);
nand U9881 (N_9881,N_9758,N_9659);
nor U9882 (N_9882,N_9776,N_9692);
nor U9883 (N_9883,N_9648,N_9711);
nand U9884 (N_9884,N_9647,N_9771);
nor U9885 (N_9885,N_9600,N_9669);
and U9886 (N_9886,N_9642,N_9785);
nand U9887 (N_9887,N_9761,N_9605);
or U9888 (N_9888,N_9795,N_9609);
nor U9889 (N_9889,N_9657,N_9635);
nand U9890 (N_9890,N_9732,N_9737);
and U9891 (N_9891,N_9631,N_9780);
nor U9892 (N_9892,N_9720,N_9713);
nand U9893 (N_9893,N_9602,N_9606);
or U9894 (N_9894,N_9638,N_9704);
nor U9895 (N_9895,N_9769,N_9740);
and U9896 (N_9896,N_9782,N_9632);
nor U9897 (N_9897,N_9652,N_9798);
nand U9898 (N_9898,N_9709,N_9763);
xor U9899 (N_9899,N_9617,N_9742);
and U9900 (N_9900,N_9708,N_9635);
xor U9901 (N_9901,N_9727,N_9622);
and U9902 (N_9902,N_9776,N_9756);
xor U9903 (N_9903,N_9676,N_9718);
nand U9904 (N_9904,N_9699,N_9738);
nor U9905 (N_9905,N_9739,N_9769);
xnor U9906 (N_9906,N_9623,N_9635);
or U9907 (N_9907,N_9632,N_9645);
and U9908 (N_9908,N_9782,N_9737);
and U9909 (N_9909,N_9603,N_9742);
nor U9910 (N_9910,N_9790,N_9671);
xor U9911 (N_9911,N_9653,N_9767);
or U9912 (N_9912,N_9663,N_9781);
nand U9913 (N_9913,N_9617,N_9607);
nand U9914 (N_9914,N_9764,N_9767);
nor U9915 (N_9915,N_9759,N_9606);
or U9916 (N_9916,N_9792,N_9742);
and U9917 (N_9917,N_9711,N_9733);
or U9918 (N_9918,N_9667,N_9794);
nor U9919 (N_9919,N_9748,N_9779);
xnor U9920 (N_9920,N_9781,N_9612);
nor U9921 (N_9921,N_9769,N_9782);
nor U9922 (N_9922,N_9658,N_9614);
nand U9923 (N_9923,N_9695,N_9606);
nand U9924 (N_9924,N_9705,N_9787);
nor U9925 (N_9925,N_9742,N_9645);
or U9926 (N_9926,N_9700,N_9713);
xor U9927 (N_9927,N_9712,N_9671);
or U9928 (N_9928,N_9658,N_9627);
nand U9929 (N_9929,N_9726,N_9701);
and U9930 (N_9930,N_9751,N_9730);
nand U9931 (N_9931,N_9745,N_9659);
nor U9932 (N_9932,N_9697,N_9764);
or U9933 (N_9933,N_9744,N_9780);
and U9934 (N_9934,N_9709,N_9679);
nand U9935 (N_9935,N_9673,N_9799);
and U9936 (N_9936,N_9608,N_9634);
xor U9937 (N_9937,N_9792,N_9722);
and U9938 (N_9938,N_9675,N_9752);
nor U9939 (N_9939,N_9784,N_9731);
xor U9940 (N_9940,N_9660,N_9651);
nand U9941 (N_9941,N_9732,N_9691);
xnor U9942 (N_9942,N_9743,N_9752);
or U9943 (N_9943,N_9780,N_9646);
and U9944 (N_9944,N_9738,N_9799);
xnor U9945 (N_9945,N_9662,N_9794);
or U9946 (N_9946,N_9765,N_9627);
xnor U9947 (N_9947,N_9775,N_9636);
nand U9948 (N_9948,N_9629,N_9735);
nand U9949 (N_9949,N_9618,N_9712);
and U9950 (N_9950,N_9608,N_9739);
and U9951 (N_9951,N_9640,N_9720);
and U9952 (N_9952,N_9630,N_9650);
nand U9953 (N_9953,N_9693,N_9798);
xnor U9954 (N_9954,N_9698,N_9720);
nand U9955 (N_9955,N_9632,N_9691);
and U9956 (N_9956,N_9610,N_9686);
nand U9957 (N_9957,N_9610,N_9796);
nor U9958 (N_9958,N_9772,N_9734);
nor U9959 (N_9959,N_9797,N_9612);
and U9960 (N_9960,N_9758,N_9646);
and U9961 (N_9961,N_9727,N_9696);
xnor U9962 (N_9962,N_9669,N_9769);
nand U9963 (N_9963,N_9631,N_9671);
nand U9964 (N_9964,N_9757,N_9612);
and U9965 (N_9965,N_9798,N_9625);
or U9966 (N_9966,N_9662,N_9611);
xor U9967 (N_9967,N_9744,N_9612);
nand U9968 (N_9968,N_9625,N_9760);
nor U9969 (N_9969,N_9670,N_9618);
nor U9970 (N_9970,N_9655,N_9607);
and U9971 (N_9971,N_9604,N_9768);
nor U9972 (N_9972,N_9710,N_9641);
and U9973 (N_9973,N_9696,N_9634);
xnor U9974 (N_9974,N_9716,N_9666);
nand U9975 (N_9975,N_9740,N_9717);
nand U9976 (N_9976,N_9711,N_9795);
xor U9977 (N_9977,N_9605,N_9708);
nor U9978 (N_9978,N_9717,N_9642);
nand U9979 (N_9979,N_9771,N_9646);
nor U9980 (N_9980,N_9743,N_9624);
nand U9981 (N_9981,N_9709,N_9704);
nor U9982 (N_9982,N_9630,N_9722);
xor U9983 (N_9983,N_9648,N_9788);
xor U9984 (N_9984,N_9633,N_9642);
nor U9985 (N_9985,N_9673,N_9681);
xnor U9986 (N_9986,N_9605,N_9749);
and U9987 (N_9987,N_9600,N_9784);
and U9988 (N_9988,N_9679,N_9793);
nor U9989 (N_9989,N_9749,N_9766);
xor U9990 (N_9990,N_9761,N_9620);
nor U9991 (N_9991,N_9790,N_9720);
nor U9992 (N_9992,N_9711,N_9659);
xnor U9993 (N_9993,N_9609,N_9634);
or U9994 (N_9994,N_9652,N_9744);
and U9995 (N_9995,N_9691,N_9751);
xnor U9996 (N_9996,N_9634,N_9629);
nor U9997 (N_9997,N_9767,N_9715);
nor U9998 (N_9998,N_9784,N_9632);
and U9999 (N_9999,N_9666,N_9745);
and UO_0 (O_0,N_9924,N_9995);
nor UO_1 (O_1,N_9834,N_9832);
xor UO_2 (O_2,N_9849,N_9983);
nor UO_3 (O_3,N_9926,N_9816);
and UO_4 (O_4,N_9889,N_9967);
nand UO_5 (O_5,N_9996,N_9809);
nor UO_6 (O_6,N_9878,N_9961);
xor UO_7 (O_7,N_9846,N_9979);
or UO_8 (O_8,N_9981,N_9851);
nand UO_9 (O_9,N_9930,N_9971);
or UO_10 (O_10,N_9828,N_9937);
nand UO_11 (O_11,N_9897,N_9959);
xnor UO_12 (O_12,N_9942,N_9812);
nand UO_13 (O_13,N_9974,N_9975);
and UO_14 (O_14,N_9847,N_9839);
or UO_15 (O_15,N_9892,N_9802);
nor UO_16 (O_16,N_9808,N_9820);
nor UO_17 (O_17,N_9989,N_9840);
xnor UO_18 (O_18,N_9841,N_9919);
nor UO_19 (O_19,N_9998,N_9933);
and UO_20 (O_20,N_9883,N_9817);
nor UO_21 (O_21,N_9973,N_9870);
nand UO_22 (O_22,N_9899,N_9922);
nor UO_23 (O_23,N_9944,N_9850);
nand UO_24 (O_24,N_9943,N_9913);
and UO_25 (O_25,N_9806,N_9985);
nand UO_26 (O_26,N_9845,N_9904);
xor UO_27 (O_27,N_9986,N_9852);
xor UO_28 (O_28,N_9823,N_9950);
and UO_29 (O_29,N_9821,N_9838);
xnor UO_30 (O_30,N_9928,N_9854);
nor UO_31 (O_31,N_9881,N_9934);
nor UO_32 (O_32,N_9970,N_9819);
nor UO_33 (O_33,N_9916,N_9874);
nand UO_34 (O_34,N_9826,N_9818);
or UO_35 (O_35,N_9984,N_9861);
nor UO_36 (O_36,N_9936,N_9927);
xnor UO_37 (O_37,N_9805,N_9946);
and UO_38 (O_38,N_9945,N_9992);
nor UO_39 (O_39,N_9814,N_9887);
nor UO_40 (O_40,N_9864,N_9896);
nor UO_41 (O_41,N_9910,N_9906);
nor UO_42 (O_42,N_9857,N_9925);
nand UO_43 (O_43,N_9859,N_9835);
nand UO_44 (O_44,N_9932,N_9994);
nand UO_45 (O_45,N_9949,N_9954);
or UO_46 (O_46,N_9844,N_9825);
xor UO_47 (O_47,N_9873,N_9968);
xor UO_48 (O_48,N_9856,N_9865);
nor UO_49 (O_49,N_9813,N_9914);
and UO_50 (O_50,N_9958,N_9831);
xnor UO_51 (O_51,N_9898,N_9941);
or UO_52 (O_52,N_9888,N_9929);
and UO_53 (O_53,N_9908,N_9901);
and UO_54 (O_54,N_9980,N_9885);
or UO_55 (O_55,N_9939,N_9807);
or UO_56 (O_56,N_9991,N_9977);
nor UO_57 (O_57,N_9960,N_9827);
xor UO_58 (O_58,N_9804,N_9976);
nor UO_59 (O_59,N_9911,N_9900);
nand UO_60 (O_60,N_9858,N_9947);
nor UO_61 (O_61,N_9871,N_9833);
nor UO_62 (O_62,N_9867,N_9902);
nand UO_63 (O_63,N_9921,N_9917);
xor UO_64 (O_64,N_9877,N_9955);
or UO_65 (O_65,N_9890,N_9811);
nand UO_66 (O_66,N_9956,N_9803);
and UO_67 (O_67,N_9999,N_9969);
nor UO_68 (O_68,N_9882,N_9993);
and UO_69 (O_69,N_9903,N_9951);
xnor UO_70 (O_70,N_9815,N_9810);
xnor UO_71 (O_71,N_9886,N_9907);
or UO_72 (O_72,N_9876,N_9872);
xor UO_73 (O_73,N_9836,N_9931);
or UO_74 (O_74,N_9863,N_9909);
and UO_75 (O_75,N_9895,N_9866);
xor UO_76 (O_76,N_9966,N_9972);
xor UO_77 (O_77,N_9920,N_9990);
xnor UO_78 (O_78,N_9860,N_9848);
xnor UO_79 (O_79,N_9963,N_9997);
nor UO_80 (O_80,N_9822,N_9893);
and UO_81 (O_81,N_9869,N_9862);
or UO_82 (O_82,N_9801,N_9800);
xnor UO_83 (O_83,N_9829,N_9875);
and UO_84 (O_84,N_9978,N_9957);
and UO_85 (O_85,N_9938,N_9964);
nand UO_86 (O_86,N_9824,N_9915);
nor UO_87 (O_87,N_9918,N_9843);
nand UO_88 (O_88,N_9982,N_9940);
and UO_89 (O_89,N_9948,N_9853);
nor UO_90 (O_90,N_9953,N_9935);
xor UO_91 (O_91,N_9855,N_9837);
nand UO_92 (O_92,N_9965,N_9880);
or UO_93 (O_93,N_9905,N_9987);
or UO_94 (O_94,N_9923,N_9842);
xor UO_95 (O_95,N_9988,N_9879);
xnor UO_96 (O_96,N_9894,N_9912);
or UO_97 (O_97,N_9830,N_9952);
nand UO_98 (O_98,N_9868,N_9884);
nand UO_99 (O_99,N_9891,N_9962);
and UO_100 (O_100,N_9961,N_9966);
or UO_101 (O_101,N_9869,N_9851);
xor UO_102 (O_102,N_9902,N_9828);
or UO_103 (O_103,N_9930,N_9963);
nand UO_104 (O_104,N_9966,N_9876);
nor UO_105 (O_105,N_9825,N_9994);
xnor UO_106 (O_106,N_9969,N_9952);
nor UO_107 (O_107,N_9868,N_9912);
nand UO_108 (O_108,N_9933,N_9834);
and UO_109 (O_109,N_9996,N_9911);
and UO_110 (O_110,N_9992,N_9897);
or UO_111 (O_111,N_9976,N_9805);
xnor UO_112 (O_112,N_9822,N_9912);
xor UO_113 (O_113,N_9811,N_9858);
xor UO_114 (O_114,N_9927,N_9825);
nor UO_115 (O_115,N_9857,N_9829);
nor UO_116 (O_116,N_9865,N_9834);
xor UO_117 (O_117,N_9965,N_9857);
and UO_118 (O_118,N_9931,N_9823);
and UO_119 (O_119,N_9960,N_9808);
xor UO_120 (O_120,N_9830,N_9899);
or UO_121 (O_121,N_9993,N_9843);
or UO_122 (O_122,N_9908,N_9837);
or UO_123 (O_123,N_9805,N_9807);
xor UO_124 (O_124,N_9950,N_9927);
or UO_125 (O_125,N_9920,N_9868);
or UO_126 (O_126,N_9966,N_9834);
xor UO_127 (O_127,N_9890,N_9888);
xor UO_128 (O_128,N_9908,N_9875);
nor UO_129 (O_129,N_9903,N_9978);
or UO_130 (O_130,N_9898,N_9929);
and UO_131 (O_131,N_9814,N_9927);
nor UO_132 (O_132,N_9902,N_9913);
xor UO_133 (O_133,N_9893,N_9961);
nor UO_134 (O_134,N_9998,N_9906);
nand UO_135 (O_135,N_9809,N_9831);
and UO_136 (O_136,N_9927,N_9879);
and UO_137 (O_137,N_9939,N_9956);
or UO_138 (O_138,N_9874,N_9844);
xnor UO_139 (O_139,N_9806,N_9904);
xor UO_140 (O_140,N_9932,N_9927);
nor UO_141 (O_141,N_9954,N_9881);
xor UO_142 (O_142,N_9834,N_9857);
nand UO_143 (O_143,N_9971,N_9893);
nor UO_144 (O_144,N_9860,N_9914);
xnor UO_145 (O_145,N_9810,N_9848);
and UO_146 (O_146,N_9839,N_9879);
xor UO_147 (O_147,N_9869,N_9863);
nor UO_148 (O_148,N_9961,N_9850);
xnor UO_149 (O_149,N_9836,N_9976);
nand UO_150 (O_150,N_9930,N_9972);
nor UO_151 (O_151,N_9934,N_9800);
xor UO_152 (O_152,N_9801,N_9908);
or UO_153 (O_153,N_9875,N_9889);
nand UO_154 (O_154,N_9867,N_9972);
and UO_155 (O_155,N_9965,N_9824);
xnor UO_156 (O_156,N_9955,N_9843);
or UO_157 (O_157,N_9930,N_9941);
xnor UO_158 (O_158,N_9951,N_9839);
nor UO_159 (O_159,N_9840,N_9804);
nand UO_160 (O_160,N_9970,N_9866);
and UO_161 (O_161,N_9930,N_9973);
xor UO_162 (O_162,N_9930,N_9936);
nand UO_163 (O_163,N_9883,N_9830);
xor UO_164 (O_164,N_9869,N_9809);
xnor UO_165 (O_165,N_9812,N_9826);
xnor UO_166 (O_166,N_9849,N_9996);
or UO_167 (O_167,N_9942,N_9863);
nand UO_168 (O_168,N_9911,N_9939);
or UO_169 (O_169,N_9917,N_9943);
or UO_170 (O_170,N_9970,N_9805);
and UO_171 (O_171,N_9834,N_9946);
and UO_172 (O_172,N_9821,N_9910);
xor UO_173 (O_173,N_9879,N_9962);
nor UO_174 (O_174,N_9842,N_9807);
nand UO_175 (O_175,N_9863,N_9977);
and UO_176 (O_176,N_9970,N_9846);
xor UO_177 (O_177,N_9954,N_9873);
xor UO_178 (O_178,N_9948,N_9930);
and UO_179 (O_179,N_9903,N_9860);
xnor UO_180 (O_180,N_9991,N_9902);
nor UO_181 (O_181,N_9819,N_9955);
nand UO_182 (O_182,N_9803,N_9939);
or UO_183 (O_183,N_9881,N_9807);
nand UO_184 (O_184,N_9974,N_9811);
nor UO_185 (O_185,N_9861,N_9822);
xor UO_186 (O_186,N_9982,N_9845);
or UO_187 (O_187,N_9958,N_9866);
or UO_188 (O_188,N_9996,N_9934);
nor UO_189 (O_189,N_9918,N_9804);
nand UO_190 (O_190,N_9848,N_9905);
and UO_191 (O_191,N_9909,N_9936);
and UO_192 (O_192,N_9815,N_9945);
and UO_193 (O_193,N_9933,N_9891);
xor UO_194 (O_194,N_9944,N_9912);
nand UO_195 (O_195,N_9983,N_9888);
xnor UO_196 (O_196,N_9904,N_9857);
nor UO_197 (O_197,N_9967,N_9997);
and UO_198 (O_198,N_9972,N_9932);
nor UO_199 (O_199,N_9942,N_9901);
or UO_200 (O_200,N_9898,N_9808);
or UO_201 (O_201,N_9964,N_9842);
nand UO_202 (O_202,N_9887,N_9812);
or UO_203 (O_203,N_9852,N_9933);
or UO_204 (O_204,N_9871,N_9986);
xnor UO_205 (O_205,N_9839,N_9807);
nand UO_206 (O_206,N_9909,N_9829);
or UO_207 (O_207,N_9892,N_9916);
nor UO_208 (O_208,N_9921,N_9868);
nand UO_209 (O_209,N_9997,N_9842);
nand UO_210 (O_210,N_9929,N_9985);
nand UO_211 (O_211,N_9957,N_9964);
xor UO_212 (O_212,N_9816,N_9972);
nor UO_213 (O_213,N_9986,N_9880);
or UO_214 (O_214,N_9804,N_9823);
nand UO_215 (O_215,N_9892,N_9834);
nor UO_216 (O_216,N_9961,N_9959);
nand UO_217 (O_217,N_9879,N_9830);
xnor UO_218 (O_218,N_9818,N_9807);
nand UO_219 (O_219,N_9911,N_9849);
nand UO_220 (O_220,N_9911,N_9827);
and UO_221 (O_221,N_9992,N_9867);
xor UO_222 (O_222,N_9904,N_9903);
nand UO_223 (O_223,N_9848,N_9910);
or UO_224 (O_224,N_9846,N_9852);
xnor UO_225 (O_225,N_9993,N_9881);
xnor UO_226 (O_226,N_9934,N_9900);
and UO_227 (O_227,N_9866,N_9800);
nor UO_228 (O_228,N_9918,N_9996);
or UO_229 (O_229,N_9883,N_9841);
nor UO_230 (O_230,N_9865,N_9992);
xor UO_231 (O_231,N_9965,N_9936);
nand UO_232 (O_232,N_9859,N_9801);
nand UO_233 (O_233,N_9907,N_9820);
nor UO_234 (O_234,N_9891,N_9879);
nand UO_235 (O_235,N_9819,N_9839);
nand UO_236 (O_236,N_9816,N_9909);
nand UO_237 (O_237,N_9950,N_9991);
nand UO_238 (O_238,N_9807,N_9936);
nor UO_239 (O_239,N_9869,N_9864);
nor UO_240 (O_240,N_9908,N_9835);
nor UO_241 (O_241,N_9847,N_9814);
nor UO_242 (O_242,N_9998,N_9905);
nand UO_243 (O_243,N_9964,N_9947);
and UO_244 (O_244,N_9820,N_9935);
xor UO_245 (O_245,N_9990,N_9985);
nand UO_246 (O_246,N_9943,N_9962);
nor UO_247 (O_247,N_9836,N_9969);
xor UO_248 (O_248,N_9889,N_9846);
and UO_249 (O_249,N_9816,N_9913);
xnor UO_250 (O_250,N_9852,N_9913);
or UO_251 (O_251,N_9829,N_9955);
nand UO_252 (O_252,N_9841,N_9832);
xor UO_253 (O_253,N_9891,N_9920);
and UO_254 (O_254,N_9866,N_9931);
nor UO_255 (O_255,N_9842,N_9932);
xnor UO_256 (O_256,N_9806,N_9828);
nand UO_257 (O_257,N_9839,N_9968);
or UO_258 (O_258,N_9958,N_9857);
and UO_259 (O_259,N_9876,N_9906);
nor UO_260 (O_260,N_9905,N_9861);
nor UO_261 (O_261,N_9832,N_9873);
or UO_262 (O_262,N_9953,N_9913);
and UO_263 (O_263,N_9829,N_9902);
or UO_264 (O_264,N_9919,N_9806);
and UO_265 (O_265,N_9803,N_9954);
and UO_266 (O_266,N_9892,N_9972);
and UO_267 (O_267,N_9859,N_9866);
xnor UO_268 (O_268,N_9898,N_9980);
nand UO_269 (O_269,N_9915,N_9938);
nand UO_270 (O_270,N_9979,N_9945);
or UO_271 (O_271,N_9825,N_9883);
xor UO_272 (O_272,N_9822,N_9844);
nand UO_273 (O_273,N_9898,N_9986);
xnor UO_274 (O_274,N_9875,N_9874);
nand UO_275 (O_275,N_9945,N_9919);
or UO_276 (O_276,N_9824,N_9922);
and UO_277 (O_277,N_9892,N_9897);
nor UO_278 (O_278,N_9909,N_9874);
or UO_279 (O_279,N_9932,N_9850);
xor UO_280 (O_280,N_9977,N_9952);
and UO_281 (O_281,N_9864,N_9807);
and UO_282 (O_282,N_9904,N_9828);
nor UO_283 (O_283,N_9920,N_9896);
xnor UO_284 (O_284,N_9842,N_9831);
and UO_285 (O_285,N_9906,N_9882);
or UO_286 (O_286,N_9829,N_9990);
and UO_287 (O_287,N_9918,N_9832);
xor UO_288 (O_288,N_9997,N_9864);
xnor UO_289 (O_289,N_9918,N_9830);
xor UO_290 (O_290,N_9989,N_9891);
nor UO_291 (O_291,N_9913,N_9911);
nor UO_292 (O_292,N_9974,N_9845);
and UO_293 (O_293,N_9851,N_9904);
xnor UO_294 (O_294,N_9815,N_9830);
nor UO_295 (O_295,N_9896,N_9841);
nand UO_296 (O_296,N_9979,N_9880);
and UO_297 (O_297,N_9984,N_9870);
or UO_298 (O_298,N_9882,N_9822);
xor UO_299 (O_299,N_9902,N_9883);
nand UO_300 (O_300,N_9917,N_9978);
xor UO_301 (O_301,N_9955,N_9867);
xor UO_302 (O_302,N_9944,N_9897);
and UO_303 (O_303,N_9974,N_9984);
nand UO_304 (O_304,N_9962,N_9846);
or UO_305 (O_305,N_9801,N_9897);
or UO_306 (O_306,N_9915,N_9870);
or UO_307 (O_307,N_9949,N_9887);
nor UO_308 (O_308,N_9978,N_9923);
and UO_309 (O_309,N_9926,N_9991);
and UO_310 (O_310,N_9924,N_9831);
or UO_311 (O_311,N_9901,N_9921);
nor UO_312 (O_312,N_9911,N_9940);
or UO_313 (O_313,N_9942,N_9804);
xnor UO_314 (O_314,N_9846,N_9948);
nor UO_315 (O_315,N_9930,N_9967);
xor UO_316 (O_316,N_9838,N_9899);
or UO_317 (O_317,N_9897,N_9893);
xnor UO_318 (O_318,N_9865,N_9988);
and UO_319 (O_319,N_9929,N_9801);
or UO_320 (O_320,N_9901,N_9988);
nor UO_321 (O_321,N_9978,N_9916);
nand UO_322 (O_322,N_9864,N_9886);
and UO_323 (O_323,N_9881,N_9866);
or UO_324 (O_324,N_9834,N_9916);
or UO_325 (O_325,N_9939,N_9963);
nand UO_326 (O_326,N_9947,N_9968);
nor UO_327 (O_327,N_9891,N_9969);
xor UO_328 (O_328,N_9805,N_9950);
or UO_329 (O_329,N_9934,N_9907);
or UO_330 (O_330,N_9865,N_9962);
nor UO_331 (O_331,N_9843,N_9979);
nor UO_332 (O_332,N_9824,N_9949);
nand UO_333 (O_333,N_9866,N_9938);
and UO_334 (O_334,N_9940,N_9921);
or UO_335 (O_335,N_9985,N_9936);
or UO_336 (O_336,N_9810,N_9964);
nor UO_337 (O_337,N_9991,N_9858);
nand UO_338 (O_338,N_9963,N_9937);
nand UO_339 (O_339,N_9937,N_9820);
xor UO_340 (O_340,N_9953,N_9971);
nor UO_341 (O_341,N_9804,N_9988);
nand UO_342 (O_342,N_9991,N_9919);
and UO_343 (O_343,N_9854,N_9933);
nor UO_344 (O_344,N_9914,N_9899);
xor UO_345 (O_345,N_9991,N_9882);
xor UO_346 (O_346,N_9850,N_9946);
or UO_347 (O_347,N_9859,N_9970);
and UO_348 (O_348,N_9999,N_9938);
or UO_349 (O_349,N_9973,N_9819);
xnor UO_350 (O_350,N_9835,N_9938);
nor UO_351 (O_351,N_9974,N_9823);
nand UO_352 (O_352,N_9844,N_9943);
xor UO_353 (O_353,N_9931,N_9843);
nand UO_354 (O_354,N_9915,N_9865);
and UO_355 (O_355,N_9986,N_9970);
or UO_356 (O_356,N_9961,N_9991);
and UO_357 (O_357,N_9881,N_9927);
and UO_358 (O_358,N_9894,N_9965);
or UO_359 (O_359,N_9934,N_9960);
or UO_360 (O_360,N_9800,N_9948);
and UO_361 (O_361,N_9906,N_9930);
xnor UO_362 (O_362,N_9936,N_9900);
nand UO_363 (O_363,N_9950,N_9980);
or UO_364 (O_364,N_9913,N_9835);
or UO_365 (O_365,N_9855,N_9990);
and UO_366 (O_366,N_9881,N_9802);
or UO_367 (O_367,N_9921,N_9897);
xnor UO_368 (O_368,N_9880,N_9992);
nand UO_369 (O_369,N_9974,N_9832);
or UO_370 (O_370,N_9840,N_9958);
or UO_371 (O_371,N_9927,N_9931);
nor UO_372 (O_372,N_9986,N_9857);
nor UO_373 (O_373,N_9919,N_9927);
or UO_374 (O_374,N_9979,N_9821);
xnor UO_375 (O_375,N_9848,N_9979);
or UO_376 (O_376,N_9885,N_9925);
xor UO_377 (O_377,N_9835,N_9815);
and UO_378 (O_378,N_9802,N_9860);
nor UO_379 (O_379,N_9847,N_9852);
or UO_380 (O_380,N_9968,N_9915);
nand UO_381 (O_381,N_9872,N_9931);
nand UO_382 (O_382,N_9953,N_9921);
and UO_383 (O_383,N_9952,N_9861);
xnor UO_384 (O_384,N_9824,N_9948);
xor UO_385 (O_385,N_9848,N_9964);
and UO_386 (O_386,N_9934,N_9971);
or UO_387 (O_387,N_9997,N_9866);
or UO_388 (O_388,N_9942,N_9849);
xor UO_389 (O_389,N_9887,N_9940);
nand UO_390 (O_390,N_9828,N_9947);
and UO_391 (O_391,N_9822,N_9980);
nor UO_392 (O_392,N_9963,N_9826);
nor UO_393 (O_393,N_9849,N_9870);
xor UO_394 (O_394,N_9952,N_9959);
xor UO_395 (O_395,N_9988,N_9959);
nor UO_396 (O_396,N_9833,N_9850);
or UO_397 (O_397,N_9973,N_9874);
nor UO_398 (O_398,N_9840,N_9811);
nand UO_399 (O_399,N_9921,N_9959);
xnor UO_400 (O_400,N_9976,N_9971);
nor UO_401 (O_401,N_9979,N_9825);
nor UO_402 (O_402,N_9915,N_9880);
nor UO_403 (O_403,N_9863,N_9925);
and UO_404 (O_404,N_9809,N_9863);
and UO_405 (O_405,N_9956,N_9990);
and UO_406 (O_406,N_9959,N_9847);
nand UO_407 (O_407,N_9997,N_9876);
nor UO_408 (O_408,N_9865,N_9964);
and UO_409 (O_409,N_9936,N_9812);
and UO_410 (O_410,N_9815,N_9931);
xor UO_411 (O_411,N_9980,N_9892);
or UO_412 (O_412,N_9945,N_9903);
or UO_413 (O_413,N_9855,N_9828);
xnor UO_414 (O_414,N_9998,N_9972);
or UO_415 (O_415,N_9870,N_9876);
or UO_416 (O_416,N_9944,N_9941);
nand UO_417 (O_417,N_9974,N_9939);
xor UO_418 (O_418,N_9997,N_9861);
or UO_419 (O_419,N_9984,N_9963);
nor UO_420 (O_420,N_9896,N_9877);
xnor UO_421 (O_421,N_9883,N_9854);
xnor UO_422 (O_422,N_9859,N_9895);
and UO_423 (O_423,N_9813,N_9942);
and UO_424 (O_424,N_9974,N_9969);
nand UO_425 (O_425,N_9839,N_9835);
nand UO_426 (O_426,N_9820,N_9934);
nand UO_427 (O_427,N_9897,N_9950);
nor UO_428 (O_428,N_9985,N_9801);
xor UO_429 (O_429,N_9964,N_9998);
nor UO_430 (O_430,N_9944,N_9854);
xor UO_431 (O_431,N_9877,N_9841);
nor UO_432 (O_432,N_9895,N_9991);
nor UO_433 (O_433,N_9970,N_9826);
xnor UO_434 (O_434,N_9948,N_9972);
or UO_435 (O_435,N_9945,N_9972);
nor UO_436 (O_436,N_9880,N_9968);
or UO_437 (O_437,N_9881,N_9803);
nand UO_438 (O_438,N_9937,N_9945);
or UO_439 (O_439,N_9984,N_9930);
and UO_440 (O_440,N_9930,N_9985);
xnor UO_441 (O_441,N_9903,N_9984);
nor UO_442 (O_442,N_9929,N_9978);
and UO_443 (O_443,N_9815,N_9864);
xnor UO_444 (O_444,N_9908,N_9987);
xnor UO_445 (O_445,N_9819,N_9840);
and UO_446 (O_446,N_9876,N_9847);
or UO_447 (O_447,N_9853,N_9994);
and UO_448 (O_448,N_9836,N_9899);
nor UO_449 (O_449,N_9968,N_9850);
nand UO_450 (O_450,N_9852,N_9997);
nand UO_451 (O_451,N_9907,N_9992);
nand UO_452 (O_452,N_9824,N_9940);
xor UO_453 (O_453,N_9898,N_9930);
xor UO_454 (O_454,N_9982,N_9836);
and UO_455 (O_455,N_9833,N_9828);
or UO_456 (O_456,N_9919,N_9984);
and UO_457 (O_457,N_9975,N_9874);
or UO_458 (O_458,N_9945,N_9969);
nand UO_459 (O_459,N_9973,N_9828);
and UO_460 (O_460,N_9881,N_9858);
nand UO_461 (O_461,N_9918,N_9974);
nand UO_462 (O_462,N_9980,N_9992);
nor UO_463 (O_463,N_9948,N_9909);
xor UO_464 (O_464,N_9827,N_9874);
nand UO_465 (O_465,N_9857,N_9987);
nand UO_466 (O_466,N_9825,N_9847);
or UO_467 (O_467,N_9979,N_9800);
xnor UO_468 (O_468,N_9802,N_9886);
or UO_469 (O_469,N_9803,N_9949);
and UO_470 (O_470,N_9997,N_9945);
nor UO_471 (O_471,N_9851,N_9977);
or UO_472 (O_472,N_9803,N_9915);
nor UO_473 (O_473,N_9972,N_9865);
and UO_474 (O_474,N_9990,N_9814);
nor UO_475 (O_475,N_9804,N_9993);
nand UO_476 (O_476,N_9983,N_9995);
or UO_477 (O_477,N_9955,N_9967);
nor UO_478 (O_478,N_9986,N_9987);
xnor UO_479 (O_479,N_9802,N_9925);
or UO_480 (O_480,N_9853,N_9866);
nor UO_481 (O_481,N_9823,N_9998);
xor UO_482 (O_482,N_9931,N_9869);
xnor UO_483 (O_483,N_9937,N_9995);
nor UO_484 (O_484,N_9801,N_9902);
nor UO_485 (O_485,N_9874,N_9932);
nand UO_486 (O_486,N_9906,N_9813);
or UO_487 (O_487,N_9974,N_9985);
and UO_488 (O_488,N_9925,N_9807);
nor UO_489 (O_489,N_9916,N_9982);
nor UO_490 (O_490,N_9894,N_9856);
nor UO_491 (O_491,N_9987,N_9920);
or UO_492 (O_492,N_9940,N_9955);
xor UO_493 (O_493,N_9936,N_9871);
xor UO_494 (O_494,N_9895,N_9809);
nand UO_495 (O_495,N_9818,N_9873);
nand UO_496 (O_496,N_9932,N_9845);
nor UO_497 (O_497,N_9863,N_9810);
nand UO_498 (O_498,N_9971,N_9927);
nor UO_499 (O_499,N_9956,N_9937);
xnor UO_500 (O_500,N_9930,N_9929);
nor UO_501 (O_501,N_9831,N_9907);
nand UO_502 (O_502,N_9803,N_9879);
xor UO_503 (O_503,N_9926,N_9876);
or UO_504 (O_504,N_9830,N_9970);
or UO_505 (O_505,N_9967,N_9954);
xnor UO_506 (O_506,N_9803,N_9931);
xor UO_507 (O_507,N_9890,N_9961);
or UO_508 (O_508,N_9968,N_9981);
or UO_509 (O_509,N_9891,N_9816);
nor UO_510 (O_510,N_9930,N_9895);
xnor UO_511 (O_511,N_9856,N_9827);
or UO_512 (O_512,N_9816,N_9930);
and UO_513 (O_513,N_9869,N_9924);
nand UO_514 (O_514,N_9950,N_9999);
and UO_515 (O_515,N_9828,N_9863);
or UO_516 (O_516,N_9944,N_9811);
or UO_517 (O_517,N_9836,N_9884);
or UO_518 (O_518,N_9970,N_9853);
nor UO_519 (O_519,N_9903,N_9979);
xnor UO_520 (O_520,N_9842,N_9900);
or UO_521 (O_521,N_9891,N_9863);
and UO_522 (O_522,N_9921,N_9819);
and UO_523 (O_523,N_9986,N_9817);
nor UO_524 (O_524,N_9843,N_9874);
xor UO_525 (O_525,N_9994,N_9973);
xnor UO_526 (O_526,N_9820,N_9933);
nand UO_527 (O_527,N_9946,N_9972);
or UO_528 (O_528,N_9865,N_9828);
and UO_529 (O_529,N_9926,N_9925);
nand UO_530 (O_530,N_9981,N_9840);
and UO_531 (O_531,N_9974,N_9861);
nand UO_532 (O_532,N_9972,N_9917);
or UO_533 (O_533,N_9805,N_9903);
nor UO_534 (O_534,N_9951,N_9828);
and UO_535 (O_535,N_9932,N_9981);
xnor UO_536 (O_536,N_9852,N_9875);
or UO_537 (O_537,N_9802,N_9975);
xor UO_538 (O_538,N_9867,N_9983);
or UO_539 (O_539,N_9940,N_9857);
nor UO_540 (O_540,N_9953,N_9968);
nor UO_541 (O_541,N_9901,N_9850);
nand UO_542 (O_542,N_9942,N_9878);
xnor UO_543 (O_543,N_9917,N_9925);
xor UO_544 (O_544,N_9970,N_9981);
nand UO_545 (O_545,N_9969,N_9800);
xnor UO_546 (O_546,N_9910,N_9996);
or UO_547 (O_547,N_9835,N_9933);
and UO_548 (O_548,N_9951,N_9845);
nand UO_549 (O_549,N_9842,N_9931);
nand UO_550 (O_550,N_9917,N_9970);
xor UO_551 (O_551,N_9866,N_9827);
nand UO_552 (O_552,N_9950,N_9844);
nand UO_553 (O_553,N_9820,N_9930);
and UO_554 (O_554,N_9997,N_9993);
nand UO_555 (O_555,N_9992,N_9892);
xnor UO_556 (O_556,N_9915,N_9942);
xnor UO_557 (O_557,N_9983,N_9869);
or UO_558 (O_558,N_9952,N_9819);
or UO_559 (O_559,N_9995,N_9969);
and UO_560 (O_560,N_9890,N_9840);
or UO_561 (O_561,N_9915,N_9931);
and UO_562 (O_562,N_9815,N_9808);
nand UO_563 (O_563,N_9973,N_9856);
xnor UO_564 (O_564,N_9880,N_9886);
and UO_565 (O_565,N_9943,N_9988);
or UO_566 (O_566,N_9992,N_9935);
or UO_567 (O_567,N_9906,N_9880);
or UO_568 (O_568,N_9945,N_9807);
nor UO_569 (O_569,N_9957,N_9925);
xor UO_570 (O_570,N_9923,N_9952);
nor UO_571 (O_571,N_9957,N_9997);
or UO_572 (O_572,N_9826,N_9897);
or UO_573 (O_573,N_9807,N_9938);
xnor UO_574 (O_574,N_9844,N_9907);
or UO_575 (O_575,N_9922,N_9938);
nand UO_576 (O_576,N_9846,N_9946);
xnor UO_577 (O_577,N_9963,N_9856);
and UO_578 (O_578,N_9957,N_9872);
and UO_579 (O_579,N_9894,N_9982);
xor UO_580 (O_580,N_9889,N_9870);
and UO_581 (O_581,N_9967,N_9916);
and UO_582 (O_582,N_9946,N_9801);
or UO_583 (O_583,N_9964,N_9824);
and UO_584 (O_584,N_9912,N_9801);
nor UO_585 (O_585,N_9995,N_9968);
nand UO_586 (O_586,N_9814,N_9882);
nor UO_587 (O_587,N_9965,N_9846);
and UO_588 (O_588,N_9991,N_9930);
and UO_589 (O_589,N_9940,N_9916);
nand UO_590 (O_590,N_9977,N_9825);
nand UO_591 (O_591,N_9839,N_9902);
xnor UO_592 (O_592,N_9853,N_9877);
and UO_593 (O_593,N_9980,N_9972);
and UO_594 (O_594,N_9872,N_9962);
nor UO_595 (O_595,N_9867,N_9961);
nand UO_596 (O_596,N_9848,N_9908);
xnor UO_597 (O_597,N_9973,N_9857);
xor UO_598 (O_598,N_9930,N_9828);
or UO_599 (O_599,N_9944,N_9974);
nor UO_600 (O_600,N_9818,N_9874);
nand UO_601 (O_601,N_9857,N_9983);
xnor UO_602 (O_602,N_9865,N_9868);
nor UO_603 (O_603,N_9981,N_9965);
and UO_604 (O_604,N_9956,N_9837);
nand UO_605 (O_605,N_9944,N_9920);
nand UO_606 (O_606,N_9863,N_9962);
and UO_607 (O_607,N_9868,N_9919);
nor UO_608 (O_608,N_9839,N_9881);
nor UO_609 (O_609,N_9962,N_9895);
xnor UO_610 (O_610,N_9931,N_9837);
nand UO_611 (O_611,N_9907,N_9854);
or UO_612 (O_612,N_9831,N_9975);
nand UO_613 (O_613,N_9873,N_9922);
and UO_614 (O_614,N_9992,N_9846);
xor UO_615 (O_615,N_9867,N_9875);
and UO_616 (O_616,N_9818,N_9961);
nand UO_617 (O_617,N_9802,N_9853);
nor UO_618 (O_618,N_9864,N_9862);
or UO_619 (O_619,N_9958,N_9928);
xnor UO_620 (O_620,N_9907,N_9840);
nand UO_621 (O_621,N_9964,N_9897);
and UO_622 (O_622,N_9917,N_9824);
nor UO_623 (O_623,N_9866,N_9998);
or UO_624 (O_624,N_9904,N_9875);
nor UO_625 (O_625,N_9963,N_9995);
and UO_626 (O_626,N_9889,N_9931);
nand UO_627 (O_627,N_9836,N_9905);
nand UO_628 (O_628,N_9881,N_9816);
nand UO_629 (O_629,N_9824,N_9933);
or UO_630 (O_630,N_9950,N_9910);
xor UO_631 (O_631,N_9931,N_9813);
nor UO_632 (O_632,N_9862,N_9903);
nand UO_633 (O_633,N_9878,N_9804);
and UO_634 (O_634,N_9919,N_9856);
and UO_635 (O_635,N_9879,N_9805);
and UO_636 (O_636,N_9972,N_9940);
or UO_637 (O_637,N_9853,N_9940);
or UO_638 (O_638,N_9853,N_9848);
xor UO_639 (O_639,N_9919,N_9943);
xnor UO_640 (O_640,N_9935,N_9954);
or UO_641 (O_641,N_9890,N_9923);
or UO_642 (O_642,N_9833,N_9918);
or UO_643 (O_643,N_9923,N_9802);
and UO_644 (O_644,N_9873,N_9905);
or UO_645 (O_645,N_9910,N_9933);
and UO_646 (O_646,N_9950,N_9893);
nand UO_647 (O_647,N_9988,N_9969);
or UO_648 (O_648,N_9968,N_9874);
xnor UO_649 (O_649,N_9973,N_9938);
and UO_650 (O_650,N_9821,N_9947);
and UO_651 (O_651,N_9861,N_9867);
and UO_652 (O_652,N_9899,N_9864);
or UO_653 (O_653,N_9855,N_9933);
xor UO_654 (O_654,N_9851,N_9937);
nor UO_655 (O_655,N_9933,N_9838);
nor UO_656 (O_656,N_9971,N_9892);
nand UO_657 (O_657,N_9920,N_9818);
and UO_658 (O_658,N_9995,N_9827);
and UO_659 (O_659,N_9847,N_9930);
and UO_660 (O_660,N_9976,N_9993);
and UO_661 (O_661,N_9998,N_9966);
nand UO_662 (O_662,N_9920,N_9832);
and UO_663 (O_663,N_9818,N_9810);
nand UO_664 (O_664,N_9838,N_9939);
and UO_665 (O_665,N_9817,N_9997);
nand UO_666 (O_666,N_9870,N_9810);
nand UO_667 (O_667,N_9968,N_9843);
nor UO_668 (O_668,N_9939,N_9928);
or UO_669 (O_669,N_9862,N_9863);
nand UO_670 (O_670,N_9958,N_9976);
nand UO_671 (O_671,N_9918,N_9931);
or UO_672 (O_672,N_9969,N_9966);
nand UO_673 (O_673,N_9957,N_9908);
and UO_674 (O_674,N_9810,N_9893);
xnor UO_675 (O_675,N_9917,N_9941);
or UO_676 (O_676,N_9848,N_9931);
or UO_677 (O_677,N_9860,N_9960);
and UO_678 (O_678,N_9914,N_9942);
or UO_679 (O_679,N_9830,N_9992);
or UO_680 (O_680,N_9921,N_9845);
xnor UO_681 (O_681,N_9835,N_9843);
nor UO_682 (O_682,N_9839,N_9981);
and UO_683 (O_683,N_9878,N_9880);
and UO_684 (O_684,N_9872,N_9843);
or UO_685 (O_685,N_9884,N_9876);
xnor UO_686 (O_686,N_9857,N_9897);
xor UO_687 (O_687,N_9916,N_9856);
or UO_688 (O_688,N_9950,N_9871);
xor UO_689 (O_689,N_9827,N_9901);
nor UO_690 (O_690,N_9986,N_9977);
or UO_691 (O_691,N_9921,N_9808);
and UO_692 (O_692,N_9973,N_9858);
or UO_693 (O_693,N_9969,N_9819);
nor UO_694 (O_694,N_9984,N_9937);
xnor UO_695 (O_695,N_9907,N_9927);
xnor UO_696 (O_696,N_9882,N_9936);
nor UO_697 (O_697,N_9920,N_9874);
or UO_698 (O_698,N_9850,N_9845);
and UO_699 (O_699,N_9948,N_9828);
nor UO_700 (O_700,N_9942,N_9852);
xor UO_701 (O_701,N_9897,N_9930);
xnor UO_702 (O_702,N_9987,N_9879);
nand UO_703 (O_703,N_9801,N_9998);
and UO_704 (O_704,N_9849,N_9824);
and UO_705 (O_705,N_9805,N_9810);
and UO_706 (O_706,N_9954,N_9911);
or UO_707 (O_707,N_9800,N_9883);
and UO_708 (O_708,N_9931,N_9916);
nor UO_709 (O_709,N_9817,N_9879);
or UO_710 (O_710,N_9996,N_9947);
nor UO_711 (O_711,N_9988,N_9887);
nor UO_712 (O_712,N_9985,N_9945);
xnor UO_713 (O_713,N_9902,N_9905);
xnor UO_714 (O_714,N_9812,N_9994);
or UO_715 (O_715,N_9964,N_9880);
nor UO_716 (O_716,N_9844,N_9891);
and UO_717 (O_717,N_9937,N_9807);
xor UO_718 (O_718,N_9948,N_9919);
nor UO_719 (O_719,N_9932,N_9953);
nor UO_720 (O_720,N_9995,N_9976);
xnor UO_721 (O_721,N_9844,N_9824);
xor UO_722 (O_722,N_9866,N_9963);
nand UO_723 (O_723,N_9877,N_9978);
nor UO_724 (O_724,N_9879,N_9829);
or UO_725 (O_725,N_9836,N_9949);
nand UO_726 (O_726,N_9802,N_9951);
nor UO_727 (O_727,N_9892,N_9996);
and UO_728 (O_728,N_9973,N_9899);
nor UO_729 (O_729,N_9958,N_9925);
and UO_730 (O_730,N_9843,N_9953);
nand UO_731 (O_731,N_9868,N_9864);
nand UO_732 (O_732,N_9904,N_9901);
nand UO_733 (O_733,N_9911,N_9866);
nor UO_734 (O_734,N_9886,N_9938);
and UO_735 (O_735,N_9955,N_9924);
or UO_736 (O_736,N_9918,N_9990);
or UO_737 (O_737,N_9841,N_9969);
or UO_738 (O_738,N_9966,N_9906);
nand UO_739 (O_739,N_9976,N_9910);
nand UO_740 (O_740,N_9826,N_9873);
xor UO_741 (O_741,N_9990,N_9934);
or UO_742 (O_742,N_9929,N_9806);
or UO_743 (O_743,N_9858,N_9876);
nand UO_744 (O_744,N_9801,N_9863);
xor UO_745 (O_745,N_9856,N_9934);
or UO_746 (O_746,N_9905,N_9884);
nor UO_747 (O_747,N_9930,N_9899);
nand UO_748 (O_748,N_9897,N_9851);
nor UO_749 (O_749,N_9805,N_9944);
nand UO_750 (O_750,N_9835,N_9811);
xnor UO_751 (O_751,N_9986,N_9877);
or UO_752 (O_752,N_9961,N_9899);
xor UO_753 (O_753,N_9946,N_9903);
nand UO_754 (O_754,N_9954,N_9923);
or UO_755 (O_755,N_9850,N_9998);
nand UO_756 (O_756,N_9899,N_9934);
xnor UO_757 (O_757,N_9980,N_9841);
xnor UO_758 (O_758,N_9862,N_9933);
and UO_759 (O_759,N_9873,N_9942);
nand UO_760 (O_760,N_9830,N_9856);
xnor UO_761 (O_761,N_9858,N_9907);
or UO_762 (O_762,N_9929,N_9979);
xnor UO_763 (O_763,N_9960,N_9970);
or UO_764 (O_764,N_9810,N_9812);
xor UO_765 (O_765,N_9848,N_9821);
nand UO_766 (O_766,N_9827,N_9913);
and UO_767 (O_767,N_9837,N_9909);
xor UO_768 (O_768,N_9997,N_9801);
and UO_769 (O_769,N_9938,N_9971);
nor UO_770 (O_770,N_9942,N_9897);
and UO_771 (O_771,N_9886,N_9898);
nand UO_772 (O_772,N_9969,N_9839);
nor UO_773 (O_773,N_9872,N_9927);
nand UO_774 (O_774,N_9896,N_9995);
or UO_775 (O_775,N_9883,N_9853);
or UO_776 (O_776,N_9945,N_9896);
or UO_777 (O_777,N_9846,N_9831);
nand UO_778 (O_778,N_9976,N_9826);
nor UO_779 (O_779,N_9992,N_9961);
nor UO_780 (O_780,N_9821,N_9950);
or UO_781 (O_781,N_9932,N_9826);
or UO_782 (O_782,N_9801,N_9921);
and UO_783 (O_783,N_9958,N_9859);
nand UO_784 (O_784,N_9987,N_9833);
xnor UO_785 (O_785,N_9982,N_9914);
nand UO_786 (O_786,N_9996,N_9955);
nand UO_787 (O_787,N_9927,N_9820);
nand UO_788 (O_788,N_9869,N_9881);
or UO_789 (O_789,N_9856,N_9964);
xnor UO_790 (O_790,N_9885,N_9873);
nor UO_791 (O_791,N_9873,N_9956);
nand UO_792 (O_792,N_9965,N_9967);
nand UO_793 (O_793,N_9970,N_9962);
xnor UO_794 (O_794,N_9995,N_9883);
or UO_795 (O_795,N_9816,N_9986);
and UO_796 (O_796,N_9881,N_9876);
and UO_797 (O_797,N_9883,N_9909);
nand UO_798 (O_798,N_9825,N_9856);
and UO_799 (O_799,N_9814,N_9815);
nor UO_800 (O_800,N_9988,N_9846);
xor UO_801 (O_801,N_9931,N_9989);
xor UO_802 (O_802,N_9939,N_9880);
or UO_803 (O_803,N_9879,N_9990);
or UO_804 (O_804,N_9828,N_9913);
or UO_805 (O_805,N_9959,N_9905);
and UO_806 (O_806,N_9819,N_9977);
xor UO_807 (O_807,N_9933,N_9967);
and UO_808 (O_808,N_9862,N_9909);
nor UO_809 (O_809,N_9897,N_9820);
nand UO_810 (O_810,N_9870,N_9815);
nand UO_811 (O_811,N_9844,N_9999);
and UO_812 (O_812,N_9829,N_9930);
or UO_813 (O_813,N_9855,N_9967);
nand UO_814 (O_814,N_9877,N_9882);
or UO_815 (O_815,N_9998,N_9802);
nor UO_816 (O_816,N_9832,N_9938);
nor UO_817 (O_817,N_9891,N_9843);
nand UO_818 (O_818,N_9902,N_9939);
nand UO_819 (O_819,N_9913,N_9907);
or UO_820 (O_820,N_9865,N_9980);
or UO_821 (O_821,N_9840,N_9999);
nor UO_822 (O_822,N_9830,N_9819);
xor UO_823 (O_823,N_9989,N_9983);
nor UO_824 (O_824,N_9859,N_9802);
and UO_825 (O_825,N_9828,N_9950);
and UO_826 (O_826,N_9810,N_9915);
or UO_827 (O_827,N_9894,N_9899);
and UO_828 (O_828,N_9918,N_9863);
nor UO_829 (O_829,N_9959,N_9946);
nand UO_830 (O_830,N_9833,N_9827);
and UO_831 (O_831,N_9976,N_9848);
and UO_832 (O_832,N_9823,N_9887);
and UO_833 (O_833,N_9823,N_9981);
nand UO_834 (O_834,N_9953,N_9858);
xnor UO_835 (O_835,N_9815,N_9990);
or UO_836 (O_836,N_9996,N_9801);
or UO_837 (O_837,N_9965,N_9884);
or UO_838 (O_838,N_9997,N_9987);
xnor UO_839 (O_839,N_9923,N_9906);
xnor UO_840 (O_840,N_9826,N_9823);
nor UO_841 (O_841,N_9976,N_9843);
xor UO_842 (O_842,N_9890,N_9838);
nor UO_843 (O_843,N_9930,N_9996);
nor UO_844 (O_844,N_9857,N_9859);
and UO_845 (O_845,N_9833,N_9997);
xor UO_846 (O_846,N_9872,N_9915);
or UO_847 (O_847,N_9807,N_9826);
and UO_848 (O_848,N_9982,N_9954);
or UO_849 (O_849,N_9908,N_9868);
nor UO_850 (O_850,N_9952,N_9979);
nand UO_851 (O_851,N_9852,N_9977);
nand UO_852 (O_852,N_9910,N_9832);
nor UO_853 (O_853,N_9835,N_9907);
xnor UO_854 (O_854,N_9816,N_9800);
and UO_855 (O_855,N_9972,N_9939);
or UO_856 (O_856,N_9894,N_9904);
xnor UO_857 (O_857,N_9882,N_9892);
nor UO_858 (O_858,N_9931,N_9926);
and UO_859 (O_859,N_9959,N_9842);
nor UO_860 (O_860,N_9866,N_9849);
nor UO_861 (O_861,N_9964,N_9960);
or UO_862 (O_862,N_9996,N_9901);
or UO_863 (O_863,N_9914,N_9951);
or UO_864 (O_864,N_9979,N_9869);
nand UO_865 (O_865,N_9818,N_9984);
and UO_866 (O_866,N_9816,N_9804);
and UO_867 (O_867,N_9922,N_9821);
nor UO_868 (O_868,N_9838,N_9857);
xnor UO_869 (O_869,N_9943,N_9991);
nand UO_870 (O_870,N_9807,N_9998);
or UO_871 (O_871,N_9890,N_9906);
nor UO_872 (O_872,N_9971,N_9942);
nand UO_873 (O_873,N_9875,N_9941);
xnor UO_874 (O_874,N_9951,N_9997);
xor UO_875 (O_875,N_9862,N_9854);
xnor UO_876 (O_876,N_9823,N_9814);
or UO_877 (O_877,N_9866,N_9994);
nand UO_878 (O_878,N_9856,N_9956);
nor UO_879 (O_879,N_9976,N_9895);
and UO_880 (O_880,N_9931,N_9974);
xor UO_881 (O_881,N_9920,N_9811);
nand UO_882 (O_882,N_9918,N_9904);
xnor UO_883 (O_883,N_9994,N_9880);
and UO_884 (O_884,N_9813,N_9804);
and UO_885 (O_885,N_9911,N_9830);
and UO_886 (O_886,N_9934,N_9822);
and UO_887 (O_887,N_9888,N_9921);
or UO_888 (O_888,N_9962,N_9923);
nor UO_889 (O_889,N_9953,N_9830);
nand UO_890 (O_890,N_9935,N_9803);
or UO_891 (O_891,N_9812,N_9907);
nor UO_892 (O_892,N_9866,N_9996);
nor UO_893 (O_893,N_9952,N_9804);
xnor UO_894 (O_894,N_9935,N_9871);
xnor UO_895 (O_895,N_9879,N_9906);
xor UO_896 (O_896,N_9864,N_9918);
xor UO_897 (O_897,N_9983,N_9815);
xor UO_898 (O_898,N_9977,N_9937);
nor UO_899 (O_899,N_9855,N_9899);
nor UO_900 (O_900,N_9986,N_9859);
nand UO_901 (O_901,N_9851,N_9969);
nand UO_902 (O_902,N_9862,N_9843);
nor UO_903 (O_903,N_9828,N_9956);
nand UO_904 (O_904,N_9814,N_9837);
and UO_905 (O_905,N_9936,N_9887);
and UO_906 (O_906,N_9880,N_9829);
or UO_907 (O_907,N_9976,N_9886);
or UO_908 (O_908,N_9817,N_9962);
and UO_909 (O_909,N_9855,N_9847);
and UO_910 (O_910,N_9969,N_9809);
xor UO_911 (O_911,N_9836,N_9987);
nor UO_912 (O_912,N_9945,N_9933);
xor UO_913 (O_913,N_9843,N_9971);
xnor UO_914 (O_914,N_9990,N_9884);
or UO_915 (O_915,N_9859,N_9973);
and UO_916 (O_916,N_9965,N_9832);
xor UO_917 (O_917,N_9869,N_9990);
or UO_918 (O_918,N_9895,N_9810);
nand UO_919 (O_919,N_9867,N_9920);
and UO_920 (O_920,N_9924,N_9997);
nor UO_921 (O_921,N_9809,N_9913);
nand UO_922 (O_922,N_9971,N_9929);
or UO_923 (O_923,N_9984,N_9898);
or UO_924 (O_924,N_9888,N_9903);
and UO_925 (O_925,N_9800,N_9951);
or UO_926 (O_926,N_9880,N_9815);
xor UO_927 (O_927,N_9881,N_9979);
nand UO_928 (O_928,N_9899,N_9963);
nor UO_929 (O_929,N_9924,N_9952);
xnor UO_930 (O_930,N_9962,N_9990);
or UO_931 (O_931,N_9920,N_9995);
and UO_932 (O_932,N_9995,N_9935);
or UO_933 (O_933,N_9901,N_9859);
or UO_934 (O_934,N_9986,N_9864);
xnor UO_935 (O_935,N_9813,N_9811);
nor UO_936 (O_936,N_9881,N_9859);
xnor UO_937 (O_937,N_9989,N_9814);
nor UO_938 (O_938,N_9904,N_9946);
nand UO_939 (O_939,N_9874,N_9896);
and UO_940 (O_940,N_9859,N_9843);
or UO_941 (O_941,N_9914,N_9895);
xor UO_942 (O_942,N_9816,N_9944);
nand UO_943 (O_943,N_9992,N_9816);
xor UO_944 (O_944,N_9808,N_9913);
or UO_945 (O_945,N_9858,N_9945);
and UO_946 (O_946,N_9956,N_9955);
and UO_947 (O_947,N_9817,N_9915);
or UO_948 (O_948,N_9933,N_9897);
and UO_949 (O_949,N_9987,N_9916);
and UO_950 (O_950,N_9813,N_9998);
nand UO_951 (O_951,N_9939,N_9840);
xor UO_952 (O_952,N_9968,N_9914);
nand UO_953 (O_953,N_9834,N_9954);
nor UO_954 (O_954,N_9992,N_9836);
and UO_955 (O_955,N_9897,N_9922);
nand UO_956 (O_956,N_9901,N_9865);
or UO_957 (O_957,N_9869,N_9843);
and UO_958 (O_958,N_9811,N_9969);
or UO_959 (O_959,N_9903,N_9877);
or UO_960 (O_960,N_9963,N_9891);
or UO_961 (O_961,N_9893,N_9813);
or UO_962 (O_962,N_9978,N_9837);
xor UO_963 (O_963,N_9886,N_9832);
xnor UO_964 (O_964,N_9860,N_9833);
nand UO_965 (O_965,N_9887,N_9882);
xnor UO_966 (O_966,N_9967,N_9924);
or UO_967 (O_967,N_9914,N_9888);
nor UO_968 (O_968,N_9980,N_9960);
nor UO_969 (O_969,N_9932,N_9999);
nand UO_970 (O_970,N_9993,N_9943);
xor UO_971 (O_971,N_9811,N_9980);
and UO_972 (O_972,N_9830,N_9808);
nand UO_973 (O_973,N_9894,N_9917);
nand UO_974 (O_974,N_9901,N_9813);
nor UO_975 (O_975,N_9881,N_9875);
and UO_976 (O_976,N_9860,N_9857);
nor UO_977 (O_977,N_9890,N_9857);
nor UO_978 (O_978,N_9878,N_9984);
nand UO_979 (O_979,N_9836,N_9916);
or UO_980 (O_980,N_9957,N_9893);
nand UO_981 (O_981,N_9870,N_9919);
or UO_982 (O_982,N_9825,N_9958);
nor UO_983 (O_983,N_9985,N_9948);
or UO_984 (O_984,N_9971,N_9956);
xnor UO_985 (O_985,N_9977,N_9803);
nand UO_986 (O_986,N_9907,N_9800);
or UO_987 (O_987,N_9821,N_9901);
nor UO_988 (O_988,N_9926,N_9889);
xor UO_989 (O_989,N_9828,N_9912);
nor UO_990 (O_990,N_9832,N_9905);
nor UO_991 (O_991,N_9867,N_9840);
xor UO_992 (O_992,N_9984,N_9978);
nand UO_993 (O_993,N_9977,N_9933);
xor UO_994 (O_994,N_9898,N_9889);
xor UO_995 (O_995,N_9976,N_9902);
nand UO_996 (O_996,N_9894,N_9921);
and UO_997 (O_997,N_9828,N_9878);
xnor UO_998 (O_998,N_9891,N_9881);
nor UO_999 (O_999,N_9920,N_9810);
nand UO_1000 (O_1000,N_9973,N_9941);
or UO_1001 (O_1001,N_9838,N_9846);
nor UO_1002 (O_1002,N_9803,N_9832);
or UO_1003 (O_1003,N_9836,N_9975);
nor UO_1004 (O_1004,N_9828,N_9889);
nor UO_1005 (O_1005,N_9998,N_9806);
xnor UO_1006 (O_1006,N_9916,N_9958);
or UO_1007 (O_1007,N_9810,N_9883);
nand UO_1008 (O_1008,N_9967,N_9966);
and UO_1009 (O_1009,N_9809,N_9810);
xnor UO_1010 (O_1010,N_9817,N_9940);
and UO_1011 (O_1011,N_9976,N_9917);
nor UO_1012 (O_1012,N_9843,N_9903);
nor UO_1013 (O_1013,N_9855,N_9821);
nor UO_1014 (O_1014,N_9819,N_9862);
nor UO_1015 (O_1015,N_9989,N_9966);
or UO_1016 (O_1016,N_9993,N_9844);
and UO_1017 (O_1017,N_9992,N_9895);
xnor UO_1018 (O_1018,N_9959,N_9849);
or UO_1019 (O_1019,N_9985,N_9915);
or UO_1020 (O_1020,N_9839,N_9834);
nand UO_1021 (O_1021,N_9946,N_9991);
or UO_1022 (O_1022,N_9841,N_9961);
xnor UO_1023 (O_1023,N_9956,N_9846);
nand UO_1024 (O_1024,N_9860,N_9983);
or UO_1025 (O_1025,N_9897,N_9830);
and UO_1026 (O_1026,N_9813,N_9899);
xor UO_1027 (O_1027,N_9921,N_9810);
nand UO_1028 (O_1028,N_9894,N_9835);
xor UO_1029 (O_1029,N_9975,N_9961);
nand UO_1030 (O_1030,N_9949,N_9964);
or UO_1031 (O_1031,N_9924,N_9979);
nor UO_1032 (O_1032,N_9852,N_9909);
xor UO_1033 (O_1033,N_9827,N_9889);
or UO_1034 (O_1034,N_9805,N_9947);
nand UO_1035 (O_1035,N_9899,N_9888);
nand UO_1036 (O_1036,N_9957,N_9856);
nand UO_1037 (O_1037,N_9828,N_9914);
nor UO_1038 (O_1038,N_9850,N_9912);
nand UO_1039 (O_1039,N_9939,N_9925);
or UO_1040 (O_1040,N_9999,N_9814);
xor UO_1041 (O_1041,N_9929,N_9840);
and UO_1042 (O_1042,N_9805,N_9983);
nor UO_1043 (O_1043,N_9900,N_9895);
nand UO_1044 (O_1044,N_9893,N_9892);
nand UO_1045 (O_1045,N_9877,N_9993);
and UO_1046 (O_1046,N_9832,N_9901);
and UO_1047 (O_1047,N_9812,N_9899);
nand UO_1048 (O_1048,N_9945,N_9914);
xor UO_1049 (O_1049,N_9965,N_9956);
or UO_1050 (O_1050,N_9918,N_9871);
or UO_1051 (O_1051,N_9910,N_9959);
xnor UO_1052 (O_1052,N_9954,N_9909);
nor UO_1053 (O_1053,N_9847,N_9845);
and UO_1054 (O_1054,N_9976,N_9943);
nand UO_1055 (O_1055,N_9879,N_9910);
nand UO_1056 (O_1056,N_9847,N_9887);
nor UO_1057 (O_1057,N_9803,N_9953);
and UO_1058 (O_1058,N_9906,N_9973);
or UO_1059 (O_1059,N_9926,N_9909);
nand UO_1060 (O_1060,N_9972,N_9988);
nor UO_1061 (O_1061,N_9954,N_9916);
xor UO_1062 (O_1062,N_9824,N_9830);
nand UO_1063 (O_1063,N_9911,N_9806);
or UO_1064 (O_1064,N_9886,N_9896);
nand UO_1065 (O_1065,N_9912,N_9938);
nand UO_1066 (O_1066,N_9854,N_9849);
and UO_1067 (O_1067,N_9998,N_9980);
xnor UO_1068 (O_1068,N_9887,N_9838);
xnor UO_1069 (O_1069,N_9851,N_9978);
or UO_1070 (O_1070,N_9945,N_9921);
nor UO_1071 (O_1071,N_9839,N_9904);
nor UO_1072 (O_1072,N_9994,N_9954);
nand UO_1073 (O_1073,N_9887,N_9956);
nor UO_1074 (O_1074,N_9984,N_9924);
or UO_1075 (O_1075,N_9901,N_9861);
xnor UO_1076 (O_1076,N_9956,N_9917);
nor UO_1077 (O_1077,N_9991,N_9988);
nor UO_1078 (O_1078,N_9835,N_9832);
nor UO_1079 (O_1079,N_9991,N_9819);
nand UO_1080 (O_1080,N_9802,N_9972);
nand UO_1081 (O_1081,N_9800,N_9930);
xnor UO_1082 (O_1082,N_9915,N_9800);
nand UO_1083 (O_1083,N_9934,N_9985);
or UO_1084 (O_1084,N_9959,N_9977);
xnor UO_1085 (O_1085,N_9978,N_9915);
nand UO_1086 (O_1086,N_9820,N_9904);
and UO_1087 (O_1087,N_9953,N_9951);
nor UO_1088 (O_1088,N_9921,N_9830);
xnor UO_1089 (O_1089,N_9985,N_9995);
and UO_1090 (O_1090,N_9901,N_9938);
xor UO_1091 (O_1091,N_9926,N_9901);
and UO_1092 (O_1092,N_9865,N_9934);
or UO_1093 (O_1093,N_9964,N_9807);
nand UO_1094 (O_1094,N_9936,N_9939);
xor UO_1095 (O_1095,N_9991,N_9832);
nor UO_1096 (O_1096,N_9955,N_9957);
xor UO_1097 (O_1097,N_9800,N_9926);
nor UO_1098 (O_1098,N_9887,N_9839);
or UO_1099 (O_1099,N_9928,N_9994);
and UO_1100 (O_1100,N_9912,N_9859);
nand UO_1101 (O_1101,N_9967,N_9895);
xnor UO_1102 (O_1102,N_9868,N_9840);
or UO_1103 (O_1103,N_9895,N_9922);
or UO_1104 (O_1104,N_9875,N_9887);
nor UO_1105 (O_1105,N_9921,N_9829);
and UO_1106 (O_1106,N_9999,N_9960);
and UO_1107 (O_1107,N_9964,N_9922);
xnor UO_1108 (O_1108,N_9848,N_9973);
nor UO_1109 (O_1109,N_9833,N_9934);
or UO_1110 (O_1110,N_9889,N_9820);
xnor UO_1111 (O_1111,N_9850,N_9811);
and UO_1112 (O_1112,N_9843,N_9865);
nor UO_1113 (O_1113,N_9883,N_9863);
nand UO_1114 (O_1114,N_9827,N_9948);
nor UO_1115 (O_1115,N_9941,N_9869);
xor UO_1116 (O_1116,N_9813,N_9847);
nand UO_1117 (O_1117,N_9916,N_9846);
or UO_1118 (O_1118,N_9952,N_9888);
or UO_1119 (O_1119,N_9821,N_9991);
nor UO_1120 (O_1120,N_9822,N_9815);
xnor UO_1121 (O_1121,N_9993,N_9824);
nand UO_1122 (O_1122,N_9908,N_9843);
or UO_1123 (O_1123,N_9894,N_9833);
or UO_1124 (O_1124,N_9924,N_9940);
nand UO_1125 (O_1125,N_9990,N_9927);
xor UO_1126 (O_1126,N_9974,N_9815);
or UO_1127 (O_1127,N_9847,N_9895);
nor UO_1128 (O_1128,N_9954,N_9850);
or UO_1129 (O_1129,N_9849,N_9955);
xnor UO_1130 (O_1130,N_9962,N_9878);
or UO_1131 (O_1131,N_9840,N_9984);
and UO_1132 (O_1132,N_9813,N_9937);
nor UO_1133 (O_1133,N_9964,N_9886);
and UO_1134 (O_1134,N_9852,N_9851);
nand UO_1135 (O_1135,N_9916,N_9988);
nand UO_1136 (O_1136,N_9830,N_9983);
xor UO_1137 (O_1137,N_9852,N_9886);
nand UO_1138 (O_1138,N_9893,N_9802);
xor UO_1139 (O_1139,N_9867,N_9811);
and UO_1140 (O_1140,N_9949,N_9892);
or UO_1141 (O_1141,N_9934,N_9973);
and UO_1142 (O_1142,N_9916,N_9919);
nor UO_1143 (O_1143,N_9909,N_9939);
nor UO_1144 (O_1144,N_9973,N_9945);
nand UO_1145 (O_1145,N_9936,N_9923);
nor UO_1146 (O_1146,N_9832,N_9900);
nor UO_1147 (O_1147,N_9921,N_9999);
or UO_1148 (O_1148,N_9860,N_9824);
xnor UO_1149 (O_1149,N_9867,N_9805);
or UO_1150 (O_1150,N_9921,N_9929);
nand UO_1151 (O_1151,N_9994,N_9989);
and UO_1152 (O_1152,N_9831,N_9868);
xor UO_1153 (O_1153,N_9875,N_9890);
nand UO_1154 (O_1154,N_9968,N_9927);
xor UO_1155 (O_1155,N_9867,N_9869);
and UO_1156 (O_1156,N_9837,N_9822);
nand UO_1157 (O_1157,N_9825,N_9861);
and UO_1158 (O_1158,N_9834,N_9851);
nand UO_1159 (O_1159,N_9975,N_9820);
nor UO_1160 (O_1160,N_9982,N_9882);
nand UO_1161 (O_1161,N_9803,N_9913);
xnor UO_1162 (O_1162,N_9990,N_9886);
nand UO_1163 (O_1163,N_9884,N_9831);
nor UO_1164 (O_1164,N_9967,N_9825);
or UO_1165 (O_1165,N_9976,N_9876);
xnor UO_1166 (O_1166,N_9891,N_9830);
nor UO_1167 (O_1167,N_9888,N_9900);
and UO_1168 (O_1168,N_9940,N_9966);
or UO_1169 (O_1169,N_9992,N_9904);
nor UO_1170 (O_1170,N_9888,N_9844);
or UO_1171 (O_1171,N_9898,N_9916);
xor UO_1172 (O_1172,N_9899,N_9816);
nand UO_1173 (O_1173,N_9909,N_9876);
nand UO_1174 (O_1174,N_9964,N_9854);
and UO_1175 (O_1175,N_9996,N_9917);
nor UO_1176 (O_1176,N_9909,N_9990);
xnor UO_1177 (O_1177,N_9921,N_9887);
nand UO_1178 (O_1178,N_9970,N_9831);
and UO_1179 (O_1179,N_9927,N_9856);
and UO_1180 (O_1180,N_9994,N_9851);
or UO_1181 (O_1181,N_9941,N_9832);
or UO_1182 (O_1182,N_9801,N_9862);
nand UO_1183 (O_1183,N_9964,N_9941);
nor UO_1184 (O_1184,N_9947,N_9880);
xnor UO_1185 (O_1185,N_9822,N_9894);
xnor UO_1186 (O_1186,N_9888,N_9941);
xor UO_1187 (O_1187,N_9839,N_9931);
nand UO_1188 (O_1188,N_9825,N_9939);
or UO_1189 (O_1189,N_9846,N_9876);
nand UO_1190 (O_1190,N_9823,N_9904);
or UO_1191 (O_1191,N_9814,N_9996);
nand UO_1192 (O_1192,N_9910,N_9875);
and UO_1193 (O_1193,N_9844,N_9991);
nand UO_1194 (O_1194,N_9823,N_9986);
or UO_1195 (O_1195,N_9830,N_9996);
nand UO_1196 (O_1196,N_9872,N_9800);
nor UO_1197 (O_1197,N_9982,N_9905);
xnor UO_1198 (O_1198,N_9895,N_9907);
nand UO_1199 (O_1199,N_9889,N_9984);
nor UO_1200 (O_1200,N_9943,N_9802);
nor UO_1201 (O_1201,N_9824,N_9905);
or UO_1202 (O_1202,N_9879,N_9813);
or UO_1203 (O_1203,N_9919,N_9924);
and UO_1204 (O_1204,N_9831,N_9875);
and UO_1205 (O_1205,N_9916,N_9873);
or UO_1206 (O_1206,N_9901,N_9849);
nand UO_1207 (O_1207,N_9835,N_9833);
and UO_1208 (O_1208,N_9871,N_9827);
xor UO_1209 (O_1209,N_9936,N_9897);
nor UO_1210 (O_1210,N_9911,N_9914);
or UO_1211 (O_1211,N_9989,N_9832);
nor UO_1212 (O_1212,N_9926,N_9834);
and UO_1213 (O_1213,N_9840,N_9850);
and UO_1214 (O_1214,N_9957,N_9973);
nand UO_1215 (O_1215,N_9933,N_9846);
nor UO_1216 (O_1216,N_9941,N_9871);
nor UO_1217 (O_1217,N_9841,N_9947);
and UO_1218 (O_1218,N_9987,N_9930);
or UO_1219 (O_1219,N_9892,N_9989);
nor UO_1220 (O_1220,N_9930,N_9962);
xor UO_1221 (O_1221,N_9887,N_9910);
and UO_1222 (O_1222,N_9818,N_9830);
or UO_1223 (O_1223,N_9986,N_9826);
xnor UO_1224 (O_1224,N_9914,N_9871);
nand UO_1225 (O_1225,N_9928,N_9908);
nor UO_1226 (O_1226,N_9813,N_9805);
nor UO_1227 (O_1227,N_9882,N_9864);
xnor UO_1228 (O_1228,N_9876,N_9970);
xor UO_1229 (O_1229,N_9993,N_9966);
and UO_1230 (O_1230,N_9882,N_9932);
nor UO_1231 (O_1231,N_9815,N_9989);
nor UO_1232 (O_1232,N_9855,N_9968);
and UO_1233 (O_1233,N_9948,N_9874);
nor UO_1234 (O_1234,N_9853,N_9984);
or UO_1235 (O_1235,N_9983,N_9981);
and UO_1236 (O_1236,N_9968,N_9998);
nor UO_1237 (O_1237,N_9860,N_9980);
and UO_1238 (O_1238,N_9820,N_9854);
or UO_1239 (O_1239,N_9968,N_9987);
xnor UO_1240 (O_1240,N_9826,N_9993);
and UO_1241 (O_1241,N_9853,N_9987);
nand UO_1242 (O_1242,N_9802,N_9971);
nor UO_1243 (O_1243,N_9845,N_9816);
nand UO_1244 (O_1244,N_9924,N_9926);
or UO_1245 (O_1245,N_9902,N_9875);
or UO_1246 (O_1246,N_9814,N_9875);
or UO_1247 (O_1247,N_9895,N_9911);
nand UO_1248 (O_1248,N_9962,N_9837);
nor UO_1249 (O_1249,N_9851,N_9941);
nand UO_1250 (O_1250,N_9945,N_9954);
nand UO_1251 (O_1251,N_9936,N_9885);
nand UO_1252 (O_1252,N_9982,N_9858);
and UO_1253 (O_1253,N_9965,N_9929);
xnor UO_1254 (O_1254,N_9929,N_9988);
nor UO_1255 (O_1255,N_9927,N_9956);
and UO_1256 (O_1256,N_9942,N_9925);
and UO_1257 (O_1257,N_9923,N_9987);
nand UO_1258 (O_1258,N_9999,N_9833);
nand UO_1259 (O_1259,N_9976,N_9913);
nand UO_1260 (O_1260,N_9883,N_9809);
xor UO_1261 (O_1261,N_9969,N_9967);
or UO_1262 (O_1262,N_9929,N_9992);
nand UO_1263 (O_1263,N_9950,N_9857);
and UO_1264 (O_1264,N_9890,N_9881);
and UO_1265 (O_1265,N_9894,N_9968);
nand UO_1266 (O_1266,N_9996,N_9909);
nand UO_1267 (O_1267,N_9952,N_9872);
and UO_1268 (O_1268,N_9805,N_9851);
and UO_1269 (O_1269,N_9837,N_9901);
nor UO_1270 (O_1270,N_9858,N_9826);
and UO_1271 (O_1271,N_9843,N_9814);
xnor UO_1272 (O_1272,N_9962,N_9940);
or UO_1273 (O_1273,N_9954,N_9809);
and UO_1274 (O_1274,N_9961,N_9861);
xor UO_1275 (O_1275,N_9840,N_9987);
and UO_1276 (O_1276,N_9892,N_9839);
or UO_1277 (O_1277,N_9937,N_9909);
nand UO_1278 (O_1278,N_9825,N_9966);
and UO_1279 (O_1279,N_9905,N_9841);
or UO_1280 (O_1280,N_9897,N_9947);
nor UO_1281 (O_1281,N_9865,N_9809);
and UO_1282 (O_1282,N_9859,N_9872);
or UO_1283 (O_1283,N_9958,N_9864);
xnor UO_1284 (O_1284,N_9936,N_9969);
nor UO_1285 (O_1285,N_9996,N_9975);
and UO_1286 (O_1286,N_9919,N_9875);
nand UO_1287 (O_1287,N_9988,N_9852);
or UO_1288 (O_1288,N_9953,N_9816);
or UO_1289 (O_1289,N_9929,N_9802);
nand UO_1290 (O_1290,N_9910,N_9947);
and UO_1291 (O_1291,N_9854,N_9974);
xnor UO_1292 (O_1292,N_9985,N_9808);
nor UO_1293 (O_1293,N_9949,N_9952);
and UO_1294 (O_1294,N_9904,N_9964);
xor UO_1295 (O_1295,N_9894,N_9815);
and UO_1296 (O_1296,N_9804,N_9907);
or UO_1297 (O_1297,N_9892,N_9948);
xnor UO_1298 (O_1298,N_9900,N_9869);
and UO_1299 (O_1299,N_9980,N_9842);
or UO_1300 (O_1300,N_9844,N_9967);
xor UO_1301 (O_1301,N_9805,N_9850);
nand UO_1302 (O_1302,N_9939,N_9831);
or UO_1303 (O_1303,N_9913,N_9900);
nand UO_1304 (O_1304,N_9813,N_9866);
nand UO_1305 (O_1305,N_9806,N_9971);
nand UO_1306 (O_1306,N_9896,N_9919);
nor UO_1307 (O_1307,N_9828,N_9933);
and UO_1308 (O_1308,N_9878,N_9883);
and UO_1309 (O_1309,N_9912,N_9966);
and UO_1310 (O_1310,N_9808,N_9814);
nand UO_1311 (O_1311,N_9800,N_9991);
nand UO_1312 (O_1312,N_9815,N_9910);
nor UO_1313 (O_1313,N_9952,N_9848);
nor UO_1314 (O_1314,N_9948,N_9931);
xor UO_1315 (O_1315,N_9980,N_9852);
xnor UO_1316 (O_1316,N_9937,N_9920);
xnor UO_1317 (O_1317,N_9988,N_9994);
nor UO_1318 (O_1318,N_9896,N_9855);
xnor UO_1319 (O_1319,N_9881,N_9857);
nand UO_1320 (O_1320,N_9991,N_9852);
xor UO_1321 (O_1321,N_9949,N_9976);
xnor UO_1322 (O_1322,N_9834,N_9891);
nand UO_1323 (O_1323,N_9807,N_9871);
or UO_1324 (O_1324,N_9809,N_9956);
nand UO_1325 (O_1325,N_9849,N_9878);
nand UO_1326 (O_1326,N_9968,N_9919);
xor UO_1327 (O_1327,N_9951,N_9813);
nor UO_1328 (O_1328,N_9860,N_9854);
nor UO_1329 (O_1329,N_9892,N_9956);
nor UO_1330 (O_1330,N_9819,N_9963);
and UO_1331 (O_1331,N_9949,N_9810);
nor UO_1332 (O_1332,N_9939,N_9869);
nand UO_1333 (O_1333,N_9884,N_9995);
and UO_1334 (O_1334,N_9835,N_9857);
or UO_1335 (O_1335,N_9950,N_9915);
nor UO_1336 (O_1336,N_9994,N_9845);
nor UO_1337 (O_1337,N_9858,N_9915);
xor UO_1338 (O_1338,N_9957,N_9838);
nand UO_1339 (O_1339,N_9804,N_9926);
nand UO_1340 (O_1340,N_9856,N_9901);
or UO_1341 (O_1341,N_9984,N_9981);
or UO_1342 (O_1342,N_9845,N_9811);
xnor UO_1343 (O_1343,N_9869,N_9801);
xor UO_1344 (O_1344,N_9960,N_9857);
nand UO_1345 (O_1345,N_9912,N_9863);
or UO_1346 (O_1346,N_9802,N_9882);
or UO_1347 (O_1347,N_9897,N_9868);
and UO_1348 (O_1348,N_9990,N_9819);
nor UO_1349 (O_1349,N_9923,N_9823);
and UO_1350 (O_1350,N_9830,N_9886);
xor UO_1351 (O_1351,N_9879,N_9958);
nand UO_1352 (O_1352,N_9992,N_9821);
nor UO_1353 (O_1353,N_9928,N_9873);
or UO_1354 (O_1354,N_9817,N_9973);
xnor UO_1355 (O_1355,N_9954,N_9965);
or UO_1356 (O_1356,N_9900,N_9951);
nor UO_1357 (O_1357,N_9980,N_9819);
nand UO_1358 (O_1358,N_9980,N_9886);
nor UO_1359 (O_1359,N_9979,N_9942);
or UO_1360 (O_1360,N_9896,N_9819);
nand UO_1361 (O_1361,N_9867,N_9842);
and UO_1362 (O_1362,N_9976,N_9840);
nand UO_1363 (O_1363,N_9919,N_9805);
xor UO_1364 (O_1364,N_9944,N_9885);
or UO_1365 (O_1365,N_9825,N_9866);
or UO_1366 (O_1366,N_9877,N_9865);
nor UO_1367 (O_1367,N_9867,N_9974);
nor UO_1368 (O_1368,N_9941,N_9935);
nand UO_1369 (O_1369,N_9821,N_9837);
nand UO_1370 (O_1370,N_9802,N_9927);
xnor UO_1371 (O_1371,N_9936,N_9806);
nand UO_1372 (O_1372,N_9974,N_9960);
and UO_1373 (O_1373,N_9940,N_9890);
nand UO_1374 (O_1374,N_9828,N_9873);
nand UO_1375 (O_1375,N_9967,N_9852);
and UO_1376 (O_1376,N_9938,N_9899);
nor UO_1377 (O_1377,N_9879,N_9866);
nor UO_1378 (O_1378,N_9878,N_9843);
nand UO_1379 (O_1379,N_9866,N_9839);
or UO_1380 (O_1380,N_9936,N_9841);
nand UO_1381 (O_1381,N_9842,N_9922);
xnor UO_1382 (O_1382,N_9849,N_9951);
or UO_1383 (O_1383,N_9939,N_9823);
nand UO_1384 (O_1384,N_9986,N_9827);
or UO_1385 (O_1385,N_9914,N_9915);
nand UO_1386 (O_1386,N_9915,N_9936);
xor UO_1387 (O_1387,N_9828,N_9864);
nand UO_1388 (O_1388,N_9872,N_9932);
or UO_1389 (O_1389,N_9982,N_9998);
or UO_1390 (O_1390,N_9830,N_9969);
or UO_1391 (O_1391,N_9823,N_9896);
and UO_1392 (O_1392,N_9947,N_9998);
or UO_1393 (O_1393,N_9991,N_9918);
xor UO_1394 (O_1394,N_9998,N_9920);
and UO_1395 (O_1395,N_9984,N_9933);
nor UO_1396 (O_1396,N_9966,N_9847);
nor UO_1397 (O_1397,N_9956,N_9845);
nand UO_1398 (O_1398,N_9969,N_9928);
nor UO_1399 (O_1399,N_9929,N_9826);
nand UO_1400 (O_1400,N_9951,N_9912);
or UO_1401 (O_1401,N_9894,N_9823);
xnor UO_1402 (O_1402,N_9889,N_9907);
or UO_1403 (O_1403,N_9947,N_9842);
and UO_1404 (O_1404,N_9990,N_9901);
and UO_1405 (O_1405,N_9830,N_9964);
or UO_1406 (O_1406,N_9935,N_9819);
nand UO_1407 (O_1407,N_9824,N_9976);
and UO_1408 (O_1408,N_9870,N_9883);
and UO_1409 (O_1409,N_9918,N_9806);
nand UO_1410 (O_1410,N_9961,N_9981);
nor UO_1411 (O_1411,N_9814,N_9835);
or UO_1412 (O_1412,N_9837,N_9942);
or UO_1413 (O_1413,N_9929,N_9878);
xnor UO_1414 (O_1414,N_9972,N_9885);
and UO_1415 (O_1415,N_9912,N_9985);
or UO_1416 (O_1416,N_9883,N_9941);
nor UO_1417 (O_1417,N_9857,N_9903);
and UO_1418 (O_1418,N_9950,N_9922);
nor UO_1419 (O_1419,N_9807,N_9950);
and UO_1420 (O_1420,N_9897,N_9978);
or UO_1421 (O_1421,N_9991,N_9966);
nor UO_1422 (O_1422,N_9946,N_9888);
and UO_1423 (O_1423,N_9937,N_9801);
nor UO_1424 (O_1424,N_9916,N_9928);
nand UO_1425 (O_1425,N_9815,N_9936);
nand UO_1426 (O_1426,N_9955,N_9946);
or UO_1427 (O_1427,N_9989,N_9999);
or UO_1428 (O_1428,N_9892,N_9832);
xnor UO_1429 (O_1429,N_9987,N_9990);
xor UO_1430 (O_1430,N_9899,N_9941);
or UO_1431 (O_1431,N_9998,N_9921);
and UO_1432 (O_1432,N_9999,N_9986);
nand UO_1433 (O_1433,N_9812,N_9898);
and UO_1434 (O_1434,N_9836,N_9921);
and UO_1435 (O_1435,N_9991,N_9927);
nor UO_1436 (O_1436,N_9984,N_9922);
xnor UO_1437 (O_1437,N_9943,N_9804);
or UO_1438 (O_1438,N_9832,N_9916);
xnor UO_1439 (O_1439,N_9855,N_9834);
and UO_1440 (O_1440,N_9981,N_9874);
nand UO_1441 (O_1441,N_9922,N_9911);
and UO_1442 (O_1442,N_9837,N_9878);
and UO_1443 (O_1443,N_9852,N_9945);
nand UO_1444 (O_1444,N_9935,N_9869);
nor UO_1445 (O_1445,N_9844,N_9883);
or UO_1446 (O_1446,N_9880,N_9953);
nand UO_1447 (O_1447,N_9858,N_9823);
xnor UO_1448 (O_1448,N_9824,N_9987);
or UO_1449 (O_1449,N_9963,N_9864);
xnor UO_1450 (O_1450,N_9991,N_9866);
or UO_1451 (O_1451,N_9994,N_9992);
nand UO_1452 (O_1452,N_9813,N_9913);
xnor UO_1453 (O_1453,N_9845,N_9966);
and UO_1454 (O_1454,N_9870,N_9850);
xor UO_1455 (O_1455,N_9959,N_9920);
and UO_1456 (O_1456,N_9981,N_9958);
nand UO_1457 (O_1457,N_9840,N_9957);
nand UO_1458 (O_1458,N_9822,N_9998);
and UO_1459 (O_1459,N_9811,N_9869);
xnor UO_1460 (O_1460,N_9981,N_9845);
nand UO_1461 (O_1461,N_9962,N_9977);
or UO_1462 (O_1462,N_9866,N_9908);
nor UO_1463 (O_1463,N_9832,N_9978);
nor UO_1464 (O_1464,N_9884,N_9800);
or UO_1465 (O_1465,N_9966,N_9806);
xnor UO_1466 (O_1466,N_9910,N_9836);
nand UO_1467 (O_1467,N_9836,N_9813);
and UO_1468 (O_1468,N_9855,N_9835);
nor UO_1469 (O_1469,N_9869,N_9813);
xnor UO_1470 (O_1470,N_9964,N_9875);
nand UO_1471 (O_1471,N_9801,N_9936);
xnor UO_1472 (O_1472,N_9983,N_9897);
nor UO_1473 (O_1473,N_9881,N_9840);
or UO_1474 (O_1474,N_9995,N_9890);
and UO_1475 (O_1475,N_9811,N_9832);
and UO_1476 (O_1476,N_9989,N_9947);
or UO_1477 (O_1477,N_9822,N_9966);
or UO_1478 (O_1478,N_9828,N_9858);
or UO_1479 (O_1479,N_9890,N_9996);
or UO_1480 (O_1480,N_9984,N_9934);
nand UO_1481 (O_1481,N_9835,N_9868);
nor UO_1482 (O_1482,N_9984,N_9832);
or UO_1483 (O_1483,N_9854,N_9800);
nor UO_1484 (O_1484,N_9899,N_9999);
or UO_1485 (O_1485,N_9837,N_9914);
nand UO_1486 (O_1486,N_9826,N_9920);
nor UO_1487 (O_1487,N_9919,N_9862);
or UO_1488 (O_1488,N_9911,N_9844);
nand UO_1489 (O_1489,N_9987,N_9962);
nor UO_1490 (O_1490,N_9909,N_9929);
nor UO_1491 (O_1491,N_9814,N_9941);
nor UO_1492 (O_1492,N_9913,N_9959);
xor UO_1493 (O_1493,N_9964,N_9859);
nor UO_1494 (O_1494,N_9890,N_9926);
xnor UO_1495 (O_1495,N_9866,N_9865);
nor UO_1496 (O_1496,N_9898,N_9955);
nor UO_1497 (O_1497,N_9930,N_9939);
xor UO_1498 (O_1498,N_9961,N_9956);
and UO_1499 (O_1499,N_9909,N_9962);
endmodule