module basic_2500_25000_3000_5_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_2331,In_1089);
nand U1 (N_1,In_1741,In_1194);
nand U2 (N_2,In_166,In_2487);
or U3 (N_3,In_610,In_87);
and U4 (N_4,In_514,In_795);
nor U5 (N_5,In_2248,In_778);
nand U6 (N_6,In_1158,In_1857);
or U7 (N_7,In_2389,In_2313);
and U8 (N_8,In_1858,In_1892);
nand U9 (N_9,In_2268,In_1161);
and U10 (N_10,In_937,In_2381);
or U11 (N_11,In_2163,In_2214);
or U12 (N_12,In_32,In_1203);
nand U13 (N_13,In_225,In_1528);
and U14 (N_14,In_326,In_1129);
and U15 (N_15,In_773,In_705);
nor U16 (N_16,In_1980,In_1647);
or U17 (N_17,In_940,In_132);
nor U18 (N_18,In_53,In_267);
and U19 (N_19,In_1295,In_998);
nand U20 (N_20,In_1767,In_2024);
and U21 (N_21,In_608,In_962);
nand U22 (N_22,In_879,In_1077);
nand U23 (N_23,In_2178,In_1974);
and U24 (N_24,In_40,In_766);
and U25 (N_25,In_1587,In_1135);
and U26 (N_26,In_241,In_896);
nor U27 (N_27,In_868,In_2022);
or U28 (N_28,In_1464,In_1398);
nand U29 (N_29,In_1111,In_487);
and U30 (N_30,In_1227,In_1414);
and U31 (N_31,In_299,In_1137);
and U32 (N_32,In_2458,In_2485);
and U33 (N_33,In_1032,In_29);
nor U34 (N_34,In_392,In_2252);
and U35 (N_35,In_2049,In_2475);
or U36 (N_36,In_1967,In_1621);
nand U37 (N_37,In_855,In_353);
or U38 (N_38,In_1831,In_1010);
or U39 (N_39,In_1037,In_61);
nand U40 (N_40,In_1677,In_447);
and U41 (N_41,In_2366,In_370);
nand U42 (N_42,In_2488,In_1512);
or U43 (N_43,In_1029,In_1814);
nand U44 (N_44,In_1257,In_154);
nand U45 (N_45,In_618,In_995);
nand U46 (N_46,In_741,In_967);
nor U47 (N_47,In_537,In_849);
and U48 (N_48,In_1365,In_546);
nand U49 (N_49,In_2016,In_494);
or U50 (N_50,In_1067,In_1164);
nor U51 (N_51,In_1792,In_697);
or U52 (N_52,In_170,In_1810);
or U53 (N_53,In_1875,In_942);
nand U54 (N_54,In_151,In_456);
or U55 (N_55,In_760,In_2284);
nand U56 (N_56,In_1688,In_1175);
nor U57 (N_57,In_759,In_2136);
nor U58 (N_58,In_2028,In_880);
and U59 (N_59,In_383,In_851);
and U60 (N_60,In_1769,In_1726);
nand U61 (N_61,In_1494,In_804);
nand U62 (N_62,In_1133,In_2274);
and U63 (N_63,In_1933,In_1446);
or U64 (N_64,In_2186,In_2143);
nor U65 (N_65,In_2081,In_8);
nand U66 (N_66,In_1379,In_934);
nand U67 (N_67,In_417,In_1460);
or U68 (N_68,In_2399,In_708);
nand U69 (N_69,In_2251,In_191);
nand U70 (N_70,In_1599,In_2020);
and U71 (N_71,In_347,In_289);
nand U72 (N_72,In_2447,In_144);
nor U73 (N_73,In_1901,In_1330);
and U74 (N_74,In_346,In_2121);
or U75 (N_75,In_905,In_526);
nor U76 (N_76,In_1056,In_109);
or U77 (N_77,In_2111,In_1333);
nor U78 (N_78,In_683,In_70);
nand U79 (N_79,In_1160,In_2319);
and U80 (N_80,In_1180,In_914);
nor U81 (N_81,In_0,In_156);
nor U82 (N_82,In_418,In_1830);
or U83 (N_83,In_949,In_1283);
nand U84 (N_84,In_1562,In_2437);
and U85 (N_85,In_452,In_801);
nor U86 (N_86,In_727,In_925);
nor U87 (N_87,In_1438,In_2308);
or U88 (N_88,In_31,In_1594);
and U89 (N_89,In_1361,In_739);
nand U90 (N_90,In_1261,In_1612);
nand U91 (N_91,In_2005,In_1115);
and U92 (N_92,In_1793,In_1891);
nor U93 (N_93,In_1760,In_567);
and U94 (N_94,In_2289,In_1791);
nor U95 (N_95,In_1863,In_2237);
or U96 (N_96,In_438,In_1656);
or U97 (N_97,In_2117,In_826);
nand U98 (N_98,In_1013,In_1313);
xor U99 (N_99,In_627,In_997);
nor U100 (N_100,In_1480,In_2066);
or U101 (N_101,In_839,In_4);
and U102 (N_102,In_823,In_1752);
or U103 (N_103,In_1452,In_1976);
and U104 (N_104,In_510,In_195);
nand U105 (N_105,In_460,In_827);
or U106 (N_106,In_1396,In_374);
nand U107 (N_107,In_2046,In_2135);
nor U108 (N_108,In_2341,In_990);
or U109 (N_109,In_2131,In_348);
nor U110 (N_110,In_677,In_2346);
and U111 (N_111,In_127,In_396);
nor U112 (N_112,In_571,In_883);
xnor U113 (N_113,In_954,In_2188);
and U114 (N_114,In_1615,In_128);
nor U115 (N_115,In_1215,In_55);
nor U116 (N_116,In_1420,In_2041);
nand U117 (N_117,In_405,In_490);
nor U118 (N_118,In_2469,In_1201);
nand U119 (N_119,In_163,In_1531);
or U120 (N_120,In_1335,In_2197);
and U121 (N_121,In_798,In_116);
nor U122 (N_122,In_290,In_2013);
or U123 (N_123,In_2257,In_1385);
nand U124 (N_124,In_1181,In_1711);
nor U125 (N_125,In_72,In_743);
or U126 (N_126,In_1900,In_1950);
and U127 (N_127,In_733,In_1883);
xor U128 (N_128,In_122,In_384);
nor U129 (N_129,In_312,In_330);
or U130 (N_130,In_1795,In_202);
nor U131 (N_131,In_1329,In_139);
nand U132 (N_132,In_1345,In_1870);
or U133 (N_133,In_1008,In_10);
or U134 (N_134,In_2004,In_714);
nand U135 (N_135,In_2153,In_1747);
nor U136 (N_136,In_696,In_2281);
nor U137 (N_137,In_785,In_2333);
or U138 (N_138,In_1202,In_1785);
nor U139 (N_139,In_853,In_797);
nor U140 (N_140,In_2420,In_1788);
or U141 (N_141,In_2150,In_2269);
nand U142 (N_142,In_479,In_367);
nand U143 (N_143,In_1255,In_2369);
nand U144 (N_144,In_1191,In_2361);
or U145 (N_145,In_820,In_782);
or U146 (N_146,In_616,In_219);
or U147 (N_147,In_2061,In_1461);
nor U148 (N_148,In_1300,In_2222);
or U149 (N_149,In_953,In_1282);
nand U150 (N_150,In_2109,In_544);
or U151 (N_151,In_2423,In_520);
nor U152 (N_152,In_2255,In_588);
nor U153 (N_153,In_1849,In_310);
nand U154 (N_154,In_483,In_898);
nor U155 (N_155,In_331,In_1616);
and U156 (N_156,In_1510,In_1211);
or U157 (N_157,In_1888,In_2037);
and U158 (N_158,In_56,In_2076);
or U159 (N_159,In_506,In_1312);
and U160 (N_160,In_1144,In_1679);
or U161 (N_161,In_11,In_388);
nor U162 (N_162,In_1840,In_2134);
or U163 (N_163,In_1664,In_253);
nand U164 (N_164,In_1811,In_278);
nand U165 (N_165,In_1694,In_2450);
or U166 (N_166,In_1479,In_889);
and U167 (N_167,In_1435,In_687);
nor U168 (N_168,In_1439,In_2315);
and U169 (N_169,In_266,In_1733);
and U170 (N_170,In_1039,In_2021);
or U171 (N_171,In_583,In_1896);
nand U172 (N_172,In_956,In_297);
or U173 (N_173,In_379,In_524);
and U174 (N_174,In_1455,In_287);
nand U175 (N_175,In_1861,In_1258);
or U176 (N_176,In_1337,In_1910);
nand U177 (N_177,In_1586,In_448);
or U178 (N_178,In_539,In_357);
xor U179 (N_179,In_115,In_1756);
nand U180 (N_180,In_1824,In_295);
nor U181 (N_181,In_1798,In_78);
nand U182 (N_182,In_1513,In_1514);
or U183 (N_183,In_2064,In_1604);
or U184 (N_184,In_763,In_651);
and U185 (N_185,In_817,In_319);
nor U186 (N_186,In_2035,In_265);
xor U187 (N_187,In_1815,In_2082);
nand U188 (N_188,In_1190,In_82);
and U189 (N_189,In_1443,In_1865);
and U190 (N_190,In_1,In_1122);
nand U191 (N_191,In_499,In_2164);
and U192 (N_192,In_716,In_196);
and U193 (N_193,In_179,In_1212);
or U194 (N_194,In_2386,In_2260);
nor U195 (N_195,In_796,In_1881);
nor U196 (N_196,In_1557,In_437);
nor U197 (N_197,In_863,In_1065);
and U198 (N_198,In_292,In_375);
and U199 (N_199,In_2122,In_1341);
or U200 (N_200,In_469,In_1059);
or U201 (N_201,In_135,In_1851);
or U202 (N_202,In_1736,In_1620);
nand U203 (N_203,In_865,In_948);
or U204 (N_204,In_1526,In_790);
or U205 (N_205,In_543,In_1041);
or U206 (N_206,In_811,In_233);
or U207 (N_207,In_1958,In_650);
nor U208 (N_208,In_21,In_1197);
nand U209 (N_209,In_1961,In_1034);
and U210 (N_210,In_1825,In_598);
and U211 (N_211,In_933,In_1229);
nand U212 (N_212,In_1252,In_736);
and U213 (N_213,In_108,In_1001);
or U214 (N_214,In_2261,In_908);
and U215 (N_215,In_1102,In_1787);
nand U216 (N_216,In_393,In_877);
nand U217 (N_217,In_1306,In_1318);
and U218 (N_218,In_723,In_625);
nand U219 (N_219,In_1482,In_2492);
nor U220 (N_220,In_1305,In_525);
and U221 (N_221,In_1167,In_1775);
or U222 (N_222,In_916,In_2123);
xor U223 (N_223,In_1240,In_83);
nor U224 (N_224,In_2091,In_2193);
and U225 (N_225,In_919,In_198);
nor U226 (N_226,In_400,In_1299);
or U227 (N_227,In_1912,In_2031);
nand U228 (N_228,In_1263,In_1713);
nor U229 (N_229,In_664,In_1945);
and U230 (N_230,In_1874,In_935);
and U231 (N_231,In_57,In_1689);
or U232 (N_232,In_986,In_275);
and U233 (N_233,In_2471,In_888);
nor U234 (N_234,In_1107,In_1415);
nor U235 (N_235,In_1275,In_614);
xnor U236 (N_236,In_1062,In_2050);
and U237 (N_237,In_1497,In_239);
and U238 (N_238,In_693,In_1907);
and U239 (N_239,In_467,In_836);
and U240 (N_240,In_726,In_1718);
or U241 (N_241,In_1436,In_1651);
xor U242 (N_242,In_1925,In_1998);
nand U243 (N_243,In_609,In_1987);
or U244 (N_244,In_646,In_2065);
nor U245 (N_245,In_459,In_1241);
nand U246 (N_246,In_1902,In_2154);
or U247 (N_247,In_2415,In_1570);
nand U248 (N_248,In_1988,In_1082);
nor U249 (N_249,In_3,In_2069);
nor U250 (N_250,In_1459,In_1071);
nand U251 (N_251,In_209,In_1533);
nor U252 (N_252,In_768,In_1649);
nor U253 (N_253,In_2406,In_407);
nand U254 (N_254,In_1289,In_1448);
nor U255 (N_255,In_2497,In_2232);
or U256 (N_256,In_498,In_1710);
nand U257 (N_257,In_1388,In_2451);
and U258 (N_258,In_1908,In_2208);
or U259 (N_259,In_1611,In_1696);
nor U260 (N_260,In_2092,In_2132);
nor U261 (N_261,In_362,In_1408);
nor U262 (N_262,In_737,In_2337);
nand U263 (N_263,In_495,In_378);
nand U264 (N_264,In_1050,In_2342);
nor U265 (N_265,In_1310,In_2089);
and U266 (N_266,In_1198,In_114);
nor U267 (N_267,In_1035,In_2396);
or U268 (N_268,In_965,In_423);
or U269 (N_269,In_1165,In_1284);
and U270 (N_270,In_812,In_957);
xnor U271 (N_271,In_762,In_837);
or U272 (N_272,In_2039,In_694);
nor U273 (N_273,In_703,In_277);
or U274 (N_274,In_1847,In_2491);
nand U275 (N_275,In_951,In_1880);
nor U276 (N_276,In_634,In_780);
nor U277 (N_277,In_1622,In_2280);
and U278 (N_278,In_332,In_2336);
or U279 (N_279,In_1639,In_1394);
or U280 (N_280,In_2340,In_1618);
or U281 (N_281,In_2171,In_1384);
or U282 (N_282,In_2124,In_234);
or U283 (N_283,In_745,In_1672);
nand U284 (N_284,In_232,In_1937);
nand U285 (N_285,In_2431,In_1975);
nand U286 (N_286,In_1632,In_799);
and U287 (N_287,In_2201,In_1027);
and U288 (N_288,In_2427,In_2168);
nor U289 (N_289,In_1952,In_2086);
or U290 (N_290,In_2419,In_893);
nand U291 (N_291,In_38,In_787);
or U292 (N_292,In_591,In_186);
nand U293 (N_293,In_2120,In_2263);
or U294 (N_294,In_471,In_1321);
nand U295 (N_295,In_1078,In_1500);
xor U296 (N_296,In_803,In_1703);
nand U297 (N_297,In_770,In_556);
or U298 (N_298,In_1488,In_977);
nor U299 (N_299,In_1100,In_1354);
xnor U300 (N_300,In_1231,In_1422);
nand U301 (N_301,In_1182,In_248);
and U302 (N_302,In_692,In_203);
nand U303 (N_303,In_2101,In_1572);
xor U304 (N_304,In_1214,In_1977);
nor U305 (N_305,In_1614,In_1105);
nand U306 (N_306,In_79,In_1650);
and U307 (N_307,In_590,In_1272);
nand U308 (N_308,In_800,In_515);
or U309 (N_309,In_806,In_1924);
and U310 (N_310,In_488,In_1501);
nor U311 (N_311,In_1508,In_1021);
or U312 (N_312,In_2177,In_831);
and U313 (N_313,In_991,In_527);
nor U314 (N_314,In_324,In_2138);
nor U315 (N_315,In_1023,In_1555);
and U316 (N_316,In_1237,In_298);
nor U317 (N_317,In_1890,In_1338);
or U318 (N_318,In_861,In_2058);
or U319 (N_319,In_1173,In_718);
nor U320 (N_320,In_171,In_2395);
and U321 (N_321,In_1085,In_496);
and U322 (N_322,In_1274,In_1151);
nor U323 (N_323,In_874,In_1685);
nor U324 (N_324,In_1364,In_476);
and U325 (N_325,In_22,In_403);
or U326 (N_326,In_1625,In_1123);
nor U327 (N_327,In_7,In_23);
and U328 (N_328,In_915,In_1728);
nand U329 (N_329,In_1166,In_913);
nand U330 (N_330,In_141,In_1049);
nor U331 (N_331,In_1324,In_660);
nand U332 (N_332,In_1866,In_1682);
nor U333 (N_333,In_2436,In_112);
nand U334 (N_334,In_895,In_2080);
or U335 (N_335,In_601,In_848);
nor U336 (N_336,In_1496,In_2302);
or U337 (N_337,In_2026,In_607);
or U338 (N_338,In_2115,In_307);
or U339 (N_339,In_2094,In_1302);
nor U340 (N_340,In_1644,In_386);
nand U341 (N_341,In_1964,In_1206);
or U342 (N_342,In_140,In_2235);
and U343 (N_343,In_2464,In_486);
and U344 (N_344,In_564,In_1566);
or U345 (N_345,In_103,In_2438);
and U346 (N_346,In_2225,In_2481);
or U347 (N_347,In_2435,In_256);
or U348 (N_348,In_1771,In_931);
xor U349 (N_349,In_238,In_1705);
and U350 (N_350,In_221,In_1954);
and U351 (N_351,In_200,In_1259);
or U352 (N_352,In_124,In_981);
nor U353 (N_353,In_1737,In_779);
and U354 (N_354,In_30,In_1162);
nor U355 (N_355,In_2303,In_1447);
nand U356 (N_356,In_2465,In_1442);
nor U357 (N_357,In_1568,In_1233);
and U358 (N_358,In_1405,In_1727);
and U359 (N_359,In_2353,In_628);
nand U360 (N_360,In_1906,In_258);
nand U361 (N_361,In_1139,In_1574);
and U362 (N_362,In_2063,In_969);
or U363 (N_363,In_13,In_2157);
nor U364 (N_364,In_1483,In_2334);
and U365 (N_365,In_80,In_2459);
nor U366 (N_366,In_1174,In_1404);
and U367 (N_367,In_629,In_581);
nor U368 (N_368,In_380,In_1163);
nand U369 (N_369,In_2452,In_2314);
and U370 (N_370,In_2417,In_1999);
nand U371 (N_371,In_2118,In_1005);
nor U372 (N_372,In_1380,In_257);
nor U373 (N_373,In_1934,In_767);
nand U374 (N_374,In_1245,In_453);
and U375 (N_375,In_1040,In_1953);
nor U376 (N_376,In_301,In_389);
nor U377 (N_377,In_71,In_81);
nand U378 (N_378,In_279,In_2070);
and U379 (N_379,In_2011,In_1783);
or U380 (N_380,In_2180,In_512);
and U381 (N_381,In_104,In_1235);
or U382 (N_382,In_1402,In_1652);
and U383 (N_383,In_833,In_864);
and U384 (N_384,In_603,In_784);
and U385 (N_385,In_1521,In_887);
or U386 (N_386,In_769,In_2279);
or U387 (N_387,In_254,In_1228);
nand U388 (N_388,In_2098,In_268);
nor U389 (N_389,In_2062,In_2329);
xor U390 (N_390,In_1707,In_2116);
and U391 (N_391,In_1764,In_2462);
and U392 (N_392,In_1602,In_1375);
nand U393 (N_393,In_33,In_223);
nand U394 (N_394,In_1445,In_2047);
nor U395 (N_395,In_36,In_1308);
nor U396 (N_396,In_706,In_1853);
nand U397 (N_397,In_305,In_1178);
nand U398 (N_398,In_722,In_2467);
nor U399 (N_399,In_1018,In_356);
nor U400 (N_400,In_1749,In_1561);
nor U401 (N_401,In_412,In_316);
nand U402 (N_402,In_449,In_2466);
or U403 (N_403,In_335,In_2344);
and U404 (N_404,In_1592,In_1267);
nand U405 (N_405,In_1316,In_2311);
or U406 (N_406,In_489,In_2205);
nor U407 (N_407,In_1800,In_1583);
nor U408 (N_408,In_783,In_2128);
and U409 (N_409,In_1556,In_871);
or U410 (N_410,In_1236,In_1803);
and U411 (N_411,In_441,In_398);
nand U412 (N_412,In_409,In_1700);
or U413 (N_413,In_1350,In_1667);
xor U414 (N_414,In_427,In_2290);
or U415 (N_415,In_1894,In_1362);
and U416 (N_416,In_2448,In_130);
nand U417 (N_417,In_2495,In_434);
or U418 (N_418,In_2218,In_2317);
or U419 (N_419,In_1843,In_1581);
nand U420 (N_420,In_1025,In_2213);
nand U421 (N_421,In_648,In_1841);
or U422 (N_422,In_1079,In_867);
and U423 (N_423,In_983,In_2159);
nand U424 (N_424,In_1758,In_1216);
nor U425 (N_425,In_1673,In_917);
nor U426 (N_426,In_158,In_1844);
nor U427 (N_427,In_2392,In_2189);
or U428 (N_428,In_2141,In_1186);
or U429 (N_429,In_758,In_270);
nand U430 (N_430,In_1797,In_1484);
nand U431 (N_431,In_1817,In_1732);
xor U432 (N_432,In_182,In_507);
nor U433 (N_433,In_586,In_695);
nor U434 (N_434,In_1991,In_824);
or U435 (N_435,In_2038,In_1820);
or U436 (N_436,In_2084,In_344);
nand U437 (N_437,In_832,In_2191);
and U438 (N_438,In_1486,In_1932);
or U439 (N_439,In_633,In_549);
nor U440 (N_440,In_1406,In_1774);
nor U441 (N_441,In_710,In_243);
nand U442 (N_442,In_358,In_342);
or U443 (N_443,In_2158,In_1168);
nand U444 (N_444,In_2221,In_894);
and U445 (N_445,In_584,In_1061);
and U446 (N_446,In_884,In_435);
or U447 (N_447,In_462,In_1823);
and U448 (N_448,In_1850,In_1692);
and U449 (N_449,In_734,In_1715);
or U450 (N_450,In_2287,In_2402);
nor U451 (N_451,In_966,In_772);
or U452 (N_452,In_2209,In_74);
and U453 (N_453,In_939,In_505);
and U454 (N_454,In_250,In_214);
nand U455 (N_455,In_1642,In_136);
or U456 (N_456,In_2383,In_1030);
or U457 (N_457,In_2348,In_2434);
or U458 (N_458,In_465,In_1346);
and U459 (N_459,In_1829,In_580);
nand U460 (N_460,In_174,In_408);
or U461 (N_461,In_318,In_2053);
nor U462 (N_462,In_272,In_1262);
or U463 (N_463,In_1899,In_261);
nand U464 (N_464,In_2190,In_1326);
or U465 (N_465,In_216,In_1268);
nor U466 (N_466,In_363,In_50);
nand U467 (N_467,In_1332,In_2085);
nand U468 (N_468,In_1453,In_1947);
and U469 (N_469,In_674,In_1805);
or U470 (N_470,In_2277,In_903);
or U471 (N_471,In_1670,In_1813);
nand U472 (N_472,In_2107,In_1550);
or U473 (N_473,In_1596,In_1544);
nand U474 (N_474,In_475,In_1256);
and U475 (N_475,In_876,In_315);
nor U476 (N_476,In_351,In_1294);
or U477 (N_477,In_1011,In_2113);
nand U478 (N_478,In_2127,In_1982);
and U479 (N_479,In_1303,In_1224);
and U480 (N_480,In_2234,In_818);
and U481 (N_481,In_1426,In_2439);
nand U482 (N_482,In_242,In_1745);
nand U483 (N_483,In_125,In_1681);
nor U484 (N_484,In_540,In_2033);
nand U485 (N_485,In_1893,In_881);
or U486 (N_486,In_1949,In_1753);
nor U487 (N_487,In_2099,In_1152);
nor U488 (N_488,In_1470,In_1686);
and U489 (N_489,In_439,In_2421);
xnor U490 (N_490,In_2278,In_1327);
and U491 (N_491,In_1099,In_2322);
or U492 (N_492,In_943,In_2199);
nor U493 (N_493,In_1918,In_645);
nor U494 (N_494,In_805,In_317);
nand U495 (N_495,In_667,In_431);
nor U496 (N_496,In_1370,In_1200);
nor U497 (N_497,In_1648,In_1789);
nand U498 (N_498,In_1293,In_1449);
nor U499 (N_499,In_1565,In_2430);
nor U500 (N_500,In_982,In_2242);
nor U501 (N_501,In_404,In_280);
and U502 (N_502,In_2007,In_680);
nand U503 (N_503,In_1757,In_548);
or U504 (N_504,In_2429,In_1898);
nand U505 (N_505,In_2025,In_1802);
nor U506 (N_506,In_1369,In_1645);
or U507 (N_507,In_1087,In_492);
and U508 (N_508,In_1022,In_1608);
or U509 (N_509,In_1605,In_1489);
or U510 (N_510,In_1585,In_1979);
nor U511 (N_511,In_578,In_1659);
or U512 (N_512,In_989,In_194);
or U513 (N_513,In_602,In_1377);
or U514 (N_514,In_184,In_75);
and U515 (N_515,In_2102,In_466);
nor U516 (N_516,In_123,In_1885);
nor U517 (N_517,In_2270,In_1780);
nor U518 (N_518,In_328,In_1524);
nor U519 (N_519,In_808,In_1560);
and U520 (N_520,In_2343,In_996);
and U521 (N_521,In_207,In_968);
nand U522 (N_522,In_519,In_1996);
nor U523 (N_523,In_77,In_1428);
xnor U524 (N_524,In_89,In_51);
nand U525 (N_525,In_1413,In_1909);
nand U526 (N_526,In_137,In_1712);
nand U527 (N_527,In_1141,In_1238);
nand U528 (N_528,In_2352,In_2262);
nor U529 (N_529,In_2489,In_561);
nand U530 (N_530,In_2215,In_657);
nor U531 (N_531,In_518,In_1535);
nor U532 (N_532,In_1244,In_2184);
and U533 (N_533,In_251,In_39);
and U534 (N_534,In_1019,In_185);
or U535 (N_535,In_1717,In_2477);
or U536 (N_536,In_2145,In_576);
nand U537 (N_537,In_678,In_2172);
and U538 (N_538,In_1142,In_24);
nor U539 (N_539,In_1383,In_929);
nand U540 (N_540,In_978,In_269);
nand U541 (N_541,In_2354,In_1125);
nor U542 (N_542,In_813,In_497);
and U543 (N_543,In_1119,In_160);
nor U544 (N_544,In_2140,In_624);
and U545 (N_545,In_976,In_1623);
and U546 (N_546,In_1522,In_834);
nor U547 (N_547,In_1495,In_302);
or U548 (N_548,In_2227,In_2265);
and U549 (N_549,In_1609,In_1702);
and U550 (N_550,In_161,In_1015);
nor U551 (N_551,In_1624,In_921);
nor U552 (N_552,In_49,In_1897);
nor U553 (N_553,In_2008,In_1088);
nor U554 (N_554,In_1835,In_461);
nor U555 (N_555,In_1093,In_2388);
nand U556 (N_556,In_890,In_1355);
nand U557 (N_557,In_789,In_1580);
nand U558 (N_558,In_259,In_410);
nor U559 (N_559,In_426,In_1818);
xor U560 (N_560,In_1914,In_1440);
and U561 (N_561,In_558,In_2236);
and U562 (N_562,In_1051,In_2097);
nand U563 (N_563,In_1114,In_900);
and U564 (N_564,In_2241,In_1411);
and U565 (N_565,In_821,In_700);
and U566 (N_566,In_1334,In_1916);
nand U567 (N_567,In_1269,In_2240);
or U568 (N_568,In_5,In_2418);
and U569 (N_569,In_1832,In_2440);
nor U570 (N_570,In_2137,In_188);
nand U571 (N_571,In_1873,In_1666);
nand U572 (N_572,In_938,In_445);
or U573 (N_573,In_193,In_1734);
nand U574 (N_574,In_2359,In_511);
and U575 (N_575,In_670,In_669);
nor U576 (N_576,In_273,In_926);
nand U577 (N_577,In_1220,In_1080);
nor U578 (N_578,In_464,In_240);
nor U579 (N_579,In_177,In_1809);
and U580 (N_580,In_183,In_1113);
nor U581 (N_581,In_415,In_1136);
nor U582 (N_582,In_99,In_649);
or U583 (N_583,In_1962,In_1516);
and U584 (N_584,In_1487,In_143);
xor U585 (N_585,In_1532,In_2282);
nor U586 (N_586,In_666,In_1739);
and U587 (N_587,In_753,In_1209);
and U588 (N_588,In_1610,In_952);
or U589 (N_589,In_455,In_2468);
nor U590 (N_590,In_2296,In_2250);
nor U591 (N_591,In_992,In_1778);
or U592 (N_592,In_1264,In_1721);
nand U593 (N_593,In_1315,In_1864);
nor U594 (N_594,In_1765,In_336);
nand U595 (N_595,In_662,In_673);
and U596 (N_596,In_686,In_885);
and U597 (N_597,In_654,In_432);
or U598 (N_598,In_1349,In_1147);
and U599 (N_599,In_2034,In_1351);
nor U600 (N_600,In_1399,In_213);
or U601 (N_601,In_2195,In_120);
and U602 (N_602,In_2075,In_1352);
nand U603 (N_603,In_1108,In_698);
nor U604 (N_604,In_866,In_2339);
nand U605 (N_605,In_1467,In_1121);
nand U606 (N_606,In_425,In_596);
or U607 (N_607,In_1276,In_1931);
or U608 (N_608,In_440,In_2360);
nor U609 (N_609,In_1393,In_1421);
nand U610 (N_610,In_2207,In_1643);
or U611 (N_611,In_1878,In_325);
nand U612 (N_612,In_133,In_2181);
and U613 (N_613,In_1336,In_1678);
nor U614 (N_614,In_1669,In_825);
nand U615 (N_615,In_1140,In_1504);
or U616 (N_616,In_1766,In_429);
and U617 (N_617,In_1607,In_101);
nor U618 (N_618,In_728,In_704);
and U619 (N_619,In_368,In_2023);
nor U620 (N_620,In_134,In_1007);
nor U621 (N_621,In_1397,In_493);
nor U622 (N_622,In_1983,In_1786);
nor U623 (N_623,In_1185,In_457);
nor U624 (N_624,In_1076,In_1882);
and U625 (N_625,In_1286,In_390);
nor U626 (N_626,In_399,In_164);
and U627 (N_627,In_1097,In_294);
and U628 (N_628,In_541,In_1978);
and U629 (N_629,In_1095,In_1277);
nand U630 (N_630,In_218,In_2088);
and U631 (N_631,In_359,In_777);
nor U632 (N_632,In_2351,In_1946);
and U633 (N_633,In_947,In_1475);
nor U634 (N_634,In_604,In_1799);
and U635 (N_635,In_661,In_142);
or U636 (N_636,In_1149,In_1590);
nor U637 (N_637,In_320,In_2297);
or U638 (N_638,In_2455,In_1434);
and U639 (N_639,In_2238,In_1716);
or U640 (N_640,In_2044,In_572);
and U641 (N_641,In_1417,In_6);
nor U642 (N_642,In_1348,In_592);
nor U643 (N_643,In_621,In_1768);
nor U644 (N_644,In_1344,In_1928);
xor U645 (N_645,In_2324,In_2444);
and U646 (N_646,In_1730,In_451);
nand U647 (N_647,In_1655,In_1498);
and U648 (N_648,In_513,In_503);
nand U649 (N_649,In_2224,In_1081);
nand U650 (N_650,In_1942,In_647);
nor U651 (N_651,In_612,In_2149);
and U652 (N_652,In_1207,In_1287);
nor U653 (N_653,In_1424,In_1390);
and U654 (N_654,In_964,In_2147);
nand U655 (N_655,In_2332,In_681);
nand U656 (N_656,In_282,In_473);
or U657 (N_657,In_1777,In_1204);
or U658 (N_658,In_886,In_1628);
nand U659 (N_659,In_1834,In_1098);
and U660 (N_660,In_2043,In_48);
nand U661 (N_661,In_2072,In_875);
nor U662 (N_662,In_2165,In_640);
xor U663 (N_663,In_2416,In_988);
and U664 (N_664,In_377,In_788);
and U665 (N_665,In_1593,In_1538);
nand U666 (N_666,In_313,In_2243);
or U667 (N_667,In_2216,In_2286);
and U668 (N_668,In_1342,In_2156);
and U669 (N_669,In_1743,In_458);
nor U670 (N_670,In_2057,In_1995);
or U671 (N_671,In_2019,In_110);
and U672 (N_672,In_663,In_1060);
or U673 (N_673,In_1409,In_1569);
and U674 (N_674,In_732,In_28);
nor U675 (N_675,In_1564,In_731);
or U676 (N_676,In_2408,In_2087);
or U677 (N_677,In_1761,In_1325);
or U678 (N_678,In_2494,In_638);
nand U679 (N_679,In_707,In_701);
or U680 (N_680,In_1304,In_2106);
or U681 (N_681,In_858,In_892);
nor U682 (N_682,In_2305,In_231);
or U683 (N_683,In_478,In_2010);
nand U684 (N_684,In_1812,In_2295);
or U685 (N_685,In_873,In_781);
or U686 (N_686,In_2474,In_149);
nor U687 (N_687,In_303,In_12);
nor U688 (N_688,In_1539,In_595);
or U689 (N_689,In_1701,In_2056);
and U690 (N_690,In_1359,In_391);
or U691 (N_691,In_1187,In_529);
xnor U692 (N_692,In_1441,In_872);
or U693 (N_693,In_2404,In_111);
xnor U694 (N_694,In_2187,In_204);
nor U695 (N_695,In_559,In_2245);
or U696 (N_696,In_971,In_1963);
or U697 (N_697,In_1391,In_1955);
nor U698 (N_698,In_593,In_1278);
nand U699 (N_699,In_2443,In_1507);
or U700 (N_700,In_167,In_936);
or U701 (N_701,In_807,In_1179);
nor U702 (N_702,In_2129,In_2460);
or U703 (N_703,In_2312,In_1177);
and U704 (N_704,In_1213,In_47);
and U705 (N_705,In_244,In_2298);
nor U706 (N_706,In_2175,In_1038);
and U707 (N_707,In_2357,In_1661);
and U708 (N_708,In_2433,In_682);
and U709 (N_709,In_1110,In_2445);
nand U710 (N_710,In_1243,In_1848);
or U711 (N_711,In_2126,In_755);
nand U712 (N_712,In_343,In_2204);
nor U713 (N_713,In_1456,In_354);
nand U714 (N_714,In_1086,In_1382);
nor U715 (N_715,In_62,In_1680);
nand U716 (N_716,In_1750,In_2259);
xor U717 (N_717,In_2079,In_1189);
and U718 (N_718,In_2030,In_2217);
nand U719 (N_719,In_42,In_2233);
nor U720 (N_720,In_1886,In_2441);
nor U721 (N_721,In_2384,In_2130);
or U722 (N_722,In_1852,In_1270);
nor U723 (N_723,In_1176,In_345);
or U724 (N_724,In_636,In_1156);
nor U725 (N_725,In_1219,In_1033);
or U726 (N_726,In_859,In_107);
nand U727 (N_727,In_2006,In_260);
nand U728 (N_728,In_689,In_394);
nor U729 (N_729,In_162,In_754);
nor U730 (N_730,In_155,In_1744);
nor U731 (N_731,In_565,In_1773);
nand U732 (N_732,In_852,In_178);
or U733 (N_733,In_463,In_1003);
nand U734 (N_734,In_1432,In_2338);
nor U735 (N_735,In_1116,In_309);
or U736 (N_736,In_1444,In_176);
nand U737 (N_737,In_2486,In_2067);
or U738 (N_738,In_2493,In_2472);
or U739 (N_739,In_59,In_1668);
nand U740 (N_740,In_746,In_236);
nand U741 (N_741,In_1320,In_1965);
nand U742 (N_742,In_1493,In_1230);
nor U743 (N_743,In_1536,In_1485);
or U744 (N_744,In_1662,In_482);
or U745 (N_745,In_2173,In_157);
or U746 (N_746,In_2155,In_509);
nor U747 (N_747,In_1989,In_1929);
xnor U748 (N_748,In_906,In_516);
nand U749 (N_749,In_1014,In_16);
or U750 (N_750,In_970,In_735);
and U751 (N_751,In_1754,In_2160);
nand U752 (N_752,In_2275,In_1499);
or U753 (N_753,In_941,In_2461);
nor U754 (N_754,In_1537,In_416);
or U755 (N_755,In_1006,In_14);
or U756 (N_756,In_2327,In_752);
nor U757 (N_757,In_2119,In_2198);
nor U758 (N_758,In_150,In_1416);
nor U759 (N_759,In_212,In_1462);
nand U760 (N_760,In_2307,In_146);
or U761 (N_761,In_1208,In_1366);
or U762 (N_762,In_829,In_870);
xor U763 (N_763,In_517,In_387);
and U764 (N_764,In_897,In_835);
nand U765 (N_765,In_985,In_1751);
or U766 (N_766,In_1148,In_2400);
or U767 (N_767,In_306,In_446);
and U768 (N_768,In_2425,In_1856);
or U769 (N_769,In_1969,In_1911);
nor U770 (N_770,In_1372,In_2114);
nand U771 (N_771,In_2385,In_2219);
and U772 (N_772,In_1630,In_2398);
or U773 (N_773,In_980,In_126);
and U774 (N_774,In_329,In_2470);
nand U775 (N_775,In_1239,In_1846);
and U776 (N_776,In_2073,In_1690);
and U777 (N_777,In_1709,In_1112);
or U778 (N_778,In_720,In_1706);
nor U779 (N_779,In_1927,In_414);
nand U780 (N_780,In_1872,In_1992);
or U781 (N_781,In_721,In_1083);
nand U782 (N_782,In_1309,In_1543);
or U783 (N_783,In_1868,In_1423);
nor U784 (N_784,In_27,In_1895);
nand U785 (N_785,In_2133,In_639);
nor U786 (N_786,In_652,In_2449);
and U787 (N_787,In_1704,In_655);
nor U788 (N_788,In_2394,In_1663);
nand U789 (N_789,In_2321,In_1506);
nand U790 (N_790,In_1994,In_1466);
and U791 (N_791,In_1183,In_2009);
or U792 (N_792,In_597,In_1876);
or U793 (N_793,In_1193,In_1017);
and U794 (N_794,In_928,In_1150);
and U795 (N_795,In_2211,In_2380);
nor U796 (N_796,In_1031,In_724);
nor U797 (N_797,In_1735,In_1281);
and U798 (N_798,In_113,In_484);
nand U799 (N_799,In_1691,In_847);
and U800 (N_800,In_945,In_1254);
and U801 (N_801,In_1981,In_90);
nor U802 (N_802,In_395,In_1195);
or U803 (N_803,In_45,In_569);
nor U804 (N_804,In_1132,In_1356);
xnor U805 (N_805,In_227,In_845);
or U806 (N_806,In_402,In_93);
and U807 (N_807,In_1804,In_2100);
nor U808 (N_808,In_2083,In_1842);
or U809 (N_809,In_1687,In_2068);
and U810 (N_810,In_1075,In_180);
nand U811 (N_811,In_2403,In_1070);
nor U812 (N_812,In_1492,In_2264);
nor U813 (N_813,In_2272,In_245);
nand U814 (N_814,In_485,In_1637);
and U815 (N_815,In_321,In_2054);
or U816 (N_816,In_1412,In_1822);
nor U817 (N_817,In_2162,In_355);
and U818 (N_818,In_2463,In_1993);
and U819 (N_819,In_411,In_793);
nand U820 (N_820,In_2110,In_323);
and U821 (N_821,In_152,In_1699);
and U822 (N_822,In_1009,In_1395);
nand U823 (N_823,In_1567,In_1043);
or U824 (N_824,In_1251,In_1523);
or U825 (N_825,In_850,In_1253);
and U826 (N_826,In_1465,In_96);
nor U827 (N_827,In_1260,In_1387);
or U828 (N_828,In_1357,In_172);
and U829 (N_829,In_702,In_2409);
or U830 (N_830,In_1223,In_1222);
and U831 (N_831,In_502,In_1134);
nand U832 (N_832,In_1353,In_1418);
or U833 (N_833,In_530,In_2371);
nand U834 (N_834,In_1322,In_2412);
xor U835 (N_835,In_1063,In_1530);
nand U836 (N_836,In_2125,In_1675);
nand U837 (N_837,In_249,In_2373);
and U838 (N_838,In_474,In_2457);
and U839 (N_839,In_923,In_360);
and U840 (N_840,In_1714,In_1473);
nand U841 (N_841,In_830,In_35);
or U842 (N_842,In_1926,In_1069);
and U843 (N_843,In_1064,In_91);
or U844 (N_844,In_842,In_658);
nor U845 (N_845,In_1790,In_2003);
and U846 (N_846,In_1072,In_2490);
nor U847 (N_847,In_350,In_2152);
and U848 (N_848,In_2093,In_2246);
and U849 (N_849,In_1266,In_1723);
and U850 (N_850,In_1285,In_924);
nand U851 (N_851,In_644,In_1271);
or U852 (N_852,In_1419,In_64);
and U853 (N_853,In_534,In_611);
and U854 (N_854,In_1169,In_1002);
or U855 (N_855,In_17,In_840);
nand U856 (N_856,In_2364,In_542);
nor U857 (N_857,In_1854,In_1221);
or U858 (N_858,In_2105,In_742);
nor U859 (N_859,In_1273,In_199);
nand U860 (N_860,In_1331,In_92);
xor U861 (N_861,In_1597,In_1867);
and U862 (N_862,In_535,In_304);
nand U863 (N_863,In_1903,In_1073);
nor U864 (N_864,In_641,In_2042);
and U865 (N_865,In_2372,In_2362);
nand U866 (N_866,In_2309,In_1046);
nand U867 (N_867,In_533,In_1708);
or U868 (N_868,In_719,In_600);
xnor U869 (N_869,In_2239,In_994);
or U870 (N_870,In_131,In_2060);
or U871 (N_871,In_1042,In_553);
or U872 (N_872,In_1990,In_1451);
and U873 (N_873,In_1225,In_369);
nor U874 (N_874,In_2090,In_37);
and U875 (N_875,In_1546,In_1794);
and U876 (N_876,In_1674,In_284);
nor U877 (N_877,In_340,In_1371);
or U878 (N_878,In_168,In_1559);
or U879 (N_879,In_632,In_235);
or U880 (N_880,In_1938,In_786);
or U881 (N_881,In_192,In_2014);
and U882 (N_882,In_973,In_854);
or U883 (N_883,In_1477,In_217);
and U884 (N_884,In_761,In_1054);
nor U885 (N_885,In_2368,In_1772);
and U886 (N_886,In_2355,In_792);
nor U887 (N_887,In_2048,In_774);
nor U888 (N_888,In_1957,In_1540);
nand U889 (N_889,In_1801,In_2496);
and U890 (N_890,In_1879,In_2320);
or U891 (N_891,In_1403,In_1155);
nor U892 (N_892,In_252,In_226);
nor U893 (N_893,In_1887,In_237);
and U894 (N_894,In_436,In_314);
nor U895 (N_895,In_349,In_1617);
and U896 (N_896,In_2001,In_1109);
or U897 (N_897,In_2347,In_1763);
or U898 (N_898,In_286,In_1052);
and U899 (N_899,In_1427,In_1529);
xnor U900 (N_900,In_528,In_15);
or U901 (N_901,In_2231,In_1819);
nor U902 (N_902,In_337,In_2096);
nor U903 (N_903,In_841,In_364);
nor U904 (N_904,In_1636,In_1431);
nor U905 (N_905,In_522,In_738);
or U906 (N_906,In_1816,In_605);
and U907 (N_907,In_1935,In_756);
or U908 (N_908,In_910,In_1171);
or U909 (N_909,In_1845,In_102);
or U910 (N_910,In_371,In_1634);
or U911 (N_911,In_229,In_2318);
or U912 (N_912,In_2325,In_844);
and U913 (N_913,In_987,In_912);
and U914 (N_914,In_1288,In_613);
and U915 (N_915,In_630,In_1048);
nand U916 (N_916,In_691,In_159);
xnor U917 (N_917,In_288,In_1471);
or U918 (N_918,In_575,In_1401);
nor U919 (N_919,In_1966,In_1292);
and U920 (N_920,In_2283,In_2390);
nor U921 (N_921,In_2032,In_1698);
nand U922 (N_922,In_1589,In_1024);
nand U923 (N_923,In_341,In_2422);
nor U924 (N_924,In_560,In_1646);
and U925 (N_925,In_1101,In_1463);
nor U926 (N_926,In_2254,In_1298);
nor U927 (N_927,In_623,In_208);
nor U928 (N_928,In_1084,In_333);
or U929 (N_929,In_819,In_656);
xor U930 (N_930,In_69,In_749);
and U931 (N_931,In_2328,In_1719);
and U932 (N_932,In_668,In_308);
xnor U933 (N_933,In_88,In_246);
xnor U934 (N_934,In_1153,In_653);
and U935 (N_935,In_1578,In_2483);
or U936 (N_936,In_562,In_1092);
or U937 (N_937,In_2401,In_1633);
nand U938 (N_938,In_1358,In_2349);
or U939 (N_939,In_972,In_1606);
or U940 (N_940,In_599,In_1588);
and U941 (N_941,In_2045,In_2144);
nand U942 (N_942,In_1154,In_1554);
nor U943 (N_943,In_2478,In_1956);
nand U944 (N_944,In_1859,In_2183);
nand U945 (N_945,In_1392,In_1044);
nor U946 (N_946,In_276,In_94);
and U947 (N_947,In_794,In_228);
or U948 (N_948,In_615,In_1491);
nand U949 (N_949,In_684,In_816);
nor U950 (N_950,In_215,In_197);
nor U951 (N_951,In_1138,In_1986);
nor U952 (N_952,In_1004,In_631);
nand U953 (N_953,In_1053,In_1234);
nand U954 (N_954,In_1695,In_1839);
and U955 (N_955,In_1157,In_2370);
or U956 (N_956,In_713,In_255);
nor U957 (N_957,In_2499,In_1660);
nor U958 (N_958,In_2104,In_2407);
and U959 (N_959,In_911,In_904);
nand U960 (N_960,In_1199,In_1725);
nor U961 (N_961,In_1600,In_1742);
nor U962 (N_962,In_2192,In_551);
nand U963 (N_963,In_121,In_1654);
xor U964 (N_964,In_220,In_2059);
nand U965 (N_965,In_1474,In_717);
nand U966 (N_966,In_58,In_2212);
nor U967 (N_967,In_2482,In_1549);
nand U968 (N_968,In_577,In_993);
nor U969 (N_969,In_2306,In_148);
or U970 (N_970,In_1534,In_2139);
nor U971 (N_971,In_444,In_1676);
and U972 (N_972,In_1941,In_1869);
nor U973 (N_973,In_1250,In_1923);
nand U974 (N_974,In_815,In_2256);
and U975 (N_975,In_554,In_2428);
and U976 (N_976,In_1601,In_1130);
or U977 (N_977,In_2375,In_2148);
and U978 (N_978,In_2453,In_2358);
or U979 (N_979,In_2294,In_420);
or U980 (N_980,In_857,In_1808);
nand U981 (N_981,In_1985,In_1781);
and U982 (N_982,In_802,In_1968);
nor U983 (N_983,In_2498,In_1722);
nand U984 (N_984,In_1410,In_1939);
or U985 (N_985,In_41,In_9);
nor U986 (N_986,In_1806,In_274);
or U987 (N_987,In_2074,In_1196);
nor U988 (N_988,In_1297,In_1468);
nand U989 (N_989,In_2480,In_1478);
nand U990 (N_990,In_1697,In_862);
and U991 (N_991,In_2374,In_2161);
nor U992 (N_992,In_1012,In_2273);
or U993 (N_993,In_63,In_2230);
nor U994 (N_994,In_2326,In_531);
nand U995 (N_995,In_856,In_86);
nand U996 (N_996,In_1407,In_1855);
xnor U997 (N_997,In_52,In_1106);
nor U998 (N_998,In_2017,In_1563);
nor U999 (N_999,In_1519,In_25);
nand U1000 (N_1000,In_1613,In_1381);
nor U1001 (N_1001,In_211,In_617);
nand U1002 (N_1002,In_1807,In_2244);
and U1003 (N_1003,In_536,In_1782);
nor U1004 (N_1004,In_1948,In_1036);
nor U1005 (N_1005,In_2292,In_18);
or U1006 (N_1006,In_1641,In_1889);
or U1007 (N_1007,In_1317,In_2304);
nand U1008 (N_1008,In_979,In_1389);
and U1009 (N_1009,In_1796,In_68);
nand U1010 (N_1010,In_860,In_293);
or U1011 (N_1011,In_1631,In_264);
xor U1012 (N_1012,In_2052,In_984);
nand U1013 (N_1013,In_523,In_1638);
and U1014 (N_1014,In_776,In_430);
nand U1015 (N_1015,In_1827,In_1090);
or U1016 (N_1016,In_2228,In_1433);
nor U1017 (N_1017,In_950,In_1057);
or U1018 (N_1018,In_43,In_1192);
and U1019 (N_1019,In_930,In_224);
nor U1020 (N_1020,In_963,In_105);
xor U1021 (N_1021,In_311,In_1000);
and U1022 (N_1022,In_1755,In_2170);
and U1023 (N_1023,In_922,In_1124);
and U1024 (N_1024,In_1323,In_1626);
or U1025 (N_1025,In_557,In_909);
nor U1026 (N_1026,In_828,In_1450);
nor U1027 (N_1027,In_725,In_1360);
xnor U1028 (N_1028,In_2378,In_1020);
xor U1029 (N_1029,In_587,In_1553);
or U1030 (N_1030,In_2310,In_1917);
and U1031 (N_1031,In_2391,In_67);
nor U1032 (N_1032,In_44,In_1296);
and U1033 (N_1033,In_206,In_814);
nand U1034 (N_1034,In_1517,In_322);
or U1035 (N_1035,In_2476,In_918);
and U1036 (N_1036,In_550,In_2167);
nand U1037 (N_1037,In_1671,In_1591);
and U1038 (N_1038,In_675,In_589);
or U1039 (N_1039,In_2247,In_1103);
nand U1040 (N_1040,In_1291,In_1248);
or U1041 (N_1041,In_1301,In_60);
nand U1042 (N_1042,In_190,In_2266);
nor U1043 (N_1043,In_406,In_932);
or U1044 (N_1044,In_1120,In_381);
nand U1045 (N_1045,In_552,In_958);
or U1046 (N_1046,In_2112,In_1247);
and U1047 (N_1047,In_1307,In_1511);
and U1048 (N_1048,In_1640,In_296);
nor U1049 (N_1049,In_2267,In_563);
nor U1050 (N_1050,In_2029,In_189);
nand U1051 (N_1051,In_1598,In_946);
or U1052 (N_1052,In_2174,In_1683);
or U1053 (N_1053,In_339,In_622);
nor U1054 (N_1054,In_740,In_1959);
xor U1055 (N_1055,In_283,In_891);
and U1056 (N_1056,In_1837,In_1363);
nand U1057 (N_1057,In_2454,In_1319);
nand U1058 (N_1058,In_1653,In_1131);
nand U1059 (N_1059,In_2271,In_1126);
nor U1060 (N_1060,In_397,In_338);
and U1061 (N_1061,In_165,In_1665);
nand U1062 (N_1062,In_545,In_2166);
or U1063 (N_1063,In_2210,In_2316);
and U1064 (N_1064,In_960,In_1921);
and U1065 (N_1065,In_679,In_500);
nand U1066 (N_1066,In_1454,In_1776);
or U1067 (N_1067,In_1128,In_585);
nand U1068 (N_1068,In_901,In_285);
or U1069 (N_1069,In_1367,In_547);
or U1070 (N_1070,In_659,In_1970);
and U1071 (N_1071,In_2253,In_2012);
and U1072 (N_1072,In_1368,In_1429);
and U1073 (N_1073,In_443,In_532);
nor U1074 (N_1074,In_2299,In_846);
and U1075 (N_1075,In_1542,In_2078);
nand U1076 (N_1076,In_574,In_1457);
nand U1077 (N_1077,In_975,In_2200);
or U1078 (N_1078,In_2095,In_1096);
nand U1079 (N_1079,In_2103,In_1828);
or U1080 (N_1080,In_1232,In_2367);
and U1081 (N_1081,In_1481,In_1575);
nor U1082 (N_1082,In_688,In_1217);
nand U1083 (N_1083,In_1579,In_1490);
nor U1084 (N_1084,In_771,In_2382);
or U1085 (N_1085,In_428,In_2258);
and U1086 (N_1086,In_401,In_372);
and U1087 (N_1087,In_2365,In_119);
or U1088 (N_1088,In_757,In_1740);
and U1089 (N_1089,In_1595,In_1930);
or U1090 (N_1090,In_2393,In_1343);
nor U1091 (N_1091,In_1826,In_1657);
or U1092 (N_1092,In_54,In_1860);
and U1093 (N_1093,In_97,In_899);
and U1094 (N_1094,In_106,In_1577);
and U1095 (N_1095,In_791,In_878);
nor U1096 (N_1096,In_2397,In_642);
nand U1097 (N_1097,In_1915,In_1339);
or U1098 (N_1098,In_1571,In_2379);
nand U1099 (N_1099,In_424,In_1347);
or U1100 (N_1100,In_98,In_1246);
nor U1101 (N_1101,In_2345,In_361);
nand U1102 (N_1102,In_1748,In_1265);
or U1103 (N_1103,In_300,In_2202);
nor U1104 (N_1104,In_2,In_1545);
and U1105 (N_1105,In_1746,In_2300);
and U1106 (N_1106,In_1836,In_365);
nor U1107 (N_1107,In_620,In_2363);
and U1108 (N_1108,In_1016,In_1984);
or U1109 (N_1109,In_775,In_568);
or U1110 (N_1110,In_1374,In_472);
or U1111 (N_1111,In_1833,In_2330);
nor U1112 (N_1112,In_76,In_1146);
nor U1113 (N_1113,In_672,In_907);
and U1114 (N_1114,In_382,In_1430);
or U1115 (N_1115,In_2071,In_959);
and U1116 (N_1116,In_508,In_1159);
or U1117 (N_1117,In_1973,In_1210);
nand U1118 (N_1118,In_1509,In_422);
or U1119 (N_1119,In_1476,In_1242);
nand U1120 (N_1120,In_751,In_1913);
or U1121 (N_1121,In_2414,In_1314);
nand U1122 (N_1122,In_1515,In_73);
nand U1123 (N_1123,In_665,In_334);
nand U1124 (N_1124,In_419,In_1738);
and U1125 (N_1125,In_1205,In_230);
nand U1126 (N_1126,In_1028,In_1821);
and U1127 (N_1127,In_2002,In_504);
and U1128 (N_1128,In_2432,In_201);
nor U1129 (N_1129,In_501,In_764);
nand U1130 (N_1130,In_2442,In_1731);
nand U1131 (N_1131,In_1045,In_281);
nor U1132 (N_1132,In_46,In_1469);
or U1133 (N_1133,In_117,In_1074);
nand U1134 (N_1134,In_1920,In_822);
and U1135 (N_1135,In_2484,In_1218);
nand U1136 (N_1136,In_413,In_481);
nor U1137 (N_1137,In_1724,In_1104);
nand U1138 (N_1138,In_1525,In_1762);
or U1139 (N_1139,In_1584,In_2000);
and U1140 (N_1140,In_1279,In_999);
and U1141 (N_1141,In_1693,In_95);
nor U1142 (N_1142,In_2413,In_1905);
nor U1143 (N_1143,In_2182,In_1971);
or U1144 (N_1144,In_573,In_709);
and U1145 (N_1145,In_2176,In_2179);
nand U1146 (N_1146,In_1400,In_433);
or U1147 (N_1147,In_187,In_2055);
and U1148 (N_1148,In_2206,In_2018);
and U1149 (N_1149,In_263,In_1527);
and U1150 (N_1150,In_1759,In_671);
nor U1151 (N_1151,In_2276,In_1877);
or U1152 (N_1152,In_2051,In_1172);
nor U1153 (N_1153,In_1629,In_169);
nand U1154 (N_1154,In_2151,In_2169);
and U1155 (N_1155,In_1940,In_594);
nand U1156 (N_1156,In_2249,In_84);
nor U1157 (N_1157,In_1376,In_1627);
nor U1158 (N_1158,In_637,In_454);
nor U1159 (N_1159,In_1066,In_869);
nor U1160 (N_1160,In_920,In_1720);
and U1161 (N_1161,In_521,In_1026);
nand U1162 (N_1162,In_927,In_1068);
or U1163 (N_1163,In_181,In_1862);
and U1164 (N_1164,In_715,In_385);
nand U1165 (N_1165,In_1784,In_442);
and U1166 (N_1166,In_582,In_1047);
or U1167 (N_1167,In_1573,In_2377);
nand U1168 (N_1168,In_2285,In_153);
nor U1169 (N_1169,In_34,In_2479);
and U1170 (N_1170,In_327,In_1373);
and U1171 (N_1171,In_1729,In_2203);
or U1172 (N_1172,In_2376,In_1472);
nand U1173 (N_1173,In_1226,In_711);
nor U1174 (N_1174,In_1944,In_1518);
xor U1175 (N_1175,In_1619,In_1378);
and U1176 (N_1176,In_838,In_373);
nor U1177 (N_1177,In_1340,In_2456);
and U1178 (N_1178,In_2291,In_843);
or U1179 (N_1179,In_750,In_421);
nand U1180 (N_1180,In_1541,In_470);
nor U1181 (N_1181,In_1943,In_2410);
or U1182 (N_1182,In_748,In_1635);
or U1183 (N_1183,In_810,In_2146);
and U1184 (N_1184,In_555,In_619);
nand U1185 (N_1185,In_1922,In_2411);
nand U1186 (N_1186,In_2335,In_1328);
or U1187 (N_1187,In_262,In_468);
nand U1188 (N_1188,In_2229,In_175);
nor U1189 (N_1189,In_1904,In_1576);
or U1190 (N_1190,In_1603,In_2223);
nand U1191 (N_1191,In_2196,In_118);
or U1192 (N_1192,In_712,In_477);
and U1193 (N_1193,In_1118,In_147);
and U1194 (N_1194,In_1503,In_744);
nand U1195 (N_1195,In_85,In_2424);
nor U1196 (N_1196,In_1458,In_2356);
nand U1197 (N_1197,In_2323,In_1055);
and U1198 (N_1198,In_2301,In_1997);
nand U1199 (N_1199,In_690,In_1170);
or U1200 (N_1200,In_730,In_1437);
and U1201 (N_1201,In_2194,In_1520);
nor U1202 (N_1202,In_2288,In_955);
or U1203 (N_1203,In_1684,In_205);
or U1204 (N_1204,In_1972,In_376);
or U1205 (N_1205,In_1558,In_138);
nand U1206 (N_1206,In_1936,In_100);
nand U1207 (N_1207,In_961,In_643);
nand U1208 (N_1208,In_366,In_2027);
and U1209 (N_1209,In_1311,In_20);
and U1210 (N_1210,In_291,In_902);
or U1211 (N_1211,In_1091,In_765);
nor U1212 (N_1212,In_2387,In_1505);
and U1213 (N_1213,In_2226,In_566);
and U1214 (N_1214,In_635,In_1552);
xor U1215 (N_1215,In_1871,In_1127);
or U1216 (N_1216,In_1582,In_2015);
or U1217 (N_1217,In_538,In_129);
or U1218 (N_1218,In_1280,In_1551);
nor U1219 (N_1219,In_1919,In_2185);
nor U1220 (N_1220,In_809,In_65);
nand U1221 (N_1221,In_1425,In_1117);
and U1222 (N_1222,In_1502,In_26);
nor U1223 (N_1223,In_974,In_2350);
or U1224 (N_1224,In_747,In_1094);
nor U1225 (N_1225,In_676,In_579);
or U1226 (N_1226,In_1184,In_19);
nor U1227 (N_1227,In_210,In_480);
nor U1228 (N_1228,In_247,In_606);
and U1229 (N_1229,In_1547,In_1058);
or U1230 (N_1230,In_1658,In_2446);
xnor U1231 (N_1231,In_1386,In_2220);
nor U1232 (N_1232,In_1143,In_352);
or U1233 (N_1233,In_2405,In_699);
and U1234 (N_1234,In_944,In_685);
nand U1235 (N_1235,In_1145,In_570);
nor U1236 (N_1236,In_173,In_271);
xor U1237 (N_1237,In_2036,In_2473);
or U1238 (N_1238,In_145,In_450);
xor U1239 (N_1239,In_729,In_222);
and U1240 (N_1240,In_1290,In_2040);
nor U1241 (N_1241,In_1249,In_1838);
and U1242 (N_1242,In_1884,In_2142);
xnor U1243 (N_1243,In_1188,In_66);
and U1244 (N_1244,In_1548,In_1951);
or U1245 (N_1245,In_2077,In_626);
or U1246 (N_1246,In_1770,In_1779);
and U1247 (N_1247,In_882,In_2293);
or U1248 (N_1248,In_1960,In_2426);
or U1249 (N_1249,In_491,In_2108);
nor U1250 (N_1250,In_1088,In_306);
or U1251 (N_1251,In_903,In_1402);
or U1252 (N_1252,In_755,In_331);
nor U1253 (N_1253,In_1985,In_2418);
nand U1254 (N_1254,In_2369,In_1357);
nor U1255 (N_1255,In_2254,In_991);
nor U1256 (N_1256,In_858,In_1090);
or U1257 (N_1257,In_296,In_1380);
or U1258 (N_1258,In_2133,In_2385);
nor U1259 (N_1259,In_2271,In_1257);
and U1260 (N_1260,In_480,In_912);
nor U1261 (N_1261,In_1966,In_1906);
and U1262 (N_1262,In_1435,In_1327);
nand U1263 (N_1263,In_1772,In_1184);
xor U1264 (N_1264,In_615,In_1518);
nand U1265 (N_1265,In_222,In_2453);
and U1266 (N_1266,In_2216,In_2096);
nand U1267 (N_1267,In_891,In_27);
nand U1268 (N_1268,In_1770,In_1982);
nand U1269 (N_1269,In_1450,In_2251);
nand U1270 (N_1270,In_604,In_2034);
and U1271 (N_1271,In_864,In_1206);
or U1272 (N_1272,In_582,In_617);
nor U1273 (N_1273,In_1648,In_1782);
or U1274 (N_1274,In_1167,In_1257);
and U1275 (N_1275,In_332,In_1827);
xnor U1276 (N_1276,In_950,In_386);
xor U1277 (N_1277,In_828,In_2024);
and U1278 (N_1278,In_2285,In_1945);
or U1279 (N_1279,In_353,In_1594);
nor U1280 (N_1280,In_309,In_641);
and U1281 (N_1281,In_36,In_1328);
and U1282 (N_1282,In_748,In_327);
nand U1283 (N_1283,In_2465,In_559);
nor U1284 (N_1284,In_490,In_905);
nor U1285 (N_1285,In_2235,In_416);
nand U1286 (N_1286,In_1640,In_954);
nand U1287 (N_1287,In_1960,In_983);
and U1288 (N_1288,In_874,In_1597);
and U1289 (N_1289,In_1226,In_2204);
and U1290 (N_1290,In_584,In_2434);
and U1291 (N_1291,In_683,In_364);
and U1292 (N_1292,In_1247,In_1126);
nor U1293 (N_1293,In_837,In_288);
nand U1294 (N_1294,In_1194,In_958);
nand U1295 (N_1295,In_810,In_905);
or U1296 (N_1296,In_2292,In_495);
or U1297 (N_1297,In_293,In_690);
nand U1298 (N_1298,In_1573,In_1131);
nor U1299 (N_1299,In_252,In_1155);
and U1300 (N_1300,In_1028,In_490);
or U1301 (N_1301,In_507,In_2265);
nand U1302 (N_1302,In_1968,In_974);
nand U1303 (N_1303,In_276,In_679);
and U1304 (N_1304,In_1139,In_516);
nor U1305 (N_1305,In_2386,In_488);
nor U1306 (N_1306,In_528,In_529);
or U1307 (N_1307,In_46,In_1117);
and U1308 (N_1308,In_1691,In_441);
nor U1309 (N_1309,In_200,In_1578);
nand U1310 (N_1310,In_1367,In_1197);
or U1311 (N_1311,In_678,In_1038);
nand U1312 (N_1312,In_600,In_1948);
or U1313 (N_1313,In_1593,In_156);
and U1314 (N_1314,In_1822,In_2487);
nand U1315 (N_1315,In_1273,In_861);
nor U1316 (N_1316,In_894,In_2324);
xor U1317 (N_1317,In_2466,In_2494);
nor U1318 (N_1318,In_1416,In_1700);
xnor U1319 (N_1319,In_2331,In_1442);
nand U1320 (N_1320,In_181,In_2156);
nand U1321 (N_1321,In_1361,In_1442);
and U1322 (N_1322,In_1129,In_274);
and U1323 (N_1323,In_132,In_1510);
and U1324 (N_1324,In_1683,In_194);
nand U1325 (N_1325,In_366,In_1058);
and U1326 (N_1326,In_538,In_243);
and U1327 (N_1327,In_1341,In_1543);
or U1328 (N_1328,In_1268,In_694);
nor U1329 (N_1329,In_938,In_1346);
and U1330 (N_1330,In_1825,In_1694);
or U1331 (N_1331,In_201,In_449);
nor U1332 (N_1332,In_135,In_347);
nor U1333 (N_1333,In_944,In_1492);
xor U1334 (N_1334,In_1499,In_601);
nand U1335 (N_1335,In_649,In_2300);
or U1336 (N_1336,In_1079,In_2127);
or U1337 (N_1337,In_984,In_1833);
nand U1338 (N_1338,In_10,In_1646);
nor U1339 (N_1339,In_2213,In_1040);
or U1340 (N_1340,In_664,In_545);
nor U1341 (N_1341,In_305,In_1604);
nor U1342 (N_1342,In_1482,In_1434);
and U1343 (N_1343,In_1778,In_708);
xor U1344 (N_1344,In_1948,In_2315);
or U1345 (N_1345,In_1892,In_23);
nor U1346 (N_1346,In_1919,In_1745);
xor U1347 (N_1347,In_1286,In_568);
or U1348 (N_1348,In_712,In_524);
and U1349 (N_1349,In_1749,In_585);
nand U1350 (N_1350,In_1374,In_1881);
nor U1351 (N_1351,In_1321,In_227);
nand U1352 (N_1352,In_1618,In_227);
nand U1353 (N_1353,In_2467,In_1820);
and U1354 (N_1354,In_893,In_2096);
or U1355 (N_1355,In_1833,In_100);
or U1356 (N_1356,In_1300,In_59);
xor U1357 (N_1357,In_1395,In_1340);
or U1358 (N_1358,In_430,In_2056);
nand U1359 (N_1359,In_575,In_31);
and U1360 (N_1360,In_1825,In_251);
or U1361 (N_1361,In_1592,In_830);
or U1362 (N_1362,In_1410,In_358);
nand U1363 (N_1363,In_1265,In_41);
and U1364 (N_1364,In_1883,In_1202);
nand U1365 (N_1365,In_2395,In_1779);
nand U1366 (N_1366,In_1228,In_1933);
xnor U1367 (N_1367,In_2079,In_47);
or U1368 (N_1368,In_673,In_1670);
or U1369 (N_1369,In_2207,In_1902);
nor U1370 (N_1370,In_1055,In_846);
nand U1371 (N_1371,In_1903,In_1741);
and U1372 (N_1372,In_262,In_2171);
nor U1373 (N_1373,In_2125,In_1916);
and U1374 (N_1374,In_2149,In_822);
nand U1375 (N_1375,In_708,In_907);
and U1376 (N_1376,In_461,In_1348);
or U1377 (N_1377,In_1978,In_32);
nand U1378 (N_1378,In_2230,In_547);
nor U1379 (N_1379,In_1192,In_1049);
nor U1380 (N_1380,In_1113,In_949);
nor U1381 (N_1381,In_1975,In_2332);
nor U1382 (N_1382,In_1058,In_1729);
nand U1383 (N_1383,In_1306,In_1699);
and U1384 (N_1384,In_1199,In_550);
and U1385 (N_1385,In_744,In_676);
nor U1386 (N_1386,In_1837,In_641);
and U1387 (N_1387,In_959,In_1883);
and U1388 (N_1388,In_1729,In_1823);
nand U1389 (N_1389,In_2438,In_2098);
nor U1390 (N_1390,In_26,In_516);
nor U1391 (N_1391,In_1066,In_376);
and U1392 (N_1392,In_1155,In_2401);
nand U1393 (N_1393,In_1342,In_1623);
and U1394 (N_1394,In_2340,In_261);
or U1395 (N_1395,In_1876,In_830);
nor U1396 (N_1396,In_21,In_1518);
or U1397 (N_1397,In_479,In_2345);
and U1398 (N_1398,In_108,In_1477);
and U1399 (N_1399,In_1486,In_73);
nand U1400 (N_1400,In_2374,In_1782);
and U1401 (N_1401,In_1774,In_1386);
nor U1402 (N_1402,In_1604,In_1412);
and U1403 (N_1403,In_1115,In_1662);
nand U1404 (N_1404,In_370,In_1124);
or U1405 (N_1405,In_1743,In_1610);
nor U1406 (N_1406,In_198,In_924);
or U1407 (N_1407,In_610,In_801);
and U1408 (N_1408,In_778,In_2211);
nor U1409 (N_1409,In_2130,In_1575);
nand U1410 (N_1410,In_1835,In_2014);
or U1411 (N_1411,In_308,In_2418);
nand U1412 (N_1412,In_240,In_657);
nand U1413 (N_1413,In_584,In_1158);
xor U1414 (N_1414,In_1907,In_2296);
or U1415 (N_1415,In_1439,In_1493);
xnor U1416 (N_1416,In_1745,In_614);
nor U1417 (N_1417,In_743,In_442);
nand U1418 (N_1418,In_394,In_339);
or U1419 (N_1419,In_2317,In_2015);
or U1420 (N_1420,In_1401,In_1626);
or U1421 (N_1421,In_121,In_1738);
and U1422 (N_1422,In_767,In_1945);
nand U1423 (N_1423,In_26,In_1639);
nor U1424 (N_1424,In_390,In_138);
nor U1425 (N_1425,In_2372,In_510);
nand U1426 (N_1426,In_692,In_823);
nand U1427 (N_1427,In_1853,In_1078);
and U1428 (N_1428,In_1887,In_54);
and U1429 (N_1429,In_1952,In_1407);
nor U1430 (N_1430,In_2370,In_1021);
nor U1431 (N_1431,In_1135,In_348);
and U1432 (N_1432,In_459,In_69);
and U1433 (N_1433,In_1489,In_495);
and U1434 (N_1434,In_1984,In_1337);
and U1435 (N_1435,In_195,In_837);
nor U1436 (N_1436,In_2353,In_1695);
or U1437 (N_1437,In_825,In_972);
and U1438 (N_1438,In_2441,In_1746);
nand U1439 (N_1439,In_613,In_1823);
and U1440 (N_1440,In_665,In_1009);
nand U1441 (N_1441,In_938,In_2296);
nand U1442 (N_1442,In_412,In_2423);
and U1443 (N_1443,In_325,In_2241);
nand U1444 (N_1444,In_2138,In_2000);
and U1445 (N_1445,In_1831,In_139);
nor U1446 (N_1446,In_2080,In_2346);
or U1447 (N_1447,In_1858,In_680);
xor U1448 (N_1448,In_242,In_893);
and U1449 (N_1449,In_1854,In_1432);
and U1450 (N_1450,In_813,In_1075);
nor U1451 (N_1451,In_2230,In_398);
and U1452 (N_1452,In_537,In_597);
and U1453 (N_1453,In_475,In_1682);
and U1454 (N_1454,In_1332,In_1568);
nand U1455 (N_1455,In_2275,In_742);
nand U1456 (N_1456,In_1492,In_1439);
and U1457 (N_1457,In_734,In_910);
nor U1458 (N_1458,In_182,In_2165);
nand U1459 (N_1459,In_319,In_251);
nor U1460 (N_1460,In_847,In_1796);
or U1461 (N_1461,In_169,In_373);
and U1462 (N_1462,In_424,In_2256);
or U1463 (N_1463,In_1816,In_643);
nor U1464 (N_1464,In_513,In_1897);
and U1465 (N_1465,In_1459,In_2143);
or U1466 (N_1466,In_50,In_2322);
nor U1467 (N_1467,In_1128,In_304);
xor U1468 (N_1468,In_2398,In_1299);
and U1469 (N_1469,In_2019,In_1961);
or U1470 (N_1470,In_1656,In_566);
nor U1471 (N_1471,In_1452,In_2254);
nor U1472 (N_1472,In_2261,In_1208);
or U1473 (N_1473,In_1474,In_2334);
nand U1474 (N_1474,In_2176,In_404);
or U1475 (N_1475,In_1617,In_108);
nand U1476 (N_1476,In_1341,In_2330);
or U1477 (N_1477,In_469,In_47);
or U1478 (N_1478,In_2188,In_2409);
nor U1479 (N_1479,In_1000,In_156);
or U1480 (N_1480,In_304,In_1983);
or U1481 (N_1481,In_1894,In_60);
and U1482 (N_1482,In_38,In_1036);
or U1483 (N_1483,In_1017,In_1504);
nor U1484 (N_1484,In_2204,In_1937);
nand U1485 (N_1485,In_1755,In_339);
nor U1486 (N_1486,In_1629,In_1224);
nand U1487 (N_1487,In_826,In_1713);
nand U1488 (N_1488,In_1932,In_573);
and U1489 (N_1489,In_898,In_1406);
nand U1490 (N_1490,In_1578,In_1317);
nand U1491 (N_1491,In_138,In_698);
nor U1492 (N_1492,In_2264,In_1933);
nand U1493 (N_1493,In_1314,In_2329);
nand U1494 (N_1494,In_1297,In_1458);
nor U1495 (N_1495,In_861,In_544);
nand U1496 (N_1496,In_784,In_349);
or U1497 (N_1497,In_1045,In_927);
xor U1498 (N_1498,In_445,In_1887);
or U1499 (N_1499,In_1179,In_1330);
nand U1500 (N_1500,In_1014,In_2023);
nand U1501 (N_1501,In_403,In_51);
nor U1502 (N_1502,In_2072,In_652);
and U1503 (N_1503,In_998,In_2068);
nand U1504 (N_1504,In_1829,In_164);
nor U1505 (N_1505,In_1268,In_582);
nor U1506 (N_1506,In_424,In_381);
and U1507 (N_1507,In_1595,In_771);
nor U1508 (N_1508,In_1896,In_1042);
and U1509 (N_1509,In_1864,In_1321);
nand U1510 (N_1510,In_405,In_2043);
nand U1511 (N_1511,In_50,In_1831);
and U1512 (N_1512,In_348,In_2223);
or U1513 (N_1513,In_1235,In_209);
and U1514 (N_1514,In_405,In_2203);
or U1515 (N_1515,In_1391,In_815);
and U1516 (N_1516,In_1658,In_437);
nor U1517 (N_1517,In_1050,In_840);
nor U1518 (N_1518,In_651,In_142);
or U1519 (N_1519,In_526,In_725);
nor U1520 (N_1520,In_2246,In_1044);
or U1521 (N_1521,In_310,In_243);
or U1522 (N_1522,In_2327,In_162);
and U1523 (N_1523,In_1812,In_2047);
nand U1524 (N_1524,In_672,In_1215);
and U1525 (N_1525,In_1873,In_1817);
nor U1526 (N_1526,In_1978,In_949);
and U1527 (N_1527,In_1100,In_776);
or U1528 (N_1528,In_997,In_1399);
nor U1529 (N_1529,In_1617,In_497);
or U1530 (N_1530,In_2212,In_567);
nand U1531 (N_1531,In_1348,In_2007);
and U1532 (N_1532,In_154,In_1377);
and U1533 (N_1533,In_667,In_1034);
nor U1534 (N_1534,In_267,In_623);
nor U1535 (N_1535,In_2416,In_1408);
and U1536 (N_1536,In_2445,In_1143);
and U1537 (N_1537,In_1069,In_1996);
xor U1538 (N_1538,In_1812,In_640);
and U1539 (N_1539,In_2000,In_543);
and U1540 (N_1540,In_1315,In_1102);
and U1541 (N_1541,In_1709,In_959);
nor U1542 (N_1542,In_1879,In_2137);
or U1543 (N_1543,In_1875,In_529);
nor U1544 (N_1544,In_737,In_61);
nor U1545 (N_1545,In_978,In_2228);
nand U1546 (N_1546,In_1409,In_763);
and U1547 (N_1547,In_872,In_1360);
or U1548 (N_1548,In_2326,In_2195);
nand U1549 (N_1549,In_1559,In_1008);
nand U1550 (N_1550,In_1226,In_356);
nor U1551 (N_1551,In_966,In_666);
nand U1552 (N_1552,In_785,In_1462);
nand U1553 (N_1553,In_376,In_1872);
nand U1554 (N_1554,In_790,In_2060);
nand U1555 (N_1555,In_61,In_2271);
nor U1556 (N_1556,In_1101,In_557);
or U1557 (N_1557,In_1353,In_331);
or U1558 (N_1558,In_1555,In_382);
and U1559 (N_1559,In_2286,In_598);
xor U1560 (N_1560,In_1518,In_1467);
nor U1561 (N_1561,In_1094,In_862);
and U1562 (N_1562,In_231,In_1250);
or U1563 (N_1563,In_2103,In_1400);
nand U1564 (N_1564,In_1796,In_951);
or U1565 (N_1565,In_1712,In_839);
nor U1566 (N_1566,In_2148,In_308);
or U1567 (N_1567,In_981,In_910);
or U1568 (N_1568,In_398,In_458);
and U1569 (N_1569,In_672,In_707);
and U1570 (N_1570,In_1467,In_2061);
nor U1571 (N_1571,In_2300,In_1751);
nor U1572 (N_1572,In_2071,In_184);
and U1573 (N_1573,In_1370,In_1843);
nor U1574 (N_1574,In_225,In_2085);
nor U1575 (N_1575,In_1213,In_1099);
or U1576 (N_1576,In_191,In_537);
nand U1577 (N_1577,In_711,In_1588);
nor U1578 (N_1578,In_2126,In_1244);
and U1579 (N_1579,In_922,In_2004);
xnor U1580 (N_1580,In_2053,In_897);
or U1581 (N_1581,In_2277,In_2420);
and U1582 (N_1582,In_1801,In_956);
and U1583 (N_1583,In_2166,In_907);
or U1584 (N_1584,In_30,In_108);
nand U1585 (N_1585,In_1682,In_1447);
nor U1586 (N_1586,In_1684,In_761);
and U1587 (N_1587,In_271,In_1362);
or U1588 (N_1588,In_37,In_186);
nand U1589 (N_1589,In_2022,In_801);
or U1590 (N_1590,In_1175,In_420);
nor U1591 (N_1591,In_1481,In_817);
and U1592 (N_1592,In_1975,In_1960);
or U1593 (N_1593,In_1053,In_1340);
nor U1594 (N_1594,In_676,In_2288);
nand U1595 (N_1595,In_1612,In_1549);
nor U1596 (N_1596,In_1888,In_1028);
nor U1597 (N_1597,In_273,In_1668);
or U1598 (N_1598,In_1085,In_1318);
nand U1599 (N_1599,In_14,In_387);
nand U1600 (N_1600,In_190,In_294);
or U1601 (N_1601,In_588,In_1248);
or U1602 (N_1602,In_2094,In_1811);
or U1603 (N_1603,In_1344,In_358);
nor U1604 (N_1604,In_1646,In_1995);
nor U1605 (N_1605,In_339,In_2107);
xor U1606 (N_1606,In_1539,In_1624);
or U1607 (N_1607,In_730,In_856);
or U1608 (N_1608,In_425,In_1425);
xnor U1609 (N_1609,In_1738,In_1219);
nor U1610 (N_1610,In_2344,In_1662);
or U1611 (N_1611,In_1170,In_1519);
xnor U1612 (N_1612,In_1775,In_1602);
nor U1613 (N_1613,In_691,In_1578);
nor U1614 (N_1614,In_1456,In_1017);
and U1615 (N_1615,In_2315,In_289);
or U1616 (N_1616,In_880,In_603);
nand U1617 (N_1617,In_2229,In_456);
nand U1618 (N_1618,In_1022,In_533);
nand U1619 (N_1619,In_374,In_420);
nand U1620 (N_1620,In_1555,In_2140);
nand U1621 (N_1621,In_1908,In_638);
nor U1622 (N_1622,In_263,In_1221);
nor U1623 (N_1623,In_1977,In_1182);
and U1624 (N_1624,In_860,In_2211);
and U1625 (N_1625,In_324,In_360);
and U1626 (N_1626,In_403,In_1608);
nor U1627 (N_1627,In_1298,In_206);
or U1628 (N_1628,In_1659,In_1855);
nand U1629 (N_1629,In_1193,In_1595);
and U1630 (N_1630,In_1962,In_176);
and U1631 (N_1631,In_76,In_675);
nor U1632 (N_1632,In_2464,In_1628);
nand U1633 (N_1633,In_1160,In_1343);
xnor U1634 (N_1634,In_2442,In_1991);
nor U1635 (N_1635,In_1466,In_1770);
and U1636 (N_1636,In_2065,In_1671);
nor U1637 (N_1637,In_539,In_2399);
or U1638 (N_1638,In_937,In_2277);
nand U1639 (N_1639,In_1075,In_216);
or U1640 (N_1640,In_60,In_942);
nor U1641 (N_1641,In_849,In_563);
nor U1642 (N_1642,In_681,In_1605);
nor U1643 (N_1643,In_1935,In_129);
and U1644 (N_1644,In_206,In_1163);
nand U1645 (N_1645,In_600,In_144);
xnor U1646 (N_1646,In_2276,In_1110);
xnor U1647 (N_1647,In_1538,In_1283);
nor U1648 (N_1648,In_2475,In_2040);
or U1649 (N_1649,In_963,In_1086);
or U1650 (N_1650,In_1270,In_1513);
nand U1651 (N_1651,In_2338,In_655);
or U1652 (N_1652,In_2028,In_2230);
and U1653 (N_1653,In_2351,In_1137);
or U1654 (N_1654,In_1833,In_689);
and U1655 (N_1655,In_2377,In_837);
or U1656 (N_1656,In_973,In_81);
and U1657 (N_1657,In_78,In_848);
nor U1658 (N_1658,In_2219,In_2064);
and U1659 (N_1659,In_651,In_2415);
xor U1660 (N_1660,In_1025,In_1654);
and U1661 (N_1661,In_1740,In_404);
nand U1662 (N_1662,In_2180,In_533);
and U1663 (N_1663,In_1134,In_283);
nand U1664 (N_1664,In_840,In_1841);
and U1665 (N_1665,In_1345,In_2231);
and U1666 (N_1666,In_43,In_252);
xnor U1667 (N_1667,In_2405,In_668);
nor U1668 (N_1668,In_1162,In_1499);
or U1669 (N_1669,In_1400,In_1424);
nor U1670 (N_1670,In_1436,In_1083);
nor U1671 (N_1671,In_407,In_1246);
or U1672 (N_1672,In_370,In_213);
or U1673 (N_1673,In_1103,In_55);
nor U1674 (N_1674,In_465,In_2460);
and U1675 (N_1675,In_818,In_943);
nor U1676 (N_1676,In_1900,In_25);
or U1677 (N_1677,In_2143,In_2370);
and U1678 (N_1678,In_199,In_507);
or U1679 (N_1679,In_1968,In_606);
nand U1680 (N_1680,In_78,In_1693);
and U1681 (N_1681,In_91,In_1454);
nor U1682 (N_1682,In_2170,In_861);
nor U1683 (N_1683,In_872,In_946);
or U1684 (N_1684,In_1998,In_884);
nor U1685 (N_1685,In_2185,In_1917);
or U1686 (N_1686,In_1568,In_1613);
and U1687 (N_1687,In_2255,In_559);
xor U1688 (N_1688,In_2061,In_677);
and U1689 (N_1689,In_900,In_1352);
xor U1690 (N_1690,In_1404,In_1568);
nand U1691 (N_1691,In_1395,In_2242);
or U1692 (N_1692,In_819,In_1413);
and U1693 (N_1693,In_80,In_1211);
or U1694 (N_1694,In_1304,In_55);
xnor U1695 (N_1695,In_1209,In_2242);
or U1696 (N_1696,In_401,In_282);
and U1697 (N_1697,In_1091,In_533);
and U1698 (N_1698,In_1317,In_1641);
nor U1699 (N_1699,In_174,In_31);
nor U1700 (N_1700,In_2031,In_429);
nor U1701 (N_1701,In_1590,In_1603);
nor U1702 (N_1702,In_1686,In_1409);
xor U1703 (N_1703,In_2487,In_342);
nor U1704 (N_1704,In_1357,In_562);
and U1705 (N_1705,In_2130,In_820);
or U1706 (N_1706,In_1274,In_662);
or U1707 (N_1707,In_113,In_2375);
nor U1708 (N_1708,In_188,In_2362);
nor U1709 (N_1709,In_1841,In_479);
nor U1710 (N_1710,In_2045,In_1421);
and U1711 (N_1711,In_2485,In_2075);
or U1712 (N_1712,In_153,In_419);
and U1713 (N_1713,In_347,In_2305);
and U1714 (N_1714,In_1056,In_1268);
and U1715 (N_1715,In_1717,In_2017);
nand U1716 (N_1716,In_1190,In_1953);
nor U1717 (N_1717,In_1699,In_269);
and U1718 (N_1718,In_882,In_323);
or U1719 (N_1719,In_2352,In_52);
nor U1720 (N_1720,In_564,In_1098);
or U1721 (N_1721,In_1200,In_1838);
nor U1722 (N_1722,In_1502,In_928);
nand U1723 (N_1723,In_569,In_1052);
nor U1724 (N_1724,In_1136,In_1775);
or U1725 (N_1725,In_1808,In_986);
or U1726 (N_1726,In_338,In_429);
nor U1727 (N_1727,In_1354,In_1637);
nor U1728 (N_1728,In_1057,In_1146);
nand U1729 (N_1729,In_1462,In_952);
nor U1730 (N_1730,In_259,In_2487);
nand U1731 (N_1731,In_1873,In_2420);
nor U1732 (N_1732,In_942,In_803);
and U1733 (N_1733,In_1755,In_2077);
and U1734 (N_1734,In_1566,In_1987);
and U1735 (N_1735,In_403,In_902);
or U1736 (N_1736,In_1833,In_1661);
nand U1737 (N_1737,In_2482,In_147);
nor U1738 (N_1738,In_2253,In_1130);
and U1739 (N_1739,In_686,In_678);
nor U1740 (N_1740,In_1164,In_946);
nor U1741 (N_1741,In_554,In_1732);
nor U1742 (N_1742,In_277,In_516);
xor U1743 (N_1743,In_1019,In_159);
nand U1744 (N_1744,In_1115,In_1137);
and U1745 (N_1745,In_603,In_190);
nor U1746 (N_1746,In_465,In_2004);
or U1747 (N_1747,In_998,In_517);
and U1748 (N_1748,In_304,In_1317);
or U1749 (N_1749,In_1659,In_1988);
and U1750 (N_1750,In_976,In_2201);
and U1751 (N_1751,In_897,In_1929);
nor U1752 (N_1752,In_858,In_936);
nand U1753 (N_1753,In_1832,In_427);
nand U1754 (N_1754,In_1487,In_29);
nand U1755 (N_1755,In_845,In_785);
and U1756 (N_1756,In_2293,In_2391);
and U1757 (N_1757,In_120,In_587);
and U1758 (N_1758,In_534,In_1902);
xor U1759 (N_1759,In_2303,In_1639);
and U1760 (N_1760,In_1497,In_180);
nand U1761 (N_1761,In_657,In_829);
nor U1762 (N_1762,In_1558,In_2384);
or U1763 (N_1763,In_491,In_199);
or U1764 (N_1764,In_213,In_2277);
nand U1765 (N_1765,In_1760,In_188);
and U1766 (N_1766,In_606,In_2360);
nand U1767 (N_1767,In_400,In_1601);
or U1768 (N_1768,In_2227,In_1282);
nor U1769 (N_1769,In_994,In_1018);
or U1770 (N_1770,In_1031,In_248);
nand U1771 (N_1771,In_1914,In_1185);
nand U1772 (N_1772,In_2448,In_2216);
nor U1773 (N_1773,In_193,In_1599);
nand U1774 (N_1774,In_194,In_1576);
and U1775 (N_1775,In_1228,In_555);
nor U1776 (N_1776,In_1898,In_2257);
nand U1777 (N_1777,In_1725,In_248);
or U1778 (N_1778,In_1100,In_47);
and U1779 (N_1779,In_554,In_851);
nand U1780 (N_1780,In_1498,In_1275);
xnor U1781 (N_1781,In_511,In_1248);
nand U1782 (N_1782,In_794,In_1774);
and U1783 (N_1783,In_169,In_1004);
nor U1784 (N_1784,In_1,In_385);
nor U1785 (N_1785,In_2316,In_2137);
nor U1786 (N_1786,In_1017,In_935);
nor U1787 (N_1787,In_2310,In_509);
and U1788 (N_1788,In_1295,In_1115);
nor U1789 (N_1789,In_2180,In_341);
and U1790 (N_1790,In_2264,In_1690);
and U1791 (N_1791,In_2373,In_2069);
nand U1792 (N_1792,In_351,In_1085);
or U1793 (N_1793,In_2497,In_2309);
or U1794 (N_1794,In_441,In_2012);
or U1795 (N_1795,In_2290,In_1229);
and U1796 (N_1796,In_2484,In_1614);
and U1797 (N_1797,In_289,In_2464);
or U1798 (N_1798,In_784,In_544);
nand U1799 (N_1799,In_426,In_1692);
nor U1800 (N_1800,In_182,In_1549);
or U1801 (N_1801,In_1294,In_1036);
nor U1802 (N_1802,In_138,In_777);
nor U1803 (N_1803,In_1838,In_1639);
or U1804 (N_1804,In_1295,In_2449);
and U1805 (N_1805,In_277,In_1405);
or U1806 (N_1806,In_2215,In_1396);
or U1807 (N_1807,In_1613,In_1096);
nor U1808 (N_1808,In_176,In_1957);
nand U1809 (N_1809,In_828,In_82);
nand U1810 (N_1810,In_1546,In_1869);
or U1811 (N_1811,In_1294,In_469);
and U1812 (N_1812,In_1386,In_786);
nor U1813 (N_1813,In_2231,In_2329);
or U1814 (N_1814,In_25,In_129);
or U1815 (N_1815,In_441,In_1596);
xor U1816 (N_1816,In_1696,In_460);
nor U1817 (N_1817,In_203,In_995);
nor U1818 (N_1818,In_526,In_16);
or U1819 (N_1819,In_29,In_1860);
nor U1820 (N_1820,In_2426,In_1765);
or U1821 (N_1821,In_1553,In_1897);
and U1822 (N_1822,In_2016,In_1224);
nor U1823 (N_1823,In_2155,In_259);
xnor U1824 (N_1824,In_502,In_1138);
nand U1825 (N_1825,In_1152,In_788);
or U1826 (N_1826,In_992,In_522);
or U1827 (N_1827,In_2051,In_1403);
and U1828 (N_1828,In_1538,In_1465);
and U1829 (N_1829,In_373,In_774);
or U1830 (N_1830,In_1457,In_880);
or U1831 (N_1831,In_1916,In_2479);
nor U1832 (N_1832,In_479,In_2059);
nor U1833 (N_1833,In_2020,In_764);
nand U1834 (N_1834,In_371,In_2097);
or U1835 (N_1835,In_958,In_1599);
nand U1836 (N_1836,In_1073,In_1197);
or U1837 (N_1837,In_553,In_516);
or U1838 (N_1838,In_1579,In_1133);
and U1839 (N_1839,In_1190,In_1721);
or U1840 (N_1840,In_476,In_416);
nor U1841 (N_1841,In_1235,In_117);
nand U1842 (N_1842,In_871,In_1536);
or U1843 (N_1843,In_164,In_2460);
nand U1844 (N_1844,In_1234,In_155);
nor U1845 (N_1845,In_187,In_274);
nor U1846 (N_1846,In_135,In_1668);
nor U1847 (N_1847,In_235,In_906);
and U1848 (N_1848,In_776,In_952);
or U1849 (N_1849,In_868,In_1672);
and U1850 (N_1850,In_1501,In_1029);
nand U1851 (N_1851,In_294,In_250);
nor U1852 (N_1852,In_1246,In_279);
nor U1853 (N_1853,In_857,In_960);
or U1854 (N_1854,In_1329,In_1234);
and U1855 (N_1855,In_1111,In_91);
nor U1856 (N_1856,In_1036,In_2431);
and U1857 (N_1857,In_2288,In_2342);
nor U1858 (N_1858,In_846,In_1099);
nor U1859 (N_1859,In_2112,In_2117);
nand U1860 (N_1860,In_606,In_568);
and U1861 (N_1861,In_2336,In_473);
xor U1862 (N_1862,In_1302,In_1658);
nor U1863 (N_1863,In_1975,In_1332);
and U1864 (N_1864,In_233,In_45);
or U1865 (N_1865,In_489,In_131);
nor U1866 (N_1866,In_965,In_387);
nor U1867 (N_1867,In_727,In_1708);
or U1868 (N_1868,In_2073,In_294);
or U1869 (N_1869,In_1583,In_2163);
or U1870 (N_1870,In_574,In_338);
and U1871 (N_1871,In_1904,In_1903);
nor U1872 (N_1872,In_2487,In_1069);
or U1873 (N_1873,In_2473,In_2269);
and U1874 (N_1874,In_1338,In_357);
nand U1875 (N_1875,In_1690,In_1647);
and U1876 (N_1876,In_793,In_1773);
or U1877 (N_1877,In_1877,In_1150);
nand U1878 (N_1878,In_1586,In_2004);
nand U1879 (N_1879,In_2262,In_1953);
or U1880 (N_1880,In_2309,In_2170);
or U1881 (N_1881,In_2155,In_424);
xnor U1882 (N_1882,In_1922,In_1010);
xor U1883 (N_1883,In_2485,In_1468);
nor U1884 (N_1884,In_1145,In_384);
nor U1885 (N_1885,In_1215,In_2255);
nor U1886 (N_1886,In_750,In_387);
or U1887 (N_1887,In_270,In_448);
nand U1888 (N_1888,In_1049,In_1854);
and U1889 (N_1889,In_2263,In_2031);
or U1890 (N_1890,In_914,In_347);
xor U1891 (N_1891,In_1956,In_1611);
and U1892 (N_1892,In_1169,In_388);
and U1893 (N_1893,In_790,In_464);
nand U1894 (N_1894,In_1494,In_104);
and U1895 (N_1895,In_1135,In_1740);
nor U1896 (N_1896,In_1508,In_1599);
nand U1897 (N_1897,In_1314,In_2128);
nand U1898 (N_1898,In_758,In_1494);
nor U1899 (N_1899,In_191,In_404);
nor U1900 (N_1900,In_1209,In_2263);
xnor U1901 (N_1901,In_288,In_890);
nand U1902 (N_1902,In_914,In_197);
and U1903 (N_1903,In_875,In_867);
nand U1904 (N_1904,In_1091,In_2246);
nor U1905 (N_1905,In_364,In_371);
nor U1906 (N_1906,In_1689,In_262);
or U1907 (N_1907,In_20,In_494);
nand U1908 (N_1908,In_2253,In_1660);
nor U1909 (N_1909,In_2232,In_825);
and U1910 (N_1910,In_976,In_1211);
nor U1911 (N_1911,In_1613,In_2160);
nor U1912 (N_1912,In_2267,In_1690);
or U1913 (N_1913,In_1885,In_1204);
or U1914 (N_1914,In_926,In_450);
or U1915 (N_1915,In_1169,In_1391);
nor U1916 (N_1916,In_150,In_321);
or U1917 (N_1917,In_874,In_826);
or U1918 (N_1918,In_237,In_2443);
nand U1919 (N_1919,In_1361,In_2383);
and U1920 (N_1920,In_140,In_69);
nor U1921 (N_1921,In_359,In_49);
and U1922 (N_1922,In_357,In_2495);
and U1923 (N_1923,In_245,In_210);
nand U1924 (N_1924,In_1432,In_578);
nor U1925 (N_1925,In_784,In_1800);
nand U1926 (N_1926,In_1847,In_1464);
and U1927 (N_1927,In_1505,In_266);
nor U1928 (N_1928,In_2457,In_468);
nor U1929 (N_1929,In_306,In_495);
nand U1930 (N_1930,In_612,In_41);
or U1931 (N_1931,In_2056,In_1869);
nand U1932 (N_1932,In_925,In_785);
xor U1933 (N_1933,In_160,In_844);
or U1934 (N_1934,In_2121,In_1637);
nor U1935 (N_1935,In_1030,In_275);
and U1936 (N_1936,In_598,In_2226);
nor U1937 (N_1937,In_2187,In_365);
nand U1938 (N_1938,In_1633,In_56);
or U1939 (N_1939,In_628,In_750);
nand U1940 (N_1940,In_284,In_1829);
and U1941 (N_1941,In_400,In_1253);
and U1942 (N_1942,In_2278,In_285);
and U1943 (N_1943,In_1925,In_1074);
xor U1944 (N_1944,In_798,In_2496);
or U1945 (N_1945,In_1378,In_708);
nand U1946 (N_1946,In_67,In_412);
or U1947 (N_1947,In_974,In_1861);
or U1948 (N_1948,In_2400,In_1301);
or U1949 (N_1949,In_1718,In_795);
and U1950 (N_1950,In_1435,In_305);
or U1951 (N_1951,In_1700,In_35);
nor U1952 (N_1952,In_1534,In_665);
nand U1953 (N_1953,In_1908,In_2111);
nand U1954 (N_1954,In_1656,In_310);
nand U1955 (N_1955,In_668,In_880);
and U1956 (N_1956,In_2206,In_316);
nor U1957 (N_1957,In_1076,In_2407);
or U1958 (N_1958,In_2255,In_408);
and U1959 (N_1959,In_875,In_1053);
and U1960 (N_1960,In_2108,In_763);
nor U1961 (N_1961,In_43,In_680);
nor U1962 (N_1962,In_351,In_1569);
or U1963 (N_1963,In_941,In_503);
or U1964 (N_1964,In_1507,In_1149);
or U1965 (N_1965,In_1054,In_1867);
nor U1966 (N_1966,In_281,In_802);
or U1967 (N_1967,In_934,In_834);
or U1968 (N_1968,In_527,In_1598);
xnor U1969 (N_1969,In_1271,In_1182);
or U1970 (N_1970,In_716,In_1238);
or U1971 (N_1971,In_1374,In_872);
or U1972 (N_1972,In_623,In_2499);
and U1973 (N_1973,In_2278,In_646);
or U1974 (N_1974,In_1240,In_1086);
or U1975 (N_1975,In_2499,In_385);
nor U1976 (N_1976,In_1349,In_365);
and U1977 (N_1977,In_1261,In_2194);
nand U1978 (N_1978,In_1706,In_1739);
and U1979 (N_1979,In_1421,In_2174);
and U1980 (N_1980,In_2176,In_982);
or U1981 (N_1981,In_864,In_1245);
nand U1982 (N_1982,In_2193,In_1347);
and U1983 (N_1983,In_170,In_1907);
or U1984 (N_1984,In_2054,In_1010);
or U1985 (N_1985,In_1679,In_822);
nor U1986 (N_1986,In_32,In_2259);
xnor U1987 (N_1987,In_1256,In_2345);
nor U1988 (N_1988,In_103,In_1260);
nor U1989 (N_1989,In_1255,In_2246);
xnor U1990 (N_1990,In_2079,In_1668);
nor U1991 (N_1991,In_1572,In_2192);
nand U1992 (N_1992,In_413,In_1291);
and U1993 (N_1993,In_1188,In_965);
nand U1994 (N_1994,In_1903,In_1755);
nand U1995 (N_1995,In_1349,In_2306);
nor U1996 (N_1996,In_295,In_1333);
and U1997 (N_1997,In_1416,In_2200);
and U1998 (N_1998,In_825,In_2128);
or U1999 (N_1999,In_1871,In_338);
or U2000 (N_2000,In_2107,In_1871);
or U2001 (N_2001,In_1084,In_2428);
nand U2002 (N_2002,In_822,In_2234);
nor U2003 (N_2003,In_446,In_1267);
and U2004 (N_2004,In_441,In_1343);
nand U2005 (N_2005,In_755,In_2088);
nand U2006 (N_2006,In_1688,In_2443);
or U2007 (N_2007,In_66,In_988);
nor U2008 (N_2008,In_1505,In_2384);
nand U2009 (N_2009,In_957,In_1534);
and U2010 (N_2010,In_2103,In_1401);
or U2011 (N_2011,In_579,In_1411);
or U2012 (N_2012,In_774,In_121);
or U2013 (N_2013,In_2350,In_229);
nor U2014 (N_2014,In_123,In_689);
or U2015 (N_2015,In_343,In_1620);
nand U2016 (N_2016,In_2470,In_1849);
nor U2017 (N_2017,In_1775,In_1756);
and U2018 (N_2018,In_1047,In_1108);
nand U2019 (N_2019,In_2336,In_1870);
nand U2020 (N_2020,In_610,In_583);
and U2021 (N_2021,In_722,In_526);
or U2022 (N_2022,In_1775,In_618);
or U2023 (N_2023,In_141,In_419);
or U2024 (N_2024,In_1349,In_400);
nand U2025 (N_2025,In_2056,In_1685);
or U2026 (N_2026,In_362,In_70);
nand U2027 (N_2027,In_2147,In_69);
nor U2028 (N_2028,In_2268,In_252);
and U2029 (N_2029,In_2353,In_2062);
and U2030 (N_2030,In_2021,In_2340);
and U2031 (N_2031,In_491,In_2385);
and U2032 (N_2032,In_1505,In_1625);
xor U2033 (N_2033,In_1931,In_445);
or U2034 (N_2034,In_1370,In_2208);
and U2035 (N_2035,In_564,In_987);
and U2036 (N_2036,In_368,In_875);
or U2037 (N_2037,In_1207,In_432);
or U2038 (N_2038,In_550,In_1324);
nand U2039 (N_2039,In_1349,In_1148);
nor U2040 (N_2040,In_1836,In_81);
nand U2041 (N_2041,In_1544,In_590);
and U2042 (N_2042,In_180,In_1453);
or U2043 (N_2043,In_2176,In_490);
or U2044 (N_2044,In_2450,In_950);
nor U2045 (N_2045,In_1846,In_2470);
or U2046 (N_2046,In_826,In_568);
nor U2047 (N_2047,In_1649,In_1747);
and U2048 (N_2048,In_550,In_618);
and U2049 (N_2049,In_778,In_1555);
nand U2050 (N_2050,In_1228,In_423);
and U2051 (N_2051,In_2054,In_164);
nor U2052 (N_2052,In_1883,In_2337);
nand U2053 (N_2053,In_33,In_1864);
or U2054 (N_2054,In_2351,In_1805);
or U2055 (N_2055,In_1500,In_1271);
nor U2056 (N_2056,In_508,In_498);
or U2057 (N_2057,In_1798,In_1374);
nor U2058 (N_2058,In_961,In_319);
and U2059 (N_2059,In_1520,In_2123);
or U2060 (N_2060,In_702,In_270);
and U2061 (N_2061,In_1567,In_224);
or U2062 (N_2062,In_1146,In_2361);
nor U2063 (N_2063,In_2483,In_880);
nor U2064 (N_2064,In_843,In_1368);
nor U2065 (N_2065,In_558,In_1029);
or U2066 (N_2066,In_944,In_1135);
nand U2067 (N_2067,In_103,In_2137);
and U2068 (N_2068,In_364,In_1243);
nand U2069 (N_2069,In_682,In_2185);
nand U2070 (N_2070,In_690,In_1922);
nand U2071 (N_2071,In_920,In_734);
and U2072 (N_2072,In_2194,In_1518);
nand U2073 (N_2073,In_2451,In_2170);
nor U2074 (N_2074,In_842,In_2325);
or U2075 (N_2075,In_933,In_1517);
nor U2076 (N_2076,In_596,In_600);
nand U2077 (N_2077,In_659,In_2063);
and U2078 (N_2078,In_1485,In_1626);
nand U2079 (N_2079,In_1994,In_667);
nor U2080 (N_2080,In_1305,In_2206);
nand U2081 (N_2081,In_509,In_334);
nand U2082 (N_2082,In_1144,In_2012);
nand U2083 (N_2083,In_1900,In_732);
or U2084 (N_2084,In_1834,In_2314);
nand U2085 (N_2085,In_1671,In_1284);
nor U2086 (N_2086,In_1903,In_2119);
and U2087 (N_2087,In_92,In_1149);
nand U2088 (N_2088,In_1233,In_2405);
nor U2089 (N_2089,In_680,In_307);
and U2090 (N_2090,In_316,In_1227);
or U2091 (N_2091,In_446,In_407);
and U2092 (N_2092,In_1465,In_1454);
or U2093 (N_2093,In_617,In_1030);
nor U2094 (N_2094,In_484,In_765);
and U2095 (N_2095,In_923,In_894);
and U2096 (N_2096,In_983,In_275);
nand U2097 (N_2097,In_2409,In_2325);
xor U2098 (N_2098,In_894,In_157);
or U2099 (N_2099,In_617,In_39);
nand U2100 (N_2100,In_2137,In_317);
and U2101 (N_2101,In_1297,In_813);
or U2102 (N_2102,In_29,In_1236);
or U2103 (N_2103,In_1582,In_1742);
and U2104 (N_2104,In_639,In_52);
nor U2105 (N_2105,In_539,In_54);
nand U2106 (N_2106,In_1328,In_23);
nor U2107 (N_2107,In_1678,In_1662);
nand U2108 (N_2108,In_862,In_598);
nand U2109 (N_2109,In_1694,In_1362);
or U2110 (N_2110,In_2291,In_675);
nand U2111 (N_2111,In_1436,In_432);
or U2112 (N_2112,In_1300,In_2299);
nor U2113 (N_2113,In_1036,In_710);
nand U2114 (N_2114,In_1564,In_1882);
nor U2115 (N_2115,In_2246,In_255);
nor U2116 (N_2116,In_1537,In_480);
nand U2117 (N_2117,In_1682,In_1622);
or U2118 (N_2118,In_1555,In_1017);
or U2119 (N_2119,In_2227,In_616);
nand U2120 (N_2120,In_1663,In_2334);
nor U2121 (N_2121,In_1955,In_1266);
nand U2122 (N_2122,In_2299,In_1823);
and U2123 (N_2123,In_1494,In_2195);
nand U2124 (N_2124,In_894,In_1237);
or U2125 (N_2125,In_746,In_435);
nor U2126 (N_2126,In_2074,In_2404);
nand U2127 (N_2127,In_1509,In_1484);
nand U2128 (N_2128,In_832,In_2223);
xnor U2129 (N_2129,In_455,In_929);
nor U2130 (N_2130,In_2039,In_162);
nor U2131 (N_2131,In_2083,In_482);
or U2132 (N_2132,In_1906,In_1785);
nand U2133 (N_2133,In_91,In_2188);
or U2134 (N_2134,In_1843,In_2149);
or U2135 (N_2135,In_520,In_1870);
nand U2136 (N_2136,In_450,In_1015);
nand U2137 (N_2137,In_1815,In_691);
nor U2138 (N_2138,In_606,In_1572);
nor U2139 (N_2139,In_919,In_21);
or U2140 (N_2140,In_2340,In_2282);
nor U2141 (N_2141,In_712,In_2024);
nand U2142 (N_2142,In_1443,In_1329);
or U2143 (N_2143,In_1168,In_2431);
xor U2144 (N_2144,In_276,In_478);
or U2145 (N_2145,In_686,In_434);
and U2146 (N_2146,In_1988,In_1792);
or U2147 (N_2147,In_1567,In_829);
and U2148 (N_2148,In_1336,In_1445);
or U2149 (N_2149,In_168,In_2460);
nor U2150 (N_2150,In_539,In_768);
and U2151 (N_2151,In_2461,In_866);
or U2152 (N_2152,In_333,In_581);
or U2153 (N_2153,In_1332,In_1804);
nor U2154 (N_2154,In_337,In_329);
nor U2155 (N_2155,In_1421,In_1262);
nor U2156 (N_2156,In_1295,In_793);
nor U2157 (N_2157,In_1700,In_38);
nor U2158 (N_2158,In_1864,In_2395);
xnor U2159 (N_2159,In_806,In_1515);
nor U2160 (N_2160,In_1929,In_1909);
nor U2161 (N_2161,In_2269,In_884);
nor U2162 (N_2162,In_496,In_164);
or U2163 (N_2163,In_1153,In_59);
and U2164 (N_2164,In_750,In_2490);
or U2165 (N_2165,In_623,In_1825);
nand U2166 (N_2166,In_294,In_934);
or U2167 (N_2167,In_417,In_1573);
and U2168 (N_2168,In_669,In_1382);
nand U2169 (N_2169,In_1022,In_1299);
nand U2170 (N_2170,In_1545,In_2039);
nor U2171 (N_2171,In_305,In_871);
nor U2172 (N_2172,In_1752,In_726);
nor U2173 (N_2173,In_1629,In_2259);
nor U2174 (N_2174,In_17,In_664);
nor U2175 (N_2175,In_902,In_1500);
nor U2176 (N_2176,In_1293,In_1907);
and U2177 (N_2177,In_876,In_822);
or U2178 (N_2178,In_2114,In_652);
nand U2179 (N_2179,In_631,In_754);
or U2180 (N_2180,In_132,In_1434);
or U2181 (N_2181,In_1956,In_812);
and U2182 (N_2182,In_1376,In_1135);
nand U2183 (N_2183,In_29,In_1971);
nor U2184 (N_2184,In_517,In_690);
and U2185 (N_2185,In_2371,In_1680);
nor U2186 (N_2186,In_531,In_574);
xor U2187 (N_2187,In_1344,In_2367);
nor U2188 (N_2188,In_1646,In_1309);
and U2189 (N_2189,In_388,In_992);
nand U2190 (N_2190,In_2397,In_2418);
or U2191 (N_2191,In_1895,In_81);
and U2192 (N_2192,In_1968,In_2136);
and U2193 (N_2193,In_2032,In_1376);
or U2194 (N_2194,In_1833,In_481);
or U2195 (N_2195,In_2454,In_1301);
and U2196 (N_2196,In_2305,In_1423);
and U2197 (N_2197,In_140,In_1257);
and U2198 (N_2198,In_114,In_1199);
and U2199 (N_2199,In_2186,In_1977);
and U2200 (N_2200,In_2408,In_1927);
nor U2201 (N_2201,In_690,In_800);
nor U2202 (N_2202,In_828,In_1346);
and U2203 (N_2203,In_2378,In_1983);
or U2204 (N_2204,In_1012,In_1706);
or U2205 (N_2205,In_1778,In_1681);
nor U2206 (N_2206,In_879,In_1633);
and U2207 (N_2207,In_1183,In_184);
or U2208 (N_2208,In_2016,In_958);
and U2209 (N_2209,In_1737,In_2413);
or U2210 (N_2210,In_730,In_933);
or U2211 (N_2211,In_647,In_1113);
nor U2212 (N_2212,In_1955,In_408);
nand U2213 (N_2213,In_1629,In_395);
nand U2214 (N_2214,In_2022,In_454);
nor U2215 (N_2215,In_2436,In_450);
xor U2216 (N_2216,In_2313,In_1408);
or U2217 (N_2217,In_959,In_1474);
nand U2218 (N_2218,In_1378,In_1866);
nor U2219 (N_2219,In_1510,In_830);
or U2220 (N_2220,In_1396,In_534);
and U2221 (N_2221,In_766,In_1920);
nor U2222 (N_2222,In_443,In_767);
nor U2223 (N_2223,In_1852,In_1821);
nand U2224 (N_2224,In_1209,In_1356);
nand U2225 (N_2225,In_1119,In_1535);
nand U2226 (N_2226,In_1981,In_167);
nand U2227 (N_2227,In_1253,In_2230);
or U2228 (N_2228,In_2376,In_931);
nand U2229 (N_2229,In_1340,In_879);
nand U2230 (N_2230,In_2260,In_2246);
or U2231 (N_2231,In_1971,In_1405);
and U2232 (N_2232,In_2433,In_878);
or U2233 (N_2233,In_693,In_1412);
or U2234 (N_2234,In_17,In_1923);
nor U2235 (N_2235,In_1287,In_1204);
or U2236 (N_2236,In_2375,In_1170);
nand U2237 (N_2237,In_624,In_466);
xor U2238 (N_2238,In_228,In_1384);
nor U2239 (N_2239,In_2384,In_1776);
xnor U2240 (N_2240,In_1815,In_416);
or U2241 (N_2241,In_430,In_1775);
or U2242 (N_2242,In_1514,In_2197);
and U2243 (N_2243,In_1121,In_1766);
or U2244 (N_2244,In_1697,In_585);
and U2245 (N_2245,In_453,In_293);
nand U2246 (N_2246,In_2096,In_549);
and U2247 (N_2247,In_588,In_1801);
and U2248 (N_2248,In_523,In_1769);
nand U2249 (N_2249,In_2131,In_880);
nor U2250 (N_2250,In_207,In_355);
nor U2251 (N_2251,In_260,In_574);
or U2252 (N_2252,In_1725,In_2146);
nand U2253 (N_2253,In_1543,In_1640);
and U2254 (N_2254,In_375,In_1710);
and U2255 (N_2255,In_2414,In_1892);
and U2256 (N_2256,In_2294,In_772);
or U2257 (N_2257,In_1015,In_1174);
and U2258 (N_2258,In_1388,In_1908);
nand U2259 (N_2259,In_580,In_396);
nor U2260 (N_2260,In_81,In_2278);
nor U2261 (N_2261,In_1030,In_1290);
nor U2262 (N_2262,In_148,In_732);
and U2263 (N_2263,In_2425,In_848);
nand U2264 (N_2264,In_2118,In_2146);
nand U2265 (N_2265,In_140,In_1030);
nand U2266 (N_2266,In_1128,In_287);
and U2267 (N_2267,In_2406,In_1960);
or U2268 (N_2268,In_569,In_1990);
nand U2269 (N_2269,In_1841,In_1813);
or U2270 (N_2270,In_2255,In_1255);
nor U2271 (N_2271,In_151,In_839);
nor U2272 (N_2272,In_1926,In_1080);
and U2273 (N_2273,In_2330,In_1850);
or U2274 (N_2274,In_409,In_2027);
nand U2275 (N_2275,In_1671,In_405);
nor U2276 (N_2276,In_2187,In_79);
nor U2277 (N_2277,In_1606,In_1602);
or U2278 (N_2278,In_33,In_2171);
or U2279 (N_2279,In_1423,In_971);
and U2280 (N_2280,In_2291,In_116);
nor U2281 (N_2281,In_1562,In_1992);
or U2282 (N_2282,In_1355,In_418);
nand U2283 (N_2283,In_1096,In_1720);
and U2284 (N_2284,In_2257,In_642);
or U2285 (N_2285,In_1456,In_1441);
nand U2286 (N_2286,In_232,In_134);
nor U2287 (N_2287,In_484,In_1540);
nand U2288 (N_2288,In_1573,In_2010);
nand U2289 (N_2289,In_1725,In_435);
nand U2290 (N_2290,In_1919,In_789);
nor U2291 (N_2291,In_352,In_999);
nor U2292 (N_2292,In_1500,In_708);
nand U2293 (N_2293,In_1026,In_1099);
nand U2294 (N_2294,In_61,In_1948);
or U2295 (N_2295,In_1104,In_546);
nand U2296 (N_2296,In_83,In_1105);
nor U2297 (N_2297,In_1314,In_1483);
nor U2298 (N_2298,In_2370,In_1243);
nand U2299 (N_2299,In_2007,In_97);
and U2300 (N_2300,In_261,In_1008);
or U2301 (N_2301,In_519,In_883);
nor U2302 (N_2302,In_2001,In_1324);
and U2303 (N_2303,In_2213,In_2098);
xnor U2304 (N_2304,In_1895,In_1864);
nand U2305 (N_2305,In_2394,In_200);
nand U2306 (N_2306,In_209,In_29);
and U2307 (N_2307,In_1100,In_683);
nand U2308 (N_2308,In_1690,In_294);
or U2309 (N_2309,In_957,In_758);
nor U2310 (N_2310,In_772,In_1018);
and U2311 (N_2311,In_1464,In_1067);
or U2312 (N_2312,In_1683,In_1786);
nand U2313 (N_2313,In_1497,In_704);
and U2314 (N_2314,In_696,In_417);
xnor U2315 (N_2315,In_1812,In_1980);
and U2316 (N_2316,In_2486,In_450);
nand U2317 (N_2317,In_651,In_1295);
nand U2318 (N_2318,In_1371,In_980);
nor U2319 (N_2319,In_979,In_909);
and U2320 (N_2320,In_934,In_1021);
nand U2321 (N_2321,In_2476,In_853);
nor U2322 (N_2322,In_208,In_1722);
nor U2323 (N_2323,In_829,In_1301);
or U2324 (N_2324,In_1516,In_1570);
nor U2325 (N_2325,In_315,In_1850);
and U2326 (N_2326,In_46,In_1543);
and U2327 (N_2327,In_1096,In_740);
or U2328 (N_2328,In_248,In_2132);
nor U2329 (N_2329,In_431,In_1668);
or U2330 (N_2330,In_1906,In_2220);
xor U2331 (N_2331,In_1448,In_2333);
and U2332 (N_2332,In_346,In_453);
nor U2333 (N_2333,In_2168,In_2284);
and U2334 (N_2334,In_1733,In_1648);
or U2335 (N_2335,In_2445,In_748);
nor U2336 (N_2336,In_243,In_700);
nand U2337 (N_2337,In_1739,In_984);
nor U2338 (N_2338,In_2474,In_955);
nor U2339 (N_2339,In_47,In_0);
nand U2340 (N_2340,In_1185,In_2067);
nor U2341 (N_2341,In_334,In_1088);
nor U2342 (N_2342,In_2010,In_341);
nand U2343 (N_2343,In_226,In_303);
or U2344 (N_2344,In_2463,In_755);
nand U2345 (N_2345,In_1570,In_2210);
nor U2346 (N_2346,In_1307,In_512);
or U2347 (N_2347,In_862,In_2365);
and U2348 (N_2348,In_275,In_1533);
and U2349 (N_2349,In_930,In_2328);
or U2350 (N_2350,In_1562,In_445);
nor U2351 (N_2351,In_1272,In_948);
and U2352 (N_2352,In_518,In_1359);
or U2353 (N_2353,In_1968,In_2321);
or U2354 (N_2354,In_1546,In_670);
nor U2355 (N_2355,In_325,In_2233);
and U2356 (N_2356,In_226,In_473);
or U2357 (N_2357,In_1741,In_1823);
nor U2358 (N_2358,In_61,In_2176);
or U2359 (N_2359,In_2185,In_242);
or U2360 (N_2360,In_1861,In_2302);
nor U2361 (N_2361,In_637,In_1700);
nor U2362 (N_2362,In_881,In_1521);
and U2363 (N_2363,In_23,In_1130);
nand U2364 (N_2364,In_783,In_1985);
or U2365 (N_2365,In_1126,In_104);
nand U2366 (N_2366,In_992,In_1949);
and U2367 (N_2367,In_664,In_1434);
and U2368 (N_2368,In_2191,In_704);
nand U2369 (N_2369,In_2209,In_1831);
and U2370 (N_2370,In_1,In_1550);
and U2371 (N_2371,In_2438,In_1705);
nor U2372 (N_2372,In_287,In_620);
and U2373 (N_2373,In_660,In_842);
xor U2374 (N_2374,In_2414,In_1077);
and U2375 (N_2375,In_681,In_898);
nand U2376 (N_2376,In_2367,In_803);
and U2377 (N_2377,In_746,In_560);
and U2378 (N_2378,In_1374,In_1823);
or U2379 (N_2379,In_1377,In_2310);
nor U2380 (N_2380,In_1568,In_379);
and U2381 (N_2381,In_2128,In_1520);
or U2382 (N_2382,In_1852,In_1260);
and U2383 (N_2383,In_1684,In_1071);
nor U2384 (N_2384,In_826,In_464);
nand U2385 (N_2385,In_1726,In_2005);
nor U2386 (N_2386,In_520,In_649);
xnor U2387 (N_2387,In_2375,In_785);
nand U2388 (N_2388,In_1774,In_728);
or U2389 (N_2389,In_939,In_1828);
or U2390 (N_2390,In_1839,In_1744);
or U2391 (N_2391,In_1038,In_2077);
nor U2392 (N_2392,In_749,In_147);
or U2393 (N_2393,In_1254,In_1084);
nor U2394 (N_2394,In_43,In_1132);
or U2395 (N_2395,In_1817,In_1605);
nor U2396 (N_2396,In_116,In_500);
nand U2397 (N_2397,In_2470,In_1677);
nand U2398 (N_2398,In_2493,In_2302);
nor U2399 (N_2399,In_2292,In_1237);
nand U2400 (N_2400,In_2406,In_1200);
and U2401 (N_2401,In_1118,In_1050);
nor U2402 (N_2402,In_1645,In_2197);
nand U2403 (N_2403,In_734,In_2308);
nor U2404 (N_2404,In_2267,In_296);
and U2405 (N_2405,In_652,In_2273);
or U2406 (N_2406,In_2312,In_1778);
and U2407 (N_2407,In_993,In_1699);
nand U2408 (N_2408,In_1216,In_2208);
xor U2409 (N_2409,In_2020,In_732);
or U2410 (N_2410,In_2135,In_2021);
nand U2411 (N_2411,In_2034,In_259);
nor U2412 (N_2412,In_1100,In_111);
nand U2413 (N_2413,In_2363,In_2405);
nand U2414 (N_2414,In_1294,In_541);
or U2415 (N_2415,In_2366,In_2401);
nor U2416 (N_2416,In_297,In_1918);
or U2417 (N_2417,In_517,In_2281);
or U2418 (N_2418,In_566,In_2122);
or U2419 (N_2419,In_1053,In_2416);
or U2420 (N_2420,In_1365,In_590);
nand U2421 (N_2421,In_159,In_1838);
nor U2422 (N_2422,In_78,In_1591);
nor U2423 (N_2423,In_4,In_1413);
or U2424 (N_2424,In_1714,In_36);
nand U2425 (N_2425,In_483,In_1464);
and U2426 (N_2426,In_213,In_450);
and U2427 (N_2427,In_1165,In_1764);
nor U2428 (N_2428,In_1957,In_1133);
or U2429 (N_2429,In_141,In_1946);
nor U2430 (N_2430,In_1677,In_704);
and U2431 (N_2431,In_1861,In_2294);
or U2432 (N_2432,In_2001,In_558);
or U2433 (N_2433,In_906,In_1959);
and U2434 (N_2434,In_628,In_1401);
nand U2435 (N_2435,In_1185,In_770);
or U2436 (N_2436,In_461,In_1788);
and U2437 (N_2437,In_326,In_202);
and U2438 (N_2438,In_2226,In_761);
and U2439 (N_2439,In_459,In_2357);
and U2440 (N_2440,In_2451,In_930);
nand U2441 (N_2441,In_1451,In_1576);
nor U2442 (N_2442,In_2152,In_52);
nor U2443 (N_2443,In_1657,In_2296);
or U2444 (N_2444,In_307,In_1234);
nand U2445 (N_2445,In_1310,In_1855);
or U2446 (N_2446,In_1129,In_1152);
and U2447 (N_2447,In_1100,In_1739);
nor U2448 (N_2448,In_1139,In_544);
and U2449 (N_2449,In_2139,In_1974);
nor U2450 (N_2450,In_1561,In_2308);
nor U2451 (N_2451,In_2268,In_917);
nand U2452 (N_2452,In_1805,In_2143);
nor U2453 (N_2453,In_1623,In_1220);
nand U2454 (N_2454,In_294,In_2113);
nor U2455 (N_2455,In_1037,In_1552);
nor U2456 (N_2456,In_463,In_75);
xnor U2457 (N_2457,In_465,In_1222);
and U2458 (N_2458,In_1168,In_853);
or U2459 (N_2459,In_1149,In_169);
and U2460 (N_2460,In_693,In_2191);
or U2461 (N_2461,In_871,In_1392);
nand U2462 (N_2462,In_289,In_1703);
and U2463 (N_2463,In_2404,In_1787);
or U2464 (N_2464,In_2035,In_1650);
xnor U2465 (N_2465,In_175,In_1416);
or U2466 (N_2466,In_768,In_2354);
and U2467 (N_2467,In_2482,In_705);
or U2468 (N_2468,In_1479,In_777);
and U2469 (N_2469,In_970,In_294);
nor U2470 (N_2470,In_2460,In_631);
nand U2471 (N_2471,In_1503,In_883);
or U2472 (N_2472,In_1217,In_824);
and U2473 (N_2473,In_251,In_2215);
nand U2474 (N_2474,In_60,In_1889);
nor U2475 (N_2475,In_980,In_1020);
and U2476 (N_2476,In_97,In_2419);
or U2477 (N_2477,In_2365,In_1863);
nor U2478 (N_2478,In_2340,In_1311);
and U2479 (N_2479,In_191,In_2093);
or U2480 (N_2480,In_2381,In_1428);
nor U2481 (N_2481,In_1654,In_218);
xnor U2482 (N_2482,In_806,In_661);
nand U2483 (N_2483,In_845,In_2198);
nand U2484 (N_2484,In_1679,In_1277);
nand U2485 (N_2485,In_2223,In_1711);
or U2486 (N_2486,In_1454,In_315);
nor U2487 (N_2487,In_165,In_560);
or U2488 (N_2488,In_148,In_1589);
and U2489 (N_2489,In_1171,In_1674);
nand U2490 (N_2490,In_106,In_15);
and U2491 (N_2491,In_823,In_2189);
and U2492 (N_2492,In_1156,In_1151);
or U2493 (N_2493,In_2389,In_595);
nor U2494 (N_2494,In_266,In_443);
or U2495 (N_2495,In_1279,In_302);
and U2496 (N_2496,In_114,In_876);
nor U2497 (N_2497,In_1926,In_1749);
and U2498 (N_2498,In_2082,In_2183);
and U2499 (N_2499,In_2303,In_2062);
nand U2500 (N_2500,In_1083,In_840);
or U2501 (N_2501,In_1783,In_1849);
and U2502 (N_2502,In_1334,In_268);
nand U2503 (N_2503,In_1578,In_317);
nand U2504 (N_2504,In_1523,In_1575);
or U2505 (N_2505,In_1684,In_863);
nor U2506 (N_2506,In_1643,In_510);
or U2507 (N_2507,In_502,In_727);
nor U2508 (N_2508,In_598,In_1016);
nand U2509 (N_2509,In_266,In_2087);
xnor U2510 (N_2510,In_762,In_255);
nand U2511 (N_2511,In_1911,In_2247);
or U2512 (N_2512,In_2045,In_1360);
and U2513 (N_2513,In_96,In_976);
and U2514 (N_2514,In_404,In_978);
nand U2515 (N_2515,In_1271,In_806);
or U2516 (N_2516,In_1770,In_814);
nor U2517 (N_2517,In_1653,In_257);
nand U2518 (N_2518,In_1126,In_1775);
or U2519 (N_2519,In_215,In_523);
or U2520 (N_2520,In_2102,In_1276);
nor U2521 (N_2521,In_2118,In_726);
and U2522 (N_2522,In_2109,In_939);
nand U2523 (N_2523,In_2262,In_2220);
nor U2524 (N_2524,In_1075,In_1804);
and U2525 (N_2525,In_473,In_1081);
nand U2526 (N_2526,In_1897,In_694);
or U2527 (N_2527,In_2035,In_451);
nand U2528 (N_2528,In_2499,In_1364);
and U2529 (N_2529,In_2484,In_240);
or U2530 (N_2530,In_269,In_1474);
or U2531 (N_2531,In_2085,In_1147);
and U2532 (N_2532,In_1422,In_468);
or U2533 (N_2533,In_1467,In_1515);
and U2534 (N_2534,In_1554,In_835);
nand U2535 (N_2535,In_608,In_1404);
nor U2536 (N_2536,In_1255,In_1239);
and U2537 (N_2537,In_345,In_1045);
or U2538 (N_2538,In_401,In_1507);
xnor U2539 (N_2539,In_2300,In_1059);
nor U2540 (N_2540,In_928,In_472);
nand U2541 (N_2541,In_2229,In_2353);
nor U2542 (N_2542,In_654,In_231);
or U2543 (N_2543,In_1537,In_1814);
nand U2544 (N_2544,In_967,In_901);
nand U2545 (N_2545,In_1032,In_1785);
or U2546 (N_2546,In_2072,In_1822);
or U2547 (N_2547,In_2463,In_1847);
xnor U2548 (N_2548,In_725,In_2448);
nand U2549 (N_2549,In_1136,In_2235);
or U2550 (N_2550,In_298,In_1482);
nor U2551 (N_2551,In_1142,In_2382);
and U2552 (N_2552,In_1668,In_410);
nand U2553 (N_2553,In_703,In_2296);
nand U2554 (N_2554,In_172,In_992);
or U2555 (N_2555,In_888,In_414);
or U2556 (N_2556,In_1481,In_512);
nor U2557 (N_2557,In_1434,In_111);
nor U2558 (N_2558,In_1301,In_2462);
or U2559 (N_2559,In_8,In_1328);
nor U2560 (N_2560,In_3,In_1034);
or U2561 (N_2561,In_2180,In_253);
nand U2562 (N_2562,In_1456,In_1448);
and U2563 (N_2563,In_2268,In_952);
or U2564 (N_2564,In_2019,In_106);
nand U2565 (N_2565,In_681,In_515);
nand U2566 (N_2566,In_1087,In_1686);
nor U2567 (N_2567,In_2434,In_1740);
nand U2568 (N_2568,In_423,In_1825);
or U2569 (N_2569,In_940,In_1643);
and U2570 (N_2570,In_2129,In_1288);
and U2571 (N_2571,In_1350,In_2076);
and U2572 (N_2572,In_1093,In_1671);
nor U2573 (N_2573,In_2278,In_160);
nor U2574 (N_2574,In_464,In_167);
nand U2575 (N_2575,In_275,In_1894);
nor U2576 (N_2576,In_2043,In_268);
and U2577 (N_2577,In_1168,In_1507);
xor U2578 (N_2578,In_640,In_1357);
or U2579 (N_2579,In_2270,In_2451);
nand U2580 (N_2580,In_663,In_1322);
or U2581 (N_2581,In_117,In_2061);
and U2582 (N_2582,In_1118,In_694);
xnor U2583 (N_2583,In_320,In_329);
and U2584 (N_2584,In_102,In_2083);
xnor U2585 (N_2585,In_1746,In_633);
nand U2586 (N_2586,In_2386,In_1863);
nor U2587 (N_2587,In_1506,In_583);
or U2588 (N_2588,In_502,In_626);
or U2589 (N_2589,In_373,In_955);
xor U2590 (N_2590,In_1445,In_1729);
nand U2591 (N_2591,In_488,In_66);
or U2592 (N_2592,In_2064,In_1151);
nand U2593 (N_2593,In_1286,In_27);
or U2594 (N_2594,In_118,In_767);
nand U2595 (N_2595,In_485,In_897);
nand U2596 (N_2596,In_677,In_562);
or U2597 (N_2597,In_1754,In_2229);
and U2598 (N_2598,In_299,In_1706);
nor U2599 (N_2599,In_905,In_1562);
or U2600 (N_2600,In_1186,In_189);
nor U2601 (N_2601,In_520,In_563);
and U2602 (N_2602,In_1300,In_2372);
or U2603 (N_2603,In_729,In_1177);
or U2604 (N_2604,In_552,In_2148);
or U2605 (N_2605,In_542,In_664);
or U2606 (N_2606,In_1544,In_2294);
and U2607 (N_2607,In_1757,In_1015);
nor U2608 (N_2608,In_2024,In_24);
or U2609 (N_2609,In_1434,In_2052);
xor U2610 (N_2610,In_1227,In_1341);
nor U2611 (N_2611,In_1224,In_1477);
or U2612 (N_2612,In_1925,In_1643);
or U2613 (N_2613,In_1758,In_1814);
nor U2614 (N_2614,In_492,In_561);
and U2615 (N_2615,In_1480,In_1813);
or U2616 (N_2616,In_718,In_2091);
nor U2617 (N_2617,In_1208,In_1278);
nor U2618 (N_2618,In_1173,In_2168);
nor U2619 (N_2619,In_1194,In_1081);
nor U2620 (N_2620,In_2465,In_163);
nand U2621 (N_2621,In_181,In_2281);
nor U2622 (N_2622,In_19,In_1600);
and U2623 (N_2623,In_1893,In_2340);
nand U2624 (N_2624,In_735,In_906);
nand U2625 (N_2625,In_2446,In_1077);
and U2626 (N_2626,In_1918,In_1583);
and U2627 (N_2627,In_1347,In_1719);
and U2628 (N_2628,In_2364,In_2346);
and U2629 (N_2629,In_1813,In_2194);
nand U2630 (N_2630,In_367,In_642);
and U2631 (N_2631,In_1598,In_1990);
nor U2632 (N_2632,In_1317,In_2174);
or U2633 (N_2633,In_114,In_1452);
and U2634 (N_2634,In_2198,In_1734);
nor U2635 (N_2635,In_1008,In_1641);
or U2636 (N_2636,In_1339,In_1523);
nor U2637 (N_2637,In_168,In_2029);
nand U2638 (N_2638,In_794,In_468);
xor U2639 (N_2639,In_488,In_1738);
or U2640 (N_2640,In_454,In_511);
and U2641 (N_2641,In_409,In_32);
nor U2642 (N_2642,In_1593,In_335);
nor U2643 (N_2643,In_1858,In_1806);
or U2644 (N_2644,In_1379,In_1485);
nor U2645 (N_2645,In_1261,In_1567);
nor U2646 (N_2646,In_830,In_1924);
or U2647 (N_2647,In_658,In_1342);
nand U2648 (N_2648,In_1785,In_82);
or U2649 (N_2649,In_1271,In_293);
and U2650 (N_2650,In_1805,In_1755);
or U2651 (N_2651,In_2148,In_16);
nor U2652 (N_2652,In_1085,In_892);
or U2653 (N_2653,In_1636,In_1648);
or U2654 (N_2654,In_2312,In_728);
and U2655 (N_2655,In_465,In_2219);
xor U2656 (N_2656,In_663,In_532);
or U2657 (N_2657,In_1010,In_1533);
nand U2658 (N_2658,In_2234,In_33);
nor U2659 (N_2659,In_85,In_2235);
nand U2660 (N_2660,In_1157,In_1905);
or U2661 (N_2661,In_2488,In_566);
nor U2662 (N_2662,In_1148,In_1432);
nand U2663 (N_2663,In_1349,In_2412);
and U2664 (N_2664,In_417,In_2175);
and U2665 (N_2665,In_2047,In_1885);
and U2666 (N_2666,In_1326,In_540);
nor U2667 (N_2667,In_1231,In_1085);
and U2668 (N_2668,In_2233,In_1414);
or U2669 (N_2669,In_252,In_1161);
or U2670 (N_2670,In_1897,In_816);
nand U2671 (N_2671,In_412,In_2099);
nor U2672 (N_2672,In_130,In_1029);
and U2673 (N_2673,In_1517,In_1772);
nor U2674 (N_2674,In_131,In_92);
nor U2675 (N_2675,In_777,In_2065);
nand U2676 (N_2676,In_1340,In_681);
nand U2677 (N_2677,In_376,In_1713);
or U2678 (N_2678,In_1140,In_1585);
or U2679 (N_2679,In_2289,In_1324);
or U2680 (N_2680,In_1441,In_202);
nor U2681 (N_2681,In_1500,In_2226);
nand U2682 (N_2682,In_1681,In_1976);
nand U2683 (N_2683,In_1338,In_1779);
and U2684 (N_2684,In_721,In_2000);
nand U2685 (N_2685,In_1857,In_2240);
xnor U2686 (N_2686,In_1848,In_1037);
nand U2687 (N_2687,In_1934,In_1447);
or U2688 (N_2688,In_941,In_728);
nand U2689 (N_2689,In_654,In_1718);
nor U2690 (N_2690,In_964,In_561);
nor U2691 (N_2691,In_1749,In_1562);
nor U2692 (N_2692,In_1568,In_603);
or U2693 (N_2693,In_1564,In_1441);
and U2694 (N_2694,In_699,In_1652);
nand U2695 (N_2695,In_299,In_748);
and U2696 (N_2696,In_2470,In_1856);
and U2697 (N_2697,In_452,In_2404);
and U2698 (N_2698,In_1211,In_1148);
nand U2699 (N_2699,In_1391,In_1733);
nor U2700 (N_2700,In_64,In_1473);
nand U2701 (N_2701,In_1562,In_933);
and U2702 (N_2702,In_88,In_900);
or U2703 (N_2703,In_2113,In_183);
nor U2704 (N_2704,In_1172,In_1175);
and U2705 (N_2705,In_1395,In_511);
or U2706 (N_2706,In_563,In_2165);
nor U2707 (N_2707,In_2181,In_1884);
and U2708 (N_2708,In_2159,In_2284);
nand U2709 (N_2709,In_475,In_1350);
and U2710 (N_2710,In_2004,In_1422);
and U2711 (N_2711,In_495,In_2046);
or U2712 (N_2712,In_1150,In_214);
nand U2713 (N_2713,In_389,In_1245);
and U2714 (N_2714,In_1090,In_2498);
and U2715 (N_2715,In_1897,In_712);
or U2716 (N_2716,In_400,In_1251);
or U2717 (N_2717,In_429,In_2083);
or U2718 (N_2718,In_2204,In_609);
nand U2719 (N_2719,In_1566,In_1973);
and U2720 (N_2720,In_477,In_523);
and U2721 (N_2721,In_255,In_1736);
or U2722 (N_2722,In_1243,In_430);
and U2723 (N_2723,In_1073,In_147);
nand U2724 (N_2724,In_1478,In_86);
nor U2725 (N_2725,In_1632,In_2450);
nor U2726 (N_2726,In_529,In_1770);
and U2727 (N_2727,In_2338,In_2283);
nand U2728 (N_2728,In_826,In_1050);
and U2729 (N_2729,In_865,In_998);
nand U2730 (N_2730,In_253,In_1693);
and U2731 (N_2731,In_152,In_1460);
nor U2732 (N_2732,In_1518,In_931);
xnor U2733 (N_2733,In_55,In_2221);
or U2734 (N_2734,In_582,In_1284);
or U2735 (N_2735,In_2244,In_1413);
and U2736 (N_2736,In_358,In_1312);
or U2737 (N_2737,In_2336,In_2395);
or U2738 (N_2738,In_942,In_1378);
nor U2739 (N_2739,In_10,In_1064);
nand U2740 (N_2740,In_1245,In_1430);
and U2741 (N_2741,In_397,In_1112);
xor U2742 (N_2742,In_1392,In_2070);
nand U2743 (N_2743,In_2204,In_842);
nor U2744 (N_2744,In_1241,In_587);
nand U2745 (N_2745,In_90,In_2007);
or U2746 (N_2746,In_60,In_1287);
and U2747 (N_2747,In_733,In_1634);
or U2748 (N_2748,In_728,In_743);
nand U2749 (N_2749,In_1114,In_863);
nand U2750 (N_2750,In_1397,In_2347);
and U2751 (N_2751,In_436,In_902);
and U2752 (N_2752,In_1688,In_624);
nand U2753 (N_2753,In_798,In_583);
nand U2754 (N_2754,In_2167,In_2449);
or U2755 (N_2755,In_72,In_933);
or U2756 (N_2756,In_282,In_141);
and U2757 (N_2757,In_2315,In_1139);
nor U2758 (N_2758,In_2356,In_1034);
nor U2759 (N_2759,In_2094,In_397);
or U2760 (N_2760,In_930,In_975);
nand U2761 (N_2761,In_265,In_717);
nand U2762 (N_2762,In_1644,In_563);
nand U2763 (N_2763,In_2009,In_464);
nand U2764 (N_2764,In_1625,In_1987);
nand U2765 (N_2765,In_1971,In_235);
nand U2766 (N_2766,In_939,In_804);
or U2767 (N_2767,In_746,In_2287);
nor U2768 (N_2768,In_2024,In_1623);
nand U2769 (N_2769,In_726,In_1356);
or U2770 (N_2770,In_814,In_277);
or U2771 (N_2771,In_2440,In_2438);
nor U2772 (N_2772,In_292,In_2002);
and U2773 (N_2773,In_1392,In_2175);
nor U2774 (N_2774,In_1643,In_1517);
or U2775 (N_2775,In_2363,In_1852);
nand U2776 (N_2776,In_1401,In_1046);
nand U2777 (N_2777,In_78,In_1919);
nor U2778 (N_2778,In_2300,In_666);
and U2779 (N_2779,In_2063,In_1681);
nand U2780 (N_2780,In_2018,In_1042);
nor U2781 (N_2781,In_1699,In_530);
nand U2782 (N_2782,In_2331,In_1888);
or U2783 (N_2783,In_850,In_689);
nor U2784 (N_2784,In_1965,In_416);
nor U2785 (N_2785,In_398,In_887);
and U2786 (N_2786,In_471,In_1235);
nor U2787 (N_2787,In_300,In_1173);
and U2788 (N_2788,In_1330,In_573);
and U2789 (N_2789,In_623,In_1875);
nand U2790 (N_2790,In_2408,In_2118);
or U2791 (N_2791,In_450,In_1972);
or U2792 (N_2792,In_56,In_1963);
or U2793 (N_2793,In_323,In_1876);
nand U2794 (N_2794,In_762,In_253);
and U2795 (N_2795,In_2400,In_2439);
or U2796 (N_2796,In_1424,In_476);
xor U2797 (N_2797,In_1545,In_143);
or U2798 (N_2798,In_1482,In_182);
nor U2799 (N_2799,In_2078,In_1696);
nor U2800 (N_2800,In_1974,In_1958);
and U2801 (N_2801,In_336,In_940);
nand U2802 (N_2802,In_1181,In_419);
or U2803 (N_2803,In_718,In_42);
nor U2804 (N_2804,In_1578,In_1018);
and U2805 (N_2805,In_2265,In_2380);
and U2806 (N_2806,In_1332,In_1137);
nand U2807 (N_2807,In_1149,In_2370);
and U2808 (N_2808,In_2475,In_928);
and U2809 (N_2809,In_2469,In_2496);
and U2810 (N_2810,In_970,In_904);
nand U2811 (N_2811,In_1523,In_231);
nand U2812 (N_2812,In_2308,In_1152);
nor U2813 (N_2813,In_90,In_929);
and U2814 (N_2814,In_680,In_623);
nand U2815 (N_2815,In_2385,In_716);
and U2816 (N_2816,In_1209,In_392);
and U2817 (N_2817,In_2389,In_2020);
nor U2818 (N_2818,In_344,In_2460);
nor U2819 (N_2819,In_1230,In_1628);
and U2820 (N_2820,In_1462,In_2092);
nand U2821 (N_2821,In_475,In_46);
xor U2822 (N_2822,In_2083,In_1409);
and U2823 (N_2823,In_779,In_1105);
nor U2824 (N_2824,In_2013,In_1737);
nor U2825 (N_2825,In_145,In_197);
nand U2826 (N_2826,In_567,In_171);
and U2827 (N_2827,In_773,In_1537);
and U2828 (N_2828,In_2245,In_957);
and U2829 (N_2829,In_1982,In_237);
or U2830 (N_2830,In_48,In_1647);
nand U2831 (N_2831,In_853,In_1881);
and U2832 (N_2832,In_825,In_2361);
nand U2833 (N_2833,In_1630,In_2260);
or U2834 (N_2834,In_315,In_1223);
nand U2835 (N_2835,In_11,In_524);
or U2836 (N_2836,In_882,In_1458);
nand U2837 (N_2837,In_324,In_1187);
nor U2838 (N_2838,In_1447,In_1961);
nand U2839 (N_2839,In_1725,In_2087);
nor U2840 (N_2840,In_1042,In_1143);
nor U2841 (N_2841,In_734,In_1041);
and U2842 (N_2842,In_1970,In_2052);
and U2843 (N_2843,In_1988,In_302);
nand U2844 (N_2844,In_472,In_958);
and U2845 (N_2845,In_407,In_1669);
nor U2846 (N_2846,In_1265,In_225);
or U2847 (N_2847,In_1944,In_521);
xor U2848 (N_2848,In_785,In_1052);
or U2849 (N_2849,In_327,In_1097);
or U2850 (N_2850,In_1321,In_1398);
and U2851 (N_2851,In_220,In_2484);
and U2852 (N_2852,In_431,In_1493);
or U2853 (N_2853,In_1828,In_1120);
and U2854 (N_2854,In_2219,In_1499);
nor U2855 (N_2855,In_2005,In_251);
nand U2856 (N_2856,In_1695,In_173);
nand U2857 (N_2857,In_1919,In_1182);
nor U2858 (N_2858,In_2064,In_1653);
nor U2859 (N_2859,In_1972,In_683);
and U2860 (N_2860,In_684,In_1534);
or U2861 (N_2861,In_720,In_2028);
or U2862 (N_2862,In_1334,In_218);
nor U2863 (N_2863,In_102,In_342);
nor U2864 (N_2864,In_1967,In_2384);
nand U2865 (N_2865,In_1886,In_1405);
and U2866 (N_2866,In_998,In_1480);
nor U2867 (N_2867,In_177,In_1063);
nor U2868 (N_2868,In_329,In_2041);
or U2869 (N_2869,In_1957,In_292);
or U2870 (N_2870,In_734,In_1535);
or U2871 (N_2871,In_2285,In_1773);
nand U2872 (N_2872,In_850,In_2126);
nand U2873 (N_2873,In_1810,In_1888);
nor U2874 (N_2874,In_2335,In_1786);
and U2875 (N_2875,In_376,In_1640);
nand U2876 (N_2876,In_1664,In_1921);
nand U2877 (N_2877,In_2210,In_728);
nand U2878 (N_2878,In_1333,In_1081);
nand U2879 (N_2879,In_923,In_948);
nor U2880 (N_2880,In_853,In_1338);
nand U2881 (N_2881,In_978,In_743);
nand U2882 (N_2882,In_808,In_484);
nand U2883 (N_2883,In_2137,In_2276);
nand U2884 (N_2884,In_563,In_11);
nor U2885 (N_2885,In_1853,In_2394);
and U2886 (N_2886,In_1157,In_1788);
nor U2887 (N_2887,In_153,In_1145);
xnor U2888 (N_2888,In_61,In_812);
or U2889 (N_2889,In_148,In_1706);
and U2890 (N_2890,In_1068,In_1617);
or U2891 (N_2891,In_234,In_1386);
and U2892 (N_2892,In_2146,In_653);
nor U2893 (N_2893,In_2389,In_820);
nor U2894 (N_2894,In_633,In_1859);
nand U2895 (N_2895,In_1197,In_2361);
and U2896 (N_2896,In_566,In_1685);
nor U2897 (N_2897,In_1466,In_2194);
or U2898 (N_2898,In_1976,In_1818);
and U2899 (N_2899,In_2474,In_2216);
nor U2900 (N_2900,In_2020,In_1534);
nor U2901 (N_2901,In_622,In_3);
or U2902 (N_2902,In_1125,In_780);
nor U2903 (N_2903,In_2493,In_1532);
nor U2904 (N_2904,In_178,In_603);
and U2905 (N_2905,In_627,In_1984);
nand U2906 (N_2906,In_1144,In_595);
or U2907 (N_2907,In_2151,In_1771);
and U2908 (N_2908,In_528,In_2313);
nor U2909 (N_2909,In_417,In_1187);
nor U2910 (N_2910,In_2180,In_1908);
and U2911 (N_2911,In_1944,In_1670);
nor U2912 (N_2912,In_23,In_2222);
or U2913 (N_2913,In_1395,In_1993);
and U2914 (N_2914,In_1969,In_289);
nor U2915 (N_2915,In_341,In_602);
or U2916 (N_2916,In_2204,In_1841);
and U2917 (N_2917,In_706,In_2271);
and U2918 (N_2918,In_2172,In_397);
and U2919 (N_2919,In_1772,In_321);
nor U2920 (N_2920,In_1393,In_1242);
nand U2921 (N_2921,In_351,In_2008);
and U2922 (N_2922,In_489,In_971);
nand U2923 (N_2923,In_2458,In_1049);
nand U2924 (N_2924,In_1934,In_1747);
or U2925 (N_2925,In_710,In_1699);
or U2926 (N_2926,In_1488,In_1386);
xor U2927 (N_2927,In_362,In_2343);
and U2928 (N_2928,In_2225,In_1392);
nor U2929 (N_2929,In_1729,In_1029);
and U2930 (N_2930,In_1985,In_1153);
and U2931 (N_2931,In_2076,In_2374);
nand U2932 (N_2932,In_571,In_2132);
and U2933 (N_2933,In_2107,In_1214);
and U2934 (N_2934,In_1882,In_933);
nand U2935 (N_2935,In_1800,In_2255);
nand U2936 (N_2936,In_2302,In_1574);
xnor U2937 (N_2937,In_862,In_1496);
or U2938 (N_2938,In_1751,In_1019);
nor U2939 (N_2939,In_1577,In_1205);
xnor U2940 (N_2940,In_255,In_1382);
and U2941 (N_2941,In_377,In_244);
nor U2942 (N_2942,In_179,In_1076);
or U2943 (N_2943,In_272,In_1418);
nor U2944 (N_2944,In_2392,In_843);
or U2945 (N_2945,In_466,In_2487);
or U2946 (N_2946,In_1935,In_1565);
nor U2947 (N_2947,In_1896,In_1703);
nand U2948 (N_2948,In_2060,In_518);
nor U2949 (N_2949,In_639,In_299);
and U2950 (N_2950,In_2490,In_1509);
and U2951 (N_2951,In_1575,In_1022);
and U2952 (N_2952,In_644,In_2430);
or U2953 (N_2953,In_94,In_1799);
or U2954 (N_2954,In_2208,In_281);
or U2955 (N_2955,In_600,In_2087);
or U2956 (N_2956,In_1589,In_1448);
nor U2957 (N_2957,In_111,In_616);
or U2958 (N_2958,In_48,In_1260);
nand U2959 (N_2959,In_691,In_2284);
or U2960 (N_2960,In_917,In_754);
nor U2961 (N_2961,In_914,In_300);
nor U2962 (N_2962,In_1870,In_776);
or U2963 (N_2963,In_1550,In_2160);
nand U2964 (N_2964,In_638,In_310);
nand U2965 (N_2965,In_1421,In_2224);
nand U2966 (N_2966,In_138,In_1893);
or U2967 (N_2967,In_235,In_383);
and U2968 (N_2968,In_1440,In_125);
nand U2969 (N_2969,In_1084,In_1594);
nor U2970 (N_2970,In_731,In_1811);
nand U2971 (N_2971,In_2018,In_1848);
nand U2972 (N_2972,In_754,In_926);
and U2973 (N_2973,In_2063,In_2274);
and U2974 (N_2974,In_1421,In_813);
and U2975 (N_2975,In_2130,In_147);
and U2976 (N_2976,In_552,In_2488);
nand U2977 (N_2977,In_530,In_644);
and U2978 (N_2978,In_1965,In_1761);
nand U2979 (N_2979,In_818,In_2061);
nand U2980 (N_2980,In_806,In_202);
nand U2981 (N_2981,In_1277,In_618);
and U2982 (N_2982,In_1134,In_248);
or U2983 (N_2983,In_1386,In_63);
and U2984 (N_2984,In_1272,In_2291);
nor U2985 (N_2985,In_1590,In_2135);
nor U2986 (N_2986,In_639,In_886);
nor U2987 (N_2987,In_2474,In_146);
nand U2988 (N_2988,In_1195,In_933);
and U2989 (N_2989,In_1419,In_1979);
or U2990 (N_2990,In_562,In_1772);
nand U2991 (N_2991,In_1873,In_1289);
or U2992 (N_2992,In_388,In_1962);
or U2993 (N_2993,In_988,In_696);
or U2994 (N_2994,In_1254,In_1006);
and U2995 (N_2995,In_1353,In_709);
and U2996 (N_2996,In_706,In_2366);
or U2997 (N_2997,In_643,In_1633);
nor U2998 (N_2998,In_1519,In_1999);
nand U2999 (N_2999,In_440,In_1893);
nand U3000 (N_3000,In_1338,In_1478);
and U3001 (N_3001,In_497,In_283);
or U3002 (N_3002,In_1735,In_473);
nor U3003 (N_3003,In_273,In_396);
and U3004 (N_3004,In_1913,In_814);
and U3005 (N_3005,In_859,In_510);
or U3006 (N_3006,In_1159,In_800);
or U3007 (N_3007,In_300,In_72);
nor U3008 (N_3008,In_619,In_2435);
and U3009 (N_3009,In_1151,In_213);
nand U3010 (N_3010,In_1264,In_2013);
or U3011 (N_3011,In_1005,In_2109);
or U3012 (N_3012,In_757,In_2383);
and U3013 (N_3013,In_1975,In_834);
and U3014 (N_3014,In_1,In_1903);
or U3015 (N_3015,In_2271,In_228);
and U3016 (N_3016,In_1277,In_1931);
and U3017 (N_3017,In_538,In_1124);
and U3018 (N_3018,In_297,In_862);
nor U3019 (N_3019,In_1435,In_172);
nor U3020 (N_3020,In_287,In_93);
or U3021 (N_3021,In_1201,In_1608);
or U3022 (N_3022,In_1474,In_292);
nor U3023 (N_3023,In_1395,In_304);
or U3024 (N_3024,In_1070,In_1929);
or U3025 (N_3025,In_147,In_1050);
and U3026 (N_3026,In_14,In_1364);
nand U3027 (N_3027,In_1830,In_1116);
and U3028 (N_3028,In_974,In_2283);
or U3029 (N_3029,In_2324,In_1105);
nor U3030 (N_3030,In_1808,In_1019);
nor U3031 (N_3031,In_1772,In_2017);
xnor U3032 (N_3032,In_408,In_1258);
or U3033 (N_3033,In_1889,In_2242);
nand U3034 (N_3034,In_1101,In_1772);
nand U3035 (N_3035,In_65,In_2372);
nor U3036 (N_3036,In_943,In_1563);
and U3037 (N_3037,In_2276,In_1850);
and U3038 (N_3038,In_1169,In_1226);
nor U3039 (N_3039,In_300,In_437);
nor U3040 (N_3040,In_2119,In_1353);
or U3041 (N_3041,In_2023,In_1591);
nor U3042 (N_3042,In_240,In_361);
and U3043 (N_3043,In_154,In_872);
or U3044 (N_3044,In_667,In_1175);
nand U3045 (N_3045,In_1377,In_1524);
nor U3046 (N_3046,In_1218,In_137);
or U3047 (N_3047,In_2297,In_2434);
nor U3048 (N_3048,In_650,In_978);
nor U3049 (N_3049,In_1004,In_72);
and U3050 (N_3050,In_26,In_1982);
and U3051 (N_3051,In_480,In_1958);
nor U3052 (N_3052,In_1226,In_1523);
and U3053 (N_3053,In_245,In_1387);
and U3054 (N_3054,In_1411,In_993);
nor U3055 (N_3055,In_616,In_2140);
nand U3056 (N_3056,In_295,In_1689);
nor U3057 (N_3057,In_2469,In_925);
and U3058 (N_3058,In_2283,In_1044);
and U3059 (N_3059,In_1626,In_2477);
xnor U3060 (N_3060,In_516,In_1603);
and U3061 (N_3061,In_2325,In_1843);
nand U3062 (N_3062,In_70,In_1916);
nor U3063 (N_3063,In_1208,In_2304);
nor U3064 (N_3064,In_1803,In_295);
and U3065 (N_3065,In_2043,In_395);
and U3066 (N_3066,In_1589,In_2373);
or U3067 (N_3067,In_2332,In_1687);
nand U3068 (N_3068,In_1253,In_1081);
and U3069 (N_3069,In_1101,In_2048);
nand U3070 (N_3070,In_1791,In_1073);
nor U3071 (N_3071,In_265,In_607);
and U3072 (N_3072,In_1896,In_2302);
or U3073 (N_3073,In_1841,In_197);
nor U3074 (N_3074,In_137,In_214);
or U3075 (N_3075,In_1221,In_1563);
nor U3076 (N_3076,In_1478,In_2343);
or U3077 (N_3077,In_2281,In_420);
and U3078 (N_3078,In_2108,In_237);
nor U3079 (N_3079,In_2205,In_2005);
or U3080 (N_3080,In_503,In_1582);
nand U3081 (N_3081,In_1930,In_2369);
nand U3082 (N_3082,In_2157,In_1626);
nor U3083 (N_3083,In_2153,In_157);
and U3084 (N_3084,In_1073,In_164);
nand U3085 (N_3085,In_1303,In_1330);
nor U3086 (N_3086,In_849,In_713);
or U3087 (N_3087,In_234,In_713);
or U3088 (N_3088,In_2391,In_1117);
and U3089 (N_3089,In_69,In_2053);
xor U3090 (N_3090,In_1059,In_2480);
or U3091 (N_3091,In_65,In_404);
nor U3092 (N_3092,In_196,In_897);
and U3093 (N_3093,In_1289,In_2181);
nor U3094 (N_3094,In_1815,In_2193);
nor U3095 (N_3095,In_2465,In_551);
nor U3096 (N_3096,In_2008,In_2353);
xnor U3097 (N_3097,In_2313,In_2499);
nor U3098 (N_3098,In_2060,In_2279);
xnor U3099 (N_3099,In_2351,In_313);
or U3100 (N_3100,In_1775,In_1048);
nand U3101 (N_3101,In_2386,In_1769);
and U3102 (N_3102,In_784,In_328);
nor U3103 (N_3103,In_736,In_1970);
and U3104 (N_3104,In_564,In_2082);
nand U3105 (N_3105,In_1618,In_1331);
or U3106 (N_3106,In_515,In_1907);
or U3107 (N_3107,In_1149,In_118);
and U3108 (N_3108,In_2412,In_433);
or U3109 (N_3109,In_915,In_2491);
nand U3110 (N_3110,In_1764,In_1443);
nor U3111 (N_3111,In_1881,In_573);
nor U3112 (N_3112,In_856,In_1147);
nand U3113 (N_3113,In_1290,In_1808);
nor U3114 (N_3114,In_1598,In_2428);
and U3115 (N_3115,In_1881,In_243);
nor U3116 (N_3116,In_2085,In_1711);
nor U3117 (N_3117,In_2288,In_65);
nand U3118 (N_3118,In_972,In_2107);
nand U3119 (N_3119,In_1422,In_112);
nor U3120 (N_3120,In_1045,In_1711);
nor U3121 (N_3121,In_1379,In_1376);
xor U3122 (N_3122,In_2133,In_912);
and U3123 (N_3123,In_392,In_1805);
nor U3124 (N_3124,In_2274,In_61);
nor U3125 (N_3125,In_1782,In_1151);
nor U3126 (N_3126,In_2269,In_840);
nand U3127 (N_3127,In_341,In_1589);
or U3128 (N_3128,In_848,In_1551);
nor U3129 (N_3129,In_1116,In_1515);
nor U3130 (N_3130,In_1063,In_1087);
and U3131 (N_3131,In_1077,In_2111);
nor U3132 (N_3132,In_330,In_230);
and U3133 (N_3133,In_69,In_1166);
nand U3134 (N_3134,In_1962,In_1119);
and U3135 (N_3135,In_1446,In_1654);
nand U3136 (N_3136,In_292,In_1629);
nor U3137 (N_3137,In_1213,In_834);
nand U3138 (N_3138,In_2093,In_2420);
nand U3139 (N_3139,In_826,In_1558);
and U3140 (N_3140,In_2219,In_981);
or U3141 (N_3141,In_3,In_58);
nor U3142 (N_3142,In_2103,In_1874);
nor U3143 (N_3143,In_57,In_1736);
or U3144 (N_3144,In_73,In_1397);
and U3145 (N_3145,In_1737,In_556);
nand U3146 (N_3146,In_4,In_473);
nor U3147 (N_3147,In_1984,In_1094);
or U3148 (N_3148,In_57,In_1640);
and U3149 (N_3149,In_1197,In_1092);
nor U3150 (N_3150,In_631,In_390);
and U3151 (N_3151,In_1121,In_1559);
nand U3152 (N_3152,In_2010,In_702);
nor U3153 (N_3153,In_1556,In_1770);
and U3154 (N_3154,In_1812,In_2071);
nand U3155 (N_3155,In_2359,In_2283);
nand U3156 (N_3156,In_2351,In_457);
nor U3157 (N_3157,In_843,In_172);
or U3158 (N_3158,In_1388,In_1007);
nand U3159 (N_3159,In_935,In_1968);
and U3160 (N_3160,In_1920,In_1261);
nor U3161 (N_3161,In_2377,In_2157);
or U3162 (N_3162,In_557,In_72);
or U3163 (N_3163,In_1359,In_2085);
and U3164 (N_3164,In_963,In_130);
and U3165 (N_3165,In_74,In_763);
nand U3166 (N_3166,In_822,In_1239);
nor U3167 (N_3167,In_1189,In_121);
or U3168 (N_3168,In_1767,In_2106);
and U3169 (N_3169,In_887,In_751);
nor U3170 (N_3170,In_1544,In_748);
nor U3171 (N_3171,In_413,In_1787);
or U3172 (N_3172,In_1393,In_463);
or U3173 (N_3173,In_1300,In_1091);
and U3174 (N_3174,In_2334,In_2379);
nor U3175 (N_3175,In_147,In_959);
or U3176 (N_3176,In_1334,In_2349);
and U3177 (N_3177,In_309,In_1092);
nand U3178 (N_3178,In_2460,In_969);
or U3179 (N_3179,In_1960,In_462);
xnor U3180 (N_3180,In_899,In_881);
nand U3181 (N_3181,In_59,In_311);
or U3182 (N_3182,In_975,In_318);
nand U3183 (N_3183,In_1466,In_658);
nor U3184 (N_3184,In_1345,In_1323);
nand U3185 (N_3185,In_685,In_553);
and U3186 (N_3186,In_1275,In_1034);
and U3187 (N_3187,In_2199,In_1200);
or U3188 (N_3188,In_1810,In_1741);
nor U3189 (N_3189,In_1798,In_25);
nand U3190 (N_3190,In_1880,In_2294);
nor U3191 (N_3191,In_1345,In_928);
nor U3192 (N_3192,In_2100,In_1007);
nand U3193 (N_3193,In_1946,In_932);
or U3194 (N_3194,In_2340,In_71);
nand U3195 (N_3195,In_2243,In_506);
nor U3196 (N_3196,In_528,In_2490);
nor U3197 (N_3197,In_2499,In_929);
or U3198 (N_3198,In_15,In_1215);
or U3199 (N_3199,In_554,In_618);
or U3200 (N_3200,In_2418,In_2304);
or U3201 (N_3201,In_2227,In_833);
nor U3202 (N_3202,In_1956,In_987);
or U3203 (N_3203,In_1456,In_75);
nor U3204 (N_3204,In_350,In_884);
nand U3205 (N_3205,In_2144,In_1132);
and U3206 (N_3206,In_48,In_1532);
or U3207 (N_3207,In_1169,In_2231);
or U3208 (N_3208,In_239,In_2085);
or U3209 (N_3209,In_2481,In_665);
and U3210 (N_3210,In_2308,In_349);
and U3211 (N_3211,In_321,In_1105);
or U3212 (N_3212,In_1756,In_210);
xor U3213 (N_3213,In_701,In_1770);
or U3214 (N_3214,In_2138,In_553);
and U3215 (N_3215,In_761,In_1407);
and U3216 (N_3216,In_195,In_2396);
nor U3217 (N_3217,In_2342,In_716);
or U3218 (N_3218,In_2127,In_544);
xor U3219 (N_3219,In_1071,In_2323);
nand U3220 (N_3220,In_974,In_493);
or U3221 (N_3221,In_211,In_1555);
and U3222 (N_3222,In_2169,In_1716);
nand U3223 (N_3223,In_902,In_1441);
or U3224 (N_3224,In_500,In_2252);
and U3225 (N_3225,In_2181,In_1782);
nor U3226 (N_3226,In_2470,In_855);
nand U3227 (N_3227,In_763,In_1571);
or U3228 (N_3228,In_2226,In_1720);
or U3229 (N_3229,In_288,In_135);
or U3230 (N_3230,In_752,In_695);
and U3231 (N_3231,In_596,In_1216);
or U3232 (N_3232,In_415,In_1260);
nand U3233 (N_3233,In_956,In_929);
or U3234 (N_3234,In_1657,In_1889);
and U3235 (N_3235,In_1878,In_1651);
nand U3236 (N_3236,In_2120,In_2078);
or U3237 (N_3237,In_1003,In_820);
and U3238 (N_3238,In_311,In_1769);
or U3239 (N_3239,In_1929,In_2253);
nor U3240 (N_3240,In_1793,In_305);
or U3241 (N_3241,In_761,In_1385);
and U3242 (N_3242,In_921,In_782);
and U3243 (N_3243,In_328,In_369);
nor U3244 (N_3244,In_1728,In_1894);
and U3245 (N_3245,In_1979,In_1529);
or U3246 (N_3246,In_182,In_2009);
or U3247 (N_3247,In_1183,In_691);
nor U3248 (N_3248,In_463,In_187);
xnor U3249 (N_3249,In_72,In_940);
nor U3250 (N_3250,In_414,In_2101);
nor U3251 (N_3251,In_1834,In_1516);
and U3252 (N_3252,In_111,In_1977);
nor U3253 (N_3253,In_280,In_530);
nor U3254 (N_3254,In_2376,In_316);
or U3255 (N_3255,In_573,In_392);
nand U3256 (N_3256,In_1639,In_799);
nor U3257 (N_3257,In_1776,In_1223);
or U3258 (N_3258,In_781,In_1993);
nand U3259 (N_3259,In_186,In_496);
nand U3260 (N_3260,In_403,In_1182);
and U3261 (N_3261,In_2354,In_1377);
nor U3262 (N_3262,In_2155,In_1250);
nor U3263 (N_3263,In_2335,In_712);
nand U3264 (N_3264,In_1423,In_1654);
or U3265 (N_3265,In_45,In_739);
or U3266 (N_3266,In_787,In_2483);
and U3267 (N_3267,In_1972,In_161);
and U3268 (N_3268,In_2399,In_398);
nor U3269 (N_3269,In_277,In_2350);
and U3270 (N_3270,In_2126,In_2284);
nand U3271 (N_3271,In_317,In_77);
nor U3272 (N_3272,In_2290,In_1988);
nand U3273 (N_3273,In_2087,In_819);
nor U3274 (N_3274,In_196,In_1510);
nor U3275 (N_3275,In_462,In_672);
nand U3276 (N_3276,In_1872,In_1713);
nor U3277 (N_3277,In_613,In_63);
or U3278 (N_3278,In_1972,In_806);
and U3279 (N_3279,In_264,In_2272);
nor U3280 (N_3280,In_1850,In_1461);
nand U3281 (N_3281,In_2110,In_2384);
and U3282 (N_3282,In_103,In_109);
nor U3283 (N_3283,In_1318,In_1237);
nor U3284 (N_3284,In_1524,In_1607);
nor U3285 (N_3285,In_932,In_1088);
nand U3286 (N_3286,In_756,In_2345);
nand U3287 (N_3287,In_1357,In_2377);
and U3288 (N_3288,In_1207,In_557);
xnor U3289 (N_3289,In_2488,In_29);
nor U3290 (N_3290,In_643,In_2305);
or U3291 (N_3291,In_2128,In_2099);
and U3292 (N_3292,In_2208,In_112);
nand U3293 (N_3293,In_672,In_688);
nor U3294 (N_3294,In_1423,In_457);
nand U3295 (N_3295,In_450,In_927);
and U3296 (N_3296,In_1243,In_453);
or U3297 (N_3297,In_1100,In_731);
and U3298 (N_3298,In_544,In_845);
or U3299 (N_3299,In_980,In_2484);
or U3300 (N_3300,In_1644,In_2477);
nand U3301 (N_3301,In_690,In_2367);
or U3302 (N_3302,In_773,In_529);
nor U3303 (N_3303,In_1444,In_2399);
or U3304 (N_3304,In_2356,In_1886);
or U3305 (N_3305,In_2029,In_128);
and U3306 (N_3306,In_832,In_2420);
xor U3307 (N_3307,In_2352,In_1509);
or U3308 (N_3308,In_1029,In_427);
nand U3309 (N_3309,In_117,In_796);
and U3310 (N_3310,In_2348,In_1489);
and U3311 (N_3311,In_893,In_1132);
and U3312 (N_3312,In_2425,In_2229);
nor U3313 (N_3313,In_1391,In_1528);
nand U3314 (N_3314,In_1843,In_768);
nor U3315 (N_3315,In_454,In_1488);
or U3316 (N_3316,In_1168,In_1395);
nand U3317 (N_3317,In_1619,In_2240);
and U3318 (N_3318,In_993,In_1364);
and U3319 (N_3319,In_1876,In_1806);
and U3320 (N_3320,In_1552,In_439);
nor U3321 (N_3321,In_250,In_1740);
nor U3322 (N_3322,In_539,In_1594);
and U3323 (N_3323,In_605,In_321);
nand U3324 (N_3324,In_1000,In_1958);
or U3325 (N_3325,In_43,In_1284);
nor U3326 (N_3326,In_2230,In_1207);
nand U3327 (N_3327,In_2204,In_1636);
and U3328 (N_3328,In_2180,In_2424);
nand U3329 (N_3329,In_967,In_294);
nor U3330 (N_3330,In_2395,In_1016);
and U3331 (N_3331,In_243,In_1447);
nand U3332 (N_3332,In_389,In_117);
or U3333 (N_3333,In_100,In_25);
nand U3334 (N_3334,In_2442,In_1424);
and U3335 (N_3335,In_99,In_155);
or U3336 (N_3336,In_516,In_377);
nand U3337 (N_3337,In_14,In_2463);
and U3338 (N_3338,In_2081,In_81);
nor U3339 (N_3339,In_1155,In_2437);
or U3340 (N_3340,In_1598,In_1576);
nand U3341 (N_3341,In_1771,In_552);
nand U3342 (N_3342,In_609,In_2274);
nand U3343 (N_3343,In_621,In_985);
and U3344 (N_3344,In_2467,In_2005);
nor U3345 (N_3345,In_2160,In_30);
nor U3346 (N_3346,In_2197,In_210);
nand U3347 (N_3347,In_2444,In_1468);
and U3348 (N_3348,In_230,In_2448);
and U3349 (N_3349,In_1713,In_1260);
and U3350 (N_3350,In_278,In_683);
nor U3351 (N_3351,In_345,In_2141);
nand U3352 (N_3352,In_2411,In_153);
nor U3353 (N_3353,In_1025,In_2498);
nor U3354 (N_3354,In_2373,In_7);
or U3355 (N_3355,In_1275,In_249);
or U3356 (N_3356,In_849,In_987);
nor U3357 (N_3357,In_756,In_1331);
or U3358 (N_3358,In_1206,In_327);
and U3359 (N_3359,In_2403,In_792);
nand U3360 (N_3360,In_1319,In_1542);
or U3361 (N_3361,In_122,In_1273);
and U3362 (N_3362,In_1568,In_975);
nand U3363 (N_3363,In_399,In_818);
and U3364 (N_3364,In_1420,In_354);
xnor U3365 (N_3365,In_946,In_2231);
nor U3366 (N_3366,In_2383,In_722);
nand U3367 (N_3367,In_1713,In_396);
nand U3368 (N_3368,In_1787,In_891);
nand U3369 (N_3369,In_1136,In_1467);
and U3370 (N_3370,In_935,In_675);
or U3371 (N_3371,In_769,In_1925);
nor U3372 (N_3372,In_2329,In_619);
or U3373 (N_3373,In_1958,In_2169);
nand U3374 (N_3374,In_1083,In_2312);
or U3375 (N_3375,In_2222,In_2069);
and U3376 (N_3376,In_2425,In_864);
nand U3377 (N_3377,In_888,In_701);
nor U3378 (N_3378,In_1575,In_1845);
and U3379 (N_3379,In_938,In_2402);
or U3380 (N_3380,In_594,In_1423);
or U3381 (N_3381,In_1681,In_651);
nor U3382 (N_3382,In_2400,In_1821);
and U3383 (N_3383,In_1916,In_186);
or U3384 (N_3384,In_1967,In_1650);
and U3385 (N_3385,In_1652,In_2069);
nor U3386 (N_3386,In_1360,In_39);
or U3387 (N_3387,In_1381,In_667);
and U3388 (N_3388,In_2260,In_2071);
nor U3389 (N_3389,In_236,In_260);
or U3390 (N_3390,In_1384,In_1126);
nand U3391 (N_3391,In_202,In_152);
xnor U3392 (N_3392,In_773,In_1573);
and U3393 (N_3393,In_669,In_1503);
or U3394 (N_3394,In_2060,In_1120);
nor U3395 (N_3395,In_1036,In_73);
xnor U3396 (N_3396,In_1356,In_369);
nand U3397 (N_3397,In_691,In_1296);
or U3398 (N_3398,In_259,In_66);
or U3399 (N_3399,In_2417,In_2050);
nand U3400 (N_3400,In_2431,In_1056);
nand U3401 (N_3401,In_532,In_424);
nor U3402 (N_3402,In_1479,In_1958);
nand U3403 (N_3403,In_1925,In_247);
and U3404 (N_3404,In_1058,In_2263);
nand U3405 (N_3405,In_1929,In_1029);
and U3406 (N_3406,In_967,In_1025);
and U3407 (N_3407,In_671,In_1520);
or U3408 (N_3408,In_1528,In_63);
or U3409 (N_3409,In_2326,In_1724);
nand U3410 (N_3410,In_2401,In_1480);
nor U3411 (N_3411,In_925,In_1651);
and U3412 (N_3412,In_888,In_1717);
nand U3413 (N_3413,In_1676,In_287);
or U3414 (N_3414,In_882,In_1323);
or U3415 (N_3415,In_1287,In_712);
nor U3416 (N_3416,In_424,In_510);
nor U3417 (N_3417,In_2051,In_1863);
or U3418 (N_3418,In_1788,In_1152);
or U3419 (N_3419,In_1220,In_902);
and U3420 (N_3420,In_1283,In_1353);
nor U3421 (N_3421,In_2307,In_581);
and U3422 (N_3422,In_1606,In_2354);
or U3423 (N_3423,In_1817,In_1302);
xnor U3424 (N_3424,In_2170,In_1839);
or U3425 (N_3425,In_972,In_214);
or U3426 (N_3426,In_2178,In_1262);
or U3427 (N_3427,In_734,In_2018);
nor U3428 (N_3428,In_1253,In_2465);
xnor U3429 (N_3429,In_1105,In_1898);
nor U3430 (N_3430,In_1836,In_132);
nand U3431 (N_3431,In_1409,In_1561);
and U3432 (N_3432,In_2448,In_2079);
and U3433 (N_3433,In_451,In_1844);
nand U3434 (N_3434,In_1153,In_1348);
or U3435 (N_3435,In_1310,In_286);
nor U3436 (N_3436,In_2400,In_1172);
nor U3437 (N_3437,In_1406,In_689);
and U3438 (N_3438,In_2328,In_2026);
or U3439 (N_3439,In_364,In_86);
and U3440 (N_3440,In_677,In_221);
nand U3441 (N_3441,In_2085,In_750);
and U3442 (N_3442,In_1273,In_2320);
nor U3443 (N_3443,In_191,In_1621);
nor U3444 (N_3444,In_1120,In_224);
nor U3445 (N_3445,In_1261,In_1078);
and U3446 (N_3446,In_1899,In_1047);
nor U3447 (N_3447,In_1989,In_106);
and U3448 (N_3448,In_246,In_1141);
or U3449 (N_3449,In_2378,In_1043);
or U3450 (N_3450,In_190,In_796);
and U3451 (N_3451,In_2029,In_437);
nor U3452 (N_3452,In_931,In_748);
nand U3453 (N_3453,In_944,In_1419);
or U3454 (N_3454,In_7,In_843);
nor U3455 (N_3455,In_2104,In_174);
nor U3456 (N_3456,In_790,In_344);
nand U3457 (N_3457,In_588,In_798);
or U3458 (N_3458,In_1245,In_371);
and U3459 (N_3459,In_2288,In_857);
and U3460 (N_3460,In_156,In_1867);
and U3461 (N_3461,In_1990,In_14);
and U3462 (N_3462,In_14,In_1771);
and U3463 (N_3463,In_1182,In_93);
and U3464 (N_3464,In_1490,In_1707);
and U3465 (N_3465,In_1462,In_900);
or U3466 (N_3466,In_849,In_691);
nand U3467 (N_3467,In_467,In_2493);
nor U3468 (N_3468,In_1172,In_1689);
nand U3469 (N_3469,In_1061,In_641);
and U3470 (N_3470,In_2022,In_2317);
or U3471 (N_3471,In_135,In_892);
and U3472 (N_3472,In_403,In_2214);
nor U3473 (N_3473,In_1643,In_1467);
and U3474 (N_3474,In_2263,In_748);
nand U3475 (N_3475,In_29,In_1798);
and U3476 (N_3476,In_1813,In_147);
nand U3477 (N_3477,In_988,In_1984);
nor U3478 (N_3478,In_195,In_1310);
nand U3479 (N_3479,In_2328,In_1959);
and U3480 (N_3480,In_525,In_2001);
or U3481 (N_3481,In_1266,In_2273);
and U3482 (N_3482,In_550,In_1263);
nor U3483 (N_3483,In_1521,In_2146);
nor U3484 (N_3484,In_323,In_522);
nand U3485 (N_3485,In_1968,In_2329);
xor U3486 (N_3486,In_2049,In_996);
nand U3487 (N_3487,In_1179,In_598);
nor U3488 (N_3488,In_368,In_2212);
nand U3489 (N_3489,In_1989,In_2404);
or U3490 (N_3490,In_1493,In_866);
and U3491 (N_3491,In_1883,In_1882);
nor U3492 (N_3492,In_498,In_1558);
nor U3493 (N_3493,In_337,In_41);
nor U3494 (N_3494,In_868,In_192);
nor U3495 (N_3495,In_1800,In_1015);
nand U3496 (N_3496,In_2338,In_1208);
nand U3497 (N_3497,In_942,In_2422);
and U3498 (N_3498,In_1510,In_1324);
nand U3499 (N_3499,In_132,In_1857);
nor U3500 (N_3500,In_20,In_2242);
nand U3501 (N_3501,In_1792,In_704);
and U3502 (N_3502,In_2021,In_2183);
nand U3503 (N_3503,In_1215,In_1479);
nor U3504 (N_3504,In_677,In_1915);
or U3505 (N_3505,In_474,In_690);
and U3506 (N_3506,In_287,In_2369);
and U3507 (N_3507,In_1296,In_1340);
nor U3508 (N_3508,In_61,In_1101);
nor U3509 (N_3509,In_931,In_1752);
or U3510 (N_3510,In_676,In_327);
nand U3511 (N_3511,In_2331,In_1644);
or U3512 (N_3512,In_1956,In_97);
nand U3513 (N_3513,In_1207,In_247);
nand U3514 (N_3514,In_1629,In_61);
xnor U3515 (N_3515,In_1,In_57);
or U3516 (N_3516,In_252,In_2153);
or U3517 (N_3517,In_2299,In_1586);
or U3518 (N_3518,In_35,In_489);
nand U3519 (N_3519,In_2199,In_1634);
nor U3520 (N_3520,In_1741,In_2406);
nor U3521 (N_3521,In_1301,In_1748);
nand U3522 (N_3522,In_1345,In_185);
nor U3523 (N_3523,In_164,In_883);
nor U3524 (N_3524,In_1077,In_525);
nand U3525 (N_3525,In_164,In_814);
nand U3526 (N_3526,In_215,In_76);
and U3527 (N_3527,In_239,In_788);
or U3528 (N_3528,In_2161,In_247);
and U3529 (N_3529,In_2305,In_1695);
nand U3530 (N_3530,In_927,In_968);
nor U3531 (N_3531,In_1954,In_582);
nand U3532 (N_3532,In_1345,In_980);
xor U3533 (N_3533,In_572,In_923);
nor U3534 (N_3534,In_1846,In_904);
or U3535 (N_3535,In_971,In_1127);
and U3536 (N_3536,In_1910,In_161);
or U3537 (N_3537,In_256,In_1307);
nand U3538 (N_3538,In_839,In_1169);
or U3539 (N_3539,In_1753,In_873);
nor U3540 (N_3540,In_1531,In_295);
and U3541 (N_3541,In_1570,In_2076);
nand U3542 (N_3542,In_1284,In_1682);
nand U3543 (N_3543,In_650,In_1614);
and U3544 (N_3544,In_1996,In_355);
nand U3545 (N_3545,In_1286,In_917);
nor U3546 (N_3546,In_1991,In_2032);
nor U3547 (N_3547,In_462,In_1471);
and U3548 (N_3548,In_1888,In_1128);
nand U3549 (N_3549,In_1490,In_349);
or U3550 (N_3550,In_1710,In_886);
nor U3551 (N_3551,In_168,In_2087);
and U3552 (N_3552,In_1115,In_1367);
and U3553 (N_3553,In_711,In_1365);
and U3554 (N_3554,In_2199,In_2091);
and U3555 (N_3555,In_69,In_115);
nor U3556 (N_3556,In_2110,In_1523);
and U3557 (N_3557,In_1887,In_2362);
and U3558 (N_3558,In_583,In_1245);
and U3559 (N_3559,In_1464,In_943);
nand U3560 (N_3560,In_1303,In_2486);
nor U3561 (N_3561,In_797,In_1066);
and U3562 (N_3562,In_457,In_928);
nand U3563 (N_3563,In_2293,In_1384);
nand U3564 (N_3564,In_278,In_1097);
or U3565 (N_3565,In_716,In_836);
or U3566 (N_3566,In_996,In_40);
and U3567 (N_3567,In_434,In_1306);
and U3568 (N_3568,In_2167,In_23);
or U3569 (N_3569,In_95,In_757);
nand U3570 (N_3570,In_2014,In_1863);
and U3571 (N_3571,In_805,In_1960);
or U3572 (N_3572,In_1185,In_1290);
and U3573 (N_3573,In_1441,In_162);
nand U3574 (N_3574,In_429,In_2435);
nor U3575 (N_3575,In_1845,In_261);
and U3576 (N_3576,In_651,In_2042);
nand U3577 (N_3577,In_444,In_1177);
nand U3578 (N_3578,In_1243,In_1939);
or U3579 (N_3579,In_2172,In_1107);
nor U3580 (N_3580,In_873,In_1255);
nor U3581 (N_3581,In_470,In_1800);
and U3582 (N_3582,In_194,In_2353);
and U3583 (N_3583,In_1254,In_1333);
nor U3584 (N_3584,In_429,In_1610);
xnor U3585 (N_3585,In_1489,In_2122);
xor U3586 (N_3586,In_1584,In_2258);
nor U3587 (N_3587,In_331,In_721);
nor U3588 (N_3588,In_872,In_2388);
nor U3589 (N_3589,In_663,In_1079);
or U3590 (N_3590,In_187,In_1715);
nand U3591 (N_3591,In_1016,In_557);
or U3592 (N_3592,In_430,In_2471);
nor U3593 (N_3593,In_661,In_839);
nor U3594 (N_3594,In_137,In_1017);
xnor U3595 (N_3595,In_1588,In_808);
nor U3596 (N_3596,In_75,In_1124);
nand U3597 (N_3597,In_298,In_1442);
nand U3598 (N_3598,In_213,In_1298);
or U3599 (N_3599,In_146,In_1011);
or U3600 (N_3600,In_1512,In_1539);
or U3601 (N_3601,In_1811,In_1283);
nor U3602 (N_3602,In_2483,In_50);
nor U3603 (N_3603,In_1323,In_1248);
and U3604 (N_3604,In_1742,In_1099);
or U3605 (N_3605,In_928,In_1064);
and U3606 (N_3606,In_854,In_1335);
nand U3607 (N_3607,In_1559,In_973);
nand U3608 (N_3608,In_1810,In_684);
and U3609 (N_3609,In_2488,In_456);
or U3610 (N_3610,In_1450,In_1542);
nand U3611 (N_3611,In_280,In_2445);
xor U3612 (N_3612,In_1836,In_30);
and U3613 (N_3613,In_35,In_1335);
or U3614 (N_3614,In_1146,In_739);
or U3615 (N_3615,In_41,In_2068);
xor U3616 (N_3616,In_137,In_2390);
or U3617 (N_3617,In_1207,In_1935);
nand U3618 (N_3618,In_478,In_24);
and U3619 (N_3619,In_1483,In_2295);
and U3620 (N_3620,In_2127,In_2053);
and U3621 (N_3621,In_593,In_897);
xnor U3622 (N_3622,In_13,In_1273);
or U3623 (N_3623,In_41,In_1188);
nand U3624 (N_3624,In_219,In_1661);
and U3625 (N_3625,In_1008,In_68);
and U3626 (N_3626,In_56,In_1085);
and U3627 (N_3627,In_207,In_1857);
and U3628 (N_3628,In_378,In_1702);
and U3629 (N_3629,In_2008,In_2361);
nand U3630 (N_3630,In_1705,In_1947);
and U3631 (N_3631,In_2450,In_21);
nand U3632 (N_3632,In_1831,In_825);
nor U3633 (N_3633,In_2284,In_361);
nor U3634 (N_3634,In_128,In_229);
nand U3635 (N_3635,In_753,In_17);
nor U3636 (N_3636,In_1854,In_1748);
and U3637 (N_3637,In_587,In_714);
and U3638 (N_3638,In_377,In_2185);
nand U3639 (N_3639,In_2421,In_910);
or U3640 (N_3640,In_750,In_229);
nor U3641 (N_3641,In_193,In_2235);
nor U3642 (N_3642,In_368,In_2182);
or U3643 (N_3643,In_1384,In_1312);
and U3644 (N_3644,In_1673,In_1847);
nand U3645 (N_3645,In_181,In_160);
nand U3646 (N_3646,In_975,In_2118);
or U3647 (N_3647,In_676,In_29);
nand U3648 (N_3648,In_1394,In_1507);
nand U3649 (N_3649,In_2145,In_2058);
or U3650 (N_3650,In_890,In_1833);
or U3651 (N_3651,In_2084,In_658);
and U3652 (N_3652,In_1226,In_719);
and U3653 (N_3653,In_548,In_1697);
or U3654 (N_3654,In_456,In_235);
nor U3655 (N_3655,In_2350,In_1979);
and U3656 (N_3656,In_19,In_2178);
xnor U3657 (N_3657,In_1547,In_642);
xor U3658 (N_3658,In_1886,In_1669);
nand U3659 (N_3659,In_80,In_1139);
and U3660 (N_3660,In_2167,In_894);
nor U3661 (N_3661,In_1550,In_58);
or U3662 (N_3662,In_2092,In_169);
and U3663 (N_3663,In_2435,In_1589);
and U3664 (N_3664,In_1686,In_1370);
and U3665 (N_3665,In_732,In_884);
nand U3666 (N_3666,In_341,In_103);
nor U3667 (N_3667,In_913,In_821);
and U3668 (N_3668,In_2264,In_1338);
and U3669 (N_3669,In_1914,In_181);
and U3670 (N_3670,In_326,In_662);
and U3671 (N_3671,In_1090,In_975);
or U3672 (N_3672,In_16,In_1712);
and U3673 (N_3673,In_208,In_796);
and U3674 (N_3674,In_1512,In_217);
nand U3675 (N_3675,In_1892,In_364);
nand U3676 (N_3676,In_64,In_878);
or U3677 (N_3677,In_1575,In_1874);
nor U3678 (N_3678,In_1958,In_663);
and U3679 (N_3679,In_257,In_2457);
nor U3680 (N_3680,In_64,In_845);
and U3681 (N_3681,In_5,In_1413);
and U3682 (N_3682,In_680,In_1731);
nor U3683 (N_3683,In_1754,In_2427);
or U3684 (N_3684,In_579,In_1461);
nor U3685 (N_3685,In_492,In_1275);
nand U3686 (N_3686,In_1061,In_386);
and U3687 (N_3687,In_42,In_1121);
nor U3688 (N_3688,In_744,In_453);
or U3689 (N_3689,In_229,In_1193);
nor U3690 (N_3690,In_1971,In_2432);
and U3691 (N_3691,In_186,In_2432);
xnor U3692 (N_3692,In_1218,In_2023);
nand U3693 (N_3693,In_560,In_860);
nor U3694 (N_3694,In_1952,In_1904);
and U3695 (N_3695,In_1579,In_361);
nor U3696 (N_3696,In_328,In_1885);
nand U3697 (N_3697,In_2022,In_1107);
or U3698 (N_3698,In_435,In_495);
or U3699 (N_3699,In_1747,In_1721);
and U3700 (N_3700,In_1975,In_871);
nand U3701 (N_3701,In_2211,In_1479);
nor U3702 (N_3702,In_2028,In_2074);
nor U3703 (N_3703,In_751,In_1985);
and U3704 (N_3704,In_1479,In_2290);
or U3705 (N_3705,In_2079,In_1239);
xnor U3706 (N_3706,In_271,In_987);
or U3707 (N_3707,In_581,In_1329);
nand U3708 (N_3708,In_660,In_1880);
nor U3709 (N_3709,In_1732,In_1343);
nand U3710 (N_3710,In_2061,In_1025);
nand U3711 (N_3711,In_1283,In_1595);
nand U3712 (N_3712,In_1126,In_520);
and U3713 (N_3713,In_67,In_493);
and U3714 (N_3714,In_2220,In_2186);
or U3715 (N_3715,In_387,In_97);
and U3716 (N_3716,In_1623,In_2305);
nand U3717 (N_3717,In_798,In_720);
nor U3718 (N_3718,In_1492,In_535);
nor U3719 (N_3719,In_1699,In_1713);
nor U3720 (N_3720,In_1416,In_2493);
and U3721 (N_3721,In_1621,In_1974);
nand U3722 (N_3722,In_687,In_1618);
nor U3723 (N_3723,In_122,In_1818);
and U3724 (N_3724,In_1538,In_2155);
nand U3725 (N_3725,In_1375,In_2377);
nand U3726 (N_3726,In_627,In_188);
nor U3727 (N_3727,In_190,In_2396);
nor U3728 (N_3728,In_1946,In_643);
or U3729 (N_3729,In_2225,In_1283);
and U3730 (N_3730,In_2325,In_1445);
nand U3731 (N_3731,In_802,In_32);
nor U3732 (N_3732,In_1928,In_1114);
nand U3733 (N_3733,In_1384,In_118);
or U3734 (N_3734,In_2287,In_1520);
nor U3735 (N_3735,In_2002,In_479);
and U3736 (N_3736,In_2185,In_965);
and U3737 (N_3737,In_873,In_1685);
nor U3738 (N_3738,In_889,In_1764);
xnor U3739 (N_3739,In_10,In_1365);
nor U3740 (N_3740,In_791,In_1425);
nand U3741 (N_3741,In_1266,In_572);
or U3742 (N_3742,In_386,In_1907);
nand U3743 (N_3743,In_1733,In_702);
nor U3744 (N_3744,In_1066,In_705);
nand U3745 (N_3745,In_205,In_1937);
and U3746 (N_3746,In_2053,In_2312);
nor U3747 (N_3747,In_942,In_497);
and U3748 (N_3748,In_2329,In_1369);
or U3749 (N_3749,In_762,In_344);
and U3750 (N_3750,In_2406,In_1400);
or U3751 (N_3751,In_142,In_1585);
xor U3752 (N_3752,In_2228,In_1963);
or U3753 (N_3753,In_2316,In_2192);
nor U3754 (N_3754,In_527,In_328);
or U3755 (N_3755,In_836,In_1141);
nor U3756 (N_3756,In_2109,In_2250);
nor U3757 (N_3757,In_4,In_2283);
and U3758 (N_3758,In_1213,In_109);
nor U3759 (N_3759,In_135,In_739);
nor U3760 (N_3760,In_2201,In_2347);
nand U3761 (N_3761,In_1456,In_2381);
and U3762 (N_3762,In_261,In_2467);
nand U3763 (N_3763,In_2445,In_219);
nor U3764 (N_3764,In_89,In_1146);
or U3765 (N_3765,In_1059,In_1614);
or U3766 (N_3766,In_1018,In_1550);
nor U3767 (N_3767,In_1739,In_420);
or U3768 (N_3768,In_968,In_2113);
nand U3769 (N_3769,In_1133,In_752);
or U3770 (N_3770,In_2002,In_1973);
nand U3771 (N_3771,In_719,In_330);
and U3772 (N_3772,In_2013,In_2080);
and U3773 (N_3773,In_2054,In_1432);
and U3774 (N_3774,In_21,In_513);
nand U3775 (N_3775,In_134,In_476);
nor U3776 (N_3776,In_1535,In_1582);
nor U3777 (N_3777,In_2159,In_719);
nand U3778 (N_3778,In_1514,In_2483);
nor U3779 (N_3779,In_1098,In_1984);
and U3780 (N_3780,In_908,In_142);
nand U3781 (N_3781,In_1145,In_1346);
or U3782 (N_3782,In_448,In_118);
or U3783 (N_3783,In_1508,In_2254);
nor U3784 (N_3784,In_1560,In_2385);
nor U3785 (N_3785,In_375,In_573);
nor U3786 (N_3786,In_1237,In_281);
or U3787 (N_3787,In_416,In_228);
or U3788 (N_3788,In_594,In_1457);
or U3789 (N_3789,In_2135,In_886);
nor U3790 (N_3790,In_1591,In_1056);
nand U3791 (N_3791,In_68,In_1244);
nand U3792 (N_3792,In_2382,In_2431);
or U3793 (N_3793,In_2247,In_295);
and U3794 (N_3794,In_1873,In_277);
and U3795 (N_3795,In_2465,In_1763);
or U3796 (N_3796,In_1795,In_143);
nor U3797 (N_3797,In_1092,In_1847);
or U3798 (N_3798,In_149,In_1588);
or U3799 (N_3799,In_1513,In_658);
or U3800 (N_3800,In_539,In_224);
nor U3801 (N_3801,In_2433,In_2358);
and U3802 (N_3802,In_2176,In_685);
nand U3803 (N_3803,In_578,In_892);
nand U3804 (N_3804,In_2130,In_32);
or U3805 (N_3805,In_1653,In_849);
or U3806 (N_3806,In_2282,In_1140);
or U3807 (N_3807,In_44,In_904);
nor U3808 (N_3808,In_1387,In_1008);
or U3809 (N_3809,In_1030,In_1125);
and U3810 (N_3810,In_428,In_1684);
or U3811 (N_3811,In_741,In_606);
nor U3812 (N_3812,In_1474,In_2371);
or U3813 (N_3813,In_1389,In_1777);
or U3814 (N_3814,In_2176,In_2115);
xnor U3815 (N_3815,In_1872,In_1893);
and U3816 (N_3816,In_1620,In_483);
nor U3817 (N_3817,In_21,In_1530);
nor U3818 (N_3818,In_632,In_504);
and U3819 (N_3819,In_61,In_1263);
nand U3820 (N_3820,In_1639,In_798);
nor U3821 (N_3821,In_744,In_804);
and U3822 (N_3822,In_310,In_1492);
nor U3823 (N_3823,In_2487,In_1087);
nand U3824 (N_3824,In_894,In_1059);
and U3825 (N_3825,In_810,In_1167);
and U3826 (N_3826,In_1033,In_754);
nor U3827 (N_3827,In_2411,In_873);
xor U3828 (N_3828,In_61,In_783);
or U3829 (N_3829,In_1830,In_582);
nor U3830 (N_3830,In_1287,In_494);
nand U3831 (N_3831,In_716,In_2152);
and U3832 (N_3832,In_1108,In_815);
nand U3833 (N_3833,In_1439,In_1364);
and U3834 (N_3834,In_145,In_1305);
xor U3835 (N_3835,In_2042,In_1171);
and U3836 (N_3836,In_942,In_1598);
nand U3837 (N_3837,In_990,In_2350);
nand U3838 (N_3838,In_650,In_733);
nor U3839 (N_3839,In_451,In_2225);
nor U3840 (N_3840,In_2142,In_908);
nor U3841 (N_3841,In_2374,In_768);
nand U3842 (N_3842,In_1153,In_1827);
or U3843 (N_3843,In_1476,In_1039);
or U3844 (N_3844,In_7,In_1830);
or U3845 (N_3845,In_1329,In_136);
xor U3846 (N_3846,In_1595,In_2112);
nor U3847 (N_3847,In_730,In_982);
nand U3848 (N_3848,In_120,In_2170);
nor U3849 (N_3849,In_2089,In_2349);
xnor U3850 (N_3850,In_1383,In_1454);
nor U3851 (N_3851,In_2344,In_2484);
nand U3852 (N_3852,In_947,In_357);
nor U3853 (N_3853,In_2155,In_1054);
and U3854 (N_3854,In_595,In_964);
nand U3855 (N_3855,In_2341,In_1933);
and U3856 (N_3856,In_1939,In_1904);
and U3857 (N_3857,In_2393,In_2237);
nor U3858 (N_3858,In_1817,In_1756);
nor U3859 (N_3859,In_626,In_881);
or U3860 (N_3860,In_917,In_177);
nand U3861 (N_3861,In_1206,In_1501);
and U3862 (N_3862,In_400,In_258);
nor U3863 (N_3863,In_1666,In_239);
and U3864 (N_3864,In_552,In_1879);
or U3865 (N_3865,In_2175,In_2102);
nand U3866 (N_3866,In_85,In_767);
nor U3867 (N_3867,In_2181,In_459);
or U3868 (N_3868,In_665,In_911);
nor U3869 (N_3869,In_1525,In_651);
nor U3870 (N_3870,In_2239,In_593);
and U3871 (N_3871,In_1938,In_2268);
or U3872 (N_3872,In_853,In_2119);
nand U3873 (N_3873,In_683,In_2061);
nor U3874 (N_3874,In_396,In_2056);
and U3875 (N_3875,In_485,In_2293);
and U3876 (N_3876,In_2487,In_965);
and U3877 (N_3877,In_1438,In_1368);
nor U3878 (N_3878,In_1685,In_1811);
or U3879 (N_3879,In_1336,In_1585);
or U3880 (N_3880,In_491,In_2301);
or U3881 (N_3881,In_75,In_1822);
nand U3882 (N_3882,In_2495,In_892);
or U3883 (N_3883,In_1599,In_937);
nand U3884 (N_3884,In_2335,In_1730);
or U3885 (N_3885,In_728,In_1446);
and U3886 (N_3886,In_1123,In_1311);
nand U3887 (N_3887,In_997,In_246);
and U3888 (N_3888,In_1637,In_1355);
nor U3889 (N_3889,In_289,In_1508);
nand U3890 (N_3890,In_824,In_1987);
nor U3891 (N_3891,In_889,In_1352);
nor U3892 (N_3892,In_1827,In_2381);
nand U3893 (N_3893,In_2011,In_694);
nand U3894 (N_3894,In_18,In_2459);
nand U3895 (N_3895,In_2211,In_879);
and U3896 (N_3896,In_1423,In_1441);
or U3897 (N_3897,In_670,In_815);
nor U3898 (N_3898,In_745,In_1940);
and U3899 (N_3899,In_1262,In_684);
nor U3900 (N_3900,In_848,In_888);
or U3901 (N_3901,In_851,In_1785);
nor U3902 (N_3902,In_2489,In_1733);
nor U3903 (N_3903,In_1601,In_2371);
and U3904 (N_3904,In_1278,In_191);
and U3905 (N_3905,In_1526,In_1458);
and U3906 (N_3906,In_775,In_1743);
nand U3907 (N_3907,In_223,In_933);
nand U3908 (N_3908,In_1882,In_130);
nand U3909 (N_3909,In_2268,In_1656);
and U3910 (N_3910,In_1243,In_2464);
nor U3911 (N_3911,In_467,In_2296);
nand U3912 (N_3912,In_841,In_1105);
and U3913 (N_3913,In_1257,In_1497);
and U3914 (N_3914,In_675,In_895);
nand U3915 (N_3915,In_241,In_2341);
nor U3916 (N_3916,In_269,In_1220);
nor U3917 (N_3917,In_1743,In_892);
or U3918 (N_3918,In_1690,In_1984);
or U3919 (N_3919,In_1621,In_2212);
or U3920 (N_3920,In_1410,In_768);
or U3921 (N_3921,In_52,In_214);
and U3922 (N_3922,In_1294,In_2229);
nor U3923 (N_3923,In_2183,In_1539);
and U3924 (N_3924,In_2036,In_188);
nor U3925 (N_3925,In_1664,In_2158);
nand U3926 (N_3926,In_2328,In_759);
nand U3927 (N_3927,In_1442,In_2315);
or U3928 (N_3928,In_1170,In_2364);
and U3929 (N_3929,In_272,In_1760);
and U3930 (N_3930,In_2490,In_614);
or U3931 (N_3931,In_1558,In_809);
xor U3932 (N_3932,In_2260,In_39);
or U3933 (N_3933,In_136,In_2219);
nand U3934 (N_3934,In_1850,In_1922);
nor U3935 (N_3935,In_760,In_922);
and U3936 (N_3936,In_2334,In_561);
and U3937 (N_3937,In_2129,In_1009);
and U3938 (N_3938,In_1627,In_1748);
and U3939 (N_3939,In_1503,In_765);
nor U3940 (N_3940,In_1063,In_2045);
and U3941 (N_3941,In_1653,In_26);
nor U3942 (N_3942,In_2490,In_1340);
nor U3943 (N_3943,In_614,In_2228);
xnor U3944 (N_3944,In_2473,In_2283);
and U3945 (N_3945,In_1216,In_73);
and U3946 (N_3946,In_1621,In_493);
and U3947 (N_3947,In_2241,In_133);
and U3948 (N_3948,In_2362,In_2260);
nor U3949 (N_3949,In_2351,In_1484);
and U3950 (N_3950,In_1107,In_2084);
nor U3951 (N_3951,In_2282,In_1211);
or U3952 (N_3952,In_2136,In_1135);
nand U3953 (N_3953,In_1891,In_1021);
nand U3954 (N_3954,In_1834,In_2296);
or U3955 (N_3955,In_1231,In_1381);
nor U3956 (N_3956,In_1550,In_1422);
or U3957 (N_3957,In_1216,In_681);
nor U3958 (N_3958,In_2487,In_2038);
nor U3959 (N_3959,In_1242,In_1761);
and U3960 (N_3960,In_118,In_1578);
nand U3961 (N_3961,In_1255,In_1861);
and U3962 (N_3962,In_2138,In_1821);
nand U3963 (N_3963,In_648,In_2033);
nand U3964 (N_3964,In_2128,In_2179);
nor U3965 (N_3965,In_1551,In_623);
or U3966 (N_3966,In_1270,In_948);
and U3967 (N_3967,In_631,In_380);
or U3968 (N_3968,In_1029,In_1322);
nor U3969 (N_3969,In_63,In_2292);
xor U3970 (N_3970,In_2494,In_1167);
and U3971 (N_3971,In_2303,In_2089);
and U3972 (N_3972,In_1170,In_843);
or U3973 (N_3973,In_2154,In_2212);
nand U3974 (N_3974,In_28,In_617);
nor U3975 (N_3975,In_502,In_337);
nor U3976 (N_3976,In_1315,In_734);
nand U3977 (N_3977,In_1341,In_9);
and U3978 (N_3978,In_290,In_2297);
xnor U3979 (N_3979,In_704,In_1215);
nand U3980 (N_3980,In_329,In_300);
nor U3981 (N_3981,In_473,In_921);
nor U3982 (N_3982,In_771,In_2244);
or U3983 (N_3983,In_1885,In_2277);
nor U3984 (N_3984,In_383,In_2010);
xor U3985 (N_3985,In_2010,In_34);
nor U3986 (N_3986,In_652,In_1072);
or U3987 (N_3987,In_2139,In_136);
nand U3988 (N_3988,In_1978,In_911);
or U3989 (N_3989,In_35,In_1183);
and U3990 (N_3990,In_624,In_1584);
nor U3991 (N_3991,In_1923,In_492);
and U3992 (N_3992,In_854,In_1587);
or U3993 (N_3993,In_1404,In_1256);
or U3994 (N_3994,In_170,In_1051);
or U3995 (N_3995,In_130,In_2176);
nand U3996 (N_3996,In_672,In_616);
nor U3997 (N_3997,In_1158,In_2012);
nand U3998 (N_3998,In_547,In_2490);
or U3999 (N_3999,In_363,In_1128);
and U4000 (N_4000,In_1411,In_1636);
or U4001 (N_4001,In_1798,In_460);
or U4002 (N_4002,In_1371,In_1767);
and U4003 (N_4003,In_250,In_2420);
and U4004 (N_4004,In_2438,In_1663);
or U4005 (N_4005,In_1387,In_1513);
and U4006 (N_4006,In_1781,In_764);
and U4007 (N_4007,In_1029,In_2039);
nor U4008 (N_4008,In_584,In_340);
nor U4009 (N_4009,In_2191,In_1703);
and U4010 (N_4010,In_2051,In_1185);
and U4011 (N_4011,In_2063,In_2196);
and U4012 (N_4012,In_1682,In_1993);
nand U4013 (N_4013,In_628,In_2270);
nand U4014 (N_4014,In_1276,In_204);
or U4015 (N_4015,In_1443,In_2210);
or U4016 (N_4016,In_1390,In_1075);
and U4017 (N_4017,In_2159,In_1312);
or U4018 (N_4018,In_582,In_870);
nor U4019 (N_4019,In_1074,In_1584);
and U4020 (N_4020,In_249,In_1174);
and U4021 (N_4021,In_1856,In_997);
nand U4022 (N_4022,In_1050,In_1097);
and U4023 (N_4023,In_956,In_2063);
or U4024 (N_4024,In_271,In_352);
nor U4025 (N_4025,In_1065,In_744);
nor U4026 (N_4026,In_2047,In_1747);
nand U4027 (N_4027,In_798,In_572);
xor U4028 (N_4028,In_1813,In_1518);
nand U4029 (N_4029,In_1493,In_347);
nor U4030 (N_4030,In_70,In_2484);
and U4031 (N_4031,In_2118,In_1039);
and U4032 (N_4032,In_1017,In_1746);
and U4033 (N_4033,In_831,In_1600);
or U4034 (N_4034,In_1096,In_1460);
or U4035 (N_4035,In_245,In_1555);
nand U4036 (N_4036,In_1401,In_445);
or U4037 (N_4037,In_657,In_102);
and U4038 (N_4038,In_332,In_2354);
nand U4039 (N_4039,In_265,In_745);
nor U4040 (N_4040,In_2211,In_247);
and U4041 (N_4041,In_298,In_941);
or U4042 (N_4042,In_1540,In_1625);
or U4043 (N_4043,In_286,In_693);
nand U4044 (N_4044,In_1493,In_1910);
nand U4045 (N_4045,In_1903,In_427);
nor U4046 (N_4046,In_230,In_1001);
or U4047 (N_4047,In_91,In_2252);
nand U4048 (N_4048,In_1428,In_569);
nand U4049 (N_4049,In_2413,In_235);
and U4050 (N_4050,In_492,In_263);
nor U4051 (N_4051,In_2193,In_960);
or U4052 (N_4052,In_1591,In_66);
nor U4053 (N_4053,In_1580,In_1864);
nand U4054 (N_4054,In_160,In_2290);
nand U4055 (N_4055,In_1346,In_1136);
nor U4056 (N_4056,In_1195,In_1478);
nand U4057 (N_4057,In_1460,In_1589);
and U4058 (N_4058,In_188,In_535);
nor U4059 (N_4059,In_2230,In_1152);
nor U4060 (N_4060,In_448,In_1986);
and U4061 (N_4061,In_2241,In_492);
or U4062 (N_4062,In_1902,In_1299);
nand U4063 (N_4063,In_2482,In_1515);
nor U4064 (N_4064,In_46,In_2071);
and U4065 (N_4065,In_2240,In_1812);
and U4066 (N_4066,In_111,In_1618);
or U4067 (N_4067,In_891,In_1925);
and U4068 (N_4068,In_282,In_194);
nor U4069 (N_4069,In_1600,In_772);
or U4070 (N_4070,In_1869,In_1171);
nand U4071 (N_4071,In_238,In_249);
and U4072 (N_4072,In_2467,In_744);
nand U4073 (N_4073,In_1442,In_2230);
nor U4074 (N_4074,In_2063,In_1725);
nor U4075 (N_4075,In_523,In_2165);
nand U4076 (N_4076,In_49,In_468);
nand U4077 (N_4077,In_503,In_6);
or U4078 (N_4078,In_2368,In_1675);
or U4079 (N_4079,In_636,In_23);
nand U4080 (N_4080,In_1107,In_2238);
nand U4081 (N_4081,In_2363,In_2361);
nand U4082 (N_4082,In_2490,In_448);
nor U4083 (N_4083,In_796,In_1401);
or U4084 (N_4084,In_470,In_948);
and U4085 (N_4085,In_145,In_2006);
xnor U4086 (N_4086,In_491,In_2412);
and U4087 (N_4087,In_1167,In_927);
nand U4088 (N_4088,In_551,In_1124);
nand U4089 (N_4089,In_430,In_1966);
nand U4090 (N_4090,In_1666,In_454);
nor U4091 (N_4091,In_486,In_2378);
nor U4092 (N_4092,In_1716,In_2192);
nor U4093 (N_4093,In_100,In_1072);
nand U4094 (N_4094,In_612,In_780);
nand U4095 (N_4095,In_438,In_1558);
nand U4096 (N_4096,In_100,In_1193);
and U4097 (N_4097,In_656,In_349);
nand U4098 (N_4098,In_161,In_1824);
or U4099 (N_4099,In_2017,In_34);
nor U4100 (N_4100,In_315,In_1445);
nor U4101 (N_4101,In_215,In_2236);
and U4102 (N_4102,In_1753,In_2394);
nand U4103 (N_4103,In_2284,In_2184);
and U4104 (N_4104,In_418,In_1728);
and U4105 (N_4105,In_1274,In_2130);
and U4106 (N_4106,In_2164,In_2079);
nor U4107 (N_4107,In_1810,In_978);
nor U4108 (N_4108,In_1742,In_1869);
or U4109 (N_4109,In_311,In_2263);
or U4110 (N_4110,In_1160,In_1757);
or U4111 (N_4111,In_1434,In_1676);
nand U4112 (N_4112,In_2235,In_1451);
and U4113 (N_4113,In_1978,In_1161);
and U4114 (N_4114,In_489,In_637);
nand U4115 (N_4115,In_171,In_974);
or U4116 (N_4116,In_2348,In_386);
and U4117 (N_4117,In_2141,In_212);
nor U4118 (N_4118,In_1470,In_1065);
or U4119 (N_4119,In_662,In_1429);
nand U4120 (N_4120,In_323,In_1658);
nor U4121 (N_4121,In_2181,In_1018);
nor U4122 (N_4122,In_1843,In_1765);
or U4123 (N_4123,In_1839,In_1448);
or U4124 (N_4124,In_253,In_1622);
or U4125 (N_4125,In_946,In_274);
or U4126 (N_4126,In_25,In_868);
or U4127 (N_4127,In_902,In_2127);
and U4128 (N_4128,In_1499,In_2433);
or U4129 (N_4129,In_1753,In_1568);
nor U4130 (N_4130,In_1360,In_2124);
and U4131 (N_4131,In_2029,In_243);
and U4132 (N_4132,In_477,In_1432);
nand U4133 (N_4133,In_2479,In_1214);
or U4134 (N_4134,In_2123,In_1592);
xor U4135 (N_4135,In_2388,In_1891);
xor U4136 (N_4136,In_1600,In_2069);
or U4137 (N_4137,In_2350,In_332);
nor U4138 (N_4138,In_153,In_1184);
or U4139 (N_4139,In_1592,In_890);
and U4140 (N_4140,In_1419,In_1348);
or U4141 (N_4141,In_1303,In_1266);
and U4142 (N_4142,In_273,In_544);
nor U4143 (N_4143,In_770,In_1080);
nand U4144 (N_4144,In_35,In_956);
or U4145 (N_4145,In_87,In_864);
nor U4146 (N_4146,In_1099,In_455);
nor U4147 (N_4147,In_272,In_1335);
or U4148 (N_4148,In_1223,In_1732);
nor U4149 (N_4149,In_518,In_428);
or U4150 (N_4150,In_2024,In_1390);
nor U4151 (N_4151,In_709,In_211);
or U4152 (N_4152,In_2182,In_904);
and U4153 (N_4153,In_2161,In_714);
nand U4154 (N_4154,In_1226,In_1141);
nor U4155 (N_4155,In_1721,In_509);
or U4156 (N_4156,In_1838,In_1827);
nor U4157 (N_4157,In_594,In_1895);
and U4158 (N_4158,In_1893,In_438);
xor U4159 (N_4159,In_546,In_17);
or U4160 (N_4160,In_498,In_2156);
nor U4161 (N_4161,In_2004,In_1112);
and U4162 (N_4162,In_853,In_2225);
or U4163 (N_4163,In_67,In_245);
nor U4164 (N_4164,In_1126,In_318);
nand U4165 (N_4165,In_922,In_1320);
or U4166 (N_4166,In_156,In_789);
nor U4167 (N_4167,In_606,In_541);
and U4168 (N_4168,In_2435,In_2094);
and U4169 (N_4169,In_1746,In_1827);
and U4170 (N_4170,In_98,In_249);
or U4171 (N_4171,In_271,In_1853);
nand U4172 (N_4172,In_130,In_66);
or U4173 (N_4173,In_1341,In_1464);
or U4174 (N_4174,In_1669,In_1821);
or U4175 (N_4175,In_838,In_1382);
nand U4176 (N_4176,In_601,In_774);
or U4177 (N_4177,In_1871,In_2474);
or U4178 (N_4178,In_2009,In_655);
nand U4179 (N_4179,In_551,In_208);
nand U4180 (N_4180,In_1509,In_658);
and U4181 (N_4181,In_918,In_1361);
nand U4182 (N_4182,In_387,In_1791);
nor U4183 (N_4183,In_163,In_1568);
or U4184 (N_4184,In_1682,In_1329);
nor U4185 (N_4185,In_1583,In_545);
nor U4186 (N_4186,In_399,In_1893);
nand U4187 (N_4187,In_703,In_1948);
and U4188 (N_4188,In_1567,In_1917);
or U4189 (N_4189,In_2462,In_1841);
nand U4190 (N_4190,In_306,In_1342);
nand U4191 (N_4191,In_21,In_802);
nor U4192 (N_4192,In_2407,In_520);
and U4193 (N_4193,In_886,In_88);
nand U4194 (N_4194,In_1585,In_1580);
or U4195 (N_4195,In_286,In_991);
nand U4196 (N_4196,In_963,In_1619);
nor U4197 (N_4197,In_1617,In_98);
and U4198 (N_4198,In_420,In_1865);
nor U4199 (N_4199,In_2310,In_1872);
and U4200 (N_4200,In_52,In_2396);
nor U4201 (N_4201,In_1773,In_2341);
and U4202 (N_4202,In_182,In_1197);
and U4203 (N_4203,In_824,In_1195);
and U4204 (N_4204,In_506,In_1825);
and U4205 (N_4205,In_2284,In_1312);
nand U4206 (N_4206,In_788,In_227);
nor U4207 (N_4207,In_926,In_1274);
and U4208 (N_4208,In_2495,In_1923);
nand U4209 (N_4209,In_181,In_1296);
nand U4210 (N_4210,In_672,In_2312);
nand U4211 (N_4211,In_565,In_1064);
and U4212 (N_4212,In_2430,In_350);
and U4213 (N_4213,In_133,In_409);
nand U4214 (N_4214,In_2393,In_1408);
or U4215 (N_4215,In_599,In_1496);
and U4216 (N_4216,In_111,In_1691);
and U4217 (N_4217,In_1513,In_1546);
xnor U4218 (N_4218,In_209,In_1923);
or U4219 (N_4219,In_1994,In_1594);
and U4220 (N_4220,In_1940,In_163);
nand U4221 (N_4221,In_400,In_752);
or U4222 (N_4222,In_1028,In_1652);
nand U4223 (N_4223,In_1549,In_1559);
nor U4224 (N_4224,In_1020,In_392);
and U4225 (N_4225,In_350,In_776);
nand U4226 (N_4226,In_1170,In_1019);
xor U4227 (N_4227,In_454,In_2412);
nand U4228 (N_4228,In_626,In_1519);
or U4229 (N_4229,In_1765,In_2475);
xor U4230 (N_4230,In_1915,In_1972);
and U4231 (N_4231,In_183,In_2322);
and U4232 (N_4232,In_662,In_2483);
or U4233 (N_4233,In_731,In_1356);
nor U4234 (N_4234,In_2453,In_465);
and U4235 (N_4235,In_1811,In_1450);
nand U4236 (N_4236,In_834,In_80);
and U4237 (N_4237,In_385,In_460);
nand U4238 (N_4238,In_589,In_1397);
nor U4239 (N_4239,In_1907,In_421);
nor U4240 (N_4240,In_1617,In_2106);
and U4241 (N_4241,In_668,In_68);
or U4242 (N_4242,In_236,In_872);
nand U4243 (N_4243,In_1397,In_106);
and U4244 (N_4244,In_371,In_1748);
or U4245 (N_4245,In_1001,In_1220);
xnor U4246 (N_4246,In_456,In_179);
nor U4247 (N_4247,In_1367,In_1844);
nor U4248 (N_4248,In_76,In_1310);
xnor U4249 (N_4249,In_1912,In_509);
nor U4250 (N_4250,In_2392,In_2339);
or U4251 (N_4251,In_1956,In_738);
and U4252 (N_4252,In_2066,In_2006);
nor U4253 (N_4253,In_715,In_254);
and U4254 (N_4254,In_990,In_1676);
and U4255 (N_4255,In_1740,In_2273);
or U4256 (N_4256,In_221,In_1226);
and U4257 (N_4257,In_925,In_1574);
nand U4258 (N_4258,In_461,In_668);
nor U4259 (N_4259,In_446,In_1756);
and U4260 (N_4260,In_123,In_681);
and U4261 (N_4261,In_611,In_44);
and U4262 (N_4262,In_974,In_1041);
and U4263 (N_4263,In_1930,In_495);
and U4264 (N_4264,In_2257,In_1367);
and U4265 (N_4265,In_1279,In_1295);
nand U4266 (N_4266,In_671,In_1826);
nand U4267 (N_4267,In_208,In_583);
and U4268 (N_4268,In_129,In_859);
and U4269 (N_4269,In_82,In_1166);
nand U4270 (N_4270,In_1204,In_158);
nand U4271 (N_4271,In_651,In_1297);
nor U4272 (N_4272,In_1138,In_750);
nor U4273 (N_4273,In_1148,In_1580);
and U4274 (N_4274,In_117,In_2136);
or U4275 (N_4275,In_1264,In_20);
or U4276 (N_4276,In_1799,In_1860);
nor U4277 (N_4277,In_78,In_2208);
nor U4278 (N_4278,In_42,In_2337);
nand U4279 (N_4279,In_1165,In_761);
and U4280 (N_4280,In_1096,In_468);
and U4281 (N_4281,In_300,In_984);
nor U4282 (N_4282,In_1285,In_1894);
or U4283 (N_4283,In_2005,In_2436);
nand U4284 (N_4284,In_1066,In_1217);
nor U4285 (N_4285,In_663,In_1085);
and U4286 (N_4286,In_639,In_875);
nand U4287 (N_4287,In_1514,In_140);
nand U4288 (N_4288,In_856,In_2365);
or U4289 (N_4289,In_1340,In_2143);
nor U4290 (N_4290,In_2278,In_2378);
or U4291 (N_4291,In_1621,In_1454);
nor U4292 (N_4292,In_919,In_1154);
and U4293 (N_4293,In_2179,In_736);
or U4294 (N_4294,In_192,In_69);
nor U4295 (N_4295,In_925,In_1954);
and U4296 (N_4296,In_177,In_709);
nor U4297 (N_4297,In_143,In_2432);
or U4298 (N_4298,In_1126,In_1584);
nand U4299 (N_4299,In_1994,In_1727);
nor U4300 (N_4300,In_428,In_124);
nor U4301 (N_4301,In_1854,In_1145);
nor U4302 (N_4302,In_156,In_2257);
nand U4303 (N_4303,In_2313,In_1821);
nand U4304 (N_4304,In_354,In_681);
and U4305 (N_4305,In_549,In_784);
nor U4306 (N_4306,In_1941,In_1723);
and U4307 (N_4307,In_1533,In_1748);
nand U4308 (N_4308,In_1906,In_2334);
and U4309 (N_4309,In_1133,In_1704);
or U4310 (N_4310,In_2161,In_20);
and U4311 (N_4311,In_1699,In_1336);
nand U4312 (N_4312,In_2027,In_2264);
nand U4313 (N_4313,In_1061,In_1600);
nor U4314 (N_4314,In_118,In_1747);
nand U4315 (N_4315,In_1325,In_1687);
xnor U4316 (N_4316,In_1139,In_979);
nand U4317 (N_4317,In_274,In_2316);
nand U4318 (N_4318,In_866,In_2034);
and U4319 (N_4319,In_959,In_757);
nand U4320 (N_4320,In_651,In_1382);
and U4321 (N_4321,In_269,In_2163);
nor U4322 (N_4322,In_2160,In_1484);
nand U4323 (N_4323,In_1492,In_2446);
nand U4324 (N_4324,In_999,In_1321);
and U4325 (N_4325,In_684,In_1721);
and U4326 (N_4326,In_1669,In_873);
nand U4327 (N_4327,In_1273,In_1484);
nand U4328 (N_4328,In_1632,In_532);
or U4329 (N_4329,In_1391,In_604);
and U4330 (N_4330,In_1732,In_377);
or U4331 (N_4331,In_304,In_1857);
nor U4332 (N_4332,In_902,In_597);
nand U4333 (N_4333,In_1729,In_2396);
and U4334 (N_4334,In_2174,In_2194);
or U4335 (N_4335,In_579,In_1102);
or U4336 (N_4336,In_739,In_396);
nand U4337 (N_4337,In_1965,In_1222);
and U4338 (N_4338,In_1440,In_10);
xnor U4339 (N_4339,In_1601,In_876);
nor U4340 (N_4340,In_238,In_148);
nor U4341 (N_4341,In_670,In_1010);
and U4342 (N_4342,In_1612,In_477);
or U4343 (N_4343,In_1654,In_1828);
nand U4344 (N_4344,In_228,In_845);
nand U4345 (N_4345,In_1819,In_1716);
nand U4346 (N_4346,In_2111,In_348);
or U4347 (N_4347,In_1463,In_2234);
and U4348 (N_4348,In_511,In_621);
or U4349 (N_4349,In_1989,In_2303);
nand U4350 (N_4350,In_1506,In_479);
or U4351 (N_4351,In_1401,In_1775);
nor U4352 (N_4352,In_1340,In_1103);
and U4353 (N_4353,In_344,In_2027);
or U4354 (N_4354,In_1596,In_2060);
nand U4355 (N_4355,In_1561,In_1127);
and U4356 (N_4356,In_1866,In_1864);
nor U4357 (N_4357,In_1335,In_2433);
or U4358 (N_4358,In_2083,In_2145);
and U4359 (N_4359,In_2034,In_353);
nor U4360 (N_4360,In_1127,In_840);
and U4361 (N_4361,In_2020,In_1528);
nand U4362 (N_4362,In_47,In_1414);
nor U4363 (N_4363,In_1246,In_2457);
or U4364 (N_4364,In_181,In_2295);
nor U4365 (N_4365,In_1874,In_576);
nand U4366 (N_4366,In_1773,In_2193);
and U4367 (N_4367,In_2170,In_2352);
nor U4368 (N_4368,In_500,In_1864);
and U4369 (N_4369,In_1099,In_703);
nor U4370 (N_4370,In_1223,In_289);
or U4371 (N_4371,In_1073,In_691);
nor U4372 (N_4372,In_1820,In_1618);
nor U4373 (N_4373,In_2398,In_549);
nand U4374 (N_4374,In_1660,In_1604);
nand U4375 (N_4375,In_2419,In_399);
nand U4376 (N_4376,In_1526,In_2313);
nand U4377 (N_4377,In_1507,In_1447);
nand U4378 (N_4378,In_1999,In_2357);
xor U4379 (N_4379,In_2148,In_1464);
or U4380 (N_4380,In_473,In_2311);
nand U4381 (N_4381,In_2165,In_1071);
nor U4382 (N_4382,In_1083,In_916);
or U4383 (N_4383,In_1428,In_19);
nor U4384 (N_4384,In_1407,In_248);
or U4385 (N_4385,In_1954,In_1441);
nor U4386 (N_4386,In_2450,In_1057);
nor U4387 (N_4387,In_1629,In_2299);
or U4388 (N_4388,In_164,In_1831);
nand U4389 (N_4389,In_6,In_867);
nor U4390 (N_4390,In_1653,In_2124);
and U4391 (N_4391,In_325,In_1168);
or U4392 (N_4392,In_597,In_514);
nand U4393 (N_4393,In_1438,In_706);
nor U4394 (N_4394,In_120,In_866);
xor U4395 (N_4395,In_322,In_471);
nor U4396 (N_4396,In_184,In_2091);
or U4397 (N_4397,In_1276,In_416);
nand U4398 (N_4398,In_2255,In_1341);
or U4399 (N_4399,In_282,In_339);
and U4400 (N_4400,In_242,In_756);
nor U4401 (N_4401,In_990,In_1706);
or U4402 (N_4402,In_824,In_2298);
and U4403 (N_4403,In_500,In_1626);
and U4404 (N_4404,In_1352,In_994);
or U4405 (N_4405,In_960,In_2042);
and U4406 (N_4406,In_1912,In_399);
or U4407 (N_4407,In_1805,In_1641);
or U4408 (N_4408,In_1640,In_854);
and U4409 (N_4409,In_1757,In_1017);
nand U4410 (N_4410,In_1086,In_1893);
or U4411 (N_4411,In_1378,In_166);
nor U4412 (N_4412,In_1737,In_1931);
or U4413 (N_4413,In_56,In_1488);
or U4414 (N_4414,In_1886,In_2135);
and U4415 (N_4415,In_1653,In_2199);
xnor U4416 (N_4416,In_2239,In_2002);
nor U4417 (N_4417,In_1554,In_508);
nand U4418 (N_4418,In_1741,In_2241);
and U4419 (N_4419,In_2141,In_1562);
and U4420 (N_4420,In_1961,In_1377);
nor U4421 (N_4421,In_2245,In_1348);
and U4422 (N_4422,In_0,In_1029);
nor U4423 (N_4423,In_814,In_865);
nor U4424 (N_4424,In_41,In_1544);
nor U4425 (N_4425,In_180,In_866);
and U4426 (N_4426,In_1790,In_948);
and U4427 (N_4427,In_1079,In_1147);
nor U4428 (N_4428,In_2421,In_1720);
nand U4429 (N_4429,In_1173,In_162);
nand U4430 (N_4430,In_270,In_2400);
and U4431 (N_4431,In_1008,In_1863);
or U4432 (N_4432,In_850,In_2368);
or U4433 (N_4433,In_1034,In_605);
or U4434 (N_4434,In_1450,In_922);
or U4435 (N_4435,In_2072,In_180);
and U4436 (N_4436,In_1281,In_1398);
and U4437 (N_4437,In_549,In_768);
or U4438 (N_4438,In_1596,In_2147);
and U4439 (N_4439,In_761,In_97);
or U4440 (N_4440,In_1702,In_2100);
xor U4441 (N_4441,In_2453,In_1763);
xnor U4442 (N_4442,In_1398,In_2468);
or U4443 (N_4443,In_308,In_1566);
nand U4444 (N_4444,In_1303,In_1729);
nand U4445 (N_4445,In_188,In_683);
or U4446 (N_4446,In_2114,In_536);
nor U4447 (N_4447,In_1060,In_1931);
nand U4448 (N_4448,In_159,In_1659);
nand U4449 (N_4449,In_70,In_808);
nand U4450 (N_4450,In_2192,In_200);
or U4451 (N_4451,In_1224,In_1903);
nor U4452 (N_4452,In_1379,In_966);
or U4453 (N_4453,In_1477,In_938);
nor U4454 (N_4454,In_1860,In_300);
nor U4455 (N_4455,In_2057,In_706);
and U4456 (N_4456,In_1317,In_1261);
nor U4457 (N_4457,In_781,In_227);
and U4458 (N_4458,In_189,In_1352);
nor U4459 (N_4459,In_762,In_76);
and U4460 (N_4460,In_1507,In_1107);
and U4461 (N_4461,In_302,In_286);
or U4462 (N_4462,In_2298,In_198);
nand U4463 (N_4463,In_208,In_1176);
xnor U4464 (N_4464,In_1740,In_970);
xor U4465 (N_4465,In_1065,In_107);
nand U4466 (N_4466,In_2031,In_2271);
nand U4467 (N_4467,In_1257,In_382);
or U4468 (N_4468,In_278,In_1307);
nor U4469 (N_4469,In_1954,In_2335);
or U4470 (N_4470,In_858,In_1224);
or U4471 (N_4471,In_2332,In_1057);
and U4472 (N_4472,In_2302,In_1424);
and U4473 (N_4473,In_482,In_1263);
or U4474 (N_4474,In_215,In_1980);
nand U4475 (N_4475,In_658,In_1550);
nor U4476 (N_4476,In_1300,In_1961);
or U4477 (N_4477,In_2188,In_1455);
nor U4478 (N_4478,In_1248,In_5);
nand U4479 (N_4479,In_1943,In_2239);
nor U4480 (N_4480,In_2484,In_438);
or U4481 (N_4481,In_123,In_1259);
and U4482 (N_4482,In_2122,In_563);
nand U4483 (N_4483,In_802,In_265);
nor U4484 (N_4484,In_861,In_1129);
or U4485 (N_4485,In_1026,In_1841);
nand U4486 (N_4486,In_693,In_1762);
and U4487 (N_4487,In_2323,In_1826);
and U4488 (N_4488,In_1711,In_1080);
nand U4489 (N_4489,In_63,In_1063);
and U4490 (N_4490,In_874,In_106);
or U4491 (N_4491,In_2319,In_53);
and U4492 (N_4492,In_437,In_549);
and U4493 (N_4493,In_1153,In_1320);
nand U4494 (N_4494,In_1630,In_1399);
nand U4495 (N_4495,In_1522,In_2314);
xor U4496 (N_4496,In_1297,In_2135);
nand U4497 (N_4497,In_1546,In_47);
nor U4498 (N_4498,In_993,In_1634);
nor U4499 (N_4499,In_2317,In_1018);
and U4500 (N_4500,In_1751,In_733);
xnor U4501 (N_4501,In_1214,In_82);
nand U4502 (N_4502,In_1790,In_2166);
or U4503 (N_4503,In_2198,In_500);
and U4504 (N_4504,In_962,In_2113);
nand U4505 (N_4505,In_1197,In_792);
or U4506 (N_4506,In_1505,In_539);
nand U4507 (N_4507,In_882,In_1057);
nor U4508 (N_4508,In_2020,In_2407);
nor U4509 (N_4509,In_35,In_915);
nor U4510 (N_4510,In_282,In_97);
or U4511 (N_4511,In_422,In_720);
or U4512 (N_4512,In_62,In_780);
nor U4513 (N_4513,In_2159,In_2226);
nor U4514 (N_4514,In_1462,In_2066);
or U4515 (N_4515,In_2263,In_1382);
nand U4516 (N_4516,In_1528,In_854);
or U4517 (N_4517,In_1921,In_1642);
nor U4518 (N_4518,In_2451,In_459);
and U4519 (N_4519,In_1572,In_1186);
nor U4520 (N_4520,In_1692,In_2305);
or U4521 (N_4521,In_1294,In_970);
nand U4522 (N_4522,In_1747,In_1276);
nand U4523 (N_4523,In_1782,In_2279);
or U4524 (N_4524,In_617,In_763);
nor U4525 (N_4525,In_557,In_77);
nor U4526 (N_4526,In_1611,In_2361);
and U4527 (N_4527,In_1475,In_2451);
and U4528 (N_4528,In_165,In_2092);
and U4529 (N_4529,In_2173,In_112);
nand U4530 (N_4530,In_1181,In_2377);
and U4531 (N_4531,In_2016,In_37);
or U4532 (N_4532,In_1452,In_579);
or U4533 (N_4533,In_2290,In_1808);
nor U4534 (N_4534,In_913,In_413);
xor U4535 (N_4535,In_1834,In_2112);
nand U4536 (N_4536,In_633,In_1166);
nand U4537 (N_4537,In_2473,In_1155);
and U4538 (N_4538,In_324,In_985);
nand U4539 (N_4539,In_1500,In_1258);
nand U4540 (N_4540,In_705,In_574);
nand U4541 (N_4541,In_2285,In_717);
or U4542 (N_4542,In_1027,In_749);
and U4543 (N_4543,In_2219,In_182);
nand U4544 (N_4544,In_2247,In_226);
xnor U4545 (N_4545,In_1973,In_93);
nand U4546 (N_4546,In_32,In_331);
or U4547 (N_4547,In_736,In_787);
nor U4548 (N_4548,In_649,In_333);
or U4549 (N_4549,In_1620,In_1878);
nand U4550 (N_4550,In_1946,In_2407);
nor U4551 (N_4551,In_1929,In_111);
and U4552 (N_4552,In_163,In_2198);
nand U4553 (N_4553,In_157,In_355);
and U4554 (N_4554,In_2125,In_2345);
nand U4555 (N_4555,In_2188,In_1010);
nor U4556 (N_4556,In_538,In_438);
and U4557 (N_4557,In_2163,In_1313);
or U4558 (N_4558,In_2090,In_1408);
or U4559 (N_4559,In_839,In_2390);
and U4560 (N_4560,In_2224,In_522);
nand U4561 (N_4561,In_1524,In_445);
nand U4562 (N_4562,In_802,In_1593);
or U4563 (N_4563,In_1975,In_1466);
or U4564 (N_4564,In_240,In_1121);
nor U4565 (N_4565,In_939,In_354);
or U4566 (N_4566,In_827,In_1310);
or U4567 (N_4567,In_1881,In_2044);
or U4568 (N_4568,In_1342,In_2235);
xor U4569 (N_4569,In_1341,In_594);
or U4570 (N_4570,In_1115,In_1996);
and U4571 (N_4571,In_63,In_1820);
nand U4572 (N_4572,In_1691,In_429);
nor U4573 (N_4573,In_2493,In_455);
or U4574 (N_4574,In_2425,In_1642);
nand U4575 (N_4575,In_2461,In_1366);
nor U4576 (N_4576,In_2251,In_1716);
nor U4577 (N_4577,In_429,In_124);
or U4578 (N_4578,In_745,In_2266);
and U4579 (N_4579,In_1103,In_2044);
and U4580 (N_4580,In_273,In_777);
nand U4581 (N_4581,In_2281,In_407);
nor U4582 (N_4582,In_1507,In_1085);
or U4583 (N_4583,In_27,In_513);
nand U4584 (N_4584,In_545,In_1251);
nand U4585 (N_4585,In_1123,In_1681);
nand U4586 (N_4586,In_2414,In_1009);
nand U4587 (N_4587,In_162,In_1545);
or U4588 (N_4588,In_189,In_386);
or U4589 (N_4589,In_1667,In_18);
and U4590 (N_4590,In_485,In_2195);
nand U4591 (N_4591,In_304,In_110);
nand U4592 (N_4592,In_1704,In_164);
nand U4593 (N_4593,In_1861,In_1551);
or U4594 (N_4594,In_289,In_2138);
nor U4595 (N_4595,In_1958,In_508);
nand U4596 (N_4596,In_2063,In_2294);
and U4597 (N_4597,In_2057,In_1387);
or U4598 (N_4598,In_1051,In_2300);
nor U4599 (N_4599,In_2091,In_2195);
or U4600 (N_4600,In_1994,In_2439);
or U4601 (N_4601,In_846,In_64);
and U4602 (N_4602,In_645,In_1073);
and U4603 (N_4603,In_2074,In_1933);
or U4604 (N_4604,In_828,In_1189);
or U4605 (N_4605,In_83,In_322);
and U4606 (N_4606,In_422,In_564);
or U4607 (N_4607,In_315,In_1443);
or U4608 (N_4608,In_2391,In_1382);
nand U4609 (N_4609,In_179,In_405);
or U4610 (N_4610,In_1742,In_185);
or U4611 (N_4611,In_1447,In_2319);
nand U4612 (N_4612,In_740,In_2400);
nor U4613 (N_4613,In_2253,In_1393);
nand U4614 (N_4614,In_926,In_1167);
and U4615 (N_4615,In_968,In_1305);
nor U4616 (N_4616,In_1467,In_1700);
and U4617 (N_4617,In_1757,In_535);
or U4618 (N_4618,In_1272,In_1024);
and U4619 (N_4619,In_529,In_2348);
nor U4620 (N_4620,In_2353,In_1540);
or U4621 (N_4621,In_119,In_1209);
or U4622 (N_4622,In_965,In_239);
nand U4623 (N_4623,In_2412,In_267);
or U4624 (N_4624,In_2036,In_512);
or U4625 (N_4625,In_1087,In_1400);
nor U4626 (N_4626,In_59,In_1034);
nand U4627 (N_4627,In_455,In_277);
and U4628 (N_4628,In_641,In_938);
and U4629 (N_4629,In_1611,In_2322);
nor U4630 (N_4630,In_2251,In_1042);
or U4631 (N_4631,In_1626,In_1402);
and U4632 (N_4632,In_572,In_328);
nor U4633 (N_4633,In_1579,In_800);
nor U4634 (N_4634,In_1518,In_486);
or U4635 (N_4635,In_1626,In_982);
nand U4636 (N_4636,In_2185,In_2128);
nor U4637 (N_4637,In_1731,In_1551);
or U4638 (N_4638,In_873,In_1072);
nor U4639 (N_4639,In_2194,In_1973);
and U4640 (N_4640,In_271,In_2478);
nor U4641 (N_4641,In_645,In_1428);
nor U4642 (N_4642,In_499,In_1817);
and U4643 (N_4643,In_1229,In_2261);
or U4644 (N_4644,In_348,In_1680);
nand U4645 (N_4645,In_71,In_417);
and U4646 (N_4646,In_1302,In_526);
nand U4647 (N_4647,In_631,In_736);
xor U4648 (N_4648,In_2356,In_1249);
and U4649 (N_4649,In_1025,In_2488);
or U4650 (N_4650,In_1235,In_970);
nand U4651 (N_4651,In_1803,In_2306);
nand U4652 (N_4652,In_83,In_823);
nor U4653 (N_4653,In_2282,In_925);
nand U4654 (N_4654,In_257,In_1682);
or U4655 (N_4655,In_372,In_2021);
and U4656 (N_4656,In_968,In_747);
and U4657 (N_4657,In_1720,In_882);
nand U4658 (N_4658,In_1579,In_1058);
and U4659 (N_4659,In_1593,In_276);
nand U4660 (N_4660,In_705,In_1512);
nand U4661 (N_4661,In_803,In_1612);
or U4662 (N_4662,In_387,In_61);
nand U4663 (N_4663,In_717,In_2474);
nor U4664 (N_4664,In_2352,In_171);
or U4665 (N_4665,In_2390,In_1375);
and U4666 (N_4666,In_330,In_1664);
and U4667 (N_4667,In_1115,In_2391);
xor U4668 (N_4668,In_2014,In_2091);
or U4669 (N_4669,In_556,In_65);
nor U4670 (N_4670,In_1337,In_977);
or U4671 (N_4671,In_28,In_2210);
or U4672 (N_4672,In_973,In_1849);
nand U4673 (N_4673,In_1686,In_593);
nor U4674 (N_4674,In_1118,In_1244);
or U4675 (N_4675,In_473,In_706);
nand U4676 (N_4676,In_1810,In_2329);
nand U4677 (N_4677,In_735,In_2436);
or U4678 (N_4678,In_346,In_89);
and U4679 (N_4679,In_1978,In_1667);
and U4680 (N_4680,In_1704,In_56);
nor U4681 (N_4681,In_1528,In_107);
nor U4682 (N_4682,In_1487,In_238);
and U4683 (N_4683,In_1686,In_2214);
nor U4684 (N_4684,In_2263,In_716);
nand U4685 (N_4685,In_51,In_54);
and U4686 (N_4686,In_42,In_174);
or U4687 (N_4687,In_698,In_611);
nor U4688 (N_4688,In_2271,In_1740);
nand U4689 (N_4689,In_1054,In_1136);
nand U4690 (N_4690,In_1801,In_1747);
and U4691 (N_4691,In_450,In_563);
nand U4692 (N_4692,In_1584,In_438);
nand U4693 (N_4693,In_2466,In_729);
nand U4694 (N_4694,In_1354,In_378);
nor U4695 (N_4695,In_469,In_1998);
nor U4696 (N_4696,In_2277,In_875);
or U4697 (N_4697,In_1463,In_2434);
nand U4698 (N_4698,In_2308,In_1199);
xor U4699 (N_4699,In_916,In_1885);
nand U4700 (N_4700,In_986,In_2058);
nor U4701 (N_4701,In_2264,In_138);
nor U4702 (N_4702,In_2164,In_219);
nand U4703 (N_4703,In_2120,In_1867);
xor U4704 (N_4704,In_1320,In_601);
or U4705 (N_4705,In_1143,In_1911);
nor U4706 (N_4706,In_1346,In_1538);
or U4707 (N_4707,In_1829,In_645);
nor U4708 (N_4708,In_1509,In_353);
and U4709 (N_4709,In_1977,In_2044);
or U4710 (N_4710,In_2477,In_2445);
and U4711 (N_4711,In_1036,In_2425);
and U4712 (N_4712,In_2089,In_2251);
nand U4713 (N_4713,In_1552,In_1554);
and U4714 (N_4714,In_2219,In_1913);
nand U4715 (N_4715,In_647,In_687);
and U4716 (N_4716,In_1019,In_2334);
nor U4717 (N_4717,In_2388,In_1131);
nor U4718 (N_4718,In_723,In_1986);
nor U4719 (N_4719,In_767,In_1300);
and U4720 (N_4720,In_1521,In_930);
nand U4721 (N_4721,In_717,In_419);
nor U4722 (N_4722,In_1625,In_1190);
and U4723 (N_4723,In_258,In_1480);
and U4724 (N_4724,In_2171,In_1787);
or U4725 (N_4725,In_1723,In_382);
or U4726 (N_4726,In_1950,In_733);
nor U4727 (N_4727,In_1782,In_227);
or U4728 (N_4728,In_187,In_1802);
nor U4729 (N_4729,In_2079,In_1974);
nor U4730 (N_4730,In_229,In_384);
or U4731 (N_4731,In_243,In_553);
and U4732 (N_4732,In_268,In_2364);
nor U4733 (N_4733,In_2062,In_1644);
nand U4734 (N_4734,In_86,In_1073);
or U4735 (N_4735,In_2284,In_60);
nor U4736 (N_4736,In_1042,In_1252);
nand U4737 (N_4737,In_1491,In_2104);
nand U4738 (N_4738,In_279,In_1726);
nor U4739 (N_4739,In_2371,In_920);
xnor U4740 (N_4740,In_2015,In_304);
nand U4741 (N_4741,In_1737,In_2319);
nor U4742 (N_4742,In_830,In_835);
nor U4743 (N_4743,In_1903,In_2051);
or U4744 (N_4744,In_1134,In_731);
and U4745 (N_4745,In_602,In_514);
nor U4746 (N_4746,In_2172,In_1175);
or U4747 (N_4747,In_1725,In_1200);
xnor U4748 (N_4748,In_1823,In_1552);
nand U4749 (N_4749,In_1738,In_1816);
and U4750 (N_4750,In_1638,In_2326);
or U4751 (N_4751,In_1305,In_1902);
and U4752 (N_4752,In_1430,In_2095);
nor U4753 (N_4753,In_317,In_133);
nand U4754 (N_4754,In_1217,In_2067);
nand U4755 (N_4755,In_280,In_1559);
nand U4756 (N_4756,In_328,In_722);
xor U4757 (N_4757,In_804,In_1102);
or U4758 (N_4758,In_510,In_531);
nor U4759 (N_4759,In_1288,In_1921);
or U4760 (N_4760,In_521,In_1937);
nand U4761 (N_4761,In_1551,In_608);
or U4762 (N_4762,In_2098,In_1464);
and U4763 (N_4763,In_1148,In_1401);
nand U4764 (N_4764,In_899,In_1754);
or U4765 (N_4765,In_1037,In_1931);
nand U4766 (N_4766,In_1183,In_1298);
or U4767 (N_4767,In_626,In_533);
nand U4768 (N_4768,In_2430,In_1702);
nor U4769 (N_4769,In_632,In_1124);
and U4770 (N_4770,In_2066,In_2495);
nand U4771 (N_4771,In_1109,In_1025);
or U4772 (N_4772,In_2136,In_560);
nor U4773 (N_4773,In_2267,In_677);
nor U4774 (N_4774,In_933,In_663);
or U4775 (N_4775,In_22,In_2068);
and U4776 (N_4776,In_970,In_927);
nand U4777 (N_4777,In_2098,In_1987);
nor U4778 (N_4778,In_766,In_1554);
and U4779 (N_4779,In_1924,In_1911);
nand U4780 (N_4780,In_2247,In_1367);
nor U4781 (N_4781,In_1769,In_1687);
nor U4782 (N_4782,In_897,In_1451);
or U4783 (N_4783,In_1265,In_1416);
or U4784 (N_4784,In_2023,In_912);
or U4785 (N_4785,In_59,In_1427);
or U4786 (N_4786,In_2213,In_526);
or U4787 (N_4787,In_2275,In_287);
xor U4788 (N_4788,In_1665,In_1687);
and U4789 (N_4789,In_2190,In_781);
or U4790 (N_4790,In_1987,In_155);
nor U4791 (N_4791,In_2432,In_1146);
and U4792 (N_4792,In_2366,In_317);
nand U4793 (N_4793,In_2032,In_2164);
and U4794 (N_4794,In_1946,In_646);
nand U4795 (N_4795,In_2273,In_2339);
nor U4796 (N_4796,In_13,In_1494);
xnor U4797 (N_4797,In_1828,In_1863);
nand U4798 (N_4798,In_2429,In_1411);
or U4799 (N_4799,In_2051,In_1776);
and U4800 (N_4800,In_365,In_178);
and U4801 (N_4801,In_1551,In_653);
nor U4802 (N_4802,In_2001,In_1641);
and U4803 (N_4803,In_1324,In_265);
or U4804 (N_4804,In_1029,In_2420);
nand U4805 (N_4805,In_1087,In_2283);
and U4806 (N_4806,In_202,In_49);
and U4807 (N_4807,In_1938,In_1626);
nor U4808 (N_4808,In_35,In_218);
nand U4809 (N_4809,In_2007,In_1136);
or U4810 (N_4810,In_1324,In_908);
or U4811 (N_4811,In_1761,In_1834);
nor U4812 (N_4812,In_1015,In_614);
nand U4813 (N_4813,In_1321,In_71);
nor U4814 (N_4814,In_2357,In_1105);
nor U4815 (N_4815,In_367,In_2304);
nor U4816 (N_4816,In_817,In_950);
nand U4817 (N_4817,In_1902,In_432);
nor U4818 (N_4818,In_681,In_1456);
nand U4819 (N_4819,In_1085,In_2019);
nand U4820 (N_4820,In_842,In_507);
nand U4821 (N_4821,In_29,In_393);
and U4822 (N_4822,In_1952,In_2272);
and U4823 (N_4823,In_254,In_2238);
nand U4824 (N_4824,In_368,In_742);
nor U4825 (N_4825,In_1381,In_1236);
or U4826 (N_4826,In_369,In_1735);
nor U4827 (N_4827,In_596,In_70);
nor U4828 (N_4828,In_472,In_1760);
xnor U4829 (N_4829,In_919,In_2075);
and U4830 (N_4830,In_1881,In_2362);
or U4831 (N_4831,In_994,In_202);
or U4832 (N_4832,In_420,In_1826);
and U4833 (N_4833,In_1634,In_604);
nand U4834 (N_4834,In_2286,In_1315);
nand U4835 (N_4835,In_1290,In_1990);
nor U4836 (N_4836,In_368,In_97);
and U4837 (N_4837,In_1520,In_1978);
nand U4838 (N_4838,In_2360,In_1191);
or U4839 (N_4839,In_1389,In_118);
nand U4840 (N_4840,In_298,In_1053);
or U4841 (N_4841,In_1411,In_227);
nor U4842 (N_4842,In_605,In_2289);
nor U4843 (N_4843,In_85,In_464);
nand U4844 (N_4844,In_884,In_558);
or U4845 (N_4845,In_1669,In_2210);
nor U4846 (N_4846,In_914,In_391);
and U4847 (N_4847,In_1738,In_245);
nand U4848 (N_4848,In_1412,In_847);
or U4849 (N_4849,In_1538,In_2057);
nand U4850 (N_4850,In_1065,In_227);
or U4851 (N_4851,In_2317,In_1516);
and U4852 (N_4852,In_2445,In_1491);
xnor U4853 (N_4853,In_1798,In_1505);
nand U4854 (N_4854,In_968,In_1472);
nor U4855 (N_4855,In_1222,In_917);
nand U4856 (N_4856,In_2395,In_1699);
nor U4857 (N_4857,In_2061,In_872);
or U4858 (N_4858,In_883,In_1221);
nor U4859 (N_4859,In_119,In_1550);
or U4860 (N_4860,In_262,In_766);
and U4861 (N_4861,In_887,In_259);
or U4862 (N_4862,In_1908,In_1409);
nor U4863 (N_4863,In_848,In_2257);
nand U4864 (N_4864,In_1976,In_1231);
or U4865 (N_4865,In_1565,In_811);
and U4866 (N_4866,In_2280,In_2155);
nor U4867 (N_4867,In_1355,In_112);
nand U4868 (N_4868,In_726,In_1987);
and U4869 (N_4869,In_1845,In_1752);
and U4870 (N_4870,In_2495,In_140);
nor U4871 (N_4871,In_1344,In_128);
nand U4872 (N_4872,In_999,In_363);
nor U4873 (N_4873,In_652,In_228);
nor U4874 (N_4874,In_2261,In_1748);
or U4875 (N_4875,In_102,In_1832);
nor U4876 (N_4876,In_910,In_1480);
and U4877 (N_4877,In_1122,In_458);
xnor U4878 (N_4878,In_775,In_2368);
nor U4879 (N_4879,In_526,In_888);
or U4880 (N_4880,In_2450,In_1409);
or U4881 (N_4881,In_1705,In_109);
and U4882 (N_4882,In_304,In_96);
or U4883 (N_4883,In_1839,In_1201);
nor U4884 (N_4884,In_141,In_1737);
xnor U4885 (N_4885,In_1875,In_90);
nand U4886 (N_4886,In_2097,In_2153);
nand U4887 (N_4887,In_950,In_344);
nor U4888 (N_4888,In_294,In_977);
and U4889 (N_4889,In_1942,In_2090);
and U4890 (N_4890,In_1021,In_87);
nand U4891 (N_4891,In_1970,In_993);
nand U4892 (N_4892,In_1304,In_2375);
xnor U4893 (N_4893,In_2368,In_2318);
nand U4894 (N_4894,In_457,In_0);
nand U4895 (N_4895,In_505,In_850);
nor U4896 (N_4896,In_792,In_1378);
nor U4897 (N_4897,In_1159,In_1872);
and U4898 (N_4898,In_297,In_912);
and U4899 (N_4899,In_1427,In_993);
and U4900 (N_4900,In_1526,In_1658);
nor U4901 (N_4901,In_681,In_2005);
or U4902 (N_4902,In_1211,In_2128);
or U4903 (N_4903,In_61,In_1331);
or U4904 (N_4904,In_2011,In_542);
nand U4905 (N_4905,In_1624,In_1252);
and U4906 (N_4906,In_573,In_752);
or U4907 (N_4907,In_1149,In_46);
or U4908 (N_4908,In_1799,In_1785);
nor U4909 (N_4909,In_693,In_381);
nor U4910 (N_4910,In_1719,In_0);
nand U4911 (N_4911,In_1982,In_937);
or U4912 (N_4912,In_1489,In_2404);
and U4913 (N_4913,In_707,In_993);
nor U4914 (N_4914,In_2278,In_354);
nand U4915 (N_4915,In_2364,In_777);
or U4916 (N_4916,In_2039,In_170);
nor U4917 (N_4917,In_1375,In_2136);
nor U4918 (N_4918,In_1108,In_1344);
nor U4919 (N_4919,In_1022,In_2289);
nand U4920 (N_4920,In_310,In_59);
or U4921 (N_4921,In_106,In_1149);
nand U4922 (N_4922,In_1016,In_1373);
and U4923 (N_4923,In_1302,In_1674);
nand U4924 (N_4924,In_82,In_1891);
nand U4925 (N_4925,In_1871,In_650);
or U4926 (N_4926,In_687,In_1007);
nand U4927 (N_4927,In_2160,In_1881);
or U4928 (N_4928,In_2234,In_2489);
or U4929 (N_4929,In_401,In_2108);
nand U4930 (N_4930,In_2282,In_760);
or U4931 (N_4931,In_1544,In_190);
and U4932 (N_4932,In_272,In_1462);
or U4933 (N_4933,In_1959,In_1328);
or U4934 (N_4934,In_403,In_2141);
nor U4935 (N_4935,In_528,In_696);
or U4936 (N_4936,In_1877,In_138);
nor U4937 (N_4937,In_524,In_1904);
or U4938 (N_4938,In_1342,In_1904);
or U4939 (N_4939,In_1659,In_2346);
or U4940 (N_4940,In_1554,In_1011);
or U4941 (N_4941,In_1074,In_1995);
nand U4942 (N_4942,In_99,In_332);
and U4943 (N_4943,In_835,In_2063);
nor U4944 (N_4944,In_2155,In_77);
and U4945 (N_4945,In_1333,In_230);
or U4946 (N_4946,In_589,In_176);
and U4947 (N_4947,In_1049,In_1575);
nand U4948 (N_4948,In_620,In_2243);
and U4949 (N_4949,In_2274,In_1319);
xnor U4950 (N_4950,In_623,In_632);
nor U4951 (N_4951,In_516,In_21);
or U4952 (N_4952,In_1545,In_2086);
or U4953 (N_4953,In_11,In_1755);
nor U4954 (N_4954,In_1640,In_860);
nor U4955 (N_4955,In_1550,In_413);
or U4956 (N_4956,In_282,In_1409);
and U4957 (N_4957,In_1625,In_2463);
or U4958 (N_4958,In_2472,In_1407);
nor U4959 (N_4959,In_1620,In_364);
or U4960 (N_4960,In_1977,In_1941);
and U4961 (N_4961,In_207,In_98);
nand U4962 (N_4962,In_2377,In_2328);
or U4963 (N_4963,In_831,In_1969);
or U4964 (N_4964,In_1202,In_2235);
and U4965 (N_4965,In_1191,In_543);
or U4966 (N_4966,In_59,In_2485);
or U4967 (N_4967,In_1163,In_2312);
nor U4968 (N_4968,In_1127,In_694);
and U4969 (N_4969,In_1587,In_1357);
and U4970 (N_4970,In_2000,In_498);
and U4971 (N_4971,In_1445,In_1237);
and U4972 (N_4972,In_1732,In_891);
and U4973 (N_4973,In_767,In_565);
and U4974 (N_4974,In_1236,In_1098);
or U4975 (N_4975,In_862,In_1435);
and U4976 (N_4976,In_2027,In_2468);
and U4977 (N_4977,In_583,In_1306);
and U4978 (N_4978,In_2298,In_1139);
nand U4979 (N_4979,In_485,In_1871);
nor U4980 (N_4980,In_862,In_1645);
nor U4981 (N_4981,In_1210,In_756);
xor U4982 (N_4982,In_320,In_2219);
nor U4983 (N_4983,In_2469,In_1430);
nor U4984 (N_4984,In_323,In_1563);
or U4985 (N_4985,In_410,In_309);
nor U4986 (N_4986,In_1268,In_1504);
or U4987 (N_4987,In_2392,In_1934);
and U4988 (N_4988,In_580,In_784);
and U4989 (N_4989,In_433,In_835);
and U4990 (N_4990,In_1274,In_1266);
nand U4991 (N_4991,In_345,In_991);
nor U4992 (N_4992,In_451,In_2262);
or U4993 (N_4993,In_781,In_2280);
and U4994 (N_4994,In_343,In_1494);
nand U4995 (N_4995,In_110,In_1833);
or U4996 (N_4996,In_1894,In_135);
nor U4997 (N_4997,In_2075,In_1506);
or U4998 (N_4998,In_1971,In_1138);
nor U4999 (N_4999,In_831,In_1848);
and U5000 (N_5000,N_4512,N_424);
and U5001 (N_5001,N_3848,N_1330);
nor U5002 (N_5002,N_1042,N_4435);
nor U5003 (N_5003,N_1473,N_3905);
or U5004 (N_5004,N_3816,N_105);
or U5005 (N_5005,N_1178,N_491);
nand U5006 (N_5006,N_1173,N_322);
and U5007 (N_5007,N_4163,N_1488);
nand U5008 (N_5008,N_4220,N_1003);
nand U5009 (N_5009,N_2340,N_4426);
nor U5010 (N_5010,N_2894,N_2382);
and U5011 (N_5011,N_337,N_4318);
and U5012 (N_5012,N_4323,N_120);
and U5013 (N_5013,N_1202,N_4092);
nand U5014 (N_5014,N_3720,N_2144);
or U5015 (N_5015,N_2559,N_2577);
nand U5016 (N_5016,N_2022,N_2499);
or U5017 (N_5017,N_4589,N_3604);
nor U5018 (N_5018,N_3608,N_2047);
or U5019 (N_5019,N_877,N_800);
nand U5020 (N_5020,N_485,N_1419);
or U5021 (N_5021,N_2567,N_1892);
and U5022 (N_5022,N_4196,N_4662);
nor U5023 (N_5023,N_2890,N_249);
and U5024 (N_5024,N_2589,N_2539);
nand U5025 (N_5025,N_2722,N_3684);
nand U5026 (N_5026,N_2359,N_2760);
and U5027 (N_5027,N_3442,N_3930);
or U5028 (N_5028,N_3889,N_341);
and U5029 (N_5029,N_3430,N_4492);
nand U5030 (N_5030,N_3668,N_572);
and U5031 (N_5031,N_3323,N_1606);
nand U5032 (N_5032,N_4856,N_14);
and U5033 (N_5033,N_3853,N_4029);
nand U5034 (N_5034,N_1009,N_659);
or U5035 (N_5035,N_2247,N_3161);
or U5036 (N_5036,N_4903,N_4730);
nor U5037 (N_5037,N_4179,N_3259);
and U5038 (N_5038,N_1691,N_535);
nand U5039 (N_5039,N_1213,N_3421);
nor U5040 (N_5040,N_2717,N_2154);
nor U5041 (N_5041,N_1794,N_1571);
nand U5042 (N_5042,N_546,N_679);
or U5043 (N_5043,N_4235,N_2073);
or U5044 (N_5044,N_3039,N_1217);
or U5045 (N_5045,N_3731,N_1672);
or U5046 (N_5046,N_4591,N_2546);
and U5047 (N_5047,N_1838,N_2579);
and U5048 (N_5048,N_945,N_3948);
nor U5049 (N_5049,N_4201,N_2442);
or U5050 (N_5050,N_2414,N_4205);
nand U5051 (N_5051,N_462,N_2179);
or U5052 (N_5052,N_2751,N_4843);
nand U5053 (N_5053,N_4046,N_1519);
nor U5054 (N_5054,N_3489,N_2912);
or U5055 (N_5055,N_584,N_3630);
and U5056 (N_5056,N_2036,N_2299);
nor U5057 (N_5057,N_2484,N_3943);
nand U5058 (N_5058,N_1122,N_616);
nand U5059 (N_5059,N_1129,N_1245);
or U5060 (N_5060,N_3739,N_2593);
or U5061 (N_5061,N_2835,N_812);
nand U5062 (N_5062,N_246,N_4604);
and U5063 (N_5063,N_3013,N_194);
and U5064 (N_5064,N_329,N_2253);
nor U5065 (N_5065,N_3225,N_2415);
nand U5066 (N_5066,N_2227,N_4468);
and U5067 (N_5067,N_1558,N_4486);
xor U5068 (N_5068,N_3652,N_1048);
and U5069 (N_5069,N_3584,N_4702);
and U5070 (N_5070,N_1992,N_1452);
nor U5071 (N_5071,N_3548,N_1443);
nand U5072 (N_5072,N_4705,N_512);
nand U5073 (N_5073,N_3766,N_2586);
nor U5074 (N_5074,N_931,N_3807);
or U5075 (N_5075,N_3502,N_1136);
nor U5076 (N_5076,N_4919,N_2055);
and U5077 (N_5077,N_513,N_1996);
and U5078 (N_5078,N_4286,N_4280);
or U5079 (N_5079,N_3945,N_2748);
and U5080 (N_5080,N_2413,N_2074);
nand U5081 (N_5081,N_2294,N_1233);
nor U5082 (N_5082,N_3193,N_2426);
nor U5083 (N_5083,N_3672,N_2849);
and U5084 (N_5084,N_278,N_715);
or U5085 (N_5085,N_4792,N_4351);
or U5086 (N_5086,N_2816,N_1349);
nor U5087 (N_5087,N_743,N_4099);
nor U5088 (N_5088,N_328,N_2996);
nor U5089 (N_5089,N_676,N_69);
nor U5090 (N_5090,N_3389,N_311);
nor U5091 (N_5091,N_1195,N_4209);
nor U5092 (N_5092,N_1235,N_4578);
or U5093 (N_5093,N_2258,N_3079);
nor U5094 (N_5094,N_2892,N_1466);
or U5095 (N_5095,N_4550,N_4976);
and U5096 (N_5096,N_1528,N_3198);
nor U5097 (N_5097,N_3524,N_4757);
or U5098 (N_5098,N_2380,N_3093);
or U5099 (N_5099,N_3879,N_2251);
and U5100 (N_5100,N_3476,N_2598);
nor U5101 (N_5101,N_1295,N_2812);
and U5102 (N_5102,N_4332,N_729);
nor U5103 (N_5103,N_1924,N_2477);
or U5104 (N_5104,N_2680,N_399);
or U5105 (N_5105,N_3743,N_4453);
or U5106 (N_5106,N_3362,N_3843);
and U5107 (N_5107,N_1510,N_205);
or U5108 (N_5108,N_4375,N_4579);
nand U5109 (N_5109,N_2041,N_936);
or U5110 (N_5110,N_2053,N_4929);
nand U5111 (N_5111,N_4513,N_795);
nor U5112 (N_5112,N_4908,N_684);
nor U5113 (N_5113,N_4729,N_4783);
or U5114 (N_5114,N_3653,N_220);
nand U5115 (N_5115,N_3959,N_4500);
nor U5116 (N_5116,N_3311,N_2627);
nand U5117 (N_5117,N_4614,N_4668);
nor U5118 (N_5118,N_137,N_822);
nor U5119 (N_5119,N_2152,N_1763);
or U5120 (N_5120,N_2583,N_3304);
nor U5121 (N_5121,N_3447,N_1154);
nand U5122 (N_5122,N_1436,N_1700);
nand U5123 (N_5123,N_298,N_4664);
and U5124 (N_5124,N_4941,N_2723);
nor U5125 (N_5125,N_409,N_4768);
nand U5126 (N_5126,N_1556,N_2199);
and U5127 (N_5127,N_4683,N_4852);
nand U5128 (N_5128,N_2172,N_1657);
nand U5129 (N_5129,N_1744,N_1053);
nor U5130 (N_5130,N_1179,N_3043);
and U5131 (N_5131,N_1739,N_3497);
or U5132 (N_5132,N_717,N_3970);
and U5133 (N_5133,N_810,N_1906);
or U5134 (N_5134,N_4054,N_1250);
nand U5135 (N_5135,N_862,N_4180);
nor U5136 (N_5136,N_4674,N_1397);
and U5137 (N_5137,N_3725,N_2824);
nand U5138 (N_5138,N_2037,N_130);
or U5139 (N_5139,N_2288,N_3967);
and U5140 (N_5140,N_1870,N_1145);
nor U5141 (N_5141,N_4562,N_1320);
nor U5142 (N_5142,N_1614,N_510);
nand U5143 (N_5143,N_3368,N_1516);
and U5144 (N_5144,N_3089,N_1782);
and U5145 (N_5145,N_2787,N_3133);
nor U5146 (N_5146,N_1599,N_3852);
and U5147 (N_5147,N_1814,N_3050);
and U5148 (N_5148,N_4236,N_2241);
or U5149 (N_5149,N_4491,N_3567);
and U5150 (N_5150,N_4018,N_1465);
or U5151 (N_5151,N_1006,N_1718);
nand U5152 (N_5152,N_3159,N_4134);
and U5153 (N_5153,N_4073,N_42);
and U5154 (N_5154,N_557,N_2162);
or U5155 (N_5155,N_4467,N_4593);
nor U5156 (N_5156,N_1773,N_3446);
nand U5157 (N_5157,N_2486,N_425);
nor U5158 (N_5158,N_1044,N_2690);
or U5159 (N_5159,N_2455,N_725);
nor U5160 (N_5160,N_3735,N_4516);
nor U5161 (N_5161,N_1970,N_3427);
and U5162 (N_5162,N_3269,N_3029);
or U5163 (N_5163,N_4725,N_2272);
nor U5164 (N_5164,N_3054,N_4088);
nor U5165 (N_5165,N_2384,N_3227);
nor U5166 (N_5166,N_318,N_3629);
nand U5167 (N_5167,N_1741,N_3402);
or U5168 (N_5168,N_4350,N_4336);
and U5169 (N_5169,N_77,N_1057);
nand U5170 (N_5170,N_1896,N_282);
or U5171 (N_5171,N_2326,N_2902);
nor U5172 (N_5172,N_297,N_2908);
nor U5173 (N_5173,N_3370,N_526);
and U5174 (N_5174,N_3593,N_3886);
or U5175 (N_5175,N_3541,N_4836);
or U5176 (N_5176,N_3200,N_2121);
or U5177 (N_5177,N_44,N_1902);
or U5178 (N_5178,N_3414,N_87);
nand U5179 (N_5179,N_2328,N_1098);
nand U5180 (N_5180,N_2271,N_4653);
nor U5181 (N_5181,N_1076,N_360);
and U5182 (N_5182,N_3728,N_2524);
nor U5183 (N_5183,N_3066,N_1461);
or U5184 (N_5184,N_602,N_3018);
nand U5185 (N_5185,N_3419,N_4630);
nor U5186 (N_5186,N_4006,N_3420);
nor U5187 (N_5187,N_4921,N_2592);
nand U5188 (N_5188,N_4264,N_26);
nand U5189 (N_5189,N_3927,N_3222);
nor U5190 (N_5190,N_4410,N_334);
or U5191 (N_5191,N_3415,N_1467);
or U5192 (N_5192,N_3175,N_682);
and U5193 (N_5193,N_2361,N_1449);
or U5194 (N_5194,N_2853,N_236);
nor U5195 (N_5195,N_864,N_705);
nand U5196 (N_5196,N_1878,N_2551);
nor U5197 (N_5197,N_3697,N_1781);
nor U5198 (N_5198,N_2840,N_1161);
or U5199 (N_5199,N_3104,N_3907);
and U5200 (N_5200,N_4892,N_2907);
and U5201 (N_5201,N_1551,N_4958);
nand U5202 (N_5202,N_4389,N_131);
nand U5203 (N_5203,N_228,N_3004);
nand U5204 (N_5204,N_998,N_3971);
nor U5205 (N_5205,N_3082,N_3596);
xnor U5206 (N_5206,N_3965,N_3106);
nor U5207 (N_5207,N_2406,N_1738);
nand U5208 (N_5208,N_4273,N_798);
nand U5209 (N_5209,N_1909,N_4329);
nor U5210 (N_5210,N_2000,N_4618);
nor U5211 (N_5211,N_4671,N_3276);
nor U5212 (N_5212,N_857,N_4140);
or U5213 (N_5213,N_3473,N_1051);
nor U5214 (N_5214,N_4412,N_3020);
nand U5215 (N_5215,N_2692,N_4128);
and U5216 (N_5216,N_1618,N_4631);
nor U5217 (N_5217,N_3547,N_588);
or U5218 (N_5218,N_4447,N_880);
or U5219 (N_5219,N_1791,N_1297);
and U5220 (N_5220,N_3403,N_1568);
nand U5221 (N_5221,N_1221,N_4807);
or U5222 (N_5222,N_2847,N_4905);
nand U5223 (N_5223,N_570,N_2485);
or U5224 (N_5224,N_3859,N_1327);
nor U5225 (N_5225,N_2004,N_2839);
nand U5226 (N_5226,N_2177,N_3456);
nand U5227 (N_5227,N_3391,N_3230);
nor U5228 (N_5228,N_3857,N_27);
nand U5229 (N_5229,N_2400,N_40);
and U5230 (N_5230,N_1273,N_314);
nand U5231 (N_5231,N_2291,N_111);
nor U5232 (N_5232,N_2799,N_1212);
and U5233 (N_5233,N_4736,N_2865);
xor U5234 (N_5234,N_1958,N_3101);
or U5235 (N_5235,N_961,N_1108);
nor U5236 (N_5236,N_3815,N_4393);
xor U5237 (N_5237,N_100,N_4756);
xor U5238 (N_5238,N_884,N_3395);
and U5239 (N_5239,N_515,N_1883);
nand U5240 (N_5240,N_4990,N_3088);
nor U5241 (N_5241,N_4814,N_1380);
or U5242 (N_5242,N_2806,N_7);
or U5243 (N_5243,N_464,N_2099);
or U5244 (N_5244,N_3319,N_3519);
nor U5245 (N_5245,N_4869,N_2206);
or U5246 (N_5246,N_4753,N_1943);
and U5247 (N_5247,N_2317,N_2914);
nor U5248 (N_5248,N_3031,N_3560);
nor U5249 (N_5249,N_504,N_4857);
nor U5250 (N_5250,N_3130,N_3439);
nand U5251 (N_5251,N_2571,N_35);
or U5252 (N_5252,N_3600,N_4870);
and U5253 (N_5253,N_1430,N_3284);
and U5254 (N_5254,N_3117,N_2255);
or U5255 (N_5255,N_4483,N_4890);
nor U5256 (N_5256,N_2945,N_3796);
nand U5257 (N_5257,N_2515,N_4111);
nor U5258 (N_5258,N_2473,N_4381);
nand U5259 (N_5259,N_3721,N_281);
or U5260 (N_5260,N_4603,N_3078);
nand U5261 (N_5261,N_4392,N_3030);
or U5262 (N_5262,N_3124,N_4456);
or U5263 (N_5263,N_2572,N_1387);
or U5264 (N_5264,N_4217,N_3734);
and U5265 (N_5265,N_143,N_3564);
nand U5266 (N_5266,N_4035,N_2023);
or U5267 (N_5267,N_4896,N_3286);
and U5268 (N_5268,N_166,N_3814);
nor U5269 (N_5269,N_4413,N_1932);
and U5270 (N_5270,N_3585,N_1645);
and U5271 (N_5271,N_1208,N_802);
and U5272 (N_5272,N_4090,N_4639);
and U5273 (N_5273,N_633,N_104);
and U5274 (N_5274,N_3057,N_4176);
or U5275 (N_5275,N_1822,N_1811);
or U5276 (N_5276,N_3771,N_762);
nand U5277 (N_5277,N_3196,N_3484);
nor U5278 (N_5278,N_1746,N_4800);
or U5279 (N_5279,N_573,N_1965);
or U5280 (N_5280,N_1020,N_1824);
or U5281 (N_5281,N_4292,N_900);
nor U5282 (N_5282,N_837,N_3428);
nand U5283 (N_5283,N_4017,N_600);
nor U5284 (N_5284,N_1347,N_4522);
or U5285 (N_5285,N_3682,N_3787);
nor U5286 (N_5286,N_2028,N_2830);
and U5287 (N_5287,N_1277,N_1707);
nor U5288 (N_5288,N_4053,N_2375);
nand U5289 (N_5289,N_3330,N_828);
and U5290 (N_5290,N_1735,N_1591);
nor U5291 (N_5291,N_628,N_1316);
and U5292 (N_5292,N_4401,N_1957);
nand U5293 (N_5293,N_2611,N_2352);
nand U5294 (N_5294,N_1263,N_1663);
and U5295 (N_5295,N_1246,N_2149);
nand U5296 (N_5296,N_4815,N_1265);
and U5297 (N_5297,N_3165,N_4396);
nor U5298 (N_5298,N_3347,N_1062);
or U5299 (N_5299,N_3180,N_859);
nand U5300 (N_5300,N_2535,N_3912);
nand U5301 (N_5301,N_3932,N_3637);
and U5302 (N_5302,N_4148,N_3396);
nor U5303 (N_5303,N_579,N_4731);
and U5304 (N_5304,N_2059,N_2276);
nand U5305 (N_5305,N_2412,N_3443);
nor U5306 (N_5306,N_2664,N_1063);
nor U5307 (N_5307,N_1294,N_1);
and U5308 (N_5308,N_1312,N_833);
xor U5309 (N_5309,N_2240,N_4543);
nand U5310 (N_5310,N_3619,N_3174);
xor U5311 (N_5311,N_319,N_3021);
or U5312 (N_5312,N_129,N_735);
nor U5313 (N_5313,N_4279,N_2314);
nand U5314 (N_5314,N_2993,N_4993);
or U5315 (N_5315,N_4372,N_2309);
nor U5316 (N_5316,N_4417,N_3738);
xor U5317 (N_5317,N_3713,N_1588);
or U5318 (N_5318,N_3376,N_490);
or U5319 (N_5319,N_1755,N_4581);
or U5320 (N_5320,N_3000,N_562);
and U5321 (N_5321,N_1120,N_516);
nor U5322 (N_5322,N_2850,N_2280);
xor U5323 (N_5323,N_3090,N_1733);
xor U5324 (N_5324,N_903,N_4839);
and U5325 (N_5325,N_2715,N_1816);
nand U5326 (N_5326,N_1169,N_3621);
nand U5327 (N_5327,N_1324,N_4519);
or U5328 (N_5328,N_4656,N_4887);
or U5329 (N_5329,N_2953,N_734);
xnor U5330 (N_5330,N_3392,N_3291);
and U5331 (N_5331,N_4331,N_3867);
xor U5332 (N_5332,N_4459,N_3163);
and U5333 (N_5333,N_2783,N_1520);
nand U5334 (N_5334,N_225,N_2187);
xnor U5335 (N_5335,N_4501,N_867);
nor U5336 (N_5336,N_3969,N_3081);
nor U5337 (N_5337,N_552,N_2275);
xnor U5338 (N_5338,N_4170,N_3955);
or U5339 (N_5339,N_2540,N_1605);
and U5340 (N_5340,N_1266,N_408);
nand U5341 (N_5341,N_3658,N_4087);
and U5342 (N_5342,N_366,N_1040);
and U5343 (N_5343,N_3818,N_403);
or U5344 (N_5344,N_3753,N_3983);
and U5345 (N_5345,N_3659,N_2481);
nor U5346 (N_5346,N_4949,N_3544);
or U5347 (N_5347,N_3663,N_25);
nand U5348 (N_5348,N_1680,N_4652);
and U5349 (N_5349,N_1889,N_1160);
nand U5350 (N_5350,N_4781,N_180);
nor U5351 (N_5351,N_3906,N_1182);
or U5352 (N_5352,N_2233,N_1550);
nor U5353 (N_5353,N_4832,N_910);
or U5354 (N_5354,N_2995,N_608);
or U5355 (N_5355,N_4033,N_2286);
nand U5356 (N_5356,N_925,N_1092);
nand U5357 (N_5357,N_1868,N_1495);
nor U5358 (N_5358,N_289,N_4617);
nand U5359 (N_5359,N_4089,N_2886);
nor U5360 (N_5360,N_3002,N_309);
nand U5361 (N_5361,N_3792,N_215);
nand U5362 (N_5362,N_907,N_4060);
or U5363 (N_5363,N_2160,N_4144);
or U5364 (N_5364,N_2236,N_1190);
nor U5365 (N_5365,N_4732,N_4126);
nand U5366 (N_5366,N_1128,N_3741);
nand U5367 (N_5367,N_766,N_3958);
nor U5368 (N_5368,N_4830,N_2332);
or U5369 (N_5369,N_4735,N_3279);
and U5370 (N_5370,N_4967,N_4241);
or U5371 (N_5371,N_2209,N_2726);
nor U5372 (N_5372,N_2256,N_2098);
and U5373 (N_5373,N_3216,N_4225);
and U5374 (N_5374,N_1354,N_3322);
nor U5375 (N_5375,N_1357,N_2402);
or U5376 (N_5376,N_4635,N_1064);
or U5377 (N_5377,N_1474,N_3510);
and U5378 (N_5378,N_2290,N_469);
or U5379 (N_5379,N_3310,N_890);
nand U5380 (N_5380,N_1699,N_1784);
nand U5381 (N_5381,N_4608,N_641);
and U5382 (N_5382,N_497,N_4003);
and U5383 (N_5383,N_4463,N_187);
and U5384 (N_5384,N_839,N_1775);
and U5385 (N_5385,N_3236,N_2916);
nand U5386 (N_5386,N_3271,N_4950);
nand U5387 (N_5387,N_4971,N_242);
nor U5388 (N_5388,N_1632,N_3450);
nor U5389 (N_5389,N_495,N_4845);
nand U5390 (N_5390,N_231,N_1127);
or U5391 (N_5391,N_1884,N_1748);
nor U5392 (N_5392,N_2647,N_260);
nand U5393 (N_5393,N_4928,N_1567);
nor U5394 (N_5394,N_1462,N_3744);
nor U5395 (N_5395,N_1963,N_2058);
and U5396 (N_5396,N_125,N_3944);
xnor U5397 (N_5397,N_4495,N_819);
or U5398 (N_5398,N_1971,N_4253);
or U5399 (N_5399,N_207,N_3636);
or U5400 (N_5400,N_2463,N_3551);
or U5401 (N_5401,N_2946,N_118);
nor U5402 (N_5402,N_1439,N_866);
nor U5403 (N_5403,N_4489,N_3342);
or U5404 (N_5404,N_1271,N_4992);
and U5405 (N_5405,N_4996,N_3762);
and U5406 (N_5406,N_3015,N_1066);
nand U5407 (N_5407,N_1721,N_620);
and U5408 (N_5408,N_539,N_1840);
and U5409 (N_5409,N_3898,N_2522);
nand U5410 (N_5410,N_2861,N_1578);
and U5411 (N_5411,N_4722,N_1543);
and U5412 (N_5412,N_1774,N_1472);
nand U5413 (N_5413,N_1493,N_2196);
and U5414 (N_5414,N_1174,N_1153);
nor U5415 (N_5415,N_4551,N_4699);
or U5416 (N_5416,N_1086,N_786);
or U5417 (N_5417,N_591,N_606);
or U5418 (N_5418,N_2489,N_3351);
and U5419 (N_5419,N_1603,N_2278);
nor U5420 (N_5420,N_256,N_4998);
and U5421 (N_5421,N_3026,N_3278);
nand U5422 (N_5422,N_2124,N_2093);
and U5423 (N_5423,N_2292,N_234);
nor U5424 (N_5424,N_4481,N_2221);
and U5425 (N_5425,N_1951,N_1766);
and U5426 (N_5426,N_3777,N_2081);
nor U5427 (N_5427,N_1124,N_247);
or U5428 (N_5428,N_4438,N_949);
and U5429 (N_5429,N_4493,N_938);
xor U5430 (N_5430,N_2507,N_3752);
and U5431 (N_5431,N_2257,N_4977);
nor U5432 (N_5432,N_2681,N_2604);
and U5433 (N_5433,N_2837,N_2032);
nor U5434 (N_5434,N_3966,N_2424);
or U5435 (N_5435,N_2940,N_2900);
or U5436 (N_5436,N_952,N_897);
nand U5437 (N_5437,N_1832,N_3509);
nor U5438 (N_5438,N_665,N_4432);
and U5439 (N_5439,N_4861,N_2349);
or U5440 (N_5440,N_1821,N_3946);
and U5441 (N_5441,N_4521,N_1552);
nor U5442 (N_5442,N_1623,N_4156);
or U5443 (N_5443,N_3773,N_51);
nand U5444 (N_5444,N_2646,N_4268);
xor U5445 (N_5445,N_2158,N_4580);
nor U5446 (N_5446,N_2456,N_2786);
and U5447 (N_5447,N_894,N_4900);
and U5448 (N_5448,N_4051,N_1751);
or U5449 (N_5449,N_3793,N_2295);
and U5450 (N_5450,N_668,N_2762);
or U5451 (N_5451,N_2223,N_933);
nor U5452 (N_5452,N_3084,N_2667);
nor U5453 (N_5453,N_92,N_2355);
nor U5454 (N_5454,N_1640,N_1726);
or U5455 (N_5455,N_2465,N_1956);
nand U5456 (N_5456,N_2635,N_2417);
nor U5457 (N_5457,N_950,N_3156);
nand U5458 (N_5458,N_4421,N_2501);
nand U5459 (N_5459,N_4437,N_2947);
nand U5460 (N_5460,N_4161,N_2198);
nor U5461 (N_5461,N_78,N_1926);
xnor U5462 (N_5462,N_3614,N_3883);
or U5463 (N_5463,N_1139,N_479);
nand U5464 (N_5464,N_1315,N_3654);
and U5465 (N_5465,N_2142,N_3924);
or U5466 (N_5466,N_2620,N_2374);
nand U5467 (N_5467,N_958,N_957);
or U5468 (N_5468,N_4177,N_4898);
nor U5469 (N_5469,N_1405,N_1104);
xnor U5470 (N_5470,N_492,N_2769);
and U5471 (N_5471,N_2109,N_791);
or U5472 (N_5472,N_2495,N_121);
nor U5473 (N_5473,N_3973,N_1252);
nand U5474 (N_5474,N_1101,N_4549);
and U5475 (N_5475,N_3281,N_636);
or U5476 (N_5476,N_3918,N_972);
nor U5477 (N_5477,N_1573,N_4019);
nor U5478 (N_5478,N_2684,N_2920);
nor U5479 (N_5479,N_1017,N_2882);
and U5480 (N_5480,N_999,N_4766);
or U5481 (N_5481,N_2588,N_3894);
and U5482 (N_5482,N_3916,N_3590);
nand U5483 (N_5483,N_1593,N_1929);
nand U5484 (N_5484,N_4964,N_3253);
nor U5485 (N_5485,N_1036,N_3767);
or U5486 (N_5486,N_2756,N_4723);
and U5487 (N_5487,N_4021,N_3052);
nand U5488 (N_5488,N_407,N_3267);
or U5489 (N_5489,N_2738,N_3102);
nand U5490 (N_5490,N_640,N_1914);
nor U5491 (N_5491,N_2768,N_85);
nor U5492 (N_5492,N_3293,N_4607);
xor U5493 (N_5493,N_109,N_2141);
and U5494 (N_5494,N_4160,N_4256);
nand U5495 (N_5495,N_1547,N_2712);
nand U5496 (N_5496,N_3774,N_780);
or U5497 (N_5497,N_744,N_4628);
and U5498 (N_5498,N_1323,N_2358);
and U5499 (N_5499,N_4423,N_2025);
or U5500 (N_5500,N_685,N_3570);
xor U5501 (N_5501,N_993,N_2147);
nor U5502 (N_5502,N_4465,N_4994);
nor U5503 (N_5503,N_421,N_1938);
and U5504 (N_5504,N_4763,N_4012);
or U5505 (N_5505,N_4918,N_1444);
nand U5506 (N_5506,N_499,N_932);
or U5507 (N_5507,N_2161,N_1404);
nand U5508 (N_5508,N_1607,N_881);
nor U5509 (N_5509,N_1968,N_1300);
and U5510 (N_5510,N_2784,N_2956);
and U5511 (N_5511,N_3367,N_4365);
and U5512 (N_5512,N_3494,N_706);
nor U5513 (N_5513,N_2804,N_2077);
and U5514 (N_5514,N_1478,N_1696);
nand U5515 (N_5515,N_139,N_1328);
nand U5516 (N_5516,N_1177,N_4065);
nor U5517 (N_5517,N_178,N_4008);
or U5518 (N_5518,N_2466,N_829);
or U5519 (N_5519,N_2429,N_2871);
nand U5520 (N_5520,N_2052,N_4822);
or U5521 (N_5521,N_4081,N_4740);
or U5522 (N_5522,N_4130,N_1501);
or U5523 (N_5523,N_3345,N_1877);
xor U5524 (N_5524,N_4678,N_4221);
or U5525 (N_5525,N_4215,N_2721);
and U5526 (N_5526,N_605,N_2277);
nor U5527 (N_5527,N_992,N_3241);
nor U5528 (N_5528,N_93,N_1238);
and U5529 (N_5529,N_173,N_520);
nand U5530 (N_5530,N_790,N_4302);
nor U5531 (N_5531,N_614,N_2);
nand U5532 (N_5532,N_1232,N_3411);
nand U5533 (N_5533,N_1765,N_2301);
nand U5534 (N_5534,N_1481,N_2672);
nand U5535 (N_5535,N_4842,N_4295);
nor U5536 (N_5536,N_2963,N_3938);
and U5537 (N_5537,N_4970,N_4469);
or U5538 (N_5538,N_2046,N_4983);
or U5539 (N_5539,N_1967,N_872);
nand U5540 (N_5540,N_3219,N_4430);
nand U5541 (N_5541,N_356,N_3841);
and U5542 (N_5542,N_630,N_661);
and U5543 (N_5543,N_357,N_3703);
nor U5544 (N_5544,N_1708,N_1882);
nand U5545 (N_5545,N_868,N_1904);
nand U5546 (N_5546,N_3194,N_2613);
nor U5547 (N_5547,N_4541,N_2243);
or U5548 (N_5548,N_2859,N_41);
nor U5549 (N_5549,N_658,N_1720);
nor U5550 (N_5550,N_181,N_4545);
nor U5551 (N_5551,N_2304,N_4709);
or U5552 (N_5552,N_2960,N_711);
or U5553 (N_5553,N_722,N_2386);
and U5554 (N_5554,N_851,N_2648);
nand U5555 (N_5555,N_4716,N_4363);
nor U5556 (N_5556,N_2521,N_4770);
nor U5557 (N_5557,N_1714,N_2747);
and U5558 (N_5558,N_4893,N_254);
and U5559 (N_5559,N_2383,N_1188);
nor U5560 (N_5560,N_4625,N_899);
or U5561 (N_5561,N_3623,N_1636);
and U5562 (N_5562,N_4181,N_638);
nand U5563 (N_5563,N_2350,N_370);
or U5564 (N_5564,N_4448,N_1579);
nand U5565 (N_5565,N_758,N_1539);
xnor U5566 (N_5566,N_3890,N_2982);
or U5567 (N_5567,N_1898,N_1670);
and U5568 (N_5568,N_4296,N_3515);
nand U5569 (N_5569,N_4335,N_1695);
or U5570 (N_5570,N_3303,N_2811);
or U5571 (N_5571,N_2118,N_2653);
or U5572 (N_5572,N_3417,N_2881);
nand U5573 (N_5573,N_2194,N_3695);
and U5574 (N_5574,N_190,N_2308);
nor U5575 (N_5575,N_2702,N_3837);
nand U5576 (N_5576,N_2215,N_553);
and U5577 (N_5577,N_2928,N_2852);
nand U5578 (N_5578,N_1535,N_1367);
or U5579 (N_5579,N_1422,N_3047);
or U5580 (N_5580,N_3302,N_3055);
or U5581 (N_5581,N_2265,N_1319);
nor U5582 (N_5582,N_3201,N_3715);
or U5583 (N_5583,N_4172,N_2006);
and U5584 (N_5584,N_1850,N_2935);
or U5585 (N_5585,N_1157,N_2765);
xor U5586 (N_5586,N_4162,N_1630);
nor U5587 (N_5587,N_1321,N_524);
nand U5588 (N_5588,N_3210,N_1325);
or U5589 (N_5589,N_4366,N_753);
and U5590 (N_5590,N_124,N_3794);
nand U5591 (N_5591,N_3709,N_2710);
and U5592 (N_5592,N_576,N_4613);
and U5593 (N_5593,N_687,N_892);
nand U5594 (N_5594,N_1867,N_2800);
nand U5595 (N_5595,N_3011,N_5);
nand U5596 (N_5596,N_4173,N_432);
nand U5597 (N_5597,N_2021,N_4953);
nand U5598 (N_5598,N_1805,N_1205);
or U5599 (N_5599,N_826,N_1989);
or U5600 (N_5600,N_3850,N_433);
nand U5601 (N_5601,N_1619,N_340);
nor U5602 (N_5602,N_4957,N_4847);
or U5603 (N_5603,N_4787,N_2655);
nor U5604 (N_5604,N_1050,N_3506);
and U5605 (N_5605,N_4920,N_2807);
or U5606 (N_5606,N_2767,N_3513);
or U5607 (N_5607,N_1856,N_1442);
and U5608 (N_5608,N_90,N_612);
nand U5609 (N_5609,N_2954,N_66);
nor U5610 (N_5610,N_2016,N_4133);
nor U5611 (N_5611,N_771,N_426);
and U5612 (N_5612,N_472,N_473);
or U5613 (N_5613,N_2776,N_293);
nand U5614 (N_5614,N_122,N_542);
nand U5615 (N_5615,N_3580,N_468);
nand U5616 (N_5616,N_1954,N_3788);
nand U5617 (N_5617,N_2819,N_1710);
and U5618 (N_5618,N_474,N_1975);
and U5619 (N_5619,N_1852,N_663);
nand U5620 (N_5620,N_846,N_1383);
nor U5621 (N_5621,N_3228,N_4101);
or U5622 (N_5622,N_594,N_2305);
nand U5623 (N_5623,N_3313,N_3220);
nor U5624 (N_5624,N_3840,N_4686);
xnor U5625 (N_5625,N_3940,N_3022);
and U5626 (N_5626,N_3469,N_718);
and U5627 (N_5627,N_782,N_792);
nand U5628 (N_5628,N_923,N_98);
or U5629 (N_5629,N_1446,N_847);
or U5630 (N_5630,N_4487,N_1549);
or U5631 (N_5631,N_1742,N_3736);
nand U5632 (N_5632,N_565,N_2387);
and U5633 (N_5633,N_3445,N_1067);
nand U5634 (N_5634,N_4771,N_1167);
nand U5635 (N_5635,N_2838,N_2422);
nor U5636 (N_5636,N_18,N_2341);
xnor U5637 (N_5637,N_4285,N_2678);
and U5638 (N_5638,N_52,N_4700);
and U5639 (N_5639,N_3400,N_4833);
nand U5640 (N_5640,N_2615,N_1118);
nor U5641 (N_5641,N_20,N_343);
nand U5642 (N_5642,N_4710,N_1757);
and U5643 (N_5643,N_2553,N_2616);
nand U5644 (N_5644,N_2064,N_4989);
or U5645 (N_5645,N_4411,N_1379);
and U5646 (N_5646,N_136,N_162);
or U5647 (N_5647,N_3891,N_2883);
nand U5648 (N_5648,N_2229,N_1538);
or U5649 (N_5649,N_865,N_4877);
nor U5650 (N_5650,N_922,N_1283);
nor U5651 (N_5651,N_4093,N_455);
nor U5652 (N_5652,N_2825,N_3339);
or U5653 (N_5653,N_4605,N_1102);
nor U5654 (N_5654,N_2011,N_132);
nor U5655 (N_5655,N_2754,N_1745);
nor U5656 (N_5656,N_519,N_4059);
nor U5657 (N_5657,N_1366,N_1105);
or U5658 (N_5658,N_2034,N_820);
nor U5659 (N_5659,N_4755,N_2574);
nand U5660 (N_5660,N_172,N_2729);
nand U5661 (N_5661,N_3675,N_2879);
and U5662 (N_5662,N_89,N_4416);
nor U5663 (N_5663,N_724,N_3963);
or U5664 (N_5664,N_2201,N_674);
nand U5665 (N_5665,N_237,N_1229);
or U5666 (N_5666,N_2033,N_694);
nor U5667 (N_5667,N_4926,N_1533);
and U5668 (N_5668,N_3316,N_554);
nor U5669 (N_5669,N_1458,N_4517);
nor U5670 (N_5670,N_2862,N_3385);
nand U5671 (N_5671,N_1192,N_2437);
and U5672 (N_5672,N_1955,N_3032);
nand U5673 (N_5673,N_4010,N_3212);
nand U5674 (N_5674,N_1402,N_106);
and U5675 (N_5675,N_2955,N_2066);
and U5676 (N_5676,N_1624,N_1371);
or U5677 (N_5677,N_784,N_4049);
nor U5678 (N_5678,N_3622,N_4537);
and U5679 (N_5679,N_742,N_1692);
and U5680 (N_5680,N_1825,N_2260);
nand U5681 (N_5681,N_2120,N_4113);
and U5682 (N_5682,N_443,N_2425);
nor U5683 (N_5683,N_418,N_454);
or U5684 (N_5684,N_953,N_2836);
nand U5685 (N_5685,N_4105,N_3457);
nand U5686 (N_5686,N_2758,N_1555);
or U5687 (N_5687,N_3681,N_4004);
or U5688 (N_5688,N_3746,N_4252);
or U5689 (N_5689,N_2042,N_1203);
or U5690 (N_5690,N_4200,N_3994);
nor U5691 (N_5691,N_359,N_3355);
or U5692 (N_5692,N_1536,N_2102);
nand U5693 (N_5693,N_2632,N_1611);
nor U5694 (N_5694,N_979,N_4310);
and U5695 (N_5695,N_4028,N_1424);
nor U5696 (N_5696,N_751,N_434);
nand U5697 (N_5697,N_3926,N_3125);
nor U5698 (N_5698,N_1407,N_3247);
and U5699 (N_5699,N_250,N_16);
and U5700 (N_5700,N_1835,N_4223);
nand U5701 (N_5701,N_2703,N_2622);
and U5702 (N_5702,N_2357,N_4397);
nor U5703 (N_5703,N_3876,N_2938);
nor U5704 (N_5704,N_2428,N_4024);
and U5705 (N_5705,N_2395,N_2660);
or U5706 (N_5706,N_3528,N_1121);
or U5707 (N_5707,N_726,N_2339);
nand U5708 (N_5708,N_3218,N_416);
or U5709 (N_5709,N_558,N_4899);
nor U5710 (N_5710,N_4239,N_1166);
nand U5711 (N_5711,N_1865,N_241);
nor U5712 (N_5712,N_2346,N_3188);
or U5713 (N_5713,N_2639,N_561);
nand U5714 (N_5714,N_2640,N_1544);
or U5715 (N_5715,N_196,N_4428);
nand U5716 (N_5716,N_3340,N_4554);
or U5717 (N_5717,N_222,N_330);
nand U5718 (N_5718,N_3718,N_4924);
and U5719 (N_5719,N_2633,N_4224);
or U5720 (N_5720,N_970,N_3140);
nor U5721 (N_5721,N_969,N_2370);
nor U5722 (N_5722,N_1639,N_4388);
xor U5723 (N_5723,N_1469,N_2163);
nand U5724 (N_5724,N_578,N_974);
nand U5725 (N_5725,N_634,N_738);
and U5726 (N_5726,N_2921,N_53);
and U5727 (N_5727,N_1486,N_3780);
or U5728 (N_5728,N_4063,N_3554);
nor U5729 (N_5729,N_2170,N_245);
or U5730 (N_5730,N_4263,N_2514);
and U5731 (N_5731,N_2534,N_1249);
nor U5732 (N_5732,N_2263,N_789);
or U5733 (N_5733,N_1230,N_4610);
and U5734 (N_5734,N_362,N_3805);
nor U5735 (N_5735,N_4758,N_452);
xor U5736 (N_5736,N_905,N_3847);
nor U5737 (N_5737,N_4538,N_768);
or U5738 (N_5738,N_4007,N_4072);
or U5739 (N_5739,N_3642,N_3027);
nand U5740 (N_5740,N_1336,N_2421);
nand U5741 (N_5741,N_4611,N_3665);
nand U5742 (N_5742,N_3633,N_4786);
nand U5743 (N_5743,N_3542,N_3761);
or U5744 (N_5744,N_1925,N_2480);
nand U5745 (N_5745,N_4788,N_3205);
nand U5746 (N_5746,N_980,N_331);
nand U5747 (N_5747,N_3587,N_818);
nand U5748 (N_5748,N_1747,N_276);
nor U5749 (N_5749,N_4742,N_4378);
nand U5750 (N_5750,N_3352,N_4307);
nand U5751 (N_5751,N_1269,N_2845);
nand U5752 (N_5752,N_700,N_4115);
and U5753 (N_5753,N_1848,N_3798);
or U5754 (N_5754,N_3327,N_1688);
and U5755 (N_5755,N_695,N_3985);
or U5756 (N_5756,N_971,N_4540);
nand U5757 (N_5757,N_3044,N_401);
and U5758 (N_5758,N_1658,N_4270);
or U5759 (N_5759,N_4210,N_350);
nor U5760 (N_5760,N_937,N_2219);
nand U5761 (N_5761,N_2606,N_2563);
xnor U5762 (N_5762,N_1753,N_4681);
nor U5763 (N_5763,N_1986,N_1846);
or U5764 (N_5764,N_707,N_4956);
and U5765 (N_5765,N_204,N_750);
nand U5766 (N_5766,N_202,N_2719);
nand U5767 (N_5767,N_4885,N_1392);
and U5768 (N_5768,N_2885,N_2975);
nand U5769 (N_5769,N_288,N_4257);
and U5770 (N_5770,N_80,N_1964);
or U5771 (N_5771,N_3987,N_2267);
nor U5772 (N_5772,N_1431,N_2701);
and U5773 (N_5773,N_3656,N_185);
nor U5774 (N_5774,N_2385,N_3569);
or U5775 (N_5775,N_2512,N_545);
nand U5776 (N_5776,N_3387,N_2060);
and U5777 (N_5777,N_301,N_1204);
or U5778 (N_5778,N_2556,N_3865);
nand U5779 (N_5779,N_1284,N_3080);
nor U5780 (N_5780,N_1715,N_2228);
nand U5781 (N_5781,N_1562,N_1196);
nand U5782 (N_5782,N_3657,N_794);
and U5783 (N_5783,N_3820,N_1089);
or U5784 (N_5784,N_808,N_567);
nand U5785 (N_5785,N_1871,N_807);
nor U5786 (N_5786,N_32,N_2268);
or U5787 (N_5787,N_4691,N_4434);
nand U5788 (N_5788,N_4648,N_2504);
nand U5789 (N_5789,N_1901,N_732);
nor U5790 (N_5790,N_475,N_2057);
nand U5791 (N_5791,N_2873,N_4277);
nand U5792 (N_5792,N_1425,N_4754);
nand U5793 (N_5793,N_2508,N_3854);
nor U5794 (N_5794,N_450,N_1170);
and U5795 (N_5795,N_4520,N_3132);
nand U5796 (N_5796,N_1455,N_142);
and U5797 (N_5797,N_3825,N_984);
nor U5798 (N_5798,N_4107,N_4476);
and U5799 (N_5799,N_1000,N_2530);
or U5800 (N_5800,N_3537,N_691);
nand U5801 (N_5801,N_65,N_4823);
nor U5802 (N_5802,N_4600,N_383);
nand U5803 (N_5803,N_384,N_2310);
nor U5804 (N_5804,N_817,N_157);
nand U5805 (N_5805,N_4594,N_3120);
nor U5806 (N_5806,N_453,N_2368);
nand U5807 (N_5807,N_4247,N_3775);
nor U5808 (N_5808,N_2642,N_97);
and U5809 (N_5809,N_2087,N_3878);
or U5810 (N_5810,N_4461,N_3511);
nor U5811 (N_5811,N_1450,N_4646);
nand U5812 (N_5812,N_4341,N_3296);
and U5813 (N_5813,N_1142,N_3588);
nand U5814 (N_5814,N_2870,N_4974);
and U5815 (N_5815,N_4563,N_60);
and U5816 (N_5816,N_3264,N_3372);
or U5817 (N_5817,N_3908,N_4657);
nand U5818 (N_5818,N_2029,N_2246);
nand U5819 (N_5819,N_2097,N_2178);
nor U5820 (N_5820,N_2910,N_3540);
and U5821 (N_5821,N_3424,N_3467);
nor U5822 (N_5822,N_4510,N_3260);
and U5823 (N_5823,N_1114,N_373);
or U5824 (N_5824,N_2331,N_1787);
or U5825 (N_5825,N_4282,N_171);
nor U5826 (N_5826,N_637,N_3957);
and U5827 (N_5827,N_3802,N_3202);
nor U5828 (N_5828,N_806,N_49);
nor U5829 (N_5829,N_623,N_3048);
nor U5830 (N_5830,N_2780,N_1502);
or U5831 (N_5831,N_3724,N_4150);
or U5832 (N_5832,N_3085,N_1764);
or U5833 (N_5833,N_2133,N_302);
or U5834 (N_5834,N_3676,N_873);
nor U5835 (N_5835,N_3669,N_1296);
and U5836 (N_5836,N_2843,N_4016);
or U5837 (N_5837,N_1813,N_61);
and U5838 (N_5838,N_197,N_3160);
or U5839 (N_5839,N_677,N_1697);
and U5840 (N_5840,N_2537,N_531);
or U5841 (N_5841,N_4025,N_4219);
or U5842 (N_5842,N_1990,N_1866);
and U5843 (N_5843,N_4091,N_2365);
nand U5844 (N_5844,N_3191,N_844);
nor U5845 (N_5845,N_4891,N_2582);
nand U5846 (N_5846,N_2078,N_1393);
and U5847 (N_5847,N_1123,N_4255);
nand U5848 (N_5848,N_3169,N_4966);
nand U5849 (N_5849,N_902,N_3143);
or U5850 (N_5850,N_3012,N_4158);
or U5851 (N_5851,N_577,N_2555);
and U5852 (N_5852,N_2104,N_1621);
or U5853 (N_5853,N_1094,N_259);
or U5854 (N_5854,N_3478,N_4084);
nor U5855 (N_5855,N_1416,N_2781);
or U5856 (N_5856,N_1762,N_4715);
xnor U5857 (N_5857,N_4948,N_1032);
nand U5858 (N_5858,N_1362,N_4737);
nand U5859 (N_5859,N_1456,N_1433);
nand U5860 (N_5860,N_4694,N_723);
nor U5861 (N_5861,N_3517,N_763);
or U5862 (N_5862,N_1604,N_4458);
nor U5863 (N_5863,N_2137,N_79);
and U5864 (N_5864,N_2905,N_4193);
nand U5865 (N_5865,N_4259,N_776);
nand U5866 (N_5866,N_2926,N_1795);
or U5867 (N_5867,N_1240,N_1440);
nor U5868 (N_5868,N_2366,N_934);
and U5869 (N_5869,N_2951,N_3172);
and U5870 (N_5870,N_3375,N_1876);
nand U5871 (N_5871,N_4174,N_1358);
and U5872 (N_5872,N_4288,N_1608);
nand U5873 (N_5873,N_1740,N_1144);
nor U5874 (N_5874,N_2091,N_67);
and U5875 (N_5875,N_1353,N_963);
nor U5876 (N_5876,N_4,N_4360);
nor U5877 (N_5877,N_3942,N_1843);
nand U5878 (N_5878,N_353,N_1626);
and U5879 (N_5879,N_4311,N_3353);
and U5880 (N_5880,N_3627,N_2999);
nand U5881 (N_5881,N_3896,N_3525);
nand U5882 (N_5882,N_3374,N_1899);
nand U5883 (N_5883,N_4514,N_4805);
nand U5884 (N_5884,N_4797,N_1788);
nand U5885 (N_5885,N_1828,N_3491);
and U5886 (N_5886,N_4789,N_4369);
nand U5887 (N_5887,N_3463,N_3171);
and U5888 (N_5888,N_3337,N_1197);
or U5889 (N_5889,N_610,N_1359);
nor U5890 (N_5890,N_885,N_1662);
nor U5891 (N_5891,N_3873,N_1385);
nor U5892 (N_5892,N_3737,N_4457);
and U5893 (N_5893,N_643,N_4548);
nor U5894 (N_5894,N_2409,N_3998);
nand U5895 (N_5895,N_292,N_1307);
or U5896 (N_5896,N_1382,N_3988);
nand U5897 (N_5897,N_4685,N_1732);
nand U5898 (N_5898,N_4692,N_1572);
and U5899 (N_5899,N_1335,N_4316);
nor U5900 (N_5900,N_681,N_930);
nand U5901 (N_5901,N_3704,N_4503);
nand U5902 (N_5902,N_2487,N_2289);
nand U5903 (N_5903,N_2693,N_3759);
nand U5904 (N_5904,N_114,N_4874);
and U5905 (N_5905,N_4358,N_4290);
xnor U5906 (N_5906,N_2826,N_3297);
or U5907 (N_5907,N_1133,N_3577);
nor U5908 (N_5908,N_2987,N_1512);
and U5909 (N_5909,N_3978,N_427);
nor U5910 (N_5910,N_2649,N_646);
or U5911 (N_5911,N_4965,N_3855);
nand U5912 (N_5912,N_2868,N_4507);
nor U5913 (N_5913,N_332,N_38);
nand U5914 (N_5914,N_1928,N_170);
and U5915 (N_5915,N_1945,N_3217);
nor U5916 (N_5916,N_2697,N_632);
nor U5917 (N_5917,N_3009,N_4819);
and U5918 (N_5918,N_4071,N_1408);
and U5919 (N_5919,N_1046,N_4988);
nand U5920 (N_5920,N_2634,N_3321);
and U5921 (N_5921,N_960,N_3);
or U5922 (N_5922,N_4880,N_1879);
nor U5923 (N_5923,N_149,N_1033);
nor U5924 (N_5924,N_590,N_4713);
and U5925 (N_5925,N_1575,N_1429);
or U5926 (N_5926,N_1268,N_2111);
and U5927 (N_5927,N_697,N_4598);
nand U5928 (N_5928,N_3025,N_1953);
nor U5929 (N_5929,N_4634,N_976);
and U5930 (N_5930,N_2597,N_4724);
nand U5931 (N_5931,N_1596,N_320);
nand U5932 (N_5932,N_4070,N_3829);
nand U5933 (N_5933,N_1984,N_268);
and U5934 (N_5934,N_3976,N_1786);
and U5935 (N_5935,N_2855,N_3595);
and U5936 (N_5936,N_3126,N_4592);
and U5937 (N_5937,N_1428,N_2829);
nor U5938 (N_5938,N_2222,N_28);
or U5939 (N_5939,N_586,N_2134);
or U5940 (N_5940,N_4377,N_4023);
or U5941 (N_5941,N_4796,N_1808);
nand U5942 (N_5942,N_3040,N_4386);
nand U5943 (N_5943,N_2464,N_1286);
or U5944 (N_5944,N_198,N_3114);
and U5945 (N_5945,N_123,N_3693);
or U5946 (N_5946,N_1165,N_2736);
and U5947 (N_5947,N_720,N_4747);
and U5948 (N_5948,N_2270,N_1272);
nand U5949 (N_5949,N_1810,N_1475);
and U5950 (N_5950,N_1863,N_1231);
nor U5951 (N_5951,N_4376,N_1010);
nand U5952 (N_5952,N_4095,N_1656);
nand U5953 (N_5953,N_4524,N_2927);
and U5954 (N_5954,N_70,N_4185);
or U5955 (N_5955,N_1030,N_4647);
nand U5956 (N_5956,N_2327,N_4765);
or U5957 (N_5957,N_1661,N_928);
or U5958 (N_5958,N_1306,N_3432);
and U5959 (N_5959,N_4682,N_2777);
or U5960 (N_5960,N_3993,N_1793);
and U5961 (N_5961,N_4527,N_420);
and U5962 (N_5962,N_4494,N_3650);
nor U5963 (N_5963,N_1836,N_3320);
or U5964 (N_5964,N_2298,N_4050);
nor U5965 (N_5965,N_3128,N_4472);
nand U5966 (N_5966,N_703,N_2773);
nand U5967 (N_5967,N_4344,N_2988);
or U5968 (N_5968,N_4586,N_2774);
nand U5969 (N_5969,N_312,N_3121);
or U5970 (N_5970,N_4086,N_2180);
nor U5971 (N_5971,N_2595,N_823);
nor U5972 (N_5972,N_428,N_99);
and U5973 (N_5973,N_1610,N_2238);
and U5974 (N_5974,N_1372,N_3190);
nand U5975 (N_5975,N_3326,N_2661);
and U5976 (N_5976,N_3037,N_975);
and U5977 (N_5977,N_326,N_2354);
nor U5978 (N_5978,N_1521,N_76);
and U5979 (N_5979,N_1893,N_483);
and U5980 (N_5980,N_1140,N_2113);
and U5981 (N_5981,N_284,N_1994);
nand U5982 (N_5982,N_2880,N_913);
and U5983 (N_5983,N_652,N_1897);
or U5984 (N_5984,N_1081,N_4398);
and U5985 (N_5985,N_3144,N_2492);
nand U5986 (N_5986,N_3947,N_1082);
nor U5987 (N_5987,N_2085,N_1115);
nand U5988 (N_5988,N_748,N_3920);
or U5989 (N_5989,N_275,N_2949);
nand U5990 (N_5990,N_4052,N_2979);
or U5991 (N_5991,N_211,N_386);
nand U5992 (N_5992,N_2528,N_3583);
xnor U5993 (N_5993,N_266,N_3549);
or U5994 (N_5994,N_471,N_3315);
nand U5995 (N_5995,N_2449,N_271);
or U5996 (N_5996,N_4629,N_2991);
nor U5997 (N_5997,N_2887,N_805);
nand U5998 (N_5998,N_1804,N_3425);
nand U5999 (N_5999,N_4539,N_2585);
and U6000 (N_6000,N_161,N_3964);
or U6001 (N_6001,N_4309,N_3499);
or U6002 (N_6002,N_4064,N_4559);
or U6003 (N_6003,N_4497,N_3844);
or U6004 (N_6004,N_3545,N_3462);
nor U6005 (N_6005,N_4044,N_2923);
nand U6006 (N_6006,N_2043,N_2694);
and U6007 (N_6007,N_1675,N_1597);
nor U6008 (N_6008,N_3263,N_1862);
nor U6009 (N_6009,N_1517,N_240);
nor U6010 (N_6010,N_4444,N_1577);
and U6011 (N_6011,N_3113,N_2135);
and U6012 (N_6012,N_1919,N_4981);
and U6013 (N_6013,N_1355,N_1038);
nand U6014 (N_6014,N_4186,N_1504);
and U6015 (N_6015,N_1613,N_2460);
or U6016 (N_6016,N_1767,N_1099);
and U6017 (N_6017,N_1659,N_2303);
and U6018 (N_6018,N_2919,N_57);
or U6019 (N_6019,N_3606,N_4034);
nor U6020 (N_6020,N_2805,N_1437);
nand U6021 (N_6021,N_2225,N_1995);
nand U6022 (N_6022,N_3571,N_273);
and U6023 (N_6023,N_3493,N_294);
nor U6024 (N_6024,N_2155,N_1403);
or U6025 (N_6025,N_1147,N_2323);
and U6026 (N_6026,N_4515,N_1290);
nand U6027 (N_6027,N_2167,N_2244);
nand U6028 (N_6028,N_1360,N_2506);
nor U6029 (N_6029,N_4917,N_2854);
nor U6030 (N_6030,N_4406,N_3555);
and U6031 (N_6031,N_927,N_4741);
or U6032 (N_6032,N_2146,N_1194);
xnor U6033 (N_6033,N_2416,N_1946);
nand U6034 (N_6034,N_2813,N_3354);
nor U6035 (N_6035,N_571,N_2474);
nor U6036 (N_6036,N_2834,N_523);
nand U6037 (N_6037,N_4813,N_3897);
nor U6038 (N_6038,N_2068,N_962);
nor U6039 (N_6039,N_4597,N_2531);
nand U6040 (N_6040,N_2490,N_4445);
or U6041 (N_6041,N_3067,N_1254);
nand U6042 (N_6042,N_2254,N_95);
or U6043 (N_6043,N_2062,N_1247);
nor U6044 (N_6044,N_3254,N_3861);
or U6045 (N_6045,N_4384,N_3312);
or U6046 (N_6046,N_1262,N_2957);
or U6047 (N_6047,N_2665,N_248);
nand U6048 (N_6048,N_3558,N_1944);
nand U6049 (N_6049,N_3647,N_3638);
or U6050 (N_6050,N_3710,N_2573);
nand U6051 (N_6051,N_3561,N_2600);
and U6052 (N_6052,N_3069,N_1333);
nand U6053 (N_6053,N_3150,N_4902);
nand U6054 (N_6054,N_2423,N_3282);
nand U6055 (N_6055,N_615,N_4032);
or U6056 (N_6056,N_4301,N_2744);
or U6057 (N_6057,N_942,N_1417);
nand U6058 (N_6058,N_4226,N_2705);
nand U6059 (N_6059,N_377,N_3238);
and U6060 (N_6060,N_852,N_4585);
or U6061 (N_6061,N_1637,N_163);
nand U6062 (N_6062,N_397,N_4317);
nor U6063 (N_6063,N_4963,N_947);
or U6064 (N_6064,N_63,N_3062);
nand U6065 (N_6065,N_845,N_1847);
or U6066 (N_6066,N_2405,N_3860);
and U6067 (N_6067,N_2014,N_4164);
nand U6068 (N_6068,N_4840,N_4189);
nand U6069 (N_6069,N_3268,N_981);
nor U6070 (N_6070,N_3482,N_2547);
nor U6071 (N_6071,N_1193,N_3146);
nor U6072 (N_6072,N_3730,N_385);
nand U6073 (N_6073,N_3329,N_2404);
or U6074 (N_6074,N_3645,N_1198);
or U6075 (N_6075,N_1665,N_1917);
nand U6076 (N_6076,N_3922,N_4640);
nor U6077 (N_6077,N_869,N_4228);
and U6078 (N_6078,N_2315,N_4841);
nand U6079 (N_6079,N_3641,N_796);
or U6080 (N_6080,N_1206,N_2601);
nor U6081 (N_6081,N_4080,N_1652);
or U6082 (N_6082,N_2360,N_2538);
or U6083 (N_6083,N_3366,N_415);
nor U6084 (N_6084,N_3858,N_888);
and U6085 (N_6085,N_1253,N_4509);
and U6086 (N_6086,N_1807,N_1438);
and U6087 (N_6087,N_4136,N_3646);
and U6088 (N_6088,N_1674,N_3336);
and U6089 (N_6089,N_627,N_3490);
and U6090 (N_6090,N_2782,N_2550);
nand U6091 (N_6091,N_3660,N_698);
or U6092 (N_6092,N_3495,N_1509);
or U6093 (N_6093,N_4999,N_394);
and U6094 (N_6094,N_836,N_1923);
or U6095 (N_6095,N_3827,N_4104);
or U6096 (N_6096,N_4477,N_4622);
and U6097 (N_6097,N_745,N_625);
and U6098 (N_6098,N_3800,N_110);
or U6099 (N_6099,N_156,N_773);
or U6100 (N_6100,N_4399,N_277);
xnor U6101 (N_6101,N_2637,N_1409);
or U6102 (N_6102,N_94,N_410);
or U6103 (N_6103,N_2745,N_435);
and U6104 (N_6104,N_4596,N_1132);
or U6105 (N_6105,N_1313,N_4767);
and U6106 (N_6106,N_1350,N_3426);
and U6107 (N_6107,N_1683,N_1895);
and U6108 (N_6108,N_2321,N_781);
and U6109 (N_6109,N_405,N_666);
nor U6110 (N_6110,N_4137,N_3910);
nand U6111 (N_6111,N_3250,N_2230);
and U6112 (N_6112,N_4570,N_2019);
nand U6113 (N_6113,N_4654,N_3465);
or U6114 (N_6114,N_599,N_4711);
or U6115 (N_6115,N_3153,N_1669);
or U6116 (N_6116,N_2453,N_3223);
nand U6117 (N_6117,N_459,N_3436);
nor U6118 (N_6118,N_3591,N_1557);
nor U6119 (N_6119,N_2300,N_1364);
or U6120 (N_6120,N_3189,N_2431);
and U6121 (N_6121,N_4910,N_3390);
or U6122 (N_6122,N_3397,N_1209);
nor U6123 (N_6123,N_2896,N_2677);
or U6124 (N_6124,N_2644,N_941);
nor U6125 (N_6125,N_2771,N_2148);
and U6126 (N_6126,N_1483,N_3687);
nor U6127 (N_6127,N_3842,N_1244);
or U6128 (N_6128,N_4868,N_487);
or U6129 (N_6129,N_2496,N_4979);
nand U6130 (N_6130,N_2324,N_622);
xor U6131 (N_6131,N_3019,N_921);
nor U6132 (N_6132,N_4057,N_4068);
nor U6133 (N_6133,N_2518,N_3398);
or U6134 (N_6134,N_3272,N_261);
or U6135 (N_6135,N_830,N_2750);
or U6136 (N_6136,N_4037,N_4860);
nor U6137 (N_6137,N_994,N_3832);
nand U6138 (N_6138,N_4473,N_3999);
and U6139 (N_6139,N_585,N_4991);
nor U6140 (N_6140,N_448,N_613);
nand U6141 (N_6141,N_2396,N_537);
or U6142 (N_6142,N_3136,N_871);
and U6143 (N_6143,N_4582,N_2408);
and U6144 (N_6144,N_2612,N_1523);
or U6145 (N_6145,N_4913,N_2520);
nor U6146 (N_6146,N_2284,N_3328);
and U6147 (N_6147,N_1100,N_218);
nand U6148 (N_6148,N_3707,N_4390);
nand U6149 (N_6149,N_189,N_1239);
or U6150 (N_6150,N_1026,N_4243);
nor U6151 (N_6151,N_609,N_4074);
nor U6152 (N_6152,N_2725,N_1448);
or U6153 (N_6153,N_1565,N_3435);
or U6154 (N_6154,N_4014,N_4818);
and U6155 (N_6155,N_1985,N_117);
nand U6156 (N_6156,N_2791,N_3157);
nand U6157 (N_6157,N_3452,N_3215);
nor U6158 (N_6158,N_3689,N_498);
or U6159 (N_6159,N_227,N_4712);
nand U6160 (N_6160,N_1241,N_1858);
or U6161 (N_6161,N_3154,N_2732);
nor U6162 (N_6162,N_4884,N_2079);
and U6163 (N_6163,N_3698,N_1819);
nand U6164 (N_6164,N_4227,N_4169);
nand U6165 (N_6165,N_2391,N_4986);
and U6166 (N_6166,N_2101,N_2191);
nor U6167 (N_6167,N_45,N_2394);
nor U6168 (N_6168,N_4362,N_2185);
and U6169 (N_6169,N_647,N_1541);
nor U6170 (N_6170,N_3790,N_4564);
nor U6171 (N_6171,N_1942,N_3300);
and U6172 (N_6172,N_1015,N_3711);
or U6173 (N_6173,N_929,N_1278);
and U6174 (N_6174,N_4355,N_3416);
or U6175 (N_6175,N_4441,N_2145);
nor U6176 (N_6176,N_4734,N_1609);
or U6177 (N_6177,N_3864,N_4659);
or U6178 (N_6178,N_317,N_2401);
or U6179 (N_6179,N_3880,N_1800);
nor U6180 (N_6180,N_863,N_2114);
nor U6181 (N_6181,N_2992,N_3058);
and U6182 (N_6182,N_3974,N_154);
nor U6183 (N_6183,N_2117,N_3256);
nand U6184 (N_6184,N_3492,N_1780);
nand U6185 (N_6185,N_4442,N_3934);
nand U6186 (N_6186,N_2967,N_1005);
nand U6187 (N_6187,N_3705,N_4688);
or U6188 (N_6188,N_3892,N_1616);
or U6189 (N_6189,N_1496,N_1043);
nand U6190 (N_6190,N_2643,N_1464);
nor U6191 (N_6191,N_2273,N_2630);
and U6192 (N_6192,N_683,N_4944);
and U6193 (N_6193,N_2005,N_3246);
or U6194 (N_6194,N_8,N_1356);
nand U6195 (N_6195,N_1019,N_2080);
or U6196 (N_6196,N_991,N_3001);
nand U6197 (N_6197,N_987,N_1833);
and U6198 (N_6198,N_3045,N_3098);
xor U6199 (N_6199,N_112,N_2126);
nand U6200 (N_6200,N_3338,N_4746);
nand U6201 (N_6201,N_2976,N_3868);
and U6202 (N_6202,N_3913,N_870);
or U6203 (N_6203,N_778,N_4114);
or U6204 (N_6204,N_3685,N_2293);
or U6205 (N_6205,N_1368,N_699);
or U6206 (N_6206,N_3016,N_4165);
nor U6207 (N_6207,N_3831,N_391);
and U6208 (N_6208,N_4782,N_2966);
and U6209 (N_6209,N_1829,N_1370);
or U6210 (N_6210,N_3539,N_182);
nand U6211 (N_6211,N_3603,N_4278);
or U6212 (N_6212,N_575,N_3662);
nand U6213 (N_6213,N_1770,N_883);
nor U6214 (N_6214,N_4166,N_2864);
nand U6215 (N_6215,N_1749,N_2915);
nor U6216 (N_6216,N_3782,N_731);
or U6217 (N_6217,N_1905,N_2944);
nor U6218 (N_6218,N_159,N_1014);
nor U6219 (N_6219,N_690,N_4636);
or U6220 (N_6220,N_4462,N_3226);
nor U6221 (N_6221,N_4706,N_378);
or U6222 (N_6222,N_2092,N_838);
nand U6223 (N_6223,N_3579,N_1432);
nand U6224 (N_6224,N_2898,N_2795);
and U6225 (N_6225,N_1785,N_2318);
nor U6226 (N_6226,N_2841,N_10);
nor U6227 (N_6227,N_4036,N_2407);
and U6228 (N_6228,N_440,N_4687);
or U6229 (N_6229,N_501,N_3111);
or U6230 (N_6230,N_3640,N_3866);
and U6231 (N_6231,N_1080,N_3601);
nor U6232 (N_6232,N_1713,N_4357);
and U6233 (N_6233,N_4146,N_3137);
or U6234 (N_6234,N_1934,N_1959);
and U6235 (N_6235,N_482,N_1117);
or U6236 (N_6236,N_1736,N_2609);
or U6237 (N_6237,N_2755,N_1476);
nand U6238 (N_6238,N_736,N_4313);
and U6239 (N_6239,N_2857,N_1109);
nor U6240 (N_6240,N_4030,N_2013);
and U6241 (N_6241,N_2165,N_4056);
and U6242 (N_6242,N_4078,N_3783);
nor U6243 (N_6243,N_2204,N_2663);
or U6244 (N_6244,N_3203,N_84);
and U6245 (N_6245,N_4951,N_3632);
nor U6246 (N_6246,N_3059,N_103);
nor U6247 (N_6247,N_2990,N_2833);
or U6248 (N_6248,N_1734,N_1927);
and U6249 (N_6249,N_4267,N_2679);
or U6250 (N_6250,N_1587,N_3655);
or U6251 (N_6251,N_2962,N_3686);
or U6252 (N_6252,N_402,N_629);
nand U6253 (N_6253,N_338,N_3757);
and U6254 (N_6254,N_4888,N_4083);
or U6255 (N_6255,N_951,N_967);
and U6256 (N_6256,N_449,N_1103);
nor U6257 (N_6257,N_3903,N_1031);
or U6258 (N_6258,N_2026,N_3003);
nand U6259 (N_6259,N_4182,N_596);
and U6260 (N_6260,N_1275,N_4139);
or U6261 (N_6261,N_47,N_4431);
nor U6262 (N_6262,N_3975,N_4925);
nor U6263 (N_6263,N_4587,N_2766);
nand U6264 (N_6264,N_2494,N_3817);
and U6265 (N_6265,N_607,N_4930);
nor U6266 (N_6266,N_2638,N_3498);
and U6267 (N_6267,N_506,N_1978);
nand U6268 (N_6268,N_107,N_4199);
nand U6269 (N_6269,N_611,N_4914);
nand U6270 (N_6270,N_1489,N_503);
or U6271 (N_6271,N_3677,N_4809);
or U6272 (N_6272,N_153,N_290);
nor U6273 (N_6273,N_714,N_429);
nand U6274 (N_6274,N_3350,N_4466);
nor U6275 (N_6275,N_770,N_4414);
nand U6276 (N_6276,N_968,N_3064);
and U6277 (N_6277,N_618,N_3950);
nor U6278 (N_6278,N_3285,N_4798);
and U6279 (N_6279,N_514,N_3749);
and U6280 (N_6280,N_4475,N_1702);
xor U6281 (N_6281,N_4698,N_3393);
nor U6282 (N_6282,N_1671,N_879);
and U6283 (N_6283,N_3073,N_3862);
and U6284 (N_6284,N_1717,N_3381);
or U6285 (N_6285,N_4644,N_1480);
xnor U6286 (N_6286,N_4194,N_2893);
nor U6287 (N_6287,N_1518,N_458);
nor U6288 (N_6288,N_1799,N_128);
or U6289 (N_6289,N_2624,N_2175);
nand U6290 (N_6290,N_2590,N_4420);
xor U6291 (N_6291,N_1564,N_3639);
nand U6292 (N_6292,N_4777,N_569);
nand U6293 (N_6293,N_1389,N_702);
or U6294 (N_6294,N_1091,N_1993);
or U6295 (N_6295,N_3348,N_1933);
or U6296 (N_6296,N_1375,N_3870);
or U6297 (N_6297,N_2475,N_3765);
nand U6298 (N_6298,N_3936,N_1650);
nor U6299 (N_6299,N_827,N_1617);
nand U6300 (N_6300,N_2313,N_2607);
nor U6301 (N_6301,N_1666,N_2454);
or U6302 (N_6302,N_3929,N_3507);
nor U6303 (N_6303,N_1991,N_1792);
or U6304 (N_6304,N_1224,N_589);
nor U6305 (N_6305,N_1598,N_595);
or U6306 (N_6306,N_2451,N_1227);
nand U6307 (N_6307,N_3470,N_62);
nand U6308 (N_6308,N_2207,N_3209);
or U6309 (N_6309,N_4284,N_3609);
xnor U6310 (N_6310,N_904,N_119);
or U6311 (N_6311,N_3197,N_158);
nand U6312 (N_6312,N_4658,N_4403);
nor U6313 (N_6313,N_2371,N_1903);
nor U6314 (N_6314,N_2183,N_4238);
nor U6315 (N_6315,N_396,N_898);
or U6316 (N_6316,N_3309,N_1969);
nor U6317 (N_6317,N_4038,N_3589);
nor U6318 (N_6318,N_1508,N_2772);
and U6319 (N_6319,N_1654,N_4745);
nor U6320 (N_6320,N_2764,N_2296);
nor U6321 (N_6321,N_4615,N_1479);
nor U6322 (N_6322,N_1667,N_671);
nand U6323 (N_6323,N_4828,N_1768);
nand U6324 (N_6324,N_4203,N_4946);
or U6325 (N_6325,N_372,N_2334);
nor U6326 (N_6326,N_3931,N_2285);
or U6327 (N_6327,N_33,N_4623);
nor U6328 (N_6328,N_4504,N_219);
nor U6329 (N_6329,N_2090,N_1332);
nor U6330 (N_6330,N_4670,N_1873);
and U6331 (N_6331,N_1920,N_4879);
nor U6332 (N_6332,N_3956,N_39);
and U6333 (N_6333,N_4429,N_1980);
and U6334 (N_6334,N_3346,N_3582);
or U6335 (N_6335,N_2336,N_3333);
or U6336 (N_6336,N_4556,N_2261);
nand U6337 (N_6337,N_2009,N_4590);
nor U6338 (N_6338,N_1705,N_598);
or U6339 (N_6339,N_3365,N_1236);
nand U6340 (N_6340,N_3869,N_2203);
and U6341 (N_6341,N_4749,N_4975);
nor U6342 (N_6342,N_708,N_3233);
nor U6343 (N_6343,N_1685,N_145);
or U6344 (N_6344,N_1112,N_1386);
and U6345 (N_6345,N_1972,N_4364);
and U6346 (N_6346,N_2434,N_1346);
or U6347 (N_6347,N_9,N_3167);
and U6348 (N_6348,N_2351,N_3335);
nand U6349 (N_6349,N_544,N_1218);
xnor U6350 (N_6350,N_439,N_269);
and U6351 (N_6351,N_1690,N_4744);
and U6352 (N_6352,N_3318,N_3358);
nor U6353 (N_6353,N_854,N_4304);
or U6354 (N_6354,N_4707,N_2968);
nor U6355 (N_6355,N_2010,N_2156);
and U6356 (N_6356,N_339,N_2157);
nor U6357 (N_6357,N_4528,N_4937);
or U6358 (N_6358,N_1820,N_1913);
nand U6359 (N_6359,N_1463,N_457);
and U6360 (N_6360,N_1600,N_1363);
and U6361 (N_6361,N_1982,N_447);
and U6362 (N_6362,N_3404,N_1299);
and U6363 (N_6363,N_3529,N_388);
nor U6364 (N_6364,N_2115,N_4801);
nor U6365 (N_6365,N_96,N_1168);
nor U6366 (N_6366,N_4568,N_1113);
and U6367 (N_6367,N_1491,N_1854);
and U6368 (N_6368,N_3893,N_582);
xnor U6369 (N_6369,N_4794,N_2872);
and U6370 (N_6370,N_3785,N_3438);
or U6371 (N_6371,N_1570,N_4117);
nand U6372 (N_6372,N_4427,N_1138);
and U6373 (N_6373,N_2054,N_1255);
nand U6374 (N_6374,N_765,N_4962);
nand U6375 (N_6375,N_1922,N_4859);
and U6376 (N_6376,N_2443,N_1484);
nor U6377 (N_6377,N_3758,N_1716);
nor U6378 (N_6378,N_3512,N_4973);
or U6379 (N_6379,N_127,N_2998);
and U6380 (N_6380,N_4002,N_1894);
or U6381 (N_6381,N_3729,N_2447);
and U6382 (N_6382,N_3488,N_1999);
nor U6383 (N_6383,N_2614,N_4935);
or U6384 (N_6384,N_538,N_315);
nor U6385 (N_6385,N_229,N_4779);
and U6386 (N_6386,N_4751,N_2731);
xnor U6387 (N_6387,N_4655,N_488);
and U6388 (N_6388,N_2683,N_2989);
nor U6389 (N_6389,N_3828,N_3207);
and U6390 (N_6390,N_4367,N_2969);
nand U6391 (N_6391,N_1542,N_2197);
or U6392 (N_6392,N_2056,N_1857);
nor U6393 (N_6393,N_1633,N_746);
nor U6394 (N_6394,N_4330,N_1806);
nor U6395 (N_6395,N_1052,N_1724);
nand U6396 (N_6396,N_4633,N_2040);
nand U6397 (N_6397,N_208,N_1130);
nor U6398 (N_6398,N_966,N_3575);
and U6399 (N_6399,N_2186,N_1420);
or U6400 (N_6400,N_1345,N_3914);
xor U6401 (N_6401,N_2798,N_3480);
xor U6402 (N_6402,N_4001,N_4934);
nor U6403 (N_6403,N_559,N_1684);
nor U6404 (N_6404,N_2345,N_1184);
or U6405 (N_6405,N_4206,N_4334);
and U6406 (N_6406,N_476,N_3270);
nor U6407 (N_6407,N_4127,N_3485);
or U6408 (N_6408,N_1340,N_4502);
or U6409 (N_6409,N_1314,N_1627);
nand U6410 (N_6410,N_1790,N_1421);
nand U6411 (N_6411,N_3086,N_2224);
nand U6412 (N_6412,N_4349,N_175);
nand U6413 (N_6413,N_3412,N_3670);
and U6414 (N_6414,N_4761,N_4145);
nand U6415 (N_6415,N_4829,N_505);
or U6416 (N_6416,N_1778,N_3968);
or U6417 (N_6417,N_4577,N_1199);
xor U6418 (N_6418,N_3566,N_4452);
or U6419 (N_6419,N_224,N_1507);
and U6420 (N_6420,N_310,N_3503);
xnor U6421 (N_6421,N_1016,N_4496);
and U6422 (N_6422,N_1988,N_4480);
nor U6423 (N_6423,N_1931,N_1352);
nand U6424 (N_6424,N_1365,N_3423);
or U6425 (N_6425,N_3754,N_1008);
nor U6426 (N_6426,N_1395,N_1394);
nand U6427 (N_6427,N_1293,N_3992);
and U6428 (N_6428,N_1529,N_13);
nor U6429 (N_6429,N_3231,N_4109);
nand U6430 (N_6430,N_3458,N_4690);
or U6431 (N_6431,N_4915,N_3607);
and U6432 (N_6432,N_4719,N_1141);
and U6433 (N_6433,N_3851,N_4812);
and U6434 (N_6434,N_2457,N_3487);
or U6435 (N_6435,N_4039,N_3145);
nor U6436 (N_6436,N_1837,N_2711);
nor U6437 (N_6437,N_4258,N_2718);
nor U6438 (N_6438,N_2675,N_4506);
nor U6439 (N_6439,N_4978,N_258);
nand U6440 (N_6440,N_3434,N_4066);
nor U6441 (N_6441,N_3211,N_3243);
nor U6442 (N_6442,N_3056,N_3077);
nor U6443 (N_6443,N_188,N_959);
nor U6444 (N_6444,N_1150,N_1698);
or U6445 (N_6445,N_583,N_2467);
nand U6446 (N_6446,N_4987,N_133);
and U6447 (N_6447,N_165,N_689);
nand U6448 (N_6448,N_1506,N_4959);
nor U6449 (N_6449,N_3295,N_272);
nor U6450 (N_6450,N_4407,N_2659);
and U6451 (N_6451,N_3716,N_3823);
nor U6452 (N_6452,N_4606,N_3074);
nor U6453 (N_6453,N_2901,N_82);
or U6454 (N_6454,N_1126,N_1911);
nand U6455 (N_6455,N_1660,N_2828);
nor U6456 (N_6456,N_3289,N_184);
nor U6457 (N_6457,N_2779,N_4750);
nor U6458 (N_6458,N_3733,N_1390);
and U6459 (N_6459,N_3535,N_3521);
and U6460 (N_6460,N_3380,N_1331);
nor U6461 (N_6461,N_144,N_4147);
nor U6462 (N_6462,N_4283,N_719);
nand U6463 (N_6463,N_1628,N_1351);
or U6464 (N_6464,N_3183,N_3692);
nand U6465 (N_6465,N_3813,N_2753);
and U6466 (N_6466,N_484,N_3431);
nand U6467 (N_6467,N_4098,N_3986);
and U6468 (N_6468,N_2250,N_3624);
nand U6469 (N_6469,N_3299,N_540);
and U6470 (N_6470,N_4211,N_4356);
and U6471 (N_6471,N_4846,N_1722);
nand U6472 (N_6472,N_4873,N_4308);
nand U6473 (N_6473,N_2911,N_1874);
nand U6474 (N_6474,N_2237,N_3576);
nor U6475 (N_6475,N_2895,N_445);
or U6476 (N_6476,N_279,N_1183);
nand U6477 (N_6477,N_489,N_2306);
nor U6478 (N_6478,N_4153,N_2994);
or U6479 (N_6479,N_2264,N_230);
nand U6480 (N_6480,N_2497,N_2335);
nand U6481 (N_6481,N_1930,N_4337);
or U6482 (N_6482,N_2173,N_4325);
or U6483 (N_6483,N_3162,N_4320);
nor U6484 (N_6484,N_1849,N_2502);
or U6485 (N_6485,N_756,N_2511);
and U6486 (N_6486,N_481,N_203);
or U6487 (N_6487,N_152,N_2789);
or U6488 (N_6488,N_3394,N_4261);
nand U6489 (N_6489,N_4439,N_1546);
and U6490 (N_6490,N_1679,N_4802);
or U6491 (N_6491,N_1888,N_4536);
nand U6492 (N_6492,N_212,N_81);
or U6493 (N_6493,N_4878,N_2116);
nand U6494 (N_6494,N_4245,N_191);
nor U6495 (N_6495,N_4720,N_3413);
nor U6496 (N_6496,N_548,N_3152);
or U6497 (N_6497,N_494,N_1083);
or U6498 (N_6498,N_4045,N_2965);
and U6499 (N_6499,N_2020,N_1007);
and U6500 (N_6500,N_1590,N_3373);
or U6501 (N_6501,N_1522,N_1940);
and U6502 (N_6502,N_775,N_3722);
or U6503 (N_6503,N_1172,N_1304);
and U6504 (N_6504,N_4569,N_4776);
or U6505 (N_6505,N_371,N_2983);
nor U6506 (N_6506,N_3557,N_496);
nand U6507 (N_6507,N_2566,N_2700);
nand U6508 (N_6508,N_760,N_2689);
and U6509 (N_6509,N_91,N_799);
and U6510 (N_6510,N_430,N_1887);
or U6511 (N_6511,N_3454,N_2977);
nor U6512 (N_6512,N_265,N_1651);
nor U6513 (N_6513,N_4327,N_2888);
xnor U6514 (N_6514,N_955,N_2670);
nand U6515 (N_6515,N_777,N_4632);
nand U6516 (N_6516,N_4026,N_3605);
nor U6517 (N_6517,N_551,N_101);
or U6518 (N_6518,N_4231,N_4820);
nand U6519 (N_6519,N_4424,N_2529);
or U6520 (N_6520,N_4339,N_1155);
and U6521 (N_6521,N_1503,N_1189);
and U6522 (N_6522,N_580,N_1149);
and U6523 (N_6523,N_4889,N_493);
or U6524 (N_6524,N_22,N_2432);
nand U6525 (N_6525,N_1004,N_4167);
and U6526 (N_6526,N_2132,N_2015);
nor U6527 (N_6527,N_3797,N_3925);
nand U6528 (N_6528,N_2410,N_3103);
nand U6529 (N_6529,N_4696,N_4875);
nand U6530 (N_6530,N_2195,N_709);
and U6531 (N_6531,N_2200,N_874);
nor U6532 (N_6532,N_1270,N_4922);
xnor U6533 (N_6533,N_3536,N_1779);
nor U6534 (N_6534,N_1841,N_2393);
and U6535 (N_6535,N_2302,N_2792);
and U6536 (N_6536,N_264,N_3620);
nand U6537 (N_6537,N_1797,N_3789);
nand U6538 (N_6538,N_2364,N_4151);
and U6539 (N_6539,N_2379,N_624);
and U6540 (N_6540,N_1445,N_4272);
or U6541 (N_6541,N_4612,N_4995);
nor U6542 (N_6542,N_3661,N_4969);
xor U6543 (N_6543,N_680,N_2418);
and U6544 (N_6544,N_3923,N_2030);
nand U6545 (N_6545,N_1303,N_3915);
and U6546 (N_6546,N_1548,N_1090);
and U6547 (N_6547,N_3070,N_1361);
and U6548 (N_6548,N_1024,N_4040);
nor U6549 (N_6549,N_4865,N_876);
or U6550 (N_6550,N_657,N_1505);
nor U6551 (N_6551,N_1677,N_1916);
nor U6552 (N_6552,N_4638,N_2096);
nand U6553 (N_6553,N_4912,N_701);
nand U6554 (N_6554,N_3092,N_4571);
nor U6555 (N_6555,N_1950,N_4565);
nand U6556 (N_6556,N_4361,N_4125);
nor U6557 (N_6557,N_1952,N_2168);
nor U6558 (N_6558,N_2875,N_4374);
nand U6559 (N_6559,N_3613,N_233);
or U6560 (N_6560,N_3546,N_3863);
nand U6561 (N_6561,N_1532,N_2462);
xnor U6562 (N_6562,N_2433,N_3479);
nor U6563 (N_6563,N_3010,N_376);
or U6564 (N_6564,N_2048,N_4154);
and U6565 (N_6565,N_895,N_1200);
nand U6566 (N_6566,N_946,N_2548);
nor U6567 (N_6567,N_4168,N_406);
and U6568 (N_6568,N_2472,N_4129);
nor U6569 (N_6569,N_2903,N_1595);
and U6570 (N_6570,N_3115,N_3565);
and U6571 (N_6571,N_4997,N_3568);
and U6572 (N_6572,N_4827,N_3982);
and U6573 (N_6573,N_4909,N_2978);
or U6574 (N_6574,N_1207,N_3904);
or U6575 (N_6575,N_4588,N_2050);
nor U6576 (N_6576,N_4535,N_1223);
and U6577 (N_6577,N_2626,N_4573);
nand U6578 (N_6578,N_2740,N_4244);
and U6579 (N_6579,N_4106,N_740);
nor U6580 (N_6580,N_3357,N_4102);
or U6581 (N_6581,N_1941,N_816);
or U6582 (N_6582,N_1310,N_155);
nand U6583 (N_6583,N_2654,N_1171);
or U6584 (N_6584,N_2860,N_3523);
or U6585 (N_6585,N_906,N_4305);
or U6586 (N_6586,N_4985,N_2662);
and U6587 (N_6587,N_1152,N_2188);
and U6588 (N_6588,N_4000,N_704);
nand U6589 (N_6589,N_56,N_3251);
nor U6590 (N_6590,N_1497,N_2933);
and U6591 (N_6591,N_4775,N_4395);
and U6592 (N_6592,N_1260,N_3468);
or U6593 (N_6593,N_1574,N_667);
nor U6594 (N_6594,N_1589,N_3688);
and U6595 (N_6595,N_825,N_692);
nor U6596 (N_6596,N_3122,N_1676);
nand U6597 (N_6597,N_3363,N_2685);
nand U6598 (N_6598,N_4436,N_1049);
and U6599 (N_6599,N_3901,N_1625);
xnor U6600 (N_6600,N_1309,N_4848);
nand U6601 (N_6601,N_4508,N_4911);
or U6602 (N_6602,N_772,N_3902);
or U6603 (N_6603,N_3804,N_3096);
nor U6604 (N_6604,N_2645,N_3597);
xor U6605 (N_6605,N_686,N_1566);
nor U6606 (N_6606,N_3791,N_4762);
and U6607 (N_6607,N_965,N_3134);
nand U6608 (N_6608,N_461,N_4347);
nor U6609 (N_6609,N_4619,N_19);
and U6610 (N_6610,N_243,N_2169);
nor U6611 (N_6611,N_2505,N_642);
nor U6612 (N_6612,N_2012,N_4212);
nor U6613 (N_6613,N_4689,N_1629);
or U6614 (N_6614,N_186,N_3060);
nand U6615 (N_6615,N_4195,N_2139);
nor U6616 (N_6616,N_4620,N_3317);
or U6617 (N_6617,N_2651,N_1279);
and U6618 (N_6618,N_1499,N_251);
nor U6619 (N_6619,N_3410,N_2086);
nor U6620 (N_6620,N_2130,N_4907);
nand U6621 (N_6621,N_15,N_3164);
nor U6622 (N_6622,N_4112,N_4669);
nand U6623 (N_6623,N_3097,N_2527);
and U6624 (N_6624,N_803,N_2796);
nand U6625 (N_6625,N_1756,N_4460);
nand U6626 (N_6626,N_2367,N_832);
and U6627 (N_6627,N_4816,N_2691);
xor U6628 (N_6628,N_4482,N_2932);
or U6629 (N_6629,N_1281,N_232);
or U6630 (N_6630,N_3118,N_4984);
or U6631 (N_6631,N_4418,N_3667);
and U6632 (N_6632,N_1045,N_3885);
nand U6633 (N_6633,N_1694,N_2344);
or U6634 (N_6634,N_239,N_1302);
or U6635 (N_6635,N_4806,N_3184);
nor U6636 (N_6636,N_323,N_1642);
nand U6637 (N_6637,N_621,N_4020);
and U6638 (N_6638,N_2778,N_174);
nor U6639 (N_6639,N_1459,N_1451);
nand U6640 (N_6640,N_1936,N_3699);
xnor U6641 (N_6641,N_4661,N_2381);
nor U6642 (N_6642,N_3921,N_1156);
nor U6643 (N_6643,N_4940,N_755);
nor U6644 (N_6644,N_3108,N_1131);
nor U6645 (N_6645,N_412,N_3626);
and U6646 (N_6646,N_2743,N_29);
nand U6647 (N_6647,N_2974,N_4218);
nand U6648 (N_6648,N_3344,N_2542);
and U6649 (N_6649,N_1460,N_1815);
nor U6650 (N_6650,N_3221,N_4240);
nor U6651 (N_6651,N_1058,N_2543);
nand U6652 (N_6652,N_1037,N_834);
or U6653 (N_6653,N_4876,N_4837);
nor U6654 (N_6654,N_656,N_2832);
and U6655 (N_6655,N_1056,N_848);
nor U6656 (N_6656,N_2471,N_3149);
xor U6657 (N_6657,N_597,N_2192);
and U6658 (N_6658,N_4027,N_2815);
or U6659 (N_6659,N_1966,N_1029);
and U6660 (N_6660,N_4855,N_2714);
nor U6661 (N_6661,N_3083,N_3035);
and U6662 (N_6662,N_2823,N_4094);
nand U6663 (N_6663,N_1935,N_1802);
and U6664 (N_6664,N_4673,N_486);
or U6665 (N_6665,N_3732,N_4013);
nor U6666 (N_6666,N_4945,N_255);
or U6667 (N_6667,N_285,N_226);
nor U6668 (N_6668,N_4923,N_2581);
nand U6669 (N_6669,N_1668,N_948);
nand U6670 (N_6670,N_983,N_1106);
nand U6671 (N_6671,N_3314,N_2972);
or U6672 (N_6672,N_4260,N_3799);
or U6673 (N_6673,N_843,N_721);
nor U6674 (N_6674,N_4159,N_4511);
nand U6675 (N_6675,N_108,N_3472);
nor U6676 (N_6676,N_2212,N_4760);
or U6677 (N_6677,N_3208,N_2082);
and U6678 (N_6678,N_3034,N_3917);
and U6679 (N_6679,N_2580,N_3386);
and U6680 (N_6680,N_3666,N_2002);
nand U6681 (N_6681,N_3334,N_4778);
nor U6682 (N_6682,N_4621,N_1289);
nor U6683 (N_6683,N_138,N_2716);
nand U6684 (N_6684,N_654,N_1384);
xor U6685 (N_6685,N_3486,N_4385);
and U6686 (N_6686,N_3937,N_4342);
nor U6687 (N_6687,N_463,N_2602);
or U6688 (N_6688,N_648,N_2727);
and U6689 (N_6689,N_2035,N_1783);
or U6690 (N_6690,N_1569,N_2430);
nor U6691 (N_6691,N_2820,N_916);
or U6692 (N_6692,N_2761,N_4560);
nor U6693 (N_6693,N_2929,N_2095);
or U6694 (N_6694,N_853,N_3331);
nand U6695 (N_6695,N_2392,N_2319);
nand U6696 (N_6696,N_3072,N_2557);
and U6697 (N_6697,N_2017,N_1998);
and U6698 (N_6698,N_737,N_2214);
nor U6699 (N_6699,N_511,N_3138);
or U6700 (N_6700,N_3708,N_649);
nor U6701 (N_6701,N_3065,N_2184);
nand U6702 (N_6702,N_1148,N_3895);
nand U6703 (N_6703,N_1406,N_563);
or U6704 (N_6704,N_626,N_1682);
or U6705 (N_6705,N_2842,N_1576);
or U6706 (N_6706,N_2930,N_4108);
or U6707 (N_6707,N_4135,N_3292);
nor U6708 (N_6708,N_3712,N_769);
nand U6709 (N_6709,N_267,N_4149);
nand U6710 (N_6710,N_2713,N_824);
nand U6711 (N_6711,N_2658,N_1949);
nand U6712 (N_6712,N_4287,N_2971);
nand U6713 (N_6713,N_2125,N_4793);
and U6714 (N_6714,N_550,N_2631);
and U6715 (N_6715,N_2316,N_3612);
nand U6716 (N_6716,N_404,N_4433);
and U6717 (N_6717,N_918,N_3781);
nand U6718 (N_6718,N_1834,N_2347);
nor U6719 (N_6719,N_1653,N_3933);
and U6720 (N_6720,N_1242,N_1886);
nand U6721 (N_6721,N_3178,N_1704);
and U6722 (N_6722,N_887,N_3935);
and U6723 (N_6723,N_3229,N_3433);
and U6724 (N_6724,N_3135,N_2817);
and U6725 (N_6725,N_4484,N_517);
and U6726 (N_6726,N_349,N_547);
nor U6727 (N_6727,N_4348,N_2904);
nor U6728 (N_6728,N_1910,N_3881);
or U6729 (N_6729,N_1035,N_2797);
nor U6730 (N_6730,N_2970,N_200);
or U6731 (N_6731,N_3280,N_3068);
nand U6732 (N_6732,N_4666,N_1534);
nor U6733 (N_6733,N_3581,N_774);
and U6734 (N_6734,N_4141,N_4804);
nor U6735 (N_6735,N_1801,N_2307);
or U6736 (N_6736,N_3578,N_4672);
or U6737 (N_6737,N_4645,N_4345);
nor U6738 (N_6738,N_1412,N_206);
or U6739 (N_6739,N_4602,N_2283);
and U6740 (N_6740,N_1175,N_2671);
nand U6741 (N_6741,N_4251,N_3520);
nor U6742 (N_6742,N_2159,N_2688);
nor U6743 (N_6743,N_34,N_4082);
or U6744 (N_6744,N_3531,N_2150);
or U6745 (N_6745,N_3834,N_423);
nor U6746 (N_6746,N_995,N_564);
nand U6747 (N_6747,N_2687,N_3997);
xor U6748 (N_6748,N_4572,N_55);
nor U6749 (N_6749,N_3696,N_4679);
or U6750 (N_6750,N_1055,N_4530);
nand U6751 (N_6751,N_1859,N_4402);
nor U6752 (N_6752,N_788,N_2075);
or U6753 (N_6753,N_4933,N_886);
nor U6754 (N_6754,N_3691,N_2605);
nor U6755 (N_6755,N_761,N_2913);
nand U6756 (N_6756,N_1011,N_1435);
nand U6757 (N_6757,N_441,N_1908);
nor U6758 (N_6758,N_4808,N_3100);
or U6759 (N_6759,N_1453,N_1525);
and U6760 (N_6760,N_4650,N_83);
and U6761 (N_6761,N_2591,N_280);
nor U6762 (N_6762,N_2770,N_2001);
or U6763 (N_6763,N_4254,N_4380);
nor U6764 (N_6764,N_3909,N_1869);
and U6765 (N_6765,N_574,N_4191);
or U6766 (N_6766,N_1498,N_1907);
or U6767 (N_6767,N_811,N_2007);
nor U6768 (N_6768,N_2045,N_1264);
or U6769 (N_6769,N_560,N_2950);
and U6770 (N_6770,N_4275,N_2808);
and U6771 (N_6771,N_2274,N_2065);
nor U6772 (N_6772,N_1513,N_2446);
nand U6773 (N_6773,N_1377,N_3651);
nand U6774 (N_6774,N_1186,N_1515);
nor U6775 (N_6775,N_313,N_2128);
nand U6776 (N_6776,N_1225,N_2939);
nand U6777 (N_6777,N_3628,N_1844);
or U6778 (N_6778,N_3252,N_1210);
and U6779 (N_6779,N_850,N_1664);
or U6780 (N_6780,N_456,N_115);
or U6781 (N_6781,N_2757,N_1018);
nor U6782 (N_6782,N_291,N_3041);
or U6783 (N_6783,N_3275,N_3714);
nor U6784 (N_6784,N_527,N_2809);
nor U6785 (N_6785,N_1678,N_3874);
nor U6786 (N_6786,N_146,N_1646);
nand U6787 (N_6787,N_3949,N_1398);
nor U6788 (N_6788,N_2248,N_2123);
or U6789 (N_6789,N_2107,N_252);
and U6790 (N_6790,N_4748,N_336);
nor U6791 (N_6791,N_2739,N_1073);
and U6792 (N_6792,N_4175,N_1410);
or U6793 (N_6793,N_1280,N_3008);
and U6794 (N_6794,N_754,N_1388);
and U6795 (N_6795,N_1842,N_3690);
or U6796 (N_6796,N_2587,N_444);
and U6797 (N_6797,N_1769,N_2445);
and U6798 (N_6798,N_4553,N_1317);
nand U6799 (N_6799,N_4982,N_601);
nor U6800 (N_6800,N_3719,N_3664);
and U6801 (N_6801,N_4677,N_4246);
nand U6802 (N_6802,N_2788,N_4183);
nor U6803 (N_6803,N_4667,N_4882);
nand U6804 (N_6804,N_3237,N_4942);
or U6805 (N_6805,N_2674,N_4216);
and U6806 (N_6806,N_831,N_4872);
nor U6807 (N_6807,N_713,N_257);
nor U6808 (N_6808,N_1530,N_3778);
nor U6809 (N_6809,N_1047,N_2287);
or U6810 (N_6810,N_4383,N_619);
or U6811 (N_6811,N_3694,N_555);
or U6812 (N_6812,N_4838,N_2869);
and U6813 (N_6813,N_177,N_1291);
nor U6814 (N_6814,N_1890,N_4152);
nor U6815 (N_6815,N_1447,N_3747);
nor U6816 (N_6816,N_1494,N_2448);
nor U6817 (N_6817,N_1758,N_3599);
nand U6818 (N_6818,N_4382,N_74);
nand U6819 (N_6819,N_387,N_393);
or U6820 (N_6820,N_2794,N_4886);
and U6821 (N_6821,N_64,N_529);
nor U6822 (N_6822,N_1823,N_672);
and U6823 (N_6823,N_4772,N_2353);
nand U6824 (N_6824,N_4866,N_2208);
or U6825 (N_6825,N_4100,N_914);
nor U6826 (N_6826,N_3239,N_3248);
or U6827 (N_6827,N_964,N_2569);
and U6828 (N_6828,N_4862,N_3053);
nor U6829 (N_6829,N_2061,N_4601);
and U6830 (N_6830,N_1054,N_3356);
or U6831 (N_6831,N_335,N_4784);
nor U6832 (N_6832,N_1647,N_1256);
nor U6833 (N_6833,N_3977,N_4319);
or U6834 (N_6834,N_593,N_3552);
nor U6835 (N_6835,N_2964,N_3206);
and U6836 (N_6836,N_4289,N_2763);
nor U6837 (N_6837,N_1027,N_4780);
or U6838 (N_6838,N_1649,N_307);
and U6839 (N_6839,N_4854,N_3846);
or U6840 (N_6840,N_779,N_1110);
or U6841 (N_6841,N_3422,N_1754);
and U6842 (N_6842,N_2202,N_3182);
nor U6843 (N_6843,N_2311,N_2138);
or U6844 (N_6844,N_878,N_4022);
nand U6845 (N_6845,N_733,N_355);
and U6846 (N_6846,N_2468,N_1376);
nor U6847 (N_6847,N_201,N_1719);
or U6848 (N_6848,N_4743,N_210);
or U6849 (N_6849,N_4192,N_4370);
nor U6850 (N_6850,N_148,N_395);
nand U6851 (N_6851,N_3244,N_3701);
nand U6852 (N_6852,N_2858,N_693);
nand U6853 (N_6853,N_1471,N_893);
and U6854 (N_6854,N_4096,N_2844);
nand U6855 (N_6855,N_3989,N_2469);
or U6856 (N_6856,N_3441,N_2039);
nor U6857 (N_6857,N_4353,N_2599);
nor U6858 (N_6858,N_3532,N_1592);
or U6859 (N_6859,N_2119,N_2617);
nand U6860 (N_6860,N_2936,N_1181);
and U6861 (N_6861,N_4901,N_1918);
nor U6862 (N_6862,N_3378,N_2372);
nor U6863 (N_6863,N_4773,N_50);
and U6864 (N_6864,N_3186,N_793);
or U6865 (N_6865,N_2749,N_3014);
and U6866 (N_6866,N_1427,N_342);
or U6867 (N_6867,N_4864,N_2909);
and U6868 (N_6868,N_2704,N_3996);
and U6869 (N_6869,N_3516,N_2031);
nand U6870 (N_6870,N_1477,N_4299);
nand U6871 (N_6871,N_1583,N_477);
nand U6872 (N_6872,N_244,N_4858);
and U6873 (N_6873,N_2541,N_4269);
or U6874 (N_6874,N_4961,N_2575);
and U6875 (N_6875,N_1267,N_1219);
nand U6876 (N_6876,N_653,N_4298);
nor U6877 (N_6877,N_909,N_1391);
nand U6878 (N_6878,N_522,N_4157);
and U6879 (N_6879,N_375,N_1602);
nor U6880 (N_6880,N_2103,N_3979);
or U6881 (N_6881,N_804,N_944);
nand U6882 (N_6882,N_4637,N_1830);
or U6883 (N_6883,N_2827,N_2322);
or U6884 (N_6884,N_4266,N_3257);
nand U6885 (N_6885,N_3573,N_3028);
or U6886 (N_6886,N_3559,N_4188);
and U6887 (N_6887,N_4047,N_4894);
or U6888 (N_6888,N_3527,N_3838);
and U6889 (N_6889,N_3168,N_1146);
and U6890 (N_6890,N_3249,N_213);
xor U6891 (N_6891,N_4303,N_1237);
and U6892 (N_6892,N_2623,N_2226);
nor U6893 (N_6893,N_3795,N_3634);
and U6894 (N_6894,N_4774,N_541);
nand U6895 (N_6895,N_344,N_2552);
nand U6896 (N_6896,N_3680,N_3648);
or U6897 (N_6897,N_3294,N_3369);
nand U6898 (N_6898,N_75,N_2500);
nor U6899 (N_6899,N_2578,N_2245);
and U6900 (N_6900,N_3899,N_4721);
nor U6901 (N_6901,N_2733,N_675);
nor U6902 (N_6902,N_442,N_4333);
and U6903 (N_6903,N_3635,N_2686);
and U6904 (N_6904,N_3671,N_2924);
nand U6905 (N_6905,N_3618,N_300);
nand U6906 (N_6906,N_169,N_48);
nor U6907 (N_6907,N_2164,N_1257);
nor U6908 (N_6908,N_1727,N_346);
and U6909 (N_6909,N_783,N_1563);
or U6910 (N_6910,N_2213,N_1803);
nand U6911 (N_6911,N_2657,N_351);
nor U6912 (N_6912,N_113,N_4233);
nand U6913 (N_6913,N_2049,N_3242);
or U6914 (N_6914,N_2513,N_2636);
nand U6915 (N_6915,N_4695,N_1962);
or U6916 (N_6916,N_2562,N_1601);
nor U6917 (N_6917,N_2329,N_2564);
or U6918 (N_6918,N_1434,N_2076);
nor U6919 (N_6919,N_4294,N_858);
and U6920 (N_6920,N_2984,N_3283);
and U6921 (N_6921,N_4131,N_460);
or U6922 (N_6922,N_1071,N_1454);
nor U6923 (N_6923,N_4850,N_747);
and U6924 (N_6924,N_988,N_150);
xor U6925 (N_6925,N_4041,N_592);
and U6926 (N_6926,N_4379,N_176);
and U6927 (N_6927,N_1187,N_411);
nor U6928 (N_6928,N_3625,N_801);
nand U6929 (N_6929,N_3107,N_2094);
or U6930 (N_6930,N_3483,N_4076);
and U6931 (N_6931,N_1022,N_23);
or U6932 (N_6932,N_3360,N_2775);
and U6933 (N_6933,N_3444,N_1673);
and U6934 (N_6934,N_2981,N_1084);
and U6935 (N_6935,N_2650,N_4595);
or U6936 (N_6936,N_2934,N_1228);
or U6937 (N_6937,N_4314,N_4916);
and U6938 (N_6938,N_4825,N_466);
nand U6939 (N_6939,N_3530,N_1401);
nor U6940 (N_6940,N_2403,N_381);
nand U6941 (N_6941,N_2190,N_86);
or U6942 (N_6942,N_3129,N_797);
nand U6943 (N_6943,N_1761,N_1851);
nand U6944 (N_6944,N_2730,N_4315);
or U6945 (N_6945,N_3308,N_2259);
nor U6946 (N_6946,N_727,N_4980);
nand U6947 (N_6947,N_4546,N_4077);
or U6948 (N_6948,N_2519,N_3179);
nor U6949 (N_6949,N_2252,N_3288);
and U6950 (N_6950,N_3877,N_4824);
or U6951 (N_6951,N_3307,N_3543);
nor U6952 (N_6952,N_764,N_1818);
and U6953 (N_6953,N_1097,N_1731);
or U6954 (N_6954,N_3459,N_3273);
xnor U6955 (N_6955,N_3952,N_3460);
nor U6956 (N_6956,N_3181,N_2189);
and U6957 (N_6957,N_1135,N_1948);
or U6958 (N_6958,N_368,N_4340);
nor U6959 (N_6959,N_1338,N_4097);
nor U6960 (N_6960,N_982,N_1615);
nor U6961 (N_6961,N_3437,N_4248);
or U6962 (N_6962,N_1581,N_3768);
nand U6963 (N_6963,N_1025,N_2803);
nand U6964 (N_6964,N_4015,N_4561);
nand U6965 (N_6965,N_2279,N_3772);
nand U6966 (N_6966,N_4415,N_3265);
nor U6967 (N_6967,N_3830,N_4566);
or U6968 (N_6968,N_908,N_352);
nor U6969 (N_6969,N_4547,N_1258);
and U6970 (N_6970,N_321,N_88);
and U6971 (N_6971,N_2072,N_3401);
or U6972 (N_6972,N_3526,N_1077);
and U6973 (N_6973,N_1013,N_2131);
nor U6974 (N_6974,N_935,N_996);
nor U6975 (N_6975,N_3872,N_2584);
or U6976 (N_6976,N_2831,N_305);
nor U6977 (N_6977,N_2176,N_4371);
or U6978 (N_6978,N_480,N_556);
nor U6979 (N_6979,N_1248,N_2089);
and U6980 (N_6980,N_4575,N_3071);
and U6981 (N_6981,N_30,N_4835);
and U6982 (N_6982,N_1643,N_533);
or U6983 (N_6983,N_4338,N_2876);
or U6984 (N_6984,N_1750,N_4120);
nand U6985 (N_6985,N_2985,N_4697);
and U6986 (N_6986,N_3451,N_1777);
nand U6987 (N_6987,N_253,N_3099);
nor U6988 (N_6988,N_4405,N_1686);
or U6989 (N_6989,N_2420,N_2628);
nor U6990 (N_6990,N_3418,N_4534);
and U6991 (N_6991,N_6,N_3505);
nor U6992 (N_6992,N_3046,N_2151);
nor U6993 (N_6993,N_2707,N_1997);
nor U6994 (N_6994,N_1947,N_1305);
or U6995 (N_6995,N_238,N_4609);
nand U6996 (N_6996,N_3166,N_1622);
and U6997 (N_6997,N_4262,N_3518);
nor U6998 (N_6998,N_4075,N_274);
and U6999 (N_6999,N_1937,N_4326);
nor U7000 (N_7000,N_4387,N_1855);
or U7001 (N_7001,N_4790,N_1812);
nand U7002 (N_7002,N_1418,N_4831);
nand U7003 (N_7003,N_4680,N_1553);
or U7004 (N_7004,N_3742,N_1400);
or U7005 (N_7005,N_1796,N_1961);
nand U7006 (N_7006,N_3586,N_2696);
and U7007 (N_7007,N_3776,N_2362);
nor U7008 (N_7008,N_11,N_1939);
xor U7009 (N_7009,N_4455,N_4479);
or U7010 (N_7010,N_369,N_2706);
and U7011 (N_7011,N_3240,N_3939);
xor U7012 (N_7012,N_3500,N_4531);
and U7013 (N_7013,N_4826,N_650);
nor U7014 (N_7014,N_54,N_3332);
nand U7015 (N_7015,N_3204,N_3377);
and U7016 (N_7016,N_4470,N_1582);
nor U7017 (N_7017,N_3871,N_1960);
nand U7018 (N_7018,N_4811,N_4058);
nor U7019 (N_7019,N_507,N_3824);
or U7020 (N_7020,N_3305,N_3643);
or U7021 (N_7021,N_1413,N_3173);
xnor U7022 (N_7022,N_1983,N_2220);
nor U7023 (N_7023,N_1243,N_1069);
nor U7024 (N_7024,N_2897,N_543);
and U7025 (N_7025,N_2621,N_4717);
and U7026 (N_7026,N_3812,N_392);
nand U7027 (N_7027,N_1912,N_1021);
xor U7028 (N_7028,N_3049,N_1396);
or U7029 (N_7029,N_3954,N_327);
and U7030 (N_7030,N_710,N_2140);
or U7031 (N_7031,N_436,N_364);
nand U7032 (N_7032,N_4474,N_3139);
xnor U7033 (N_7033,N_4419,N_2937);
and U7034 (N_7034,N_4471,N_3678);
or U7035 (N_7035,N_508,N_4293);
nor U7036 (N_7036,N_4234,N_2629);
or U7037 (N_7037,N_4542,N_4739);
nand U7038 (N_7038,N_2376,N_4229);
or U7039 (N_7039,N_4863,N_741);
and U7040 (N_7040,N_940,N_358);
nor U7041 (N_7041,N_3900,N_3550);
nand U7042 (N_7042,N_3142,N_3266);
and U7043 (N_7043,N_2343,N_1111);
nor U7044 (N_7044,N_2503,N_1648);
and U7045 (N_7045,N_2110,N_4955);
or U7046 (N_7046,N_1641,N_4297);
nand U7047 (N_7047,N_785,N_2440);
and U7048 (N_7048,N_2741,N_270);
xnor U7049 (N_7049,N_363,N_3673);
nand U7050 (N_7050,N_2373,N_841);
nor U7051 (N_7051,N_2891,N_4810);
nand U7052 (N_7052,N_568,N_199);
and U7053 (N_7053,N_3235,N_4849);
nor U7054 (N_7054,N_2709,N_379);
nor U7055 (N_7055,N_4213,N_1151);
and U7056 (N_7056,N_2129,N_4237);
and U7057 (N_7057,N_855,N_2878);
and U7058 (N_7058,N_193,N_3745);
and U7059 (N_7059,N_4684,N_943);
xor U7060 (N_7060,N_2008,N_528);
or U7061 (N_7061,N_1537,N_3324);
nand U7062 (N_7062,N_1107,N_4518);
and U7063 (N_7063,N_1222,N_3801);
and U7064 (N_7064,N_1976,N_382);
and U7065 (N_7065,N_1974,N_1921);
xor U7066 (N_7066,N_2231,N_2746);
and U7067 (N_7067,N_882,N_2399);
and U7068 (N_7068,N_2205,N_3408);
or U7069 (N_7069,N_1586,N_1470);
nor U7070 (N_7070,N_4274,N_3075);
nand U7071 (N_7071,N_3453,N_4738);
nor U7072 (N_7072,N_678,N_4498);
or U7073 (N_7073,N_398,N_2570);
or U7074 (N_7074,N_3382,N_1337);
or U7075 (N_7075,N_4478,N_4883);
nand U7076 (N_7076,N_587,N_1540);
nand U7077 (N_7077,N_4069,N_4488);
nand U7078 (N_7078,N_2398,N_306);
nand U7079 (N_7079,N_1729,N_4343);
or U7080 (N_7080,N_3962,N_3383);
and U7081 (N_7081,N_1311,N_509);
xnor U7082 (N_7082,N_1308,N_3262);
nand U7083 (N_7083,N_3819,N_3361);
or U7084 (N_7084,N_3836,N_43);
or U7085 (N_7085,N_3301,N_603);
and U7086 (N_7086,N_2742,N_2533);
and U7087 (N_7087,N_3833,N_147);
and U7088 (N_7088,N_1378,N_990);
or U7089 (N_7089,N_3683,N_4708);
nand U7090 (N_7090,N_3429,N_354);
and U7091 (N_7091,N_2899,N_521);
or U7092 (N_7092,N_1631,N_4642);
nor U7093 (N_7093,N_2801,N_4803);
nand U7094 (N_7094,N_1760,N_367);
nor U7095 (N_7095,N_1891,N_1096);
nand U7096 (N_7096,N_4532,N_500);
nand U7097 (N_7097,N_835,N_2673);
or U7098 (N_7098,N_3471,N_4197);
or U7099 (N_7099,N_2363,N_235);
and U7100 (N_7100,N_3822,N_3461);
nand U7101 (N_7101,N_2027,N_1845);
or U7102 (N_7102,N_2821,N_1095);
and U7103 (N_7103,N_1162,N_1381);
nor U7104 (N_7104,N_2561,N_1872);
and U7105 (N_7105,N_465,N_3170);
nand U7106 (N_7106,N_1560,N_4394);
nand U7107 (N_7107,N_1737,N_2544);
nand U7108 (N_7108,N_151,N_1981);
and U7109 (N_7109,N_3803,N_4190);
nor U7110 (N_7110,N_2438,N_3051);
and U7111 (N_7111,N_4490,N_141);
nor U7112 (N_7112,N_126,N_2656);
or U7113 (N_7113,N_116,N_4943);
and U7114 (N_7114,N_134,N_4123);
nand U7115 (N_7115,N_3984,N_2682);
or U7116 (N_7116,N_21,N_3141);
nand U7117 (N_7117,N_1487,N_3475);
nor U7118 (N_7118,N_4752,N_2491);
nor U7119 (N_7119,N_1041,N_4954);
or U7120 (N_7120,N_1817,N_333);
nor U7121 (N_7121,N_4676,N_2906);
and U7122 (N_7122,N_4085,N_3572);
or U7123 (N_7123,N_2479,N_2846);
nor U7124 (N_7124,N_1526,N_2856);
and U7125 (N_7125,N_4062,N_4947);
nor U7126 (N_7126,N_2088,N_1594);
nor U7127 (N_7127,N_3972,N_840);
or U7128 (N_7128,N_3779,N_2439);
and U7129 (N_7129,N_4785,N_1861);
or U7130 (N_7130,N_4952,N_3980);
nor U7131 (N_7131,N_3514,N_4627);
nand U7132 (N_7132,N_860,N_4574);
nor U7133 (N_7133,N_4799,N_4440);
or U7134 (N_7134,N_1612,N_2452);
or U7135 (N_7135,N_4276,N_2478);
nand U7136 (N_7136,N_2874,N_2282);
nor U7137 (N_7137,N_891,N_4844);
nand U7138 (N_7138,N_3371,N_1703);
nor U7139 (N_7139,N_2262,N_2067);
nand U7140 (N_7140,N_437,N_4249);
xnor U7141 (N_7141,N_4184,N_380);
nand U7142 (N_7142,N_1158,N_3119);
and U7143 (N_7143,N_316,N_4306);
or U7144 (N_7144,N_4103,N_4110);
or U7145 (N_7145,N_2610,N_1482);
nand U7146 (N_7146,N_3245,N_4851);
nor U7147 (N_7147,N_3187,N_3810);
xor U7148 (N_7148,N_3477,N_1344);
and U7149 (N_7149,N_4544,N_2943);
xor U7150 (N_7150,N_1119,N_3131);
or U7151 (N_7151,N_2509,N_549);
and U7152 (N_7152,N_4584,N_1411);
nor U7153 (N_7153,N_3809,N_59);
nor U7154 (N_7154,N_1693,N_2069);
nand U7155 (N_7155,N_3562,N_3195);
nand U7156 (N_7156,N_518,N_214);
or U7157 (N_7157,N_917,N_1220);
xnor U7158 (N_7158,N_2549,N_365);
nand U7159 (N_7159,N_4204,N_3928);
or U7160 (N_7160,N_1885,N_3388);
nor U7161 (N_7161,N_3127,N_2848);
xor U7162 (N_7162,N_1288,N_2470);
nand U7163 (N_7163,N_221,N_3941);
nor U7164 (N_7164,N_821,N_1511);
or U7165 (N_7165,N_3574,N_3990);
or U7166 (N_7166,N_1085,N_217);
or U7167 (N_7167,N_4718,N_3717);
and U7168 (N_7168,N_478,N_345);
and U7169 (N_7169,N_4660,N_2523);
and U7170 (N_7170,N_2266,N_2917);
nand U7171 (N_7171,N_2348,N_4927);
nand U7172 (N_7172,N_2232,N_71);
or U7173 (N_7173,N_4043,N_2619);
nor U7174 (N_7174,N_3409,N_4009);
nand U7175 (N_7175,N_1180,N_2980);
and U7176 (N_7176,N_2959,N_3277);
nor U7177 (N_7177,N_1028,N_3405);
and U7178 (N_7178,N_4936,N_3109);
or U7179 (N_7179,N_135,N_1875);
xnor U7180 (N_7180,N_660,N_2676);
nand U7181 (N_7181,N_3095,N_645);
and U7182 (N_7182,N_3723,N_4422);
and U7183 (N_7183,N_2397,N_1259);
nand U7184 (N_7184,N_1689,N_670);
nand U7185 (N_7185,N_2814,N_422);
nor U7186 (N_7186,N_4881,N_2596);
nand U7187 (N_7187,N_3343,N_4624);
and U7188 (N_7188,N_4557,N_1987);
or U7189 (N_7189,N_4328,N_1292);
xor U7190 (N_7190,N_3706,N_2181);
nand U7191 (N_7191,N_1261,N_68);
and U7192 (N_7192,N_389,N_2333);
nor U7193 (N_7193,N_2669,N_3960);
or U7194 (N_7194,N_655,N_2986);
and U7195 (N_7195,N_1580,N_4312);
xor U7196 (N_7196,N_4834,N_2122);
nand U7197 (N_7197,N_2641,N_889);
nor U7198 (N_7198,N_3533,N_3598);
and U7199 (N_7199,N_2958,N_639);
and U7200 (N_7200,N_1711,N_2083);
nand U7201 (N_7201,N_1116,N_2889);
or U7202 (N_7202,N_2411,N_3232);
or U7203 (N_7203,N_2024,N_2217);
and U7204 (N_7204,N_3702,N_1485);
nor U7205 (N_7205,N_662,N_3961);
nor U7206 (N_7206,N_3610,N_3700);
or U7207 (N_7207,N_160,N_1078);
and U7208 (N_7208,N_3727,N_716);
or U7209 (N_7209,N_3763,N_4505);
nand U7210 (N_7210,N_4714,N_2127);
and U7211 (N_7211,N_3856,N_216);
nand U7212 (N_7212,N_3644,N_536);
and U7213 (N_7213,N_12,N_2249);
nor U7214 (N_7214,N_308,N_1827);
nand U7215 (N_7215,N_1880,N_1201);
nor U7216 (N_7216,N_3726,N_2618);
or U7217 (N_7217,N_2737,N_2517);
nor U7218 (N_7218,N_2851,N_4207);
nor U7219 (N_7219,N_2952,N_4764);
and U7220 (N_7220,N_2193,N_1973);
nand U7221 (N_7221,N_4552,N_4599);
nand U7222 (N_7222,N_4643,N_997);
nand U7223 (N_7223,N_4124,N_1490);
nor U7224 (N_7224,N_502,N_3185);
or U7225 (N_7225,N_978,N_2884);
xor U7226 (N_7226,N_2390,N_4533);
nand U7227 (N_7227,N_2652,N_3508);
nand U7228 (N_7228,N_3538,N_2084);
nand U7229 (N_7229,N_3501,N_446);
or U7230 (N_7230,N_673,N_4048);
or U7231 (N_7231,N_325,N_4626);
and U7232 (N_7232,N_1809,N_3087);
nor U7233 (N_7233,N_749,N_296);
and U7234 (N_7234,N_2459,N_4443);
or U7235 (N_7235,N_262,N_4576);
and U7236 (N_7236,N_2922,N_1326);
nor U7237 (N_7237,N_4558,N_1881);
and U7238 (N_7238,N_3751,N_4675);
nand U7239 (N_7239,N_3274,N_2070);
or U7240 (N_7240,N_604,N_4132);
nor U7241 (N_7241,N_374,N_2698);
or U7242 (N_7242,N_2108,N_2941);
nand U7243 (N_7243,N_3806,N_4960);
and U7244 (N_7244,N_3033,N_1545);
nor U7245 (N_7245,N_17,N_4450);
or U7246 (N_7246,N_3821,N_0);
nand U7247 (N_7247,N_767,N_4005);
nor U7248 (N_7248,N_3466,N_2444);
nand U7249 (N_7249,N_1164,N_4727);
nor U7250 (N_7250,N_2450,N_4116);
nor U7251 (N_7251,N_1900,N_4409);
nor U7252 (N_7252,N_1620,N_4583);
nor U7253 (N_7253,N_532,N_919);
and U7254 (N_7254,N_4906,N_3808);
or U7255 (N_7255,N_2458,N_3151);
or U7256 (N_7256,N_1234,N_4222);
nand U7257 (N_7257,N_2560,N_3036);
nor U7258 (N_7258,N_669,N_1318);
or U7259 (N_7259,N_4525,N_2925);
nand U7260 (N_7260,N_1061,N_2752);
nor U7261 (N_7261,N_1282,N_4665);
and U7262 (N_7262,N_1426,N_1176);
nand U7263 (N_7263,N_4663,N_4178);
or U7264 (N_7264,N_4119,N_1725);
or U7265 (N_7265,N_1301,N_1343);
nor U7266 (N_7266,N_920,N_3649);
nand U7267 (N_7267,N_4641,N_1531);
and U7268 (N_7268,N_2961,N_2100);
or U7269 (N_7269,N_2931,N_4817);
or U7270 (N_7270,N_3440,N_3784);
and U7271 (N_7271,N_2281,N_4932);
nor U7272 (N_7272,N_1864,N_263);
and U7273 (N_7273,N_3631,N_757);
xnor U7274 (N_7274,N_3750,N_413);
nand U7275 (N_7275,N_361,N_2211);
nand U7276 (N_7276,N_1373,N_2003);
nand U7277 (N_7277,N_4704,N_195);
or U7278 (N_7278,N_4529,N_3448);
and U7279 (N_7279,N_728,N_530);
nor U7280 (N_7280,N_644,N_4931);
or U7281 (N_7281,N_3594,N_3024);
nand U7282 (N_7282,N_3953,N_2476);
nand U7283 (N_7283,N_1723,N_3740);
xor U7284 (N_7284,N_3786,N_3455);
nor U7285 (N_7285,N_973,N_3255);
nor U7286 (N_7286,N_2699,N_4726);
or U7287 (N_7287,N_1752,N_4281);
or U7288 (N_7288,N_4939,N_4871);
and U7289 (N_7289,N_3234,N_4138);
or U7290 (N_7290,N_4404,N_3261);
or U7291 (N_7291,N_1709,N_1143);
and U7292 (N_7292,N_4555,N_4693);
nor U7293 (N_7293,N_651,N_2389);
or U7294 (N_7294,N_1776,N_3379);
nor U7295 (N_7295,N_295,N_2378);
nor U7296 (N_7296,N_2337,N_1023);
nor U7297 (N_7297,N_1216,N_1524);
or U7298 (N_7298,N_2038,N_915);
nand U7299 (N_7299,N_688,N_985);
or U7300 (N_7300,N_2427,N_2312);
or U7301 (N_7301,N_2174,N_1334);
or U7302 (N_7302,N_3023,N_4733);
nand U7303 (N_7303,N_4142,N_431);
nor U7304 (N_7304,N_3911,N_1074);
or U7305 (N_7305,N_2320,N_4346);
nand U7306 (N_7306,N_2866,N_1065);
and U7307 (N_7307,N_1374,N_1635);
xor U7308 (N_7308,N_179,N_4198);
or U7309 (N_7309,N_1728,N_1322);
or U7310 (N_7310,N_1789,N_2369);
or U7311 (N_7311,N_46,N_2554);
xor U7312 (N_7312,N_856,N_3464);
nand U7313 (N_7313,N_348,N_759);
or U7314 (N_7314,N_3017,N_1743);
nor U7315 (N_7315,N_3845,N_2436);
nand U7316 (N_7316,N_2532,N_2018);
nor U7317 (N_7317,N_4321,N_1274);
and U7318 (N_7318,N_286,N_1839);
and U7319 (N_7319,N_4155,N_1853);
or U7320 (N_7320,N_1772,N_2242);
nand U7321 (N_7321,N_2818,N_2790);
and U7322 (N_7322,N_1831,N_4079);
or U7323 (N_7323,N_4143,N_4067);
or U7324 (N_7324,N_1329,N_1701);
nor U7325 (N_7325,N_4250,N_4795);
and U7326 (N_7326,N_1251,N_3399);
and U7327 (N_7327,N_4373,N_4499);
nor U7328 (N_7328,N_3888,N_1087);
nand U7329 (N_7329,N_3007,N_4651);
or U7330 (N_7330,N_896,N_223);
nor U7331 (N_7331,N_31,N_1399);
nand U7332 (N_7332,N_192,N_1226);
nand U7333 (N_7333,N_3481,N_2182);
or U7334 (N_7334,N_815,N_664);
or U7335 (N_7335,N_1561,N_2493);
nor U7336 (N_7336,N_1559,N_2482);
nor U7337 (N_7337,N_2112,N_2867);
nand U7338 (N_7338,N_3770,N_2510);
and U7339 (N_7339,N_2695,N_1163);
nor U7340 (N_7340,N_417,N_3474);
or U7341 (N_7341,N_3826,N_3504);
or U7342 (N_7342,N_2297,N_4271);
and U7343 (N_7343,N_4324,N_2106);
and U7344 (N_7344,N_4769,N_4400);
nor U7345 (N_7345,N_3384,N_3123);
nor U7346 (N_7346,N_1060,N_4242);
and U7347 (N_7347,N_525,N_3341);
nand U7348 (N_7348,N_3155,N_3147);
and U7349 (N_7349,N_3592,N_4230);
and U7350 (N_7350,N_3258,N_2234);
nand U7351 (N_7351,N_635,N_4759);
or U7352 (N_7352,N_2044,N_1079);
or U7353 (N_7353,N_3364,N_2166);
xor U7354 (N_7354,N_3556,N_2071);
and U7355 (N_7355,N_4728,N_3224);
and U7356 (N_7356,N_956,N_2576);
and U7357 (N_7357,N_1075,N_1638);
or U7358 (N_7358,N_1584,N_849);
or U7359 (N_7359,N_2759,N_1771);
nand U7360 (N_7360,N_3213,N_3407);
nand U7361 (N_7361,N_2594,N_1860);
nand U7362 (N_7362,N_4265,N_1644);
and U7363 (N_7363,N_3112,N_730);
or U7364 (N_7364,N_2441,N_1369);
and U7365 (N_7365,N_2488,N_1215);
or U7366 (N_7366,N_926,N_4616);
nand U7367 (N_7367,N_3042,N_3349);
nor U7368 (N_7368,N_901,N_1214);
or U7369 (N_7369,N_1527,N_2942);
nand U7370 (N_7370,N_4368,N_2568);
or U7371 (N_7371,N_2918,N_58);
and U7372 (N_7372,N_3298,N_3006);
xnor U7373 (N_7373,N_3875,N_1191);
xnor U7374 (N_7374,N_1002,N_534);
nand U7375 (N_7375,N_3760,N_1276);
and U7376 (N_7376,N_2545,N_2356);
nor U7377 (N_7377,N_4523,N_1492);
nand U7378 (N_7378,N_3995,N_3991);
or U7379 (N_7379,N_4968,N_4972);
nor U7380 (N_7380,N_2668,N_2105);
xnor U7381 (N_7381,N_1706,N_814);
xor U7382 (N_7382,N_2724,N_2435);
nand U7383 (N_7383,N_3192,N_467);
or U7384 (N_7384,N_809,N_4454);
and U7385 (N_7385,N_3359,N_4171);
nand U7386 (N_7386,N_2526,N_73);
nor U7387 (N_7387,N_989,N_3764);
nor U7388 (N_7388,N_3611,N_140);
nor U7389 (N_7389,N_3884,N_3325);
and U7390 (N_7390,N_4214,N_1423);
and U7391 (N_7391,N_2325,N_2802);
nand U7392 (N_7392,N_4904,N_1634);
nand U7393 (N_7393,N_324,N_4354);
nand U7394 (N_7394,N_1088,N_304);
nor U7395 (N_7395,N_4042,N_3617);
or U7396 (N_7396,N_1500,N_1093);
and U7397 (N_7397,N_283,N_939);
and U7398 (N_7398,N_3287,N_2136);
nor U7399 (N_7399,N_3553,N_102);
or U7400 (N_7400,N_4567,N_4938);
nor U7401 (N_7401,N_977,N_3496);
or U7402 (N_7402,N_3674,N_390);
or U7403 (N_7403,N_954,N_4446);
or U7404 (N_7404,N_4011,N_4055);
or U7405 (N_7405,N_4208,N_1712);
or U7406 (N_7406,N_4821,N_3290);
nand U7407 (N_7407,N_2625,N_924);
or U7408 (N_7408,N_2388,N_4291);
nor U7409 (N_7409,N_1125,N_2153);
nor U7410 (N_7410,N_842,N_2720);
or U7411 (N_7411,N_3063,N_1072);
nand U7412 (N_7412,N_4322,N_3748);
or U7413 (N_7413,N_986,N_3755);
nor U7414 (N_7414,N_3094,N_2793);
and U7415 (N_7415,N_1341,N_1159);
nor U7416 (N_7416,N_3158,N_1348);
or U7417 (N_7417,N_2608,N_1977);
and U7418 (N_7418,N_36,N_2051);
or U7419 (N_7419,N_3091,N_2735);
nor U7420 (N_7420,N_4703,N_4300);
or U7421 (N_7421,N_3005,N_414);
and U7422 (N_7422,N_2536,N_1001);
and U7423 (N_7423,N_3951,N_4118);
nor U7424 (N_7424,N_912,N_183);
nand U7425 (N_7425,N_2558,N_2525);
or U7426 (N_7426,N_2377,N_1034);
or U7427 (N_7427,N_1342,N_3811);
nand U7428 (N_7428,N_164,N_2666);
and U7429 (N_7429,N_4701,N_438);
xor U7430 (N_7430,N_3563,N_617);
nand U7431 (N_7431,N_1514,N_72);
and U7432 (N_7432,N_813,N_1285);
or U7433 (N_7433,N_631,N_1441);
or U7434 (N_7434,N_4391,N_1070);
nand U7435 (N_7435,N_287,N_3919);
and U7436 (N_7436,N_299,N_3602);
and U7437 (N_7437,N_4867,N_3882);
nor U7438 (N_7438,N_861,N_1915);
nor U7439 (N_7439,N_1730,N_2973);
or U7440 (N_7440,N_303,N_696);
and U7441 (N_7441,N_4791,N_3679);
nor U7442 (N_7442,N_2708,N_1759);
and U7443 (N_7443,N_4187,N_4031);
or U7444 (N_7444,N_1012,N_24);
nor U7445 (N_7445,N_3038,N_3176);
or U7446 (N_7446,N_911,N_4352);
nor U7447 (N_7447,N_3981,N_167);
nor U7448 (N_7448,N_1059,N_1585);
nand U7449 (N_7449,N_2997,N_2810);
nor U7450 (N_7450,N_787,N_2063);
nor U7451 (N_7451,N_3076,N_2565);
nand U7452 (N_7452,N_752,N_566);
xnor U7453 (N_7453,N_4451,N_1287);
and U7454 (N_7454,N_1414,N_1655);
or U7455 (N_7455,N_4408,N_470);
and U7456 (N_7456,N_1211,N_3835);
nand U7457 (N_7457,N_451,N_3616);
nor U7458 (N_7458,N_3615,N_347);
nor U7459 (N_7459,N_1457,N_4526);
and U7460 (N_7460,N_2822,N_4485);
nor U7461 (N_7461,N_2948,N_3449);
nor U7462 (N_7462,N_2143,N_2877);
nor U7463 (N_7463,N_2171,N_4359);
and U7464 (N_7464,N_3839,N_4061);
or U7465 (N_7465,N_3887,N_1137);
or U7466 (N_7466,N_1681,N_712);
or U7467 (N_7467,N_3116,N_2330);
nor U7468 (N_7468,N_4232,N_1039);
or U7469 (N_7469,N_1687,N_2218);
or U7470 (N_7470,N_3306,N_2269);
nor U7471 (N_7471,N_3769,N_4853);
nand U7472 (N_7472,N_4121,N_2239);
or U7473 (N_7473,N_4425,N_3110);
or U7474 (N_7474,N_1415,N_3849);
or U7475 (N_7475,N_4895,N_168);
or U7476 (N_7476,N_2728,N_3534);
nor U7477 (N_7477,N_1798,N_1979);
nor U7478 (N_7478,N_2338,N_4464);
nor U7479 (N_7479,N_2603,N_2235);
nand U7480 (N_7480,N_2210,N_4122);
or U7481 (N_7481,N_1554,N_3177);
nand U7482 (N_7482,N_4649,N_2498);
nand U7483 (N_7483,N_419,N_2863);
nand U7484 (N_7484,N_4449,N_1468);
or U7485 (N_7485,N_2342,N_3756);
and U7486 (N_7486,N_209,N_3406);
and U7487 (N_7487,N_400,N_2216);
nor U7488 (N_7488,N_3214,N_1185);
or U7489 (N_7489,N_3199,N_4202);
nor U7490 (N_7490,N_3148,N_3522);
or U7491 (N_7491,N_2734,N_2516);
nand U7492 (N_7492,N_1339,N_581);
and U7493 (N_7493,N_1826,N_3105);
nand U7494 (N_7494,N_1298,N_2461);
or U7495 (N_7495,N_2483,N_875);
nor U7496 (N_7496,N_739,N_2419);
nand U7497 (N_7497,N_1134,N_4897);
nor U7498 (N_7498,N_3061,N_37);
nand U7499 (N_7499,N_2785,N_1068);
and U7500 (N_7500,N_673,N_4070);
or U7501 (N_7501,N_437,N_1684);
or U7502 (N_7502,N_999,N_1363);
nand U7503 (N_7503,N_1453,N_1227);
xor U7504 (N_7504,N_10,N_1149);
or U7505 (N_7505,N_1006,N_4176);
xnor U7506 (N_7506,N_3476,N_124);
nand U7507 (N_7507,N_2670,N_1047);
and U7508 (N_7508,N_295,N_1164);
nand U7509 (N_7509,N_4507,N_2946);
nand U7510 (N_7510,N_1946,N_1901);
and U7511 (N_7511,N_2887,N_3949);
nor U7512 (N_7512,N_665,N_3631);
nor U7513 (N_7513,N_4505,N_2090);
nand U7514 (N_7514,N_408,N_1699);
and U7515 (N_7515,N_2728,N_373);
and U7516 (N_7516,N_3910,N_359);
or U7517 (N_7517,N_4651,N_3789);
or U7518 (N_7518,N_1893,N_3314);
and U7519 (N_7519,N_1466,N_740);
and U7520 (N_7520,N_3859,N_329);
nor U7521 (N_7521,N_148,N_1253);
or U7522 (N_7522,N_2552,N_4961);
or U7523 (N_7523,N_3769,N_3881);
or U7524 (N_7524,N_2850,N_4152);
nand U7525 (N_7525,N_89,N_4238);
nor U7526 (N_7526,N_4370,N_3704);
or U7527 (N_7527,N_3243,N_4524);
nand U7528 (N_7528,N_115,N_3210);
nor U7529 (N_7529,N_2493,N_1264);
nand U7530 (N_7530,N_304,N_4437);
nor U7531 (N_7531,N_979,N_3835);
and U7532 (N_7532,N_540,N_747);
nand U7533 (N_7533,N_1237,N_2446);
or U7534 (N_7534,N_1121,N_3685);
xnor U7535 (N_7535,N_1624,N_2101);
and U7536 (N_7536,N_4986,N_2089);
nor U7537 (N_7537,N_4681,N_4347);
nor U7538 (N_7538,N_971,N_4555);
and U7539 (N_7539,N_1122,N_1815);
xor U7540 (N_7540,N_1387,N_901);
nand U7541 (N_7541,N_681,N_4539);
xnor U7542 (N_7542,N_2280,N_232);
nand U7543 (N_7543,N_4729,N_707);
nor U7544 (N_7544,N_4823,N_2198);
xnor U7545 (N_7545,N_2673,N_2775);
nor U7546 (N_7546,N_271,N_2390);
nand U7547 (N_7547,N_1577,N_70);
and U7548 (N_7548,N_2981,N_616);
or U7549 (N_7549,N_2819,N_2163);
and U7550 (N_7550,N_4506,N_2007);
nor U7551 (N_7551,N_4093,N_3506);
nor U7552 (N_7552,N_2322,N_344);
nor U7553 (N_7553,N_2577,N_1535);
and U7554 (N_7554,N_1444,N_1906);
or U7555 (N_7555,N_3097,N_4591);
nand U7556 (N_7556,N_1765,N_3496);
or U7557 (N_7557,N_2960,N_1631);
nand U7558 (N_7558,N_828,N_100);
nor U7559 (N_7559,N_4146,N_358);
or U7560 (N_7560,N_92,N_2273);
nand U7561 (N_7561,N_4165,N_4328);
or U7562 (N_7562,N_1861,N_4866);
and U7563 (N_7563,N_2034,N_2100);
nor U7564 (N_7564,N_1063,N_4829);
and U7565 (N_7565,N_1841,N_1431);
and U7566 (N_7566,N_1858,N_1338);
nand U7567 (N_7567,N_1840,N_2931);
or U7568 (N_7568,N_3553,N_3246);
or U7569 (N_7569,N_253,N_4653);
nor U7570 (N_7570,N_3260,N_167);
nor U7571 (N_7571,N_2707,N_4539);
nand U7572 (N_7572,N_3235,N_2284);
nor U7573 (N_7573,N_1937,N_3583);
or U7574 (N_7574,N_1619,N_1229);
nor U7575 (N_7575,N_4887,N_2899);
nor U7576 (N_7576,N_2251,N_4847);
nor U7577 (N_7577,N_2397,N_1006);
and U7578 (N_7578,N_1346,N_827);
and U7579 (N_7579,N_2146,N_4969);
nor U7580 (N_7580,N_4180,N_43);
nor U7581 (N_7581,N_3393,N_4385);
or U7582 (N_7582,N_1592,N_775);
nand U7583 (N_7583,N_3936,N_1565);
nand U7584 (N_7584,N_827,N_2988);
and U7585 (N_7585,N_420,N_4804);
and U7586 (N_7586,N_3838,N_4574);
nand U7587 (N_7587,N_4126,N_3132);
nor U7588 (N_7588,N_4735,N_443);
and U7589 (N_7589,N_4507,N_4364);
and U7590 (N_7590,N_473,N_4060);
xnor U7591 (N_7591,N_3044,N_1348);
and U7592 (N_7592,N_3262,N_3098);
and U7593 (N_7593,N_1203,N_758);
nor U7594 (N_7594,N_3035,N_4754);
nand U7595 (N_7595,N_1918,N_3728);
or U7596 (N_7596,N_4559,N_2754);
or U7597 (N_7597,N_2891,N_2963);
nand U7598 (N_7598,N_4748,N_111);
and U7599 (N_7599,N_2337,N_3686);
and U7600 (N_7600,N_3346,N_3057);
nor U7601 (N_7601,N_2531,N_524);
nor U7602 (N_7602,N_4096,N_1484);
nand U7603 (N_7603,N_1580,N_418);
nand U7604 (N_7604,N_3130,N_1095);
nand U7605 (N_7605,N_4296,N_4842);
nor U7606 (N_7606,N_2311,N_4407);
and U7607 (N_7607,N_1550,N_4758);
nor U7608 (N_7608,N_4884,N_3942);
or U7609 (N_7609,N_519,N_2779);
or U7610 (N_7610,N_1028,N_4222);
and U7611 (N_7611,N_1264,N_1086);
nor U7612 (N_7612,N_53,N_793);
nand U7613 (N_7613,N_3006,N_3218);
and U7614 (N_7614,N_1521,N_3784);
or U7615 (N_7615,N_1070,N_4234);
nor U7616 (N_7616,N_109,N_1442);
nand U7617 (N_7617,N_3294,N_991);
xor U7618 (N_7618,N_4382,N_601);
nand U7619 (N_7619,N_4481,N_1007);
or U7620 (N_7620,N_4951,N_2703);
nor U7621 (N_7621,N_2162,N_3257);
nor U7622 (N_7622,N_432,N_235);
or U7623 (N_7623,N_4122,N_4303);
nand U7624 (N_7624,N_2471,N_1164);
nand U7625 (N_7625,N_706,N_2791);
nand U7626 (N_7626,N_1136,N_2663);
nand U7627 (N_7627,N_169,N_2857);
nand U7628 (N_7628,N_4786,N_3122);
and U7629 (N_7629,N_984,N_268);
nand U7630 (N_7630,N_4943,N_4428);
nor U7631 (N_7631,N_1010,N_1582);
and U7632 (N_7632,N_712,N_2562);
or U7633 (N_7633,N_4675,N_16);
nor U7634 (N_7634,N_4215,N_2723);
or U7635 (N_7635,N_267,N_4639);
and U7636 (N_7636,N_2851,N_3603);
or U7637 (N_7637,N_2424,N_1737);
nand U7638 (N_7638,N_2434,N_1388);
nor U7639 (N_7639,N_2971,N_1558);
and U7640 (N_7640,N_3159,N_1749);
or U7641 (N_7641,N_2857,N_3993);
or U7642 (N_7642,N_183,N_1845);
and U7643 (N_7643,N_3551,N_3105);
nand U7644 (N_7644,N_4575,N_954);
or U7645 (N_7645,N_135,N_1897);
or U7646 (N_7646,N_828,N_4707);
or U7647 (N_7647,N_4279,N_2699);
nand U7648 (N_7648,N_4323,N_4426);
nand U7649 (N_7649,N_566,N_4128);
nor U7650 (N_7650,N_4609,N_3934);
nor U7651 (N_7651,N_2595,N_2497);
or U7652 (N_7652,N_2597,N_3172);
nor U7653 (N_7653,N_1011,N_2002);
and U7654 (N_7654,N_2147,N_1358);
nor U7655 (N_7655,N_2243,N_1277);
or U7656 (N_7656,N_2561,N_4009);
or U7657 (N_7657,N_4976,N_1334);
nand U7658 (N_7658,N_2226,N_233);
or U7659 (N_7659,N_3264,N_328);
nand U7660 (N_7660,N_1815,N_3559);
or U7661 (N_7661,N_3657,N_601);
nor U7662 (N_7662,N_3154,N_4953);
or U7663 (N_7663,N_999,N_3975);
or U7664 (N_7664,N_152,N_2154);
or U7665 (N_7665,N_481,N_1838);
nand U7666 (N_7666,N_3082,N_2582);
and U7667 (N_7667,N_118,N_1516);
and U7668 (N_7668,N_4578,N_3552);
and U7669 (N_7669,N_3369,N_1236);
or U7670 (N_7670,N_3713,N_3606);
or U7671 (N_7671,N_407,N_952);
nand U7672 (N_7672,N_4584,N_1317);
or U7673 (N_7673,N_1314,N_4663);
nor U7674 (N_7674,N_3542,N_2904);
and U7675 (N_7675,N_65,N_2485);
and U7676 (N_7676,N_2685,N_2373);
or U7677 (N_7677,N_842,N_2618);
and U7678 (N_7678,N_478,N_2059);
nand U7679 (N_7679,N_4706,N_819);
nor U7680 (N_7680,N_3761,N_2093);
nor U7681 (N_7681,N_806,N_738);
or U7682 (N_7682,N_1574,N_3341);
xor U7683 (N_7683,N_1421,N_3089);
or U7684 (N_7684,N_4066,N_2188);
or U7685 (N_7685,N_1685,N_3423);
nand U7686 (N_7686,N_2830,N_64);
and U7687 (N_7687,N_4573,N_4000);
and U7688 (N_7688,N_4860,N_2523);
xor U7689 (N_7689,N_751,N_3931);
or U7690 (N_7690,N_2810,N_1585);
nor U7691 (N_7691,N_466,N_560);
nand U7692 (N_7692,N_4479,N_2948);
nand U7693 (N_7693,N_716,N_1530);
xnor U7694 (N_7694,N_2079,N_332);
and U7695 (N_7695,N_2361,N_31);
and U7696 (N_7696,N_4794,N_4672);
nor U7697 (N_7697,N_2562,N_2969);
nor U7698 (N_7698,N_3969,N_3745);
nor U7699 (N_7699,N_1433,N_342);
or U7700 (N_7700,N_1723,N_1434);
and U7701 (N_7701,N_335,N_3568);
nand U7702 (N_7702,N_3256,N_590);
nor U7703 (N_7703,N_4311,N_2746);
nor U7704 (N_7704,N_620,N_1567);
nor U7705 (N_7705,N_4563,N_1559);
and U7706 (N_7706,N_1067,N_160);
or U7707 (N_7707,N_4002,N_3119);
or U7708 (N_7708,N_551,N_4500);
nand U7709 (N_7709,N_1498,N_1736);
or U7710 (N_7710,N_534,N_1077);
nand U7711 (N_7711,N_4516,N_703);
or U7712 (N_7712,N_3913,N_3785);
nand U7713 (N_7713,N_3505,N_2756);
nand U7714 (N_7714,N_3499,N_3791);
or U7715 (N_7715,N_4710,N_1632);
nor U7716 (N_7716,N_1698,N_4965);
and U7717 (N_7717,N_1570,N_2055);
nor U7718 (N_7718,N_4196,N_1496);
nor U7719 (N_7719,N_4782,N_4024);
nand U7720 (N_7720,N_3015,N_4360);
and U7721 (N_7721,N_1686,N_2015);
nor U7722 (N_7722,N_3272,N_1083);
nand U7723 (N_7723,N_4328,N_3615);
nor U7724 (N_7724,N_3233,N_4616);
nor U7725 (N_7725,N_51,N_4798);
and U7726 (N_7726,N_3105,N_2676);
and U7727 (N_7727,N_2357,N_3276);
and U7728 (N_7728,N_1417,N_829);
and U7729 (N_7729,N_447,N_108);
nor U7730 (N_7730,N_4320,N_1029);
nand U7731 (N_7731,N_4565,N_1381);
nand U7732 (N_7732,N_2022,N_1124);
or U7733 (N_7733,N_2399,N_1354);
nor U7734 (N_7734,N_273,N_2406);
nor U7735 (N_7735,N_3379,N_3794);
or U7736 (N_7736,N_4609,N_2467);
nand U7737 (N_7737,N_747,N_2608);
nor U7738 (N_7738,N_227,N_3778);
and U7739 (N_7739,N_1787,N_615);
nor U7740 (N_7740,N_1098,N_792);
nor U7741 (N_7741,N_2729,N_3794);
nand U7742 (N_7742,N_3536,N_2522);
nand U7743 (N_7743,N_3488,N_3763);
nor U7744 (N_7744,N_3141,N_4760);
or U7745 (N_7745,N_3931,N_1828);
nor U7746 (N_7746,N_4648,N_824);
nor U7747 (N_7747,N_470,N_1133);
nand U7748 (N_7748,N_4608,N_2846);
nor U7749 (N_7749,N_2108,N_1862);
xnor U7750 (N_7750,N_823,N_4171);
and U7751 (N_7751,N_4024,N_4930);
nor U7752 (N_7752,N_2308,N_1767);
nor U7753 (N_7753,N_2990,N_2116);
and U7754 (N_7754,N_2108,N_2948);
nand U7755 (N_7755,N_2151,N_1819);
nand U7756 (N_7756,N_2790,N_1548);
and U7757 (N_7757,N_3705,N_792);
or U7758 (N_7758,N_2585,N_999);
and U7759 (N_7759,N_4383,N_4324);
and U7760 (N_7760,N_4617,N_470);
and U7761 (N_7761,N_3337,N_981);
nand U7762 (N_7762,N_3274,N_2552);
nand U7763 (N_7763,N_3727,N_1539);
and U7764 (N_7764,N_25,N_4118);
nor U7765 (N_7765,N_2987,N_611);
nand U7766 (N_7766,N_918,N_4765);
or U7767 (N_7767,N_3033,N_3328);
or U7768 (N_7768,N_4418,N_3584);
nand U7769 (N_7769,N_1281,N_4700);
or U7770 (N_7770,N_2515,N_3635);
or U7771 (N_7771,N_1326,N_4788);
or U7772 (N_7772,N_1541,N_4528);
nand U7773 (N_7773,N_1792,N_2155);
xnor U7774 (N_7774,N_3597,N_1677);
nand U7775 (N_7775,N_3436,N_4337);
nand U7776 (N_7776,N_2573,N_3730);
or U7777 (N_7777,N_1525,N_1340);
nor U7778 (N_7778,N_181,N_2477);
nand U7779 (N_7779,N_3197,N_4760);
or U7780 (N_7780,N_328,N_2325);
nor U7781 (N_7781,N_4039,N_3292);
and U7782 (N_7782,N_695,N_206);
or U7783 (N_7783,N_2895,N_3556);
and U7784 (N_7784,N_831,N_2722);
and U7785 (N_7785,N_2320,N_1554);
nor U7786 (N_7786,N_1551,N_1822);
nand U7787 (N_7787,N_2988,N_3172);
or U7788 (N_7788,N_693,N_4791);
and U7789 (N_7789,N_55,N_4970);
nand U7790 (N_7790,N_3489,N_4411);
nor U7791 (N_7791,N_2836,N_1633);
or U7792 (N_7792,N_3176,N_1210);
nand U7793 (N_7793,N_1036,N_694);
nor U7794 (N_7794,N_1494,N_2125);
nor U7795 (N_7795,N_3212,N_3874);
nand U7796 (N_7796,N_919,N_4048);
nor U7797 (N_7797,N_1746,N_1526);
nand U7798 (N_7798,N_2824,N_1422);
or U7799 (N_7799,N_534,N_2275);
nand U7800 (N_7800,N_1448,N_2768);
nor U7801 (N_7801,N_3839,N_1788);
or U7802 (N_7802,N_161,N_4222);
and U7803 (N_7803,N_1639,N_4566);
or U7804 (N_7804,N_2023,N_4464);
nand U7805 (N_7805,N_2951,N_3221);
and U7806 (N_7806,N_3411,N_838);
nor U7807 (N_7807,N_3587,N_149);
nand U7808 (N_7808,N_3758,N_2376);
and U7809 (N_7809,N_3210,N_3271);
nand U7810 (N_7810,N_4090,N_4915);
or U7811 (N_7811,N_2038,N_2659);
or U7812 (N_7812,N_3968,N_2552);
nor U7813 (N_7813,N_788,N_2268);
nor U7814 (N_7814,N_1654,N_3369);
or U7815 (N_7815,N_2204,N_4465);
nand U7816 (N_7816,N_1856,N_4706);
nand U7817 (N_7817,N_4650,N_3915);
and U7818 (N_7818,N_62,N_351);
and U7819 (N_7819,N_1959,N_3471);
or U7820 (N_7820,N_2906,N_4264);
nor U7821 (N_7821,N_4170,N_1319);
nor U7822 (N_7822,N_3000,N_4650);
nor U7823 (N_7823,N_3229,N_4455);
nand U7824 (N_7824,N_1400,N_732);
and U7825 (N_7825,N_1879,N_1213);
or U7826 (N_7826,N_4745,N_2727);
nand U7827 (N_7827,N_2796,N_896);
or U7828 (N_7828,N_2665,N_478);
nand U7829 (N_7829,N_2867,N_1621);
and U7830 (N_7830,N_205,N_3767);
nand U7831 (N_7831,N_1672,N_4676);
or U7832 (N_7832,N_1889,N_213);
nand U7833 (N_7833,N_1464,N_1484);
nand U7834 (N_7834,N_1464,N_709);
and U7835 (N_7835,N_3561,N_3402);
xor U7836 (N_7836,N_3846,N_3228);
nand U7837 (N_7837,N_448,N_4196);
nand U7838 (N_7838,N_485,N_2092);
or U7839 (N_7839,N_1220,N_4794);
and U7840 (N_7840,N_2927,N_3401);
nand U7841 (N_7841,N_636,N_249);
xor U7842 (N_7842,N_3603,N_2513);
and U7843 (N_7843,N_3211,N_1136);
and U7844 (N_7844,N_3276,N_3766);
or U7845 (N_7845,N_961,N_3703);
nor U7846 (N_7846,N_330,N_459);
or U7847 (N_7847,N_4119,N_4904);
and U7848 (N_7848,N_2950,N_3813);
nand U7849 (N_7849,N_3356,N_807);
nand U7850 (N_7850,N_552,N_3554);
and U7851 (N_7851,N_2542,N_2668);
and U7852 (N_7852,N_3620,N_4734);
nor U7853 (N_7853,N_797,N_2984);
and U7854 (N_7854,N_2003,N_598);
nand U7855 (N_7855,N_2110,N_4553);
and U7856 (N_7856,N_1965,N_4226);
nand U7857 (N_7857,N_3163,N_1140);
and U7858 (N_7858,N_643,N_2056);
nand U7859 (N_7859,N_2007,N_2901);
and U7860 (N_7860,N_388,N_534);
or U7861 (N_7861,N_2430,N_1746);
nor U7862 (N_7862,N_3123,N_1618);
and U7863 (N_7863,N_147,N_200);
and U7864 (N_7864,N_4373,N_4078);
nand U7865 (N_7865,N_4842,N_886);
and U7866 (N_7866,N_3588,N_1030);
nand U7867 (N_7867,N_3482,N_1965);
or U7868 (N_7868,N_2542,N_4388);
nor U7869 (N_7869,N_4575,N_1418);
nor U7870 (N_7870,N_266,N_464);
and U7871 (N_7871,N_3375,N_865);
and U7872 (N_7872,N_861,N_4650);
nand U7873 (N_7873,N_4400,N_1414);
nor U7874 (N_7874,N_4585,N_1719);
nor U7875 (N_7875,N_798,N_291);
or U7876 (N_7876,N_3956,N_189);
nand U7877 (N_7877,N_2760,N_3535);
nor U7878 (N_7878,N_3830,N_4567);
nand U7879 (N_7879,N_2126,N_3230);
nand U7880 (N_7880,N_468,N_4887);
or U7881 (N_7881,N_499,N_4874);
xnor U7882 (N_7882,N_706,N_3297);
nor U7883 (N_7883,N_724,N_3251);
nor U7884 (N_7884,N_2300,N_4819);
nand U7885 (N_7885,N_2356,N_3413);
or U7886 (N_7886,N_4793,N_711);
or U7887 (N_7887,N_4447,N_4314);
or U7888 (N_7888,N_836,N_179);
nor U7889 (N_7889,N_1894,N_3748);
or U7890 (N_7890,N_2679,N_3977);
nand U7891 (N_7891,N_2834,N_3570);
or U7892 (N_7892,N_1675,N_2413);
nand U7893 (N_7893,N_178,N_4622);
nor U7894 (N_7894,N_733,N_2215);
or U7895 (N_7895,N_1045,N_78);
or U7896 (N_7896,N_1364,N_3045);
or U7897 (N_7897,N_4719,N_3590);
nor U7898 (N_7898,N_3041,N_2139);
or U7899 (N_7899,N_4930,N_1446);
and U7900 (N_7900,N_1192,N_73);
nand U7901 (N_7901,N_2739,N_1535);
nand U7902 (N_7902,N_4556,N_3698);
nor U7903 (N_7903,N_2172,N_4629);
nor U7904 (N_7904,N_4573,N_4635);
and U7905 (N_7905,N_2661,N_2175);
nor U7906 (N_7906,N_1180,N_1841);
nor U7907 (N_7907,N_3663,N_1754);
nand U7908 (N_7908,N_4035,N_3851);
nor U7909 (N_7909,N_603,N_3282);
nand U7910 (N_7910,N_3714,N_2245);
or U7911 (N_7911,N_4685,N_1790);
and U7912 (N_7912,N_3210,N_2179);
nand U7913 (N_7913,N_4900,N_4878);
or U7914 (N_7914,N_2479,N_2446);
and U7915 (N_7915,N_2336,N_415);
nand U7916 (N_7916,N_3618,N_1778);
and U7917 (N_7917,N_2550,N_1633);
nand U7918 (N_7918,N_4097,N_424);
nor U7919 (N_7919,N_482,N_1666);
nand U7920 (N_7920,N_1443,N_1342);
and U7921 (N_7921,N_3649,N_3462);
nor U7922 (N_7922,N_552,N_4390);
nor U7923 (N_7923,N_3705,N_98);
nand U7924 (N_7924,N_1755,N_4286);
or U7925 (N_7925,N_2190,N_1659);
or U7926 (N_7926,N_3520,N_2703);
or U7927 (N_7927,N_1348,N_981);
or U7928 (N_7928,N_1696,N_1467);
nor U7929 (N_7929,N_3497,N_393);
nor U7930 (N_7930,N_281,N_1959);
or U7931 (N_7931,N_3891,N_994);
nand U7932 (N_7932,N_2719,N_1345);
nor U7933 (N_7933,N_2686,N_1386);
or U7934 (N_7934,N_2273,N_4333);
nor U7935 (N_7935,N_110,N_4824);
or U7936 (N_7936,N_2436,N_1975);
nor U7937 (N_7937,N_1083,N_4913);
nor U7938 (N_7938,N_1437,N_4240);
nand U7939 (N_7939,N_1455,N_1623);
nor U7940 (N_7940,N_969,N_1290);
or U7941 (N_7941,N_4112,N_813);
or U7942 (N_7942,N_96,N_4645);
or U7943 (N_7943,N_4834,N_3189);
nor U7944 (N_7944,N_2384,N_4054);
and U7945 (N_7945,N_3229,N_794);
nor U7946 (N_7946,N_3418,N_759);
and U7947 (N_7947,N_2529,N_2322);
and U7948 (N_7948,N_3651,N_2192);
or U7949 (N_7949,N_282,N_1148);
xnor U7950 (N_7950,N_1456,N_581);
nor U7951 (N_7951,N_4563,N_44);
nor U7952 (N_7952,N_1541,N_433);
and U7953 (N_7953,N_232,N_3420);
nand U7954 (N_7954,N_946,N_1047);
and U7955 (N_7955,N_1042,N_1343);
nor U7956 (N_7956,N_325,N_3775);
nor U7957 (N_7957,N_717,N_4733);
nor U7958 (N_7958,N_3070,N_1029);
nand U7959 (N_7959,N_1747,N_1949);
or U7960 (N_7960,N_4564,N_2925);
or U7961 (N_7961,N_4690,N_1733);
and U7962 (N_7962,N_1993,N_3809);
and U7963 (N_7963,N_3398,N_2645);
or U7964 (N_7964,N_1345,N_1088);
nand U7965 (N_7965,N_4940,N_1933);
nand U7966 (N_7966,N_1747,N_2756);
nor U7967 (N_7967,N_435,N_1783);
nor U7968 (N_7968,N_4416,N_2510);
nand U7969 (N_7969,N_4376,N_762);
nor U7970 (N_7970,N_2171,N_4950);
nor U7971 (N_7971,N_4154,N_4327);
nor U7972 (N_7972,N_839,N_988);
or U7973 (N_7973,N_3285,N_1291);
and U7974 (N_7974,N_3973,N_4891);
and U7975 (N_7975,N_1893,N_1909);
nand U7976 (N_7976,N_4856,N_3267);
and U7977 (N_7977,N_2134,N_3265);
or U7978 (N_7978,N_33,N_1485);
nor U7979 (N_7979,N_2983,N_2698);
and U7980 (N_7980,N_1596,N_4330);
nand U7981 (N_7981,N_1955,N_2678);
nand U7982 (N_7982,N_2622,N_491);
nor U7983 (N_7983,N_2721,N_2522);
nor U7984 (N_7984,N_405,N_3275);
and U7985 (N_7985,N_3723,N_3435);
nor U7986 (N_7986,N_1358,N_3905);
nor U7987 (N_7987,N_945,N_4275);
nand U7988 (N_7988,N_2399,N_3676);
nand U7989 (N_7989,N_1003,N_112);
or U7990 (N_7990,N_2953,N_2011);
nand U7991 (N_7991,N_3832,N_2599);
nand U7992 (N_7992,N_2498,N_4397);
or U7993 (N_7993,N_2604,N_908);
nand U7994 (N_7994,N_3333,N_248);
nand U7995 (N_7995,N_740,N_864);
or U7996 (N_7996,N_52,N_2);
nor U7997 (N_7997,N_3496,N_4426);
nand U7998 (N_7998,N_1815,N_3421);
or U7999 (N_7999,N_3916,N_1620);
nor U8000 (N_8000,N_865,N_2837);
xnor U8001 (N_8001,N_1116,N_4043);
and U8002 (N_8002,N_4093,N_604);
and U8003 (N_8003,N_2668,N_1714);
nand U8004 (N_8004,N_2466,N_630);
nor U8005 (N_8005,N_3659,N_2321);
and U8006 (N_8006,N_4979,N_1865);
nand U8007 (N_8007,N_4355,N_4078);
or U8008 (N_8008,N_1158,N_75);
and U8009 (N_8009,N_1715,N_3623);
nor U8010 (N_8010,N_1025,N_120);
nand U8011 (N_8011,N_3197,N_502);
nand U8012 (N_8012,N_1407,N_816);
nor U8013 (N_8013,N_4568,N_2331);
nor U8014 (N_8014,N_2911,N_4089);
or U8015 (N_8015,N_2146,N_2342);
or U8016 (N_8016,N_4732,N_4226);
or U8017 (N_8017,N_339,N_2423);
xor U8018 (N_8018,N_2617,N_213);
or U8019 (N_8019,N_4517,N_114);
nor U8020 (N_8020,N_4778,N_3121);
and U8021 (N_8021,N_3538,N_2878);
or U8022 (N_8022,N_1067,N_4993);
nor U8023 (N_8023,N_4596,N_3161);
nand U8024 (N_8024,N_3466,N_23);
and U8025 (N_8025,N_3995,N_3286);
or U8026 (N_8026,N_3806,N_3678);
nor U8027 (N_8027,N_4582,N_2148);
and U8028 (N_8028,N_1936,N_2337);
xor U8029 (N_8029,N_3111,N_4076);
and U8030 (N_8030,N_33,N_2900);
nand U8031 (N_8031,N_4920,N_1880);
and U8032 (N_8032,N_1450,N_4359);
nand U8033 (N_8033,N_123,N_1491);
nor U8034 (N_8034,N_4788,N_4879);
nand U8035 (N_8035,N_1723,N_3065);
or U8036 (N_8036,N_2119,N_3437);
nor U8037 (N_8037,N_284,N_4927);
or U8038 (N_8038,N_4458,N_1177);
nor U8039 (N_8039,N_1803,N_3054);
nor U8040 (N_8040,N_565,N_1176);
nor U8041 (N_8041,N_4857,N_4939);
and U8042 (N_8042,N_1420,N_3834);
or U8043 (N_8043,N_3886,N_1635);
and U8044 (N_8044,N_3282,N_4257);
or U8045 (N_8045,N_3040,N_96);
nor U8046 (N_8046,N_3059,N_4994);
nor U8047 (N_8047,N_1194,N_4191);
and U8048 (N_8048,N_1320,N_705);
nor U8049 (N_8049,N_3076,N_3534);
nor U8050 (N_8050,N_4308,N_2193);
and U8051 (N_8051,N_3329,N_2504);
or U8052 (N_8052,N_1353,N_3509);
nand U8053 (N_8053,N_39,N_1990);
nor U8054 (N_8054,N_132,N_4705);
nor U8055 (N_8055,N_2825,N_2555);
nand U8056 (N_8056,N_333,N_2185);
nor U8057 (N_8057,N_1430,N_503);
and U8058 (N_8058,N_869,N_380);
nand U8059 (N_8059,N_427,N_3159);
or U8060 (N_8060,N_2680,N_4861);
nor U8061 (N_8061,N_299,N_542);
nand U8062 (N_8062,N_1680,N_2160);
and U8063 (N_8063,N_1913,N_2651);
or U8064 (N_8064,N_2243,N_4646);
nor U8065 (N_8065,N_2929,N_4257);
or U8066 (N_8066,N_3097,N_4104);
nand U8067 (N_8067,N_3230,N_2043);
and U8068 (N_8068,N_1110,N_1734);
and U8069 (N_8069,N_4418,N_4993);
and U8070 (N_8070,N_45,N_1533);
and U8071 (N_8071,N_3814,N_1889);
and U8072 (N_8072,N_1315,N_3182);
nand U8073 (N_8073,N_3293,N_4710);
nand U8074 (N_8074,N_4744,N_1005);
or U8075 (N_8075,N_4671,N_3205);
or U8076 (N_8076,N_3205,N_2097);
or U8077 (N_8077,N_2757,N_4023);
and U8078 (N_8078,N_606,N_2438);
and U8079 (N_8079,N_4483,N_1792);
and U8080 (N_8080,N_2496,N_2770);
nand U8081 (N_8081,N_4226,N_513);
or U8082 (N_8082,N_4966,N_1083);
nand U8083 (N_8083,N_4328,N_2090);
nor U8084 (N_8084,N_653,N_2432);
nand U8085 (N_8085,N_1112,N_4078);
nand U8086 (N_8086,N_266,N_262);
nand U8087 (N_8087,N_4053,N_4895);
nor U8088 (N_8088,N_2738,N_2483);
nor U8089 (N_8089,N_4689,N_4461);
nand U8090 (N_8090,N_4011,N_4975);
nand U8091 (N_8091,N_3629,N_2735);
nor U8092 (N_8092,N_4114,N_3800);
nor U8093 (N_8093,N_519,N_1790);
or U8094 (N_8094,N_4185,N_889);
and U8095 (N_8095,N_4822,N_2085);
nand U8096 (N_8096,N_1489,N_2608);
nand U8097 (N_8097,N_317,N_1062);
nand U8098 (N_8098,N_1742,N_138);
nor U8099 (N_8099,N_2012,N_4887);
and U8100 (N_8100,N_2010,N_590);
or U8101 (N_8101,N_1338,N_4123);
or U8102 (N_8102,N_751,N_3231);
and U8103 (N_8103,N_506,N_3572);
nor U8104 (N_8104,N_4175,N_1799);
or U8105 (N_8105,N_4608,N_667);
nand U8106 (N_8106,N_156,N_4077);
nand U8107 (N_8107,N_2194,N_105);
or U8108 (N_8108,N_127,N_3700);
and U8109 (N_8109,N_3402,N_1687);
or U8110 (N_8110,N_3347,N_2520);
nor U8111 (N_8111,N_2948,N_4113);
nand U8112 (N_8112,N_1600,N_1322);
nor U8113 (N_8113,N_3311,N_3607);
or U8114 (N_8114,N_4992,N_1603);
xnor U8115 (N_8115,N_4001,N_2783);
nor U8116 (N_8116,N_3090,N_1683);
or U8117 (N_8117,N_468,N_533);
or U8118 (N_8118,N_2705,N_1386);
nor U8119 (N_8119,N_2848,N_3058);
nor U8120 (N_8120,N_4550,N_590);
or U8121 (N_8121,N_4778,N_1723);
nor U8122 (N_8122,N_1109,N_2856);
and U8123 (N_8123,N_3870,N_1140);
nand U8124 (N_8124,N_2749,N_4352);
and U8125 (N_8125,N_3030,N_697);
and U8126 (N_8126,N_3233,N_1793);
nor U8127 (N_8127,N_665,N_4576);
nor U8128 (N_8128,N_1703,N_684);
and U8129 (N_8129,N_3613,N_3040);
nand U8130 (N_8130,N_1335,N_4357);
nand U8131 (N_8131,N_2437,N_1141);
and U8132 (N_8132,N_283,N_105);
or U8133 (N_8133,N_351,N_408);
and U8134 (N_8134,N_1951,N_3442);
nand U8135 (N_8135,N_731,N_1414);
nand U8136 (N_8136,N_1615,N_3227);
nand U8137 (N_8137,N_4059,N_2741);
xnor U8138 (N_8138,N_4715,N_3783);
nor U8139 (N_8139,N_4354,N_1346);
nand U8140 (N_8140,N_4555,N_4741);
and U8141 (N_8141,N_2127,N_1975);
nor U8142 (N_8142,N_3060,N_1251);
or U8143 (N_8143,N_3072,N_3690);
nand U8144 (N_8144,N_1097,N_2757);
nand U8145 (N_8145,N_612,N_2344);
or U8146 (N_8146,N_3820,N_1425);
xnor U8147 (N_8147,N_2796,N_1204);
and U8148 (N_8148,N_2156,N_4078);
xnor U8149 (N_8149,N_108,N_1785);
nor U8150 (N_8150,N_3328,N_1572);
and U8151 (N_8151,N_3474,N_696);
nor U8152 (N_8152,N_253,N_764);
nand U8153 (N_8153,N_2992,N_4256);
and U8154 (N_8154,N_822,N_1007);
nor U8155 (N_8155,N_4372,N_2661);
and U8156 (N_8156,N_3141,N_3217);
nor U8157 (N_8157,N_1182,N_4204);
nand U8158 (N_8158,N_368,N_1173);
and U8159 (N_8159,N_3344,N_3761);
and U8160 (N_8160,N_4681,N_4586);
or U8161 (N_8161,N_3543,N_2718);
or U8162 (N_8162,N_4674,N_4438);
nand U8163 (N_8163,N_571,N_1715);
nor U8164 (N_8164,N_4400,N_1678);
nor U8165 (N_8165,N_1075,N_778);
nand U8166 (N_8166,N_441,N_1152);
xor U8167 (N_8167,N_2636,N_1334);
nor U8168 (N_8168,N_4628,N_3229);
or U8169 (N_8169,N_4347,N_2248);
nand U8170 (N_8170,N_4784,N_2306);
nor U8171 (N_8171,N_4299,N_2676);
or U8172 (N_8172,N_780,N_1549);
nand U8173 (N_8173,N_2464,N_322);
nor U8174 (N_8174,N_4956,N_3009);
or U8175 (N_8175,N_1212,N_3538);
nor U8176 (N_8176,N_4130,N_1963);
or U8177 (N_8177,N_2458,N_2140);
nor U8178 (N_8178,N_762,N_831);
or U8179 (N_8179,N_3876,N_1582);
and U8180 (N_8180,N_4001,N_3525);
and U8181 (N_8181,N_4265,N_3036);
and U8182 (N_8182,N_4803,N_3140);
nor U8183 (N_8183,N_1179,N_2310);
and U8184 (N_8184,N_1010,N_4047);
or U8185 (N_8185,N_4900,N_4584);
and U8186 (N_8186,N_4316,N_2855);
and U8187 (N_8187,N_1805,N_4395);
nand U8188 (N_8188,N_286,N_4630);
and U8189 (N_8189,N_3238,N_580);
and U8190 (N_8190,N_3395,N_3257);
nor U8191 (N_8191,N_3094,N_4269);
or U8192 (N_8192,N_1918,N_3193);
xor U8193 (N_8193,N_991,N_3004);
or U8194 (N_8194,N_3148,N_3489);
or U8195 (N_8195,N_4741,N_2709);
or U8196 (N_8196,N_4753,N_3445);
or U8197 (N_8197,N_2999,N_3407);
and U8198 (N_8198,N_4887,N_3553);
nand U8199 (N_8199,N_4565,N_1110);
nor U8200 (N_8200,N_2950,N_2190);
or U8201 (N_8201,N_1869,N_924);
xnor U8202 (N_8202,N_1281,N_2008);
nand U8203 (N_8203,N_1629,N_483);
or U8204 (N_8204,N_3810,N_2397);
nand U8205 (N_8205,N_1917,N_4735);
or U8206 (N_8206,N_733,N_2885);
nor U8207 (N_8207,N_1542,N_955);
or U8208 (N_8208,N_1713,N_3814);
nor U8209 (N_8209,N_2644,N_3013);
nand U8210 (N_8210,N_1139,N_3121);
nor U8211 (N_8211,N_943,N_2061);
nor U8212 (N_8212,N_1728,N_505);
or U8213 (N_8213,N_4334,N_467);
nand U8214 (N_8214,N_3047,N_384);
or U8215 (N_8215,N_739,N_1900);
nand U8216 (N_8216,N_4417,N_4063);
nor U8217 (N_8217,N_2735,N_4450);
nand U8218 (N_8218,N_2199,N_2432);
or U8219 (N_8219,N_2001,N_319);
nor U8220 (N_8220,N_1095,N_1034);
and U8221 (N_8221,N_4666,N_1824);
or U8222 (N_8222,N_316,N_321);
nand U8223 (N_8223,N_3600,N_2336);
nand U8224 (N_8224,N_119,N_2332);
and U8225 (N_8225,N_2549,N_2412);
or U8226 (N_8226,N_2923,N_2480);
and U8227 (N_8227,N_873,N_1527);
and U8228 (N_8228,N_1078,N_3956);
and U8229 (N_8229,N_342,N_258);
or U8230 (N_8230,N_1954,N_2599);
or U8231 (N_8231,N_2704,N_4794);
and U8232 (N_8232,N_2511,N_4529);
nand U8233 (N_8233,N_1330,N_3755);
nor U8234 (N_8234,N_2488,N_4953);
nand U8235 (N_8235,N_730,N_2690);
or U8236 (N_8236,N_1025,N_4894);
or U8237 (N_8237,N_101,N_1623);
nand U8238 (N_8238,N_2825,N_3645);
or U8239 (N_8239,N_1962,N_1369);
and U8240 (N_8240,N_621,N_3785);
nand U8241 (N_8241,N_3243,N_1370);
nand U8242 (N_8242,N_3776,N_3355);
or U8243 (N_8243,N_3206,N_2400);
nor U8244 (N_8244,N_3748,N_4489);
nand U8245 (N_8245,N_1607,N_4407);
nand U8246 (N_8246,N_3104,N_1090);
nand U8247 (N_8247,N_3863,N_1320);
nor U8248 (N_8248,N_2370,N_3930);
nor U8249 (N_8249,N_3398,N_2652);
or U8250 (N_8250,N_1293,N_2076);
or U8251 (N_8251,N_4139,N_3543);
nand U8252 (N_8252,N_1186,N_2632);
xnor U8253 (N_8253,N_4703,N_4293);
or U8254 (N_8254,N_1936,N_4575);
nand U8255 (N_8255,N_4960,N_3359);
nand U8256 (N_8256,N_1961,N_955);
nand U8257 (N_8257,N_3408,N_1881);
nand U8258 (N_8258,N_1799,N_229);
or U8259 (N_8259,N_4283,N_428);
and U8260 (N_8260,N_2936,N_1787);
nor U8261 (N_8261,N_3933,N_3895);
nand U8262 (N_8262,N_2388,N_1775);
nand U8263 (N_8263,N_4348,N_4201);
nand U8264 (N_8264,N_1276,N_59);
nand U8265 (N_8265,N_1981,N_3866);
nor U8266 (N_8266,N_1951,N_1686);
or U8267 (N_8267,N_1184,N_2278);
nand U8268 (N_8268,N_1500,N_307);
and U8269 (N_8269,N_2535,N_1273);
nor U8270 (N_8270,N_819,N_1235);
or U8271 (N_8271,N_3335,N_3740);
and U8272 (N_8272,N_3395,N_62);
or U8273 (N_8273,N_2674,N_1017);
and U8274 (N_8274,N_3338,N_4275);
nor U8275 (N_8275,N_4316,N_1040);
nor U8276 (N_8276,N_2584,N_2057);
or U8277 (N_8277,N_2857,N_2215);
xor U8278 (N_8278,N_2264,N_927);
and U8279 (N_8279,N_4105,N_78);
or U8280 (N_8280,N_424,N_1885);
nand U8281 (N_8281,N_2407,N_4861);
and U8282 (N_8282,N_1335,N_4995);
or U8283 (N_8283,N_2014,N_2007);
nand U8284 (N_8284,N_4306,N_172);
nor U8285 (N_8285,N_3507,N_697);
or U8286 (N_8286,N_3833,N_3250);
nor U8287 (N_8287,N_3824,N_1271);
nor U8288 (N_8288,N_3384,N_425);
nand U8289 (N_8289,N_3815,N_1859);
nand U8290 (N_8290,N_1737,N_4764);
nor U8291 (N_8291,N_703,N_1902);
or U8292 (N_8292,N_3225,N_4232);
or U8293 (N_8293,N_2396,N_1566);
nand U8294 (N_8294,N_1787,N_1993);
and U8295 (N_8295,N_565,N_2153);
xor U8296 (N_8296,N_1441,N_4296);
nand U8297 (N_8297,N_3197,N_2993);
or U8298 (N_8298,N_1250,N_1272);
nand U8299 (N_8299,N_575,N_3334);
or U8300 (N_8300,N_4030,N_4283);
nor U8301 (N_8301,N_1972,N_435);
or U8302 (N_8302,N_1007,N_836);
and U8303 (N_8303,N_1230,N_4004);
nand U8304 (N_8304,N_4875,N_2651);
xnor U8305 (N_8305,N_3563,N_418);
nor U8306 (N_8306,N_4151,N_465);
nor U8307 (N_8307,N_1616,N_4937);
or U8308 (N_8308,N_3353,N_3432);
or U8309 (N_8309,N_1504,N_2460);
nand U8310 (N_8310,N_4381,N_1338);
nor U8311 (N_8311,N_2825,N_944);
nor U8312 (N_8312,N_2763,N_253);
nand U8313 (N_8313,N_1588,N_2304);
nand U8314 (N_8314,N_3567,N_4510);
nor U8315 (N_8315,N_4001,N_504);
and U8316 (N_8316,N_2203,N_2461);
and U8317 (N_8317,N_4700,N_439);
or U8318 (N_8318,N_411,N_2579);
or U8319 (N_8319,N_4396,N_4189);
or U8320 (N_8320,N_1202,N_3502);
or U8321 (N_8321,N_1181,N_202);
and U8322 (N_8322,N_2513,N_1385);
or U8323 (N_8323,N_2803,N_3865);
or U8324 (N_8324,N_342,N_3323);
or U8325 (N_8325,N_3695,N_4199);
nand U8326 (N_8326,N_1498,N_848);
nand U8327 (N_8327,N_1232,N_385);
nor U8328 (N_8328,N_3473,N_1587);
nor U8329 (N_8329,N_3638,N_894);
and U8330 (N_8330,N_1968,N_3412);
nor U8331 (N_8331,N_3072,N_1187);
and U8332 (N_8332,N_1455,N_519);
or U8333 (N_8333,N_2166,N_119);
nand U8334 (N_8334,N_713,N_3951);
nor U8335 (N_8335,N_1311,N_2331);
nor U8336 (N_8336,N_2523,N_942);
or U8337 (N_8337,N_2918,N_4021);
and U8338 (N_8338,N_234,N_896);
and U8339 (N_8339,N_4117,N_4203);
or U8340 (N_8340,N_1855,N_1807);
nand U8341 (N_8341,N_4430,N_2801);
and U8342 (N_8342,N_4679,N_3721);
nor U8343 (N_8343,N_2821,N_1134);
nor U8344 (N_8344,N_3592,N_4655);
or U8345 (N_8345,N_4594,N_667);
nand U8346 (N_8346,N_3847,N_1376);
or U8347 (N_8347,N_3637,N_253);
or U8348 (N_8348,N_2617,N_1192);
or U8349 (N_8349,N_2559,N_4431);
or U8350 (N_8350,N_4942,N_1728);
and U8351 (N_8351,N_24,N_1484);
nand U8352 (N_8352,N_880,N_4391);
or U8353 (N_8353,N_1741,N_4291);
nand U8354 (N_8354,N_2586,N_4340);
nand U8355 (N_8355,N_2405,N_1820);
and U8356 (N_8356,N_1826,N_1712);
and U8357 (N_8357,N_268,N_3276);
nor U8358 (N_8358,N_3082,N_983);
or U8359 (N_8359,N_4951,N_775);
or U8360 (N_8360,N_3634,N_1640);
and U8361 (N_8361,N_1456,N_2790);
nor U8362 (N_8362,N_2850,N_2317);
nor U8363 (N_8363,N_4248,N_3241);
nor U8364 (N_8364,N_1165,N_674);
nor U8365 (N_8365,N_712,N_2783);
nand U8366 (N_8366,N_2366,N_3987);
and U8367 (N_8367,N_4240,N_779);
nand U8368 (N_8368,N_1752,N_1048);
nand U8369 (N_8369,N_321,N_3605);
nor U8370 (N_8370,N_648,N_2962);
nand U8371 (N_8371,N_1048,N_1514);
or U8372 (N_8372,N_2314,N_376);
and U8373 (N_8373,N_1966,N_1034);
and U8374 (N_8374,N_3139,N_676);
or U8375 (N_8375,N_4777,N_1636);
and U8376 (N_8376,N_1885,N_1431);
or U8377 (N_8377,N_825,N_2598);
or U8378 (N_8378,N_4882,N_3988);
and U8379 (N_8379,N_261,N_4338);
or U8380 (N_8380,N_4288,N_967);
nand U8381 (N_8381,N_576,N_1403);
or U8382 (N_8382,N_2407,N_2113);
or U8383 (N_8383,N_1399,N_3718);
and U8384 (N_8384,N_2037,N_4005);
nor U8385 (N_8385,N_1176,N_1284);
nand U8386 (N_8386,N_4271,N_51);
nand U8387 (N_8387,N_4712,N_3670);
nor U8388 (N_8388,N_1084,N_4636);
nor U8389 (N_8389,N_1157,N_2497);
and U8390 (N_8390,N_2449,N_4285);
and U8391 (N_8391,N_1820,N_792);
nand U8392 (N_8392,N_2366,N_2521);
and U8393 (N_8393,N_2079,N_4340);
or U8394 (N_8394,N_893,N_4025);
and U8395 (N_8395,N_2165,N_1201);
nand U8396 (N_8396,N_932,N_2210);
nor U8397 (N_8397,N_531,N_824);
or U8398 (N_8398,N_1522,N_864);
nand U8399 (N_8399,N_1950,N_4160);
or U8400 (N_8400,N_2186,N_3990);
nand U8401 (N_8401,N_2824,N_1726);
or U8402 (N_8402,N_2378,N_1174);
and U8403 (N_8403,N_4865,N_3073);
xnor U8404 (N_8404,N_4003,N_1837);
or U8405 (N_8405,N_2951,N_3552);
nor U8406 (N_8406,N_540,N_3677);
nor U8407 (N_8407,N_1769,N_571);
and U8408 (N_8408,N_3663,N_3300);
nor U8409 (N_8409,N_564,N_4609);
or U8410 (N_8410,N_192,N_1752);
nor U8411 (N_8411,N_2047,N_1133);
nand U8412 (N_8412,N_1756,N_3671);
or U8413 (N_8413,N_4918,N_4295);
nor U8414 (N_8414,N_4904,N_1014);
or U8415 (N_8415,N_3801,N_4692);
and U8416 (N_8416,N_3238,N_4830);
xor U8417 (N_8417,N_1788,N_4196);
or U8418 (N_8418,N_2916,N_1695);
or U8419 (N_8419,N_1665,N_3515);
nor U8420 (N_8420,N_373,N_559);
nand U8421 (N_8421,N_1971,N_3633);
nand U8422 (N_8422,N_2451,N_2196);
and U8423 (N_8423,N_3613,N_3515);
nor U8424 (N_8424,N_4483,N_431);
or U8425 (N_8425,N_4773,N_3983);
nor U8426 (N_8426,N_332,N_3874);
or U8427 (N_8427,N_2301,N_1249);
nor U8428 (N_8428,N_4476,N_934);
or U8429 (N_8429,N_1225,N_3009);
and U8430 (N_8430,N_103,N_195);
nand U8431 (N_8431,N_972,N_2652);
nor U8432 (N_8432,N_3104,N_1050);
nor U8433 (N_8433,N_4234,N_4688);
xnor U8434 (N_8434,N_2670,N_4297);
nand U8435 (N_8435,N_3185,N_1322);
nor U8436 (N_8436,N_3271,N_384);
and U8437 (N_8437,N_4934,N_2635);
or U8438 (N_8438,N_641,N_820);
nand U8439 (N_8439,N_984,N_3049);
nand U8440 (N_8440,N_1286,N_1479);
nor U8441 (N_8441,N_4291,N_976);
nand U8442 (N_8442,N_3688,N_3944);
nor U8443 (N_8443,N_3146,N_3913);
and U8444 (N_8444,N_872,N_3358);
nor U8445 (N_8445,N_627,N_2290);
nand U8446 (N_8446,N_4090,N_558);
nor U8447 (N_8447,N_3742,N_4428);
nor U8448 (N_8448,N_3522,N_4000);
nor U8449 (N_8449,N_3486,N_4252);
nor U8450 (N_8450,N_1164,N_4118);
nor U8451 (N_8451,N_1981,N_4664);
nand U8452 (N_8452,N_1684,N_2805);
or U8453 (N_8453,N_1535,N_1029);
nor U8454 (N_8454,N_2550,N_271);
nor U8455 (N_8455,N_1095,N_3699);
nor U8456 (N_8456,N_2121,N_4465);
and U8457 (N_8457,N_885,N_1140);
nand U8458 (N_8458,N_2736,N_4863);
nand U8459 (N_8459,N_646,N_76);
or U8460 (N_8460,N_3454,N_3823);
or U8461 (N_8461,N_4507,N_1671);
nand U8462 (N_8462,N_4489,N_3378);
nand U8463 (N_8463,N_4312,N_2580);
and U8464 (N_8464,N_2603,N_3783);
and U8465 (N_8465,N_1742,N_4880);
or U8466 (N_8466,N_1653,N_705);
and U8467 (N_8467,N_2327,N_2865);
or U8468 (N_8468,N_3561,N_3201);
nand U8469 (N_8469,N_834,N_2358);
or U8470 (N_8470,N_634,N_2846);
nor U8471 (N_8471,N_4899,N_1046);
and U8472 (N_8472,N_1793,N_898);
and U8473 (N_8473,N_580,N_1004);
and U8474 (N_8474,N_1391,N_2758);
or U8475 (N_8475,N_686,N_3012);
nor U8476 (N_8476,N_2772,N_1648);
or U8477 (N_8477,N_1975,N_3564);
or U8478 (N_8478,N_411,N_3446);
or U8479 (N_8479,N_3883,N_1103);
nor U8480 (N_8480,N_352,N_2881);
nor U8481 (N_8481,N_2366,N_2867);
or U8482 (N_8482,N_4485,N_2192);
nand U8483 (N_8483,N_3450,N_2212);
nor U8484 (N_8484,N_1610,N_2211);
and U8485 (N_8485,N_4445,N_2234);
or U8486 (N_8486,N_1922,N_113);
or U8487 (N_8487,N_189,N_1272);
nor U8488 (N_8488,N_687,N_839);
nand U8489 (N_8489,N_3606,N_3792);
nor U8490 (N_8490,N_1689,N_4340);
nor U8491 (N_8491,N_2524,N_1494);
nor U8492 (N_8492,N_1324,N_1734);
or U8493 (N_8493,N_3963,N_135);
or U8494 (N_8494,N_493,N_354);
or U8495 (N_8495,N_4772,N_1905);
or U8496 (N_8496,N_3537,N_4447);
or U8497 (N_8497,N_4427,N_2701);
and U8498 (N_8498,N_3872,N_4268);
nor U8499 (N_8499,N_1125,N_1595);
and U8500 (N_8500,N_4491,N_855);
and U8501 (N_8501,N_390,N_2056);
or U8502 (N_8502,N_1711,N_1938);
nand U8503 (N_8503,N_2858,N_1260);
and U8504 (N_8504,N_4419,N_1606);
nor U8505 (N_8505,N_2462,N_1262);
nand U8506 (N_8506,N_4955,N_3743);
or U8507 (N_8507,N_887,N_3277);
and U8508 (N_8508,N_3979,N_4025);
nor U8509 (N_8509,N_709,N_3121);
nor U8510 (N_8510,N_3213,N_1354);
and U8511 (N_8511,N_695,N_4640);
and U8512 (N_8512,N_4599,N_2633);
and U8513 (N_8513,N_2281,N_1330);
nor U8514 (N_8514,N_2757,N_446);
nand U8515 (N_8515,N_722,N_761);
and U8516 (N_8516,N_4570,N_3781);
and U8517 (N_8517,N_251,N_2259);
nor U8518 (N_8518,N_4424,N_3904);
nor U8519 (N_8519,N_261,N_1300);
nand U8520 (N_8520,N_796,N_4594);
or U8521 (N_8521,N_4350,N_2876);
nor U8522 (N_8522,N_2148,N_386);
or U8523 (N_8523,N_2431,N_4773);
or U8524 (N_8524,N_2060,N_1417);
and U8525 (N_8525,N_11,N_3646);
nand U8526 (N_8526,N_640,N_2068);
nand U8527 (N_8527,N_3842,N_742);
nand U8528 (N_8528,N_3891,N_2553);
nand U8529 (N_8529,N_2304,N_4968);
and U8530 (N_8530,N_3262,N_1457);
or U8531 (N_8531,N_3027,N_2631);
and U8532 (N_8532,N_578,N_831);
or U8533 (N_8533,N_2905,N_4839);
nand U8534 (N_8534,N_1474,N_1914);
nand U8535 (N_8535,N_1362,N_3569);
nor U8536 (N_8536,N_2869,N_3262);
and U8537 (N_8537,N_3055,N_1260);
and U8538 (N_8538,N_2024,N_1271);
or U8539 (N_8539,N_2510,N_167);
nand U8540 (N_8540,N_1874,N_409);
xor U8541 (N_8541,N_1505,N_4856);
or U8542 (N_8542,N_3437,N_3447);
nand U8543 (N_8543,N_3682,N_1014);
or U8544 (N_8544,N_4966,N_2401);
nor U8545 (N_8545,N_4430,N_2693);
nand U8546 (N_8546,N_1113,N_2782);
nand U8547 (N_8547,N_1609,N_4053);
and U8548 (N_8548,N_3110,N_2127);
nor U8549 (N_8549,N_668,N_2250);
nand U8550 (N_8550,N_3666,N_769);
xnor U8551 (N_8551,N_1967,N_1256);
nand U8552 (N_8552,N_3425,N_60);
or U8553 (N_8553,N_3034,N_4420);
and U8554 (N_8554,N_51,N_4706);
and U8555 (N_8555,N_1219,N_2223);
nand U8556 (N_8556,N_4513,N_139);
and U8557 (N_8557,N_4009,N_2661);
and U8558 (N_8558,N_3819,N_1547);
and U8559 (N_8559,N_2990,N_4170);
and U8560 (N_8560,N_2187,N_4798);
nand U8561 (N_8561,N_280,N_3771);
and U8562 (N_8562,N_3817,N_3787);
nor U8563 (N_8563,N_174,N_4123);
or U8564 (N_8564,N_3266,N_2076);
nor U8565 (N_8565,N_3927,N_3439);
and U8566 (N_8566,N_93,N_4134);
and U8567 (N_8567,N_2103,N_3573);
nor U8568 (N_8568,N_3806,N_3320);
nand U8569 (N_8569,N_2252,N_275);
or U8570 (N_8570,N_1640,N_3934);
or U8571 (N_8571,N_3197,N_4764);
nand U8572 (N_8572,N_4361,N_3389);
nor U8573 (N_8573,N_197,N_2268);
nand U8574 (N_8574,N_3513,N_3609);
nor U8575 (N_8575,N_3253,N_1170);
nor U8576 (N_8576,N_705,N_4334);
or U8577 (N_8577,N_2623,N_2721);
and U8578 (N_8578,N_648,N_2415);
and U8579 (N_8579,N_239,N_36);
nor U8580 (N_8580,N_4144,N_1704);
or U8581 (N_8581,N_3834,N_3315);
or U8582 (N_8582,N_3863,N_1033);
xnor U8583 (N_8583,N_1294,N_3851);
and U8584 (N_8584,N_703,N_706);
and U8585 (N_8585,N_4507,N_3441);
nor U8586 (N_8586,N_2626,N_4773);
or U8587 (N_8587,N_1023,N_4426);
nor U8588 (N_8588,N_225,N_216);
and U8589 (N_8589,N_2099,N_3359);
nor U8590 (N_8590,N_524,N_2072);
and U8591 (N_8591,N_2624,N_3984);
and U8592 (N_8592,N_480,N_2544);
nand U8593 (N_8593,N_4848,N_2670);
nand U8594 (N_8594,N_544,N_4349);
and U8595 (N_8595,N_2830,N_4277);
nor U8596 (N_8596,N_3623,N_3564);
nor U8597 (N_8597,N_3118,N_4941);
and U8598 (N_8598,N_4426,N_1479);
or U8599 (N_8599,N_1103,N_2218);
nor U8600 (N_8600,N_3451,N_3528);
or U8601 (N_8601,N_1309,N_1567);
or U8602 (N_8602,N_4179,N_691);
and U8603 (N_8603,N_318,N_695);
nand U8604 (N_8604,N_4925,N_722);
and U8605 (N_8605,N_957,N_3999);
xnor U8606 (N_8606,N_2735,N_4852);
nand U8607 (N_8607,N_901,N_352);
nor U8608 (N_8608,N_1747,N_1283);
or U8609 (N_8609,N_2000,N_0);
nand U8610 (N_8610,N_2405,N_2678);
or U8611 (N_8611,N_4612,N_202);
xor U8612 (N_8612,N_1175,N_3679);
nor U8613 (N_8613,N_3295,N_4206);
nor U8614 (N_8614,N_1667,N_2497);
nor U8615 (N_8615,N_4203,N_753);
and U8616 (N_8616,N_4419,N_4397);
nand U8617 (N_8617,N_1837,N_1931);
nor U8618 (N_8618,N_3280,N_3867);
and U8619 (N_8619,N_1137,N_1676);
nand U8620 (N_8620,N_819,N_1924);
and U8621 (N_8621,N_1635,N_4802);
or U8622 (N_8622,N_3521,N_4622);
or U8623 (N_8623,N_758,N_2573);
nand U8624 (N_8624,N_2245,N_2501);
nand U8625 (N_8625,N_4706,N_3190);
nand U8626 (N_8626,N_3517,N_2501);
and U8627 (N_8627,N_1540,N_2246);
nor U8628 (N_8628,N_647,N_4104);
nand U8629 (N_8629,N_69,N_2390);
and U8630 (N_8630,N_745,N_1904);
nor U8631 (N_8631,N_3977,N_1938);
or U8632 (N_8632,N_4030,N_4717);
or U8633 (N_8633,N_4711,N_3621);
nand U8634 (N_8634,N_3261,N_2638);
or U8635 (N_8635,N_3777,N_173);
nor U8636 (N_8636,N_1438,N_3029);
nor U8637 (N_8637,N_199,N_1872);
and U8638 (N_8638,N_508,N_1626);
nor U8639 (N_8639,N_93,N_1480);
and U8640 (N_8640,N_2563,N_2237);
nor U8641 (N_8641,N_2309,N_2039);
or U8642 (N_8642,N_1546,N_2443);
nor U8643 (N_8643,N_1034,N_4440);
nand U8644 (N_8644,N_2784,N_887);
and U8645 (N_8645,N_3458,N_3804);
nand U8646 (N_8646,N_1553,N_4717);
nor U8647 (N_8647,N_2626,N_276);
or U8648 (N_8648,N_2551,N_4212);
or U8649 (N_8649,N_3953,N_4257);
nand U8650 (N_8650,N_462,N_3145);
nand U8651 (N_8651,N_2408,N_3698);
and U8652 (N_8652,N_3118,N_2031);
nor U8653 (N_8653,N_1545,N_3536);
nand U8654 (N_8654,N_959,N_2970);
xor U8655 (N_8655,N_3678,N_1283);
nand U8656 (N_8656,N_2960,N_2329);
and U8657 (N_8657,N_2846,N_2806);
nand U8658 (N_8658,N_1311,N_2287);
or U8659 (N_8659,N_3687,N_2110);
and U8660 (N_8660,N_2737,N_4200);
nor U8661 (N_8661,N_4305,N_2700);
nand U8662 (N_8662,N_3633,N_1088);
and U8663 (N_8663,N_2201,N_3129);
or U8664 (N_8664,N_2924,N_2063);
and U8665 (N_8665,N_1029,N_876);
nand U8666 (N_8666,N_1848,N_1103);
nor U8667 (N_8667,N_1068,N_1936);
nor U8668 (N_8668,N_4084,N_4033);
and U8669 (N_8669,N_4819,N_4583);
nand U8670 (N_8670,N_616,N_1018);
or U8671 (N_8671,N_4476,N_1788);
xnor U8672 (N_8672,N_1254,N_2413);
and U8673 (N_8673,N_762,N_4207);
or U8674 (N_8674,N_3593,N_1026);
nor U8675 (N_8675,N_674,N_332);
and U8676 (N_8676,N_3398,N_4422);
or U8677 (N_8677,N_2664,N_2598);
or U8678 (N_8678,N_3390,N_2561);
or U8679 (N_8679,N_3892,N_2679);
nand U8680 (N_8680,N_1833,N_4535);
nor U8681 (N_8681,N_3388,N_84);
nor U8682 (N_8682,N_4086,N_1703);
and U8683 (N_8683,N_2818,N_263);
and U8684 (N_8684,N_4958,N_3887);
or U8685 (N_8685,N_1386,N_817);
and U8686 (N_8686,N_3789,N_2288);
nand U8687 (N_8687,N_2537,N_4577);
nor U8688 (N_8688,N_1953,N_3635);
nor U8689 (N_8689,N_1070,N_4293);
nor U8690 (N_8690,N_486,N_3558);
nor U8691 (N_8691,N_3830,N_2451);
and U8692 (N_8692,N_4476,N_4134);
nor U8693 (N_8693,N_3669,N_1921);
nor U8694 (N_8694,N_3898,N_3217);
nand U8695 (N_8695,N_3810,N_772);
nand U8696 (N_8696,N_2894,N_3515);
or U8697 (N_8697,N_856,N_3220);
nor U8698 (N_8698,N_757,N_671);
nand U8699 (N_8699,N_2044,N_1345);
nand U8700 (N_8700,N_2281,N_4971);
or U8701 (N_8701,N_2745,N_3770);
nor U8702 (N_8702,N_3864,N_4074);
nor U8703 (N_8703,N_3720,N_1072);
nor U8704 (N_8704,N_1857,N_3001);
nand U8705 (N_8705,N_1896,N_589);
and U8706 (N_8706,N_1958,N_1355);
or U8707 (N_8707,N_1741,N_842);
nand U8708 (N_8708,N_4508,N_4313);
or U8709 (N_8709,N_629,N_469);
and U8710 (N_8710,N_3732,N_3784);
nand U8711 (N_8711,N_3425,N_2154);
nor U8712 (N_8712,N_3007,N_3772);
and U8713 (N_8713,N_3144,N_1035);
or U8714 (N_8714,N_1246,N_4641);
and U8715 (N_8715,N_3788,N_3536);
xor U8716 (N_8716,N_391,N_957);
and U8717 (N_8717,N_4799,N_4655);
nand U8718 (N_8718,N_867,N_1926);
nor U8719 (N_8719,N_2115,N_136);
nand U8720 (N_8720,N_69,N_4538);
nor U8721 (N_8721,N_3816,N_494);
nand U8722 (N_8722,N_547,N_2065);
and U8723 (N_8723,N_1263,N_2085);
nand U8724 (N_8724,N_4426,N_3838);
or U8725 (N_8725,N_294,N_4231);
or U8726 (N_8726,N_4232,N_1430);
and U8727 (N_8727,N_268,N_3529);
and U8728 (N_8728,N_2380,N_1258);
nand U8729 (N_8729,N_3955,N_457);
nor U8730 (N_8730,N_1975,N_807);
and U8731 (N_8731,N_4388,N_1905);
and U8732 (N_8732,N_4352,N_3789);
nor U8733 (N_8733,N_2566,N_3013);
xor U8734 (N_8734,N_913,N_3789);
nor U8735 (N_8735,N_1576,N_2471);
and U8736 (N_8736,N_3303,N_3353);
nor U8737 (N_8737,N_1107,N_2766);
and U8738 (N_8738,N_1411,N_4029);
nand U8739 (N_8739,N_1827,N_1067);
or U8740 (N_8740,N_4317,N_4261);
nor U8741 (N_8741,N_4052,N_4780);
or U8742 (N_8742,N_4220,N_2169);
nand U8743 (N_8743,N_1369,N_2759);
nor U8744 (N_8744,N_2402,N_883);
nand U8745 (N_8745,N_4335,N_734);
nor U8746 (N_8746,N_4717,N_461);
nand U8747 (N_8747,N_608,N_4226);
nor U8748 (N_8748,N_4203,N_3596);
and U8749 (N_8749,N_2745,N_977);
and U8750 (N_8750,N_2222,N_1368);
and U8751 (N_8751,N_2359,N_1533);
and U8752 (N_8752,N_4197,N_501);
nor U8753 (N_8753,N_2162,N_2332);
or U8754 (N_8754,N_2682,N_2031);
nor U8755 (N_8755,N_3746,N_19);
and U8756 (N_8756,N_3165,N_3763);
nand U8757 (N_8757,N_4966,N_368);
and U8758 (N_8758,N_771,N_3879);
nor U8759 (N_8759,N_2368,N_3564);
or U8760 (N_8760,N_612,N_3324);
or U8761 (N_8761,N_89,N_964);
or U8762 (N_8762,N_910,N_1215);
and U8763 (N_8763,N_4344,N_390);
and U8764 (N_8764,N_2920,N_672);
nor U8765 (N_8765,N_2570,N_3286);
xor U8766 (N_8766,N_828,N_3780);
nor U8767 (N_8767,N_3208,N_431);
or U8768 (N_8768,N_99,N_3738);
nor U8769 (N_8769,N_3656,N_1351);
nor U8770 (N_8770,N_4575,N_1536);
or U8771 (N_8771,N_1026,N_4151);
nand U8772 (N_8772,N_3990,N_2266);
and U8773 (N_8773,N_4088,N_2539);
or U8774 (N_8774,N_4405,N_1481);
nand U8775 (N_8775,N_1651,N_1485);
or U8776 (N_8776,N_911,N_3008);
or U8777 (N_8777,N_3950,N_4699);
and U8778 (N_8778,N_4037,N_2494);
nand U8779 (N_8779,N_579,N_495);
and U8780 (N_8780,N_3523,N_332);
nor U8781 (N_8781,N_3691,N_63);
and U8782 (N_8782,N_1265,N_3480);
or U8783 (N_8783,N_2072,N_4768);
nor U8784 (N_8784,N_1571,N_4334);
and U8785 (N_8785,N_2922,N_2447);
xnor U8786 (N_8786,N_3297,N_1242);
nor U8787 (N_8787,N_827,N_2558);
nand U8788 (N_8788,N_4559,N_4188);
nor U8789 (N_8789,N_2890,N_2882);
and U8790 (N_8790,N_864,N_2218);
and U8791 (N_8791,N_375,N_1250);
or U8792 (N_8792,N_4837,N_608);
or U8793 (N_8793,N_91,N_3566);
and U8794 (N_8794,N_57,N_1701);
nor U8795 (N_8795,N_3604,N_3790);
nor U8796 (N_8796,N_2769,N_718);
and U8797 (N_8797,N_1378,N_4001);
and U8798 (N_8798,N_4337,N_2303);
xnor U8799 (N_8799,N_175,N_3202);
or U8800 (N_8800,N_3351,N_3034);
or U8801 (N_8801,N_2417,N_4987);
or U8802 (N_8802,N_4616,N_2933);
and U8803 (N_8803,N_3102,N_399);
or U8804 (N_8804,N_2125,N_3546);
or U8805 (N_8805,N_340,N_1013);
or U8806 (N_8806,N_866,N_4689);
and U8807 (N_8807,N_877,N_149);
or U8808 (N_8808,N_4638,N_1709);
or U8809 (N_8809,N_2251,N_1899);
or U8810 (N_8810,N_2939,N_1109);
nand U8811 (N_8811,N_192,N_3500);
and U8812 (N_8812,N_2619,N_4788);
nand U8813 (N_8813,N_3653,N_2160);
nand U8814 (N_8814,N_1556,N_3197);
and U8815 (N_8815,N_2620,N_259);
nor U8816 (N_8816,N_2698,N_3907);
nand U8817 (N_8817,N_3732,N_2252);
nor U8818 (N_8818,N_3692,N_1815);
nor U8819 (N_8819,N_3636,N_2529);
xor U8820 (N_8820,N_1914,N_972);
nor U8821 (N_8821,N_4183,N_3779);
nor U8822 (N_8822,N_3557,N_4898);
or U8823 (N_8823,N_4610,N_2086);
or U8824 (N_8824,N_2641,N_1510);
nor U8825 (N_8825,N_1208,N_4644);
nand U8826 (N_8826,N_1958,N_2832);
nor U8827 (N_8827,N_678,N_1604);
or U8828 (N_8828,N_3398,N_3376);
nand U8829 (N_8829,N_1535,N_2449);
and U8830 (N_8830,N_3360,N_4338);
nand U8831 (N_8831,N_4433,N_4774);
nor U8832 (N_8832,N_1097,N_3388);
and U8833 (N_8833,N_4577,N_981);
nand U8834 (N_8834,N_113,N_3946);
nand U8835 (N_8835,N_941,N_2406);
and U8836 (N_8836,N_1180,N_695);
nor U8837 (N_8837,N_4133,N_3890);
nor U8838 (N_8838,N_4769,N_985);
nand U8839 (N_8839,N_443,N_2517);
and U8840 (N_8840,N_2491,N_4272);
and U8841 (N_8841,N_1437,N_4751);
or U8842 (N_8842,N_1511,N_2674);
nand U8843 (N_8843,N_938,N_1081);
nand U8844 (N_8844,N_697,N_1469);
nand U8845 (N_8845,N_3681,N_435);
and U8846 (N_8846,N_2341,N_4065);
nand U8847 (N_8847,N_1970,N_288);
or U8848 (N_8848,N_2985,N_1191);
nand U8849 (N_8849,N_2166,N_1894);
or U8850 (N_8850,N_3014,N_689);
nand U8851 (N_8851,N_1553,N_463);
or U8852 (N_8852,N_1789,N_2505);
or U8853 (N_8853,N_1817,N_4539);
or U8854 (N_8854,N_1590,N_2944);
and U8855 (N_8855,N_2983,N_3714);
or U8856 (N_8856,N_560,N_708);
xor U8857 (N_8857,N_3982,N_4311);
or U8858 (N_8858,N_2664,N_2379);
nand U8859 (N_8859,N_1243,N_3088);
nor U8860 (N_8860,N_2540,N_132);
and U8861 (N_8861,N_2084,N_3841);
nor U8862 (N_8862,N_2999,N_2321);
or U8863 (N_8863,N_1331,N_3780);
nand U8864 (N_8864,N_85,N_3767);
nand U8865 (N_8865,N_3732,N_4581);
nand U8866 (N_8866,N_3365,N_618);
nor U8867 (N_8867,N_4825,N_2626);
and U8868 (N_8868,N_3813,N_2840);
nor U8869 (N_8869,N_652,N_2031);
or U8870 (N_8870,N_4022,N_1450);
nor U8871 (N_8871,N_468,N_453);
and U8872 (N_8872,N_4725,N_682);
and U8873 (N_8873,N_1707,N_2842);
xor U8874 (N_8874,N_831,N_2397);
or U8875 (N_8875,N_1098,N_355);
nand U8876 (N_8876,N_1147,N_3348);
and U8877 (N_8877,N_301,N_3021);
and U8878 (N_8878,N_2484,N_3503);
or U8879 (N_8879,N_3087,N_4413);
nand U8880 (N_8880,N_1201,N_2348);
nand U8881 (N_8881,N_3706,N_1133);
and U8882 (N_8882,N_872,N_2826);
and U8883 (N_8883,N_180,N_3773);
or U8884 (N_8884,N_4945,N_3369);
or U8885 (N_8885,N_4185,N_3542);
nor U8886 (N_8886,N_1436,N_3075);
nor U8887 (N_8887,N_3911,N_4163);
and U8888 (N_8888,N_3777,N_503);
and U8889 (N_8889,N_1192,N_408);
or U8890 (N_8890,N_4503,N_2508);
and U8891 (N_8891,N_1797,N_3959);
and U8892 (N_8892,N_708,N_1770);
nor U8893 (N_8893,N_3299,N_856);
and U8894 (N_8894,N_4066,N_2311);
nand U8895 (N_8895,N_3567,N_1073);
nor U8896 (N_8896,N_3452,N_4066);
nand U8897 (N_8897,N_4946,N_2338);
and U8898 (N_8898,N_3624,N_62);
and U8899 (N_8899,N_3654,N_3262);
nand U8900 (N_8900,N_3534,N_3183);
and U8901 (N_8901,N_1788,N_1537);
nor U8902 (N_8902,N_4841,N_1814);
nor U8903 (N_8903,N_4970,N_4379);
or U8904 (N_8904,N_3776,N_640);
or U8905 (N_8905,N_1045,N_2529);
or U8906 (N_8906,N_4036,N_1914);
and U8907 (N_8907,N_1529,N_2283);
or U8908 (N_8908,N_1578,N_1163);
and U8909 (N_8909,N_3121,N_3278);
nand U8910 (N_8910,N_397,N_115);
nand U8911 (N_8911,N_2628,N_1528);
nand U8912 (N_8912,N_565,N_3995);
and U8913 (N_8913,N_3573,N_771);
nor U8914 (N_8914,N_4139,N_1351);
and U8915 (N_8915,N_3480,N_2643);
or U8916 (N_8916,N_1388,N_2462);
and U8917 (N_8917,N_4227,N_651);
and U8918 (N_8918,N_169,N_442);
and U8919 (N_8919,N_270,N_1901);
and U8920 (N_8920,N_801,N_2190);
nor U8921 (N_8921,N_1001,N_697);
and U8922 (N_8922,N_1899,N_2456);
nand U8923 (N_8923,N_1967,N_3039);
nor U8924 (N_8924,N_2118,N_62);
and U8925 (N_8925,N_1886,N_4707);
nor U8926 (N_8926,N_2638,N_156);
nand U8927 (N_8927,N_280,N_1900);
nand U8928 (N_8928,N_2190,N_4412);
nand U8929 (N_8929,N_3063,N_3995);
nor U8930 (N_8930,N_973,N_1546);
nor U8931 (N_8931,N_901,N_2959);
or U8932 (N_8932,N_4080,N_997);
and U8933 (N_8933,N_4995,N_3000);
nand U8934 (N_8934,N_1403,N_2122);
and U8935 (N_8935,N_2757,N_2788);
or U8936 (N_8936,N_2561,N_4828);
and U8937 (N_8937,N_4441,N_1962);
nor U8938 (N_8938,N_1926,N_1721);
xor U8939 (N_8939,N_49,N_36);
nor U8940 (N_8940,N_4027,N_3525);
nand U8941 (N_8941,N_4434,N_3419);
nand U8942 (N_8942,N_4829,N_1188);
or U8943 (N_8943,N_4554,N_4422);
nand U8944 (N_8944,N_1433,N_3816);
nor U8945 (N_8945,N_3479,N_732);
and U8946 (N_8946,N_1315,N_4002);
or U8947 (N_8947,N_3827,N_1925);
or U8948 (N_8948,N_335,N_330);
nand U8949 (N_8949,N_330,N_1313);
nand U8950 (N_8950,N_4426,N_2610);
nor U8951 (N_8951,N_3362,N_3947);
nand U8952 (N_8952,N_65,N_3448);
nor U8953 (N_8953,N_3185,N_2861);
or U8954 (N_8954,N_4138,N_228);
or U8955 (N_8955,N_1509,N_1078);
and U8956 (N_8956,N_4062,N_2060);
nor U8957 (N_8957,N_4807,N_2344);
nand U8958 (N_8958,N_1021,N_4490);
or U8959 (N_8959,N_2903,N_1754);
or U8960 (N_8960,N_3356,N_955);
or U8961 (N_8961,N_1795,N_55);
xor U8962 (N_8962,N_1508,N_4090);
and U8963 (N_8963,N_1113,N_2288);
nor U8964 (N_8964,N_523,N_679);
nor U8965 (N_8965,N_288,N_346);
nand U8966 (N_8966,N_4652,N_3240);
xor U8967 (N_8967,N_1312,N_3009);
nor U8968 (N_8968,N_4146,N_1174);
nor U8969 (N_8969,N_2090,N_2983);
nor U8970 (N_8970,N_3631,N_4574);
nor U8971 (N_8971,N_2565,N_3012);
or U8972 (N_8972,N_4367,N_317);
or U8973 (N_8973,N_3305,N_130);
or U8974 (N_8974,N_3632,N_1911);
nand U8975 (N_8975,N_3350,N_3935);
nor U8976 (N_8976,N_3176,N_1908);
nor U8977 (N_8977,N_4933,N_707);
and U8978 (N_8978,N_196,N_1044);
and U8979 (N_8979,N_4396,N_1726);
and U8980 (N_8980,N_516,N_86);
and U8981 (N_8981,N_3830,N_1371);
nand U8982 (N_8982,N_2232,N_3844);
and U8983 (N_8983,N_3532,N_2059);
nor U8984 (N_8984,N_2234,N_3521);
nand U8985 (N_8985,N_1888,N_300);
nand U8986 (N_8986,N_703,N_3101);
and U8987 (N_8987,N_3011,N_2635);
and U8988 (N_8988,N_56,N_4377);
or U8989 (N_8989,N_1017,N_1764);
nor U8990 (N_8990,N_4762,N_2017);
nor U8991 (N_8991,N_1699,N_4727);
nand U8992 (N_8992,N_1512,N_571);
nor U8993 (N_8993,N_3606,N_4055);
nand U8994 (N_8994,N_3143,N_862);
or U8995 (N_8995,N_3745,N_255);
and U8996 (N_8996,N_2378,N_2999);
or U8997 (N_8997,N_2055,N_2971);
xor U8998 (N_8998,N_3457,N_3412);
and U8999 (N_8999,N_3314,N_1805);
nor U9000 (N_9000,N_3866,N_113);
nand U9001 (N_9001,N_2224,N_893);
nor U9002 (N_9002,N_3039,N_2343);
or U9003 (N_9003,N_777,N_2628);
and U9004 (N_9004,N_1270,N_504);
nor U9005 (N_9005,N_1858,N_570);
nand U9006 (N_9006,N_526,N_859);
nand U9007 (N_9007,N_920,N_104);
nand U9008 (N_9008,N_4596,N_4844);
nand U9009 (N_9009,N_3310,N_106);
nor U9010 (N_9010,N_2583,N_10);
and U9011 (N_9011,N_1083,N_898);
or U9012 (N_9012,N_229,N_3511);
and U9013 (N_9013,N_2804,N_2732);
nor U9014 (N_9014,N_3074,N_1099);
nand U9015 (N_9015,N_1886,N_4810);
and U9016 (N_9016,N_1315,N_3137);
nor U9017 (N_9017,N_2955,N_635);
and U9018 (N_9018,N_4333,N_1507);
or U9019 (N_9019,N_577,N_2553);
or U9020 (N_9020,N_3240,N_4943);
and U9021 (N_9021,N_1561,N_3884);
and U9022 (N_9022,N_3109,N_3035);
or U9023 (N_9023,N_4202,N_2282);
nor U9024 (N_9024,N_4261,N_3672);
and U9025 (N_9025,N_3964,N_646);
nor U9026 (N_9026,N_4706,N_1691);
and U9027 (N_9027,N_1204,N_3940);
nand U9028 (N_9028,N_2777,N_4123);
and U9029 (N_9029,N_487,N_1488);
and U9030 (N_9030,N_4070,N_1895);
nor U9031 (N_9031,N_65,N_4743);
or U9032 (N_9032,N_1133,N_655);
nand U9033 (N_9033,N_3622,N_4670);
nand U9034 (N_9034,N_1256,N_863);
or U9035 (N_9035,N_2632,N_3332);
or U9036 (N_9036,N_4592,N_355);
nand U9037 (N_9037,N_3981,N_3361);
and U9038 (N_9038,N_1004,N_111);
and U9039 (N_9039,N_904,N_1151);
nand U9040 (N_9040,N_4964,N_585);
nand U9041 (N_9041,N_2420,N_3691);
nor U9042 (N_9042,N_1661,N_2894);
nor U9043 (N_9043,N_1886,N_4300);
nor U9044 (N_9044,N_3628,N_3581);
or U9045 (N_9045,N_3710,N_3109);
and U9046 (N_9046,N_4458,N_4622);
nand U9047 (N_9047,N_4739,N_2293);
and U9048 (N_9048,N_460,N_4149);
nand U9049 (N_9049,N_167,N_2881);
nand U9050 (N_9050,N_1731,N_1469);
nor U9051 (N_9051,N_1345,N_1199);
and U9052 (N_9052,N_2979,N_1442);
or U9053 (N_9053,N_1236,N_3409);
or U9054 (N_9054,N_3138,N_3716);
and U9055 (N_9055,N_4087,N_4252);
nand U9056 (N_9056,N_4759,N_2288);
nand U9057 (N_9057,N_138,N_1917);
nor U9058 (N_9058,N_2612,N_1274);
and U9059 (N_9059,N_437,N_4470);
or U9060 (N_9060,N_3394,N_3758);
or U9061 (N_9061,N_4790,N_2854);
or U9062 (N_9062,N_1541,N_4408);
nor U9063 (N_9063,N_200,N_2213);
and U9064 (N_9064,N_2024,N_1675);
nand U9065 (N_9065,N_2115,N_636);
nand U9066 (N_9066,N_4482,N_3247);
nor U9067 (N_9067,N_2214,N_3724);
or U9068 (N_9068,N_1414,N_1339);
nand U9069 (N_9069,N_2541,N_3841);
nand U9070 (N_9070,N_2674,N_1979);
nand U9071 (N_9071,N_4234,N_2217);
or U9072 (N_9072,N_1872,N_1131);
or U9073 (N_9073,N_3549,N_3556);
nand U9074 (N_9074,N_3144,N_1438);
and U9075 (N_9075,N_833,N_1691);
nand U9076 (N_9076,N_1258,N_2422);
or U9077 (N_9077,N_4859,N_1955);
and U9078 (N_9078,N_2754,N_2715);
nor U9079 (N_9079,N_3911,N_4997);
or U9080 (N_9080,N_1540,N_3325);
and U9081 (N_9081,N_3622,N_3798);
nor U9082 (N_9082,N_1465,N_2055);
or U9083 (N_9083,N_1775,N_193);
or U9084 (N_9084,N_1581,N_2464);
nor U9085 (N_9085,N_3812,N_3263);
nand U9086 (N_9086,N_262,N_725);
and U9087 (N_9087,N_3031,N_2325);
or U9088 (N_9088,N_2676,N_2030);
nor U9089 (N_9089,N_4946,N_3494);
or U9090 (N_9090,N_4972,N_3565);
nor U9091 (N_9091,N_2715,N_3584);
xnor U9092 (N_9092,N_2690,N_3111);
nand U9093 (N_9093,N_3304,N_2306);
and U9094 (N_9094,N_4462,N_3313);
and U9095 (N_9095,N_1857,N_967);
nand U9096 (N_9096,N_2931,N_145);
nand U9097 (N_9097,N_1080,N_613);
and U9098 (N_9098,N_2978,N_4756);
nor U9099 (N_9099,N_4465,N_2885);
or U9100 (N_9100,N_2580,N_4158);
and U9101 (N_9101,N_3,N_3820);
or U9102 (N_9102,N_832,N_2882);
nor U9103 (N_9103,N_2782,N_4350);
nor U9104 (N_9104,N_3154,N_313);
nand U9105 (N_9105,N_1883,N_4987);
nor U9106 (N_9106,N_3355,N_2923);
or U9107 (N_9107,N_1519,N_2110);
and U9108 (N_9108,N_544,N_4489);
nor U9109 (N_9109,N_3668,N_4013);
or U9110 (N_9110,N_2604,N_1693);
nor U9111 (N_9111,N_4266,N_4990);
nand U9112 (N_9112,N_352,N_763);
nor U9113 (N_9113,N_1168,N_4630);
nand U9114 (N_9114,N_202,N_3612);
and U9115 (N_9115,N_4222,N_2075);
and U9116 (N_9116,N_1510,N_3614);
or U9117 (N_9117,N_2108,N_2763);
or U9118 (N_9118,N_1991,N_749);
nor U9119 (N_9119,N_137,N_2354);
nor U9120 (N_9120,N_171,N_624);
or U9121 (N_9121,N_691,N_2494);
or U9122 (N_9122,N_4514,N_302);
nand U9123 (N_9123,N_85,N_3206);
and U9124 (N_9124,N_2081,N_4554);
nor U9125 (N_9125,N_954,N_2743);
and U9126 (N_9126,N_1851,N_4190);
xnor U9127 (N_9127,N_1560,N_2607);
nor U9128 (N_9128,N_4765,N_4441);
nor U9129 (N_9129,N_444,N_1923);
nor U9130 (N_9130,N_3442,N_4332);
or U9131 (N_9131,N_2830,N_3628);
and U9132 (N_9132,N_2739,N_572);
nor U9133 (N_9133,N_1557,N_3500);
nor U9134 (N_9134,N_3343,N_4816);
nor U9135 (N_9135,N_1183,N_3070);
or U9136 (N_9136,N_3086,N_4513);
nor U9137 (N_9137,N_1789,N_3863);
and U9138 (N_9138,N_1107,N_512);
and U9139 (N_9139,N_2442,N_4109);
or U9140 (N_9140,N_1500,N_4966);
nor U9141 (N_9141,N_35,N_4135);
nor U9142 (N_9142,N_3489,N_3670);
nor U9143 (N_9143,N_594,N_1858);
or U9144 (N_9144,N_2296,N_1912);
nor U9145 (N_9145,N_3673,N_852);
nand U9146 (N_9146,N_3753,N_3648);
xnor U9147 (N_9147,N_3607,N_3452);
nor U9148 (N_9148,N_661,N_3353);
nor U9149 (N_9149,N_3629,N_4000);
nand U9150 (N_9150,N_4644,N_1700);
or U9151 (N_9151,N_645,N_1330);
and U9152 (N_9152,N_2560,N_3687);
nor U9153 (N_9153,N_977,N_1644);
nand U9154 (N_9154,N_1587,N_1244);
or U9155 (N_9155,N_3998,N_2583);
or U9156 (N_9156,N_1705,N_2219);
nor U9157 (N_9157,N_3190,N_231);
nor U9158 (N_9158,N_2228,N_4215);
nand U9159 (N_9159,N_2937,N_2266);
and U9160 (N_9160,N_1188,N_3914);
and U9161 (N_9161,N_2193,N_752);
and U9162 (N_9162,N_4681,N_3057);
and U9163 (N_9163,N_594,N_606);
nor U9164 (N_9164,N_4674,N_1137);
nand U9165 (N_9165,N_2939,N_2075);
nand U9166 (N_9166,N_3494,N_3680);
nor U9167 (N_9167,N_2858,N_4301);
nor U9168 (N_9168,N_403,N_4340);
and U9169 (N_9169,N_3442,N_2800);
nand U9170 (N_9170,N_819,N_4289);
and U9171 (N_9171,N_3979,N_4033);
and U9172 (N_9172,N_3966,N_3086);
nand U9173 (N_9173,N_2587,N_84);
nand U9174 (N_9174,N_2930,N_4428);
nand U9175 (N_9175,N_1249,N_2495);
and U9176 (N_9176,N_2039,N_2193);
and U9177 (N_9177,N_2424,N_893);
and U9178 (N_9178,N_2649,N_3551);
or U9179 (N_9179,N_734,N_1992);
nand U9180 (N_9180,N_1219,N_143);
or U9181 (N_9181,N_2616,N_918);
nand U9182 (N_9182,N_3297,N_348);
nor U9183 (N_9183,N_3747,N_4310);
or U9184 (N_9184,N_3920,N_779);
nand U9185 (N_9185,N_2171,N_3772);
nand U9186 (N_9186,N_859,N_2777);
and U9187 (N_9187,N_3936,N_2760);
nor U9188 (N_9188,N_3182,N_942);
and U9189 (N_9189,N_3608,N_664);
nand U9190 (N_9190,N_1301,N_4442);
nand U9191 (N_9191,N_4076,N_3782);
nand U9192 (N_9192,N_3309,N_4720);
or U9193 (N_9193,N_3193,N_3917);
nand U9194 (N_9194,N_3026,N_3213);
and U9195 (N_9195,N_1409,N_4385);
and U9196 (N_9196,N_3876,N_2572);
or U9197 (N_9197,N_3620,N_4489);
and U9198 (N_9198,N_498,N_2661);
and U9199 (N_9199,N_2262,N_799);
and U9200 (N_9200,N_482,N_4110);
and U9201 (N_9201,N_3624,N_3354);
nand U9202 (N_9202,N_4165,N_3094);
and U9203 (N_9203,N_147,N_3818);
nand U9204 (N_9204,N_4894,N_2765);
or U9205 (N_9205,N_4172,N_3059);
nor U9206 (N_9206,N_4038,N_1151);
nand U9207 (N_9207,N_2337,N_4679);
nor U9208 (N_9208,N_3294,N_806);
nor U9209 (N_9209,N_3591,N_3673);
nor U9210 (N_9210,N_1189,N_1835);
or U9211 (N_9211,N_3309,N_3022);
nand U9212 (N_9212,N_399,N_855);
or U9213 (N_9213,N_4091,N_1955);
nor U9214 (N_9214,N_280,N_2176);
or U9215 (N_9215,N_256,N_1550);
and U9216 (N_9216,N_1572,N_1848);
nor U9217 (N_9217,N_3799,N_2935);
or U9218 (N_9218,N_2569,N_4186);
nand U9219 (N_9219,N_1786,N_2279);
or U9220 (N_9220,N_57,N_4140);
nand U9221 (N_9221,N_3085,N_4352);
or U9222 (N_9222,N_1821,N_725);
or U9223 (N_9223,N_1290,N_1989);
or U9224 (N_9224,N_4709,N_2954);
nor U9225 (N_9225,N_1079,N_3802);
nand U9226 (N_9226,N_1087,N_377);
nor U9227 (N_9227,N_1988,N_2517);
nor U9228 (N_9228,N_2523,N_2639);
or U9229 (N_9229,N_3554,N_3560);
or U9230 (N_9230,N_3897,N_3007);
and U9231 (N_9231,N_2480,N_3104);
or U9232 (N_9232,N_1601,N_683);
nor U9233 (N_9233,N_2787,N_4508);
and U9234 (N_9234,N_394,N_1809);
nor U9235 (N_9235,N_4369,N_4103);
nor U9236 (N_9236,N_4813,N_4763);
or U9237 (N_9237,N_4565,N_2868);
nor U9238 (N_9238,N_824,N_3910);
or U9239 (N_9239,N_2904,N_1829);
nor U9240 (N_9240,N_2432,N_1305);
nor U9241 (N_9241,N_954,N_3918);
nand U9242 (N_9242,N_1020,N_826);
nor U9243 (N_9243,N_1249,N_618);
nor U9244 (N_9244,N_1474,N_1224);
nor U9245 (N_9245,N_4355,N_1603);
nor U9246 (N_9246,N_870,N_2086);
or U9247 (N_9247,N_901,N_50);
and U9248 (N_9248,N_718,N_3771);
or U9249 (N_9249,N_4592,N_2360);
nand U9250 (N_9250,N_1368,N_4053);
nand U9251 (N_9251,N_1906,N_3210);
or U9252 (N_9252,N_1229,N_4684);
nand U9253 (N_9253,N_2766,N_4883);
and U9254 (N_9254,N_117,N_2783);
nand U9255 (N_9255,N_432,N_3816);
nor U9256 (N_9256,N_3083,N_3521);
or U9257 (N_9257,N_4926,N_1937);
nand U9258 (N_9258,N_1120,N_4768);
or U9259 (N_9259,N_1188,N_771);
or U9260 (N_9260,N_2410,N_3703);
nor U9261 (N_9261,N_86,N_2382);
nor U9262 (N_9262,N_4763,N_2779);
or U9263 (N_9263,N_4129,N_4187);
or U9264 (N_9264,N_3323,N_1679);
and U9265 (N_9265,N_4097,N_1621);
nor U9266 (N_9266,N_4701,N_4886);
or U9267 (N_9267,N_4273,N_4660);
nand U9268 (N_9268,N_2058,N_4346);
nor U9269 (N_9269,N_4336,N_1803);
nand U9270 (N_9270,N_2427,N_3156);
nor U9271 (N_9271,N_612,N_2935);
and U9272 (N_9272,N_870,N_2867);
nor U9273 (N_9273,N_536,N_4722);
nand U9274 (N_9274,N_1569,N_4490);
xor U9275 (N_9275,N_4183,N_1142);
or U9276 (N_9276,N_4322,N_162);
and U9277 (N_9277,N_3931,N_3034);
nor U9278 (N_9278,N_2715,N_840);
nand U9279 (N_9279,N_1816,N_3068);
or U9280 (N_9280,N_3507,N_4495);
and U9281 (N_9281,N_3678,N_3878);
nor U9282 (N_9282,N_3921,N_2454);
or U9283 (N_9283,N_4585,N_4798);
nor U9284 (N_9284,N_1491,N_416);
nor U9285 (N_9285,N_2072,N_1601);
or U9286 (N_9286,N_13,N_1178);
nand U9287 (N_9287,N_1398,N_1088);
or U9288 (N_9288,N_2652,N_916);
nand U9289 (N_9289,N_3000,N_2051);
or U9290 (N_9290,N_1391,N_4972);
or U9291 (N_9291,N_2834,N_2688);
or U9292 (N_9292,N_2147,N_3846);
and U9293 (N_9293,N_1391,N_4850);
nor U9294 (N_9294,N_3636,N_4927);
or U9295 (N_9295,N_4710,N_2689);
and U9296 (N_9296,N_882,N_1662);
nand U9297 (N_9297,N_4608,N_710);
and U9298 (N_9298,N_304,N_550);
and U9299 (N_9299,N_779,N_2600);
nor U9300 (N_9300,N_3949,N_1925);
nor U9301 (N_9301,N_2525,N_1570);
and U9302 (N_9302,N_1167,N_3017);
and U9303 (N_9303,N_3077,N_1747);
or U9304 (N_9304,N_1021,N_3374);
or U9305 (N_9305,N_53,N_4499);
nor U9306 (N_9306,N_2864,N_3890);
xor U9307 (N_9307,N_1023,N_3220);
nor U9308 (N_9308,N_972,N_3104);
nor U9309 (N_9309,N_2278,N_3522);
and U9310 (N_9310,N_1055,N_4979);
and U9311 (N_9311,N_1844,N_504);
nor U9312 (N_9312,N_3484,N_2530);
nor U9313 (N_9313,N_3749,N_1978);
and U9314 (N_9314,N_2674,N_2043);
and U9315 (N_9315,N_4344,N_3553);
xnor U9316 (N_9316,N_655,N_1122);
and U9317 (N_9317,N_16,N_1279);
or U9318 (N_9318,N_2943,N_44);
nor U9319 (N_9319,N_3086,N_1130);
or U9320 (N_9320,N_3519,N_1719);
or U9321 (N_9321,N_1954,N_2985);
nor U9322 (N_9322,N_4811,N_3111);
nor U9323 (N_9323,N_3219,N_139);
and U9324 (N_9324,N_3811,N_2863);
nand U9325 (N_9325,N_3148,N_2362);
nand U9326 (N_9326,N_65,N_2295);
or U9327 (N_9327,N_525,N_1163);
or U9328 (N_9328,N_451,N_1257);
nand U9329 (N_9329,N_2810,N_4641);
nor U9330 (N_9330,N_3208,N_1766);
and U9331 (N_9331,N_4687,N_4265);
or U9332 (N_9332,N_899,N_2553);
and U9333 (N_9333,N_4423,N_3184);
nand U9334 (N_9334,N_3990,N_515);
nand U9335 (N_9335,N_4836,N_3386);
nand U9336 (N_9336,N_1030,N_1426);
xor U9337 (N_9337,N_3220,N_1984);
or U9338 (N_9338,N_4894,N_4191);
nand U9339 (N_9339,N_3934,N_2177);
nor U9340 (N_9340,N_3824,N_499);
nor U9341 (N_9341,N_837,N_1241);
or U9342 (N_9342,N_1739,N_2162);
or U9343 (N_9343,N_4066,N_4443);
nand U9344 (N_9344,N_1174,N_2877);
nor U9345 (N_9345,N_2578,N_3279);
and U9346 (N_9346,N_2259,N_1360);
and U9347 (N_9347,N_4238,N_79);
nand U9348 (N_9348,N_4230,N_4560);
and U9349 (N_9349,N_1550,N_445);
or U9350 (N_9350,N_3450,N_463);
nor U9351 (N_9351,N_1663,N_4683);
and U9352 (N_9352,N_2100,N_3091);
nor U9353 (N_9353,N_1245,N_815);
and U9354 (N_9354,N_2985,N_2468);
and U9355 (N_9355,N_643,N_4069);
and U9356 (N_9356,N_1016,N_304);
or U9357 (N_9357,N_1828,N_3785);
nor U9358 (N_9358,N_2990,N_2871);
and U9359 (N_9359,N_4623,N_99);
nor U9360 (N_9360,N_636,N_3780);
and U9361 (N_9361,N_3379,N_4922);
nand U9362 (N_9362,N_2872,N_4081);
nand U9363 (N_9363,N_3754,N_553);
nand U9364 (N_9364,N_1035,N_2741);
nand U9365 (N_9365,N_3406,N_16);
or U9366 (N_9366,N_1691,N_1411);
nand U9367 (N_9367,N_2749,N_3009);
or U9368 (N_9368,N_3529,N_603);
and U9369 (N_9369,N_4100,N_3794);
and U9370 (N_9370,N_3908,N_2579);
nand U9371 (N_9371,N_2096,N_579);
and U9372 (N_9372,N_1033,N_3935);
or U9373 (N_9373,N_2631,N_795);
or U9374 (N_9374,N_1385,N_1573);
nand U9375 (N_9375,N_4146,N_1325);
and U9376 (N_9376,N_646,N_3427);
or U9377 (N_9377,N_3818,N_1868);
nand U9378 (N_9378,N_2015,N_3084);
nand U9379 (N_9379,N_891,N_3757);
nand U9380 (N_9380,N_667,N_3244);
and U9381 (N_9381,N_2355,N_2766);
nand U9382 (N_9382,N_1162,N_4698);
nor U9383 (N_9383,N_2040,N_4159);
and U9384 (N_9384,N_3931,N_351);
nor U9385 (N_9385,N_141,N_372);
or U9386 (N_9386,N_2901,N_1802);
nand U9387 (N_9387,N_2599,N_1023);
nand U9388 (N_9388,N_796,N_2940);
nor U9389 (N_9389,N_1469,N_3552);
or U9390 (N_9390,N_3415,N_1320);
and U9391 (N_9391,N_878,N_3929);
and U9392 (N_9392,N_761,N_126);
nand U9393 (N_9393,N_4798,N_1577);
xor U9394 (N_9394,N_2204,N_596);
or U9395 (N_9395,N_3600,N_678);
nand U9396 (N_9396,N_449,N_920);
and U9397 (N_9397,N_108,N_2104);
or U9398 (N_9398,N_3058,N_3021);
and U9399 (N_9399,N_4147,N_4308);
nor U9400 (N_9400,N_354,N_1144);
xnor U9401 (N_9401,N_637,N_1915);
and U9402 (N_9402,N_2982,N_387);
nand U9403 (N_9403,N_4217,N_4328);
and U9404 (N_9404,N_3016,N_996);
nor U9405 (N_9405,N_4621,N_1652);
or U9406 (N_9406,N_4582,N_85);
and U9407 (N_9407,N_3407,N_3054);
and U9408 (N_9408,N_460,N_4675);
or U9409 (N_9409,N_2596,N_1364);
and U9410 (N_9410,N_2260,N_4879);
and U9411 (N_9411,N_4315,N_2817);
nor U9412 (N_9412,N_4708,N_3871);
nor U9413 (N_9413,N_548,N_3481);
or U9414 (N_9414,N_1216,N_1000);
nor U9415 (N_9415,N_4790,N_499);
or U9416 (N_9416,N_2598,N_2273);
or U9417 (N_9417,N_3440,N_4720);
or U9418 (N_9418,N_1249,N_1530);
and U9419 (N_9419,N_220,N_4483);
and U9420 (N_9420,N_4490,N_3499);
nand U9421 (N_9421,N_1953,N_203);
and U9422 (N_9422,N_4570,N_1507);
or U9423 (N_9423,N_1951,N_4003);
nand U9424 (N_9424,N_117,N_549);
nand U9425 (N_9425,N_1386,N_4495);
nand U9426 (N_9426,N_2805,N_2305);
and U9427 (N_9427,N_3968,N_4993);
nor U9428 (N_9428,N_1603,N_1848);
nor U9429 (N_9429,N_2646,N_658);
nor U9430 (N_9430,N_4319,N_318);
nand U9431 (N_9431,N_1653,N_4);
nor U9432 (N_9432,N_1085,N_3147);
nand U9433 (N_9433,N_1949,N_1880);
nor U9434 (N_9434,N_2682,N_3067);
xnor U9435 (N_9435,N_3541,N_3661);
and U9436 (N_9436,N_3268,N_4539);
and U9437 (N_9437,N_3133,N_1468);
or U9438 (N_9438,N_4263,N_2128);
or U9439 (N_9439,N_3840,N_818);
and U9440 (N_9440,N_2368,N_4139);
nand U9441 (N_9441,N_3400,N_3818);
nor U9442 (N_9442,N_4499,N_1450);
nor U9443 (N_9443,N_945,N_3203);
nand U9444 (N_9444,N_2267,N_2887);
nor U9445 (N_9445,N_2178,N_926);
and U9446 (N_9446,N_1118,N_4505);
and U9447 (N_9447,N_2901,N_3072);
nand U9448 (N_9448,N_1719,N_2116);
and U9449 (N_9449,N_2616,N_3924);
nand U9450 (N_9450,N_4639,N_4945);
nor U9451 (N_9451,N_4480,N_1683);
and U9452 (N_9452,N_3017,N_106);
xnor U9453 (N_9453,N_1371,N_2017);
or U9454 (N_9454,N_3943,N_4901);
or U9455 (N_9455,N_3509,N_2947);
xor U9456 (N_9456,N_3068,N_1368);
nor U9457 (N_9457,N_268,N_3102);
or U9458 (N_9458,N_3133,N_2604);
xor U9459 (N_9459,N_547,N_4795);
and U9460 (N_9460,N_369,N_2440);
nand U9461 (N_9461,N_2234,N_3143);
or U9462 (N_9462,N_2642,N_1053);
and U9463 (N_9463,N_4283,N_2424);
nor U9464 (N_9464,N_549,N_2726);
nand U9465 (N_9465,N_3101,N_3482);
and U9466 (N_9466,N_3594,N_269);
or U9467 (N_9467,N_3117,N_901);
nor U9468 (N_9468,N_2203,N_1549);
xnor U9469 (N_9469,N_4231,N_3632);
or U9470 (N_9470,N_1833,N_714);
or U9471 (N_9471,N_4722,N_2999);
and U9472 (N_9472,N_1152,N_3064);
and U9473 (N_9473,N_331,N_1876);
or U9474 (N_9474,N_410,N_2959);
nand U9475 (N_9475,N_2994,N_2257);
or U9476 (N_9476,N_2637,N_1013);
and U9477 (N_9477,N_581,N_3499);
nor U9478 (N_9478,N_3333,N_3209);
nand U9479 (N_9479,N_3810,N_4285);
nor U9480 (N_9480,N_2,N_3275);
or U9481 (N_9481,N_1392,N_4856);
or U9482 (N_9482,N_2545,N_4596);
xnor U9483 (N_9483,N_3785,N_1999);
and U9484 (N_9484,N_2146,N_1237);
xnor U9485 (N_9485,N_3504,N_4169);
nor U9486 (N_9486,N_1532,N_179);
nor U9487 (N_9487,N_1753,N_4975);
nor U9488 (N_9488,N_359,N_984);
nand U9489 (N_9489,N_3934,N_3482);
nor U9490 (N_9490,N_4941,N_462);
or U9491 (N_9491,N_3578,N_3904);
and U9492 (N_9492,N_2790,N_1672);
nand U9493 (N_9493,N_1855,N_1979);
and U9494 (N_9494,N_2248,N_4433);
nand U9495 (N_9495,N_2463,N_957);
or U9496 (N_9496,N_784,N_3015);
and U9497 (N_9497,N_862,N_2414);
nand U9498 (N_9498,N_1637,N_1556);
nor U9499 (N_9499,N_2629,N_2410);
and U9500 (N_9500,N_4190,N_4327);
xor U9501 (N_9501,N_1790,N_786);
nand U9502 (N_9502,N_1704,N_1305);
nor U9503 (N_9503,N_654,N_1487);
or U9504 (N_9504,N_2488,N_442);
and U9505 (N_9505,N_1195,N_4340);
or U9506 (N_9506,N_802,N_4964);
nor U9507 (N_9507,N_1005,N_3228);
and U9508 (N_9508,N_3985,N_3429);
or U9509 (N_9509,N_2846,N_1409);
and U9510 (N_9510,N_151,N_3717);
or U9511 (N_9511,N_2817,N_318);
and U9512 (N_9512,N_3856,N_4174);
or U9513 (N_9513,N_2662,N_1828);
and U9514 (N_9514,N_2889,N_1472);
and U9515 (N_9515,N_175,N_4620);
nor U9516 (N_9516,N_67,N_773);
nor U9517 (N_9517,N_916,N_3112);
or U9518 (N_9518,N_3204,N_4835);
and U9519 (N_9519,N_904,N_3320);
nand U9520 (N_9520,N_2613,N_370);
or U9521 (N_9521,N_195,N_2052);
nor U9522 (N_9522,N_4150,N_180);
nand U9523 (N_9523,N_3167,N_2681);
and U9524 (N_9524,N_870,N_3739);
and U9525 (N_9525,N_378,N_4895);
or U9526 (N_9526,N_4747,N_3719);
nand U9527 (N_9527,N_3988,N_1150);
or U9528 (N_9528,N_2887,N_640);
and U9529 (N_9529,N_3302,N_3372);
nand U9530 (N_9530,N_4466,N_558);
nor U9531 (N_9531,N_4495,N_2379);
nor U9532 (N_9532,N_1160,N_2537);
nand U9533 (N_9533,N_4065,N_1379);
and U9534 (N_9534,N_2587,N_1390);
or U9535 (N_9535,N_246,N_1338);
nor U9536 (N_9536,N_2738,N_4494);
or U9537 (N_9537,N_1003,N_2196);
and U9538 (N_9538,N_2071,N_4655);
nor U9539 (N_9539,N_3548,N_4948);
or U9540 (N_9540,N_2801,N_2027);
or U9541 (N_9541,N_4647,N_3884);
nand U9542 (N_9542,N_3125,N_446);
and U9543 (N_9543,N_4022,N_2776);
nand U9544 (N_9544,N_2166,N_4845);
nor U9545 (N_9545,N_4374,N_4389);
or U9546 (N_9546,N_2027,N_3651);
or U9547 (N_9547,N_3679,N_1732);
or U9548 (N_9548,N_3901,N_1180);
or U9549 (N_9549,N_2817,N_1388);
or U9550 (N_9550,N_3217,N_1141);
and U9551 (N_9551,N_238,N_4018);
nor U9552 (N_9552,N_4724,N_2529);
and U9553 (N_9553,N_4860,N_600);
or U9554 (N_9554,N_2559,N_4214);
nor U9555 (N_9555,N_64,N_1622);
nand U9556 (N_9556,N_4952,N_4299);
or U9557 (N_9557,N_1051,N_3842);
nand U9558 (N_9558,N_138,N_1549);
nand U9559 (N_9559,N_4514,N_3602);
and U9560 (N_9560,N_2697,N_3278);
or U9561 (N_9561,N_4958,N_1331);
nor U9562 (N_9562,N_4348,N_3427);
nand U9563 (N_9563,N_1117,N_4460);
or U9564 (N_9564,N_1600,N_4032);
nand U9565 (N_9565,N_113,N_799);
nand U9566 (N_9566,N_1160,N_1337);
nor U9567 (N_9567,N_4846,N_3762);
and U9568 (N_9568,N_4549,N_4707);
or U9569 (N_9569,N_215,N_440);
or U9570 (N_9570,N_1427,N_1760);
or U9571 (N_9571,N_4278,N_517);
or U9572 (N_9572,N_3253,N_2627);
nor U9573 (N_9573,N_1185,N_3084);
nand U9574 (N_9574,N_1473,N_2574);
and U9575 (N_9575,N_1469,N_4263);
nand U9576 (N_9576,N_1979,N_4664);
nor U9577 (N_9577,N_1760,N_3647);
and U9578 (N_9578,N_1821,N_3725);
nand U9579 (N_9579,N_3209,N_2077);
nand U9580 (N_9580,N_4183,N_2316);
nand U9581 (N_9581,N_1050,N_693);
or U9582 (N_9582,N_2450,N_1473);
nand U9583 (N_9583,N_2045,N_1523);
nor U9584 (N_9584,N_44,N_1009);
nand U9585 (N_9585,N_320,N_4836);
nor U9586 (N_9586,N_2576,N_308);
nor U9587 (N_9587,N_4864,N_2350);
nand U9588 (N_9588,N_785,N_1387);
nor U9589 (N_9589,N_1900,N_463);
or U9590 (N_9590,N_1107,N_3683);
nand U9591 (N_9591,N_682,N_110);
and U9592 (N_9592,N_4666,N_230);
nor U9593 (N_9593,N_2296,N_2682);
nor U9594 (N_9594,N_3626,N_4991);
nand U9595 (N_9595,N_4430,N_4252);
nor U9596 (N_9596,N_4367,N_4936);
nor U9597 (N_9597,N_4326,N_3571);
nor U9598 (N_9598,N_2976,N_1451);
nand U9599 (N_9599,N_3569,N_3752);
nor U9600 (N_9600,N_2204,N_733);
or U9601 (N_9601,N_3962,N_1277);
or U9602 (N_9602,N_4799,N_3624);
nor U9603 (N_9603,N_3749,N_2797);
or U9604 (N_9604,N_4934,N_1930);
nand U9605 (N_9605,N_1022,N_871);
and U9606 (N_9606,N_823,N_2860);
or U9607 (N_9607,N_4862,N_989);
or U9608 (N_9608,N_2508,N_4341);
nand U9609 (N_9609,N_2590,N_2230);
and U9610 (N_9610,N_135,N_3294);
or U9611 (N_9611,N_1448,N_2070);
nand U9612 (N_9612,N_577,N_2925);
nand U9613 (N_9613,N_1090,N_4072);
and U9614 (N_9614,N_2795,N_1346);
nor U9615 (N_9615,N_1634,N_3735);
and U9616 (N_9616,N_2083,N_996);
or U9617 (N_9617,N_2721,N_656);
nand U9618 (N_9618,N_1869,N_4466);
or U9619 (N_9619,N_484,N_1999);
and U9620 (N_9620,N_867,N_1330);
nor U9621 (N_9621,N_1351,N_1662);
or U9622 (N_9622,N_336,N_224);
nand U9623 (N_9623,N_3883,N_1781);
and U9624 (N_9624,N_371,N_3273);
nand U9625 (N_9625,N_240,N_28);
and U9626 (N_9626,N_778,N_2833);
nand U9627 (N_9627,N_438,N_316);
and U9628 (N_9628,N_4739,N_3904);
or U9629 (N_9629,N_841,N_471);
nor U9630 (N_9630,N_1962,N_1923);
or U9631 (N_9631,N_4843,N_2549);
nand U9632 (N_9632,N_1546,N_656);
or U9633 (N_9633,N_2939,N_2424);
and U9634 (N_9634,N_2219,N_279);
or U9635 (N_9635,N_3966,N_3850);
or U9636 (N_9636,N_3330,N_2701);
nor U9637 (N_9637,N_4054,N_4718);
nor U9638 (N_9638,N_1865,N_3733);
nand U9639 (N_9639,N_1018,N_3827);
nor U9640 (N_9640,N_4874,N_2273);
nand U9641 (N_9641,N_2617,N_202);
or U9642 (N_9642,N_4797,N_3408);
nor U9643 (N_9643,N_448,N_2818);
and U9644 (N_9644,N_2077,N_978);
or U9645 (N_9645,N_545,N_931);
nor U9646 (N_9646,N_2371,N_2260);
or U9647 (N_9647,N_4732,N_1205);
or U9648 (N_9648,N_1801,N_4425);
nor U9649 (N_9649,N_2294,N_2458);
or U9650 (N_9650,N_3603,N_130);
or U9651 (N_9651,N_1498,N_4544);
nand U9652 (N_9652,N_3841,N_2611);
or U9653 (N_9653,N_1846,N_428);
or U9654 (N_9654,N_1398,N_1453);
nor U9655 (N_9655,N_3869,N_82);
and U9656 (N_9656,N_4823,N_4638);
nand U9657 (N_9657,N_3952,N_566);
and U9658 (N_9658,N_3087,N_3540);
and U9659 (N_9659,N_2383,N_3503);
nor U9660 (N_9660,N_3900,N_656);
nor U9661 (N_9661,N_3096,N_336);
nand U9662 (N_9662,N_711,N_445);
or U9663 (N_9663,N_1161,N_2881);
and U9664 (N_9664,N_3837,N_2844);
or U9665 (N_9665,N_3830,N_4315);
xnor U9666 (N_9666,N_1073,N_993);
and U9667 (N_9667,N_1067,N_397);
or U9668 (N_9668,N_1658,N_4379);
and U9669 (N_9669,N_1293,N_3793);
and U9670 (N_9670,N_2803,N_57);
and U9671 (N_9671,N_2491,N_2366);
nand U9672 (N_9672,N_3398,N_3909);
and U9673 (N_9673,N_3446,N_4077);
or U9674 (N_9674,N_3194,N_2446);
or U9675 (N_9675,N_953,N_2160);
nand U9676 (N_9676,N_4404,N_1096);
or U9677 (N_9677,N_3566,N_2056);
nor U9678 (N_9678,N_1633,N_2610);
nor U9679 (N_9679,N_2080,N_4201);
nand U9680 (N_9680,N_4654,N_65);
xor U9681 (N_9681,N_3643,N_207);
nor U9682 (N_9682,N_2741,N_2622);
nor U9683 (N_9683,N_3359,N_3764);
nand U9684 (N_9684,N_104,N_977);
and U9685 (N_9685,N_1523,N_2256);
nand U9686 (N_9686,N_811,N_1992);
nor U9687 (N_9687,N_725,N_715);
nand U9688 (N_9688,N_2494,N_1937);
and U9689 (N_9689,N_1463,N_3353);
nor U9690 (N_9690,N_4920,N_837);
nor U9691 (N_9691,N_2700,N_4150);
and U9692 (N_9692,N_2294,N_1045);
and U9693 (N_9693,N_688,N_396);
nor U9694 (N_9694,N_3234,N_2220);
or U9695 (N_9695,N_1586,N_199);
or U9696 (N_9696,N_4223,N_4318);
or U9697 (N_9697,N_874,N_2668);
or U9698 (N_9698,N_1716,N_4291);
nand U9699 (N_9699,N_3090,N_1979);
nor U9700 (N_9700,N_1240,N_2454);
and U9701 (N_9701,N_365,N_195);
nor U9702 (N_9702,N_1156,N_1386);
xor U9703 (N_9703,N_2278,N_4137);
or U9704 (N_9704,N_1506,N_616);
nand U9705 (N_9705,N_2573,N_1943);
nor U9706 (N_9706,N_1521,N_4477);
nor U9707 (N_9707,N_2904,N_1933);
nand U9708 (N_9708,N_4595,N_16);
nor U9709 (N_9709,N_4798,N_571);
nand U9710 (N_9710,N_4753,N_2645);
or U9711 (N_9711,N_1865,N_2444);
nor U9712 (N_9712,N_3587,N_4981);
or U9713 (N_9713,N_4893,N_4605);
and U9714 (N_9714,N_1027,N_896);
nor U9715 (N_9715,N_4572,N_2567);
and U9716 (N_9716,N_4038,N_3350);
nand U9717 (N_9717,N_197,N_2152);
or U9718 (N_9718,N_4476,N_1517);
or U9719 (N_9719,N_498,N_256);
nor U9720 (N_9720,N_3737,N_1555);
nor U9721 (N_9721,N_139,N_2175);
nand U9722 (N_9722,N_1818,N_451);
nand U9723 (N_9723,N_323,N_4627);
or U9724 (N_9724,N_4875,N_3783);
nand U9725 (N_9725,N_3249,N_1206);
nor U9726 (N_9726,N_2434,N_37);
nand U9727 (N_9727,N_2816,N_3045);
nor U9728 (N_9728,N_1161,N_1011);
nor U9729 (N_9729,N_2549,N_3977);
nor U9730 (N_9730,N_999,N_2186);
and U9731 (N_9731,N_3572,N_1618);
nand U9732 (N_9732,N_2333,N_3882);
or U9733 (N_9733,N_3473,N_2225);
nor U9734 (N_9734,N_2645,N_1537);
nor U9735 (N_9735,N_3607,N_3771);
and U9736 (N_9736,N_4464,N_1066);
nor U9737 (N_9737,N_4495,N_2721);
nor U9738 (N_9738,N_1203,N_3474);
nand U9739 (N_9739,N_3402,N_3777);
nor U9740 (N_9740,N_4586,N_2151);
or U9741 (N_9741,N_3547,N_1122);
nor U9742 (N_9742,N_3620,N_2104);
nand U9743 (N_9743,N_3293,N_3077);
and U9744 (N_9744,N_4244,N_1970);
nor U9745 (N_9745,N_1116,N_1420);
and U9746 (N_9746,N_1076,N_944);
nand U9747 (N_9747,N_708,N_4820);
nand U9748 (N_9748,N_1061,N_1652);
and U9749 (N_9749,N_129,N_3340);
nand U9750 (N_9750,N_3392,N_4269);
or U9751 (N_9751,N_4439,N_3552);
or U9752 (N_9752,N_4959,N_985);
nand U9753 (N_9753,N_605,N_1991);
nand U9754 (N_9754,N_772,N_4522);
or U9755 (N_9755,N_1271,N_4536);
nand U9756 (N_9756,N_2703,N_3922);
nor U9757 (N_9757,N_878,N_2321);
nor U9758 (N_9758,N_4552,N_4868);
or U9759 (N_9759,N_4963,N_3721);
or U9760 (N_9760,N_730,N_3097);
and U9761 (N_9761,N_622,N_59);
nor U9762 (N_9762,N_1328,N_248);
nor U9763 (N_9763,N_2646,N_1843);
nor U9764 (N_9764,N_1485,N_2040);
nor U9765 (N_9765,N_1262,N_3538);
and U9766 (N_9766,N_49,N_3311);
nand U9767 (N_9767,N_4937,N_3226);
and U9768 (N_9768,N_166,N_3027);
or U9769 (N_9769,N_3903,N_2153);
nand U9770 (N_9770,N_283,N_3624);
xnor U9771 (N_9771,N_4364,N_1427);
nand U9772 (N_9772,N_1305,N_3130);
nand U9773 (N_9773,N_4418,N_1022);
and U9774 (N_9774,N_4527,N_1083);
nor U9775 (N_9775,N_4138,N_2371);
nor U9776 (N_9776,N_2861,N_1880);
nor U9777 (N_9777,N_4892,N_3995);
and U9778 (N_9778,N_4748,N_4517);
and U9779 (N_9779,N_50,N_174);
nor U9780 (N_9780,N_198,N_3135);
and U9781 (N_9781,N_4392,N_987);
or U9782 (N_9782,N_2155,N_3509);
and U9783 (N_9783,N_2030,N_1347);
or U9784 (N_9784,N_1902,N_2212);
nand U9785 (N_9785,N_4523,N_2460);
and U9786 (N_9786,N_920,N_621);
and U9787 (N_9787,N_4399,N_1934);
or U9788 (N_9788,N_1087,N_4121);
nand U9789 (N_9789,N_3360,N_4689);
or U9790 (N_9790,N_4575,N_4868);
nand U9791 (N_9791,N_4577,N_4084);
and U9792 (N_9792,N_3471,N_4723);
and U9793 (N_9793,N_4811,N_584);
nor U9794 (N_9794,N_3206,N_1670);
nor U9795 (N_9795,N_1778,N_2274);
and U9796 (N_9796,N_4607,N_1635);
or U9797 (N_9797,N_4716,N_203);
or U9798 (N_9798,N_3173,N_4848);
or U9799 (N_9799,N_4962,N_4390);
nand U9800 (N_9800,N_814,N_4478);
nand U9801 (N_9801,N_3139,N_3008);
and U9802 (N_9802,N_4931,N_3260);
and U9803 (N_9803,N_4822,N_587);
xnor U9804 (N_9804,N_2516,N_1933);
nor U9805 (N_9805,N_2771,N_322);
xor U9806 (N_9806,N_2725,N_2569);
and U9807 (N_9807,N_2144,N_1875);
and U9808 (N_9808,N_813,N_647);
nor U9809 (N_9809,N_4178,N_4133);
or U9810 (N_9810,N_2462,N_775);
nor U9811 (N_9811,N_3236,N_2420);
nor U9812 (N_9812,N_3363,N_1074);
nand U9813 (N_9813,N_800,N_3175);
nor U9814 (N_9814,N_4123,N_4465);
nand U9815 (N_9815,N_4413,N_4927);
nand U9816 (N_9816,N_840,N_1344);
nand U9817 (N_9817,N_3871,N_1236);
nor U9818 (N_9818,N_2824,N_2884);
nor U9819 (N_9819,N_4472,N_4711);
nor U9820 (N_9820,N_3687,N_3401);
nand U9821 (N_9821,N_3896,N_3999);
or U9822 (N_9822,N_2126,N_1569);
nor U9823 (N_9823,N_3702,N_4368);
or U9824 (N_9824,N_1913,N_4137);
or U9825 (N_9825,N_4558,N_3766);
nor U9826 (N_9826,N_174,N_658);
or U9827 (N_9827,N_627,N_4550);
nand U9828 (N_9828,N_378,N_3608);
nand U9829 (N_9829,N_520,N_4529);
or U9830 (N_9830,N_1213,N_4442);
or U9831 (N_9831,N_2902,N_1947);
or U9832 (N_9832,N_3173,N_3786);
nor U9833 (N_9833,N_2777,N_597);
or U9834 (N_9834,N_4917,N_4983);
xnor U9835 (N_9835,N_3104,N_4592);
or U9836 (N_9836,N_4235,N_486);
and U9837 (N_9837,N_1610,N_2253);
nand U9838 (N_9838,N_3186,N_3734);
nand U9839 (N_9839,N_4112,N_1981);
and U9840 (N_9840,N_3485,N_4948);
or U9841 (N_9841,N_3287,N_2272);
or U9842 (N_9842,N_4793,N_1794);
or U9843 (N_9843,N_1924,N_4651);
nor U9844 (N_9844,N_684,N_3162);
xor U9845 (N_9845,N_1569,N_3466);
or U9846 (N_9846,N_676,N_3003);
and U9847 (N_9847,N_284,N_784);
nand U9848 (N_9848,N_3874,N_3942);
nor U9849 (N_9849,N_2329,N_4778);
and U9850 (N_9850,N_1960,N_1204);
and U9851 (N_9851,N_872,N_2916);
and U9852 (N_9852,N_3928,N_2055);
nor U9853 (N_9853,N_4104,N_1478);
nand U9854 (N_9854,N_3788,N_938);
or U9855 (N_9855,N_3610,N_3835);
and U9856 (N_9856,N_4840,N_544);
or U9857 (N_9857,N_2988,N_4316);
or U9858 (N_9858,N_2711,N_871);
nand U9859 (N_9859,N_2800,N_4446);
and U9860 (N_9860,N_685,N_1026);
or U9861 (N_9861,N_991,N_757);
and U9862 (N_9862,N_4751,N_804);
nor U9863 (N_9863,N_1233,N_2737);
and U9864 (N_9864,N_4384,N_1296);
nand U9865 (N_9865,N_495,N_1397);
or U9866 (N_9866,N_3052,N_1395);
or U9867 (N_9867,N_584,N_1334);
and U9868 (N_9868,N_3697,N_4232);
or U9869 (N_9869,N_1991,N_545);
or U9870 (N_9870,N_4394,N_4761);
nand U9871 (N_9871,N_4134,N_4894);
and U9872 (N_9872,N_2316,N_4390);
or U9873 (N_9873,N_539,N_979);
and U9874 (N_9874,N_4139,N_2613);
or U9875 (N_9875,N_3763,N_101);
or U9876 (N_9876,N_1481,N_314);
and U9877 (N_9877,N_4037,N_500);
and U9878 (N_9878,N_1085,N_4234);
and U9879 (N_9879,N_4127,N_1491);
nand U9880 (N_9880,N_2165,N_178);
nand U9881 (N_9881,N_3788,N_3187);
nand U9882 (N_9882,N_2039,N_3945);
nor U9883 (N_9883,N_3794,N_495);
nor U9884 (N_9884,N_1619,N_3862);
or U9885 (N_9885,N_1711,N_2458);
nand U9886 (N_9886,N_3639,N_2875);
nand U9887 (N_9887,N_2168,N_1608);
xnor U9888 (N_9888,N_4173,N_3639);
nand U9889 (N_9889,N_1375,N_4191);
nor U9890 (N_9890,N_2208,N_1265);
nor U9891 (N_9891,N_166,N_2481);
nand U9892 (N_9892,N_3577,N_1963);
or U9893 (N_9893,N_3379,N_2033);
nor U9894 (N_9894,N_4613,N_690);
or U9895 (N_9895,N_3954,N_3700);
nor U9896 (N_9896,N_3178,N_2183);
nor U9897 (N_9897,N_830,N_4097);
nand U9898 (N_9898,N_255,N_2849);
nor U9899 (N_9899,N_2971,N_2282);
nor U9900 (N_9900,N_747,N_2547);
nand U9901 (N_9901,N_2077,N_123);
or U9902 (N_9902,N_4279,N_1776);
or U9903 (N_9903,N_4927,N_781);
nor U9904 (N_9904,N_2051,N_1343);
and U9905 (N_9905,N_46,N_430);
nor U9906 (N_9906,N_418,N_4014);
nor U9907 (N_9907,N_2572,N_804);
and U9908 (N_9908,N_4913,N_350);
or U9909 (N_9909,N_125,N_418);
nand U9910 (N_9910,N_1005,N_865);
nor U9911 (N_9911,N_1643,N_166);
nor U9912 (N_9912,N_4555,N_1021);
and U9913 (N_9913,N_648,N_4174);
or U9914 (N_9914,N_668,N_2996);
nand U9915 (N_9915,N_3898,N_3730);
and U9916 (N_9916,N_906,N_3199);
and U9917 (N_9917,N_4428,N_3777);
nand U9918 (N_9918,N_1910,N_1242);
or U9919 (N_9919,N_4716,N_2159);
xnor U9920 (N_9920,N_1936,N_1656);
nor U9921 (N_9921,N_3219,N_872);
or U9922 (N_9922,N_3532,N_2843);
nand U9923 (N_9923,N_2936,N_1224);
or U9924 (N_9924,N_4895,N_1520);
or U9925 (N_9925,N_144,N_3739);
and U9926 (N_9926,N_4013,N_837);
and U9927 (N_9927,N_1139,N_2261);
nand U9928 (N_9928,N_227,N_2567);
nor U9929 (N_9929,N_3265,N_2289);
or U9930 (N_9930,N_3877,N_436);
nor U9931 (N_9931,N_2465,N_3792);
or U9932 (N_9932,N_3603,N_3321);
nor U9933 (N_9933,N_133,N_1967);
nor U9934 (N_9934,N_1097,N_4278);
nor U9935 (N_9935,N_4023,N_2214);
and U9936 (N_9936,N_4072,N_1286);
or U9937 (N_9937,N_1077,N_3361);
and U9938 (N_9938,N_591,N_4854);
xor U9939 (N_9939,N_803,N_1090);
nand U9940 (N_9940,N_2700,N_4129);
xnor U9941 (N_9941,N_4602,N_2863);
nand U9942 (N_9942,N_1134,N_4941);
nand U9943 (N_9943,N_4535,N_3000);
or U9944 (N_9944,N_3823,N_2529);
nand U9945 (N_9945,N_4003,N_4139);
or U9946 (N_9946,N_3338,N_3794);
nor U9947 (N_9947,N_851,N_4475);
and U9948 (N_9948,N_2940,N_259);
and U9949 (N_9949,N_2455,N_410);
nor U9950 (N_9950,N_861,N_2217);
and U9951 (N_9951,N_1528,N_3325);
or U9952 (N_9952,N_626,N_4768);
xor U9953 (N_9953,N_1034,N_529);
nand U9954 (N_9954,N_581,N_2551);
nor U9955 (N_9955,N_4447,N_849);
nand U9956 (N_9956,N_1468,N_2295);
or U9957 (N_9957,N_3664,N_4171);
or U9958 (N_9958,N_456,N_1525);
or U9959 (N_9959,N_1639,N_1661);
nor U9960 (N_9960,N_3501,N_1718);
or U9961 (N_9961,N_592,N_1279);
nor U9962 (N_9962,N_614,N_4111);
nand U9963 (N_9963,N_1783,N_3545);
and U9964 (N_9964,N_174,N_135);
nor U9965 (N_9965,N_3283,N_1947);
nor U9966 (N_9966,N_3000,N_1467);
or U9967 (N_9967,N_2390,N_2304);
and U9968 (N_9968,N_1409,N_3022);
nand U9969 (N_9969,N_1389,N_1578);
nand U9970 (N_9970,N_950,N_337);
nor U9971 (N_9971,N_3365,N_4561);
nor U9972 (N_9972,N_3573,N_3736);
nand U9973 (N_9973,N_2823,N_2927);
nor U9974 (N_9974,N_2901,N_3697);
nand U9975 (N_9975,N_1739,N_2033);
nand U9976 (N_9976,N_3420,N_3331);
or U9977 (N_9977,N_2224,N_2705);
nand U9978 (N_9978,N_2305,N_3404);
nor U9979 (N_9979,N_1373,N_1770);
nor U9980 (N_9980,N_3347,N_3603);
nand U9981 (N_9981,N_74,N_3957);
and U9982 (N_9982,N_749,N_1079);
nor U9983 (N_9983,N_3586,N_4731);
and U9984 (N_9984,N_315,N_1620);
nand U9985 (N_9985,N_4380,N_1654);
and U9986 (N_9986,N_3813,N_4803);
nand U9987 (N_9987,N_4764,N_3342);
nand U9988 (N_9988,N_3705,N_2864);
nand U9989 (N_9989,N_1660,N_2300);
and U9990 (N_9990,N_2414,N_4858);
or U9991 (N_9991,N_3930,N_2468);
nor U9992 (N_9992,N_4738,N_2775);
or U9993 (N_9993,N_276,N_876);
or U9994 (N_9994,N_4624,N_1484);
and U9995 (N_9995,N_2223,N_4498);
nand U9996 (N_9996,N_3167,N_110);
nand U9997 (N_9997,N_1641,N_1347);
nor U9998 (N_9998,N_2908,N_510);
or U9999 (N_9999,N_580,N_3759);
and U10000 (N_10000,N_5114,N_6929);
and U10001 (N_10001,N_6108,N_8554);
nor U10002 (N_10002,N_7835,N_5727);
and U10003 (N_10003,N_6401,N_6615);
nand U10004 (N_10004,N_6416,N_8252);
nor U10005 (N_10005,N_9651,N_6136);
or U10006 (N_10006,N_7136,N_9935);
nand U10007 (N_10007,N_8332,N_5030);
nand U10008 (N_10008,N_9597,N_5264);
nor U10009 (N_10009,N_7623,N_7668);
nor U10010 (N_10010,N_6697,N_8747);
nor U10011 (N_10011,N_5321,N_6088);
or U10012 (N_10012,N_7893,N_5444);
nand U10013 (N_10013,N_5363,N_6489);
or U10014 (N_10014,N_7114,N_9835);
or U10015 (N_10015,N_6117,N_5620);
and U10016 (N_10016,N_6154,N_6557);
nor U10017 (N_10017,N_7305,N_7041);
nand U10018 (N_10018,N_6734,N_7141);
or U10019 (N_10019,N_8294,N_5557);
nor U10020 (N_10020,N_8160,N_6314);
and U10021 (N_10021,N_7675,N_8094);
nor U10022 (N_10022,N_6083,N_9296);
nand U10023 (N_10023,N_6335,N_7162);
nand U10024 (N_10024,N_9929,N_8658);
and U10025 (N_10025,N_5927,N_5919);
nor U10026 (N_10026,N_5377,N_9174);
and U10027 (N_10027,N_9314,N_6054);
nor U10028 (N_10028,N_5222,N_5379);
nor U10029 (N_10029,N_8320,N_7147);
nand U10030 (N_10030,N_9812,N_6232);
or U10031 (N_10031,N_9680,N_8907);
nand U10032 (N_10032,N_6101,N_9841);
and U10033 (N_10033,N_8020,N_6607);
nand U10034 (N_10034,N_5277,N_9939);
nor U10035 (N_10035,N_6479,N_6482);
nor U10036 (N_10036,N_9095,N_7303);
or U10037 (N_10037,N_7727,N_5064);
or U10038 (N_10038,N_6327,N_5443);
xor U10039 (N_10039,N_7090,N_6063);
nand U10040 (N_10040,N_9354,N_7638);
nand U10041 (N_10041,N_5245,N_9747);
or U10042 (N_10042,N_7430,N_6141);
xnor U10043 (N_10043,N_5118,N_9467);
or U10044 (N_10044,N_6069,N_5068);
and U10045 (N_10045,N_7327,N_8274);
and U10046 (N_10046,N_9344,N_5661);
nor U10047 (N_10047,N_5348,N_7076);
or U10048 (N_10048,N_8607,N_5767);
or U10049 (N_10049,N_6642,N_8847);
xor U10050 (N_10050,N_5232,N_9601);
and U10051 (N_10051,N_8060,N_5105);
nand U10052 (N_10052,N_9479,N_9988);
or U10053 (N_10053,N_5844,N_6654);
nand U10054 (N_10054,N_6725,N_9434);
and U10055 (N_10055,N_8901,N_9888);
or U10056 (N_10056,N_6409,N_9688);
nand U10057 (N_10057,N_9047,N_8871);
nor U10058 (N_10058,N_9053,N_6098);
nand U10059 (N_10059,N_6427,N_8626);
nor U10060 (N_10060,N_9829,N_5129);
or U10061 (N_10061,N_6002,N_5853);
nor U10062 (N_10062,N_6723,N_7115);
and U10063 (N_10063,N_6149,N_9243);
and U10064 (N_10064,N_8667,N_8707);
and U10065 (N_10065,N_9015,N_9216);
xnor U10066 (N_10066,N_7463,N_6158);
and U10067 (N_10067,N_5812,N_5580);
nand U10068 (N_10068,N_8326,N_9814);
nand U10069 (N_10069,N_9778,N_9474);
and U10070 (N_10070,N_7067,N_7832);
nand U10071 (N_10071,N_8042,N_6562);
or U10072 (N_10072,N_8727,N_9007);
nor U10073 (N_10073,N_6528,N_9782);
nand U10074 (N_10074,N_6741,N_7402);
nor U10075 (N_10075,N_8759,N_5044);
or U10076 (N_10076,N_6031,N_6168);
nand U10077 (N_10077,N_6797,N_5378);
nand U10078 (N_10078,N_9683,N_8786);
or U10079 (N_10079,N_6790,N_6203);
and U10080 (N_10080,N_5122,N_5588);
or U10081 (N_10081,N_8186,N_9693);
nand U10082 (N_10082,N_8258,N_7592);
nand U10083 (N_10083,N_8187,N_8022);
or U10084 (N_10084,N_6955,N_7802);
xor U10085 (N_10085,N_5438,N_5263);
nor U10086 (N_10086,N_5560,N_9868);
and U10087 (N_10087,N_5611,N_6922);
and U10088 (N_10088,N_8900,N_6784);
and U10089 (N_10089,N_5704,N_7302);
nand U10090 (N_10090,N_5709,N_5230);
nor U10091 (N_10091,N_8849,N_7806);
nand U10092 (N_10092,N_5052,N_5539);
nand U10093 (N_10093,N_7070,N_7493);
nor U10094 (N_10094,N_7601,N_5080);
or U10095 (N_10095,N_9709,N_9412);
nor U10096 (N_10096,N_5799,N_9126);
nand U10097 (N_10097,N_6817,N_5644);
and U10098 (N_10098,N_7709,N_6605);
or U10099 (N_10099,N_6079,N_8710);
nand U10100 (N_10100,N_8764,N_5858);
nand U10101 (N_10101,N_9227,N_7036);
and U10102 (N_10102,N_7961,N_5914);
or U10103 (N_10103,N_8247,N_6791);
and U10104 (N_10104,N_9067,N_9366);
xnor U10105 (N_10105,N_6833,N_6333);
or U10106 (N_10106,N_8107,N_8008);
or U10107 (N_10107,N_8348,N_6286);
nand U10108 (N_10108,N_9886,N_7932);
nor U10109 (N_10109,N_9637,N_6926);
xnor U10110 (N_10110,N_6344,N_9538);
and U10111 (N_10111,N_5106,N_7117);
xnor U10112 (N_10112,N_8176,N_8814);
nor U10113 (N_10113,N_8261,N_9926);
nor U10114 (N_10114,N_7234,N_7843);
and U10115 (N_10115,N_5651,N_8561);
or U10116 (N_10116,N_9838,N_7164);
nor U10117 (N_10117,N_5745,N_5559);
and U10118 (N_10118,N_7864,N_8706);
nor U10119 (N_10119,N_5362,N_6755);
nor U10120 (N_10120,N_7670,N_5434);
and U10121 (N_10121,N_7973,N_7989);
or U10122 (N_10122,N_7145,N_9490);
nand U10123 (N_10123,N_9547,N_8374);
or U10124 (N_10124,N_8859,N_7081);
nand U10125 (N_10125,N_6614,N_6988);
nor U10126 (N_10126,N_9981,N_5094);
or U10127 (N_10127,N_5375,N_9225);
and U10128 (N_10128,N_5946,N_9566);
nand U10129 (N_10129,N_8352,N_5574);
nand U10130 (N_10130,N_8054,N_7074);
nor U10131 (N_10131,N_5173,N_9898);
or U10132 (N_10132,N_7200,N_9508);
nand U10133 (N_10133,N_6558,N_6771);
nor U10134 (N_10134,N_9417,N_9735);
nor U10135 (N_10135,N_7683,N_5325);
nand U10136 (N_10136,N_9327,N_7772);
or U10137 (N_10137,N_9828,N_6356);
or U10138 (N_10138,N_9658,N_8182);
nor U10139 (N_10139,N_8991,N_8314);
nand U10140 (N_10140,N_7744,N_6392);
and U10141 (N_10141,N_7272,N_7578);
or U10142 (N_10142,N_7982,N_6243);
and U10143 (N_10143,N_8582,N_7176);
nand U10144 (N_10144,N_6729,N_8244);
nor U10145 (N_10145,N_8618,N_5784);
nand U10146 (N_10146,N_6431,N_9920);
or U10147 (N_10147,N_5758,N_5857);
nor U10148 (N_10148,N_5600,N_8532);
or U10149 (N_10149,N_7531,N_6980);
and U10150 (N_10150,N_5616,N_8510);
and U10151 (N_10151,N_8179,N_7049);
nand U10152 (N_10152,N_8192,N_9050);
nand U10153 (N_10153,N_9757,N_6722);
nand U10154 (N_10154,N_5630,N_9671);
nor U10155 (N_10155,N_7376,N_9315);
and U10156 (N_10156,N_6318,N_8905);
or U10157 (N_10157,N_7016,N_6399);
nor U10158 (N_10158,N_8389,N_6381);
nand U10159 (N_10159,N_6444,N_9144);
and U10160 (N_10160,N_8406,N_8290);
nor U10161 (N_10161,N_5934,N_8169);
nand U10162 (N_10162,N_8584,N_5199);
nor U10163 (N_10163,N_5386,N_7833);
or U10164 (N_10164,N_9745,N_7439);
and U10165 (N_10165,N_5452,N_8307);
or U10166 (N_10166,N_8789,N_7228);
nand U10167 (N_10167,N_8875,N_7552);
nand U10168 (N_10168,N_9294,N_8914);
nand U10169 (N_10169,N_6897,N_8181);
nand U10170 (N_10170,N_8830,N_8453);
or U10171 (N_10171,N_8629,N_6024);
or U10172 (N_10172,N_5387,N_6257);
or U10173 (N_10173,N_9101,N_6801);
or U10174 (N_10174,N_7087,N_6813);
xnor U10175 (N_10175,N_9178,N_5982);
nand U10176 (N_10176,N_8185,N_5200);
nand U10177 (N_10177,N_9990,N_8865);
nor U10178 (N_10178,N_5150,N_5806);
or U10179 (N_10179,N_9332,N_8306);
and U10180 (N_10180,N_8207,N_5132);
nor U10181 (N_10181,N_5191,N_7227);
nor U10182 (N_10182,N_5111,N_5728);
nand U10183 (N_10183,N_9030,N_9065);
or U10184 (N_10184,N_7357,N_5936);
nand U10185 (N_10185,N_9617,N_7572);
nand U10186 (N_10186,N_6183,N_6347);
nand U10187 (N_10187,N_8180,N_8354);
nand U10188 (N_10188,N_9020,N_7192);
nand U10189 (N_10189,N_7970,N_6857);
nor U10190 (N_10190,N_9131,N_5318);
or U10191 (N_10191,N_8044,N_6402);
nand U10192 (N_10192,N_6421,N_8709);
xnor U10193 (N_10193,N_5022,N_7980);
and U10194 (N_10194,N_7766,N_7025);
nand U10195 (N_10195,N_6586,N_9940);
nor U10196 (N_10196,N_9529,N_5324);
or U10197 (N_10197,N_6037,N_6685);
and U10198 (N_10198,N_9567,N_6084);
nand U10199 (N_10199,N_9060,N_7570);
and U10200 (N_10200,N_7129,N_9260);
and U10201 (N_10201,N_6550,N_5592);
nor U10202 (N_10202,N_5859,N_9207);
or U10203 (N_10203,N_8072,N_7914);
nor U10204 (N_10204,N_9739,N_9188);
or U10205 (N_10205,N_9179,N_8704);
nand U10206 (N_10206,N_6704,N_7134);
and U10207 (N_10207,N_6360,N_6923);
nand U10208 (N_10208,N_6345,N_8712);
nand U10209 (N_10209,N_7705,N_9117);
xor U10210 (N_10210,N_9218,N_5718);
or U10211 (N_10211,N_8965,N_6390);
or U10212 (N_10212,N_7786,N_9644);
nand U10213 (N_10213,N_6748,N_5097);
nand U10214 (N_10214,N_8347,N_6008);
nor U10215 (N_10215,N_5698,N_6361);
nand U10216 (N_10216,N_8587,N_6966);
and U10217 (N_10217,N_8446,N_8810);
or U10218 (N_10218,N_7886,N_8911);
nand U10219 (N_10219,N_8735,N_6800);
nand U10220 (N_10220,N_8249,N_9203);
nor U10221 (N_10221,N_9469,N_5506);
nand U10222 (N_10222,N_5912,N_8264);
nand U10223 (N_10223,N_9071,N_6250);
nor U10224 (N_10224,N_6716,N_7512);
or U10225 (N_10225,N_7437,N_7538);
or U10226 (N_10226,N_7329,N_7651);
or U10227 (N_10227,N_9970,N_7157);
nor U10228 (N_10228,N_8489,N_8550);
nand U10229 (N_10229,N_7776,N_9682);
or U10230 (N_10230,N_8482,N_5167);
nand U10231 (N_10231,N_8571,N_7729);
or U10232 (N_10232,N_9702,N_5170);
nand U10233 (N_10233,N_8864,N_8337);
nor U10234 (N_10234,N_9790,N_7276);
or U10235 (N_10235,N_8619,N_8127);
nand U10236 (N_10236,N_5025,N_5641);
nor U10237 (N_10237,N_6004,N_5038);
or U10238 (N_10238,N_5637,N_6611);
xnor U10239 (N_10239,N_9026,N_9480);
nor U10240 (N_10240,N_8038,N_8139);
or U10241 (N_10241,N_5259,N_7896);
and U10242 (N_10242,N_9403,N_8994);
or U10243 (N_10243,N_9191,N_9621);
or U10244 (N_10244,N_8271,N_6028);
and U10245 (N_10245,N_5138,N_8670);
nor U10246 (N_10246,N_7356,N_7678);
and U10247 (N_10247,N_5107,N_7880);
or U10248 (N_10248,N_5903,N_7490);
nand U10249 (N_10249,N_5370,N_7354);
or U10250 (N_10250,N_5127,N_8310);
nor U10251 (N_10251,N_9370,N_5341);
nand U10252 (N_10252,N_9011,N_8442);
nor U10253 (N_10253,N_8867,N_6446);
and U10254 (N_10254,N_5531,N_5490);
or U10255 (N_10255,N_5124,N_5313);
or U10256 (N_10256,N_9805,N_6698);
nor U10257 (N_10257,N_8818,N_9168);
and U10258 (N_10258,N_6694,N_8535);
or U10259 (N_10259,N_8476,N_9088);
nor U10260 (N_10260,N_5078,N_9731);
and U10261 (N_10261,N_5954,N_7604);
nor U10262 (N_10262,N_9789,N_7722);
and U10263 (N_10263,N_9686,N_9699);
or U10264 (N_10264,N_9119,N_9404);
and U10265 (N_10265,N_7960,N_5904);
and U10266 (N_10266,N_9595,N_5890);
and U10267 (N_10267,N_5461,N_5652);
nand U10268 (N_10268,N_7353,N_8408);
and U10269 (N_10269,N_8073,N_7718);
nor U10270 (N_10270,N_9994,N_7467);
nand U10271 (N_10271,N_8080,N_6161);
or U10272 (N_10272,N_6169,N_7630);
nor U10273 (N_10273,N_7173,N_6921);
nand U10274 (N_10274,N_9295,N_5713);
or U10275 (N_10275,N_5149,N_5163);
or U10276 (N_10276,N_6012,N_6653);
nor U10277 (N_10277,N_9608,N_9389);
or U10278 (N_10278,N_6320,N_6543);
nand U10279 (N_10279,N_8597,N_6647);
nand U10280 (N_10280,N_9733,N_9063);
and U10281 (N_10281,N_6513,N_5683);
nand U10282 (N_10282,N_9411,N_8518);
nand U10283 (N_10283,N_5034,N_8769);
or U10284 (N_10284,N_7548,N_6567);
nand U10285 (N_10285,N_7794,N_9717);
or U10286 (N_10286,N_5162,N_5000);
xnor U10287 (N_10287,N_5270,N_6452);
or U10288 (N_10288,N_8996,N_5288);
nor U10289 (N_10289,N_5763,N_9276);
and U10290 (N_10290,N_9158,N_8763);
nor U10291 (N_10291,N_7023,N_8303);
nor U10292 (N_10292,N_7213,N_9330);
and U10293 (N_10293,N_8342,N_5194);
nand U10294 (N_10294,N_8196,N_7253);
nor U10295 (N_10295,N_8552,N_9380);
or U10296 (N_10296,N_8205,N_6827);
and U10297 (N_10297,N_6093,N_8633);
nor U10298 (N_10298,N_5005,N_7805);
nand U10299 (N_10299,N_7998,N_9570);
xor U10300 (N_10300,N_7486,N_6096);
nor U10301 (N_10301,N_8108,N_9130);
xor U10302 (N_10302,N_9541,N_9152);
nand U10303 (N_10303,N_7361,N_9077);
and U10304 (N_10304,N_9204,N_7482);
and U10305 (N_10305,N_7244,N_6125);
nand U10306 (N_10306,N_8239,N_5887);
nor U10307 (N_10307,N_8572,N_8775);
nand U10308 (N_10308,N_6739,N_8212);
nand U10309 (N_10309,N_8464,N_5441);
or U10310 (N_10310,N_5722,N_8642);
nor U10311 (N_10311,N_8330,N_7316);
or U10312 (N_10312,N_7257,N_9664);
or U10313 (N_10313,N_8019,N_8887);
nor U10314 (N_10314,N_8988,N_9073);
or U10315 (N_10315,N_8266,N_7250);
nor U10316 (N_10316,N_8088,N_9925);
and U10317 (N_10317,N_9362,N_9445);
nand U10318 (N_10318,N_7518,N_6112);
nor U10319 (N_10319,N_9718,N_6309);
nand U10320 (N_10320,N_5468,N_9599);
nand U10321 (N_10321,N_7990,N_7195);
nand U10322 (N_10322,N_7814,N_9794);
or U10323 (N_10323,N_9714,N_6295);
or U10324 (N_10324,N_9748,N_7922);
nand U10325 (N_10325,N_8715,N_9464);
nand U10326 (N_10326,N_9409,N_9236);
nor U10327 (N_10327,N_9918,N_5888);
and U10328 (N_10328,N_8652,N_6786);
or U10329 (N_10329,N_6672,N_8774);
nand U10330 (N_10330,N_9230,N_6041);
or U10331 (N_10331,N_8257,N_7241);
nand U10332 (N_10332,N_7274,N_8158);
nor U10333 (N_10333,N_8190,N_8079);
or U10334 (N_10334,N_9522,N_8195);
nor U10335 (N_10335,N_5885,N_8673);
and U10336 (N_10336,N_7608,N_6764);
nand U10337 (N_10337,N_7889,N_6167);
nor U10338 (N_10338,N_5175,N_7908);
nor U10339 (N_10339,N_8897,N_7645);
nand U10340 (N_10340,N_7819,N_8492);
or U10341 (N_10341,N_5793,N_9750);
nor U10342 (N_10342,N_6463,N_7046);
and U10343 (N_10343,N_7554,N_5555);
or U10344 (N_10344,N_6525,N_7974);
and U10345 (N_10345,N_6864,N_7054);
and U10346 (N_10346,N_7730,N_5602);
and U10347 (N_10347,N_5514,N_5762);
or U10348 (N_10348,N_5673,N_6546);
nor U10349 (N_10349,N_7954,N_6200);
nor U10350 (N_10350,N_7428,N_6821);
or U10351 (N_10351,N_7334,N_5322);
nand U10352 (N_10352,N_7897,N_6754);
nor U10353 (N_10353,N_9674,N_5096);
nor U10354 (N_10354,N_9321,N_5234);
nand U10355 (N_10355,N_9725,N_7348);
nor U10356 (N_10356,N_8889,N_8375);
nand U10357 (N_10357,N_5835,N_6506);
nand U10358 (N_10358,N_5723,N_7101);
nand U10359 (N_10359,N_7196,N_7745);
nand U10360 (N_10360,N_5686,N_9081);
or U10361 (N_10361,N_5100,N_6204);
and U10362 (N_10362,N_9105,N_8409);
or U10363 (N_10363,N_8308,N_5846);
and U10364 (N_10364,N_8784,N_5818);
and U10365 (N_10365,N_5119,N_6695);
and U10366 (N_10366,N_7643,N_9313);
and U10367 (N_10367,N_5821,N_5586);
nor U10368 (N_10368,N_8119,N_6820);
and U10369 (N_10369,N_5569,N_5448);
or U10370 (N_10370,N_6035,N_6999);
nor U10371 (N_10371,N_6175,N_5057);
nor U10372 (N_10372,N_6102,N_9099);
or U10373 (N_10373,N_7323,N_7541);
or U10374 (N_10374,N_5629,N_6325);
nand U10375 (N_10375,N_9799,N_6619);
or U10376 (N_10376,N_6376,N_9211);
nand U10377 (N_10377,N_9952,N_9684);
and U10378 (N_10378,N_6027,N_6227);
nand U10379 (N_10379,N_8002,N_8318);
and U10380 (N_10380,N_6106,N_5649);
or U10381 (N_10381,N_8516,N_8245);
or U10382 (N_10382,N_8113,N_8728);
nor U10383 (N_10383,N_9571,N_9549);
and U10384 (N_10384,N_9390,N_9496);
and U10385 (N_10385,N_6889,N_6851);
nor U10386 (N_10386,N_8220,N_7442);
and U10387 (N_10387,N_5613,N_6850);
nor U10388 (N_10388,N_8100,N_5480);
and U10389 (N_10389,N_6991,N_8285);
nand U10390 (N_10390,N_6588,N_5014);
nand U10391 (N_10391,N_6599,N_9233);
nand U10392 (N_10392,N_9863,N_8105);
and U10393 (N_10393,N_5524,N_9420);
nor U10394 (N_10394,N_8566,N_9641);
and U10395 (N_10395,N_7952,N_6042);
nand U10396 (N_10396,N_5986,N_6290);
nand U10397 (N_10397,N_8070,N_7471);
nand U10398 (N_10398,N_7803,N_6738);
nand U10399 (N_10399,N_9269,N_8263);
nand U10400 (N_10400,N_8349,N_5258);
and U10401 (N_10401,N_9051,N_9226);
nand U10402 (N_10402,N_5892,N_8369);
nor U10403 (N_10403,N_8420,N_7462);
or U10404 (N_10404,N_8890,N_7539);
or U10405 (N_10405,N_8421,N_6901);
nor U10406 (N_10406,N_5523,N_8678);
or U10407 (N_10407,N_8504,N_7171);
nor U10408 (N_10408,N_8544,N_5721);
nand U10409 (N_10409,N_7262,N_7060);
nand U10410 (N_10410,N_9044,N_5367);
or U10411 (N_10411,N_6089,N_6673);
xnor U10412 (N_10412,N_9447,N_7965);
and U10413 (N_10413,N_8857,N_6792);
nand U10414 (N_10414,N_6499,N_7288);
and U10415 (N_10415,N_5248,N_6278);
nor U10416 (N_10416,N_6486,N_6420);
and U10417 (N_10417,N_9628,N_6856);
or U10418 (N_10418,N_9033,N_5478);
nor U10419 (N_10419,N_8843,N_8280);
xor U10420 (N_10420,N_7975,N_5371);
or U10421 (N_10421,N_6266,N_9758);
nand U10422 (N_10422,N_7149,N_9763);
nor U10423 (N_10423,N_6000,N_9086);
nand U10424 (N_10424,N_5732,N_6458);
nand U10425 (N_10425,N_9610,N_9552);
nor U10426 (N_10426,N_8688,N_6223);
or U10427 (N_10427,N_7088,N_6964);
nor U10428 (N_10428,N_5414,N_5393);
and U10429 (N_10429,N_9631,N_5210);
nand U10430 (N_10430,N_5016,N_5749);
and U10431 (N_10431,N_8522,N_9328);
nand U10432 (N_10432,N_9183,N_5518);
nor U10433 (N_10433,N_7861,N_6386);
or U10434 (N_10434,N_8570,N_5561);
nand U10435 (N_10435,N_8436,N_5423);
nor U10436 (N_10436,N_9210,N_7579);
and U10437 (N_10437,N_8242,N_5071);
nor U10438 (N_10438,N_6293,N_7092);
or U10439 (N_10439,N_8173,N_9110);
nand U10440 (N_10440,N_6366,N_6828);
or U10441 (N_10441,N_7315,N_8809);
and U10442 (N_10442,N_6689,N_8831);
nand U10443 (N_10443,N_8077,N_7432);
and U10444 (N_10444,N_5553,N_7130);
and U10445 (N_10445,N_7091,N_6811);
nand U10446 (N_10446,N_7169,N_5121);
or U10447 (N_10447,N_9924,N_5027);
nor U10448 (N_10448,N_6371,N_7947);
nor U10449 (N_10449,N_6329,N_9859);
nor U10450 (N_10450,N_7717,N_8665);
nor U10451 (N_10451,N_7589,N_7199);
nand U10452 (N_10452,N_6709,N_7505);
nor U10453 (N_10453,N_6571,N_9652);
xnor U10454 (N_10454,N_6807,N_7905);
nor U10455 (N_10455,N_7594,N_6467);
nand U10456 (N_10456,N_6737,N_7161);
or U10457 (N_10457,N_9826,N_6835);
nand U10458 (N_10458,N_8846,N_8718);
and U10459 (N_10459,N_5719,N_7930);
nor U10460 (N_10460,N_5664,N_9079);
nand U10461 (N_10461,N_9300,N_9115);
nand U10462 (N_10462,N_9869,N_5999);
and U10463 (N_10463,N_8423,N_7454);
nor U10464 (N_10464,N_7816,N_6812);
and U10465 (N_10465,N_8917,N_5372);
and U10466 (N_10466,N_6869,N_5233);
nand U10467 (N_10467,N_6221,N_6814);
nand U10468 (N_10468,N_7218,N_8376);
and U10469 (N_10469,N_9930,N_5931);
nand U10470 (N_10470,N_9998,N_8794);
nand U10471 (N_10471,N_8136,N_9944);
and U10472 (N_10472,N_5220,N_5457);
and U10473 (N_10473,N_8526,N_7798);
or U10474 (N_10474,N_5881,N_6520);
nand U10475 (N_10475,N_7118,N_9452);
and U10476 (N_10476,N_9304,N_5069);
or U10477 (N_10477,N_7618,N_5421);
and U10478 (N_10478,N_9726,N_6603);
nor U10479 (N_10479,N_6690,N_8654);
nand U10480 (N_10480,N_9292,N_5843);
nor U10481 (N_10481,N_8366,N_9329);
and U10482 (N_10482,N_7089,N_7494);
nand U10483 (N_10483,N_8201,N_9979);
nor U10484 (N_10484,N_7193,N_8432);
xor U10485 (N_10485,N_9374,N_6981);
and U10486 (N_10486,N_7821,N_8145);
and U10487 (N_10487,N_8651,N_8426);
or U10488 (N_10488,N_7155,N_9816);
nand U10489 (N_10489,N_7993,N_7544);
xor U10490 (N_10490,N_5204,N_7808);
nor U10491 (N_10491,N_7152,N_5939);
and U10492 (N_10492,N_9734,N_7923);
xnor U10493 (N_10493,N_9556,N_9796);
nor U10494 (N_10494,N_7211,N_8361);
nor U10495 (N_10495,N_7953,N_9883);
and U10496 (N_10496,N_9677,N_6968);
nand U10497 (N_10497,N_7981,N_5527);
and U10498 (N_10498,N_7720,N_6246);
and U10499 (N_10499,N_5612,N_5023);
nand U10500 (N_10500,N_8997,N_5739);
or U10501 (N_10501,N_5413,N_6013);
nand U10502 (N_10502,N_7966,N_5201);
or U10503 (N_10503,N_6066,N_6395);
nand U10504 (N_10504,N_9845,N_9128);
or U10505 (N_10505,N_6408,N_9710);
or U10506 (N_10506,N_7292,N_5275);
nor U10507 (N_10507,N_9359,N_5823);
nor U10508 (N_10508,N_5212,N_6214);
and U10509 (N_10509,N_5312,N_6116);
nand U10510 (N_10510,N_5225,N_5469);
nand U10511 (N_10511,N_6618,N_6488);
or U10512 (N_10512,N_9217,N_9807);
nor U10513 (N_10513,N_8740,N_5813);
and U10514 (N_10514,N_9833,N_5394);
nand U10515 (N_10515,N_7167,N_7962);
nand U10516 (N_10516,N_9629,N_8780);
nor U10517 (N_10517,N_5384,N_5929);
nand U10518 (N_10518,N_8174,N_9879);
and U10519 (N_10519,N_7656,N_6132);
nand U10520 (N_10520,N_7921,N_5898);
or U10521 (N_10521,N_5778,N_8329);
or U10522 (N_10522,N_6606,N_9423);
or U10523 (N_10523,N_5872,N_7456);
nor U10524 (N_10524,N_7109,N_7511);
nor U10525 (N_10525,N_9408,N_8690);
or U10526 (N_10526,N_6776,N_5507);
or U10527 (N_10527,N_6773,N_9061);
or U10528 (N_10528,N_9159,N_7687);
or U10529 (N_10529,N_9375,N_8255);
nor U10530 (N_10530,N_7321,N_8156);
nor U10531 (N_10531,N_5740,N_9909);
nand U10532 (N_10532,N_5925,N_8048);
and U10533 (N_10533,N_9536,N_5143);
or U10534 (N_10534,N_7862,N_7841);
or U10535 (N_10535,N_7634,N_9336);
nor U10536 (N_10536,N_9546,N_5422);
and U10537 (N_10537,N_7300,N_8229);
nand U10538 (N_10538,N_5766,N_5980);
or U10539 (N_10539,N_9715,N_8703);
or U10540 (N_10540,N_5416,N_7865);
nand U10541 (N_10541,N_9881,N_9766);
and U10542 (N_10542,N_6504,N_6663);
and U10543 (N_10543,N_8799,N_7820);
xor U10544 (N_10544,N_6404,N_6670);
or U10545 (N_10545,N_8480,N_5356);
nand U10546 (N_10546,N_5847,N_6691);
or U10547 (N_10547,N_9820,N_7688);
and U10548 (N_10548,N_6505,N_9986);
nor U10549 (N_10549,N_6808,N_6403);
nand U10550 (N_10550,N_5614,N_9742);
and U10551 (N_10551,N_9850,N_6992);
nand U10552 (N_10552,N_6338,N_5832);
xor U10553 (N_10553,N_5789,N_5460);
or U10554 (N_10554,N_6058,N_6118);
nand U10555 (N_10555,N_9724,N_6628);
and U10556 (N_10556,N_7751,N_5998);
or U10557 (N_10557,N_8569,N_6536);
nand U10558 (N_10558,N_7423,N_9908);
nor U10559 (N_10559,N_6336,N_7613);
nor U10560 (N_10560,N_9153,N_9554);
or U10561 (N_10561,N_8881,N_7750);
and U10562 (N_10562,N_6579,N_9035);
nand U10563 (N_10563,N_9421,N_6524);
nor U10564 (N_10564,N_9842,N_5439);
nand U10565 (N_10565,N_8194,N_6919);
and U10566 (N_10566,N_7684,N_5975);
nand U10567 (N_10567,N_5228,N_6255);
nor U10568 (N_10568,N_5577,N_5581);
nand U10569 (N_10569,N_5601,N_5817);
nand U10570 (N_10570,N_9520,N_5015);
nand U10571 (N_10571,N_5188,N_7278);
and U10572 (N_10572,N_7753,N_6906);
nor U10573 (N_10573,N_8978,N_7254);
or U10574 (N_10574,N_6534,N_6022);
nand U10575 (N_10575,N_5737,N_5746);
nand U10576 (N_10576,N_9106,N_5962);
or U10577 (N_10577,N_6794,N_5177);
and U10578 (N_10578,N_5195,N_7264);
nand U10579 (N_10579,N_9193,N_7170);
or U10580 (N_10580,N_5063,N_7660);
xnor U10581 (N_10581,N_7414,N_9592);
nor U10582 (N_10582,N_5864,N_9271);
nor U10583 (N_10583,N_9082,N_7148);
and U10584 (N_10584,N_7112,N_7191);
nor U10585 (N_10585,N_6388,N_5305);
nand U10586 (N_10586,N_9055,N_7606);
and U10587 (N_10587,N_7230,N_6418);
nand U10588 (N_10588,N_7568,N_7810);
nor U10589 (N_10589,N_8487,N_5726);
xor U10590 (N_10590,N_7163,N_6779);
xor U10591 (N_10591,N_9864,N_7530);
or U10592 (N_10592,N_8081,N_9264);
or U10593 (N_10593,N_8672,N_8806);
or U10594 (N_10594,N_6241,N_5109);
and U10595 (N_10595,N_5902,N_5236);
nor U10596 (N_10596,N_6945,N_5807);
or U10597 (N_10597,N_9577,N_7299);
nor U10598 (N_10598,N_7464,N_7723);
nor U10599 (N_10599,N_7602,N_5590);
or U10600 (N_10600,N_8793,N_5529);
nand U10601 (N_10601,N_8204,N_7079);
and U10602 (N_10602,N_9885,N_6184);
or U10603 (N_10603,N_7759,N_6898);
nand U10604 (N_10604,N_7116,N_7069);
or U10605 (N_10605,N_5435,N_6448);
nand U10606 (N_10606,N_8863,N_6492);
nor U10607 (N_10607,N_8581,N_5058);
nand U10608 (N_10608,N_5113,N_9346);
nor U10609 (N_10609,N_6507,N_6609);
nand U10610 (N_10610,N_6902,N_9273);
nor U10611 (N_10611,N_8101,N_5943);
nor U10612 (N_10612,N_7917,N_5791);
nand U10613 (N_10613,N_8679,N_8430);
and U10614 (N_10614,N_7510,N_7206);
nor U10615 (N_10615,N_9316,N_9510);
xor U10616 (N_10616,N_7096,N_8473);
nor U10617 (N_10617,N_6429,N_7680);
nand U10618 (N_10618,N_8339,N_8284);
xor U10619 (N_10619,N_8798,N_9756);
xor U10620 (N_10620,N_6860,N_6449);
or U10621 (N_10621,N_5395,N_8371);
or U10622 (N_10622,N_6303,N_9603);
and U10623 (N_10623,N_8097,N_5689);
nand U10624 (N_10624,N_7328,N_8017);
and U10625 (N_10625,N_6891,N_6206);
or U10626 (N_10626,N_9148,N_6852);
nand U10627 (N_10627,N_7249,N_6720);
and U10628 (N_10628,N_9847,N_6038);
nand U10629 (N_10629,N_9494,N_6358);
nor U10630 (N_10630,N_8995,N_7281);
and U10631 (N_10631,N_5408,N_6264);
or U10632 (N_10632,N_9456,N_6631);
nand U10633 (N_10633,N_9381,N_8828);
and U10634 (N_10634,N_5065,N_6781);
and U10635 (N_10635,N_6359,N_5369);
nand U10636 (N_10636,N_5070,N_9482);
nand U10637 (N_10637,N_9713,N_8608);
or U10638 (N_10638,N_6556,N_8214);
nand U10639 (N_10639,N_7878,N_9252);
or U10640 (N_10640,N_6047,N_7410);
nor U10641 (N_10641,N_8219,N_5033);
and U10642 (N_10642,N_7500,N_8452);
or U10643 (N_10643,N_5973,N_8218);
xnor U10644 (N_10644,N_6190,N_5255);
nor U10645 (N_10645,N_5345,N_5309);
nor U10646 (N_10646,N_8443,N_6568);
nand U10647 (N_10647,N_6052,N_6861);
nand U10648 (N_10648,N_8699,N_9162);
or U10649 (N_10649,N_7858,N_6760);
nor U10650 (N_10650,N_5272,N_6155);
nor U10651 (N_10651,N_6211,N_5035);
nand U10652 (N_10652,N_7240,N_6675);
nor U10653 (N_10653,N_5772,N_6572);
and U10654 (N_10654,N_7142,N_8049);
and U10655 (N_10655,N_8043,N_7409);
nor U10656 (N_10656,N_5102,N_9372);
nor U10657 (N_10657,N_8756,N_9238);
or U10658 (N_10658,N_6016,N_7906);
or U10659 (N_10659,N_5407,N_8327);
or U10660 (N_10660,N_6306,N_7562);
or U10661 (N_10661,N_7536,N_8977);
and U10662 (N_10662,N_6056,N_5428);
xor U10663 (N_10663,N_6364,N_8711);
or U10664 (N_10664,N_5048,N_7469);
or U10665 (N_10665,N_5502,N_5690);
or U10666 (N_10666,N_6355,N_5403);
and U10667 (N_10667,N_7337,N_5298);
or U10668 (N_10668,N_9517,N_8431);
or U10669 (N_10669,N_9242,N_5125);
and U10670 (N_10670,N_6332,N_8708);
nor U10671 (N_10671,N_6730,N_9402);
nor U10672 (N_10672,N_7346,N_8854);
and U10673 (N_10673,N_5653,N_6745);
nand U10674 (N_10674,N_6238,N_6300);
nand U10675 (N_10675,N_8983,N_9668);
or U10676 (N_10676,N_9419,N_7392);
and U10677 (N_10677,N_8893,N_7769);
nor U10678 (N_10678,N_7026,N_8221);
nor U10679 (N_10679,N_5663,N_5306);
nand U10680 (N_10680,N_5640,N_6805);
or U10681 (N_10681,N_8211,N_7673);
xnor U10682 (N_10682,N_8062,N_5049);
nor U10683 (N_10683,N_6627,N_9848);
or U10684 (N_10684,N_7295,N_6752);
nor U10685 (N_10685,N_8472,N_7202);
and U10686 (N_10686,N_5928,N_9014);
xnor U10687 (N_10687,N_5754,N_9560);
or U10688 (N_10688,N_5715,N_5960);
and U10689 (N_10689,N_9351,N_8766);
and U10690 (N_10690,N_5347,N_7030);
and U10691 (N_10691,N_5335,N_5583);
nor U10692 (N_10692,N_9342,N_9853);
or U10693 (N_10693,N_5638,N_6806);
nor U10694 (N_10694,N_7733,N_8910);
and U10695 (N_10695,N_8300,N_5084);
nor U10696 (N_10696,N_6245,N_5090);
or U10697 (N_10697,N_9527,N_9416);
nor U10698 (N_10698,N_7277,N_6383);
nor U10699 (N_10699,N_8947,N_7209);
or U10700 (N_10700,N_9377,N_9904);
and U10701 (N_10701,N_5755,N_8661);
nand U10702 (N_10702,N_5187,N_6530);
nand U10703 (N_10703,N_7185,N_9176);
and U10704 (N_10704,N_5184,N_7029);
nand U10705 (N_10705,N_8161,N_8178);
or U10706 (N_10706,N_5873,N_8191);
or U10707 (N_10707,N_7201,N_5066);
or U10708 (N_10708,N_7859,N_5165);
or U10709 (N_10709,N_5521,N_9645);
nor U10710 (N_10710,N_7028,N_7706);
or U10711 (N_10711,N_5351,N_5702);
nand U10712 (N_10712,N_9614,N_8596);
nor U10713 (N_10713,N_9737,N_6025);
or U10714 (N_10714,N_8412,N_8855);
nand U10715 (N_10715,N_7359,N_6733);
nand U10716 (N_10716,N_7256,N_7543);
nand U10717 (N_10717,N_6990,N_9876);
nor U10718 (N_10718,N_7042,N_5952);
nand U10719 (N_10719,N_8058,N_7696);
nand U10720 (N_10720,N_9830,N_6578);
or U10721 (N_10721,N_8750,N_6146);
nor U10722 (N_10722,N_8268,N_7738);
or U10723 (N_10723,N_7314,N_5147);
nor U10724 (N_10724,N_7949,N_5582);
and U10725 (N_10725,N_7123,N_9224);
and U10726 (N_10726,N_6522,N_5226);
xnor U10727 (N_10727,N_6711,N_7800);
and U10728 (N_10728,N_7637,N_8051);
nor U10729 (N_10729,N_8804,N_6229);
and U10730 (N_10730,N_9956,N_7540);
and U10731 (N_10731,N_8149,N_9291);
xnor U10732 (N_10732,N_5285,N_8979);
and U10733 (N_10733,N_5037,N_9576);
or U10734 (N_10734,N_5656,N_9201);
or U10735 (N_10735,N_9997,N_8934);
and U10736 (N_10736,N_6128,N_9137);
and U10737 (N_10737,N_5319,N_8980);
nor U10738 (N_10738,N_8873,N_9383);
nand U10739 (N_10739,N_5152,N_7019);
nor U10740 (N_10740,N_5360,N_9523);
and U10741 (N_10741,N_8919,N_7285);
nor U10742 (N_10742,N_7449,N_8237);
or U10743 (N_10743,N_8719,N_7559);
or U10744 (N_10744,N_8741,N_8834);
nor U10745 (N_10745,N_5429,N_5227);
nor U10746 (N_10746,N_8114,N_6585);
nand U10747 (N_10747,N_5672,N_8009);
nand U10748 (N_10748,N_5160,N_6055);
nand U10749 (N_10749,N_5522,N_5752);
xor U10750 (N_10750,N_9116,N_8018);
or U10751 (N_10751,N_8331,N_5747);
and U10752 (N_10752,N_8413,N_9596);
or U10753 (N_10753,N_5814,N_8289);
or U10754 (N_10754,N_8796,N_7397);
and U10755 (N_10755,N_9989,N_7065);
or U10756 (N_10756,N_7676,N_6270);
nand U10757 (N_10757,N_9973,N_8091);
nand U10758 (N_10758,N_5886,N_9430);
nor U10759 (N_10759,N_5028,N_7024);
nor U10760 (N_10760,N_8951,N_8035);
and U10761 (N_10761,N_5894,N_9132);
and U10762 (N_10762,N_6310,N_8069);
or U10763 (N_10763,N_6163,N_9045);
nor U10764 (N_10764,N_6459,N_5499);
and U10765 (N_10765,N_6077,N_5850);
or U10766 (N_10766,N_9676,N_7520);
or U10767 (N_10767,N_7537,N_8466);
or U10768 (N_10768,N_6382,N_9484);
or U10769 (N_10769,N_6177,N_6050);
nand U10770 (N_10770,N_8842,N_8686);
and U10771 (N_10771,N_9440,N_9036);
and U10772 (N_10772,N_8116,N_7818);
or U10773 (N_10773,N_7458,N_7979);
nand U10774 (N_10774,N_9730,N_6198);
nor U10775 (N_10775,N_7689,N_5951);
nand U10776 (N_10776,N_7870,N_6893);
nor U10777 (N_10777,N_9307,N_6021);
or U10778 (N_10778,N_5411,N_8783);
nand U10779 (N_10779,N_7693,N_7894);
nor U10780 (N_10780,N_6215,N_8567);
or U10781 (N_10781,N_9360,N_9278);
or U10782 (N_10782,N_6236,N_6848);
or U10783 (N_10783,N_5819,N_7556);
nand U10784 (N_10784,N_5012,N_8397);
nand U10785 (N_10785,N_6617,N_7120);
and U10786 (N_10786,N_8010,N_6143);
xnor U10787 (N_10787,N_8954,N_9518);
nor U10788 (N_10788,N_6085,N_6057);
and U10789 (N_10789,N_8573,N_8964);
nor U10790 (N_10790,N_7021,N_9921);
nor U10791 (N_10791,N_6712,N_7313);
xnor U10792 (N_10792,N_7611,N_8669);
and U10793 (N_10793,N_8296,N_5491);
or U10794 (N_10794,N_6139,N_7597);
xnor U10795 (N_10795,N_5376,N_7855);
or U10796 (N_10796,N_7752,N_5585);
nand U10797 (N_10797,N_8171,N_8985);
nand U10798 (N_10798,N_5575,N_7848);
and U10799 (N_10799,N_8316,N_7985);
nand U10800 (N_10800,N_5970,N_7996);
nor U10801 (N_10801,N_8753,N_6292);
nand U10802 (N_10802,N_6064,N_9586);
nor U10803 (N_10803,N_6570,N_9205);
nor U10804 (N_10804,N_5445,N_6126);
nand U10805 (N_10805,N_5838,N_7154);
xor U10806 (N_10806,N_6468,N_9437);
or U10807 (N_10807,N_6406,N_9453);
and U10808 (N_10808,N_6514,N_8729);
or U10809 (N_10809,N_7403,N_5417);
and U10810 (N_10810,N_9272,N_7887);
nor U10811 (N_10811,N_6877,N_7452);
or U10812 (N_10812,N_8370,N_7177);
nand U10813 (N_10813,N_6625,N_7742);
and U10814 (N_10814,N_7052,N_6235);
and U10815 (N_10815,N_9854,N_6517);
and U10816 (N_10816,N_7627,N_6900);
and U10817 (N_10817,N_8013,N_7100);
and U10818 (N_10818,N_8826,N_6884);
nand U10819 (N_10819,N_9991,N_6879);
or U10820 (N_10820,N_8527,N_5108);
nor U10821 (N_10821,N_6702,N_8427);
xnor U10822 (N_10822,N_9602,N_6944);
and U10823 (N_10823,N_5475,N_8283);
and U10824 (N_10824,N_8998,N_6197);
and U10825 (N_10825,N_7526,N_5390);
or U10826 (N_10826,N_6831,N_6304);
nor U10827 (N_10827,N_6460,N_8695);
and U10828 (N_10828,N_9967,N_6260);
nand U10829 (N_10829,N_9743,N_8501);
or U10830 (N_10830,N_6140,N_9971);
nor U10831 (N_10831,N_8888,N_9701);
and U10832 (N_10832,N_5598,N_5549);
and U10833 (N_10833,N_9785,N_7061);
xor U10834 (N_10834,N_7884,N_9459);
nand U10835 (N_10835,N_9400,N_5291);
nand U10836 (N_10836,N_8134,N_9667);
or U10837 (N_10837,N_8465,N_6009);
xor U10838 (N_10838,N_6535,N_9513);
or U10839 (N_10839,N_7926,N_6751);
and U10840 (N_10840,N_6878,N_7817);
nor U10841 (N_10841,N_6648,N_8143);
xnor U10842 (N_10842,N_8411,N_9764);
or U10843 (N_10843,N_7555,N_6707);
and U10844 (N_10844,N_7804,N_6896);
nand U10845 (N_10845,N_6967,N_5148);
nand U10846 (N_10846,N_5606,N_5011);
nor U10847 (N_10847,N_5449,N_5430);
or U10848 (N_10848,N_5922,N_8961);
nor U10849 (N_10849,N_5699,N_6462);
and U10850 (N_10850,N_9475,N_8189);
nor U10851 (N_10851,N_6133,N_7341);
nand U10852 (N_10852,N_9647,N_7657);
xor U10853 (N_10853,N_7260,N_9804);
and U10854 (N_10854,N_5282,N_5682);
and U10855 (N_10855,N_9320,N_6836);
nand U10856 (N_10856,N_6151,N_5257);
nor U10857 (N_10857,N_7617,N_9286);
nand U10858 (N_10858,N_6540,N_9305);
nor U10859 (N_10859,N_8338,N_5062);
nand U10860 (N_10860,N_9801,N_7652);
or U10861 (N_10861,N_8309,N_6630);
and U10862 (N_10862,N_8512,N_5576);
and U10863 (N_10863,N_9187,N_6389);
or U10864 (N_10864,N_9882,N_6796);
and U10865 (N_10865,N_7331,N_9927);
or U10866 (N_10866,N_7851,N_6216);
and U10867 (N_10867,N_9208,N_9186);
nor U10868 (N_10868,N_9301,N_5545);
and U10869 (N_10869,N_5398,N_5007);
nand U10870 (N_10870,N_7131,N_6494);
nand U10871 (N_10871,N_9455,N_6271);
and U10872 (N_10872,N_9533,N_5307);
nor U10873 (N_10873,N_8345,N_9964);
nand U10874 (N_10874,N_9942,N_7307);
nand U10875 (N_10875,N_8236,N_6596);
or U10876 (N_10876,N_8358,N_6391);
nor U10877 (N_10877,N_7015,N_6453);
nor U10878 (N_10878,N_7099,N_9246);
nand U10879 (N_10879,N_9251,N_9149);
nand U10880 (N_10880,N_9947,N_6142);
or U10881 (N_10881,N_5547,N_8884);
or U10882 (N_10882,N_5254,N_7420);
nor U10883 (N_10883,N_6785,N_8970);
nand U10884 (N_10884,N_8912,N_5466);
nand U10885 (N_10885,N_5942,N_9878);
and U10886 (N_10886,N_7489,N_8639);
or U10887 (N_10887,N_8021,N_5047);
and U10888 (N_10888,N_9818,N_5515);
and U10889 (N_10889,N_9955,N_5396);
or U10890 (N_10890,N_5117,N_9912);
nor U10891 (N_10891,N_9127,N_6342);
xor U10892 (N_10892,N_9135,N_6934);
nor U10893 (N_10893,N_9995,N_8215);
or U10894 (N_10894,N_9574,N_5945);
nand U10895 (N_10895,N_7984,N_6067);
or U10896 (N_10896,N_5761,N_5642);
and U10897 (N_10897,N_5700,N_6885);
or U10898 (N_10898,N_9783,N_8302);
nand U10899 (N_10899,N_7913,N_6687);
and U10900 (N_10900,N_9363,N_5453);
or U10901 (N_10901,N_6718,N_7582);
or U10902 (N_10902,N_6466,N_8952);
and U10903 (N_10903,N_5330,N_9234);
nand U10904 (N_10904,N_5093,N_5061);
nand U10905 (N_10905,N_6228,N_6483);
or U10906 (N_10906,N_9906,N_5116);
nand U10907 (N_10907,N_7672,N_6708);
and U10908 (N_10908,N_5290,N_8118);
or U10909 (N_10909,N_8694,N_6931);
nand U10910 (N_10910,N_8545,N_6377);
or U10911 (N_10911,N_7535,N_7373);
or U10912 (N_10912,N_6413,N_8240);
xnor U10913 (N_10913,N_8225,N_6301);
or U10914 (N_10914,N_6633,N_6903);
nand U10915 (N_10915,N_8317,N_5297);
nand U10916 (N_10916,N_9615,N_7047);
or U10917 (N_10917,N_7784,N_7749);
and U10918 (N_10918,N_9143,N_9123);
nor U10919 (N_10919,N_8334,N_7083);
and U10920 (N_10920,N_9762,N_5639);
nor U10921 (N_10921,N_7497,N_8491);
nor U10922 (N_10922,N_6935,N_9875);
or U10923 (N_10923,N_6894,N_6268);
nand U10924 (N_10924,N_8429,N_5436);
and U10925 (N_10925,N_6219,N_6011);
and U10926 (N_10926,N_6224,N_8821);
and U10927 (N_10927,N_6859,N_9890);
nor U10928 (N_10928,N_5159,N_8055);
or U10929 (N_10929,N_9993,N_9983);
and U10930 (N_10930,N_5497,N_7221);
nor U10931 (N_10931,N_7144,N_6363);
nor U10932 (N_10932,N_7160,N_8944);
and U10933 (N_10933,N_9540,N_7415);
nor U10934 (N_10934,N_8364,N_5274);
or U10935 (N_10935,N_9449,N_6445);
nand U10936 (N_10936,N_8685,N_7639);
nand U10937 (N_10937,N_7215,N_5172);
or U10938 (N_10938,N_9505,N_5865);
and U10939 (N_10939,N_5142,N_6478);
nand U10940 (N_10940,N_9299,N_5717);
and U10941 (N_10941,N_9436,N_8380);
nand U10942 (N_10942,N_7936,N_8460);
nand U10943 (N_10943,N_9181,N_7596);
nor U10944 (N_10944,N_7967,N_6761);
and U10945 (N_10945,N_8514,N_5043);
nor U10946 (N_10946,N_6425,N_9198);
xor U10947 (N_10947,N_9487,N_5735);
nand U10948 (N_10948,N_8455,N_8790);
nor U10949 (N_10949,N_6331,N_8166);
nand U10950 (N_10950,N_9928,N_6288);
xor U10951 (N_10951,N_6819,N_7394);
and U10952 (N_10952,N_6804,N_5244);
nand U10953 (N_10953,N_9125,N_5292);
nor U10954 (N_10954,N_9704,N_7703);
xnor U10955 (N_10955,N_9163,N_9585);
nand U10956 (N_10956,N_7080,N_6978);
and U10957 (N_10957,N_6422,N_6218);
nor U10958 (N_10958,N_5060,N_7951);
nand U10959 (N_10959,N_6759,N_5072);
and U10960 (N_10960,N_5024,N_8962);
nor U10961 (N_10961,N_7725,N_6289);
or U10962 (N_10962,N_5554,N_7944);
or U10963 (N_10963,N_5868,N_6191);
and U10964 (N_10964,N_8383,N_5486);
nand U10965 (N_10965,N_9199,N_6634);
nand U10966 (N_10966,N_8359,N_6247);
and U10967 (N_10967,N_8130,N_9958);
nor U10968 (N_10968,N_7849,N_9635);
nor U10969 (N_10969,N_9551,N_8990);
nand U10970 (N_10970,N_5280,N_7362);
nand U10971 (N_10971,N_5383,N_5947);
nand U10972 (N_10972,N_6592,N_5537);
or U10973 (N_10973,N_8976,N_8213);
and U10974 (N_10974,N_8368,N_9663);
nand U10975 (N_10975,N_6539,N_9184);
nor U10976 (N_10976,N_9526,N_8177);
nand U10977 (N_10977,N_6946,N_9657);
and U10978 (N_10978,N_9424,N_8539);
and U10979 (N_10979,N_5535,N_8982);
nor U10980 (N_10980,N_8151,N_7686);
and U10981 (N_10981,N_7002,N_6287);
nand U10982 (N_10982,N_5567,N_5800);
nand U10983 (N_10983,N_5705,N_7610);
nand U10984 (N_10984,N_7071,N_8612);
nor U10985 (N_10985,N_5158,N_6357);
and U10986 (N_10986,N_6916,N_8103);
and U10987 (N_10987,N_7567,N_8691);
nor U10988 (N_10988,N_6491,N_6417);
or U10989 (N_10989,N_9290,N_5889);
or U10990 (N_10990,N_9857,N_8922);
nor U10991 (N_10991,N_9140,N_7010);
nor U10992 (N_10992,N_6584,N_7708);
or U10993 (N_10993,N_8050,N_9170);
nor U10994 (N_10994,N_6294,N_7231);
nand U10995 (N_10995,N_8015,N_6230);
nand U10996 (N_10996,N_7137,N_9934);
nor U10997 (N_10997,N_8047,N_8632);
nor U10998 (N_10998,N_6843,N_6455);
or U10999 (N_10999,N_7903,N_9873);
or U11000 (N_11000,N_8485,N_5026);
nor U11001 (N_11001,N_6124,N_8131);
nor U11002 (N_11002,N_8531,N_6872);
nand U11003 (N_11003,N_6302,N_7546);
nor U11004 (N_11004,N_7877,N_8384);
and U11005 (N_11005,N_9435,N_8975);
or U11006 (N_11006,N_5829,N_7842);
nand U11007 (N_11007,N_8636,N_9666);
or U11008 (N_11008,N_8896,N_5092);
nand U11009 (N_11009,N_6501,N_9771);
or U11010 (N_11010,N_5190,N_7268);
nand U11011 (N_11011,N_7710,N_8614);
and U11012 (N_11012,N_8850,N_9960);
nor U11013 (N_11013,N_7916,N_7375);
nor U11014 (N_11014,N_7506,N_9815);
or U11015 (N_11015,N_9248,N_5953);
nand U11016 (N_11016,N_5687,N_6855);
and U11017 (N_11017,N_8388,N_8344);
nor U11018 (N_11018,N_7885,N_7987);
nand U11019 (N_11019,N_6284,N_7955);
or U11020 (N_11020,N_9542,N_7517);
nor U11021 (N_11021,N_9938,N_8424);
and U11022 (N_11022,N_5771,N_9911);
nor U11023 (N_11023,N_8154,N_6749);
nor U11024 (N_11024,N_6643,N_6362);
and U11025 (N_11025,N_7038,N_7626);
nand U11026 (N_11026,N_8456,N_6757);
and U11027 (N_11027,N_5834,N_8754);
nand U11028 (N_11028,N_8099,N_7073);
or U11029 (N_11029,N_7294,N_7839);
nand U11030 (N_11030,N_7846,N_7436);
nor U11031 (N_11031,N_5076,N_5660);
nor U11032 (N_11032,N_9028,N_6908);
or U11033 (N_11033,N_8858,N_7699);
nand U11034 (N_11034,N_7957,N_7728);
nand U11035 (N_11035,N_8202,N_9945);
nand U11036 (N_11036,N_8981,N_7549);
nor U11037 (N_11037,N_9150,N_7583);
nand U11038 (N_11038,N_5785,N_7935);
nor U11039 (N_11039,N_5670,N_5594);
nor U11040 (N_11040,N_8563,N_8851);
nor U11041 (N_11041,N_7182,N_6982);
or U11042 (N_11042,N_5250,N_8410);
or U11043 (N_11043,N_8470,N_8815);
nor U11044 (N_11044,N_7399,N_9495);
xnor U11045 (N_11045,N_7166,N_6984);
nand U11046 (N_11046,N_7925,N_6545);
nor U11047 (N_11047,N_9564,N_6799);
nand U11048 (N_11048,N_9884,N_6495);
and U11049 (N_11049,N_7721,N_7732);
and U11050 (N_11050,N_8521,N_6590);
and U11051 (N_11051,N_7103,N_8335);
nand U11052 (N_11052,N_9650,N_8346);
nand U11053 (N_11053,N_9221,N_9094);
xor U11054 (N_11054,N_5808,N_9414);
nor U11055 (N_11055,N_9626,N_9070);
and U11056 (N_11056,N_6886,N_7135);
or U11057 (N_11057,N_6956,N_8254);
or U11058 (N_11058,N_8515,N_5420);
nor U11059 (N_11059,N_9543,N_8210);
or U11060 (N_11060,N_6099,N_7551);
xnor U11061 (N_11061,N_6575,N_8731);
nor U11062 (N_11062,N_8056,N_9866);
nand U11063 (N_11063,N_9379,N_8676);
nand U11064 (N_11064,N_8395,N_7523);
or U11065 (N_11065,N_9969,N_8394);
and U11066 (N_11066,N_5564,N_8200);
or U11067 (N_11067,N_5877,N_7387);
nor U11068 (N_11068,N_9386,N_5511);
nand U11069 (N_11069,N_5571,N_5716);
and U11070 (N_11070,N_5810,N_5530);
or U11071 (N_11071,N_8869,N_9703);
or U11072 (N_11072,N_7239,N_6581);
and U11073 (N_11073,N_5219,N_9497);
or U11074 (N_11074,N_9019,N_7386);
and U11075 (N_11075,N_5353,N_5628);
and U11076 (N_11076,N_5073,N_9827);
and U11077 (N_11077,N_5548,N_9289);
or U11078 (N_11078,N_8468,N_8785);
nor U11079 (N_11079,N_6005,N_8519);
or U11080 (N_11080,N_5077,N_8634);
nor U11081 (N_11081,N_5694,N_5913);
nor U11082 (N_11082,N_6071,N_8469);
nand U11083 (N_11083,N_7747,N_7158);
or U11084 (N_11084,N_6472,N_8744);
nand U11085 (N_11085,N_5883,N_9166);
or U11086 (N_11086,N_8716,N_6185);
and U11087 (N_11087,N_6237,N_8958);
and U11088 (N_11088,N_6135,N_6768);
nor U11089 (N_11089,N_7174,N_7907);
nand U11090 (N_11090,N_8923,N_9722);
nand U11091 (N_11091,N_9761,N_9946);
nand U11092 (N_11092,N_5311,N_8801);
nand U11093 (N_11093,N_5921,N_9950);
or U11094 (N_11094,N_6130,N_9433);
nor U11095 (N_11095,N_6082,N_9568);
or U11096 (N_11096,N_6503,N_9338);
and U11097 (N_11097,N_9172,N_6498);
nor U11098 (N_11098,N_5786,N_8551);
nand U11099 (N_11099,N_8277,N_6762);
nor U11100 (N_11100,N_8012,N_7032);
and U11101 (N_11101,N_8671,N_9232);
nand U11102 (N_11102,N_9237,N_7831);
or U11103 (N_11103,N_7455,N_5380);
nor U11104 (N_11104,N_6688,N_5243);
nand U11105 (N_11105,N_7352,N_5154);
and U11106 (N_11106,N_7576,N_9669);
and U11107 (N_11107,N_9809,N_6469);
nor U11108 (N_11108,N_8623,N_7132);
nor U11109 (N_11109,N_8643,N_8524);
nand U11110 (N_11110,N_8495,N_5676);
nand U11111 (N_11111,N_6188,N_7105);
and U11112 (N_11112,N_5753,N_6972);
nand U11113 (N_11113,N_6624,N_5296);
or U11114 (N_11114,N_7251,N_9711);
nand U11115 (N_11115,N_5884,N_5681);
nor U11116 (N_11116,N_6847,N_8792);
nor U11117 (N_11117,N_5650,N_5267);
or U11118 (N_11118,N_9325,N_8248);
nor U11119 (N_11119,N_8530,N_7339);
nor U11120 (N_11120,N_7525,N_8278);
nor U11121 (N_11121,N_6954,N_6174);
or U11122 (N_11122,N_8112,N_5059);
or U11123 (N_11123,N_7598,N_9000);
nand U11124 (N_11124,N_9151,N_9537);
and U11125 (N_11125,N_5992,N_8984);
and U11126 (N_11126,N_8666,N_5253);
or U11127 (N_11127,N_6700,N_8993);
nor U11128 (N_11128,N_5769,N_8434);
nand U11129 (N_11129,N_9133,N_8023);
and U11130 (N_11130,N_8276,N_8037);
nor U11131 (N_11131,N_9639,N_5738);
nor U11132 (N_11132,N_7741,N_9887);
and U11133 (N_11133,N_8839,N_9623);
nor U11134 (N_11134,N_7644,N_9974);
nor U11135 (N_11135,N_5137,N_5415);
or U11136 (N_11136,N_6645,N_7697);
nand U11137 (N_11137,N_5880,N_8760);
nor U11138 (N_11138,N_6846,N_8477);
nor U11139 (N_11139,N_6888,N_7027);
and U11140 (N_11140,N_8565,N_9501);
and U11141 (N_11141,N_8613,N_5284);
or U11142 (N_11142,N_8698,N_6111);
nor U11143 (N_11143,N_5679,N_6352);
nand U11144 (N_11144,N_9874,N_7599);
or U11145 (N_11145,N_6457,N_6353);
xor U11146 (N_11146,N_8425,N_6213);
and U11147 (N_11147,N_8001,N_9773);
nand U11148 (N_11148,N_9806,N_8915);
and U11149 (N_11149,N_5798,N_7521);
and U11150 (N_11150,N_7377,N_5293);
nor U11151 (N_11151,N_9142,N_5089);
or U11152 (N_11152,N_6680,N_5842);
nor U11153 (N_11153,N_5691,N_8045);
nand U11154 (N_11154,N_6983,N_7445);
nor U11155 (N_11155,N_8751,N_8609);
or U11156 (N_11156,N_8771,N_8894);
nor U11157 (N_11157,N_5487,N_5316);
xor U11158 (N_11158,N_7591,N_5045);
or U11159 (N_11159,N_6109,N_9779);
nor U11160 (N_11160,N_7391,N_9046);
nand U11161 (N_11161,N_6917,N_9274);
and U11162 (N_11162,N_7388,N_8146);
nand U11163 (N_11163,N_8650,N_9720);
or U11164 (N_11164,N_9024,N_6305);
nand U11165 (N_11165,N_9109,N_7312);
and U11166 (N_11166,N_8577,N_7856);
and U11167 (N_11167,N_5711,N_6100);
or U11168 (N_11168,N_7633,N_9084);
or U11169 (N_11169,N_9406,N_9395);
xor U11170 (N_11170,N_5891,N_6941);
nor U11171 (N_11171,N_7764,N_8092);
nor U11172 (N_11172,N_7791,N_9643);
and U11173 (N_11173,N_5426,N_7508);
and U11174 (N_11174,N_8311,N_8223);
nand U11175 (N_11175,N_7360,N_6951);
or U11176 (N_11176,N_7406,N_5552);
and U11177 (N_11177,N_6316,N_6635);
nor U11178 (N_11178,N_7662,N_9182);
and U11179 (N_11179,N_8448,N_6267);
nor U11180 (N_11180,N_8602,N_6769);
nor U11181 (N_11181,N_6034,N_9333);
and U11182 (N_11182,N_5040,N_8407);
nor U11183 (N_11183,N_8543,N_8197);
and U11184 (N_11184,N_7208,N_5039);
and U11185 (N_11185,N_8405,N_9368);
nor U11186 (N_11186,N_7600,N_5338);
xnor U11187 (N_11187,N_7702,N_9001);
nor U11188 (N_11188,N_6782,N_5815);
or U11189 (N_11189,N_8848,N_5941);
nor U11190 (N_11190,N_8579,N_6587);
and U11191 (N_11191,N_8653,N_9266);
nor U11192 (N_11192,N_5281,N_9369);
nor U11193 (N_11193,N_7168,N_9941);
nand U11194 (N_11194,N_7005,N_8390);
and U11195 (N_11195,N_6275,N_5231);
or U11196 (N_11196,N_5317,N_8968);
or U11197 (N_11197,N_5828,N_7372);
nand U11198 (N_11198,N_6526,N_7700);
and U11199 (N_11199,N_9446,N_8808);
nand U11200 (N_11200,N_9074,N_9054);
nand U11201 (N_11201,N_6532,N_7876);
nor U11202 (N_11202,N_6849,N_6952);
or U11203 (N_11203,N_7762,N_8305);
nor U11204 (N_11204,N_6070,N_5937);
or U11205 (N_11205,N_7854,N_6950);
xnor U11206 (N_11206,N_9959,N_7815);
nor U11207 (N_11207,N_7756,N_8098);
and U11208 (N_11208,N_8768,N_6258);
or U11209 (N_11209,N_9665,N_7416);
and U11210 (N_11210,N_8657,N_6020);
or U11211 (N_11211,N_8486,N_9090);
or U11212 (N_11212,N_6986,N_7018);
nand U11213 (N_11213,N_9439,N_8066);
and U11214 (N_11214,N_5851,N_7740);
and U11215 (N_11215,N_5578,N_5783);
and U11216 (N_11216,N_9049,N_6162);
nand U11217 (N_11217,N_9948,N_5909);
nand U11218 (N_11218,N_5082,N_5021);
nand U11219 (N_11219,N_9843,N_7872);
nand U11220 (N_11220,N_5495,N_8734);
nor U11221 (N_11221,N_9048,N_7628);
or U11222 (N_11222,N_7003,N_5211);
nand U11223 (N_11223,N_8398,N_9803);
nor U11224 (N_11224,N_7485,N_7224);
or U11225 (N_11225,N_6825,N_7007);
nand U11226 (N_11226,N_5329,N_7184);
nand U11227 (N_11227,N_9062,N_8511);
nand U11228 (N_11228,N_7267,N_9458);
xor U11229 (N_11229,N_8135,N_9002);
or U11230 (N_11230,N_9016,N_7444);
or U11231 (N_11231,N_5391,N_7850);
nand U11232 (N_11232,N_9937,N_6887);
and U11233 (N_11233,N_6802,N_9951);
nand U11234 (N_11234,N_5520,N_9555);
or U11235 (N_11235,N_5374,N_9917);
xor U11236 (N_11236,N_5820,N_6844);
nand U11237 (N_11237,N_8445,N_5446);
xnor U11238 (N_11238,N_8955,N_7545);
and U11239 (N_11239,N_7447,N_8559);
nor U11240 (N_11240,N_6580,N_9256);
nor U11241 (N_11241,N_6876,N_8084);
nor U11242 (N_11242,N_8323,N_6313);
nor U11243 (N_11243,N_9708,N_9107);
nand U11244 (N_11244,N_5544,N_8797);
nor U11245 (N_11245,N_8203,N_6032);
or U11246 (N_11246,N_7695,N_6994);
nor U11247 (N_11247,N_5627,N_6090);
and U11248 (N_11248,N_6816,N_9837);
and U11249 (N_11249,N_8542,N_5974);
and U11250 (N_11250,N_8684,N_7140);
nor U11251 (N_11251,N_6636,N_8343);
nor U11252 (N_11252,N_5708,N_7991);
or U11253 (N_11253,N_6475,N_8820);
and U11254 (N_11254,N_6743,N_5433);
nor U11255 (N_11255,N_8909,N_9618);
nand U11256 (N_11256,N_8360,N_6396);
nand U11257 (N_11257,N_5203,N_9382);
nor U11258 (N_11258,N_5431,N_9802);
nor U11259 (N_11259,N_5079,N_7094);
and U11260 (N_11260,N_6870,N_6840);
nor U11261 (N_11261,N_9481,N_5193);
or U11262 (N_11262,N_9422,N_5146);
or U11263 (N_11263,N_7438,N_8272);
or U11264 (N_11264,N_8246,N_7690);
or U11265 (N_11265,N_6279,N_7075);
or U11266 (N_11266,N_7495,N_6285);
and U11267 (N_11267,N_7476,N_6985);
and U11268 (N_11268,N_7053,N_6639);
or U11269 (N_11269,N_6649,N_8611);
xnor U11270 (N_11270,N_8039,N_7942);
nor U11271 (N_11271,N_7183,N_7719);
nand U11272 (N_11272,N_6075,N_9032);
nand U11273 (N_11273,N_7840,N_7068);
or U11274 (N_11274,N_7450,N_9340);
nor U11275 (N_11275,N_5751,N_7175);
or U11276 (N_11276,N_6282,N_9813);
nor U11277 (N_11277,N_6280,N_5563);
nand U11278 (N_11278,N_5217,N_9933);
nor U11279 (N_11279,N_7563,N_7320);
nand U11280 (N_11280,N_9605,N_9976);
and U11281 (N_11281,N_8175,N_8812);
nor U11282 (N_11282,N_6078,N_5950);
xor U11283 (N_11283,N_6544,N_5392);
nor U11284 (N_11284,N_9531,N_9262);
nor U11285 (N_11285,N_5801,N_6049);
nor U11286 (N_11286,N_7237,N_9880);
and U11287 (N_11287,N_8649,N_6350);
and U11288 (N_11288,N_9160,N_5805);
and U11289 (N_11289,N_6810,N_5328);
nand U11290 (N_11290,N_5459,N_6942);
nand U11291 (N_11291,N_9612,N_8068);
nor U11292 (N_11292,N_9394,N_5920);
nand U11293 (N_11293,N_7106,N_9932);
nand U11294 (N_11294,N_9339,N_8377);
and U11295 (N_11295,N_6920,N_8733);
and U11296 (N_11296,N_8087,N_6839);
or U11297 (N_11297,N_6975,N_8689);
nor U11298 (N_11298,N_5189,N_5500);
nand U11299 (N_11299,N_8297,N_8835);
and U11300 (N_11300,N_5202,N_6914);
or U11301 (N_11301,N_8700,N_6481);
nand U11302 (N_11302,N_7483,N_5197);
nand U11303 (N_11303,N_8549,N_8226);
and U11304 (N_11304,N_6343,N_9695);
nor U11305 (N_11305,N_6621,N_9124);
nor U11306 (N_11306,N_9923,N_5568);
nand U11307 (N_11307,N_6895,N_9772);
and U11308 (N_11308,N_5764,N_9578);
and U11309 (N_11309,N_5906,N_7533);
and U11310 (N_11310,N_6719,N_5848);
or U11311 (N_11311,N_7813,N_5631);
and U11312 (N_11312,N_6803,N_9147);
and U11313 (N_11313,N_8231,N_5540);
nand U11314 (N_11314,N_6541,N_9343);
and U11315 (N_11315,N_6717,N_9367);
or U11316 (N_11316,N_5450,N_7504);
nor U11317 (N_11317,N_6461,N_5693);
nand U11318 (N_11318,N_7045,N_9122);
nand U11319 (N_11319,N_6144,N_8724);
and U11320 (N_11320,N_7665,N_9302);
nand U11321 (N_11321,N_5133,N_7825);
and U11322 (N_11322,N_9840,N_8767);
nor U11323 (N_11323,N_5725,N_5830);
nand U11324 (N_11324,N_7304,N_5168);
nand U11325 (N_11325,N_5295,N_5344);
and U11326 (N_11326,N_8506,N_7350);
or U11327 (N_11327,N_5995,N_6315);
nand U11328 (N_11328,N_7499,N_9753);
nand U11329 (N_11329,N_9465,N_5703);
and U11330 (N_11330,N_9288,N_6783);
nor U11331 (N_11331,N_6509,N_7909);
xor U11332 (N_11332,N_5634,N_7964);
nand U11333 (N_11333,N_9009,N_6368);
nand U11334 (N_11334,N_7648,N_6433);
nor U11335 (N_11335,N_9759,N_8913);
nand U11336 (N_11336,N_9871,N_8351);
nor U11337 (N_11337,N_7205,N_5541);
nor U11338 (N_11338,N_5238,N_6222);
and U11339 (N_11339,N_6194,N_6756);
nand U11340 (N_11340,N_5685,N_7097);
nor U11341 (N_11341,N_9229,N_7421);
nand U11342 (N_11342,N_7153,N_8660);
nand U11343 (N_11343,N_8631,N_7838);
or U11344 (N_11344,N_8170,N_8416);
nand U11345 (N_11345,N_5565,N_6918);
and U11346 (N_11346,N_7265,N_7661);
nand U11347 (N_11347,N_9511,N_6705);
nand U11348 (N_11348,N_8111,N_8628);
and U11349 (N_11349,N_9797,N_7674);
or U11350 (N_11350,N_9373,N_7866);
nand U11351 (N_11351,N_8499,N_6307);
and U11352 (N_11352,N_6225,N_7620);
or U11353 (N_11353,N_5482,N_8438);
nand U11354 (N_11354,N_5734,N_8450);
and U11355 (N_11355,N_9899,N_6881);
xor U11356 (N_11356,N_8564,N_5773);
and U11357 (N_11357,N_7289,N_7475);
nand U11358 (N_11358,N_9811,N_8041);
nor U11359 (N_11359,N_7107,N_8167);
and U11360 (N_11360,N_9355,N_9418);
and U11361 (N_11361,N_7210,N_9784);
nor U11362 (N_11362,N_8948,N_9535);
nor U11363 (N_11363,N_7774,N_8825);
nor U11364 (N_11364,N_6977,N_5774);
nand U11365 (N_11365,N_7126,N_5241);
nand U11366 (N_11366,N_6296,N_9575);
nor U11367 (N_11367,N_8030,N_5618);
and U11368 (N_11368,N_7892,N_9769);
nand U11369 (N_11369,N_9249,N_7585);
nor U11370 (N_11370,N_5981,N_9627);
and U11371 (N_11371,N_6051,N_6263);
nor U11372 (N_11372,N_9253,N_6030);
nor U11373 (N_11373,N_9284,N_6370);
and U11374 (N_11374,N_7271,N_8227);
nor U11375 (N_11375,N_8106,N_5905);
nand U11376 (N_11376,N_7603,N_8270);
and U11377 (N_11377,N_7077,N_8128);
nor U11378 (N_11378,N_7319,N_6770);
nor U11379 (N_11379,N_6424,N_7565);
nand U11380 (N_11380,N_9461,N_7796);
or U11381 (N_11381,N_9670,N_6269);
or U11382 (N_11382,N_5781,N_5440);
nor U11383 (N_11383,N_8882,N_7711);
or U11384 (N_11384,N_8286,N_8451);
or U11385 (N_11385,N_7082,N_9171);
xnor U11386 (N_11386,N_9865,N_5001);
or U11387 (N_11387,N_5591,N_7976);
nor U11388 (N_11388,N_9705,N_7370);
or U11389 (N_11389,N_5013,N_6165);
and U11390 (N_11390,N_9491,N_8921);
nor U11391 (N_11391,N_5185,N_6298);
and U11392 (N_11392,N_8895,N_7624);
and U11393 (N_11393,N_6379,N_7033);
or U11394 (N_11394,N_8132,N_8505);
or U11395 (N_11395,N_6750,N_6131);
nor U11396 (N_11396,N_8555,N_5935);
and U11397 (N_11397,N_5870,N_7385);
and U11398 (N_11398,N_6428,N_8184);
and U11399 (N_11399,N_7248,N_8216);
and U11400 (N_11400,N_8959,N_7507);
nand U11401 (N_11401,N_9795,N_9091);
or U11402 (N_11402,N_6582,N_5918);
or U11403 (N_11403,N_9169,N_8986);
nor U11404 (N_11404,N_8133,N_8585);
or U11405 (N_11405,N_6542,N_8637);
nand U11406 (N_11406,N_7396,N_8293);
nand U11407 (N_11407,N_7619,N_5856);
and U11408 (N_11408,N_9819,N_5827);
xor U11409 (N_11409,N_6620,N_8591);
or U11410 (N_11410,N_6397,N_5893);
nor U11411 (N_11411,N_6426,N_5525);
nand U11412 (N_11412,N_6650,N_8011);
nor U11413 (N_11413,N_9352,N_8662);
or U11414 (N_11414,N_5969,N_7502);
or U11415 (N_11415,N_7968,N_5803);
and U11416 (N_11416,N_7379,N_7425);
nand U11417 (N_11417,N_7044,N_7770);
xor U11418 (N_11418,N_7997,N_5854);
and U11419 (N_11419,N_7063,N_8697);
or U11420 (N_11420,N_6940,N_5364);
xor U11421 (N_11421,N_8291,N_6552);
and U11422 (N_11422,N_6036,N_7178);
xnor U11423 (N_11423,N_5983,N_7424);
nand U11424 (N_11424,N_5957,N_9413);
or U11425 (N_11425,N_6415,N_7110);
and U11426 (N_11426,N_5085,N_8391);
xnor U11427 (N_11427,N_7927,N_5366);
or U11428 (N_11428,N_7405,N_7151);
nor U11429 (N_11429,N_7279,N_6152);
nand U11430 (N_11430,N_7235,N_5215);
and U11431 (N_11431,N_7891,N_8401);
xor U11432 (N_11432,N_8916,N_6793);
or U11433 (N_11433,N_7763,N_8299);
and U11434 (N_11434,N_6721,N_6531);
or U11435 (N_11435,N_9649,N_8945);
nor U11436 (N_11436,N_8742,N_7780);
nor U11437 (N_11437,N_9387,N_6610);
nor U11438 (N_11438,N_7731,N_6234);
or U11439 (N_11439,N_8872,N_5382);
nor U11440 (N_11440,N_8382,N_7734);
nand U11441 (N_11441,N_9648,N_5862);
and U11442 (N_11442,N_5655,N_8874);
and U11443 (N_11443,N_5246,N_9297);
nand U11444 (N_11444,N_8036,N_7411);
xnor U11445 (N_11445,N_9716,N_6960);
nor U11446 (N_11446,N_6512,N_8046);
nand U11447 (N_11447,N_8720,N_6765);
nor U11448 (N_11448,N_6679,N_6251);
nand U11449 (N_11449,N_6677,N_7111);
nand U11450 (N_11450,N_9075,N_8576);
xor U11451 (N_11451,N_6244,N_8899);
nor U11452 (N_11452,N_8583,N_5671);
and U11453 (N_11453,N_7707,N_5357);
nand U11454 (N_11454,N_8053,N_8599);
nand U11455 (N_11455,N_7912,N_5968);
nand U11456 (N_11456,N_8435,N_8630);
nand U11457 (N_11457,N_7778,N_6465);
nor U11458 (N_11458,N_9348,N_7297);
nor U11459 (N_11459,N_8805,N_6626);
or U11460 (N_11460,N_5804,N_8687);
nand U11461 (N_11461,N_7658,N_7322);
nand U11462 (N_11462,N_7429,N_7789);
nand U11463 (N_11463,N_9066,N_8275);
nand U11464 (N_11464,N_8404,N_8027);
nand U11465 (N_11465,N_5625,N_7797);
and U11466 (N_11466,N_5251,N_5358);
nor U11467 (N_11467,N_9903,N_8987);
and U11468 (N_11468,N_9378,N_5287);
nand U11469 (N_11469,N_6533,N_5776);
and U11470 (N_11470,N_7574,N_6080);
nor U11471 (N_11471,N_6464,N_7904);
and U11472 (N_11472,N_5279,N_7004);
and U11473 (N_11473,N_8209,N_6321);
nand U11474 (N_11474,N_8971,N_7958);
or U11475 (N_11475,N_7006,N_8461);
and U11476 (N_11476,N_5326,N_6281);
and U11477 (N_11477,N_5916,N_5879);
and U11478 (N_11478,N_8386,N_5304);
nand U11479 (N_11479,N_7587,N_8926);
nand U11480 (N_11480,N_7233,N_8562);
nand U11481 (N_11481,N_7034,N_5032);
and U11482 (N_11482,N_5334,N_5566);
nand U11483 (N_11483,N_9093,N_8490);
and U11484 (N_11484,N_5871,N_9085);
nand U11485 (N_11485,N_8003,N_9692);
and U11486 (N_11486,N_8553,N_8595);
nand U11487 (N_11487,N_8852,N_8819);
nand U11488 (N_11488,N_6454,N_9822);
nand U11489 (N_11489,N_5933,N_7480);
nor U11490 (N_11490,N_7412,N_6471);
and U11491 (N_11491,N_9821,N_5361);
nand U11492 (N_11492,N_9588,N_6045);
or U11493 (N_11493,N_8957,N_6113);
nor U11494 (N_11494,N_8536,N_5008);
nor U11495 (N_11495,N_7058,N_9239);
nor U11496 (N_11496,N_6830,N_6928);
and U11497 (N_11497,N_5103,N_9384);
nor U11498 (N_11498,N_5930,N_9831);
and U11499 (N_11499,N_9364,N_5050);
and U11500 (N_11500,N_9057,N_5095);
nor U11501 (N_11501,N_7448,N_8601);
xor U11502 (N_11502,N_9867,N_9021);
nand U11503 (N_11503,N_7641,N_7515);
and U11504 (N_11504,N_6182,N_6858);
and U11505 (N_11505,N_9298,N_9222);
or U11506 (N_11506,N_5235,N_6890);
and U11507 (N_11507,N_6699,N_5418);
or U11508 (N_11508,N_6189,N_6447);
nand U11509 (N_11509,N_8817,N_9190);
nor U11510 (N_11510,N_9319,N_7460);
nor U11511 (N_11511,N_5839,N_6485);
nor U11512 (N_11512,N_5112,N_5550);
xor U11513 (N_11513,N_9468,N_6091);
xor U11514 (N_11514,N_9255,N_9642);
or U11515 (N_11515,N_8749,N_8415);
or U11516 (N_11516,N_6795,N_5029);
and U11517 (N_11517,N_6410,N_5352);
nor U11518 (N_11518,N_9723,N_6641);
nor U11519 (N_11519,N_5797,N_9425);
nand U11520 (N_11520,N_8973,N_9059);
nand U11521 (N_11521,N_5795,N_5635);
nand U11522 (N_11522,N_7569,N_6423);
xor U11523 (N_11523,N_6854,N_6959);
nor U11524 (N_11524,N_9265,N_6273);
or U11525 (N_11525,N_9624,N_5519);
and U11526 (N_11526,N_5266,N_8513);
or U11527 (N_11527,N_9870,N_8029);
and U11528 (N_11528,N_7229,N_7108);
xnor U11529 (N_11529,N_8883,N_7498);
or U11530 (N_11530,N_8057,N_8788);
and U11531 (N_11531,N_6787,N_9138);
nand U11532 (N_11532,N_5213,N_7767);
nor U11533 (N_11533,N_9371,N_6040);
and U11534 (N_11534,N_9485,N_8262);
nand U11535 (N_11535,N_9282,N_7095);
nand U11536 (N_11536,N_9860,N_5787);
nand U11537 (N_11537,N_6073,N_5221);
or U11538 (N_11538,N_7828,N_6832);
or U11539 (N_11539,N_9729,N_7503);
or U11540 (N_11540,N_7557,N_8075);
or U11541 (N_11541,N_8928,N_6094);
or U11542 (N_11542,N_7389,N_7622);
nor U11543 (N_11543,N_6122,N_9466);
nand U11544 (N_11544,N_8605,N_9040);
and U11545 (N_11545,N_8746,N_9322);
or U11546 (N_11546,N_5899,N_6713);
and U11547 (N_11547,N_7593,N_7470);
nor U11548 (N_11548,N_9987,N_8449);
or U11549 (N_11549,N_8224,N_5156);
and U11550 (N_11550,N_6394,N_7214);
nand U11551 (N_11551,N_6516,N_9164);
or U11552 (N_11552,N_5944,N_5979);
nor U11553 (N_11553,N_6684,N_9027);
nor U11554 (N_11554,N_7883,N_6789);
nand U11555 (N_11555,N_9514,N_7431);
nor U11556 (N_11556,N_5714,N_8497);
and U11557 (N_11557,N_6074,N_5470);
or U11558 (N_11558,N_5536,N_9121);
and U11559 (N_11559,N_5665,N_7999);
and U11560 (N_11560,N_7325,N_6595);
or U11561 (N_11561,N_8967,N_8578);
nand U11562 (N_11562,N_7496,N_9905);
nand U11563 (N_11563,N_9633,N_9323);
nor U11564 (N_11564,N_8906,N_9167);
nand U11565 (N_11565,N_7844,N_7085);
nand U11566 (N_11566,N_6924,N_9161);
or U11567 (N_11567,N_5976,N_7056);
and U11568 (N_11568,N_5346,N_8414);
or U11569 (N_11569,N_6949,N_7472);
and U11570 (N_11570,N_5966,N_7008);
nor U11571 (N_11571,N_7983,N_6196);
and U11572 (N_11572,N_5517,N_6682);
or U11573 (N_11573,N_9486,N_5675);
or U11574 (N_11574,N_8065,N_5512);
nor U11575 (N_11575,N_6554,N_7575);
nor U11576 (N_11576,N_9744,N_8208);
nor U11577 (N_11577,N_9707,N_9287);
or U11578 (N_11578,N_8138,N_5489);
and U11579 (N_11579,N_6574,N_8095);
nand U11580 (N_11580,N_7236,N_5240);
and U11581 (N_11581,N_6932,N_9058);
or U11582 (N_11582,N_7345,N_8655);
and U11583 (N_11583,N_7139,N_9681);
or U11584 (N_11584,N_9261,N_6476);
nand U11585 (N_11585,N_7963,N_6330);
nor U11586 (N_11586,N_5140,N_7773);
or U11587 (N_11587,N_6480,N_5327);
nand U11588 (N_11588,N_9607,N_7159);
or U11589 (N_11589,N_8935,N_5183);
nor U11590 (N_11590,N_6933,N_8222);
nand U11591 (N_11591,N_8574,N_5406);
or U11592 (N_11592,N_5624,N_9679);
nor U11593 (N_11593,N_6150,N_5083);
or U11594 (N_11594,N_9755,N_5861);
nor U11595 (N_11595,N_9025,N_8147);
nand U11596 (N_11596,N_8726,N_7663);
nand U11597 (N_11597,N_5350,N_7899);
nand U11598 (N_11598,N_8494,N_8946);
nor U11599 (N_11599,N_9579,N_9228);
and U11600 (N_11600,N_6744,N_9259);
and U11601 (N_11601,N_5031,N_6778);
and U11602 (N_11602,N_7261,N_6939);
nor U11603 (N_11603,N_9029,N_5993);
nor U11604 (N_11604,N_6597,N_8301);
or U11605 (N_11605,N_6405,N_5101);
and U11606 (N_11606,N_5472,N_7898);
or U11607 (N_11607,N_7779,N_6115);
nand U11608 (N_11608,N_9004,N_7768);
nor U11609 (N_11609,N_9760,N_6989);
nor U11610 (N_11610,N_9862,N_9326);
or U11611 (N_11611,N_5956,N_8757);
nand U11612 (N_11612,N_9889,N_9008);
xnor U11613 (N_11613,N_6671,N_8765);
and U11614 (N_11614,N_5551,N_5958);
or U11615 (N_11615,N_5381,N_5961);
nand U11616 (N_11616,N_9949,N_9112);
and U11617 (N_11617,N_7888,N_7992);
nor U11618 (N_11618,N_5018,N_7929);
or U11619 (N_11619,N_5701,N_7433);
or U11620 (N_11620,N_6181,N_5901);
nor U11621 (N_11621,N_7031,N_5926);
or U11622 (N_11622,N_7127,N_8800);
and U11623 (N_11623,N_7017,N_5645);
nor U11624 (N_11624,N_9100,N_8493);
and U11625 (N_11625,N_9572,N_8773);
nand U11626 (N_11626,N_6120,N_5359);
nor U11627 (N_11627,N_7748,N_7698);
nand U11628 (N_11628,N_9515,N_5822);
nor U11629 (N_11629,N_5299,N_8548);
or U11630 (N_11630,N_9365,N_7785);
nor U11631 (N_11631,N_7128,N_8558);
nand U11632 (N_11632,N_9189,N_7713);
xnor U11633 (N_11633,N_5837,N_9532);
nor U11634 (N_11634,N_9502,N_8381);
nor U11635 (N_11635,N_5308,N_6815);
or U11636 (N_11636,N_7712,N_7704);
nor U11637 (N_11637,N_7584,N_6384);
and U11638 (N_11638,N_8102,N_6947);
and U11639 (N_11639,N_8974,N_7050);
nand U11640 (N_11640,N_7895,N_9235);
and U11641 (N_11641,N_8005,N_5562);
nand U11642 (N_11642,N_9397,N_6173);
or U11643 (N_11643,N_5668,N_5128);
nand U11644 (N_11644,N_5179,N_8924);
nor U11645 (N_11645,N_9562,N_5402);
nand U11646 (N_11646,N_7401,N_7614);
or U11647 (N_11647,N_6323,N_5437);
or U11648 (N_11648,N_7682,N_9558);
xnor U11649 (N_11649,N_5412,N_6537);
or U11650 (N_11650,N_9438,N_5332);
nand U11651 (N_11651,N_8645,N_8777);
or U11652 (N_11652,N_6123,N_9361);
nor U11653 (N_11653,N_9306,N_5824);
and U11654 (N_11654,N_7459,N_5840);
nor U11655 (N_11655,N_9982,N_8336);
nand U11656 (N_11656,N_5115,N_8152);
or U11657 (N_11657,N_6910,N_5169);
or U11658 (N_11658,N_6127,N_6436);
xnor U11659 (N_11659,N_8811,N_8743);
nor U11660 (N_11660,N_6818,N_9919);
or U11661 (N_11661,N_6412,N_5997);
nor U11662 (N_11662,N_7419,N_8459);
or U11663 (N_11663,N_6927,N_8441);
or U11664 (N_11664,N_7492,N_6735);
nor U11665 (N_11665,N_5855,N_7417);
xor U11666 (N_11666,N_7692,N_8141);
or U11667 (N_11667,N_9197,N_5915);
nand U11668 (N_11668,N_9792,N_9872);
nor U11669 (N_11669,N_7755,N_9894);
nor U11670 (N_11670,N_6326,N_5780);
nor U11671 (N_11671,N_7020,N_8444);
or U11672 (N_11672,N_5067,N_9173);
and U11673 (N_11673,N_9594,N_9103);
and U11674 (N_11674,N_5971,N_9751);
nand U11675 (N_11675,N_6317,N_8006);
nand U11676 (N_11676,N_5736,N_5385);
nor U11677 (N_11677,N_5744,N_8594);
xnor U11678 (N_11678,N_5485,N_6948);
nor U11679 (N_11679,N_8517,N_5648);
nor U11680 (N_11680,N_9519,N_9965);
nor U11681 (N_11681,N_7995,N_6442);
nand U11682 (N_11682,N_8885,N_5509);
nand U11683 (N_11683,N_5196,N_8779);
and U11684 (N_11684,N_6259,N_6441);
nor U11685 (N_11685,N_5610,N_7367);
and U11686 (N_11686,N_9240,N_9194);
or U11687 (N_11687,N_9584,N_9900);
nor U11688 (N_11688,N_6600,N_9565);
and U11689 (N_11689,N_5455,N_9968);
nand U11690 (N_11690,N_9192,N_8155);
nor U11691 (N_11691,N_7138,N_8680);
nand U11692 (N_11692,N_9503,N_7795);
nor U11693 (N_11693,N_9660,N_8538);
nand U11694 (N_11694,N_9984,N_8723);
nor U11695 (N_11695,N_9241,N_8702);
nor U11696 (N_11696,N_8034,N_6646);
nor U11697 (N_11697,N_8399,N_7086);
and U11698 (N_11698,N_6511,N_9957);
or U11699 (N_11699,N_7451,N_7344);
and U11700 (N_11700,N_5276,N_6995);
or U11701 (N_11701,N_8481,N_8428);
and U11702 (N_11702,N_5505,N_8340);
and U11703 (N_11703,N_8250,N_6822);
and U11704 (N_11704,N_8722,N_5462);
or U11705 (N_11705,N_5198,N_7826);
nor U11706 (N_11706,N_6365,N_9498);
and U11707 (N_11707,N_6731,N_6740);
nor U11708 (N_11708,N_7811,N_8115);
and U11709 (N_11709,N_5790,N_7527);
and U11710 (N_11710,N_6061,N_8031);
and U11711 (N_11711,N_9728,N_6661);
nand U11712 (N_11712,N_5697,N_9006);
and U11713 (N_11713,N_8795,N_6936);
nor U11714 (N_11714,N_5224,N_5144);
and U11715 (N_11715,N_6824,N_9277);
or U11716 (N_11716,N_5965,N_9765);
and U11717 (N_11717,N_9443,N_6551);
or U11718 (N_11718,N_5074,N_5869);
nand U11719 (N_11719,N_9111,N_7853);
or U11720 (N_11720,N_6233,N_6640);
or U11721 (N_11721,N_7629,N_8902);
or U11722 (N_11722,N_6252,N_8500);
nand U11723 (N_11723,N_5262,N_5546);
nor U11724 (N_11724,N_6913,N_8972);
nor U11725 (N_11725,N_6961,N_7418);
and U11726 (N_11726,N_7522,N_5104);
or U11727 (N_11727,N_7986,N_8198);
or U11728 (N_11728,N_8557,N_5268);
and U11729 (N_11729,N_8163,N_5796);
nor U11730 (N_11730,N_8090,N_5609);
and U11731 (N_11731,N_5315,N_5401);
nand U11732 (N_11732,N_7834,N_6515);
nand U11733 (N_11733,N_5208,N_6087);
or U11734 (N_11734,N_5053,N_7338);
and U11735 (N_11735,N_7143,N_5866);
nand U11736 (N_11736,N_7332,N_5532);
and U11737 (N_11737,N_7309,N_6979);
nand U11738 (N_11738,N_6938,N_9972);
nand U11739 (N_11739,N_5161,N_6871);
and U11740 (N_11740,N_5605,N_7238);
nor U11741 (N_11741,N_9042,N_8488);
nor U11742 (N_11742,N_6033,N_7263);
or U11743 (N_11743,N_7775,N_5409);
and U11744 (N_11744,N_5456,N_7296);
or U11745 (N_11745,N_5017,N_9013);
nor U11746 (N_11746,N_7837,N_9118);
nor U11747 (N_11747,N_5157,N_9736);
and U11748 (N_11748,N_6502,N_8162);
and U11749 (N_11749,N_8737,N_9341);
and U11750 (N_11750,N_8004,N_9694);
nand U11751 (N_11751,N_8281,N_7701);
nor U11752 (N_11752,N_6272,N_8365);
and U11753 (N_11753,N_8028,N_7920);
or U11754 (N_11754,N_6339,N_8273);
nor U11755 (N_11755,N_5153,N_8714);
nand U11756 (N_11756,N_6880,N_8319);
nand U11757 (N_11757,N_8498,N_6659);
or U11758 (N_11758,N_5214,N_5209);
nand U11759 (N_11759,N_8422,N_7172);
nand U11760 (N_11760,N_5967,N_6208);
nor U11761 (N_11761,N_5218,N_5599);
and U11762 (N_11762,N_6519,N_9824);
and U11763 (N_11763,N_5674,N_9961);
or U11764 (N_11764,N_5442,N_6681);
nand U11765 (N_11765,N_6217,N_7812);
nor U11766 (N_11766,N_8509,N_9334);
or U11767 (N_11767,N_6179,N_5963);
nor U11768 (N_11768,N_6104,N_6419);
or U11769 (N_11769,N_9593,N_6166);
or U11770 (N_11770,N_9598,N_5932);
nor U11771 (N_11771,N_5009,N_9817);
nor U11772 (N_11772,N_6043,N_9506);
or U11773 (N_11773,N_6638,N_7481);
nor U11774 (N_11774,N_7343,N_6060);
nand U11775 (N_11775,N_7561,N_6997);
or U11776 (N_11776,N_7355,N_5573);
and U11777 (N_11777,N_7586,N_9613);
or U11778 (N_11778,N_6963,N_9257);
xnor U11779 (N_11779,N_8541,N_7365);
nand U11780 (N_11780,N_9268,N_6882);
nand U11781 (N_11781,N_6602,N_9347);
nor U11782 (N_11782,N_8963,N_6374);
and U11783 (N_11783,N_6678,N_6565);
or U11784 (N_11784,N_5938,N_5302);
nor U11785 (N_11785,N_9591,N_6875);
nand U11786 (N_11786,N_8638,N_6297);
nand U11787 (N_11787,N_8600,N_9018);
nor U11788 (N_11788,N_6337,N_9500);
nor U11789 (N_11789,N_5669,N_7040);
nor U11790 (N_11790,N_8829,N_5180);
or U11791 (N_11791,N_8853,N_7659);
and U11792 (N_11792,N_6774,N_6137);
or U11793 (N_11793,N_6311,N_7124);
nor U11794 (N_11794,N_7743,N_9177);
nand U11795 (N_11795,N_7534,N_5467);
nor U11796 (N_11796,N_7595,N_6837);
nor U11797 (N_11797,N_5825,N_6693);
or U11798 (N_11798,N_9810,N_6965);
nor U11799 (N_11799,N_5831,N_6703);
xor U11800 (N_11800,N_6351,N_6925);
nor U11801 (N_11801,N_5623,N_8528);
and U11802 (N_11802,N_6226,N_7931);
and U11803 (N_11803,N_8137,N_9270);
or U11804 (N_11804,N_9619,N_9219);
and U11805 (N_11805,N_6538,N_8471);
nor U11806 (N_11806,N_6559,N_8484);
or U11807 (N_11807,N_7093,N_8458);
nand U11808 (N_11808,N_9358,N_5991);
or U11809 (N_11809,N_8841,N_8124);
nor U11810 (N_11810,N_9640,N_5724);
nand U11811 (N_11811,N_9396,N_7642);
nor U11812 (N_11812,N_9659,N_6019);
and U11813 (N_11813,N_6026,N_5720);
and U11814 (N_11814,N_5471,N_9625);
and U11815 (N_11815,N_8758,N_5949);
and U11816 (N_11816,N_7671,N_7226);
or U11817 (N_11817,N_7919,N_8357);
and U11818 (N_11818,N_9195,N_9962);
and U11819 (N_11819,N_5658,N_9673);
nor U11820 (N_11820,N_7890,N_6829);
and U11821 (N_11821,N_5479,N_8076);
nand U11822 (N_11822,N_8439,N_5680);
and U11823 (N_11823,N_9391,N_7636);
or U11824 (N_11824,N_6667,N_6601);
nand U11825 (N_11825,N_6527,N_5136);
or U11826 (N_11826,N_5730,N_6443);
nor U11827 (N_11827,N_8533,N_7243);
and U11828 (N_11828,N_5036,N_5917);
nor U11829 (N_11829,N_7654,N_7757);
or U11830 (N_11830,N_8621,N_5775);
and U11831 (N_11831,N_6589,N_6969);
or U11832 (N_11832,N_7194,N_6669);
and U11833 (N_11833,N_9129,N_9913);
and U11834 (N_11834,N_5256,N_5809);
nand U11835 (N_11835,N_9017,N_5619);
or U11836 (N_11836,N_9214,N_7937);
or U11837 (N_11837,N_9697,N_8761);
nor U11838 (N_11838,N_7577,N_9293);
or U11839 (N_11839,N_7336,N_6971);
and U11840 (N_11840,N_7524,N_5677);
nand U11841 (N_11841,N_6686,N_6398);
nand U11842 (N_11842,N_5526,N_6593);
nand U11843 (N_11843,N_5373,N_8942);
nand U11844 (N_11844,N_7736,N_5882);
nand U11845 (N_11845,N_6904,N_7631);
xnor U11846 (N_11846,N_5558,N_5110);
or U11847 (N_11847,N_9200,N_7716);
or U11848 (N_11848,N_8093,N_7318);
or U11849 (N_11849,N_8372,N_6710);
or U11850 (N_11850,N_9223,N_7057);
and U11851 (N_11851,N_5425,N_8063);
and U11852 (N_11852,N_7514,N_7938);
and U11853 (N_11853,N_9281,N_9442);
nor U11854 (N_11854,N_6157,N_9472);
nor U11855 (N_11855,N_7197,N_9685);
and U11856 (N_11856,N_7735,N_9337);
and U11857 (N_11857,N_5570,N_7868);
nor U11858 (N_11858,N_7000,N_9448);
xnor U11859 (N_11859,N_6207,N_8738);
and U11860 (N_11860,N_8260,N_9312);
nor U11861 (N_11861,N_7972,N_8385);
and U11862 (N_11862,N_5171,N_9548);
nand U11863 (N_11863,N_9582,N_5731);
and U11864 (N_11864,N_9139,N_9185);
and U11865 (N_11865,N_5343,N_9489);
nor U11866 (N_11866,N_8026,N_9345);
and U11867 (N_11867,N_9428,N_6842);
or U11868 (N_11868,N_6728,N_8110);
nor U11869 (N_11869,N_9721,N_7125);
nor U11870 (N_11870,N_7443,N_6437);
or U11871 (N_11871,N_8603,N_6943);
nand U11872 (N_11872,N_6508,N_7867);
nor U11873 (N_11873,N_7435,N_6496);
nor U11874 (N_11874,N_7616,N_5283);
nor U11875 (N_11875,N_7252,N_5261);
or U11876 (N_11876,N_5474,N_7349);
nor U11877 (N_11877,N_9076,N_9895);
or U11878 (N_11878,N_5684,N_7165);
nand U11879 (N_11879,N_5131,N_8878);
nand U11880 (N_11880,N_5139,N_8845);
nand U11881 (N_11881,N_7393,N_5477);
or U11882 (N_11882,N_7478,N_8713);
or U11883 (N_11883,N_7928,N_9064);
or U11884 (N_11884,N_9068,N_6451);
and U11885 (N_11885,N_7358,N_7255);
or U11886 (N_11886,N_7477,N_8234);
and U11887 (N_11887,N_5205,N_9331);
or U11888 (N_11888,N_8625,N_9317);
nor U11889 (N_11889,N_6974,N_9244);
and U11890 (N_11890,N_7440,N_8586);
and U11891 (N_11891,N_8419,N_8322);
or U11892 (N_11892,N_9206,N_7284);
xnor U11893 (N_11893,N_9788,N_9675);
nor U11894 (N_11894,N_5845,N_5010);
nor U11895 (N_11895,N_8675,N_5216);
and U11896 (N_11896,N_8188,N_9897);
or U11897 (N_11897,N_6907,N_6651);
or U11898 (N_11898,N_8876,N_5617);
nand U11899 (N_11899,N_6068,N_6899);
and U11900 (N_11900,N_9604,N_9727);
nor U11901 (N_11901,N_5451,N_9915);
or U11902 (N_11902,N_9858,N_9154);
nand U11903 (N_11903,N_9696,N_7290);
and U11904 (N_11904,N_8157,N_8120);
nor U11905 (N_11905,N_6632,N_7553);
nand U11906 (N_11906,N_5516,N_9622);
nor U11907 (N_11907,N_9072,N_9097);
and U11908 (N_11908,N_6560,N_6727);
nor U11909 (N_11909,N_9741,N_8355);
or U11910 (N_11910,N_6777,N_6766);
nor U11911 (N_11911,N_7380,N_9672);
nand U11912 (N_11912,N_8616,N_7441);
nor U11913 (N_11913,N_5875,N_6010);
and U11914 (N_11914,N_9600,N_9043);
and U11915 (N_11915,N_7977,N_7368);
xor U11916 (N_11916,N_9303,N_5543);
nor U11917 (N_11917,N_8082,N_8144);
xor U11918 (N_11918,N_7649,N_8253);
nand U11919 (N_11919,N_9896,N_6726);
and U11920 (N_11920,N_9836,N_7306);
and U11921 (N_11921,N_8148,N_7043);
nand U11922 (N_11922,N_8085,N_7340);
nand U11923 (N_11923,N_6239,N_6604);
or U11924 (N_11924,N_8235,N_8730);
and U11925 (N_11925,N_9083,N_9092);
or U11926 (N_11926,N_6930,N_8159);
nand U11927 (N_11927,N_7104,N_9544);
and U11928 (N_11928,N_8941,N_8778);
or U11929 (N_11929,N_5542,N_6432);
or U11930 (N_11930,N_9457,N_5410);
nand U11931 (N_11931,N_8168,N_7948);
or U11932 (N_11932,N_8682,N_8502);
xor U11933 (N_11933,N_7308,N_9450);
or U11934 (N_11934,N_8172,N_6853);
nand U11935 (N_11935,N_8802,N_7607);
and U11936 (N_11936,N_9557,N_9732);
and U11937 (N_11937,N_8403,N_7066);
xor U11938 (N_11938,N_7324,N_9460);
and U11939 (N_11939,N_9444,N_6996);
nand U11940 (N_11940,N_6658,N_7941);
and U11941 (N_11941,N_8933,N_5289);
nor U11942 (N_11942,N_9620,N_7259);
nand U11943 (N_11943,N_5310,N_9844);
and U11944 (N_11944,N_9039,N_6874);
or U11945 (N_11945,N_8467,N_7971);
and U11946 (N_11946,N_6274,N_7666);
and U11947 (N_11947,N_5126,N_8507);
or U11948 (N_11948,N_7945,N_5908);
nor U11949 (N_11949,N_6665,N_9787);
or U11950 (N_11950,N_6261,N_5151);
or U11951 (N_11951,N_8356,N_6003);
or U11952 (N_11952,N_7395,N_8827);
and U11953 (N_11953,N_6039,N_6706);
or U11954 (N_11954,N_8931,N_5404);
or U11955 (N_11955,N_8927,N_6210);
nor U11956 (N_11956,N_7847,N_9318);
nand U11957 (N_11957,N_9263,N_7347);
or U11958 (N_11958,N_9606,N_8025);
nand U11959 (N_11959,N_5984,N_6732);
and U11960 (N_11960,N_7739,N_8325);
or U11961 (N_11961,N_9213,N_7900);
or U11962 (N_11962,N_8739,N_8898);
or U11963 (N_11963,N_5454,N_6014);
or U11964 (N_11964,N_5294,N_9534);
or U11965 (N_11965,N_5355,N_5959);
nand U11966 (N_11966,N_8960,N_6209);
nand U11967 (N_11967,N_8298,N_6767);
nand U11968 (N_11968,N_7588,N_6121);
nand U11969 (N_11969,N_9691,N_8483);
xnor U11970 (N_11970,N_7037,N_7564);
or U11971 (N_11971,N_8755,N_5841);
nor U11972 (N_11972,N_6308,N_8575);
nor U11973 (N_11973,N_7933,N_8546);
nand U11974 (N_11974,N_8233,N_6834);
nand U11975 (N_11975,N_9832,N_8787);
nand U11976 (N_11976,N_7461,N_8705);
nand U11977 (N_11977,N_5508,N_6655);
xor U11978 (N_11978,N_9113,N_7220);
or U11979 (N_11979,N_8659,N_9902);
or U11980 (N_11980,N_5473,N_9559);
nand U11981 (N_11981,N_7466,N_7956);
and U11982 (N_11982,N_6841,N_7787);
or U11983 (N_11983,N_8078,N_7488);
and U11984 (N_11984,N_7988,N_9215);
nor U11985 (N_11985,N_9165,N_7001);
xnor U11986 (N_11986,N_7369,N_7685);
or U11987 (N_11987,N_8624,N_8206);
or U11988 (N_11988,N_9893,N_8886);
or U11989 (N_11989,N_5604,N_5340);
or U11990 (N_11990,N_6072,N_6385);
and U11991 (N_11991,N_6248,N_8523);
nand U11992 (N_11992,N_6378,N_8837);
and U11993 (N_11993,N_5533,N_6563);
or U11994 (N_11994,N_5476,N_5336);
nand U11995 (N_11995,N_5989,N_8123);
nand U11996 (N_11996,N_8540,N_9441);
nor U11997 (N_11997,N_9931,N_8610);
or U11998 (N_11998,N_5365,N_6201);
nand U11999 (N_11999,N_6103,N_5041);
nor U12000 (N_12000,N_5484,N_9999);
nor U12001 (N_12001,N_8150,N_6015);
or U12002 (N_12002,N_7667,N_9376);
nand U12003 (N_12003,N_8129,N_5046);
and U12004 (N_12004,N_5863,N_8568);
or U12005 (N_12005,N_8228,N_5633);
nand U12006 (N_12006,N_6523,N_5896);
or U12007 (N_12007,N_5239,N_6018);
or U12008 (N_12008,N_7064,N_8333);
and U12009 (N_12009,N_9493,N_5654);
nand U12010 (N_12010,N_5895,N_7098);
nand U12011 (N_12011,N_9856,N_6529);
or U12012 (N_12012,N_6138,N_9031);
nand U12013 (N_12013,N_8644,N_6637);
nand U12014 (N_12014,N_6490,N_9678);
nor U12015 (N_12015,N_9849,N_7950);
nand U12016 (N_12016,N_9478,N_5331);
nor U12017 (N_12017,N_8938,N_7298);
nand U12018 (N_12018,N_7216,N_9910);
nand U12019 (N_12019,N_7198,N_7342);
and U12020 (N_12020,N_7801,N_7793);
and U12021 (N_12021,N_7809,N_6202);
or U12022 (N_12022,N_7873,N_6583);
nand U12023 (N_12023,N_8647,N_8862);
and U12024 (N_12024,N_8836,N_5504);
and U12025 (N_12025,N_7901,N_5657);
or U12026 (N_12026,N_7836,N_6500);
nand U12027 (N_12027,N_7484,N_6958);
and U12028 (N_12028,N_8016,N_7714);
or U12029 (N_12029,N_6046,N_6324);
and U12030 (N_12030,N_9175,N_9477);
nor U12031 (N_12031,N_8379,N_6905);
or U12032 (N_12032,N_6059,N_6172);
nor U12033 (N_12033,N_7404,N_5696);
and U12034 (N_12034,N_9963,N_8880);
and U12035 (N_12035,N_5659,N_8232);
nand U12036 (N_12036,N_5768,N_9516);
nand U12037 (N_12037,N_7119,N_9776);
or U12038 (N_12038,N_6868,N_7823);
nand U12039 (N_12039,N_9398,N_6753);
or U12040 (N_12040,N_8648,N_7869);
nand U12041 (N_12041,N_8251,N_8992);
nand U12042 (N_12042,N_8447,N_7301);
nor U12043 (N_12043,N_7491,N_8725);
nor U12044 (N_12044,N_8508,N_7055);
nor U12045 (N_12045,N_8918,N_5249);
or U12046 (N_12046,N_9524,N_7761);
or U12047 (N_12047,N_7581,N_5481);
nor U12048 (N_12048,N_6380,N_9146);
or U12049 (N_12049,N_7398,N_6387);
nor U12050 (N_12050,N_7291,N_8547);
or U12051 (N_12051,N_9512,N_6231);
nand U12052 (N_12052,N_5320,N_5300);
nand U12053 (N_12053,N_8791,N_5368);
and U12054 (N_12054,N_7590,N_9936);
nor U12055 (N_12055,N_5695,N_5339);
and U12056 (N_12056,N_9010,N_7012);
and U12057 (N_12057,N_6862,N_5002);
nor U12058 (N_12058,N_8692,N_9034);
nor U12059 (N_12059,N_5342,N_7381);
and U12060 (N_12060,N_6119,N_9003);
nand U12061 (N_12061,N_8259,N_5020);
and U12062 (N_12062,N_6199,N_9231);
nand U12063 (N_12063,N_9781,N_6048);
and U12064 (N_12064,N_6564,N_8362);
or U12065 (N_12065,N_6192,N_9834);
and U12066 (N_12066,N_7566,N_7737);
or U12067 (N_12067,N_9415,N_7783);
and U12068 (N_12068,N_9258,N_7122);
and U12069 (N_12069,N_8315,N_8748);
nand U12070 (N_12070,N_5091,N_7048);
and U12071 (N_12071,N_8387,N_5260);
and U12072 (N_12072,N_6736,N_5004);
nor U12073 (N_12073,N_9892,N_5337);
and U12074 (N_12074,N_8071,N_6569);
nor U12075 (N_12075,N_6195,N_6838);
and U12076 (N_12076,N_5750,N_5923);
and U12077 (N_12077,N_9429,N_5712);
nor U12078 (N_12078,N_5743,N_7875);
or U12079 (N_12079,N_8122,N_8615);
and U12080 (N_12080,N_7400,N_9357);
xnor U12081 (N_12081,N_9350,N_6555);
or U12082 (N_12082,N_7468,N_9653);
nand U12083 (N_12083,N_9245,N_5706);
or U12084 (N_12084,N_9825,N_6912);
or U12085 (N_12085,N_7874,N_7413);
or U12086 (N_12086,N_9309,N_9632);
or U12087 (N_12087,N_6319,N_5278);
or U12088 (N_12088,N_6823,N_7270);
or U12089 (N_12089,N_6863,N_6623);
nand U12090 (N_12090,N_5733,N_6276);
and U12091 (N_12091,N_7225,N_5166);
and U12092 (N_12092,N_5134,N_5273);
and U12093 (N_12093,N_7266,N_6883);
xnor U12094 (N_12094,N_9104,N_5757);
and U12095 (N_12095,N_9561,N_7679);
nand U12096 (N_12096,N_7434,N_5878);
and U12097 (N_12097,N_6487,N_7247);
nand U12098 (N_12098,N_8781,N_7011);
nand U12099 (N_12099,N_5314,N_5349);
nor U12100 (N_12100,N_8677,N_7282);
and U12101 (N_12101,N_9037,N_9746);
nand U12102 (N_12102,N_5003,N_5086);
or U12103 (N_12103,N_8238,N_5513);
and U12104 (N_12104,N_5286,N_6957);
or U12105 (N_12105,N_5593,N_8592);
nand U12106 (N_12106,N_7516,N_5223);
or U12107 (N_12107,N_7232,N_9311);
nor U12108 (N_12108,N_9712,N_8282);
or U12109 (N_12109,N_7378,N_6354);
or U12110 (N_12110,N_9471,N_7422);
or U12111 (N_12111,N_8606,N_9609);
nor U12112 (N_12112,N_5626,N_6763);
and U12113 (N_12113,N_5155,N_9839);
and U12114 (N_12114,N_8217,N_5940);
nor U12115 (N_12115,N_9247,N_7446);
nand U12116 (N_12116,N_6044,N_5206);
and U12117 (N_12117,N_5603,N_8109);
xor U12118 (N_12118,N_9476,N_6521);
nand U12119 (N_12119,N_8061,N_9267);
nor U12120 (N_12120,N_9638,N_6400);
or U12121 (N_12121,N_6372,N_9012);
nor U12122 (N_12122,N_7146,N_7280);
nor U12123 (N_12123,N_8693,N_8866);
nand U12124 (N_12124,N_7807,N_8265);
nor U12125 (N_12125,N_8598,N_9069);
nor U12126 (N_12126,N_5123,N_8683);
nor U12127 (N_12127,N_6518,N_9507);
nor U12128 (N_12128,N_5688,N_7084);
nor U12129 (N_12129,N_5528,N_7547);
nand U12130 (N_12130,N_6937,N_9275);
nor U12131 (N_12131,N_9080,N_6107);
nor U12132 (N_12132,N_9096,N_8593);
or U12133 (N_12133,N_5608,N_7121);
nand U12134 (N_12134,N_7223,N_7640);
or U12135 (N_12135,N_9922,N_6187);
nor U12136 (N_12136,N_6160,N_8943);
nor U12137 (N_12137,N_7283,N_5498);
and U12138 (N_12138,N_8256,N_9980);
and U12139 (N_12139,N_5493,N_9846);
or U12140 (N_12140,N_7207,N_8350);
or U12141 (N_12141,N_8877,N_9798);
nand U12142 (N_12142,N_5867,N_8832);
or U12143 (N_12143,N_9569,N_9700);
nor U12144 (N_12144,N_9349,N_8525);
or U12145 (N_12145,N_8183,N_9022);
nor U12146 (N_12146,N_5756,N_6656);
or U12147 (N_12147,N_7664,N_8321);
nand U12148 (N_12148,N_5174,N_5494);
or U12149 (N_12149,N_6193,N_8879);
and U12150 (N_12150,N_9689,N_6328);
and U12151 (N_12151,N_5399,N_9877);
and U12152 (N_12152,N_7188,N_6742);
nand U12153 (N_12153,N_6205,N_9220);
and U12154 (N_12154,N_6892,N_9738);
and U12155 (N_12155,N_6865,N_6001);
or U12156 (N_12156,N_6962,N_7246);
nor U12157 (N_12157,N_8940,N_5666);
and U12158 (N_12158,N_7181,N_6662);
and U12159 (N_12159,N_7426,N_7635);
or U12160 (N_12160,N_7799,N_6746);
nor U12161 (N_12161,N_8378,N_6176);
and U12162 (N_12162,N_8745,N_8086);
and U12163 (N_12163,N_8772,N_9740);
and U12164 (N_12164,N_8353,N_8033);
nand U12165 (N_12165,N_7915,N_6696);
nand U12166 (N_12166,N_7632,N_7881);
nor U12167 (N_12167,N_9749,N_9985);
nor U12168 (N_12168,N_6573,N_5729);
or U12169 (N_12169,N_7203,N_9038);
and U12170 (N_12170,N_8269,N_6548);
or U12171 (N_12171,N_6973,N_8949);
nor U12172 (N_12172,N_5621,N_8230);
nand U12173 (N_12173,N_8126,N_8936);
and U12174 (N_12174,N_9583,N_5186);
nand U12175 (N_12175,N_7621,N_5135);
nand U12176 (N_12176,N_9254,N_7615);
and U12177 (N_12177,N_7364,N_5990);
xor U12178 (N_12178,N_7822,N_7330);
and U12179 (N_12179,N_8668,N_7542);
or U12180 (N_12180,N_6414,N_9545);
and U12181 (N_12181,N_6007,N_5088);
or U12182 (N_12182,N_9499,N_5792);
nand U12183 (N_12183,N_7326,N_8052);
or U12184 (N_12184,N_9786,N_5836);
and U12185 (N_12185,N_8000,N_7457);
or U12186 (N_12186,N_8520,N_7580);
nand U12187 (N_12187,N_8024,N_8892);
or U12188 (N_12188,N_5874,N_6747);
and U12189 (N_12189,N_6407,N_6953);
nand U12190 (N_12190,N_6629,N_8969);
and U12191 (N_12191,N_6758,N_7335);
nor U12192 (N_12192,N_6473,N_5860);
nor U12193 (N_12193,N_8953,N_6608);
nand U12194 (N_12194,N_8904,N_7258);
nand U12195 (N_12195,N_8328,N_9975);
and U12196 (N_12196,N_9687,N_9953);
and U12197 (N_12197,N_8313,N_9706);
or U12198 (N_12198,N_8861,N_9393);
or U12199 (N_12199,N_9356,N_7217);
and U12200 (N_12200,N_7062,N_7879);
nor U12201 (N_12201,N_5816,N_8279);
or U12202 (N_12202,N_9308,N_9581);
or U12203 (N_12203,N_6715,N_5779);
xnor U12204 (N_12204,N_7918,N_7150);
nor U12205 (N_12205,N_5182,N_9180);
or U12206 (N_12206,N_6017,N_8752);
nand U12207 (N_12207,N_7647,N_7035);
or U12208 (N_12208,N_7655,N_7852);
nand U12209 (N_12209,N_7273,N_8295);
or U12210 (N_12210,N_6873,N_7022);
nor U12211 (N_12211,N_6497,N_7924);
or U12212 (N_12212,N_7453,N_9800);
nand U12213 (N_12213,N_7625,N_5458);
and U12214 (N_12214,N_6145,N_8193);
xor U12215 (N_12215,N_5955,N_5419);
nor U12216 (N_12216,N_8040,N_7969);
nor U12217 (N_12217,N_9504,N_7078);
nand U12218 (N_12218,N_6692,N_8999);
or U12219 (N_12219,N_8950,N_5465);
or U12220 (N_12220,N_5178,N_6993);
or U12221 (N_12221,N_9539,N_5333);
nor U12222 (N_12222,N_9914,N_8930);
and U12223 (N_12223,N_7532,N_9310);
or U12224 (N_12224,N_6826,N_9041);
and U12225 (N_12225,N_9521,N_9563);
nand U12226 (N_12226,N_5759,N_7474);
nand U12227 (N_12227,N_8696,N_8903);
nand U12228 (N_12228,N_7560,N_6866);
nor U12229 (N_12229,N_6780,N_5770);
nand U12230 (N_12230,N_6775,N_8776);
and U12231 (N_12231,N_8908,N_7333);
or U12232 (N_12232,N_9966,N_5615);
or U12233 (N_12233,N_5782,N_6095);
or U12234 (N_12234,N_8475,N_8641);
nand U12235 (N_12235,N_8824,N_8833);
nand U12236 (N_12236,N_9630,N_8856);
nor U12237 (N_12237,N_7190,N_9754);
and U12238 (N_12238,N_7382,N_5794);
nor U12239 (N_12239,N_7479,N_5075);
nand U12240 (N_12240,N_6434,N_9078);
nand U12241 (N_12241,N_6341,N_8241);
nor U12242 (N_12242,N_7113,N_7857);
nand U12243 (N_12243,N_5483,N_7528);
nor U12244 (N_12244,N_8635,N_8721);
or U12245 (N_12245,N_9611,N_5242);
nor U12246 (N_12246,N_6312,N_9767);
nor U12247 (N_12247,N_6369,N_7902);
and U12248 (N_12248,N_9553,N_5632);
and U12249 (N_12249,N_8153,N_7646);
or U12250 (N_12250,N_5572,N_5130);
nor U12251 (N_12251,N_7287,N_5556);
nand U12252 (N_12252,N_5692,N_8400);
nor U12253 (N_12253,N_5964,N_9470);
nand U12254 (N_12254,N_5707,N_9385);
nand U12255 (N_12255,N_5994,N_8646);
nor U12256 (N_12256,N_6652,N_9823);
nor U12257 (N_12257,N_6086,N_7860);
nor U12258 (N_12258,N_5924,N_5503);
nor U12259 (N_12259,N_6657,N_9768);
nor U12260 (N_12260,N_5833,N_8674);
or U12261 (N_12261,N_9023,N_9196);
nor U12262 (N_12262,N_7978,N_6484);
nor U12263 (N_12263,N_9136,N_7363);
and U12264 (N_12264,N_7245,N_5269);
and U12265 (N_12265,N_6349,N_7219);
and U12266 (N_12266,N_8142,N_9155);
or U12267 (N_12267,N_5463,N_7788);
nand U12268 (N_12268,N_8324,N_6242);
nor U12269 (N_12269,N_7605,N_6156);
and U12270 (N_12270,N_7222,N_5247);
and U12271 (N_12271,N_8312,N_8014);
or U12272 (N_12272,N_6612,N_5488);
xnor U12273 (N_12273,N_6212,N_9431);
nor U12274 (N_12274,N_6976,N_8937);
nor U12275 (N_12275,N_8537,N_5534);
and U12276 (N_12276,N_7013,N_6809);
or U12277 (N_12277,N_5741,N_7571);
xor U12278 (N_12278,N_9509,N_7771);
or U12279 (N_12279,N_9087,N_7275);
or U12280 (N_12280,N_9462,N_5622);
nand U12281 (N_12281,N_6006,N_5597);
nor U12282 (N_12282,N_9698,N_7293);
nand U12283 (N_12283,N_7501,N_7310);
nand U12284 (N_12284,N_5662,N_5777);
nor U12285 (N_12285,N_5056,N_7550);
nor U12286 (N_12286,N_9978,N_8534);
nor U12287 (N_12287,N_8287,N_5099);
nor U12288 (N_12288,N_5054,N_5042);
nor U12289 (N_12289,N_8920,N_6477);
nand U12290 (N_12290,N_8367,N_7519);
or U12291 (N_12291,N_6277,N_5424);
or U12292 (N_12292,N_5145,N_8701);
and U12293 (N_12293,N_7694,N_7758);
nand U12294 (N_12294,N_9492,N_5389);
nand U12295 (N_12295,N_9209,N_9120);
nor U12296 (N_12296,N_6911,N_7558);
and U12297 (N_12297,N_6591,N_6577);
nand U12298 (N_12298,N_6668,N_6598);
or U12299 (N_12299,N_8474,N_5496);
nor U12300 (N_12300,N_7427,N_6262);
nor U12301 (N_12301,N_8125,N_5647);
or U12302 (N_12302,N_6798,N_8373);
nor U12303 (N_12303,N_6249,N_6254);
and U12304 (N_12304,N_7317,N_5579);
or U12305 (N_12305,N_5229,N_9102);
or U12306 (N_12306,N_7792,N_8844);
or U12307 (N_12307,N_8932,N_8663);
or U12308 (N_12308,N_7212,N_9392);
and U12309 (N_12309,N_7863,N_8462);
or U12310 (N_12310,N_5081,N_7681);
and U12311 (N_12311,N_6256,N_7072);
or U12312 (N_12312,N_6683,N_8478);
nand U12313 (N_12313,N_5181,N_7465);
nor U12314 (N_12314,N_9996,N_9752);
and U12315 (N_12315,N_5447,N_7911);
nor U12316 (N_12316,N_8840,N_9901);
or U12317 (N_12317,N_5742,N_6220);
nand U12318 (N_12318,N_5996,N_5271);
nand U12319 (N_12319,N_6594,N_7691);
and U12320 (N_12320,N_8104,N_9861);
nor U12321 (N_12321,N_7371,N_6998);
nand U12322 (N_12322,N_6171,N_5265);
nor U12323 (N_12323,N_5584,N_9463);
nand U12324 (N_12324,N_9108,N_8457);
or U12325 (N_12325,N_7882,N_8479);
nor U12326 (N_12326,N_8966,N_5192);
nor U12327 (N_12327,N_7487,N_7189);
nand U12328 (N_12328,N_5501,N_7242);
and U12329 (N_12329,N_6178,N_7726);
and U12330 (N_12330,N_8556,N_8074);
nor U12331 (N_12331,N_9852,N_9280);
or U12332 (N_12332,N_5019,N_7845);
and U12333 (N_12333,N_9808,N_9690);
and U12334 (N_12334,N_7830,N_9775);
and U12335 (N_12335,N_7669,N_5596);
nor U12336 (N_12336,N_5852,N_8402);
and U12337 (N_12337,N_8392,N_7782);
nor U12338 (N_12338,N_5164,N_8463);
and U12339 (N_12339,N_7940,N_8717);
and U12340 (N_12340,N_8267,N_9089);
and U12341 (N_12341,N_6470,N_5207);
xor U12342 (N_12342,N_7102,N_8089);
nand U12343 (N_12343,N_8891,N_8059);
and U12344 (N_12344,N_7790,N_9454);
nand U12345 (N_12345,N_6076,N_5876);
nand U12346 (N_12346,N_8437,N_6097);
and U12347 (N_12347,N_6970,N_7573);
and U12348 (N_12348,N_6438,N_9780);
and U12349 (N_12349,N_6439,N_6613);
nor U12350 (N_12350,N_8064,N_8823);
nor U12351 (N_12351,N_5492,N_7039);
and U12352 (N_12352,N_9655,N_8732);
or U12353 (N_12353,N_9855,N_7910);
or U12354 (N_12354,N_9646,N_9587);
and U12355 (N_12355,N_7994,N_5646);
and U12356 (N_12356,N_8813,N_6367);
nor U12357 (N_12357,N_7366,N_6701);
nor U12358 (N_12358,N_8989,N_9432);
or U12359 (N_12359,N_9451,N_5595);
or U12360 (N_12360,N_7408,N_5252);
and U12361 (N_12361,N_8503,N_5405);
nand U12362 (N_12362,N_8083,N_9719);
and U12363 (N_12363,N_6159,N_7677);
and U12364 (N_12364,N_8822,N_9052);
nor U12365 (N_12365,N_9992,N_7612);
nor U12366 (N_12366,N_5303,N_7513);
nand U12367 (N_12367,N_9056,N_6549);
and U12368 (N_12368,N_5788,N_7765);
and U12369 (N_12369,N_6772,N_6440);
and U12370 (N_12370,N_6456,N_8925);
nor U12371 (N_12371,N_6373,N_8956);
nand U12372 (N_12372,N_8589,N_9636);
nand U12373 (N_12373,N_7959,N_8560);
nand U12374 (N_12374,N_6153,N_5678);
nand U12375 (N_12375,N_8304,N_8803);
or U12376 (N_12376,N_6253,N_8121);
nand U12377 (N_12377,N_6053,N_5760);
nor U12378 (N_12378,N_7473,N_6547);
nand U12379 (N_12379,N_9590,N_6915);
or U12380 (N_12380,N_6435,N_6170);
nand U12381 (N_12381,N_8807,N_8664);
xor U12382 (N_12382,N_9114,N_8860);
nor U12383 (N_12383,N_8939,N_6164);
and U12384 (N_12384,N_7186,N_6340);
or U12385 (N_12385,N_8816,N_9212);
nor U12386 (N_12386,N_7939,N_6114);
and U12387 (N_12387,N_8067,N_9324);
nor U12388 (N_12388,N_9550,N_5087);
or U12389 (N_12389,N_9483,N_6666);
nand U12390 (N_12390,N_5978,N_6576);
nor U12391 (N_12391,N_8396,N_6474);
and U12392 (N_12392,N_9907,N_5907);
and U12393 (N_12393,N_5176,N_9528);
nand U12394 (N_12394,N_8140,N_8627);
or U12395 (N_12395,N_7407,N_8117);
or U12396 (N_12396,N_6147,N_6788);
and U12397 (N_12397,N_9156,N_7934);
or U12398 (N_12398,N_8838,N_8243);
or U12399 (N_12399,N_5051,N_7351);
nand U12400 (N_12400,N_5826,N_9954);
and U12401 (N_12401,N_8529,N_8288);
and U12402 (N_12402,N_5977,N_8096);
or U12403 (N_12403,N_9654,N_7390);
and U12404 (N_12404,N_9410,N_6346);
nor U12405 (N_12405,N_8929,N_6240);
nor U12406 (N_12406,N_6660,N_5710);
and U12407 (N_12407,N_9427,N_5354);
nor U12408 (N_12408,N_8418,N_7653);
nand U12409 (N_12409,N_5667,N_7384);
or U12410 (N_12410,N_9916,N_6299);
nor U12411 (N_12411,N_9530,N_8590);
or U12412 (N_12412,N_8736,N_7051);
nand U12413 (N_12413,N_5301,N_7754);
nor U12414 (N_12414,N_6023,N_9851);
nand U12415 (N_12415,N_5900,N_6909);
and U12416 (N_12416,N_6081,N_5849);
and U12417 (N_12417,N_5802,N_6065);
and U12418 (N_12418,N_5607,N_8640);
and U12419 (N_12419,N_6291,N_7650);
nor U12420 (N_12420,N_9285,N_8588);
nor U12421 (N_12421,N_6987,N_9426);
nand U12422 (N_12422,N_5323,N_6186);
nand U12423 (N_12423,N_5120,N_5972);
nor U12424 (N_12424,N_7871,N_5400);
nor U12425 (N_12425,N_7187,N_5006);
nand U12426 (N_12426,N_6180,N_6348);
nand U12427 (N_12427,N_5948,N_9589);
nand U12428 (N_12428,N_5985,N_6616);
and U12429 (N_12429,N_7204,N_6510);
nor U12430 (N_12430,N_9580,N_8454);
or U12431 (N_12431,N_9134,N_5643);
or U12432 (N_12432,N_8622,N_6334);
and U12433 (N_12433,N_7179,N_9943);
or U12434 (N_12434,N_8617,N_8580);
and U12435 (N_12435,N_5748,N_9634);
and U12436 (N_12436,N_9279,N_8782);
and U12437 (N_12437,N_7269,N_9793);
or U12438 (N_12438,N_8656,N_7014);
xor U12439 (N_12439,N_5910,N_9770);
or U12440 (N_12440,N_7509,N_6105);
or U12441 (N_12441,N_7943,N_5388);
nand U12442 (N_12442,N_7383,N_9661);
nand U12443 (N_12443,N_9005,N_8199);
and U12444 (N_12444,N_8440,N_6129);
nand U12445 (N_12445,N_9405,N_5587);
nand U12446 (N_12446,N_6265,N_5765);
and U12447 (N_12447,N_5988,N_6553);
or U12448 (N_12448,N_9473,N_5098);
nor U12449 (N_12449,N_8393,N_5987);
and U12450 (N_12450,N_8604,N_9098);
nor U12451 (N_12451,N_9616,N_6676);
or U12452 (N_12452,N_6644,N_9399);
and U12453 (N_12453,N_8032,N_6493);
or U12454 (N_12454,N_5397,N_7156);
or U12455 (N_12455,N_7529,N_7311);
nor U12456 (N_12456,N_6322,N_9388);
nand U12457 (N_12457,N_7715,N_6411);
and U12458 (N_12458,N_8341,N_7760);
or U12459 (N_12459,N_6062,N_8681);
and U12460 (N_12460,N_7059,N_8165);
and U12461 (N_12461,N_9777,N_8868);
or U12462 (N_12462,N_7946,N_6430);
or U12463 (N_12463,N_9977,N_8164);
and U12464 (N_12464,N_7781,N_8417);
and U12465 (N_12465,N_5811,N_9157);
nor U12466 (N_12466,N_6450,N_9488);
or U12467 (N_12467,N_6867,N_8433);
nand U12468 (N_12468,N_6110,N_5141);
xnor U12469 (N_12469,N_6375,N_5510);
nand U12470 (N_12470,N_8762,N_6092);
and U12471 (N_12471,N_5897,N_7180);
nor U12472 (N_12472,N_6283,N_5427);
nor U12473 (N_12473,N_6134,N_9573);
xor U12474 (N_12474,N_9353,N_8292);
nand U12475 (N_12475,N_6714,N_7827);
nand U12476 (N_12476,N_8870,N_9401);
nor U12477 (N_12477,N_7829,N_5055);
nor U12478 (N_12478,N_8770,N_7777);
or U12479 (N_12479,N_7133,N_8496);
and U12480 (N_12480,N_9335,N_9145);
nor U12481 (N_12481,N_6561,N_6724);
nand U12482 (N_12482,N_9250,N_5432);
or U12483 (N_12483,N_5911,N_8363);
nor U12484 (N_12484,N_9791,N_8007);
nor U12485 (N_12485,N_9891,N_7746);
nor U12486 (N_12486,N_7286,N_7374);
and U12487 (N_12487,N_6148,N_5538);
and U12488 (N_12488,N_6393,N_9662);
or U12489 (N_12489,N_6622,N_7609);
nor U12490 (N_12490,N_6845,N_5636);
nor U12491 (N_12491,N_9656,N_9774);
nor U12492 (N_12492,N_9202,N_8620);
nor U12493 (N_12493,N_5464,N_7009);
nor U12494 (N_12494,N_9141,N_6566);
nor U12495 (N_12495,N_6664,N_9525);
nand U12496 (N_12496,N_9407,N_6674);
or U12497 (N_12497,N_7724,N_5237);
and U12498 (N_12498,N_7824,N_6029);
nor U12499 (N_12499,N_5589,N_9283);
nor U12500 (N_12500,N_5119,N_8455);
and U12501 (N_12501,N_8378,N_8077);
nand U12502 (N_12502,N_6803,N_9003);
or U12503 (N_12503,N_5088,N_7135);
and U12504 (N_12504,N_7826,N_8309);
or U12505 (N_12505,N_6152,N_6793);
or U12506 (N_12506,N_8518,N_7506);
and U12507 (N_12507,N_6833,N_6975);
and U12508 (N_12508,N_6116,N_7662);
and U12509 (N_12509,N_6821,N_6773);
and U12510 (N_12510,N_6040,N_7702);
nor U12511 (N_12511,N_6037,N_6827);
or U12512 (N_12512,N_9028,N_8473);
or U12513 (N_12513,N_5223,N_5159);
nand U12514 (N_12514,N_7376,N_7543);
nor U12515 (N_12515,N_6894,N_9509);
and U12516 (N_12516,N_5638,N_9821);
or U12517 (N_12517,N_9795,N_9748);
nor U12518 (N_12518,N_7078,N_5865);
nor U12519 (N_12519,N_5893,N_7717);
nand U12520 (N_12520,N_9227,N_8115);
and U12521 (N_12521,N_6635,N_5543);
or U12522 (N_12522,N_5663,N_9557);
and U12523 (N_12523,N_7756,N_9812);
nor U12524 (N_12524,N_6688,N_8988);
nor U12525 (N_12525,N_8146,N_6224);
and U12526 (N_12526,N_8623,N_7768);
nand U12527 (N_12527,N_6932,N_7417);
xnor U12528 (N_12528,N_6083,N_9007);
or U12529 (N_12529,N_9108,N_5188);
nor U12530 (N_12530,N_9418,N_8408);
or U12531 (N_12531,N_5576,N_9009);
or U12532 (N_12532,N_6088,N_5959);
nand U12533 (N_12533,N_9785,N_8305);
nand U12534 (N_12534,N_9504,N_5443);
nand U12535 (N_12535,N_5645,N_5002);
and U12536 (N_12536,N_7658,N_5589);
nor U12537 (N_12537,N_7456,N_7987);
nor U12538 (N_12538,N_7312,N_6322);
or U12539 (N_12539,N_5615,N_6103);
or U12540 (N_12540,N_5711,N_7157);
or U12541 (N_12541,N_6814,N_9413);
nand U12542 (N_12542,N_9382,N_6737);
xor U12543 (N_12543,N_6640,N_8823);
or U12544 (N_12544,N_8505,N_6698);
and U12545 (N_12545,N_9053,N_5520);
nand U12546 (N_12546,N_7264,N_8566);
or U12547 (N_12547,N_5706,N_8357);
or U12548 (N_12548,N_8977,N_5371);
and U12549 (N_12549,N_8032,N_7293);
or U12550 (N_12550,N_5708,N_8778);
and U12551 (N_12551,N_9603,N_6928);
xnor U12552 (N_12552,N_5474,N_5915);
and U12553 (N_12553,N_5098,N_7655);
and U12554 (N_12554,N_5961,N_7789);
or U12555 (N_12555,N_6069,N_7506);
and U12556 (N_12556,N_8506,N_5276);
and U12557 (N_12557,N_5922,N_6553);
nor U12558 (N_12558,N_9021,N_9154);
nand U12559 (N_12559,N_7242,N_7524);
and U12560 (N_12560,N_5301,N_5456);
or U12561 (N_12561,N_6037,N_8580);
or U12562 (N_12562,N_7330,N_9447);
and U12563 (N_12563,N_5650,N_5433);
or U12564 (N_12564,N_7927,N_6013);
nand U12565 (N_12565,N_6980,N_5042);
or U12566 (N_12566,N_8428,N_9984);
and U12567 (N_12567,N_5818,N_9272);
or U12568 (N_12568,N_5458,N_6930);
nor U12569 (N_12569,N_7186,N_9452);
nand U12570 (N_12570,N_7171,N_5731);
nand U12571 (N_12571,N_7995,N_6492);
and U12572 (N_12572,N_6514,N_8251);
nand U12573 (N_12573,N_6810,N_6525);
nor U12574 (N_12574,N_7789,N_8956);
and U12575 (N_12575,N_5580,N_8951);
or U12576 (N_12576,N_5427,N_5114);
and U12577 (N_12577,N_9505,N_7160);
and U12578 (N_12578,N_7695,N_6238);
or U12579 (N_12579,N_9913,N_8461);
and U12580 (N_12580,N_5157,N_8392);
or U12581 (N_12581,N_5702,N_7442);
nand U12582 (N_12582,N_7708,N_7638);
nand U12583 (N_12583,N_9023,N_8068);
nand U12584 (N_12584,N_5595,N_9015);
or U12585 (N_12585,N_7635,N_8885);
nand U12586 (N_12586,N_9139,N_7039);
or U12587 (N_12587,N_6981,N_6681);
nand U12588 (N_12588,N_9403,N_5622);
nand U12589 (N_12589,N_7406,N_5231);
or U12590 (N_12590,N_8988,N_5404);
nand U12591 (N_12591,N_7223,N_8458);
nor U12592 (N_12592,N_9467,N_9767);
or U12593 (N_12593,N_6064,N_9303);
nor U12594 (N_12594,N_9244,N_9757);
nand U12595 (N_12595,N_5285,N_8087);
nor U12596 (N_12596,N_9753,N_9685);
and U12597 (N_12597,N_9719,N_5715);
and U12598 (N_12598,N_9243,N_6470);
nand U12599 (N_12599,N_7627,N_9309);
and U12600 (N_12600,N_9421,N_8766);
or U12601 (N_12601,N_5764,N_8781);
nand U12602 (N_12602,N_5175,N_8973);
and U12603 (N_12603,N_6284,N_7895);
nand U12604 (N_12604,N_7485,N_8249);
nand U12605 (N_12605,N_8587,N_5863);
nor U12606 (N_12606,N_6447,N_7500);
and U12607 (N_12607,N_7715,N_8043);
nand U12608 (N_12608,N_6868,N_6744);
or U12609 (N_12609,N_8661,N_7839);
nand U12610 (N_12610,N_8088,N_6063);
and U12611 (N_12611,N_9783,N_9185);
nor U12612 (N_12612,N_8897,N_5224);
nor U12613 (N_12613,N_6858,N_8581);
xnor U12614 (N_12614,N_8641,N_7298);
nand U12615 (N_12615,N_5490,N_8566);
nor U12616 (N_12616,N_7483,N_6133);
or U12617 (N_12617,N_7893,N_8438);
or U12618 (N_12618,N_9200,N_7595);
nand U12619 (N_12619,N_6348,N_5122);
nor U12620 (N_12620,N_6762,N_5879);
nor U12621 (N_12621,N_5652,N_9855);
nand U12622 (N_12622,N_9191,N_8822);
nor U12623 (N_12623,N_7356,N_8946);
or U12624 (N_12624,N_5022,N_9707);
and U12625 (N_12625,N_6821,N_7239);
and U12626 (N_12626,N_8212,N_5828);
nor U12627 (N_12627,N_9273,N_6658);
nor U12628 (N_12628,N_7730,N_5368);
and U12629 (N_12629,N_5764,N_9846);
or U12630 (N_12630,N_8396,N_8351);
xor U12631 (N_12631,N_5384,N_8578);
or U12632 (N_12632,N_7330,N_7368);
and U12633 (N_12633,N_6505,N_8459);
or U12634 (N_12634,N_5185,N_5745);
nor U12635 (N_12635,N_6675,N_6432);
or U12636 (N_12636,N_7627,N_8427);
and U12637 (N_12637,N_7630,N_8715);
and U12638 (N_12638,N_6202,N_6567);
nand U12639 (N_12639,N_7476,N_9834);
nand U12640 (N_12640,N_9820,N_9925);
and U12641 (N_12641,N_5412,N_5536);
and U12642 (N_12642,N_6683,N_9579);
nor U12643 (N_12643,N_9815,N_6576);
nand U12644 (N_12644,N_7784,N_9402);
and U12645 (N_12645,N_6840,N_8957);
or U12646 (N_12646,N_9902,N_6901);
nor U12647 (N_12647,N_6412,N_5519);
and U12648 (N_12648,N_8247,N_8129);
or U12649 (N_12649,N_9759,N_5783);
and U12650 (N_12650,N_7581,N_5057);
and U12651 (N_12651,N_5960,N_8783);
nor U12652 (N_12652,N_5139,N_9966);
xor U12653 (N_12653,N_8135,N_9690);
nand U12654 (N_12654,N_7901,N_7107);
nor U12655 (N_12655,N_5641,N_6419);
and U12656 (N_12656,N_6999,N_5539);
and U12657 (N_12657,N_6969,N_9127);
nor U12658 (N_12658,N_9443,N_5990);
and U12659 (N_12659,N_5372,N_9510);
nor U12660 (N_12660,N_7830,N_5976);
nand U12661 (N_12661,N_5842,N_6715);
xor U12662 (N_12662,N_6339,N_5986);
or U12663 (N_12663,N_6158,N_8596);
and U12664 (N_12664,N_8186,N_7397);
and U12665 (N_12665,N_9951,N_6509);
nor U12666 (N_12666,N_5093,N_9316);
nand U12667 (N_12667,N_6243,N_8372);
nand U12668 (N_12668,N_7712,N_8873);
nand U12669 (N_12669,N_9501,N_5404);
or U12670 (N_12670,N_8193,N_9913);
and U12671 (N_12671,N_7280,N_9670);
nand U12672 (N_12672,N_7046,N_7967);
nor U12673 (N_12673,N_9229,N_7821);
nor U12674 (N_12674,N_9228,N_6698);
or U12675 (N_12675,N_5909,N_6881);
or U12676 (N_12676,N_6666,N_7722);
or U12677 (N_12677,N_6927,N_9596);
nand U12678 (N_12678,N_9332,N_8205);
or U12679 (N_12679,N_5894,N_7054);
and U12680 (N_12680,N_8173,N_7043);
nand U12681 (N_12681,N_5491,N_6156);
or U12682 (N_12682,N_5470,N_6869);
and U12683 (N_12683,N_5170,N_9225);
or U12684 (N_12684,N_8845,N_9862);
or U12685 (N_12685,N_9388,N_8834);
or U12686 (N_12686,N_6118,N_9421);
nor U12687 (N_12687,N_5718,N_6687);
nor U12688 (N_12688,N_6430,N_7080);
and U12689 (N_12689,N_9139,N_7610);
nand U12690 (N_12690,N_7004,N_6524);
nand U12691 (N_12691,N_9950,N_6986);
or U12692 (N_12692,N_5721,N_5177);
nand U12693 (N_12693,N_6912,N_9658);
nor U12694 (N_12694,N_5750,N_7033);
nand U12695 (N_12695,N_8964,N_6074);
nand U12696 (N_12696,N_9937,N_5322);
and U12697 (N_12697,N_9340,N_9481);
or U12698 (N_12698,N_5516,N_5193);
nand U12699 (N_12699,N_7906,N_9017);
nand U12700 (N_12700,N_7953,N_5548);
nand U12701 (N_12701,N_7748,N_9067);
nor U12702 (N_12702,N_5463,N_8219);
nor U12703 (N_12703,N_7555,N_8697);
nand U12704 (N_12704,N_5069,N_5697);
nor U12705 (N_12705,N_6621,N_6182);
nand U12706 (N_12706,N_8973,N_9093);
or U12707 (N_12707,N_6492,N_8288);
and U12708 (N_12708,N_7084,N_8227);
nand U12709 (N_12709,N_9051,N_9130);
nand U12710 (N_12710,N_6377,N_8925);
xor U12711 (N_12711,N_7449,N_9139);
or U12712 (N_12712,N_6978,N_5329);
or U12713 (N_12713,N_7204,N_8820);
or U12714 (N_12714,N_8124,N_9681);
nor U12715 (N_12715,N_7193,N_9763);
or U12716 (N_12716,N_7602,N_5002);
nor U12717 (N_12717,N_8505,N_7720);
or U12718 (N_12718,N_5608,N_5043);
xnor U12719 (N_12719,N_8925,N_7583);
and U12720 (N_12720,N_6219,N_6908);
nor U12721 (N_12721,N_5802,N_9196);
nand U12722 (N_12722,N_8866,N_8686);
and U12723 (N_12723,N_6896,N_8729);
nand U12724 (N_12724,N_9064,N_6266);
and U12725 (N_12725,N_6793,N_6689);
nor U12726 (N_12726,N_6172,N_9157);
nor U12727 (N_12727,N_5094,N_9955);
and U12728 (N_12728,N_9792,N_7839);
nor U12729 (N_12729,N_7638,N_5319);
nor U12730 (N_12730,N_8186,N_9206);
or U12731 (N_12731,N_8232,N_9584);
and U12732 (N_12732,N_6762,N_5507);
nor U12733 (N_12733,N_8317,N_5194);
nand U12734 (N_12734,N_7277,N_7115);
or U12735 (N_12735,N_5792,N_7561);
xnor U12736 (N_12736,N_6357,N_7524);
xnor U12737 (N_12737,N_7393,N_7238);
or U12738 (N_12738,N_8590,N_9044);
nor U12739 (N_12739,N_9282,N_6718);
or U12740 (N_12740,N_8990,N_8293);
nand U12741 (N_12741,N_8617,N_5644);
and U12742 (N_12742,N_8325,N_6585);
or U12743 (N_12743,N_7776,N_6182);
nand U12744 (N_12744,N_5043,N_8340);
nand U12745 (N_12745,N_5677,N_8072);
nor U12746 (N_12746,N_7762,N_7051);
nor U12747 (N_12747,N_7951,N_7943);
nand U12748 (N_12748,N_5050,N_5017);
or U12749 (N_12749,N_7732,N_9871);
or U12750 (N_12750,N_7463,N_5904);
and U12751 (N_12751,N_7146,N_7417);
and U12752 (N_12752,N_9677,N_7097);
and U12753 (N_12753,N_5700,N_5340);
or U12754 (N_12754,N_5784,N_9567);
nor U12755 (N_12755,N_7593,N_8390);
and U12756 (N_12756,N_5626,N_7597);
or U12757 (N_12757,N_8131,N_7670);
nand U12758 (N_12758,N_9004,N_6719);
and U12759 (N_12759,N_9817,N_7008);
nor U12760 (N_12760,N_8073,N_5540);
or U12761 (N_12761,N_6148,N_6244);
nor U12762 (N_12762,N_8027,N_9603);
nand U12763 (N_12763,N_9548,N_9996);
and U12764 (N_12764,N_8043,N_7354);
and U12765 (N_12765,N_8397,N_7637);
nand U12766 (N_12766,N_7115,N_5115);
nand U12767 (N_12767,N_8756,N_6559);
or U12768 (N_12768,N_8567,N_7503);
nor U12769 (N_12769,N_5393,N_5696);
nor U12770 (N_12770,N_9890,N_6356);
and U12771 (N_12771,N_9036,N_6668);
nand U12772 (N_12772,N_9090,N_8840);
nand U12773 (N_12773,N_7985,N_8953);
or U12774 (N_12774,N_5357,N_7667);
nand U12775 (N_12775,N_7567,N_6458);
or U12776 (N_12776,N_7517,N_7241);
and U12777 (N_12777,N_8467,N_7094);
or U12778 (N_12778,N_7276,N_8117);
or U12779 (N_12779,N_7640,N_6831);
xnor U12780 (N_12780,N_5839,N_6834);
xor U12781 (N_12781,N_8689,N_9716);
or U12782 (N_12782,N_6889,N_7964);
or U12783 (N_12783,N_8261,N_7917);
nor U12784 (N_12784,N_5442,N_5274);
or U12785 (N_12785,N_6649,N_5977);
and U12786 (N_12786,N_7081,N_6034);
or U12787 (N_12787,N_6267,N_5833);
or U12788 (N_12788,N_8280,N_5716);
nand U12789 (N_12789,N_7996,N_7100);
nor U12790 (N_12790,N_6288,N_7692);
nor U12791 (N_12791,N_8472,N_7946);
nor U12792 (N_12792,N_5624,N_8667);
nor U12793 (N_12793,N_5246,N_7128);
and U12794 (N_12794,N_5688,N_6018);
nor U12795 (N_12795,N_9020,N_9483);
nand U12796 (N_12796,N_7522,N_6509);
nand U12797 (N_12797,N_8914,N_8018);
and U12798 (N_12798,N_5902,N_5945);
nand U12799 (N_12799,N_5678,N_7590);
and U12800 (N_12800,N_9133,N_6887);
nor U12801 (N_12801,N_6669,N_7451);
or U12802 (N_12802,N_7612,N_5925);
and U12803 (N_12803,N_7956,N_6089);
or U12804 (N_12804,N_7566,N_6574);
nor U12805 (N_12805,N_7200,N_9694);
nor U12806 (N_12806,N_5306,N_5502);
or U12807 (N_12807,N_8065,N_7302);
or U12808 (N_12808,N_7928,N_6006);
or U12809 (N_12809,N_6344,N_6382);
or U12810 (N_12810,N_9638,N_9027);
nor U12811 (N_12811,N_5865,N_7826);
nor U12812 (N_12812,N_5336,N_8728);
and U12813 (N_12813,N_6444,N_8633);
nor U12814 (N_12814,N_9528,N_7396);
or U12815 (N_12815,N_6064,N_7495);
nand U12816 (N_12816,N_6503,N_6115);
and U12817 (N_12817,N_7495,N_9712);
or U12818 (N_12818,N_6500,N_8835);
and U12819 (N_12819,N_9608,N_9524);
nor U12820 (N_12820,N_6879,N_5346);
nand U12821 (N_12821,N_6855,N_5530);
or U12822 (N_12822,N_5525,N_5792);
xnor U12823 (N_12823,N_7405,N_6065);
nand U12824 (N_12824,N_8029,N_8632);
and U12825 (N_12825,N_5440,N_5771);
nand U12826 (N_12826,N_9507,N_9236);
or U12827 (N_12827,N_9247,N_9592);
nor U12828 (N_12828,N_8048,N_5108);
nand U12829 (N_12829,N_7129,N_6045);
nor U12830 (N_12830,N_8173,N_7205);
or U12831 (N_12831,N_8955,N_7958);
nand U12832 (N_12832,N_9311,N_9437);
and U12833 (N_12833,N_6428,N_8325);
nor U12834 (N_12834,N_5940,N_7124);
nand U12835 (N_12835,N_7092,N_8917);
nor U12836 (N_12836,N_9527,N_5005);
or U12837 (N_12837,N_6903,N_9950);
and U12838 (N_12838,N_5496,N_8018);
or U12839 (N_12839,N_8845,N_7578);
nand U12840 (N_12840,N_5536,N_9509);
and U12841 (N_12841,N_7861,N_6088);
nor U12842 (N_12842,N_9127,N_6116);
and U12843 (N_12843,N_8301,N_8466);
nand U12844 (N_12844,N_7095,N_9147);
and U12845 (N_12845,N_8745,N_8387);
nand U12846 (N_12846,N_5495,N_8759);
nor U12847 (N_12847,N_8165,N_9592);
nand U12848 (N_12848,N_9462,N_5408);
or U12849 (N_12849,N_9279,N_8326);
nand U12850 (N_12850,N_8838,N_6569);
or U12851 (N_12851,N_9594,N_7817);
and U12852 (N_12852,N_9677,N_7535);
nor U12853 (N_12853,N_9078,N_6685);
nand U12854 (N_12854,N_7407,N_5710);
nor U12855 (N_12855,N_7768,N_6839);
nand U12856 (N_12856,N_9213,N_5925);
or U12857 (N_12857,N_8847,N_9716);
or U12858 (N_12858,N_8843,N_5732);
nand U12859 (N_12859,N_9183,N_9577);
or U12860 (N_12860,N_9455,N_7523);
nand U12861 (N_12861,N_7563,N_6842);
nor U12862 (N_12862,N_6110,N_6761);
nand U12863 (N_12863,N_6151,N_9541);
or U12864 (N_12864,N_6277,N_5904);
nand U12865 (N_12865,N_5559,N_9871);
nor U12866 (N_12866,N_6051,N_8619);
or U12867 (N_12867,N_7397,N_9478);
and U12868 (N_12868,N_8396,N_9486);
and U12869 (N_12869,N_7860,N_9272);
and U12870 (N_12870,N_8640,N_9265);
nor U12871 (N_12871,N_7574,N_6943);
and U12872 (N_12872,N_5804,N_9260);
and U12873 (N_12873,N_6049,N_7121);
nand U12874 (N_12874,N_9836,N_5381);
nand U12875 (N_12875,N_7537,N_5921);
nor U12876 (N_12876,N_8643,N_8054);
nand U12877 (N_12877,N_5606,N_9169);
nand U12878 (N_12878,N_5345,N_9990);
and U12879 (N_12879,N_7149,N_8663);
xor U12880 (N_12880,N_9969,N_6714);
nor U12881 (N_12881,N_5350,N_8096);
nand U12882 (N_12882,N_5825,N_5457);
or U12883 (N_12883,N_5422,N_9820);
xor U12884 (N_12884,N_6031,N_5326);
and U12885 (N_12885,N_9138,N_9127);
and U12886 (N_12886,N_7806,N_7832);
nand U12887 (N_12887,N_8197,N_8850);
or U12888 (N_12888,N_9439,N_9933);
and U12889 (N_12889,N_9938,N_8784);
nor U12890 (N_12890,N_6107,N_5338);
nor U12891 (N_12891,N_5222,N_9472);
nor U12892 (N_12892,N_9316,N_7292);
or U12893 (N_12893,N_7990,N_8390);
or U12894 (N_12894,N_6723,N_7245);
or U12895 (N_12895,N_9208,N_6495);
nand U12896 (N_12896,N_5785,N_5535);
nor U12897 (N_12897,N_8994,N_6512);
or U12898 (N_12898,N_9685,N_9374);
and U12899 (N_12899,N_5828,N_5889);
nor U12900 (N_12900,N_9058,N_6252);
and U12901 (N_12901,N_5063,N_9554);
nand U12902 (N_12902,N_7490,N_8152);
nor U12903 (N_12903,N_8113,N_5541);
and U12904 (N_12904,N_6996,N_9505);
nor U12905 (N_12905,N_7298,N_8285);
nand U12906 (N_12906,N_5619,N_5528);
and U12907 (N_12907,N_6638,N_6736);
nor U12908 (N_12908,N_7226,N_8308);
and U12909 (N_12909,N_9315,N_7011);
nor U12910 (N_12910,N_9324,N_6094);
or U12911 (N_12911,N_5488,N_7936);
or U12912 (N_12912,N_8838,N_5505);
or U12913 (N_12913,N_5882,N_7473);
and U12914 (N_12914,N_9052,N_6203);
xnor U12915 (N_12915,N_9741,N_6118);
nand U12916 (N_12916,N_5528,N_5423);
nor U12917 (N_12917,N_8458,N_8442);
or U12918 (N_12918,N_7869,N_5098);
or U12919 (N_12919,N_7036,N_6664);
nand U12920 (N_12920,N_5036,N_5658);
or U12921 (N_12921,N_8462,N_8449);
nand U12922 (N_12922,N_5567,N_5342);
or U12923 (N_12923,N_5912,N_5960);
nor U12924 (N_12924,N_8872,N_7249);
nor U12925 (N_12925,N_5633,N_5101);
and U12926 (N_12926,N_5674,N_5170);
nand U12927 (N_12927,N_8462,N_8784);
or U12928 (N_12928,N_5561,N_7587);
nand U12929 (N_12929,N_6186,N_8560);
nor U12930 (N_12930,N_9293,N_5717);
or U12931 (N_12931,N_7588,N_6748);
nand U12932 (N_12932,N_9213,N_9625);
nand U12933 (N_12933,N_5498,N_6008);
nand U12934 (N_12934,N_7055,N_9884);
and U12935 (N_12935,N_6477,N_7680);
and U12936 (N_12936,N_8159,N_5370);
nand U12937 (N_12937,N_6677,N_8512);
nor U12938 (N_12938,N_6315,N_5895);
nand U12939 (N_12939,N_5818,N_8413);
and U12940 (N_12940,N_8534,N_6278);
nor U12941 (N_12941,N_8024,N_8282);
nor U12942 (N_12942,N_9617,N_5695);
or U12943 (N_12943,N_7768,N_7883);
or U12944 (N_12944,N_9944,N_7272);
and U12945 (N_12945,N_6437,N_9152);
nand U12946 (N_12946,N_6518,N_5536);
and U12947 (N_12947,N_7360,N_7954);
and U12948 (N_12948,N_7463,N_9114);
or U12949 (N_12949,N_6432,N_7180);
nand U12950 (N_12950,N_7768,N_7674);
or U12951 (N_12951,N_9603,N_5068);
nand U12952 (N_12952,N_5039,N_6537);
nand U12953 (N_12953,N_7348,N_8055);
or U12954 (N_12954,N_7410,N_9670);
and U12955 (N_12955,N_7269,N_6109);
nand U12956 (N_12956,N_7277,N_7178);
nand U12957 (N_12957,N_8374,N_5003);
nor U12958 (N_12958,N_6672,N_9644);
or U12959 (N_12959,N_5512,N_7981);
or U12960 (N_12960,N_7927,N_6843);
nor U12961 (N_12961,N_5822,N_5683);
and U12962 (N_12962,N_5139,N_6849);
nor U12963 (N_12963,N_8199,N_6328);
and U12964 (N_12964,N_5297,N_5569);
and U12965 (N_12965,N_7981,N_6023);
nand U12966 (N_12966,N_6420,N_7681);
and U12967 (N_12967,N_5718,N_8879);
or U12968 (N_12968,N_8922,N_8196);
nand U12969 (N_12969,N_9024,N_7785);
nand U12970 (N_12970,N_6178,N_6502);
and U12971 (N_12971,N_8524,N_9686);
and U12972 (N_12972,N_6906,N_5127);
or U12973 (N_12973,N_6560,N_9194);
nand U12974 (N_12974,N_6071,N_8658);
nor U12975 (N_12975,N_9813,N_8514);
nand U12976 (N_12976,N_6130,N_5623);
and U12977 (N_12977,N_8406,N_8966);
and U12978 (N_12978,N_6096,N_9352);
xnor U12979 (N_12979,N_6530,N_5988);
and U12980 (N_12980,N_6357,N_8398);
or U12981 (N_12981,N_9158,N_5812);
and U12982 (N_12982,N_7305,N_9981);
or U12983 (N_12983,N_5671,N_5555);
and U12984 (N_12984,N_5492,N_9502);
nor U12985 (N_12985,N_5107,N_6397);
and U12986 (N_12986,N_7853,N_8918);
and U12987 (N_12987,N_8850,N_5654);
nand U12988 (N_12988,N_9842,N_9859);
nand U12989 (N_12989,N_7343,N_9093);
xnor U12990 (N_12990,N_8324,N_5853);
nand U12991 (N_12991,N_9520,N_8184);
and U12992 (N_12992,N_9182,N_5504);
and U12993 (N_12993,N_6930,N_7666);
nor U12994 (N_12994,N_5158,N_6361);
nand U12995 (N_12995,N_8391,N_6949);
or U12996 (N_12996,N_9093,N_6390);
nand U12997 (N_12997,N_7331,N_8939);
or U12998 (N_12998,N_8417,N_8826);
or U12999 (N_12999,N_9780,N_7963);
nand U13000 (N_13000,N_8039,N_9869);
or U13001 (N_13001,N_6089,N_5551);
or U13002 (N_13002,N_5621,N_7092);
or U13003 (N_13003,N_5058,N_5202);
and U13004 (N_13004,N_5695,N_8937);
or U13005 (N_13005,N_7197,N_5607);
nor U13006 (N_13006,N_8103,N_6623);
nor U13007 (N_13007,N_7784,N_9534);
nor U13008 (N_13008,N_9137,N_7087);
nor U13009 (N_13009,N_6285,N_5185);
and U13010 (N_13010,N_5510,N_7928);
and U13011 (N_13011,N_6924,N_5803);
and U13012 (N_13012,N_5875,N_6718);
nand U13013 (N_13013,N_9105,N_9844);
or U13014 (N_13014,N_8747,N_5724);
nor U13015 (N_13015,N_8400,N_7446);
or U13016 (N_13016,N_6932,N_8679);
nand U13017 (N_13017,N_5793,N_8042);
and U13018 (N_13018,N_9336,N_6041);
and U13019 (N_13019,N_8422,N_5854);
and U13020 (N_13020,N_5825,N_5592);
or U13021 (N_13021,N_8406,N_7320);
or U13022 (N_13022,N_9922,N_9009);
or U13023 (N_13023,N_7177,N_5096);
or U13024 (N_13024,N_7289,N_7610);
nor U13025 (N_13025,N_6794,N_8450);
nor U13026 (N_13026,N_7348,N_7561);
and U13027 (N_13027,N_8269,N_8622);
nor U13028 (N_13028,N_7407,N_8483);
and U13029 (N_13029,N_9775,N_9852);
nor U13030 (N_13030,N_5553,N_6090);
nor U13031 (N_13031,N_5357,N_6062);
nand U13032 (N_13032,N_8549,N_6377);
nor U13033 (N_13033,N_7934,N_8356);
xor U13034 (N_13034,N_8701,N_5583);
or U13035 (N_13035,N_9282,N_9750);
nor U13036 (N_13036,N_9106,N_5260);
nand U13037 (N_13037,N_7608,N_8241);
or U13038 (N_13038,N_9885,N_9958);
or U13039 (N_13039,N_8474,N_7022);
and U13040 (N_13040,N_8196,N_8908);
nand U13041 (N_13041,N_5746,N_9880);
or U13042 (N_13042,N_9753,N_5688);
nor U13043 (N_13043,N_6657,N_5396);
nand U13044 (N_13044,N_6928,N_8280);
and U13045 (N_13045,N_8214,N_6700);
nor U13046 (N_13046,N_6665,N_6227);
and U13047 (N_13047,N_5236,N_6242);
nor U13048 (N_13048,N_7588,N_5723);
and U13049 (N_13049,N_7381,N_8365);
nand U13050 (N_13050,N_6771,N_8748);
nor U13051 (N_13051,N_8594,N_9044);
nor U13052 (N_13052,N_5213,N_8729);
nor U13053 (N_13053,N_5360,N_6498);
and U13054 (N_13054,N_7614,N_7972);
and U13055 (N_13055,N_6465,N_6368);
and U13056 (N_13056,N_5144,N_9586);
nand U13057 (N_13057,N_8312,N_9218);
nand U13058 (N_13058,N_9465,N_7742);
nor U13059 (N_13059,N_5596,N_6126);
or U13060 (N_13060,N_5965,N_8228);
or U13061 (N_13061,N_5279,N_9113);
nor U13062 (N_13062,N_9849,N_5394);
nor U13063 (N_13063,N_8981,N_9449);
nor U13064 (N_13064,N_5125,N_6919);
or U13065 (N_13065,N_6955,N_6809);
nor U13066 (N_13066,N_8670,N_9643);
nor U13067 (N_13067,N_6169,N_5958);
or U13068 (N_13068,N_5074,N_6840);
and U13069 (N_13069,N_9036,N_8038);
nor U13070 (N_13070,N_9341,N_8908);
or U13071 (N_13071,N_8692,N_8842);
or U13072 (N_13072,N_9757,N_5989);
nand U13073 (N_13073,N_5844,N_6985);
xnor U13074 (N_13074,N_6355,N_9009);
or U13075 (N_13075,N_7712,N_5671);
nor U13076 (N_13076,N_9522,N_7713);
and U13077 (N_13077,N_6196,N_6516);
nand U13078 (N_13078,N_8502,N_6822);
or U13079 (N_13079,N_5765,N_6116);
nand U13080 (N_13080,N_8052,N_6584);
and U13081 (N_13081,N_9178,N_8588);
or U13082 (N_13082,N_5267,N_7434);
and U13083 (N_13083,N_7959,N_9837);
nor U13084 (N_13084,N_6961,N_9698);
nand U13085 (N_13085,N_8237,N_5818);
nand U13086 (N_13086,N_5067,N_9722);
nand U13087 (N_13087,N_7569,N_6835);
and U13088 (N_13088,N_5929,N_5315);
or U13089 (N_13089,N_8630,N_9754);
or U13090 (N_13090,N_6891,N_7774);
and U13091 (N_13091,N_8179,N_6995);
nand U13092 (N_13092,N_8063,N_9482);
nor U13093 (N_13093,N_7190,N_8984);
nor U13094 (N_13094,N_8923,N_6083);
or U13095 (N_13095,N_8285,N_7588);
nor U13096 (N_13096,N_5680,N_6052);
nand U13097 (N_13097,N_8766,N_5097);
and U13098 (N_13098,N_7039,N_5305);
or U13099 (N_13099,N_8459,N_9928);
nand U13100 (N_13100,N_9128,N_6316);
and U13101 (N_13101,N_9964,N_5642);
and U13102 (N_13102,N_8451,N_6800);
xnor U13103 (N_13103,N_5217,N_6562);
nand U13104 (N_13104,N_6906,N_5056);
nand U13105 (N_13105,N_9947,N_6460);
nand U13106 (N_13106,N_8413,N_9162);
nand U13107 (N_13107,N_9063,N_8942);
or U13108 (N_13108,N_9883,N_6174);
nor U13109 (N_13109,N_7110,N_8889);
nand U13110 (N_13110,N_8915,N_9174);
nand U13111 (N_13111,N_5285,N_7197);
nand U13112 (N_13112,N_9549,N_5611);
nand U13113 (N_13113,N_7210,N_8721);
and U13114 (N_13114,N_6415,N_5544);
nor U13115 (N_13115,N_9635,N_8324);
or U13116 (N_13116,N_9651,N_6277);
and U13117 (N_13117,N_6720,N_8874);
and U13118 (N_13118,N_9724,N_9532);
nor U13119 (N_13119,N_6014,N_7425);
and U13120 (N_13120,N_6337,N_9961);
nor U13121 (N_13121,N_7735,N_7880);
nand U13122 (N_13122,N_6465,N_9665);
nor U13123 (N_13123,N_9468,N_7872);
xnor U13124 (N_13124,N_6330,N_6596);
or U13125 (N_13125,N_7076,N_5362);
nand U13126 (N_13126,N_9318,N_6495);
or U13127 (N_13127,N_8901,N_5697);
nor U13128 (N_13128,N_5587,N_9326);
nand U13129 (N_13129,N_9400,N_9098);
nor U13130 (N_13130,N_8507,N_8083);
nand U13131 (N_13131,N_8524,N_8455);
and U13132 (N_13132,N_9390,N_7684);
or U13133 (N_13133,N_5786,N_6268);
nor U13134 (N_13134,N_6567,N_9839);
nor U13135 (N_13135,N_7864,N_9572);
nor U13136 (N_13136,N_9527,N_7021);
and U13137 (N_13137,N_8990,N_5330);
nor U13138 (N_13138,N_8267,N_6395);
or U13139 (N_13139,N_6594,N_6041);
nand U13140 (N_13140,N_6467,N_8880);
and U13141 (N_13141,N_9929,N_6910);
and U13142 (N_13142,N_6454,N_8062);
and U13143 (N_13143,N_7654,N_7840);
nand U13144 (N_13144,N_6229,N_5285);
nor U13145 (N_13145,N_5529,N_7797);
and U13146 (N_13146,N_7042,N_7530);
or U13147 (N_13147,N_9269,N_7609);
nand U13148 (N_13148,N_8527,N_7925);
or U13149 (N_13149,N_5720,N_8360);
nor U13150 (N_13150,N_7372,N_5989);
or U13151 (N_13151,N_6223,N_9645);
and U13152 (N_13152,N_6383,N_6746);
xor U13153 (N_13153,N_7520,N_7637);
or U13154 (N_13154,N_6765,N_6982);
nand U13155 (N_13155,N_9437,N_5866);
nand U13156 (N_13156,N_7046,N_8652);
or U13157 (N_13157,N_6956,N_5833);
nand U13158 (N_13158,N_7461,N_6534);
or U13159 (N_13159,N_6413,N_5067);
or U13160 (N_13160,N_6156,N_6607);
xor U13161 (N_13161,N_8646,N_8482);
and U13162 (N_13162,N_9343,N_9377);
or U13163 (N_13163,N_7539,N_6231);
nand U13164 (N_13164,N_9210,N_5329);
and U13165 (N_13165,N_9242,N_9824);
xor U13166 (N_13166,N_7383,N_5203);
nand U13167 (N_13167,N_9984,N_7085);
or U13168 (N_13168,N_6160,N_5128);
nand U13169 (N_13169,N_6606,N_5650);
and U13170 (N_13170,N_7921,N_9500);
and U13171 (N_13171,N_5577,N_5020);
or U13172 (N_13172,N_8237,N_6228);
nand U13173 (N_13173,N_8020,N_6407);
or U13174 (N_13174,N_7429,N_9439);
nor U13175 (N_13175,N_9711,N_5440);
or U13176 (N_13176,N_5192,N_5366);
or U13177 (N_13177,N_7047,N_7045);
and U13178 (N_13178,N_6046,N_7958);
nor U13179 (N_13179,N_5096,N_9067);
and U13180 (N_13180,N_9483,N_6553);
or U13181 (N_13181,N_8123,N_7807);
nand U13182 (N_13182,N_8058,N_7941);
nor U13183 (N_13183,N_7289,N_7792);
and U13184 (N_13184,N_9561,N_5044);
nand U13185 (N_13185,N_5511,N_6774);
or U13186 (N_13186,N_6613,N_9429);
nand U13187 (N_13187,N_8224,N_6691);
nand U13188 (N_13188,N_6319,N_5349);
and U13189 (N_13189,N_7186,N_6379);
and U13190 (N_13190,N_8828,N_6839);
and U13191 (N_13191,N_6493,N_9449);
nor U13192 (N_13192,N_5038,N_6694);
or U13193 (N_13193,N_6724,N_8634);
nand U13194 (N_13194,N_6732,N_8526);
nand U13195 (N_13195,N_8287,N_8598);
nor U13196 (N_13196,N_5935,N_7445);
nand U13197 (N_13197,N_9512,N_9987);
or U13198 (N_13198,N_8635,N_5964);
nor U13199 (N_13199,N_5241,N_9363);
and U13200 (N_13200,N_8020,N_5909);
and U13201 (N_13201,N_5914,N_5680);
nor U13202 (N_13202,N_5497,N_7942);
or U13203 (N_13203,N_5097,N_7299);
or U13204 (N_13204,N_6690,N_5251);
nor U13205 (N_13205,N_5503,N_8799);
and U13206 (N_13206,N_8186,N_9436);
or U13207 (N_13207,N_6991,N_8627);
nor U13208 (N_13208,N_7829,N_9650);
or U13209 (N_13209,N_5762,N_5412);
or U13210 (N_13210,N_9382,N_6522);
and U13211 (N_13211,N_9535,N_7827);
nor U13212 (N_13212,N_6741,N_8319);
nand U13213 (N_13213,N_9964,N_5794);
and U13214 (N_13214,N_6564,N_6201);
nand U13215 (N_13215,N_5127,N_7906);
nor U13216 (N_13216,N_7210,N_6939);
or U13217 (N_13217,N_8101,N_6421);
and U13218 (N_13218,N_9091,N_7939);
nor U13219 (N_13219,N_8968,N_8836);
nor U13220 (N_13220,N_9327,N_6914);
or U13221 (N_13221,N_8015,N_7761);
or U13222 (N_13222,N_6517,N_8009);
nand U13223 (N_13223,N_7002,N_5405);
or U13224 (N_13224,N_6004,N_5023);
or U13225 (N_13225,N_7255,N_5828);
and U13226 (N_13226,N_9292,N_7986);
nor U13227 (N_13227,N_7844,N_9222);
nand U13228 (N_13228,N_8424,N_5188);
and U13229 (N_13229,N_8441,N_8573);
or U13230 (N_13230,N_5544,N_9762);
and U13231 (N_13231,N_8338,N_6502);
or U13232 (N_13232,N_7503,N_9584);
or U13233 (N_13233,N_9702,N_8740);
nor U13234 (N_13234,N_5506,N_5654);
nand U13235 (N_13235,N_5918,N_5409);
nor U13236 (N_13236,N_8006,N_9742);
and U13237 (N_13237,N_8086,N_7808);
nor U13238 (N_13238,N_8102,N_6797);
and U13239 (N_13239,N_9528,N_7126);
and U13240 (N_13240,N_7389,N_9743);
or U13241 (N_13241,N_9183,N_9112);
and U13242 (N_13242,N_6410,N_7234);
nand U13243 (N_13243,N_8798,N_7119);
nand U13244 (N_13244,N_7497,N_9892);
xnor U13245 (N_13245,N_6826,N_7692);
nand U13246 (N_13246,N_8465,N_7328);
nand U13247 (N_13247,N_7968,N_9560);
nor U13248 (N_13248,N_8400,N_9434);
nand U13249 (N_13249,N_6951,N_9332);
nor U13250 (N_13250,N_8568,N_9087);
nand U13251 (N_13251,N_9026,N_9439);
nand U13252 (N_13252,N_6961,N_9226);
or U13253 (N_13253,N_8407,N_7919);
and U13254 (N_13254,N_9672,N_5515);
nand U13255 (N_13255,N_7721,N_7139);
and U13256 (N_13256,N_5657,N_5738);
nor U13257 (N_13257,N_5967,N_5870);
nor U13258 (N_13258,N_7278,N_7431);
nand U13259 (N_13259,N_9313,N_7989);
and U13260 (N_13260,N_9155,N_8332);
or U13261 (N_13261,N_7669,N_6891);
nor U13262 (N_13262,N_5639,N_6361);
and U13263 (N_13263,N_8815,N_6202);
and U13264 (N_13264,N_6036,N_5645);
and U13265 (N_13265,N_9049,N_8883);
nor U13266 (N_13266,N_9720,N_5159);
and U13267 (N_13267,N_9379,N_8304);
nand U13268 (N_13268,N_7093,N_9880);
or U13269 (N_13269,N_9017,N_9466);
and U13270 (N_13270,N_5378,N_6555);
nor U13271 (N_13271,N_7377,N_8054);
and U13272 (N_13272,N_6601,N_5478);
and U13273 (N_13273,N_7384,N_5693);
or U13274 (N_13274,N_9981,N_9753);
or U13275 (N_13275,N_6292,N_9018);
or U13276 (N_13276,N_9066,N_7500);
nand U13277 (N_13277,N_6789,N_5360);
or U13278 (N_13278,N_5409,N_6285);
nor U13279 (N_13279,N_7043,N_8551);
or U13280 (N_13280,N_8818,N_6732);
and U13281 (N_13281,N_6281,N_6965);
nor U13282 (N_13282,N_9871,N_9853);
and U13283 (N_13283,N_7729,N_5700);
and U13284 (N_13284,N_8543,N_8399);
or U13285 (N_13285,N_9629,N_5498);
nand U13286 (N_13286,N_9509,N_7714);
and U13287 (N_13287,N_7772,N_8940);
and U13288 (N_13288,N_9957,N_7566);
nor U13289 (N_13289,N_7480,N_7727);
nand U13290 (N_13290,N_8417,N_5318);
and U13291 (N_13291,N_7413,N_7623);
nand U13292 (N_13292,N_7391,N_9235);
nand U13293 (N_13293,N_7071,N_6127);
and U13294 (N_13294,N_6404,N_8410);
and U13295 (N_13295,N_7496,N_8925);
nand U13296 (N_13296,N_5497,N_7939);
or U13297 (N_13297,N_6900,N_9722);
or U13298 (N_13298,N_7433,N_5726);
and U13299 (N_13299,N_8561,N_9389);
and U13300 (N_13300,N_8221,N_5243);
and U13301 (N_13301,N_7570,N_7857);
nand U13302 (N_13302,N_5941,N_9184);
nand U13303 (N_13303,N_9157,N_7342);
nor U13304 (N_13304,N_5899,N_9355);
nor U13305 (N_13305,N_9245,N_6906);
and U13306 (N_13306,N_7644,N_6752);
xor U13307 (N_13307,N_6271,N_8425);
nor U13308 (N_13308,N_7528,N_7053);
nand U13309 (N_13309,N_8280,N_6291);
and U13310 (N_13310,N_8161,N_7996);
nand U13311 (N_13311,N_8103,N_9856);
or U13312 (N_13312,N_6735,N_9974);
nor U13313 (N_13313,N_7198,N_5229);
and U13314 (N_13314,N_6854,N_5482);
nand U13315 (N_13315,N_9118,N_6123);
nand U13316 (N_13316,N_9264,N_6619);
nor U13317 (N_13317,N_5360,N_9104);
nand U13318 (N_13318,N_8389,N_5450);
nand U13319 (N_13319,N_6571,N_7990);
and U13320 (N_13320,N_9699,N_8231);
nand U13321 (N_13321,N_7170,N_8387);
xnor U13322 (N_13322,N_6301,N_9750);
nor U13323 (N_13323,N_7171,N_8028);
nor U13324 (N_13324,N_9441,N_8811);
or U13325 (N_13325,N_9267,N_9977);
nand U13326 (N_13326,N_7801,N_5858);
or U13327 (N_13327,N_6224,N_5798);
or U13328 (N_13328,N_7788,N_8171);
nand U13329 (N_13329,N_8404,N_5469);
or U13330 (N_13330,N_6014,N_7799);
and U13331 (N_13331,N_6875,N_5823);
xor U13332 (N_13332,N_6385,N_8421);
nor U13333 (N_13333,N_6787,N_9069);
nand U13334 (N_13334,N_7116,N_5422);
and U13335 (N_13335,N_7219,N_8590);
and U13336 (N_13336,N_9297,N_5342);
nand U13337 (N_13337,N_9620,N_8038);
and U13338 (N_13338,N_5004,N_5134);
or U13339 (N_13339,N_6209,N_8184);
nor U13340 (N_13340,N_6549,N_8936);
and U13341 (N_13341,N_5465,N_9451);
nor U13342 (N_13342,N_9611,N_5365);
nor U13343 (N_13343,N_6279,N_8287);
or U13344 (N_13344,N_8151,N_5761);
and U13345 (N_13345,N_8391,N_5277);
or U13346 (N_13346,N_6909,N_9248);
nand U13347 (N_13347,N_5929,N_9626);
and U13348 (N_13348,N_5359,N_9381);
or U13349 (N_13349,N_8424,N_9923);
or U13350 (N_13350,N_7850,N_6152);
nand U13351 (N_13351,N_5270,N_7285);
nand U13352 (N_13352,N_8715,N_8215);
nand U13353 (N_13353,N_9503,N_5361);
nor U13354 (N_13354,N_5395,N_5270);
or U13355 (N_13355,N_5224,N_9868);
nand U13356 (N_13356,N_5720,N_7684);
nand U13357 (N_13357,N_9715,N_9162);
and U13358 (N_13358,N_9307,N_6571);
and U13359 (N_13359,N_6295,N_6331);
nor U13360 (N_13360,N_6115,N_8978);
xor U13361 (N_13361,N_5230,N_5545);
or U13362 (N_13362,N_8883,N_8500);
nor U13363 (N_13363,N_9672,N_8298);
nand U13364 (N_13364,N_8876,N_5072);
nand U13365 (N_13365,N_7420,N_7625);
nor U13366 (N_13366,N_7584,N_5357);
nand U13367 (N_13367,N_8631,N_5127);
nand U13368 (N_13368,N_5804,N_9198);
nor U13369 (N_13369,N_7171,N_7688);
or U13370 (N_13370,N_5534,N_6156);
or U13371 (N_13371,N_9658,N_7974);
nand U13372 (N_13372,N_7299,N_8358);
nand U13373 (N_13373,N_6125,N_8289);
and U13374 (N_13374,N_6434,N_7576);
nand U13375 (N_13375,N_7682,N_5945);
nand U13376 (N_13376,N_9522,N_9983);
or U13377 (N_13377,N_7270,N_7916);
and U13378 (N_13378,N_6383,N_9573);
nand U13379 (N_13379,N_8401,N_6416);
and U13380 (N_13380,N_5572,N_8667);
nor U13381 (N_13381,N_7605,N_8721);
and U13382 (N_13382,N_7482,N_7907);
or U13383 (N_13383,N_7419,N_9775);
and U13384 (N_13384,N_5767,N_5157);
or U13385 (N_13385,N_8649,N_5393);
or U13386 (N_13386,N_7355,N_8424);
nand U13387 (N_13387,N_9435,N_6924);
or U13388 (N_13388,N_7988,N_7861);
or U13389 (N_13389,N_5417,N_5135);
or U13390 (N_13390,N_9584,N_8826);
nor U13391 (N_13391,N_8734,N_5133);
nor U13392 (N_13392,N_8256,N_8819);
nand U13393 (N_13393,N_9672,N_9445);
and U13394 (N_13394,N_9442,N_7400);
nor U13395 (N_13395,N_8123,N_5888);
and U13396 (N_13396,N_5054,N_7901);
or U13397 (N_13397,N_9811,N_9959);
nand U13398 (N_13398,N_9105,N_9968);
or U13399 (N_13399,N_7018,N_9564);
or U13400 (N_13400,N_5543,N_6947);
nor U13401 (N_13401,N_5229,N_5468);
nand U13402 (N_13402,N_9957,N_9780);
or U13403 (N_13403,N_6550,N_7896);
nor U13404 (N_13404,N_9139,N_8801);
or U13405 (N_13405,N_6514,N_8486);
nor U13406 (N_13406,N_8413,N_5127);
or U13407 (N_13407,N_9397,N_5240);
nand U13408 (N_13408,N_9118,N_9185);
xnor U13409 (N_13409,N_5552,N_5030);
nand U13410 (N_13410,N_8810,N_9314);
nor U13411 (N_13411,N_8997,N_9372);
nand U13412 (N_13412,N_6654,N_8903);
and U13413 (N_13413,N_8470,N_9672);
and U13414 (N_13414,N_9436,N_9836);
nor U13415 (N_13415,N_7363,N_8787);
and U13416 (N_13416,N_8836,N_9998);
and U13417 (N_13417,N_8887,N_9989);
and U13418 (N_13418,N_9774,N_9616);
and U13419 (N_13419,N_9863,N_8323);
nand U13420 (N_13420,N_9531,N_9960);
nand U13421 (N_13421,N_6347,N_7112);
nor U13422 (N_13422,N_6991,N_7275);
and U13423 (N_13423,N_9801,N_8935);
or U13424 (N_13424,N_8083,N_8508);
or U13425 (N_13425,N_7440,N_9206);
and U13426 (N_13426,N_9094,N_8184);
and U13427 (N_13427,N_7492,N_7305);
and U13428 (N_13428,N_8547,N_7722);
and U13429 (N_13429,N_7789,N_7301);
or U13430 (N_13430,N_7594,N_9778);
and U13431 (N_13431,N_6339,N_8814);
and U13432 (N_13432,N_9521,N_5668);
and U13433 (N_13433,N_5844,N_5806);
and U13434 (N_13434,N_7871,N_8249);
nor U13435 (N_13435,N_8721,N_6326);
nor U13436 (N_13436,N_5368,N_9091);
or U13437 (N_13437,N_8485,N_5362);
and U13438 (N_13438,N_7930,N_7718);
nand U13439 (N_13439,N_6455,N_9634);
or U13440 (N_13440,N_5168,N_7633);
nor U13441 (N_13441,N_8915,N_8913);
nor U13442 (N_13442,N_9348,N_5626);
nor U13443 (N_13443,N_5457,N_7583);
and U13444 (N_13444,N_5358,N_9447);
nand U13445 (N_13445,N_7740,N_7161);
nor U13446 (N_13446,N_8347,N_8251);
or U13447 (N_13447,N_9859,N_9536);
nand U13448 (N_13448,N_8699,N_8901);
nand U13449 (N_13449,N_7071,N_8796);
nand U13450 (N_13450,N_5300,N_6777);
nand U13451 (N_13451,N_7302,N_6804);
nor U13452 (N_13452,N_5221,N_8575);
or U13453 (N_13453,N_8573,N_9308);
nand U13454 (N_13454,N_6348,N_7656);
nand U13455 (N_13455,N_6532,N_5786);
nor U13456 (N_13456,N_9171,N_6542);
and U13457 (N_13457,N_7426,N_6004);
and U13458 (N_13458,N_9183,N_5751);
and U13459 (N_13459,N_7519,N_5227);
nand U13460 (N_13460,N_7785,N_7552);
and U13461 (N_13461,N_5945,N_6595);
and U13462 (N_13462,N_5386,N_5059);
nand U13463 (N_13463,N_9537,N_5108);
nand U13464 (N_13464,N_6023,N_9347);
nor U13465 (N_13465,N_8948,N_7262);
and U13466 (N_13466,N_8305,N_7283);
nand U13467 (N_13467,N_9825,N_5198);
and U13468 (N_13468,N_8408,N_8271);
nor U13469 (N_13469,N_7850,N_8674);
nand U13470 (N_13470,N_8536,N_7877);
nand U13471 (N_13471,N_5857,N_7505);
and U13472 (N_13472,N_9256,N_6793);
and U13473 (N_13473,N_7341,N_9143);
and U13474 (N_13474,N_8207,N_9476);
nor U13475 (N_13475,N_7080,N_9900);
nor U13476 (N_13476,N_5744,N_8787);
or U13477 (N_13477,N_9822,N_8799);
and U13478 (N_13478,N_6332,N_8262);
and U13479 (N_13479,N_6854,N_6373);
nor U13480 (N_13480,N_7647,N_6846);
or U13481 (N_13481,N_5050,N_9785);
nand U13482 (N_13482,N_6972,N_8431);
or U13483 (N_13483,N_5837,N_7885);
nand U13484 (N_13484,N_5770,N_9477);
nor U13485 (N_13485,N_6196,N_9671);
or U13486 (N_13486,N_8583,N_5833);
or U13487 (N_13487,N_6387,N_6336);
or U13488 (N_13488,N_5511,N_5894);
nor U13489 (N_13489,N_5091,N_8477);
or U13490 (N_13490,N_9794,N_9054);
and U13491 (N_13491,N_8151,N_8627);
nor U13492 (N_13492,N_5496,N_8338);
and U13493 (N_13493,N_8238,N_5467);
nor U13494 (N_13494,N_8450,N_9363);
nand U13495 (N_13495,N_5605,N_7164);
nor U13496 (N_13496,N_9915,N_8641);
nor U13497 (N_13497,N_6982,N_9388);
and U13498 (N_13498,N_6501,N_6469);
nand U13499 (N_13499,N_6975,N_9099);
and U13500 (N_13500,N_9049,N_9564);
nand U13501 (N_13501,N_7268,N_6193);
nand U13502 (N_13502,N_8898,N_8427);
nor U13503 (N_13503,N_5901,N_6257);
nand U13504 (N_13504,N_5984,N_9657);
nand U13505 (N_13505,N_9561,N_7018);
or U13506 (N_13506,N_6396,N_8884);
nor U13507 (N_13507,N_7761,N_8525);
xnor U13508 (N_13508,N_5511,N_9970);
nor U13509 (N_13509,N_6640,N_8738);
nor U13510 (N_13510,N_8333,N_5525);
or U13511 (N_13511,N_6101,N_9509);
nand U13512 (N_13512,N_9240,N_6164);
nor U13513 (N_13513,N_6581,N_5563);
xnor U13514 (N_13514,N_7792,N_6866);
or U13515 (N_13515,N_5762,N_9157);
nor U13516 (N_13516,N_6175,N_9254);
nor U13517 (N_13517,N_8369,N_6652);
nand U13518 (N_13518,N_8527,N_7894);
or U13519 (N_13519,N_7013,N_5417);
nand U13520 (N_13520,N_6889,N_6485);
nand U13521 (N_13521,N_5297,N_7843);
or U13522 (N_13522,N_5417,N_6462);
and U13523 (N_13523,N_7308,N_8392);
nand U13524 (N_13524,N_9670,N_5855);
and U13525 (N_13525,N_9600,N_6252);
nor U13526 (N_13526,N_9222,N_6601);
and U13527 (N_13527,N_5652,N_9623);
or U13528 (N_13528,N_8641,N_9100);
or U13529 (N_13529,N_7777,N_6301);
nor U13530 (N_13530,N_8791,N_9379);
or U13531 (N_13531,N_9173,N_8171);
and U13532 (N_13532,N_9491,N_7031);
and U13533 (N_13533,N_7159,N_7723);
nor U13534 (N_13534,N_7585,N_5779);
nor U13535 (N_13535,N_5331,N_6060);
or U13536 (N_13536,N_8182,N_7181);
nor U13537 (N_13537,N_8188,N_9690);
nor U13538 (N_13538,N_8720,N_8846);
and U13539 (N_13539,N_5555,N_6061);
and U13540 (N_13540,N_5593,N_8712);
nand U13541 (N_13541,N_7261,N_6491);
nand U13542 (N_13542,N_5402,N_6312);
nand U13543 (N_13543,N_7114,N_5742);
and U13544 (N_13544,N_9986,N_7062);
and U13545 (N_13545,N_5181,N_5644);
or U13546 (N_13546,N_7318,N_6358);
nand U13547 (N_13547,N_5231,N_5772);
nand U13548 (N_13548,N_9579,N_7309);
nor U13549 (N_13549,N_7330,N_8427);
nor U13550 (N_13550,N_7237,N_6165);
and U13551 (N_13551,N_5899,N_7075);
nor U13552 (N_13552,N_6317,N_6124);
nor U13553 (N_13553,N_7929,N_7767);
and U13554 (N_13554,N_8252,N_6006);
nor U13555 (N_13555,N_9330,N_5132);
nand U13556 (N_13556,N_8959,N_8621);
nor U13557 (N_13557,N_9455,N_9806);
nor U13558 (N_13558,N_6294,N_9972);
nand U13559 (N_13559,N_9379,N_6800);
and U13560 (N_13560,N_6128,N_6762);
nor U13561 (N_13561,N_6305,N_9550);
or U13562 (N_13562,N_6991,N_5985);
nand U13563 (N_13563,N_9389,N_5128);
nand U13564 (N_13564,N_6431,N_6546);
nand U13565 (N_13565,N_7112,N_6142);
or U13566 (N_13566,N_6243,N_8305);
nand U13567 (N_13567,N_7608,N_9605);
nand U13568 (N_13568,N_6214,N_6100);
and U13569 (N_13569,N_7953,N_5821);
and U13570 (N_13570,N_5362,N_9866);
nand U13571 (N_13571,N_8915,N_5648);
or U13572 (N_13572,N_8066,N_6957);
nand U13573 (N_13573,N_8166,N_9899);
nand U13574 (N_13574,N_6490,N_6056);
nor U13575 (N_13575,N_7043,N_7589);
or U13576 (N_13576,N_7661,N_8296);
or U13577 (N_13577,N_9542,N_5489);
nand U13578 (N_13578,N_6975,N_5644);
nor U13579 (N_13579,N_8444,N_9505);
nor U13580 (N_13580,N_8681,N_8730);
nand U13581 (N_13581,N_8299,N_9067);
or U13582 (N_13582,N_7718,N_9090);
or U13583 (N_13583,N_7346,N_8149);
and U13584 (N_13584,N_8074,N_6732);
nand U13585 (N_13585,N_7092,N_8704);
or U13586 (N_13586,N_8264,N_7471);
xnor U13587 (N_13587,N_9282,N_7978);
nor U13588 (N_13588,N_7178,N_7473);
nor U13589 (N_13589,N_6530,N_5733);
nor U13590 (N_13590,N_9098,N_8929);
nor U13591 (N_13591,N_8737,N_5762);
or U13592 (N_13592,N_5143,N_9750);
and U13593 (N_13593,N_6451,N_6581);
and U13594 (N_13594,N_9100,N_6758);
nor U13595 (N_13595,N_8290,N_8678);
nor U13596 (N_13596,N_8115,N_5438);
and U13597 (N_13597,N_9968,N_9201);
or U13598 (N_13598,N_8889,N_8368);
or U13599 (N_13599,N_7280,N_7158);
nor U13600 (N_13600,N_9480,N_8884);
or U13601 (N_13601,N_7356,N_7109);
or U13602 (N_13602,N_9156,N_7556);
nor U13603 (N_13603,N_9697,N_7615);
and U13604 (N_13604,N_8921,N_8278);
and U13605 (N_13605,N_9335,N_7200);
or U13606 (N_13606,N_7836,N_8909);
or U13607 (N_13607,N_6073,N_7159);
and U13608 (N_13608,N_7799,N_8026);
nand U13609 (N_13609,N_5289,N_6048);
and U13610 (N_13610,N_7965,N_9562);
nor U13611 (N_13611,N_5884,N_6466);
or U13612 (N_13612,N_8968,N_9986);
or U13613 (N_13613,N_9792,N_6158);
nand U13614 (N_13614,N_7468,N_6304);
or U13615 (N_13615,N_9385,N_9173);
nand U13616 (N_13616,N_8502,N_8518);
nor U13617 (N_13617,N_6009,N_5255);
or U13618 (N_13618,N_9896,N_6911);
nor U13619 (N_13619,N_6419,N_7127);
nand U13620 (N_13620,N_5309,N_5136);
and U13621 (N_13621,N_8523,N_7189);
nor U13622 (N_13622,N_5110,N_8410);
nand U13623 (N_13623,N_9107,N_9503);
and U13624 (N_13624,N_7028,N_7239);
nor U13625 (N_13625,N_9044,N_8877);
or U13626 (N_13626,N_8510,N_5985);
or U13627 (N_13627,N_6885,N_8429);
and U13628 (N_13628,N_8260,N_6797);
nand U13629 (N_13629,N_9763,N_8324);
nand U13630 (N_13630,N_7529,N_9739);
nand U13631 (N_13631,N_5158,N_5878);
or U13632 (N_13632,N_9947,N_8059);
nor U13633 (N_13633,N_7503,N_5534);
xor U13634 (N_13634,N_8479,N_6654);
or U13635 (N_13635,N_9442,N_8480);
nand U13636 (N_13636,N_7435,N_7474);
xnor U13637 (N_13637,N_6352,N_8075);
or U13638 (N_13638,N_9450,N_6698);
or U13639 (N_13639,N_7523,N_5338);
nand U13640 (N_13640,N_5544,N_9464);
or U13641 (N_13641,N_6507,N_7555);
and U13642 (N_13642,N_6699,N_9674);
and U13643 (N_13643,N_6690,N_5556);
xor U13644 (N_13644,N_8544,N_8796);
and U13645 (N_13645,N_7014,N_6311);
or U13646 (N_13646,N_8663,N_7174);
nand U13647 (N_13647,N_9970,N_5363);
nor U13648 (N_13648,N_5053,N_7065);
or U13649 (N_13649,N_9281,N_6401);
nand U13650 (N_13650,N_8807,N_8520);
and U13651 (N_13651,N_7544,N_8801);
or U13652 (N_13652,N_7998,N_9879);
nand U13653 (N_13653,N_9281,N_7053);
and U13654 (N_13654,N_9267,N_9733);
nor U13655 (N_13655,N_7189,N_9936);
and U13656 (N_13656,N_7289,N_5797);
nor U13657 (N_13657,N_8862,N_7119);
nand U13658 (N_13658,N_5904,N_7007);
or U13659 (N_13659,N_7078,N_5665);
and U13660 (N_13660,N_7281,N_8941);
and U13661 (N_13661,N_8430,N_9168);
nand U13662 (N_13662,N_5649,N_7262);
or U13663 (N_13663,N_8982,N_8228);
nand U13664 (N_13664,N_6708,N_6049);
nor U13665 (N_13665,N_5599,N_8149);
nor U13666 (N_13666,N_6560,N_7967);
and U13667 (N_13667,N_7484,N_5074);
or U13668 (N_13668,N_7160,N_9335);
or U13669 (N_13669,N_9795,N_7668);
and U13670 (N_13670,N_8783,N_6342);
or U13671 (N_13671,N_9079,N_6207);
nor U13672 (N_13672,N_6195,N_6835);
or U13673 (N_13673,N_6306,N_8850);
or U13674 (N_13674,N_7063,N_8337);
or U13675 (N_13675,N_9515,N_5413);
or U13676 (N_13676,N_5697,N_6468);
or U13677 (N_13677,N_7220,N_7377);
nor U13678 (N_13678,N_6949,N_7576);
nand U13679 (N_13679,N_8439,N_8470);
or U13680 (N_13680,N_7049,N_7849);
or U13681 (N_13681,N_9426,N_5773);
or U13682 (N_13682,N_7608,N_5810);
nand U13683 (N_13683,N_5122,N_7284);
and U13684 (N_13684,N_7329,N_5851);
or U13685 (N_13685,N_6840,N_9262);
or U13686 (N_13686,N_9061,N_8686);
and U13687 (N_13687,N_9401,N_9522);
nand U13688 (N_13688,N_5143,N_8813);
nand U13689 (N_13689,N_9702,N_6688);
and U13690 (N_13690,N_5593,N_9862);
and U13691 (N_13691,N_9626,N_5807);
or U13692 (N_13692,N_6639,N_5638);
or U13693 (N_13693,N_6788,N_8340);
or U13694 (N_13694,N_5206,N_8319);
and U13695 (N_13695,N_7826,N_9641);
and U13696 (N_13696,N_8363,N_9948);
nor U13697 (N_13697,N_6598,N_7379);
or U13698 (N_13698,N_6967,N_7209);
and U13699 (N_13699,N_5789,N_8363);
nand U13700 (N_13700,N_5092,N_9710);
and U13701 (N_13701,N_7444,N_7959);
or U13702 (N_13702,N_8662,N_8654);
or U13703 (N_13703,N_7516,N_8077);
nor U13704 (N_13704,N_7622,N_7151);
xnor U13705 (N_13705,N_6778,N_5564);
or U13706 (N_13706,N_5632,N_5439);
or U13707 (N_13707,N_6213,N_5490);
nor U13708 (N_13708,N_8393,N_8838);
nand U13709 (N_13709,N_7969,N_6321);
and U13710 (N_13710,N_9622,N_7557);
nor U13711 (N_13711,N_8417,N_7269);
or U13712 (N_13712,N_7731,N_6016);
nand U13713 (N_13713,N_5819,N_6109);
and U13714 (N_13714,N_9140,N_6487);
nor U13715 (N_13715,N_6231,N_7846);
nand U13716 (N_13716,N_7196,N_7936);
or U13717 (N_13717,N_9610,N_9044);
nor U13718 (N_13718,N_7170,N_6764);
nor U13719 (N_13719,N_7437,N_6566);
and U13720 (N_13720,N_7712,N_5232);
or U13721 (N_13721,N_6592,N_9642);
nand U13722 (N_13722,N_7375,N_5514);
nor U13723 (N_13723,N_9009,N_5090);
nor U13724 (N_13724,N_6088,N_8860);
or U13725 (N_13725,N_8234,N_9546);
nand U13726 (N_13726,N_7978,N_9511);
and U13727 (N_13727,N_9329,N_7913);
nand U13728 (N_13728,N_8929,N_8958);
or U13729 (N_13729,N_9962,N_5920);
and U13730 (N_13730,N_8603,N_7233);
nor U13731 (N_13731,N_6762,N_8794);
xor U13732 (N_13732,N_8577,N_6283);
or U13733 (N_13733,N_7899,N_8921);
or U13734 (N_13734,N_6324,N_8516);
nor U13735 (N_13735,N_7320,N_5495);
nor U13736 (N_13736,N_8546,N_8314);
nor U13737 (N_13737,N_5691,N_5531);
nor U13738 (N_13738,N_6027,N_8853);
nand U13739 (N_13739,N_9128,N_9213);
nor U13740 (N_13740,N_6959,N_8412);
nand U13741 (N_13741,N_9868,N_6958);
nor U13742 (N_13742,N_6296,N_8037);
and U13743 (N_13743,N_5476,N_9026);
nor U13744 (N_13744,N_7779,N_6162);
or U13745 (N_13745,N_7417,N_5724);
and U13746 (N_13746,N_9219,N_6837);
nand U13747 (N_13747,N_9185,N_8146);
nor U13748 (N_13748,N_9576,N_8418);
and U13749 (N_13749,N_9622,N_8654);
or U13750 (N_13750,N_8371,N_5644);
nor U13751 (N_13751,N_8447,N_5512);
and U13752 (N_13752,N_9115,N_8849);
and U13753 (N_13753,N_5305,N_8977);
nor U13754 (N_13754,N_5987,N_5910);
and U13755 (N_13755,N_9522,N_5337);
nand U13756 (N_13756,N_8706,N_5127);
nor U13757 (N_13757,N_8015,N_5307);
nand U13758 (N_13758,N_8771,N_8748);
or U13759 (N_13759,N_5779,N_5300);
nor U13760 (N_13760,N_5010,N_8539);
nand U13761 (N_13761,N_7610,N_6906);
and U13762 (N_13762,N_7293,N_6712);
and U13763 (N_13763,N_5517,N_8012);
nand U13764 (N_13764,N_9603,N_7332);
or U13765 (N_13765,N_7825,N_6934);
nand U13766 (N_13766,N_8624,N_8249);
nor U13767 (N_13767,N_9344,N_6621);
or U13768 (N_13768,N_9768,N_5257);
nor U13769 (N_13769,N_5136,N_9358);
nand U13770 (N_13770,N_7114,N_8477);
or U13771 (N_13771,N_8651,N_8739);
nand U13772 (N_13772,N_8749,N_5366);
or U13773 (N_13773,N_9188,N_6578);
and U13774 (N_13774,N_6469,N_7396);
and U13775 (N_13775,N_7295,N_9803);
or U13776 (N_13776,N_9003,N_9587);
xnor U13777 (N_13777,N_8280,N_8176);
and U13778 (N_13778,N_9612,N_9943);
and U13779 (N_13779,N_5071,N_8126);
nor U13780 (N_13780,N_5742,N_5052);
nand U13781 (N_13781,N_5877,N_9064);
or U13782 (N_13782,N_8673,N_8750);
xor U13783 (N_13783,N_9824,N_8865);
nor U13784 (N_13784,N_5897,N_9149);
or U13785 (N_13785,N_8349,N_7378);
nor U13786 (N_13786,N_7290,N_5065);
and U13787 (N_13787,N_9851,N_8396);
nor U13788 (N_13788,N_9336,N_6312);
and U13789 (N_13789,N_6536,N_8743);
or U13790 (N_13790,N_9845,N_6699);
or U13791 (N_13791,N_6472,N_7190);
and U13792 (N_13792,N_6841,N_6957);
or U13793 (N_13793,N_6789,N_6863);
or U13794 (N_13794,N_8140,N_6994);
nor U13795 (N_13795,N_9823,N_7119);
and U13796 (N_13796,N_6082,N_8422);
or U13797 (N_13797,N_9734,N_7421);
and U13798 (N_13798,N_7528,N_7482);
nor U13799 (N_13799,N_6693,N_6756);
nand U13800 (N_13800,N_5826,N_5289);
nor U13801 (N_13801,N_8001,N_5459);
or U13802 (N_13802,N_9689,N_5323);
nand U13803 (N_13803,N_6892,N_5769);
nor U13804 (N_13804,N_9674,N_9671);
and U13805 (N_13805,N_9447,N_5847);
nor U13806 (N_13806,N_5727,N_8977);
nand U13807 (N_13807,N_8176,N_7645);
and U13808 (N_13808,N_8708,N_7555);
nand U13809 (N_13809,N_7230,N_7415);
nand U13810 (N_13810,N_6748,N_9692);
nand U13811 (N_13811,N_7708,N_9531);
nor U13812 (N_13812,N_6591,N_5621);
or U13813 (N_13813,N_5226,N_8693);
nand U13814 (N_13814,N_8524,N_6127);
or U13815 (N_13815,N_5199,N_8758);
nor U13816 (N_13816,N_7128,N_7866);
nand U13817 (N_13817,N_5740,N_8458);
or U13818 (N_13818,N_8464,N_6617);
and U13819 (N_13819,N_6507,N_5840);
or U13820 (N_13820,N_6856,N_9060);
or U13821 (N_13821,N_6717,N_6933);
nand U13822 (N_13822,N_7771,N_6428);
and U13823 (N_13823,N_5172,N_6117);
xnor U13824 (N_13824,N_8698,N_8562);
or U13825 (N_13825,N_9655,N_5558);
or U13826 (N_13826,N_9953,N_7532);
nor U13827 (N_13827,N_5213,N_8335);
nand U13828 (N_13828,N_9415,N_8431);
nand U13829 (N_13829,N_5768,N_9452);
xor U13830 (N_13830,N_8739,N_5667);
nand U13831 (N_13831,N_6213,N_9695);
nor U13832 (N_13832,N_8912,N_6233);
or U13833 (N_13833,N_5240,N_9782);
nand U13834 (N_13834,N_5731,N_5898);
and U13835 (N_13835,N_7070,N_8050);
or U13836 (N_13836,N_8846,N_9171);
and U13837 (N_13837,N_5864,N_7431);
nor U13838 (N_13838,N_8698,N_5710);
nand U13839 (N_13839,N_6486,N_7094);
nor U13840 (N_13840,N_7628,N_5069);
or U13841 (N_13841,N_5977,N_5718);
and U13842 (N_13842,N_8363,N_5730);
nor U13843 (N_13843,N_8292,N_5470);
nand U13844 (N_13844,N_9736,N_6373);
or U13845 (N_13845,N_8453,N_5938);
or U13846 (N_13846,N_5192,N_6936);
and U13847 (N_13847,N_6322,N_5318);
nand U13848 (N_13848,N_5247,N_6540);
nand U13849 (N_13849,N_8361,N_8521);
or U13850 (N_13850,N_7186,N_7031);
and U13851 (N_13851,N_6350,N_9614);
nand U13852 (N_13852,N_7874,N_8484);
or U13853 (N_13853,N_6840,N_7549);
or U13854 (N_13854,N_5787,N_7324);
nor U13855 (N_13855,N_5053,N_7899);
nand U13856 (N_13856,N_7922,N_8028);
nand U13857 (N_13857,N_8735,N_7969);
and U13858 (N_13858,N_5771,N_7562);
and U13859 (N_13859,N_8155,N_5473);
nand U13860 (N_13860,N_7047,N_6678);
and U13861 (N_13861,N_9907,N_7074);
nor U13862 (N_13862,N_9343,N_9326);
nand U13863 (N_13863,N_5740,N_9133);
and U13864 (N_13864,N_9195,N_9294);
and U13865 (N_13865,N_6401,N_5209);
or U13866 (N_13866,N_9888,N_5111);
nand U13867 (N_13867,N_8842,N_6305);
and U13868 (N_13868,N_8355,N_8702);
nor U13869 (N_13869,N_5448,N_5592);
or U13870 (N_13870,N_9647,N_9362);
and U13871 (N_13871,N_6476,N_9192);
or U13872 (N_13872,N_7411,N_6424);
xnor U13873 (N_13873,N_7938,N_6932);
nor U13874 (N_13874,N_5082,N_8953);
xor U13875 (N_13875,N_8607,N_8117);
nor U13876 (N_13876,N_7961,N_7841);
or U13877 (N_13877,N_7901,N_9991);
or U13878 (N_13878,N_5450,N_9846);
nor U13879 (N_13879,N_6624,N_7034);
or U13880 (N_13880,N_6330,N_7922);
nor U13881 (N_13881,N_7801,N_7693);
nand U13882 (N_13882,N_5654,N_5152);
or U13883 (N_13883,N_5695,N_9995);
nor U13884 (N_13884,N_7720,N_9705);
or U13885 (N_13885,N_6381,N_5670);
nor U13886 (N_13886,N_7910,N_5735);
nand U13887 (N_13887,N_6011,N_9157);
nor U13888 (N_13888,N_5221,N_6152);
and U13889 (N_13889,N_8807,N_7458);
nor U13890 (N_13890,N_8059,N_9225);
and U13891 (N_13891,N_5665,N_8399);
nor U13892 (N_13892,N_5421,N_5885);
nand U13893 (N_13893,N_6886,N_6318);
and U13894 (N_13894,N_8351,N_6954);
nand U13895 (N_13895,N_6183,N_9944);
and U13896 (N_13896,N_9233,N_7849);
nor U13897 (N_13897,N_6509,N_8647);
or U13898 (N_13898,N_7247,N_7581);
nor U13899 (N_13899,N_7055,N_7699);
nand U13900 (N_13900,N_6223,N_9011);
nor U13901 (N_13901,N_8968,N_8075);
nand U13902 (N_13902,N_7367,N_9040);
nand U13903 (N_13903,N_6894,N_9415);
or U13904 (N_13904,N_8830,N_6228);
nand U13905 (N_13905,N_6370,N_8548);
nand U13906 (N_13906,N_8088,N_9070);
nand U13907 (N_13907,N_6174,N_9851);
nor U13908 (N_13908,N_5040,N_6713);
nand U13909 (N_13909,N_7172,N_7933);
nand U13910 (N_13910,N_7749,N_6716);
xor U13911 (N_13911,N_7448,N_5071);
and U13912 (N_13912,N_6364,N_7550);
nand U13913 (N_13913,N_5487,N_8210);
or U13914 (N_13914,N_7184,N_8601);
or U13915 (N_13915,N_6179,N_6762);
and U13916 (N_13916,N_6254,N_5275);
nand U13917 (N_13917,N_5535,N_6083);
nor U13918 (N_13918,N_9192,N_6233);
nand U13919 (N_13919,N_6548,N_7861);
and U13920 (N_13920,N_8720,N_6231);
and U13921 (N_13921,N_6869,N_5184);
or U13922 (N_13922,N_5794,N_5783);
nor U13923 (N_13923,N_6102,N_6776);
and U13924 (N_13924,N_8679,N_9093);
and U13925 (N_13925,N_7466,N_7397);
and U13926 (N_13926,N_5346,N_7909);
or U13927 (N_13927,N_8819,N_5541);
or U13928 (N_13928,N_6800,N_5072);
and U13929 (N_13929,N_5287,N_6338);
nand U13930 (N_13930,N_7700,N_7164);
or U13931 (N_13931,N_6407,N_5960);
or U13932 (N_13932,N_7824,N_5816);
nand U13933 (N_13933,N_9579,N_8975);
nand U13934 (N_13934,N_5941,N_9443);
nand U13935 (N_13935,N_6071,N_7478);
nor U13936 (N_13936,N_7172,N_9183);
nand U13937 (N_13937,N_9767,N_7728);
or U13938 (N_13938,N_8111,N_9673);
nand U13939 (N_13939,N_8329,N_7454);
nand U13940 (N_13940,N_9444,N_6693);
nand U13941 (N_13941,N_6716,N_7683);
or U13942 (N_13942,N_8667,N_9682);
nand U13943 (N_13943,N_5230,N_5817);
nand U13944 (N_13944,N_8046,N_6329);
nor U13945 (N_13945,N_8666,N_5846);
nor U13946 (N_13946,N_5103,N_8089);
nor U13947 (N_13947,N_7027,N_6881);
nand U13948 (N_13948,N_6024,N_9015);
or U13949 (N_13949,N_7672,N_5579);
and U13950 (N_13950,N_9742,N_6171);
nor U13951 (N_13951,N_5921,N_7499);
nand U13952 (N_13952,N_6458,N_9477);
nor U13953 (N_13953,N_6757,N_5894);
or U13954 (N_13954,N_5982,N_9379);
nand U13955 (N_13955,N_7086,N_6427);
or U13956 (N_13956,N_5871,N_9631);
nand U13957 (N_13957,N_6010,N_5305);
nand U13958 (N_13958,N_6712,N_6799);
or U13959 (N_13959,N_5721,N_6883);
nand U13960 (N_13960,N_6011,N_8618);
nor U13961 (N_13961,N_8469,N_9565);
and U13962 (N_13962,N_9998,N_8252);
or U13963 (N_13963,N_9033,N_6585);
and U13964 (N_13964,N_7247,N_6467);
and U13965 (N_13965,N_9015,N_7179);
nand U13966 (N_13966,N_5011,N_7262);
nor U13967 (N_13967,N_6619,N_8389);
and U13968 (N_13968,N_8170,N_5355);
and U13969 (N_13969,N_6340,N_8348);
nand U13970 (N_13970,N_5889,N_5851);
nand U13971 (N_13971,N_6841,N_9893);
or U13972 (N_13972,N_5776,N_7492);
nand U13973 (N_13973,N_6222,N_8288);
nand U13974 (N_13974,N_7807,N_5007);
and U13975 (N_13975,N_8670,N_5460);
nor U13976 (N_13976,N_7202,N_7492);
nor U13977 (N_13977,N_7482,N_9946);
and U13978 (N_13978,N_7029,N_7323);
nand U13979 (N_13979,N_9744,N_5779);
or U13980 (N_13980,N_6800,N_8178);
nand U13981 (N_13981,N_6460,N_7509);
nor U13982 (N_13982,N_6575,N_6313);
and U13983 (N_13983,N_5010,N_5609);
nand U13984 (N_13984,N_7143,N_6233);
nand U13985 (N_13985,N_6612,N_6424);
and U13986 (N_13986,N_6679,N_8074);
nor U13987 (N_13987,N_8665,N_7554);
nand U13988 (N_13988,N_9510,N_8303);
nand U13989 (N_13989,N_5161,N_6548);
or U13990 (N_13990,N_8240,N_7935);
nor U13991 (N_13991,N_7179,N_5764);
and U13992 (N_13992,N_8538,N_7738);
and U13993 (N_13993,N_9899,N_8948);
nand U13994 (N_13994,N_9120,N_5336);
or U13995 (N_13995,N_7985,N_5827);
and U13996 (N_13996,N_6205,N_9904);
and U13997 (N_13997,N_7138,N_8332);
nor U13998 (N_13998,N_8040,N_5705);
nor U13999 (N_13999,N_8255,N_9078);
nand U14000 (N_14000,N_8201,N_7310);
and U14001 (N_14001,N_9271,N_9525);
or U14002 (N_14002,N_5059,N_9266);
or U14003 (N_14003,N_6453,N_7745);
nand U14004 (N_14004,N_8960,N_7976);
nor U14005 (N_14005,N_7349,N_5441);
or U14006 (N_14006,N_6185,N_8243);
nand U14007 (N_14007,N_6738,N_6813);
and U14008 (N_14008,N_8924,N_5358);
or U14009 (N_14009,N_8139,N_8342);
nand U14010 (N_14010,N_6381,N_7790);
nor U14011 (N_14011,N_7765,N_8494);
nand U14012 (N_14012,N_6239,N_6017);
nor U14013 (N_14013,N_6184,N_5523);
and U14014 (N_14014,N_9297,N_8104);
nor U14015 (N_14015,N_6908,N_9027);
or U14016 (N_14016,N_5914,N_9176);
and U14017 (N_14017,N_8341,N_9553);
nand U14018 (N_14018,N_6383,N_6389);
and U14019 (N_14019,N_5071,N_5013);
and U14020 (N_14020,N_6606,N_5307);
or U14021 (N_14021,N_5786,N_6534);
nand U14022 (N_14022,N_5774,N_6917);
or U14023 (N_14023,N_7765,N_6432);
or U14024 (N_14024,N_7071,N_8658);
xnor U14025 (N_14025,N_7162,N_8459);
nand U14026 (N_14026,N_8611,N_6248);
nand U14027 (N_14027,N_8135,N_7585);
and U14028 (N_14028,N_5491,N_7181);
and U14029 (N_14029,N_6258,N_6484);
and U14030 (N_14030,N_5053,N_8046);
and U14031 (N_14031,N_9365,N_9625);
nor U14032 (N_14032,N_5740,N_9994);
or U14033 (N_14033,N_8947,N_6180);
and U14034 (N_14034,N_8581,N_5045);
nor U14035 (N_14035,N_6668,N_7503);
and U14036 (N_14036,N_7511,N_7064);
nand U14037 (N_14037,N_7662,N_6883);
nor U14038 (N_14038,N_7316,N_7581);
and U14039 (N_14039,N_7975,N_6012);
or U14040 (N_14040,N_6852,N_6127);
or U14041 (N_14041,N_5414,N_9056);
or U14042 (N_14042,N_7885,N_6783);
or U14043 (N_14043,N_5991,N_5322);
nor U14044 (N_14044,N_9722,N_7807);
and U14045 (N_14045,N_7399,N_9942);
nor U14046 (N_14046,N_7407,N_6287);
or U14047 (N_14047,N_6996,N_8446);
nor U14048 (N_14048,N_6586,N_5829);
nand U14049 (N_14049,N_8997,N_8156);
or U14050 (N_14050,N_9508,N_6874);
nand U14051 (N_14051,N_6745,N_7876);
nand U14052 (N_14052,N_5146,N_5919);
nand U14053 (N_14053,N_8802,N_5397);
or U14054 (N_14054,N_7529,N_8019);
nand U14055 (N_14055,N_7451,N_8154);
nand U14056 (N_14056,N_6848,N_5613);
and U14057 (N_14057,N_7024,N_7044);
nand U14058 (N_14058,N_9918,N_7968);
or U14059 (N_14059,N_6971,N_9200);
nand U14060 (N_14060,N_9289,N_8399);
and U14061 (N_14061,N_5127,N_9898);
and U14062 (N_14062,N_9360,N_9407);
nand U14063 (N_14063,N_9182,N_9675);
and U14064 (N_14064,N_7184,N_5246);
nand U14065 (N_14065,N_6251,N_9541);
nor U14066 (N_14066,N_9380,N_5998);
nand U14067 (N_14067,N_5555,N_9799);
nand U14068 (N_14068,N_8841,N_9850);
nand U14069 (N_14069,N_7986,N_5220);
and U14070 (N_14070,N_7085,N_5856);
nand U14071 (N_14071,N_7673,N_6597);
or U14072 (N_14072,N_6581,N_9689);
nor U14073 (N_14073,N_7186,N_7244);
nand U14074 (N_14074,N_5140,N_5268);
nand U14075 (N_14075,N_6937,N_5674);
nand U14076 (N_14076,N_7267,N_7985);
nand U14077 (N_14077,N_9661,N_9289);
or U14078 (N_14078,N_6534,N_5903);
or U14079 (N_14079,N_7428,N_9324);
nor U14080 (N_14080,N_8844,N_9312);
or U14081 (N_14081,N_6997,N_6641);
and U14082 (N_14082,N_5323,N_8505);
nand U14083 (N_14083,N_6339,N_6718);
and U14084 (N_14084,N_7445,N_6066);
and U14085 (N_14085,N_5201,N_9981);
or U14086 (N_14086,N_6496,N_7896);
or U14087 (N_14087,N_5518,N_9904);
or U14088 (N_14088,N_9575,N_9269);
or U14089 (N_14089,N_9237,N_8998);
nor U14090 (N_14090,N_5687,N_8311);
or U14091 (N_14091,N_9578,N_8888);
nor U14092 (N_14092,N_5919,N_8490);
and U14093 (N_14093,N_9448,N_7574);
or U14094 (N_14094,N_9703,N_7017);
nor U14095 (N_14095,N_8676,N_6111);
and U14096 (N_14096,N_7746,N_9443);
or U14097 (N_14097,N_7449,N_6465);
or U14098 (N_14098,N_7410,N_6701);
and U14099 (N_14099,N_6287,N_8712);
nor U14100 (N_14100,N_8662,N_8570);
nand U14101 (N_14101,N_8895,N_8898);
and U14102 (N_14102,N_7291,N_9004);
or U14103 (N_14103,N_8356,N_5464);
nand U14104 (N_14104,N_7070,N_8169);
nor U14105 (N_14105,N_7110,N_7031);
nor U14106 (N_14106,N_8795,N_8149);
nand U14107 (N_14107,N_7608,N_9290);
and U14108 (N_14108,N_5239,N_7066);
or U14109 (N_14109,N_6583,N_7119);
and U14110 (N_14110,N_8550,N_8825);
nand U14111 (N_14111,N_5851,N_8617);
or U14112 (N_14112,N_5690,N_8672);
and U14113 (N_14113,N_8618,N_6221);
and U14114 (N_14114,N_9547,N_9602);
nor U14115 (N_14115,N_7389,N_7168);
and U14116 (N_14116,N_6313,N_6064);
nor U14117 (N_14117,N_9884,N_8629);
nor U14118 (N_14118,N_5990,N_9750);
xnor U14119 (N_14119,N_8372,N_8034);
nand U14120 (N_14120,N_7847,N_6897);
nand U14121 (N_14121,N_7845,N_8539);
nand U14122 (N_14122,N_9150,N_8986);
nor U14123 (N_14123,N_7850,N_8871);
or U14124 (N_14124,N_5550,N_5376);
and U14125 (N_14125,N_5961,N_6489);
or U14126 (N_14126,N_6977,N_9560);
or U14127 (N_14127,N_6964,N_9244);
nand U14128 (N_14128,N_5601,N_7179);
nand U14129 (N_14129,N_7156,N_9847);
nor U14130 (N_14130,N_6477,N_6679);
or U14131 (N_14131,N_8747,N_8759);
or U14132 (N_14132,N_5131,N_6217);
nand U14133 (N_14133,N_5948,N_9788);
nand U14134 (N_14134,N_8112,N_9995);
and U14135 (N_14135,N_8367,N_8973);
nand U14136 (N_14136,N_7461,N_7457);
nand U14137 (N_14137,N_6360,N_8553);
nor U14138 (N_14138,N_5142,N_9367);
and U14139 (N_14139,N_7989,N_7680);
and U14140 (N_14140,N_7687,N_9787);
nand U14141 (N_14141,N_9175,N_7646);
nand U14142 (N_14142,N_5939,N_8079);
and U14143 (N_14143,N_7821,N_5632);
and U14144 (N_14144,N_7194,N_9863);
nand U14145 (N_14145,N_8638,N_7851);
and U14146 (N_14146,N_8866,N_5678);
nor U14147 (N_14147,N_8307,N_8967);
nor U14148 (N_14148,N_9518,N_5796);
nand U14149 (N_14149,N_9266,N_9705);
or U14150 (N_14150,N_6437,N_7250);
or U14151 (N_14151,N_7797,N_7956);
and U14152 (N_14152,N_8207,N_8372);
or U14153 (N_14153,N_5174,N_7835);
nand U14154 (N_14154,N_5739,N_8378);
and U14155 (N_14155,N_5861,N_9734);
and U14156 (N_14156,N_6445,N_6718);
nand U14157 (N_14157,N_9760,N_8458);
nor U14158 (N_14158,N_9498,N_9065);
xnor U14159 (N_14159,N_8540,N_9770);
nor U14160 (N_14160,N_8725,N_7037);
or U14161 (N_14161,N_5762,N_5693);
or U14162 (N_14162,N_9959,N_7073);
or U14163 (N_14163,N_5241,N_8185);
and U14164 (N_14164,N_5406,N_9671);
nand U14165 (N_14165,N_9003,N_5208);
and U14166 (N_14166,N_5178,N_5365);
and U14167 (N_14167,N_8079,N_8409);
or U14168 (N_14168,N_5311,N_6627);
or U14169 (N_14169,N_8816,N_9107);
or U14170 (N_14170,N_6254,N_5857);
and U14171 (N_14171,N_6508,N_8934);
and U14172 (N_14172,N_7100,N_8392);
nand U14173 (N_14173,N_5442,N_7404);
or U14174 (N_14174,N_8134,N_6899);
and U14175 (N_14175,N_6570,N_5881);
or U14176 (N_14176,N_5459,N_7380);
and U14177 (N_14177,N_9179,N_7076);
or U14178 (N_14178,N_8753,N_8876);
nand U14179 (N_14179,N_6419,N_9820);
or U14180 (N_14180,N_8005,N_7813);
nor U14181 (N_14181,N_5431,N_7905);
or U14182 (N_14182,N_8189,N_5520);
and U14183 (N_14183,N_9670,N_6966);
and U14184 (N_14184,N_5193,N_6488);
nor U14185 (N_14185,N_9306,N_8752);
nor U14186 (N_14186,N_5114,N_8640);
nor U14187 (N_14187,N_8639,N_5545);
nor U14188 (N_14188,N_6777,N_6870);
nor U14189 (N_14189,N_7153,N_9863);
or U14190 (N_14190,N_9297,N_6740);
or U14191 (N_14191,N_9794,N_9579);
and U14192 (N_14192,N_8082,N_7382);
nand U14193 (N_14193,N_6706,N_6786);
nand U14194 (N_14194,N_8287,N_7309);
or U14195 (N_14195,N_8134,N_7288);
nor U14196 (N_14196,N_9227,N_7502);
nor U14197 (N_14197,N_9138,N_7525);
nand U14198 (N_14198,N_6764,N_8268);
nand U14199 (N_14199,N_5162,N_6371);
nand U14200 (N_14200,N_8286,N_6159);
nor U14201 (N_14201,N_8778,N_6074);
and U14202 (N_14202,N_7467,N_8183);
nand U14203 (N_14203,N_7761,N_5207);
and U14204 (N_14204,N_5425,N_7997);
or U14205 (N_14205,N_6160,N_5642);
and U14206 (N_14206,N_8307,N_9776);
and U14207 (N_14207,N_9508,N_5072);
nor U14208 (N_14208,N_6011,N_5399);
or U14209 (N_14209,N_7874,N_6295);
and U14210 (N_14210,N_8858,N_6420);
and U14211 (N_14211,N_9477,N_9390);
nor U14212 (N_14212,N_5657,N_8142);
nand U14213 (N_14213,N_6012,N_9320);
or U14214 (N_14214,N_6981,N_6798);
nand U14215 (N_14215,N_7375,N_7432);
nor U14216 (N_14216,N_9599,N_8196);
nand U14217 (N_14217,N_8345,N_9732);
nor U14218 (N_14218,N_9869,N_5273);
and U14219 (N_14219,N_7600,N_6590);
xnor U14220 (N_14220,N_8716,N_6337);
and U14221 (N_14221,N_8187,N_9463);
and U14222 (N_14222,N_6395,N_8562);
or U14223 (N_14223,N_5451,N_8612);
nand U14224 (N_14224,N_9276,N_9057);
and U14225 (N_14225,N_5217,N_8895);
nor U14226 (N_14226,N_9913,N_8646);
or U14227 (N_14227,N_9393,N_8307);
and U14228 (N_14228,N_7481,N_5959);
or U14229 (N_14229,N_6166,N_8114);
and U14230 (N_14230,N_6438,N_7818);
nor U14231 (N_14231,N_7490,N_7959);
or U14232 (N_14232,N_7391,N_7814);
nand U14233 (N_14233,N_5100,N_9394);
or U14234 (N_14234,N_7786,N_5423);
or U14235 (N_14235,N_6298,N_8779);
nand U14236 (N_14236,N_7697,N_8426);
and U14237 (N_14237,N_6307,N_5249);
or U14238 (N_14238,N_9904,N_8148);
or U14239 (N_14239,N_6332,N_7971);
nor U14240 (N_14240,N_6354,N_9208);
or U14241 (N_14241,N_5972,N_8318);
and U14242 (N_14242,N_6405,N_8940);
or U14243 (N_14243,N_7967,N_8493);
nand U14244 (N_14244,N_9980,N_7629);
and U14245 (N_14245,N_9423,N_6033);
nor U14246 (N_14246,N_6799,N_7060);
and U14247 (N_14247,N_6898,N_7950);
nor U14248 (N_14248,N_5150,N_5686);
nor U14249 (N_14249,N_8738,N_7095);
nand U14250 (N_14250,N_9992,N_5724);
nor U14251 (N_14251,N_6744,N_6016);
or U14252 (N_14252,N_6253,N_7127);
nor U14253 (N_14253,N_9170,N_5014);
nand U14254 (N_14254,N_7640,N_6993);
or U14255 (N_14255,N_6518,N_5328);
xor U14256 (N_14256,N_9298,N_7911);
or U14257 (N_14257,N_8081,N_9979);
nand U14258 (N_14258,N_8714,N_5640);
and U14259 (N_14259,N_8124,N_6168);
or U14260 (N_14260,N_8876,N_8222);
nor U14261 (N_14261,N_8141,N_8663);
xnor U14262 (N_14262,N_9276,N_5514);
nor U14263 (N_14263,N_9251,N_7287);
nor U14264 (N_14264,N_7684,N_5580);
or U14265 (N_14265,N_5328,N_9082);
nor U14266 (N_14266,N_5248,N_8459);
nand U14267 (N_14267,N_7248,N_6197);
nor U14268 (N_14268,N_6043,N_7085);
nor U14269 (N_14269,N_7414,N_9008);
nor U14270 (N_14270,N_9474,N_9789);
nand U14271 (N_14271,N_7420,N_8630);
nor U14272 (N_14272,N_8635,N_9784);
and U14273 (N_14273,N_7453,N_7404);
nand U14274 (N_14274,N_6632,N_7546);
nor U14275 (N_14275,N_8940,N_7037);
nand U14276 (N_14276,N_6408,N_5937);
or U14277 (N_14277,N_6995,N_9774);
or U14278 (N_14278,N_8456,N_7845);
or U14279 (N_14279,N_9389,N_5565);
nand U14280 (N_14280,N_5692,N_8330);
or U14281 (N_14281,N_7544,N_8530);
or U14282 (N_14282,N_8276,N_6711);
or U14283 (N_14283,N_9706,N_8208);
and U14284 (N_14284,N_6948,N_7146);
and U14285 (N_14285,N_8939,N_6455);
nand U14286 (N_14286,N_7277,N_5770);
nor U14287 (N_14287,N_8903,N_9334);
or U14288 (N_14288,N_7350,N_7774);
or U14289 (N_14289,N_8071,N_9033);
nor U14290 (N_14290,N_8803,N_6776);
or U14291 (N_14291,N_8422,N_9997);
or U14292 (N_14292,N_8698,N_8905);
and U14293 (N_14293,N_6815,N_5846);
nand U14294 (N_14294,N_5732,N_8745);
nor U14295 (N_14295,N_6127,N_6896);
nor U14296 (N_14296,N_7690,N_9435);
nand U14297 (N_14297,N_5674,N_9290);
or U14298 (N_14298,N_9294,N_8661);
or U14299 (N_14299,N_9021,N_7862);
or U14300 (N_14300,N_6313,N_7334);
nand U14301 (N_14301,N_7993,N_5103);
nor U14302 (N_14302,N_8515,N_5851);
or U14303 (N_14303,N_7152,N_9037);
or U14304 (N_14304,N_9825,N_8274);
or U14305 (N_14305,N_6381,N_5461);
and U14306 (N_14306,N_7704,N_9174);
nor U14307 (N_14307,N_7163,N_6519);
nor U14308 (N_14308,N_8632,N_5977);
or U14309 (N_14309,N_9231,N_9507);
or U14310 (N_14310,N_9710,N_9621);
nor U14311 (N_14311,N_5027,N_5943);
and U14312 (N_14312,N_8267,N_5660);
xor U14313 (N_14313,N_9329,N_6012);
and U14314 (N_14314,N_7936,N_9607);
and U14315 (N_14315,N_7955,N_6067);
or U14316 (N_14316,N_7506,N_8676);
or U14317 (N_14317,N_6889,N_8195);
and U14318 (N_14318,N_8813,N_5424);
nor U14319 (N_14319,N_9613,N_5186);
nor U14320 (N_14320,N_6078,N_9822);
xor U14321 (N_14321,N_7484,N_6019);
or U14322 (N_14322,N_5072,N_7605);
nand U14323 (N_14323,N_7687,N_7334);
nor U14324 (N_14324,N_7731,N_8523);
nand U14325 (N_14325,N_6437,N_6280);
and U14326 (N_14326,N_6060,N_5351);
nand U14327 (N_14327,N_9539,N_7370);
nand U14328 (N_14328,N_8253,N_8965);
and U14329 (N_14329,N_7271,N_5664);
and U14330 (N_14330,N_7667,N_9721);
or U14331 (N_14331,N_5141,N_7799);
nor U14332 (N_14332,N_7127,N_8940);
or U14333 (N_14333,N_9193,N_9237);
nor U14334 (N_14334,N_7367,N_8504);
nor U14335 (N_14335,N_6040,N_5885);
nor U14336 (N_14336,N_8414,N_8807);
nand U14337 (N_14337,N_6889,N_9762);
nor U14338 (N_14338,N_6281,N_6823);
and U14339 (N_14339,N_7782,N_6063);
or U14340 (N_14340,N_6298,N_9363);
or U14341 (N_14341,N_7127,N_6601);
nor U14342 (N_14342,N_6631,N_8661);
and U14343 (N_14343,N_6101,N_7995);
or U14344 (N_14344,N_7070,N_7972);
nor U14345 (N_14345,N_8460,N_9101);
nand U14346 (N_14346,N_8006,N_5524);
and U14347 (N_14347,N_8347,N_7800);
nor U14348 (N_14348,N_5439,N_7390);
or U14349 (N_14349,N_9371,N_9448);
and U14350 (N_14350,N_9672,N_6563);
nor U14351 (N_14351,N_6963,N_6641);
or U14352 (N_14352,N_6210,N_7003);
nand U14353 (N_14353,N_9192,N_8537);
nor U14354 (N_14354,N_8588,N_5695);
nor U14355 (N_14355,N_5968,N_9985);
nor U14356 (N_14356,N_5133,N_9155);
nor U14357 (N_14357,N_9593,N_5031);
and U14358 (N_14358,N_7482,N_5241);
nor U14359 (N_14359,N_9995,N_5406);
or U14360 (N_14360,N_6495,N_5286);
and U14361 (N_14361,N_6510,N_7779);
and U14362 (N_14362,N_7207,N_8640);
nand U14363 (N_14363,N_5842,N_7229);
nor U14364 (N_14364,N_9630,N_8007);
nand U14365 (N_14365,N_6182,N_5778);
nor U14366 (N_14366,N_6615,N_6447);
or U14367 (N_14367,N_6341,N_9271);
or U14368 (N_14368,N_8243,N_9042);
and U14369 (N_14369,N_6570,N_6956);
nor U14370 (N_14370,N_7721,N_8904);
and U14371 (N_14371,N_8415,N_5301);
nand U14372 (N_14372,N_6373,N_9252);
and U14373 (N_14373,N_9166,N_6686);
and U14374 (N_14374,N_9464,N_5935);
nor U14375 (N_14375,N_6883,N_7156);
and U14376 (N_14376,N_9404,N_6275);
or U14377 (N_14377,N_6564,N_9181);
or U14378 (N_14378,N_9304,N_9548);
nor U14379 (N_14379,N_7112,N_5003);
xor U14380 (N_14380,N_8114,N_8521);
or U14381 (N_14381,N_9906,N_8760);
or U14382 (N_14382,N_5991,N_6965);
nor U14383 (N_14383,N_5440,N_9997);
or U14384 (N_14384,N_6473,N_7065);
nor U14385 (N_14385,N_9378,N_9421);
and U14386 (N_14386,N_5618,N_7663);
nor U14387 (N_14387,N_8296,N_7452);
and U14388 (N_14388,N_7238,N_6351);
or U14389 (N_14389,N_8868,N_7956);
or U14390 (N_14390,N_7034,N_6960);
or U14391 (N_14391,N_5527,N_9587);
nand U14392 (N_14392,N_5727,N_8473);
nor U14393 (N_14393,N_9870,N_8015);
and U14394 (N_14394,N_8708,N_9173);
or U14395 (N_14395,N_6235,N_9578);
nor U14396 (N_14396,N_6583,N_6635);
nor U14397 (N_14397,N_8648,N_6687);
nor U14398 (N_14398,N_6465,N_7037);
and U14399 (N_14399,N_9487,N_5155);
or U14400 (N_14400,N_5074,N_6078);
and U14401 (N_14401,N_9712,N_7466);
nor U14402 (N_14402,N_7731,N_5873);
and U14403 (N_14403,N_7824,N_8210);
and U14404 (N_14404,N_7299,N_9897);
nor U14405 (N_14405,N_5359,N_7359);
and U14406 (N_14406,N_7778,N_6587);
nor U14407 (N_14407,N_6111,N_5696);
nor U14408 (N_14408,N_9015,N_8463);
or U14409 (N_14409,N_6076,N_9317);
and U14410 (N_14410,N_6007,N_9742);
nand U14411 (N_14411,N_6191,N_5520);
nor U14412 (N_14412,N_9704,N_5808);
and U14413 (N_14413,N_6917,N_8531);
nor U14414 (N_14414,N_8090,N_9066);
nor U14415 (N_14415,N_7576,N_7854);
or U14416 (N_14416,N_8781,N_6516);
nor U14417 (N_14417,N_6247,N_7522);
and U14418 (N_14418,N_5186,N_8572);
and U14419 (N_14419,N_9602,N_6461);
and U14420 (N_14420,N_9010,N_7623);
and U14421 (N_14421,N_8560,N_8873);
nor U14422 (N_14422,N_5637,N_6655);
or U14423 (N_14423,N_8057,N_6610);
xor U14424 (N_14424,N_8565,N_7264);
or U14425 (N_14425,N_9841,N_8512);
or U14426 (N_14426,N_9504,N_8291);
nor U14427 (N_14427,N_9805,N_7208);
and U14428 (N_14428,N_5924,N_6282);
nor U14429 (N_14429,N_5018,N_9765);
and U14430 (N_14430,N_9614,N_9044);
nor U14431 (N_14431,N_7836,N_5009);
nand U14432 (N_14432,N_6648,N_8085);
and U14433 (N_14433,N_5746,N_8570);
or U14434 (N_14434,N_7980,N_9126);
nand U14435 (N_14435,N_9664,N_9731);
and U14436 (N_14436,N_5560,N_7028);
and U14437 (N_14437,N_5334,N_9216);
nor U14438 (N_14438,N_5249,N_9715);
or U14439 (N_14439,N_7350,N_9832);
and U14440 (N_14440,N_9311,N_8628);
or U14441 (N_14441,N_6736,N_8917);
nand U14442 (N_14442,N_9224,N_5298);
and U14443 (N_14443,N_5142,N_7403);
nor U14444 (N_14444,N_7426,N_9887);
nand U14445 (N_14445,N_8438,N_8081);
nand U14446 (N_14446,N_5035,N_6245);
and U14447 (N_14447,N_5122,N_5220);
or U14448 (N_14448,N_5169,N_7999);
or U14449 (N_14449,N_6662,N_7036);
or U14450 (N_14450,N_5084,N_6211);
nor U14451 (N_14451,N_5648,N_8564);
or U14452 (N_14452,N_7958,N_6027);
nor U14453 (N_14453,N_5945,N_9170);
nand U14454 (N_14454,N_8522,N_7014);
nor U14455 (N_14455,N_5876,N_5920);
nand U14456 (N_14456,N_9969,N_5518);
nand U14457 (N_14457,N_5514,N_9983);
nor U14458 (N_14458,N_7907,N_8193);
and U14459 (N_14459,N_6521,N_5842);
nand U14460 (N_14460,N_5539,N_9011);
xnor U14461 (N_14461,N_9756,N_6235);
and U14462 (N_14462,N_8036,N_7959);
and U14463 (N_14463,N_6901,N_9279);
or U14464 (N_14464,N_9914,N_7042);
and U14465 (N_14465,N_7358,N_8916);
and U14466 (N_14466,N_9889,N_7714);
nand U14467 (N_14467,N_9419,N_5677);
or U14468 (N_14468,N_6512,N_5536);
and U14469 (N_14469,N_5367,N_9836);
nand U14470 (N_14470,N_5815,N_5916);
nor U14471 (N_14471,N_6204,N_9649);
nor U14472 (N_14472,N_6044,N_5705);
nor U14473 (N_14473,N_5177,N_5760);
nand U14474 (N_14474,N_8447,N_9039);
nand U14475 (N_14475,N_7948,N_5743);
or U14476 (N_14476,N_7640,N_8701);
and U14477 (N_14477,N_7976,N_8068);
and U14478 (N_14478,N_8720,N_6199);
nor U14479 (N_14479,N_5384,N_6962);
and U14480 (N_14480,N_5958,N_9623);
nor U14481 (N_14481,N_8432,N_5177);
and U14482 (N_14482,N_8640,N_5372);
and U14483 (N_14483,N_8984,N_9255);
nor U14484 (N_14484,N_8699,N_5920);
and U14485 (N_14485,N_8390,N_5395);
and U14486 (N_14486,N_5613,N_7669);
nor U14487 (N_14487,N_9422,N_7185);
and U14488 (N_14488,N_8648,N_5390);
and U14489 (N_14489,N_9960,N_7982);
nor U14490 (N_14490,N_5448,N_5439);
and U14491 (N_14491,N_8447,N_6331);
and U14492 (N_14492,N_8653,N_6536);
nor U14493 (N_14493,N_5371,N_9639);
or U14494 (N_14494,N_9236,N_8913);
xnor U14495 (N_14495,N_5416,N_5604);
and U14496 (N_14496,N_5892,N_5079);
nand U14497 (N_14497,N_9355,N_9955);
and U14498 (N_14498,N_9050,N_8394);
nand U14499 (N_14499,N_6223,N_9486);
and U14500 (N_14500,N_9672,N_5622);
nand U14501 (N_14501,N_5815,N_6306);
or U14502 (N_14502,N_6674,N_6322);
xor U14503 (N_14503,N_9690,N_8291);
nand U14504 (N_14504,N_8880,N_9173);
and U14505 (N_14505,N_7365,N_5501);
and U14506 (N_14506,N_5802,N_5348);
nor U14507 (N_14507,N_9931,N_9572);
and U14508 (N_14508,N_8226,N_7122);
or U14509 (N_14509,N_7808,N_5167);
or U14510 (N_14510,N_8337,N_7267);
or U14511 (N_14511,N_9235,N_5405);
and U14512 (N_14512,N_9439,N_5127);
and U14513 (N_14513,N_5337,N_7089);
or U14514 (N_14514,N_6938,N_8119);
nor U14515 (N_14515,N_7034,N_6874);
nor U14516 (N_14516,N_8397,N_7694);
or U14517 (N_14517,N_7245,N_5909);
and U14518 (N_14518,N_7578,N_9428);
and U14519 (N_14519,N_8573,N_7122);
nor U14520 (N_14520,N_7692,N_6251);
nor U14521 (N_14521,N_8371,N_9819);
nand U14522 (N_14522,N_7755,N_6873);
and U14523 (N_14523,N_6141,N_7035);
and U14524 (N_14524,N_7326,N_8967);
xnor U14525 (N_14525,N_7781,N_7017);
nor U14526 (N_14526,N_7146,N_8573);
nor U14527 (N_14527,N_7462,N_5079);
nor U14528 (N_14528,N_5082,N_7761);
nand U14529 (N_14529,N_9167,N_7748);
nor U14530 (N_14530,N_7616,N_6795);
nor U14531 (N_14531,N_5991,N_9126);
nor U14532 (N_14532,N_8002,N_6481);
nand U14533 (N_14533,N_5869,N_5442);
nand U14534 (N_14534,N_9317,N_5223);
nand U14535 (N_14535,N_8304,N_8727);
nand U14536 (N_14536,N_9928,N_9043);
nor U14537 (N_14537,N_6102,N_7208);
nor U14538 (N_14538,N_9549,N_8609);
or U14539 (N_14539,N_9820,N_7547);
and U14540 (N_14540,N_9815,N_8553);
nor U14541 (N_14541,N_6843,N_6095);
and U14542 (N_14542,N_9328,N_7374);
or U14543 (N_14543,N_6626,N_9715);
or U14544 (N_14544,N_5589,N_6142);
nand U14545 (N_14545,N_6653,N_6270);
nand U14546 (N_14546,N_6828,N_5765);
nand U14547 (N_14547,N_7013,N_6202);
or U14548 (N_14548,N_6920,N_9746);
nor U14549 (N_14549,N_8525,N_9943);
nor U14550 (N_14550,N_9649,N_9887);
or U14551 (N_14551,N_6712,N_7645);
and U14552 (N_14552,N_7853,N_6915);
nand U14553 (N_14553,N_9413,N_7603);
nor U14554 (N_14554,N_9885,N_9924);
nand U14555 (N_14555,N_5208,N_6732);
or U14556 (N_14556,N_7636,N_6278);
and U14557 (N_14557,N_5195,N_6712);
and U14558 (N_14558,N_7245,N_5531);
and U14559 (N_14559,N_9058,N_9075);
and U14560 (N_14560,N_7291,N_8945);
nand U14561 (N_14561,N_7517,N_9286);
and U14562 (N_14562,N_9685,N_6514);
nand U14563 (N_14563,N_7350,N_7783);
or U14564 (N_14564,N_7804,N_6229);
nand U14565 (N_14565,N_5520,N_7049);
nor U14566 (N_14566,N_9086,N_6434);
and U14567 (N_14567,N_8709,N_9341);
nor U14568 (N_14568,N_8727,N_9131);
nor U14569 (N_14569,N_7069,N_7365);
or U14570 (N_14570,N_6288,N_5779);
xnor U14571 (N_14571,N_8445,N_6167);
or U14572 (N_14572,N_6612,N_6910);
and U14573 (N_14573,N_7156,N_8637);
or U14574 (N_14574,N_9878,N_8053);
and U14575 (N_14575,N_8930,N_9024);
and U14576 (N_14576,N_5013,N_6116);
nand U14577 (N_14577,N_5428,N_8471);
and U14578 (N_14578,N_6942,N_9656);
nor U14579 (N_14579,N_9168,N_6320);
or U14580 (N_14580,N_9052,N_8161);
and U14581 (N_14581,N_9013,N_6584);
and U14582 (N_14582,N_8239,N_9532);
nor U14583 (N_14583,N_8571,N_7735);
or U14584 (N_14584,N_8897,N_9478);
or U14585 (N_14585,N_5804,N_8293);
and U14586 (N_14586,N_8452,N_8920);
or U14587 (N_14587,N_5891,N_9633);
and U14588 (N_14588,N_7272,N_8765);
nor U14589 (N_14589,N_5451,N_6868);
nand U14590 (N_14590,N_5290,N_6477);
nand U14591 (N_14591,N_7735,N_7669);
and U14592 (N_14592,N_6993,N_5627);
or U14593 (N_14593,N_7305,N_9942);
and U14594 (N_14594,N_9182,N_6106);
or U14595 (N_14595,N_7314,N_6282);
nand U14596 (N_14596,N_7378,N_9325);
or U14597 (N_14597,N_5731,N_7389);
and U14598 (N_14598,N_8896,N_8501);
nand U14599 (N_14599,N_8494,N_5947);
or U14600 (N_14600,N_6574,N_7067);
and U14601 (N_14601,N_9617,N_5330);
nand U14602 (N_14602,N_7136,N_9331);
or U14603 (N_14603,N_6940,N_5626);
and U14604 (N_14604,N_6399,N_6975);
nor U14605 (N_14605,N_9136,N_7668);
nor U14606 (N_14606,N_7571,N_9673);
nand U14607 (N_14607,N_7138,N_7914);
nor U14608 (N_14608,N_9511,N_7772);
nor U14609 (N_14609,N_5660,N_9938);
nor U14610 (N_14610,N_5315,N_7661);
nor U14611 (N_14611,N_9206,N_8280);
nor U14612 (N_14612,N_8983,N_5792);
or U14613 (N_14613,N_9615,N_9445);
nor U14614 (N_14614,N_8832,N_5118);
xnor U14615 (N_14615,N_6202,N_8179);
or U14616 (N_14616,N_6500,N_9690);
nand U14617 (N_14617,N_8157,N_5337);
nand U14618 (N_14618,N_9090,N_6471);
nor U14619 (N_14619,N_9714,N_8062);
nor U14620 (N_14620,N_9942,N_8589);
nand U14621 (N_14621,N_7363,N_8578);
nor U14622 (N_14622,N_8661,N_9984);
or U14623 (N_14623,N_8915,N_7810);
and U14624 (N_14624,N_9899,N_5306);
nor U14625 (N_14625,N_8350,N_9656);
and U14626 (N_14626,N_5209,N_8127);
xnor U14627 (N_14627,N_8594,N_6375);
or U14628 (N_14628,N_6691,N_7575);
nor U14629 (N_14629,N_5446,N_9710);
nor U14630 (N_14630,N_6867,N_9872);
and U14631 (N_14631,N_7256,N_7965);
nand U14632 (N_14632,N_7937,N_8925);
xor U14633 (N_14633,N_5730,N_7079);
nor U14634 (N_14634,N_5782,N_9224);
or U14635 (N_14635,N_8812,N_6457);
nand U14636 (N_14636,N_9007,N_7513);
and U14637 (N_14637,N_6989,N_6749);
and U14638 (N_14638,N_5323,N_8361);
nand U14639 (N_14639,N_7473,N_8201);
and U14640 (N_14640,N_7546,N_9825);
or U14641 (N_14641,N_7881,N_7555);
or U14642 (N_14642,N_8870,N_5232);
and U14643 (N_14643,N_9490,N_9849);
or U14644 (N_14644,N_7425,N_6425);
and U14645 (N_14645,N_5432,N_6281);
or U14646 (N_14646,N_7143,N_6348);
and U14647 (N_14647,N_8502,N_6133);
and U14648 (N_14648,N_9565,N_8435);
and U14649 (N_14649,N_8837,N_9574);
nand U14650 (N_14650,N_7560,N_7656);
or U14651 (N_14651,N_5384,N_5953);
and U14652 (N_14652,N_9789,N_6772);
nand U14653 (N_14653,N_9675,N_6939);
or U14654 (N_14654,N_9667,N_7961);
nor U14655 (N_14655,N_8487,N_5353);
and U14656 (N_14656,N_7087,N_6375);
and U14657 (N_14657,N_8422,N_6510);
and U14658 (N_14658,N_5794,N_6512);
nor U14659 (N_14659,N_9659,N_6168);
nand U14660 (N_14660,N_8731,N_9922);
or U14661 (N_14661,N_8358,N_8290);
or U14662 (N_14662,N_8445,N_9470);
or U14663 (N_14663,N_5472,N_5036);
or U14664 (N_14664,N_8711,N_9662);
nor U14665 (N_14665,N_8272,N_7807);
nor U14666 (N_14666,N_9691,N_8237);
or U14667 (N_14667,N_5740,N_8294);
nand U14668 (N_14668,N_6651,N_5866);
and U14669 (N_14669,N_9404,N_6070);
or U14670 (N_14670,N_9772,N_8526);
xor U14671 (N_14671,N_8302,N_6103);
nor U14672 (N_14672,N_9879,N_8871);
and U14673 (N_14673,N_7626,N_5655);
and U14674 (N_14674,N_6182,N_8456);
or U14675 (N_14675,N_5247,N_5275);
and U14676 (N_14676,N_9903,N_6917);
nand U14677 (N_14677,N_5735,N_9228);
or U14678 (N_14678,N_7647,N_6163);
or U14679 (N_14679,N_5949,N_7704);
nand U14680 (N_14680,N_5538,N_9144);
nand U14681 (N_14681,N_8102,N_6752);
nor U14682 (N_14682,N_6695,N_7474);
or U14683 (N_14683,N_5789,N_8645);
and U14684 (N_14684,N_5304,N_9034);
or U14685 (N_14685,N_9305,N_5938);
and U14686 (N_14686,N_7215,N_8184);
nor U14687 (N_14687,N_6599,N_8092);
and U14688 (N_14688,N_5652,N_5890);
or U14689 (N_14689,N_9688,N_9891);
nor U14690 (N_14690,N_5994,N_8899);
nor U14691 (N_14691,N_8190,N_7968);
nand U14692 (N_14692,N_9667,N_6145);
nand U14693 (N_14693,N_8108,N_8454);
or U14694 (N_14694,N_6595,N_9590);
nand U14695 (N_14695,N_5522,N_6596);
or U14696 (N_14696,N_7172,N_6849);
nand U14697 (N_14697,N_9070,N_5211);
or U14698 (N_14698,N_9904,N_7972);
and U14699 (N_14699,N_8375,N_9503);
or U14700 (N_14700,N_5449,N_7511);
and U14701 (N_14701,N_5384,N_6877);
nand U14702 (N_14702,N_9702,N_5094);
nor U14703 (N_14703,N_7179,N_7440);
nor U14704 (N_14704,N_8683,N_5128);
nor U14705 (N_14705,N_6478,N_9677);
or U14706 (N_14706,N_9513,N_6870);
and U14707 (N_14707,N_9496,N_8400);
or U14708 (N_14708,N_7745,N_5265);
nand U14709 (N_14709,N_6410,N_6746);
nand U14710 (N_14710,N_6342,N_7844);
nor U14711 (N_14711,N_7613,N_8930);
nor U14712 (N_14712,N_5523,N_5913);
nor U14713 (N_14713,N_9836,N_6049);
nor U14714 (N_14714,N_6986,N_8875);
nand U14715 (N_14715,N_6358,N_5928);
and U14716 (N_14716,N_8794,N_6436);
and U14717 (N_14717,N_7788,N_6961);
nand U14718 (N_14718,N_5393,N_8335);
nor U14719 (N_14719,N_8584,N_8541);
nor U14720 (N_14720,N_9965,N_5217);
xnor U14721 (N_14721,N_6061,N_6086);
nand U14722 (N_14722,N_9141,N_6586);
and U14723 (N_14723,N_5404,N_6932);
nor U14724 (N_14724,N_9698,N_9169);
nor U14725 (N_14725,N_6328,N_5604);
nand U14726 (N_14726,N_8241,N_9093);
or U14727 (N_14727,N_5218,N_8982);
nand U14728 (N_14728,N_9662,N_7117);
or U14729 (N_14729,N_8671,N_6985);
or U14730 (N_14730,N_5634,N_8562);
nor U14731 (N_14731,N_6139,N_9228);
nor U14732 (N_14732,N_5373,N_5262);
or U14733 (N_14733,N_8517,N_6584);
or U14734 (N_14734,N_6294,N_9503);
nor U14735 (N_14735,N_7525,N_8721);
or U14736 (N_14736,N_6114,N_8495);
nand U14737 (N_14737,N_5576,N_5505);
and U14738 (N_14738,N_7725,N_9747);
and U14739 (N_14739,N_6318,N_8698);
or U14740 (N_14740,N_9764,N_8531);
nor U14741 (N_14741,N_6004,N_7805);
or U14742 (N_14742,N_6823,N_8745);
nand U14743 (N_14743,N_8355,N_7121);
or U14744 (N_14744,N_6978,N_6463);
or U14745 (N_14745,N_5577,N_9369);
or U14746 (N_14746,N_6941,N_8059);
or U14747 (N_14747,N_6298,N_6433);
nor U14748 (N_14748,N_9156,N_6221);
nor U14749 (N_14749,N_8357,N_8753);
or U14750 (N_14750,N_8423,N_9058);
nand U14751 (N_14751,N_6787,N_8922);
and U14752 (N_14752,N_7181,N_6765);
nor U14753 (N_14753,N_6776,N_6109);
nor U14754 (N_14754,N_7633,N_8341);
nor U14755 (N_14755,N_7716,N_8751);
nor U14756 (N_14756,N_6279,N_9641);
and U14757 (N_14757,N_8119,N_6650);
xor U14758 (N_14758,N_7016,N_8477);
nand U14759 (N_14759,N_5821,N_6421);
and U14760 (N_14760,N_5894,N_9824);
nand U14761 (N_14761,N_5408,N_7867);
and U14762 (N_14762,N_5252,N_5182);
or U14763 (N_14763,N_6580,N_5041);
nand U14764 (N_14764,N_5027,N_6385);
or U14765 (N_14765,N_8484,N_9724);
or U14766 (N_14766,N_5787,N_9367);
and U14767 (N_14767,N_5990,N_8281);
or U14768 (N_14768,N_5915,N_6488);
or U14769 (N_14769,N_8518,N_7642);
nand U14770 (N_14770,N_5977,N_7479);
xor U14771 (N_14771,N_9100,N_9396);
and U14772 (N_14772,N_5862,N_8451);
nand U14773 (N_14773,N_5453,N_9279);
nand U14774 (N_14774,N_7201,N_8823);
nor U14775 (N_14775,N_7905,N_6358);
and U14776 (N_14776,N_9132,N_8213);
nor U14777 (N_14777,N_8035,N_7015);
nand U14778 (N_14778,N_7099,N_9462);
nand U14779 (N_14779,N_5448,N_9065);
and U14780 (N_14780,N_9502,N_7489);
or U14781 (N_14781,N_6357,N_8809);
and U14782 (N_14782,N_6996,N_5923);
nor U14783 (N_14783,N_6925,N_7190);
or U14784 (N_14784,N_7892,N_8574);
or U14785 (N_14785,N_9235,N_9141);
nand U14786 (N_14786,N_6192,N_5032);
xnor U14787 (N_14787,N_6021,N_7177);
or U14788 (N_14788,N_8603,N_8380);
nor U14789 (N_14789,N_7197,N_6284);
or U14790 (N_14790,N_9650,N_5047);
or U14791 (N_14791,N_7328,N_6021);
nand U14792 (N_14792,N_6513,N_9199);
or U14793 (N_14793,N_7128,N_5251);
and U14794 (N_14794,N_6072,N_6164);
nor U14795 (N_14795,N_7589,N_5106);
nor U14796 (N_14796,N_7647,N_9715);
or U14797 (N_14797,N_9841,N_6348);
nand U14798 (N_14798,N_5420,N_7515);
nand U14799 (N_14799,N_9801,N_5548);
nand U14800 (N_14800,N_5142,N_9219);
and U14801 (N_14801,N_8661,N_6700);
and U14802 (N_14802,N_7863,N_9167);
and U14803 (N_14803,N_8429,N_5574);
and U14804 (N_14804,N_6837,N_5363);
nor U14805 (N_14805,N_5815,N_7174);
xor U14806 (N_14806,N_8362,N_7776);
nand U14807 (N_14807,N_5109,N_7843);
nand U14808 (N_14808,N_5456,N_9588);
or U14809 (N_14809,N_9170,N_5205);
nor U14810 (N_14810,N_5641,N_6203);
or U14811 (N_14811,N_6715,N_9181);
and U14812 (N_14812,N_5166,N_9856);
and U14813 (N_14813,N_5288,N_9868);
nand U14814 (N_14814,N_8359,N_9665);
or U14815 (N_14815,N_5894,N_7836);
and U14816 (N_14816,N_7180,N_8282);
nand U14817 (N_14817,N_7017,N_6261);
nand U14818 (N_14818,N_8430,N_8693);
or U14819 (N_14819,N_5192,N_7510);
and U14820 (N_14820,N_9963,N_8187);
or U14821 (N_14821,N_9746,N_8395);
nand U14822 (N_14822,N_9799,N_9427);
nor U14823 (N_14823,N_7409,N_9717);
nand U14824 (N_14824,N_8545,N_8998);
xnor U14825 (N_14825,N_6000,N_8713);
nor U14826 (N_14826,N_5589,N_8149);
nand U14827 (N_14827,N_5751,N_7239);
nand U14828 (N_14828,N_7336,N_9639);
nand U14829 (N_14829,N_9838,N_9739);
or U14830 (N_14830,N_5162,N_5009);
and U14831 (N_14831,N_8561,N_6129);
and U14832 (N_14832,N_5608,N_8573);
nor U14833 (N_14833,N_8621,N_7983);
nand U14834 (N_14834,N_6376,N_9813);
or U14835 (N_14835,N_6934,N_9652);
and U14836 (N_14836,N_6548,N_9371);
nor U14837 (N_14837,N_8002,N_9895);
nor U14838 (N_14838,N_6904,N_8236);
and U14839 (N_14839,N_5764,N_8425);
nand U14840 (N_14840,N_8446,N_5100);
or U14841 (N_14841,N_7151,N_8245);
nor U14842 (N_14842,N_5421,N_8243);
nor U14843 (N_14843,N_8044,N_8381);
nand U14844 (N_14844,N_9419,N_5643);
nand U14845 (N_14845,N_5026,N_9695);
nand U14846 (N_14846,N_7441,N_8425);
nand U14847 (N_14847,N_7365,N_6722);
nor U14848 (N_14848,N_8018,N_7889);
or U14849 (N_14849,N_6030,N_8746);
and U14850 (N_14850,N_9059,N_7501);
nand U14851 (N_14851,N_6053,N_5287);
nor U14852 (N_14852,N_8254,N_5696);
nor U14853 (N_14853,N_9644,N_7886);
or U14854 (N_14854,N_8022,N_5365);
nor U14855 (N_14855,N_9723,N_7377);
and U14856 (N_14856,N_9320,N_5619);
or U14857 (N_14857,N_7237,N_6687);
nand U14858 (N_14858,N_9787,N_9803);
and U14859 (N_14859,N_9312,N_5310);
nand U14860 (N_14860,N_6374,N_5066);
nor U14861 (N_14861,N_9650,N_5388);
nor U14862 (N_14862,N_7315,N_8192);
nand U14863 (N_14863,N_9086,N_6017);
or U14864 (N_14864,N_5093,N_5251);
xor U14865 (N_14865,N_9641,N_9057);
nor U14866 (N_14866,N_7150,N_9955);
or U14867 (N_14867,N_7606,N_7971);
or U14868 (N_14868,N_5069,N_9764);
or U14869 (N_14869,N_5673,N_8379);
nor U14870 (N_14870,N_8101,N_8452);
and U14871 (N_14871,N_5181,N_8600);
nand U14872 (N_14872,N_9005,N_9098);
and U14873 (N_14873,N_8381,N_7107);
or U14874 (N_14874,N_5766,N_8834);
nand U14875 (N_14875,N_9242,N_8443);
nand U14876 (N_14876,N_8672,N_8613);
and U14877 (N_14877,N_5154,N_8970);
nand U14878 (N_14878,N_7258,N_9137);
or U14879 (N_14879,N_5357,N_5016);
and U14880 (N_14880,N_7358,N_6762);
or U14881 (N_14881,N_5444,N_7743);
nor U14882 (N_14882,N_9363,N_9203);
nor U14883 (N_14883,N_8017,N_7961);
and U14884 (N_14884,N_5455,N_5793);
xnor U14885 (N_14885,N_5076,N_9388);
or U14886 (N_14886,N_9590,N_6155);
nor U14887 (N_14887,N_5401,N_6991);
and U14888 (N_14888,N_6548,N_8742);
nand U14889 (N_14889,N_9557,N_8717);
nand U14890 (N_14890,N_6388,N_9236);
nand U14891 (N_14891,N_9737,N_7481);
or U14892 (N_14892,N_9512,N_8409);
nand U14893 (N_14893,N_8183,N_5388);
nand U14894 (N_14894,N_7829,N_6792);
nand U14895 (N_14895,N_8088,N_5872);
nor U14896 (N_14896,N_9664,N_9892);
and U14897 (N_14897,N_7180,N_8612);
or U14898 (N_14898,N_5807,N_5668);
and U14899 (N_14899,N_9989,N_9650);
and U14900 (N_14900,N_5546,N_5324);
and U14901 (N_14901,N_9622,N_5177);
nand U14902 (N_14902,N_5567,N_6748);
nand U14903 (N_14903,N_7211,N_8781);
or U14904 (N_14904,N_8433,N_6702);
nand U14905 (N_14905,N_6691,N_5874);
nand U14906 (N_14906,N_7066,N_8282);
nand U14907 (N_14907,N_6506,N_8532);
nor U14908 (N_14908,N_5260,N_6582);
nor U14909 (N_14909,N_8427,N_5747);
and U14910 (N_14910,N_7203,N_9128);
and U14911 (N_14911,N_5365,N_5128);
nand U14912 (N_14912,N_7172,N_5788);
or U14913 (N_14913,N_5719,N_9393);
and U14914 (N_14914,N_6836,N_8528);
and U14915 (N_14915,N_8980,N_6408);
or U14916 (N_14916,N_9410,N_7295);
nor U14917 (N_14917,N_7851,N_7338);
or U14918 (N_14918,N_9010,N_9734);
nor U14919 (N_14919,N_7298,N_9165);
nand U14920 (N_14920,N_5774,N_7851);
nand U14921 (N_14921,N_8398,N_9911);
and U14922 (N_14922,N_6239,N_8745);
nand U14923 (N_14923,N_7479,N_9288);
and U14924 (N_14924,N_9478,N_7607);
or U14925 (N_14925,N_8237,N_9109);
or U14926 (N_14926,N_9554,N_9880);
nor U14927 (N_14927,N_7942,N_8427);
or U14928 (N_14928,N_5951,N_7766);
nand U14929 (N_14929,N_9166,N_5988);
or U14930 (N_14930,N_5886,N_7559);
and U14931 (N_14931,N_6962,N_7899);
or U14932 (N_14932,N_5045,N_8831);
nand U14933 (N_14933,N_9042,N_9669);
and U14934 (N_14934,N_5086,N_9991);
and U14935 (N_14935,N_6507,N_9017);
xnor U14936 (N_14936,N_8810,N_9283);
xor U14937 (N_14937,N_7843,N_9748);
and U14938 (N_14938,N_8139,N_5949);
and U14939 (N_14939,N_9168,N_8308);
nand U14940 (N_14940,N_6918,N_7354);
nand U14941 (N_14941,N_6792,N_9056);
or U14942 (N_14942,N_6171,N_9097);
and U14943 (N_14943,N_8739,N_8792);
nor U14944 (N_14944,N_8243,N_5154);
nor U14945 (N_14945,N_5818,N_7375);
or U14946 (N_14946,N_9140,N_5414);
and U14947 (N_14947,N_6444,N_6021);
or U14948 (N_14948,N_7155,N_5904);
nand U14949 (N_14949,N_8761,N_8013);
or U14950 (N_14950,N_7205,N_5449);
or U14951 (N_14951,N_6577,N_6166);
and U14952 (N_14952,N_6494,N_8512);
nor U14953 (N_14953,N_6010,N_8169);
nand U14954 (N_14954,N_7347,N_7276);
nand U14955 (N_14955,N_6610,N_7954);
or U14956 (N_14956,N_8127,N_6957);
and U14957 (N_14957,N_8950,N_5499);
or U14958 (N_14958,N_5813,N_5489);
or U14959 (N_14959,N_7656,N_5297);
or U14960 (N_14960,N_8099,N_9564);
or U14961 (N_14961,N_9411,N_9834);
nor U14962 (N_14962,N_9436,N_7880);
or U14963 (N_14963,N_7779,N_9227);
nor U14964 (N_14964,N_7735,N_5373);
and U14965 (N_14965,N_8947,N_7812);
and U14966 (N_14966,N_8073,N_7979);
and U14967 (N_14967,N_6756,N_9378);
and U14968 (N_14968,N_8959,N_5605);
and U14969 (N_14969,N_9343,N_9044);
or U14970 (N_14970,N_9740,N_8321);
or U14971 (N_14971,N_8828,N_7253);
or U14972 (N_14972,N_6255,N_7850);
nand U14973 (N_14973,N_7436,N_6604);
or U14974 (N_14974,N_6341,N_6590);
nand U14975 (N_14975,N_7249,N_8816);
and U14976 (N_14976,N_6347,N_7584);
and U14977 (N_14977,N_9290,N_6683);
nor U14978 (N_14978,N_9944,N_5609);
and U14979 (N_14979,N_7703,N_5972);
and U14980 (N_14980,N_8710,N_7946);
nor U14981 (N_14981,N_8808,N_7346);
nor U14982 (N_14982,N_7004,N_5344);
nor U14983 (N_14983,N_5541,N_5413);
nor U14984 (N_14984,N_8832,N_9782);
and U14985 (N_14985,N_7249,N_6649);
or U14986 (N_14986,N_8456,N_5804);
and U14987 (N_14987,N_7132,N_5465);
nor U14988 (N_14988,N_6874,N_6160);
nand U14989 (N_14989,N_7748,N_7946);
nand U14990 (N_14990,N_6091,N_7395);
or U14991 (N_14991,N_8974,N_5383);
nand U14992 (N_14992,N_8876,N_7256);
and U14993 (N_14993,N_9113,N_9600);
and U14994 (N_14994,N_9521,N_6303);
nor U14995 (N_14995,N_5867,N_9653);
nor U14996 (N_14996,N_5805,N_8570);
or U14997 (N_14997,N_7156,N_9239);
or U14998 (N_14998,N_6010,N_9255);
nor U14999 (N_14999,N_6265,N_8807);
or U15000 (N_15000,N_13270,N_14881);
and U15001 (N_15001,N_14826,N_10499);
nand U15002 (N_15002,N_11247,N_13142);
nand U15003 (N_15003,N_10675,N_11441);
or U15004 (N_15004,N_13569,N_11464);
nand U15005 (N_15005,N_14827,N_12158);
or U15006 (N_15006,N_13799,N_14584);
nor U15007 (N_15007,N_10546,N_12503);
nor U15008 (N_15008,N_11035,N_14149);
or U15009 (N_15009,N_14099,N_12057);
xnor U15010 (N_15010,N_12001,N_10103);
and U15011 (N_15011,N_12334,N_14474);
and U15012 (N_15012,N_13004,N_11877);
nand U15013 (N_15013,N_13212,N_12263);
or U15014 (N_15014,N_14284,N_10899);
nand U15015 (N_15015,N_12656,N_12816);
xnor U15016 (N_15016,N_12989,N_12366);
or U15017 (N_15017,N_12330,N_10667);
nor U15018 (N_15018,N_11760,N_12443);
nor U15019 (N_15019,N_14407,N_11514);
and U15020 (N_15020,N_10849,N_10114);
or U15021 (N_15021,N_12280,N_10775);
xnor U15022 (N_15022,N_10673,N_11936);
or U15023 (N_15023,N_10721,N_10293);
and U15024 (N_15024,N_12702,N_14890);
nand U15025 (N_15025,N_12274,N_10023);
nor U15026 (N_15026,N_13181,N_10662);
nor U15027 (N_15027,N_14063,N_12099);
nand U15028 (N_15028,N_12639,N_12568);
nor U15029 (N_15029,N_10030,N_12710);
or U15030 (N_15030,N_10129,N_14281);
or U15031 (N_15031,N_12582,N_11787);
nand U15032 (N_15032,N_11724,N_11453);
and U15033 (N_15033,N_11994,N_10746);
or U15034 (N_15034,N_13176,N_10484);
and U15035 (N_15035,N_14590,N_10349);
and U15036 (N_15036,N_13217,N_13797);
and U15037 (N_15037,N_14379,N_11072);
nor U15038 (N_15038,N_13612,N_13990);
or U15039 (N_15039,N_10783,N_13829);
or U15040 (N_15040,N_13676,N_10929);
or U15041 (N_15041,N_13005,N_14905);
nor U15042 (N_15042,N_11479,N_10630);
nand U15043 (N_15043,N_11949,N_13620);
nor U15044 (N_15044,N_10043,N_10756);
or U15045 (N_15045,N_11937,N_14080);
or U15046 (N_15046,N_11717,N_11652);
nor U15047 (N_15047,N_12472,N_14835);
nand U15048 (N_15048,N_10250,N_10087);
or U15049 (N_15049,N_13947,N_13890);
nor U15050 (N_15050,N_14822,N_14988);
and U15051 (N_15051,N_14721,N_13543);
xor U15052 (N_15052,N_13635,N_14567);
or U15053 (N_15053,N_14122,N_14177);
or U15054 (N_15054,N_13009,N_12002);
nand U15055 (N_15055,N_11752,N_10223);
or U15056 (N_15056,N_10866,N_14675);
nor U15057 (N_15057,N_10239,N_10346);
nor U15058 (N_15058,N_13559,N_11424);
or U15059 (N_15059,N_13775,N_11201);
and U15060 (N_15060,N_13608,N_14006);
or U15061 (N_15061,N_14949,N_11270);
or U15062 (N_15062,N_11747,N_10342);
and U15063 (N_15063,N_10928,N_10823);
and U15064 (N_15064,N_10649,N_10230);
nand U15065 (N_15065,N_12809,N_10222);
nor U15066 (N_15066,N_11767,N_11709);
nor U15067 (N_15067,N_14823,N_13241);
nand U15068 (N_15068,N_11641,N_11449);
nand U15069 (N_15069,N_14764,N_10504);
nor U15070 (N_15070,N_10085,N_10862);
nor U15071 (N_15071,N_10276,N_13630);
nor U15072 (N_15072,N_12772,N_11252);
and U15073 (N_15073,N_11896,N_13452);
nand U15074 (N_15074,N_13399,N_11154);
or U15075 (N_15075,N_10002,N_11625);
nand U15076 (N_15076,N_12345,N_10179);
and U15077 (N_15077,N_10073,N_12662);
nor U15078 (N_15078,N_12798,N_11714);
nor U15079 (N_15079,N_12153,N_10054);
and U15080 (N_15080,N_13474,N_11599);
or U15081 (N_15081,N_14683,N_11999);
and U15082 (N_15082,N_14261,N_12103);
or U15083 (N_15083,N_11681,N_12755);
nand U15084 (N_15084,N_13285,N_13973);
xnor U15085 (N_15085,N_11582,N_13624);
nand U15086 (N_15086,N_12234,N_14419);
nand U15087 (N_15087,N_14652,N_11845);
and U15088 (N_15088,N_14832,N_12232);
and U15089 (N_15089,N_14493,N_10229);
nor U15090 (N_15090,N_11023,N_11055);
and U15091 (N_15091,N_13373,N_10505);
xnor U15092 (N_15092,N_13727,N_10781);
and U15093 (N_15093,N_13506,N_14674);
or U15094 (N_15094,N_13333,N_14280);
or U15095 (N_15095,N_13747,N_14694);
or U15096 (N_15096,N_12365,N_14211);
and U15097 (N_15097,N_14882,N_12940);
nand U15098 (N_15098,N_10955,N_10100);
xor U15099 (N_15099,N_13991,N_12194);
and U15100 (N_15100,N_14530,N_13589);
or U15101 (N_15101,N_11535,N_14834);
or U15102 (N_15102,N_13438,N_12546);
or U15103 (N_15103,N_13495,N_10827);
nand U15104 (N_15104,N_10989,N_14982);
and U15105 (N_15105,N_14361,N_13822);
and U15106 (N_15106,N_13546,N_10444);
xnor U15107 (N_15107,N_13049,N_14370);
nand U15108 (N_15108,N_14517,N_14927);
or U15109 (N_15109,N_11618,N_10931);
nand U15110 (N_15110,N_11614,N_11073);
and U15111 (N_15111,N_14179,N_10733);
or U15112 (N_15112,N_10914,N_14442);
nor U15113 (N_15113,N_10300,N_10120);
nor U15114 (N_15114,N_12214,N_12992);
nor U15115 (N_15115,N_14874,N_10324);
or U15116 (N_15116,N_10824,N_13713);
and U15117 (N_15117,N_10701,N_14819);
nor U15118 (N_15118,N_10258,N_12984);
and U15119 (N_15119,N_11084,N_11696);
nand U15120 (N_15120,N_13062,N_12819);
nor U15121 (N_15121,N_12937,N_10060);
nor U15122 (N_15122,N_14998,N_11866);
or U15123 (N_15123,N_11263,N_10090);
or U15124 (N_15124,N_14718,N_13187);
and U15125 (N_15125,N_14167,N_12128);
nor U15126 (N_15126,N_13419,N_13283);
and U15127 (N_15127,N_14333,N_14313);
nor U15128 (N_15128,N_10228,N_10478);
nor U15129 (N_15129,N_12053,N_12492);
and U15130 (N_15130,N_12590,N_14685);
or U15131 (N_15131,N_11174,N_11202);
or U15132 (N_15132,N_12850,N_10902);
or U15133 (N_15133,N_10048,N_10555);
nand U15134 (N_15134,N_10353,N_10210);
nor U15135 (N_15135,N_12668,N_10692);
nand U15136 (N_15136,N_13792,N_14628);
and U15137 (N_15137,N_11275,N_14308);
or U15138 (N_15138,N_11329,N_11735);
nor U15139 (N_15139,N_10600,N_11519);
or U15140 (N_15140,N_14772,N_14305);
nor U15141 (N_15141,N_13463,N_14319);
and U15142 (N_15142,N_11269,N_11826);
and U15143 (N_15143,N_10777,N_14172);
nand U15144 (N_15144,N_13099,N_14836);
nand U15145 (N_15145,N_14723,N_11907);
nor U15146 (N_15146,N_14369,N_11506);
or U15147 (N_15147,N_10643,N_11150);
nor U15148 (N_15148,N_13958,N_12652);
nand U15149 (N_15149,N_13090,N_11560);
or U15150 (N_15150,N_10331,N_11611);
xnor U15151 (N_15151,N_11344,N_13366);
and U15152 (N_15152,N_12766,N_12764);
and U15153 (N_15153,N_12824,N_12270);
and U15154 (N_15154,N_12588,N_14456);
nor U15155 (N_15155,N_11967,N_14698);
nand U15156 (N_15156,N_13725,N_11588);
and U15157 (N_15157,N_13097,N_10415);
nand U15158 (N_15158,N_11232,N_12319);
or U15159 (N_15159,N_10235,N_14366);
and U15160 (N_15160,N_10072,N_14316);
or U15161 (N_15161,N_10295,N_11547);
and U15162 (N_15162,N_10808,N_11692);
and U15163 (N_15163,N_12032,N_11358);
nor U15164 (N_15164,N_14409,N_12219);
nand U15165 (N_15165,N_10475,N_10007);
nor U15166 (N_15166,N_12462,N_11635);
or U15167 (N_15167,N_10336,N_14522);
nor U15168 (N_15168,N_10465,N_12241);
or U15169 (N_15169,N_12341,N_12320);
and U15170 (N_15170,N_11149,N_10493);
or U15171 (N_15171,N_11012,N_12416);
or U15172 (N_15172,N_11989,N_12348);
nor U15173 (N_15173,N_10307,N_10032);
or U15174 (N_15174,N_14354,N_10556);
or U15175 (N_15175,N_14964,N_10565);
or U15176 (N_15176,N_11185,N_11505);
nand U15177 (N_15177,N_13834,N_10811);
nor U15178 (N_15178,N_13383,N_13138);
or U15179 (N_15179,N_13813,N_14645);
nor U15180 (N_15180,N_14662,N_12985);
and U15181 (N_15181,N_11995,N_10940);
and U15182 (N_15182,N_12564,N_12011);
or U15183 (N_15183,N_10577,N_11299);
or U15184 (N_15184,N_11902,N_12790);
nand U15185 (N_15185,N_10375,N_12557);
or U15186 (N_15186,N_12466,N_12998);
nand U15187 (N_15187,N_14575,N_12297);
or U15188 (N_15188,N_13454,N_12851);
or U15189 (N_15189,N_12253,N_10448);
nand U15190 (N_15190,N_10896,N_13444);
or U15191 (N_15191,N_13531,N_14779);
nand U15192 (N_15192,N_12629,N_14117);
nor U15193 (N_15193,N_11191,N_10852);
nor U15194 (N_15194,N_14376,N_10078);
and U15195 (N_15195,N_14735,N_12507);
nand U15196 (N_15196,N_11969,N_14966);
nor U15197 (N_15197,N_12430,N_11074);
nand U15198 (N_15198,N_11488,N_10839);
nor U15199 (N_15199,N_11975,N_14148);
nor U15200 (N_15200,N_10009,N_14594);
or U15201 (N_15201,N_10999,N_13875);
and U15202 (N_15202,N_11003,N_14412);
nor U15203 (N_15203,N_13206,N_11444);
nor U15204 (N_15204,N_11345,N_10867);
or U15205 (N_15205,N_11805,N_10338);
and U15206 (N_15206,N_11306,N_12182);
or U15207 (N_15207,N_12007,N_11122);
nand U15208 (N_15208,N_14453,N_11603);
or U15209 (N_15209,N_14020,N_11671);
nand U15210 (N_15210,N_12885,N_10483);
or U15211 (N_15211,N_13820,N_14644);
nor U15212 (N_15212,N_14765,N_13293);
xnor U15213 (N_15213,N_14842,N_13261);
or U15214 (N_15214,N_11629,N_11677);
or U15215 (N_15215,N_14037,N_13302);
nor U15216 (N_15216,N_12116,N_14174);
or U15217 (N_15217,N_11871,N_13355);
nor U15218 (N_15218,N_12963,N_13769);
or U15219 (N_15219,N_10587,N_14784);
xor U15220 (N_15220,N_12168,N_14257);
or U15221 (N_15221,N_10670,N_11952);
nor U15222 (N_15222,N_12536,N_14904);
nand U15223 (N_15223,N_11828,N_12831);
or U15224 (N_15224,N_10534,N_13215);
and U15225 (N_15225,N_11861,N_12948);
nor U15226 (N_15226,N_12283,N_12360);
xnor U15227 (N_15227,N_10298,N_13571);
and U15228 (N_15228,N_14898,N_11503);
or U15229 (N_15229,N_14670,N_12373);
or U15230 (N_15230,N_11580,N_11756);
or U15231 (N_15231,N_11156,N_13673);
nand U15232 (N_15232,N_10599,N_12339);
and U15233 (N_15233,N_12034,N_14506);
or U15234 (N_15234,N_14877,N_12954);
or U15235 (N_15235,N_10650,N_10612);
nor U15236 (N_15236,N_10743,N_10528);
or U15237 (N_15237,N_12732,N_11412);
and U15238 (N_15238,N_12523,N_13165);
xnor U15239 (N_15239,N_14999,N_13230);
nand U15240 (N_15240,N_12577,N_13318);
nor U15241 (N_15241,N_11274,N_12526);
and U15242 (N_15242,N_11928,N_12311);
nand U15243 (N_15243,N_14263,N_13823);
nor U15244 (N_15244,N_13964,N_12769);
and U15245 (N_15245,N_10387,N_14353);
and U15246 (N_15246,N_12121,N_12245);
or U15247 (N_15247,N_13002,N_12782);
nor U15248 (N_15248,N_12257,N_10784);
nor U15249 (N_15249,N_10189,N_13024);
nand U15250 (N_15250,N_14009,N_14061);
nor U15251 (N_15251,N_12248,N_10097);
or U15252 (N_15252,N_10402,N_11623);
nand U15253 (N_15253,N_13519,N_10146);
nand U15254 (N_15254,N_13115,N_12711);
and U15255 (N_15255,N_10330,N_10765);
or U15256 (N_15256,N_14925,N_14331);
nand U15257 (N_15257,N_10998,N_13362);
and U15258 (N_15258,N_13781,N_11892);
or U15259 (N_15259,N_14088,N_14038);
nor U15260 (N_15260,N_13104,N_10204);
nor U15261 (N_15261,N_13856,N_11331);
nor U15262 (N_15262,N_13103,N_13788);
xnor U15263 (N_15263,N_12335,N_11076);
nor U15264 (N_15264,N_12862,N_12695);
nor U15265 (N_15265,N_14075,N_10497);
nor U15266 (N_15266,N_14697,N_12789);
and U15267 (N_15267,N_13077,N_14385);
nand U15268 (N_15268,N_10814,N_11884);
and U15269 (N_15269,N_11373,N_12859);
nor U15270 (N_15270,N_10156,N_14555);
and U15271 (N_15271,N_13640,N_14098);
nand U15272 (N_15272,N_12820,N_14023);
or U15273 (N_15273,N_13521,N_14813);
xnor U15274 (N_15274,N_12213,N_14427);
and U15275 (N_15275,N_13852,N_13730);
and U15276 (N_15276,N_12312,N_14660);
or U15277 (N_15277,N_12870,N_13381);
nor U15278 (N_15278,N_14907,N_14921);
nor U15279 (N_15279,N_14750,N_12972);
or U15280 (N_15280,N_13391,N_10615);
nor U15281 (N_15281,N_10794,N_14479);
nor U15282 (N_15282,N_14841,N_10244);
and U15283 (N_15283,N_12803,N_11184);
nand U15284 (N_15284,N_12450,N_14028);
and U15285 (N_15285,N_12298,N_14649);
and U15286 (N_15286,N_10291,N_14951);
or U15287 (N_15287,N_14279,N_14895);
and U15288 (N_15288,N_13407,N_12900);
nor U15289 (N_15289,N_10385,N_10598);
and U15290 (N_15290,N_10644,N_10821);
and U15291 (N_15291,N_14844,N_10076);
and U15292 (N_15292,N_12968,N_14658);
and U15293 (N_15293,N_11883,N_11389);
nand U15294 (N_15294,N_13374,N_11546);
and U15295 (N_15295,N_10135,N_13083);
nor U15296 (N_15296,N_13485,N_11660);
or U15297 (N_15297,N_13325,N_12559);
nor U15298 (N_15298,N_10683,N_12691);
or U15299 (N_15299,N_12544,N_10725);
nor U15300 (N_15300,N_11241,N_14896);
or U15301 (N_15301,N_13209,N_13866);
or U15302 (N_15302,N_11935,N_12272);
nor U15303 (N_15303,N_13084,N_13455);
or U15304 (N_15304,N_14854,N_14993);
or U15305 (N_15305,N_13654,N_10618);
nor U15306 (N_15306,N_10218,N_13551);
nand U15307 (N_15307,N_10150,N_13584);
nor U15308 (N_15308,N_12428,N_14202);
nor U15309 (N_15309,N_14234,N_14940);
and U15310 (N_15310,N_13553,N_11164);
nor U15311 (N_15311,N_13647,N_11810);
or U15312 (N_15312,N_13783,N_14414);
and U15313 (N_15313,N_14351,N_13561);
and U15314 (N_15314,N_14397,N_13617);
or U15315 (N_15315,N_13033,N_11339);
or U15316 (N_15316,N_14087,N_10106);
nand U15317 (N_15317,N_14496,N_13233);
or U15318 (N_15318,N_13168,N_11846);
or U15319 (N_15319,N_14243,N_13914);
and U15320 (N_15320,N_12922,N_13441);
nand U15321 (N_15321,N_11411,N_13698);
xnor U15322 (N_15322,N_10786,N_11207);
or U15323 (N_15323,N_11210,N_14304);
nand U15324 (N_15324,N_14445,N_12394);
nor U15325 (N_15325,N_10715,N_14745);
nand U15326 (N_15326,N_11564,N_14036);
and U15327 (N_15327,N_10270,N_13023);
and U15328 (N_15328,N_14143,N_13190);
and U15329 (N_15329,N_10578,N_14792);
and U15330 (N_15330,N_14299,N_12268);
nor U15331 (N_15331,N_11923,N_14503);
nor U15332 (N_15332,N_12132,N_13322);
or U15333 (N_15333,N_14300,N_10638);
or U15334 (N_15334,N_13742,N_12452);
or U15335 (N_15335,N_10158,N_13805);
or U15336 (N_15336,N_13061,N_11777);
nor U15337 (N_15337,N_11098,N_11437);
xor U15338 (N_15338,N_12150,N_13672);
and U15339 (N_15339,N_11260,N_10884);
nand U15340 (N_15340,N_12172,N_12663);
nor U15341 (N_15341,N_11356,N_10635);
nor U15342 (N_15342,N_11755,N_12643);
nor U15343 (N_15343,N_13078,N_12187);
nor U15344 (N_15344,N_12949,N_13824);
or U15345 (N_15345,N_11286,N_13919);
or U15346 (N_15346,N_11016,N_11139);
nor U15347 (N_15347,N_13012,N_12793);
and U15348 (N_15348,N_13582,N_11398);
nor U15349 (N_15349,N_13307,N_14114);
nand U15350 (N_15350,N_10732,N_10904);
nor U15351 (N_15351,N_10315,N_12550);
or U15352 (N_15352,N_14116,N_10303);
or U15353 (N_15353,N_14611,N_13179);
nor U15354 (N_15354,N_14879,N_13595);
or U15355 (N_15355,N_10944,N_10540);
or U15356 (N_15356,N_10905,N_13927);
nor U15357 (N_15357,N_14521,N_10506);
and U15358 (N_15358,N_13039,N_14980);
nand U15359 (N_15359,N_12068,N_12482);
and U15360 (N_15360,N_12477,N_12898);
nand U15361 (N_15361,N_13798,N_11292);
nand U15362 (N_15362,N_12388,N_12863);
nand U15363 (N_15363,N_11462,N_11920);
and U15364 (N_15364,N_12332,N_12101);
nand U15365 (N_15365,N_11248,N_12200);
nand U15366 (N_15366,N_14971,N_13043);
and U15367 (N_15367,N_11416,N_14430);
nand U15368 (N_15368,N_12742,N_10409);
nand U15369 (N_15369,N_13281,N_14307);
nand U15370 (N_15370,N_10614,N_13906);
or U15371 (N_15371,N_13476,N_10249);
and U15372 (N_15372,N_11392,N_10633);
or U15373 (N_15373,N_13720,N_10580);
or U15374 (N_15374,N_12402,N_14719);
or U15375 (N_15375,N_13884,N_11972);
nor U15376 (N_15376,N_11667,N_14560);
nor U15377 (N_15377,N_11812,N_11419);
nand U15378 (N_15378,N_11743,N_10401);
or U15379 (N_15379,N_14511,N_14773);
nand U15380 (N_15380,N_10406,N_14033);
nand U15381 (N_15381,N_12299,N_13022);
nand U15382 (N_15382,N_13472,N_14274);
nand U15383 (N_15383,N_14540,N_13468);
and U15384 (N_15384,N_12369,N_10780);
and U15385 (N_15385,N_14145,N_10464);
nor U15386 (N_15386,N_14065,N_12527);
nor U15387 (N_15387,N_10525,N_13386);
and U15388 (N_15388,N_14965,N_12528);
nor U15389 (N_15389,N_10545,N_11357);
and U15390 (N_15390,N_10379,N_13003);
nand U15391 (N_15391,N_12750,N_14935);
nor U15392 (N_15392,N_12006,N_14686);
nor U15393 (N_15393,N_10136,N_10201);
nor U15394 (N_15394,N_13889,N_14968);
nor U15395 (N_15395,N_12911,N_10742);
nand U15396 (N_15396,N_12833,N_13710);
nand U15397 (N_15397,N_13464,N_13702);
nand U15398 (N_15398,N_12860,N_11842);
nor U15399 (N_15399,N_14207,N_11221);
nor U15400 (N_15400,N_13649,N_14358);
or U15401 (N_15401,N_11063,N_10672);
or U15402 (N_15402,N_14589,N_13684);
nand U15403 (N_15403,N_12094,N_13185);
nand U15404 (N_15404,N_10301,N_10166);
and U15405 (N_15405,N_12042,N_14219);
nor U15406 (N_15406,N_12329,N_11595);
and U15407 (N_15407,N_12930,N_13421);
nand U15408 (N_15408,N_14737,N_12399);
or U15409 (N_15409,N_14922,N_11565);
nand U15410 (N_15410,N_13743,N_10686);
and U15411 (N_15411,N_14679,N_12454);
nor U15412 (N_15412,N_13156,N_14947);
or U15413 (N_15413,N_13063,N_12328);
nor U15414 (N_15414,N_12469,N_11837);
or U15415 (N_15415,N_14634,N_11388);
xnor U15416 (N_15416,N_10011,N_10946);
and U15417 (N_15417,N_12131,N_13916);
or U15418 (N_15418,N_10278,N_13113);
nand U15419 (N_15419,N_14198,N_11266);
nor U15420 (N_15420,N_13069,N_13051);
nand U15421 (N_15421,N_11848,N_14630);
nand U15422 (N_15422,N_10413,N_14062);
or U15423 (N_15423,N_10547,N_10831);
and U15424 (N_15424,N_14421,N_10885);
nand U15425 (N_15425,N_12017,N_11673);
nand U15426 (N_15426,N_14956,N_14661);
nor U15427 (N_15427,N_12134,N_11739);
nor U15428 (N_15428,N_13790,N_13054);
or U15429 (N_15429,N_13403,N_11308);
nand U15430 (N_15430,N_12220,N_10225);
and U15431 (N_15431,N_11507,N_14785);
nand U15432 (N_15432,N_14051,N_10137);
and U15433 (N_15433,N_13456,N_14408);
or U15434 (N_15434,N_10010,N_12161);
nand U15435 (N_15435,N_11662,N_14746);
or U15436 (N_15436,N_10704,N_13257);
or U15437 (N_15437,N_10802,N_14963);
or U15438 (N_15438,N_11079,N_14296);
nor U15439 (N_15439,N_10981,N_14460);
and U15440 (N_15440,N_12731,N_11407);
and U15441 (N_15441,N_12987,N_11452);
and U15442 (N_15442,N_13922,N_11367);
or U15443 (N_15443,N_11821,N_14306);
xnor U15444 (N_15444,N_12195,N_11425);
and U15445 (N_15445,N_10154,N_10826);
nand U15446 (N_15446,N_12359,N_10741);
nor U15447 (N_15447,N_12846,N_14636);
xor U15448 (N_15448,N_13894,N_11335);
nand U15449 (N_15449,N_10762,N_14342);
and U15450 (N_15450,N_11909,N_13818);
and U15451 (N_15451,N_12260,N_11046);
nand U15452 (N_15452,N_14060,N_13193);
or U15453 (N_15453,N_11744,N_12491);
xnor U15454 (N_15454,N_12144,N_12000);
or U15455 (N_15455,N_10817,N_13242);
and U15456 (N_15456,N_10344,N_13191);
and U15457 (N_15457,N_11733,N_12368);
nand U15458 (N_15458,N_12302,N_12918);
or U15459 (N_15459,N_12786,N_11151);
or U15460 (N_15460,N_10971,N_12840);
nand U15461 (N_15461,N_12129,N_10772);
nor U15462 (N_15462,N_11251,N_14431);
xnor U15463 (N_15463,N_11982,N_10829);
or U15464 (N_15464,N_12417,N_13714);
or U15465 (N_15465,N_14958,N_11362);
nor U15466 (N_15466,N_12688,N_11377);
nand U15467 (N_15467,N_12599,N_12928);
or U15468 (N_15468,N_14232,N_10750);
nor U15469 (N_15469,N_11713,N_14021);
nor U15470 (N_15470,N_12203,N_13317);
and U15471 (N_15471,N_13974,N_14146);
and U15472 (N_15472,N_14046,N_11486);
nand U15473 (N_15473,N_10651,N_13757);
nor U15474 (N_15474,N_14903,N_12612);
nor U15475 (N_15475,N_11058,N_14559);
and U15476 (N_15476,N_10142,N_13904);
nor U15477 (N_15477,N_11303,N_14564);
nand U15478 (N_15478,N_14251,N_10573);
and U15479 (N_15479,N_13669,N_10785);
nor U15480 (N_15480,N_12160,N_14349);
xor U15481 (N_15481,N_13276,N_12265);
nor U15482 (N_15482,N_11782,N_12465);
xnor U15483 (N_15483,N_11684,N_13855);
nor U15484 (N_15484,N_10511,N_12135);
or U15485 (N_15485,N_12828,N_11439);
nor U15486 (N_15486,N_14378,N_14108);
and U15487 (N_15487,N_13999,N_13245);
and U15488 (N_15488,N_10723,N_12779);
nor U15489 (N_15489,N_10436,N_12109);
and U15490 (N_15490,N_13717,N_10461);
or U15491 (N_15491,N_13550,N_11018);
or U15492 (N_15492,N_11715,N_10522);
nand U15493 (N_15493,N_14599,N_12690);
nand U15494 (N_15494,N_14533,N_10969);
or U15495 (N_15495,N_13659,N_13915);
nor U15496 (N_15496,N_11494,N_11267);
or U15497 (N_15497,N_13445,N_11770);
nor U15498 (N_15498,N_13228,N_10842);
or U15499 (N_15499,N_14216,N_14578);
and U15500 (N_15500,N_14700,N_13804);
nor U15501 (N_15501,N_12830,N_13045);
xnor U15502 (N_15502,N_11324,N_10018);
nand U15503 (N_15503,N_14977,N_11159);
nand U15504 (N_15504,N_14541,N_12364);
nor U15505 (N_15505,N_14213,N_12781);
or U15506 (N_15506,N_10729,N_14016);
nor U15507 (N_15507,N_13031,N_11215);
or U15508 (N_15508,N_14911,N_13197);
nor U15509 (N_15509,N_12300,N_13996);
nand U15510 (N_15510,N_11596,N_11761);
nor U15511 (N_15511,N_12857,N_14931);
nor U15512 (N_15512,N_12277,N_11737);
nor U15513 (N_15513,N_13372,N_14640);
or U15514 (N_15514,N_12249,N_10753);
nand U15515 (N_15515,N_10767,N_10488);
nand U15516 (N_15516,N_13933,N_13854);
or U15517 (N_15517,N_10485,N_12321);
nor U15518 (N_15518,N_13405,N_10537);
nor U15519 (N_15519,N_11663,N_11131);
nand U15520 (N_15520,N_10642,N_13101);
xnor U15521 (N_15521,N_13048,N_13838);
or U15522 (N_15522,N_13149,N_11493);
or U15523 (N_15523,N_12440,N_12719);
or U15524 (N_15524,N_11249,N_13954);
nand U15525 (N_15525,N_10093,N_14732);
nand U15526 (N_15526,N_11647,N_12515);
nor U15527 (N_15527,N_13515,N_13970);
nor U15528 (N_15528,N_10579,N_12692);
nor U15529 (N_15529,N_13268,N_14318);
or U15530 (N_15530,N_12347,N_14338);
nor U15531 (N_15531,N_11077,N_13496);
nand U15532 (N_15532,N_12539,N_10255);
or U15533 (N_15533,N_10807,N_14173);
and U15534 (N_15534,N_10611,N_13460);
or U15535 (N_15535,N_13483,N_12142);
nor U15536 (N_15536,N_14736,N_12282);
and U15537 (N_15537,N_11970,N_10372);
or U15538 (N_15538,N_10131,N_11466);
nand U15539 (N_15539,N_13392,N_11404);
and U15540 (N_15540,N_14180,N_14348);
and U15541 (N_15541,N_14267,N_10168);
nor U15542 (N_15542,N_14368,N_12835);
nand U15543 (N_15543,N_14542,N_14112);
nand U15544 (N_15544,N_12843,N_12060);
or U15545 (N_15545,N_10795,N_12625);
nor U15546 (N_15546,N_10719,N_12810);
or U15547 (N_15547,N_10538,N_10584);
and U15548 (N_15548,N_13255,N_10176);
nor U15549 (N_15549,N_13323,N_13642);
and U15550 (N_15550,N_14598,N_10134);
and U15551 (N_15551,N_11468,N_13414);
and U15552 (N_15552,N_12609,N_13437);
and U15553 (N_15553,N_10886,N_13231);
and U15554 (N_15554,N_12877,N_10031);
nand U15555 (N_15555,N_12585,N_13475);
and U15556 (N_15556,N_11984,N_14059);
or U15557 (N_15557,N_13663,N_12861);
nand U15558 (N_15558,N_11169,N_14056);
nor U15559 (N_15559,N_10963,N_10352);
and U15560 (N_15560,N_14195,N_13117);
xnor U15561 (N_15561,N_10216,N_10013);
or U15562 (N_15562,N_14298,N_14204);
nor U15563 (N_15563,N_12407,N_10727);
nand U15564 (N_15564,N_13633,N_11051);
nor U15565 (N_15565,N_14196,N_10015);
or U15566 (N_15566,N_14337,N_12083);
or U15567 (N_15567,N_13059,N_14265);
nor U15568 (N_15568,N_14415,N_10424);
nor U15569 (N_15569,N_12982,N_14380);
or U15570 (N_15570,N_11980,N_11708);
or U15571 (N_15571,N_10252,N_11602);
nor U15572 (N_15572,N_11173,N_12983);
or U15573 (N_15573,N_13573,N_14829);
or U15574 (N_15574,N_10924,N_10042);
nor U15575 (N_15575,N_14125,N_14272);
nand U15576 (N_15576,N_12421,N_12429);
or U15577 (N_15577,N_14711,N_10143);
and U15578 (N_15578,N_12881,N_13703);
nand U15579 (N_15579,N_12751,N_14734);
or U15580 (N_15580,N_13013,N_14585);
or U15581 (N_15581,N_10717,N_10959);
nand U15582 (N_15582,N_10200,N_13555);
nor U15583 (N_15583,N_13666,N_12709);
nand U15584 (N_15584,N_10922,N_10289);
nand U15585 (N_15585,N_11509,N_12962);
or U15586 (N_15586,N_13538,N_10119);
and U15587 (N_15587,N_11591,N_11351);
nor U15588 (N_15588,N_10046,N_11123);
nor U15589 (N_15589,N_10206,N_13542);
and U15590 (N_15590,N_14945,N_14483);
nor U15591 (N_15591,N_13446,N_12041);
or U15592 (N_15592,N_13849,N_12834);
nor U15593 (N_15593,N_13184,N_10040);
nand U15594 (N_15594,N_12837,N_12389);
or U15595 (N_15595,N_13956,N_12667);
or U15596 (N_15596,N_10068,N_14786);
nor U15597 (N_15597,N_13287,N_11117);
nand U15598 (N_15598,N_11219,N_11991);
nand U15599 (N_15599,N_14163,N_11350);
nor U15600 (N_15600,N_12054,N_10659);
or U15601 (N_15601,N_11375,N_10997);
nor U15602 (N_15602,N_10543,N_13699);
or U15603 (N_15603,N_10022,N_14768);
nor U15604 (N_15604,N_13670,N_14952);
nand U15605 (N_15605,N_12594,N_12196);
and U15606 (N_15606,N_10541,N_11898);
and U15607 (N_15607,N_14141,N_13164);
nand U15608 (N_15608,N_13199,N_11803);
or U15609 (N_15609,N_11617,N_13294);
or U15610 (N_15610,N_11410,N_11478);
nor U15611 (N_15611,N_10440,N_10132);
nand U15612 (N_15612,N_11730,N_13028);
and U15613 (N_15613,N_14848,N_13118);
xnor U15614 (N_15614,N_11878,N_10730);
nor U15615 (N_15615,N_12119,N_12414);
nand U15616 (N_15616,N_10369,N_12126);
nor U15617 (N_15617,N_14875,N_12938);
or U15618 (N_15618,N_11938,N_11523);
nand U15619 (N_15619,N_12566,N_11593);
nand U15620 (N_15620,N_11136,N_13136);
nand U15621 (N_15621,N_11198,N_14115);
nand U15622 (N_15622,N_13631,N_10995);
nand U15623 (N_15623,N_10897,N_14681);
nand U15624 (N_15624,N_13388,N_10476);
and U15625 (N_15625,N_11520,N_10943);
nor U15626 (N_15626,N_12510,N_11751);
or U15627 (N_15627,N_11799,N_13511);
nor U15628 (N_15628,N_12448,N_14513);
nand U15629 (N_15629,N_12075,N_12313);
or U15630 (N_15630,N_12541,N_12082);
nand U15631 (N_15631,N_13835,N_12303);
or U15632 (N_15632,N_13639,N_12326);
or U15633 (N_15633,N_14128,N_13667);
or U15634 (N_15634,N_14441,N_13015);
nand U15635 (N_15635,N_12642,N_13901);
or U15636 (N_15636,N_10297,N_12291);
nand U15637 (N_15637,N_14389,N_11155);
nand U15638 (N_15638,N_14902,N_14897);
nand U15639 (N_15639,N_12367,N_10061);
nand U15640 (N_15640,N_12897,N_10912);
and U15641 (N_15641,N_14843,N_13275);
or U15642 (N_15642,N_14224,N_14803);
and U15643 (N_15643,N_12896,N_12524);
and U15644 (N_15644,N_14808,N_10102);
nand U15645 (N_15645,N_12171,N_10954);
nor U15646 (N_15646,N_13772,N_10122);
and U15647 (N_15647,N_12490,N_14119);
or U15648 (N_15648,N_13607,N_14582);
and U15649 (N_15649,N_14226,N_11636);
nor U15650 (N_15650,N_14692,N_14969);
or U15651 (N_15651,N_14201,N_14672);
or U15652 (N_15652,N_10028,N_13917);
nor U15653 (N_15653,N_10152,N_13172);
and U15654 (N_15654,N_10130,N_13409);
nor U15655 (N_15655,N_14553,N_11047);
and U15656 (N_15656,N_11181,N_13272);
nor U15657 (N_15657,N_13298,N_13232);
nand U15658 (N_15658,N_11304,N_12179);
or U15659 (N_15659,N_12235,N_14825);
and U15660 (N_15660,N_11319,N_13134);
nor U15661 (N_15661,N_12980,N_14132);
nor U15662 (N_15662,N_10319,N_10075);
and U15663 (N_15663,N_10870,N_14713);
and U15664 (N_15664,N_14238,N_10872);
nand U15665 (N_15665,N_11321,N_12669);
nor U15666 (N_15666,N_10423,N_13535);
nand U15667 (N_15667,N_12164,N_13610);
nor U15668 (N_15668,N_11659,N_14001);
nand U15669 (N_15669,N_10550,N_14972);
and U15670 (N_15670,N_11836,N_10113);
nand U15671 (N_15671,N_12915,N_11534);
nand U15672 (N_15672,N_14150,N_12425);
nand U15673 (N_15673,N_12531,N_10447);
nand U15674 (N_15674,N_12178,N_11119);
or U15675 (N_15675,N_14991,N_11790);
or U15676 (N_15676,N_13660,N_14990);
and U15677 (N_15677,N_11276,N_13754);
nand U15678 (N_15678,N_11111,N_14816);
and U15679 (N_15679,N_13357,N_14228);
nand U15680 (N_15680,N_13425,N_10455);
nand U15681 (N_15681,N_11533,N_14806);
xnor U15682 (N_15682,N_13135,N_12137);
or U15683 (N_15683,N_14248,N_10706);
or U15684 (N_15684,N_12033,N_12728);
and U15685 (N_15685,N_11910,N_14069);
nor U15686 (N_15686,N_10676,N_13431);
and U15687 (N_15687,N_12139,N_14892);
or U15688 (N_15688,N_14151,N_14543);
nor U15689 (N_15689,N_12522,N_12701);
nor U15690 (N_15690,N_12969,N_14103);
or U15691 (N_15691,N_10036,N_12390);
and U15692 (N_15692,N_10835,N_11282);
nand U15693 (N_15693,N_10859,N_12216);
and U15694 (N_15694,N_12547,N_10863);
and U15695 (N_15695,N_10949,N_12943);
nand U15696 (N_15696,N_12090,N_14864);
or U15697 (N_15697,N_13141,N_14025);
nand U15698 (N_15698,N_11978,N_13082);
nand U15699 (N_15699,N_10329,N_13262);
nor U15700 (N_15700,N_14470,N_12650);
nor U15701 (N_15701,N_13385,N_11973);
and U15702 (N_15702,N_14347,N_14231);
nor U15703 (N_15703,N_13052,N_13885);
nor U15704 (N_15704,N_12617,N_10139);
and U15705 (N_15705,N_14791,N_12162);
or U15706 (N_15706,N_11697,N_13936);
and U15707 (N_15707,N_13413,N_14078);
nor U15708 (N_15708,N_10806,N_13677);
and U15709 (N_15709,N_14086,N_12210);
or U15710 (N_15710,N_14203,N_11903);
and U15711 (N_15711,N_10828,N_14083);
and U15712 (N_15712,N_13032,N_10281);
and U15713 (N_15713,N_11060,N_12147);
and U15714 (N_15714,N_12761,N_12767);
or U15715 (N_15715,N_11163,N_14710);
nand U15716 (N_15716,N_10232,N_14343);
or U15717 (N_15717,N_13057,N_11532);
and U15718 (N_15718,N_12892,N_14872);
or U15719 (N_15719,N_10482,N_11859);
nor U15720 (N_15720,N_13253,N_14755);
or U15721 (N_15721,N_13347,N_13095);
and U15722 (N_15722,N_10126,N_13335);
or U15723 (N_15723,N_12601,N_14603);
nand U15724 (N_15724,N_14096,N_12338);
nor U15725 (N_15725,N_13489,N_11583);
and U15726 (N_15726,N_12071,N_14356);
or U15727 (N_15727,N_14979,N_11758);
nor U15728 (N_15728,N_10764,N_11811);
nand U15729 (N_15729,N_11006,N_14863);
nor U15730 (N_15730,N_14341,N_10690);
or U15731 (N_15731,N_10231,N_10838);
and U15732 (N_15732,N_12349,N_13959);
nor U15733 (N_15733,N_14794,N_11882);
or U15734 (N_15734,N_10937,N_11839);
and U15735 (N_15735,N_14363,N_12799);
nor U15736 (N_15736,N_14627,N_12061);
nand U15737 (N_15737,N_12866,N_11062);
and U15738 (N_15738,N_10589,N_10208);
or U15739 (N_15739,N_11813,N_13926);
nand U15740 (N_15740,N_11102,N_10052);
nor U15741 (N_15741,N_12130,N_14187);
and U15742 (N_15742,N_12903,N_11827);
and U15743 (N_15743,N_13432,N_10321);
or U15744 (N_15744,N_10332,N_12730);
xnor U15745 (N_15745,N_13971,N_12494);
nor U15746 (N_15746,N_11855,N_11895);
nor U15747 (N_15747,N_11885,N_13564);
nor U15748 (N_15748,N_11033,N_14657);
nand U15749 (N_15749,N_10173,N_14539);
or U15750 (N_15750,N_14089,N_13349);
nand U15751 (N_15751,N_14311,N_12997);
nor U15752 (N_15752,N_13602,N_13290);
and U15753 (N_15753,N_11430,N_11075);
and U15754 (N_15754,N_11570,N_10008);
nand U15755 (N_15755,N_11958,N_13845);
or U15756 (N_15756,N_11471,N_12358);
nor U15757 (N_15757,N_11824,N_14568);
nor U15758 (N_15758,N_14748,N_11922);
nand U15759 (N_15759,N_12063,N_14067);
and U15760 (N_15760,N_10133,N_12114);
and U15761 (N_15761,N_10738,N_13932);
or U15762 (N_15762,N_14583,N_12288);
or U15763 (N_15763,N_10752,N_12384);
or U15764 (N_15764,N_12333,N_12540);
xnor U15765 (N_15765,N_11302,N_14486);
nand U15766 (N_15766,N_14229,N_11807);
or U15767 (N_15767,N_14252,N_12201);
nor U15768 (N_15768,N_12412,N_11986);
and U15769 (N_15769,N_12978,N_10323);
and U15770 (N_15770,N_10275,N_10711);
nand U15771 (N_15771,N_11977,N_13177);
nand U15772 (N_15772,N_11212,N_12226);
xnor U15773 (N_15773,N_14049,N_10820);
nand U15774 (N_15774,N_11701,N_10552);
or U15775 (N_15775,N_13998,N_13886);
nor U15776 (N_15776,N_13777,N_13731);
or U15777 (N_15777,N_11092,N_10069);
nor U15778 (N_15778,N_12961,N_13704);
nand U15779 (N_15779,N_13957,N_12956);
and U15780 (N_15780,N_10282,N_13946);
nor U15781 (N_15781,N_13071,N_13085);
nand U15782 (N_15782,N_10739,N_12655);
or U15783 (N_15783,N_12567,N_10350);
or U15784 (N_15784,N_13756,N_12474);
and U15785 (N_15785,N_11825,N_14741);
nand U15786 (N_15786,N_10196,N_11780);
or U15787 (N_15787,N_13778,N_11328);
and U15788 (N_15788,N_12573,N_11243);
or U15789 (N_15789,N_13017,N_11095);
and U15790 (N_15790,N_12794,N_13046);
or U15791 (N_15791,N_10463,N_10993);
or U15792 (N_15792,N_13119,N_10053);
or U15793 (N_15793,N_11172,N_13930);
or U15794 (N_15794,N_10262,N_14392);
and U15795 (N_15795,N_13701,N_13853);
nor U15796 (N_15796,N_12736,N_11965);
or U15797 (N_15797,N_12967,N_14635);
nor U15798 (N_15798,N_12832,N_14689);
nand U15799 (N_15799,N_11968,N_12953);
or U15800 (N_15800,N_14052,N_12058);
nand U15801 (N_15801,N_13811,N_12043);
xor U15802 (N_15802,N_13105,N_10443);
and U15803 (N_15803,N_13504,N_13091);
and U15804 (N_15804,N_14709,N_10192);
xor U15805 (N_15805,N_10473,N_14024);
nand U15806 (N_15806,N_10796,N_10530);
nand U15807 (N_15807,N_13214,N_12089);
nand U15808 (N_15808,N_14457,N_13128);
or U15809 (N_15809,N_10080,N_10045);
or U15810 (N_15810,N_12530,N_10390);
or U15811 (N_15811,N_10627,N_11455);
or U15812 (N_15812,N_14946,N_14375);
nand U15813 (N_15813,N_10425,N_11934);
and U15814 (N_15814,N_11021,N_10489);
nand U15815 (N_15815,N_12045,N_10868);
nand U15816 (N_15816,N_11687,N_11706);
or U15817 (N_15817,N_12648,N_14880);
nor U15818 (N_15818,N_14085,N_12314);
and U15819 (N_15819,N_14066,N_13221);
xor U15820 (N_15820,N_12152,N_10951);
nand U15821 (N_15821,N_13311,N_13398);
nor U15822 (N_15822,N_11094,N_10883);
nor U15823 (N_15823,N_10322,N_13401);
nor U15824 (N_15824,N_14840,N_14554);
nor U15825 (N_15825,N_12973,N_12059);
nand U15826 (N_15826,N_10172,N_13692);
or U15827 (N_15827,N_14162,N_11262);
and U15828 (N_15828,N_13375,N_14934);
and U15829 (N_15829,N_12015,N_11897);
or U15830 (N_15830,N_11763,N_12644);
nand U15831 (N_15831,N_12887,N_14950);
nand U15832 (N_15832,N_13442,N_13058);
nand U15833 (N_15833,N_10570,N_10893);
and U15834 (N_15834,N_14048,N_13766);
nand U15835 (N_15835,N_14104,N_11665);
nor U15836 (N_15836,N_14708,N_14899);
or U15837 (N_15837,N_10427,N_14753);
or U15838 (N_15838,N_14433,N_14619);
nand U15839 (N_15839,N_13139,N_11011);
or U15840 (N_15840,N_11571,N_13011);
nor U15841 (N_15841,N_10144,N_13434);
nand U15842 (N_15842,N_12247,N_13127);
nand U15843 (N_15843,N_11245,N_14482);
nand U15844 (N_15844,N_12087,N_13303);
nor U15845 (N_15845,N_10408,N_13600);
or U15846 (N_15846,N_13198,N_11932);
nand U15847 (N_15847,N_14962,N_11390);
and U15848 (N_15848,N_14550,N_13416);
nand U15849 (N_15849,N_11296,N_10634);
nand U15850 (N_15850,N_11985,N_13484);
nand U15851 (N_15851,N_13516,N_10822);
or U15852 (N_15852,N_14793,N_14695);
nor U15853 (N_15853,N_12561,N_10498);
nand U15854 (N_15854,N_12411,N_11472);
or U15855 (N_15855,N_10451,N_14406);
nor U15856 (N_15856,N_14362,N_13532);
and U15857 (N_15857,N_11291,N_13893);
and U15858 (N_15858,N_13661,N_14225);
nand U15859 (N_15859,N_11029,N_11820);
nand U15860 (N_15860,N_10891,N_14525);
nand U15861 (N_15861,N_13503,N_10325);
nand U15862 (N_15862,N_10492,N_12250);
nor U15863 (N_15863,N_13334,N_14617);
nand U15864 (N_15864,N_10259,N_11010);
and U15865 (N_15865,N_14396,N_14161);
and U15866 (N_15866,N_10089,N_13847);
nand U15867 (N_15867,N_11707,N_12067);
and U15868 (N_15868,N_11054,N_14546);
or U15869 (N_15869,N_13937,N_11998);
or U15870 (N_15870,N_10843,N_11384);
or U15871 (N_15871,N_13344,N_10640);
nand U15872 (N_15872,N_14074,N_11869);
or U15873 (N_15873,N_11540,N_10939);
nand U15874 (N_15874,N_11772,N_14637);
and U15875 (N_15875,N_12721,N_13363);
nand U15876 (N_15876,N_11025,N_13249);
nor U15877 (N_15877,N_10388,N_14355);
and U15878 (N_15878,N_13315,N_13169);
or U15879 (N_15879,N_11849,N_13508);
or U15880 (N_15880,N_11454,N_11800);
nand U15881 (N_15881,N_12433,N_13237);
or U15882 (N_15882,N_14529,N_14894);
and U15883 (N_15883,N_11148,N_11014);
nand U15884 (N_15884,N_11891,N_13345);
or U15885 (N_15885,N_10393,N_12387);
and U15886 (N_15886,N_10890,N_11353);
nor U15887 (N_15887,N_10367,N_14616);
or U15888 (N_15888,N_14984,N_11796);
and U15889 (N_15889,N_11856,N_14072);
and U15890 (N_15890,N_12640,N_14462);
nor U15891 (N_15891,N_10646,N_14913);
nor U15892 (N_15892,N_12946,N_10720);
nor U15893 (N_15893,N_13619,N_13604);
or U15894 (N_15894,N_10059,N_12148);
nor U15895 (N_15895,N_14297,N_14446);
or U15896 (N_15896,N_13860,N_11137);
or U15897 (N_15897,N_14255,N_12677);
or U15898 (N_15898,N_12505,N_13320);
or U15899 (N_15899,N_11386,N_10566);
nor U15900 (N_15900,N_10217,N_11088);
and U15901 (N_15901,N_10703,N_10380);
or U15902 (N_15902,N_14758,N_12286);
nor U15903 (N_15903,N_11314,N_10376);
nand U15904 (N_15904,N_12743,N_13331);
and U15905 (N_15905,N_12426,N_14918);
nand U15906 (N_15906,N_14312,N_10934);
or U15907 (N_15907,N_14671,N_10620);
and U15908 (N_15908,N_12176,N_11208);
nor U15909 (N_15909,N_13422,N_13877);
nor U15910 (N_15910,N_14839,N_13000);
nor U15911 (N_15911,N_13994,N_12934);
and U15912 (N_15912,N_12305,N_11048);
nand U15913 (N_15913,N_13196,N_12829);
and U15914 (N_15914,N_14489,N_12264);
nand U15915 (N_15915,N_12028,N_10608);
nor U15916 (N_15916,N_12047,N_13087);
and U15917 (N_15917,N_12243,N_12442);
nand U15918 (N_15918,N_14449,N_11068);
nor U15919 (N_15919,N_12876,N_12468);
and U15920 (N_15920,N_14293,N_11843);
and U15921 (N_15921,N_12785,N_11675);
or U15922 (N_15922,N_10107,N_11397);
or U15923 (N_15923,N_14687,N_14774);
nor U15924 (N_15924,N_10665,N_12797);
and U15925 (N_15925,N_14923,N_13632);
and U15926 (N_15926,N_11893,N_11656);
nor U15927 (N_15927,N_11334,N_11110);
xor U15928 (N_15928,N_11422,N_13721);
and U15929 (N_15929,N_12838,N_12774);
and U15930 (N_15930,N_14438,N_11990);
nor U15931 (N_15931,N_13126,N_12678);
and U15932 (N_15932,N_14475,N_12726);
or U15933 (N_15933,N_13737,N_13767);
and U15934 (N_15934,N_12133,N_11091);
nand U15935 (N_15935,N_14124,N_12698);
nor U15936 (N_15936,N_14526,N_11053);
and U15937 (N_15937,N_14873,N_10716);
nor U15938 (N_15938,N_14120,N_13810);
nand U15939 (N_15939,N_11216,N_13471);
and U15940 (N_15940,N_14523,N_14986);
or U15941 (N_15941,N_14322,N_10840);
nor U15942 (N_15942,N_14461,N_11729);
nand U15943 (N_15943,N_10165,N_13912);
nor U15944 (N_15944,N_10049,N_14465);
nor U15945 (N_15945,N_13219,N_11619);
and U15946 (N_15946,N_12784,N_11538);
xnor U15947 (N_15947,N_14798,N_13312);
and U15948 (N_15948,N_13477,N_11326);
nor U15949 (N_15949,N_12717,N_10961);
or U15950 (N_15950,N_12096,N_14618);
or U15951 (N_15951,N_11363,N_12917);
nor U15952 (N_15952,N_14458,N_11774);
nor U15953 (N_15953,N_11961,N_11115);
nand U15954 (N_15954,N_14948,N_12649);
xor U15955 (N_15955,N_14027,N_12193);
or U15956 (N_15956,N_13056,N_10718);
nand U15957 (N_15957,N_12538,N_10248);
and U15958 (N_15958,N_11009,N_14615);
and U15959 (N_15959,N_14684,N_12632);
or U15960 (N_15960,N_14459,N_11567);
nand U15961 (N_15961,N_12552,N_11576);
or U15962 (N_15962,N_11204,N_12281);
nor U15963 (N_15963,N_10398,N_10098);
or U15964 (N_15964,N_11889,N_10563);
nand U15965 (N_15965,N_11581,N_13952);
nand U15966 (N_15966,N_12705,N_11065);
nor U15967 (N_15967,N_12960,N_10674);
nor U15968 (N_15968,N_11434,N_12495);
nand U15969 (N_15969,N_11551,N_11176);
nor U15970 (N_15970,N_13948,N_12016);
and U15971 (N_15971,N_10263,N_12500);
and U15972 (N_15972,N_13486,N_10695);
and U15973 (N_15973,N_11426,N_10790);
nor U15974 (N_15974,N_11594,N_13876);
nand U15975 (N_15975,N_13992,N_13691);
or U15976 (N_15976,N_12404,N_13273);
or U15977 (N_15977,N_14157,N_12852);
or U15978 (N_15978,N_10669,N_10405);
or U15979 (N_15979,N_12864,N_11513);
nand U15980 (N_15980,N_13740,N_13870);
nor U15981 (N_15981,N_14992,N_12470);
and U15982 (N_15982,N_12511,N_13997);
and U15983 (N_15983,N_13223,N_12102);
nor U15984 (N_15984,N_14996,N_13638);
nand U15985 (N_15985,N_10148,N_11956);
or U15986 (N_15986,N_12914,N_10926);
or U15987 (N_15987,N_12912,N_10936);
xor U15988 (N_15988,N_11364,N_13433);
or U15989 (N_15989,N_11942,N_12603);
nor U15990 (N_15990,N_10799,N_14008);
or U15991 (N_15991,N_14620,N_11220);
and U15992 (N_15992,N_13844,N_10198);
nor U15993 (N_15993,N_13047,N_13213);
and U15994 (N_15994,N_12920,N_12401);
nand U15995 (N_15995,N_10986,N_11736);
or U15996 (N_15996,N_10613,N_10572);
and U15997 (N_15997,N_14631,N_10115);
nand U15998 (N_15998,N_10395,N_14165);
xnor U15999 (N_15999,N_14797,N_13711);
nand U16000 (N_16000,N_13753,N_10507);
and U16001 (N_16001,N_14955,N_11939);
nor U16002 (N_16002,N_13615,N_11537);
nor U16003 (N_16003,N_13154,N_14814);
and U16004 (N_16004,N_11300,N_12942);
or U16005 (N_16005,N_11255,N_10782);
nor U16006 (N_16006,N_13942,N_11784);
and U16007 (N_16007,N_11401,N_12672);
nor U16008 (N_16008,N_10594,N_14815);
nor U16009 (N_16009,N_14113,N_13146);
nand U16010 (N_16010,N_11096,N_14500);
nor U16011 (N_16011,N_13963,N_10515);
nor U16012 (N_16012,N_11030,N_12941);
and U16013 (N_16013,N_13821,N_13380);
nand U16014 (N_16014,N_13923,N_10590);
and U16015 (N_16015,N_12030,N_12947);
and U16016 (N_16016,N_14199,N_12516);
nand U16017 (N_16017,N_10987,N_14678);
or U16018 (N_16018,N_13574,N_12441);
nor U16019 (N_16019,N_12463,N_12269);
or U16020 (N_16020,N_14079,N_14862);
nor U16021 (N_16021,N_11093,N_10145);
or U16022 (N_16022,N_13389,N_13406);
or U16023 (N_16023,N_12484,N_13218);
and U16024 (N_16024,N_10561,N_11161);
and U16025 (N_16025,N_12621,N_11783);
or U16026 (N_16026,N_11347,N_14573);
or U16027 (N_16027,N_12246,N_14608);
and U16028 (N_16028,N_10747,N_10209);
or U16029 (N_16029,N_12205,N_10180);
nand U16030 (N_16030,N_14677,N_14410);
nand U16031 (N_16031,N_10279,N_11103);
nor U16032 (N_16032,N_10562,N_14537);
and U16033 (N_16033,N_12610,N_10320);
nor U16034 (N_16034,N_12597,N_14031);
and U16035 (N_16035,N_11272,N_10419);
or U16036 (N_16036,N_11835,N_14591);
and U16037 (N_16037,N_14650,N_12294);
and U16038 (N_16038,N_11640,N_14602);
and U16039 (N_16039,N_14572,N_11558);
nor U16040 (N_16040,N_13306,N_13552);
nand U16041 (N_16041,N_10745,N_11447);
or U16042 (N_16042,N_11489,N_12700);
and U16043 (N_16043,N_10219,N_10848);
or U16044 (N_16044,N_12958,N_12296);
nor U16045 (N_16045,N_13968,N_14974);
nand U16046 (N_16046,N_14869,N_11764);
nor U16047 (N_16047,N_11613,N_11887);
or U16048 (N_16048,N_10661,N_12093);
and U16049 (N_16049,N_10112,N_14452);
and U16050 (N_16050,N_11239,N_14212);
nand U16051 (N_16051,N_12485,N_11996);
nand U16052 (N_16052,N_12572,N_11732);
nor U16053 (N_16053,N_11574,N_13578);
nand U16054 (N_16054,N_12884,N_11555);
nor U16055 (N_16055,N_11349,N_13976);
or U16056 (N_16056,N_10491,N_10020);
nand U16057 (N_16057,N_14403,N_12576);
nor U16058 (N_16058,N_10834,N_11311);
and U16059 (N_16059,N_11552,N_14387);
nor U16060 (N_16060,N_11657,N_11528);
and U16061 (N_16061,N_11283,N_12409);
nand U16062 (N_16062,N_11526,N_12775);
or U16063 (N_16063,N_14527,N_13162);
nand U16064 (N_16064,N_13724,N_13225);
nand U16065 (N_16065,N_11722,N_13068);
nor U16066 (N_16066,N_13920,N_14335);
or U16067 (N_16067,N_14519,N_13557);
and U16068 (N_16068,N_13316,N_13488);
nor U16069 (N_16069,N_13993,N_10347);
nor U16070 (N_16070,N_11214,N_10818);
nor U16071 (N_16071,N_11864,N_12447);
and U16072 (N_16072,N_13461,N_11365);
nor U16073 (N_16073,N_14715,N_10111);
or U16074 (N_16074,N_12924,N_12965);
xnor U16075 (N_16075,N_13733,N_14405);
or U16076 (N_16076,N_10757,N_11953);
or U16077 (N_16077,N_12489,N_10203);
or U16078 (N_16078,N_13863,N_10399);
nand U16079 (N_16079,N_14259,N_14802);
nand U16080 (N_16080,N_11168,N_10435);
and U16081 (N_16081,N_12673,N_14883);
or U16082 (N_16082,N_13092,N_13368);
nor U16083 (N_16083,N_14592,N_10256);
nand U16084 (N_16084,N_10974,N_11071);
or U16085 (N_16085,N_10678,N_11529);
and U16086 (N_16086,N_12574,N_10809);
and U16087 (N_16087,N_14082,N_13352);
nand U16088 (N_16088,N_13449,N_14005);
nand U16089 (N_16089,N_12768,N_12461);
or U16090 (N_16090,N_14253,N_11916);
or U16091 (N_16091,N_11549,N_12826);
and U16092 (N_16092,N_11666,N_11043);
or U16093 (N_16093,N_12616,N_13712);
and U16094 (N_16094,N_11432,N_12285);
and U16095 (N_16095,N_14524,N_10431);
nor U16096 (N_16096,N_13256,N_14551);
and U16097 (N_16097,N_11318,N_12242);
nand U16098 (N_16098,N_10460,N_11109);
nand U16099 (N_16099,N_10124,N_13786);
nand U16100 (N_16100,N_13879,N_12891);
nand U16101 (N_16101,N_14756,N_14399);
and U16102 (N_16102,N_11875,N_11323);
and U16103 (N_16103,N_11876,N_11140);
nand U16104 (N_16104,N_14437,N_11340);
or U16105 (N_16105,N_11257,N_11844);
or U16106 (N_16106,N_14302,N_10337);
xor U16107 (N_16107,N_10305,N_11322);
nor U16108 (N_16108,N_12771,N_13873);
and U16109 (N_16109,N_12403,N_13025);
nor U16110 (N_16110,N_13857,N_12385);
and U16111 (N_16111,N_10779,N_14133);
or U16112 (N_16112,N_10271,N_12397);
and U16113 (N_16113,N_10188,N_12197);
xor U16114 (N_16114,N_11312,N_10178);
nand U16115 (N_16115,N_12192,N_11361);
and U16116 (N_16116,N_11901,N_13299);
nand U16117 (N_16117,N_11645,N_10517);
nand U16118 (N_16118,N_14004,N_10972);
and U16119 (N_16119,N_10892,N_14767);
nor U16120 (N_16120,N_10290,N_10685);
or U16121 (N_16121,N_11899,N_12259);
or U16122 (N_16122,N_13808,N_10623);
nand U16123 (N_16123,N_13204,N_11948);
or U16124 (N_16124,N_14596,N_13887);
or U16125 (N_16125,N_10170,N_11816);
or U16126 (N_16126,N_13340,N_11616);
nor U16127 (N_16127,N_11823,N_13771);
or U16128 (N_16128,N_12079,N_10622);
nor U16129 (N_16129,N_14587,N_13614);
or U16130 (N_16130,N_10062,N_10006);
or U16131 (N_16131,N_13367,N_11476);
or U16132 (N_16132,N_11233,N_14920);
nand U16133 (N_16133,N_12418,N_14701);
nand U16134 (N_16134,N_13140,N_11575);
and U16135 (N_16135,N_12424,N_14070);
nor U16136 (N_16136,N_14217,N_13570);
and U16137 (N_16137,N_11822,N_12271);
and U16138 (N_16138,N_13794,N_12765);
nand U16139 (N_16139,N_12340,N_10909);
nand U16140 (N_16140,N_12670,N_10847);
and U16141 (N_16141,N_11499,N_13960);
nor U16142 (N_16142,N_10523,N_12122);
and U16143 (N_16143,N_13170,N_11674);
and U16144 (N_16144,N_10383,N_12423);
nand U16145 (N_16145,N_10581,N_12783);
and U16146 (N_16146,N_10758,N_12780);
or U16147 (N_16147,N_11237,N_13370);
nor U16148 (N_16148,N_11087,N_11921);
nor U16149 (N_16149,N_10787,N_10601);
and U16150 (N_16150,N_12571,N_14158);
and U16151 (N_16151,N_13224,N_10684);
or U16152 (N_16152,N_13491,N_10141);
or U16153 (N_16153,N_12393,N_13075);
or U16154 (N_16154,N_13770,N_11569);
nor U16155 (N_16155,N_11414,N_11070);
or U16156 (N_16156,N_10140,N_12906);
and U16157 (N_16157,N_10970,N_11742);
nand U16158 (N_16158,N_10345,N_13843);
nor U16159 (N_16159,N_11224,N_10663);
nand U16160 (N_16160,N_13918,N_13384);
nand U16161 (N_16161,N_14557,N_14481);
and U16162 (N_16162,N_12853,N_11954);
nor U16163 (N_16163,N_11686,N_11682);
nor U16164 (N_16164,N_13026,N_11005);
nand U16165 (N_16165,N_13435,N_14562);
or U16166 (N_16166,N_12653,N_11627);
and U16167 (N_16167,N_11766,N_11721);
nand U16168 (N_16168,N_12371,N_14171);
xor U16169 (N_16169,N_14625,N_12744);
or U16170 (N_16170,N_14468,N_11405);
nor U16171 (N_16171,N_12092,N_13110);
nand U16172 (N_16172,N_11370,N_13247);
or U16173 (N_16173,N_11206,N_10542);
nand U16174 (N_16174,N_11438,N_11515);
nand U16175 (N_16175,N_11456,N_14942);
or U16176 (N_16176,N_11113,N_14283);
or U16177 (N_16177,N_14576,N_14285);
and U16178 (N_16178,N_11543,N_10657);
nand U16179 (N_16179,N_10529,N_13819);
nand U16180 (N_16180,N_14448,N_11740);
nor U16181 (N_16181,N_10654,N_10591);
nand U16182 (N_16182,N_14413,N_14531);
nand U16183 (N_16183,N_12608,N_13738);
or U16184 (N_16184,N_13523,N_13353);
nand U16185 (N_16185,N_14638,N_14518);
or U16186 (N_16186,N_13301,N_12342);
nand U16187 (N_16187,N_14776,N_14330);
and U16188 (N_16188,N_10487,N_12377);
and U16189 (N_16189,N_10815,N_11496);
nor U16190 (N_16190,N_12186,N_11369);
or U16191 (N_16191,N_13412,N_13329);
nor U16192 (N_16192,N_14754,N_14622);
or U16193 (N_16193,N_14688,N_14532);
xnor U16194 (N_16194,N_10014,N_13657);
and U16195 (N_16195,N_11501,N_10714);
nor U16196 (N_16196,N_13909,N_12481);
or U16197 (N_16197,N_12085,N_13780);
and U16198 (N_16198,N_13744,N_11082);
nand U16199 (N_16199,N_11749,N_13761);
nand U16200 (N_16200,N_11604,N_13949);
xor U16201 (N_16201,N_14286,N_14197);
nor U16202 (N_16202,N_12199,N_10027);
and U16203 (N_16203,N_11226,N_13330);
nand U16204 (N_16204,N_12563,N_13418);
nand U16205 (N_16205,N_10771,N_13259);
and U16206 (N_16206,N_10418,N_12905);
or U16207 (N_16207,N_11440,N_12076);
nand U16208 (N_16208,N_11500,N_11290);
nor U16209 (N_16209,N_14301,N_11561);
nor U16210 (N_16210,N_14997,N_14870);
nand U16211 (N_16211,N_14783,N_12140);
nand U16212 (N_16212,N_14156,N_12437);
nand U16213 (N_16213,N_10185,N_10982);
or U16214 (N_16214,N_10397,N_11064);
or U16215 (N_16215,N_13260,N_11135);
or U16216 (N_16216,N_12392,N_13987);
nor U16217 (N_16217,N_13524,N_12619);
nand U16218 (N_16218,N_13377,N_13723);
nand U16219 (N_16219,N_12009,N_13540);
and U16220 (N_16220,N_13183,N_13481);
nand U16221 (N_16221,N_14011,N_14344);
and U16222 (N_16222,N_13336,N_10494);
nand U16223 (N_16223,N_13297,N_14886);
or U16224 (N_16224,N_12004,N_14654);
nor U16225 (N_16225,N_11918,N_11773);
or U16226 (N_16226,N_11873,N_13006);
and U16227 (N_16227,N_13112,N_10980);
nand U16228 (N_16228,N_14155,N_12022);
or U16229 (N_16229,N_11785,N_12951);
nand U16230 (N_16230,N_11521,N_10254);
nand U16231 (N_16231,N_14239,N_12149);
or U16232 (N_16232,N_14019,N_11152);
nor U16233 (N_16233,N_14276,N_11858);
nor U16234 (N_16234,N_14111,N_11597);
and U16235 (N_16235,N_12307,N_13277);
nor U16236 (N_16236,N_13423,N_10708);
or U16237 (N_16237,N_13514,N_14497);
xor U16238 (N_16238,N_12821,N_10074);
xor U16239 (N_16239,N_11992,N_14928);
or U16240 (N_16240,N_10264,N_11230);
or U16241 (N_16241,N_11685,N_14484);
and U16242 (N_16242,N_12304,N_13186);
and U16243 (N_16243,N_14480,N_13189);
and U16244 (N_16244,N_10776,N_13201);
or U16245 (N_16245,N_12880,N_10647);
nor U16246 (N_16246,N_11372,N_13010);
and U16247 (N_16247,N_12225,N_14221);
nor U16248 (N_16248,N_12787,N_10916);
nand U16249 (N_16249,N_12323,N_11605);
or U16250 (N_16250,N_14804,N_12177);
nor U16251 (N_16251,N_11664,N_12508);
nand U16252 (N_16252,N_14714,N_12697);
nor U16253 (N_16253,N_10871,N_14350);
nor U16254 (N_16254,N_14106,N_14610);
nor U16255 (N_16255,N_14508,N_10687);
nand U16256 (N_16256,N_11586,N_13308);
and U16257 (N_16257,N_10583,N_12635);
nor U16258 (N_16258,N_11963,N_11218);
nor U16259 (N_16259,N_10021,N_11847);
and U16260 (N_16260,N_12752,N_13825);
and U16261 (N_16261,N_12316,N_13687);
nor U16262 (N_16262,N_14478,N_10079);
nand U16263 (N_16263,N_14134,N_12535);
nand U16264 (N_16264,N_13541,N_11264);
nor U16265 (N_16265,N_11524,N_10370);
nor U16266 (N_16266,N_13304,N_13828);
nand U16267 (N_16267,N_12207,N_10930);
nand U16268 (N_16268,N_12344,N_12759);
nand U16269 (N_16269,N_10553,N_11307);
or U16270 (N_16270,N_14324,N_11863);
and U16271 (N_16271,N_11566,N_11443);
or U16272 (N_16272,N_13074,N_12578);
or U16273 (N_16273,N_14394,N_14014);
nand U16274 (N_16274,N_14246,N_14799);
and U16275 (N_16275,N_11655,N_12252);
and U16276 (N_16276,N_11183,N_12391);
nand U16277 (N_16277,N_11315,N_11694);
or U16278 (N_16278,N_13267,N_13785);
nor U16279 (N_16279,N_10549,N_12382);
nand U16280 (N_16280,N_11167,N_10302);
nand U16281 (N_16281,N_10754,N_14987);
nand U16282 (N_16282,N_12029,N_10860);
nor U16283 (N_16283,N_14077,N_12174);
and U16284 (N_16284,N_14193,N_11979);
and U16285 (N_16285,N_12351,N_11287);
or U16286 (N_16286,N_12986,N_14372);
nor U16287 (N_16287,N_10186,N_10810);
and U16288 (N_16288,N_11964,N_14770);
nor U16289 (N_16289,N_10108,N_14817);
and U16290 (N_16290,N_12050,N_10697);
and U16291 (N_16291,N_11795,N_10457);
and U16292 (N_16292,N_13222,N_11343);
nor U16293 (N_16293,N_13851,N_10832);
nor U16294 (N_16294,N_11584,N_12451);
nand U16295 (N_16295,N_10005,N_12645);
nor U16296 (N_16296,N_11554,N_12190);
and U16297 (N_16297,N_10285,N_13585);
nor U16298 (N_16298,N_10648,N_11731);
and U16299 (N_16299,N_10837,N_14771);
and U16300 (N_16300,N_11734,N_10603);
nor U16301 (N_16301,N_11945,N_12812);
nand U16302 (N_16302,N_12933,N_13888);
nor U16303 (N_16303,N_10508,N_11360);
xnor U16304 (N_16304,N_14571,N_10994);
nor U16305 (N_16305,N_14291,N_11578);
nor U16306 (N_16306,N_14569,N_12095);
nor U16307 (N_16307,N_12882,N_14439);
nor U16308 (N_16308,N_12773,N_11433);
or U16309 (N_16309,N_11097,N_13732);
or U16310 (N_16310,N_14130,N_11913);
or U16311 (N_16311,N_11470,N_11925);
nand U16312 (N_16312,N_11919,N_14884);
nor U16313 (N_16313,N_11199,N_11573);
and U16314 (N_16314,N_11718,N_14032);
nand U16315 (N_16315,N_11165,N_14495);
nand U16316 (N_16316,N_10761,N_12310);
nor U16317 (N_16317,N_10531,N_13796);
nor U16318 (N_16318,N_12805,N_14975);
or U16319 (N_16319,N_11634,N_10311);
or U16320 (N_16320,N_10227,N_14131);
nor U16321 (N_16321,N_12562,N_14451);
nand U16322 (N_16322,N_13072,N_12813);
or U16323 (N_16323,N_12913,N_12273);
nand U16324 (N_16324,N_13408,N_11962);
nand U16325 (N_16325,N_10656,N_11818);
and U16326 (N_16326,N_11639,N_13626);
nor U16327 (N_16327,N_12255,N_10927);
nor U16328 (N_16328,N_11061,N_13764);
or U16329 (N_16329,N_13314,N_14580);
nand U16330 (N_16330,N_10770,N_14367);
nor U16331 (N_16331,N_12959,N_12107);
nor U16332 (N_16332,N_10481,N_14233);
xor U16333 (N_16333,N_10495,N_13310);
and U16334 (N_16334,N_14183,N_14215);
or U16335 (N_16335,N_13774,N_14205);
nor U16336 (N_16336,N_14707,N_10576);
and U16337 (N_16337,N_14961,N_10903);
and U16338 (N_16338,N_14744,N_10841);
and U16339 (N_16339,N_12049,N_10277);
and U16340 (N_16340,N_11789,N_14663);
nand U16341 (N_16341,N_11090,N_10901);
nor U16342 (N_16342,N_11748,N_14807);
nand U16343 (N_16343,N_11668,N_10175);
and U16344 (N_16344,N_11705,N_11280);
nor U16345 (N_16345,N_10518,N_10193);
and U16346 (N_16346,N_10617,N_11915);
and U16347 (N_16347,N_13150,N_14889);
nand U16348 (N_16348,N_12261,N_11128);
and U16349 (N_16349,N_12634,N_11517);
or U16350 (N_16350,N_12498,N_11330);
and U16351 (N_16351,N_11089,N_14747);
nor U16352 (N_16352,N_13763,N_11085);
and U16353 (N_16353,N_11712,N_14831);
and U16354 (N_16354,N_10194,N_14400);
and U16355 (N_16355,N_13618,N_13361);
nand U16356 (N_16356,N_12848,N_12046);
or U16357 (N_16357,N_14282,N_11727);
or U16358 (N_16358,N_14245,N_14153);
and U16359 (N_16359,N_10830,N_10889);
nand U16360 (N_16360,N_12637,N_11223);
and U16361 (N_16361,N_10348,N_13520);
nand U16362 (N_16362,N_14015,N_14809);
nor U16363 (N_16363,N_12113,N_12191);
or U16364 (N_16364,N_10265,N_11607);
and U16365 (N_16365,N_13235,N_13921);
or U16366 (N_16366,N_10996,N_11130);
or U16367 (N_16367,N_11050,N_14041);
nor U16368 (N_16368,N_14007,N_10879);
nor U16369 (N_16369,N_10557,N_11037);
or U16370 (N_16370,N_10109,N_13364);
nor U16371 (N_16371,N_10412,N_14936);
nand U16372 (N_16372,N_10243,N_14722);
nor U16373 (N_16373,N_10067,N_13358);
and U16374 (N_16374,N_12868,N_14957);
nand U16375 (N_16375,N_13815,N_10234);
or U16376 (N_16376,N_14240,N_12012);
nand U16377 (N_16377,N_10439,N_13850);
or U16378 (N_16378,N_13266,N_14716);
or U16379 (N_16379,N_10377,N_14954);
nor U16380 (N_16380,N_10740,N_11041);
xor U16381 (N_16381,N_14326,N_13925);
nor U16382 (N_16382,N_11850,N_13924);
nor U16383 (N_16383,N_13512,N_13016);
nor U16384 (N_16384,N_14492,N_13338);
nor U16385 (N_16385,N_10734,N_14871);
nand U16386 (N_16386,N_13613,N_14912);
or U16387 (N_16387,N_10519,N_12791);
nand U16388 (N_16388,N_10247,N_13592);
nor U16389 (N_16389,N_13891,N_12112);
or U16390 (N_16390,N_12706,N_10184);
and U16391 (N_16391,N_10976,N_12040);
nand U16392 (N_16392,N_14509,N_11026);
nor U16393 (N_16393,N_14887,N_12352);
nor U16394 (N_16394,N_11415,N_11485);
and U16395 (N_16395,N_14287,N_10125);
and U16396 (N_16396,N_10070,N_14200);
and U16397 (N_16397,N_12166,N_10624);
nand U16398 (N_16398,N_10699,N_14434);
nand U16399 (N_16399,N_14985,N_13252);
nand U16400 (N_16400,N_11955,N_12055);
and U16401 (N_16401,N_10768,N_11403);
and U16402 (N_16402,N_11160,N_13018);
or U16403 (N_16403,N_11190,N_10907);
nor U16404 (N_16404,N_10925,N_13623);
or U16405 (N_16405,N_14621,N_14845);
nand U16406 (N_16406,N_10857,N_13429);
nand U16407 (N_16407,N_12361,N_11988);
nand U16408 (N_16408,N_11545,N_14035);
nor U16409 (N_16409,N_12908,N_11600);
or U16410 (N_16410,N_10513,N_13751);
xor U16411 (N_16411,N_11301,N_10702);
nand U16412 (N_16412,N_13008,N_13436);
nand U16413 (N_16413,N_12062,N_14821);
nor U16414 (N_16414,N_14868,N_14467);
and U16415 (N_16415,N_10414,N_13675);
or U16416 (N_16416,N_11078,N_10813);
and U16417 (N_16417,N_14632,N_12543);
and U16418 (N_16418,N_11804,N_12534);
nand U16419 (N_16419,N_12106,N_12110);
nand U16420 (N_16420,N_12065,N_12795);
nor U16421 (N_16421,N_13038,N_10979);
nor U16422 (N_16422,N_13752,N_13995);
nor U16423 (N_16423,N_11143,N_13202);
and U16424 (N_16424,N_10900,N_13641);
nor U16425 (N_16425,N_10918,N_10237);
and U16426 (N_16426,N_11381,N_11644);
nand U16427 (N_16427,N_10003,N_12586);
and U16428 (N_16428,N_11974,N_13291);
nor U16429 (N_16429,N_11809,N_12374);
nor U16430 (N_16430,N_11383,N_10123);
and U16431 (N_16431,N_10984,N_12127);
nor U16432 (N_16432,N_12596,N_12081);
and U16433 (N_16433,N_13940,N_10671);
or U16434 (N_16434,N_10294,N_13499);
nand U16435 (N_16435,N_14010,N_13192);
nor U16436 (N_16436,N_11959,N_12124);
nor U16437 (N_16437,N_14273,N_11643);
nor U16438 (N_16438,N_14140,N_11563);
nand U16439 (N_16439,N_11069,N_14093);
nand U16440 (N_16440,N_14262,N_14629);
nor U16441 (N_16441,N_14081,N_10722);
nand U16442 (N_16442,N_14012,N_12746);
or U16443 (N_16443,N_10844,N_11927);
or U16444 (N_16444,N_13041,N_13728);
or U16445 (N_16445,N_12738,N_14294);
nand U16446 (N_16446,N_13123,N_10760);
nand U16447 (N_16447,N_14317,N_12188);
nor U16448 (N_16448,N_14292,N_13525);
nor U16449 (N_16449,N_10437,N_12198);
nand U16450 (N_16450,N_12623,N_13178);
nor U16451 (N_16451,N_13284,N_14266);
nor U16452 (N_16452,N_13404,N_13250);
nand U16453 (N_16453,N_13321,N_13726);
nand U16454 (N_16454,N_10261,N_13883);
nor U16455 (N_16455,N_11993,N_13175);
nor U16456 (N_16456,N_10873,N_14623);
or U16457 (N_16457,N_11378,N_14068);
nor U16458 (N_16458,N_11531,N_11886);
and U16459 (N_16459,N_13116,N_13415);
and U16460 (N_16460,N_10952,N_11615);
nand U16461 (N_16461,N_14463,N_10788);
nor U16462 (N_16462,N_13133,N_13706);
or U16463 (N_16463,N_10453,N_12827);
xor U16464 (N_16464,N_13544,N_12238);
nor U16465 (N_16465,N_13784,N_11776);
nand U16466 (N_16466,N_10199,N_14030);
or U16467 (N_16467,N_11461,N_13067);
nand U16468 (N_16468,N_13951,N_12823);
nor U16469 (N_16469,N_14002,N_14315);
nand U16470 (N_16470,N_13319,N_12117);
nand U16471 (N_16471,N_12475,N_14321);
xnor U16472 (N_16472,N_13254,N_13121);
nand U16473 (N_16473,N_10597,N_11294);
nand U16474 (N_16474,N_11116,N_12856);
xor U16475 (N_16475,N_14763,N_12036);
and U16476 (N_16476,N_10400,N_14152);
or U16477 (N_16477,N_12024,N_14548);
nand U16478 (N_16478,N_12410,N_14303);
and U16479 (N_16479,N_14976,N_12502);
xor U16480 (N_16480,N_10066,N_11911);
nand U16481 (N_16481,N_11354,N_10426);
or U16482 (N_16482,N_14159,N_11409);
and U16483 (N_16483,N_12208,N_11104);
nand U16484 (N_16484,N_10698,N_14499);
and U16485 (N_16485,N_11121,N_11904);
nand U16486 (N_16486,N_11688,N_14820);
nor U16487 (N_16487,N_11101,N_12936);
nor U16488 (N_16488,N_10520,N_12206);
xor U16489 (N_16489,N_11225,N_12337);
nor U16490 (N_16490,N_13741,N_11511);
and U16491 (N_16491,N_11145,N_14728);
nand U16492 (N_16492,N_13665,N_14858);
nand U16493 (N_16493,N_14121,N_14359);
or U16494 (N_16494,N_10502,N_10983);
nand U16495 (N_16495,N_12215,N_12545);
or U16496 (N_16496,N_12598,N_13977);
nand U16497 (N_16497,N_13986,N_10312);
nand U16498 (N_16498,N_14222,N_13094);
nor U16499 (N_16499,N_10182,N_13120);
or U16500 (N_16500,N_10195,N_14762);
or U16501 (N_16501,N_11621,N_13907);
nor U16502 (N_16502,N_13981,N_10710);
xor U16503 (N_16503,N_13837,N_14743);
or U16504 (N_16504,N_14885,N_13174);
and U16505 (N_16505,N_13686,N_14761);
and U16506 (N_16506,N_14795,N_13034);
or U16507 (N_16507,N_10333,N_12222);
nor U16508 (N_16508,N_11976,N_10127);
nand U16509 (N_16509,N_14138,N_12355);
and U16510 (N_16510,N_11868,N_14110);
nor U16511 (N_16511,N_14485,N_10174);
and U16512 (N_16512,N_14828,N_13343);
or U16513 (N_16513,N_10679,N_10306);
or U16514 (N_16514,N_11211,N_11757);
nor U16515 (N_16515,N_11702,N_10632);
or U16516 (N_16516,N_11458,N_12849);
nor U16517 (N_16517,N_12886,N_14490);
nor U16518 (N_16518,N_14123,N_13536);
nor U16519 (N_16519,N_12173,N_14853);
nand U16520 (N_16520,N_11427,N_10181);
and U16521 (N_16521,N_12325,N_12665);
and U16522 (N_16522,N_10774,N_12999);
nor U16523 (N_16523,N_13180,N_10539);
nor U16524 (N_16524,N_13387,N_11536);
nand U16525 (N_16525,N_14237,N_10631);
nor U16526 (N_16526,N_12400,N_12014);
and U16527 (N_16527,N_14665,N_10466);
nor U16528 (N_16528,N_10524,N_13579);
or U16529 (N_16529,N_12336,N_12211);
xor U16530 (N_16530,N_14939,N_14851);
and U16531 (N_16531,N_12624,N_10958);
or U16532 (N_16532,N_14013,N_10527);
and U16533 (N_16533,N_12630,N_11253);
nor U16534 (N_16534,N_14510,N_14209);
and U16535 (N_16535,N_11562,N_13346);
nor U16536 (N_16536,N_13505,N_14428);
or U16537 (N_16537,N_10737,N_13722);
or U16538 (N_16538,N_12446,N_13528);
and U16539 (N_16539,N_12496,N_11271);
or U16540 (N_16540,N_13591,N_11127);
nor U16541 (N_16541,N_12613,N_11106);
nor U16542 (N_16542,N_11769,N_10268);
nor U16543 (N_16543,N_13941,N_14357);
and U16544 (N_16544,N_11492,N_10947);
or U16545 (N_16545,N_11298,N_12788);
and U16546 (N_16546,N_12817,N_11421);
xnor U16547 (N_16547,N_11118,N_11457);
or U16548 (N_16548,N_10977,N_13282);
or U16549 (N_16549,N_12770,N_10766);
nor U16550 (N_16550,N_12745,N_12707);
nand U16551 (N_16551,N_14705,N_11417);
nand U16552 (N_16552,N_12681,N_14973);
nand U16553 (N_16553,N_13668,N_11711);
and U16554 (N_16554,N_12104,N_10913);
and U16555 (N_16555,N_13265,N_11086);
nor U16556 (N_16556,N_11651,N_13674);
nand U16557 (N_16557,N_13159,N_14249);
and U16558 (N_16558,N_14176,N_11908);
or U16559 (N_16559,N_11502,N_14181);
nor U16560 (N_16560,N_11019,N_14953);
or U16561 (N_16561,N_13962,N_10266);
or U16562 (N_16562,N_12919,N_11446);
or U16563 (N_16563,N_11142,N_12529);
nor U16564 (N_16564,N_13817,N_13846);
nand U16565 (N_16565,N_11483,N_11235);
and U16566 (N_16566,N_14558,N_12878);
nor U16567 (N_16567,N_10117,N_14382);
nand U16568 (N_16568,N_13195,N_12078);
nand U16569 (N_16569,N_14393,N_10240);
or U16570 (N_16570,N_11525,N_12975);
and U16571 (N_16571,N_13945,N_14270);
nor U16572 (N_16572,N_11189,N_13841);
nand U16573 (N_16573,N_14418,N_12894);
nor U16574 (N_16574,N_12143,N_13513);
xnor U16575 (N_16575,N_13106,N_10110);
nor U16576 (N_16576,N_10359,N_10138);
nand U16577 (N_16577,N_12858,N_14017);
and U16578 (N_16578,N_11125,N_12105);
or U16579 (N_16579,N_11626,N_11840);
xnor U16580 (N_16580,N_14182,N_11020);
and U16581 (N_16581,N_11632,N_11049);
nor U16582 (N_16582,N_10606,N_13898);
and U16583 (N_16583,N_11031,N_10619);
or U16584 (N_16584,N_11393,N_11066);
or U16585 (N_16585,N_12422,N_14811);
nor U16586 (N_16586,N_10759,N_12021);
nand U16587 (N_16587,N_11888,N_13036);
and U16588 (N_16588,N_12396,N_12560);
or U16589 (N_16589,N_10677,N_14455);
nor U16590 (N_16590,N_12740,N_11518);
nand U16591 (N_16591,N_12679,N_12415);
nor U16592 (N_16592,N_11900,N_13768);
and U16593 (N_16593,N_11481,N_10501);
nand U16594 (N_16594,N_10037,N_13908);
or U16595 (N_16595,N_12703,N_10923);
nand U16596 (N_16596,N_10050,N_10462);
or U16597 (N_16597,N_13465,N_13278);
or U16598 (N_16598,N_12010,N_10363);
xnor U16599 (N_16599,N_13309,N_14512);
nor U16600 (N_16600,N_14534,N_10207);
and U16601 (N_16601,N_10224,N_12499);
xnor U16602 (N_16602,N_10391,N_10214);
nand U16603 (N_16603,N_14381,N_12278);
nor U16604 (N_16604,N_14295,N_11015);
nand U16605 (N_16605,N_12088,N_11940);
nor U16606 (N_16606,N_12845,N_12555);
or U16607 (N_16607,N_12733,N_12641);
nor U16608 (N_16608,N_10288,N_13500);
xnor U16609 (N_16609,N_10099,N_12974);
or U16610 (N_16610,N_10205,N_10688);
and U16611 (N_16611,N_12724,N_10339);
nor U16612 (N_16612,N_12202,N_14536);
and U16613 (N_16613,N_12100,N_14289);
and U16614 (N_16614,N_10361,N_10846);
and U16615 (N_16615,N_14837,N_10314);
nor U16616 (N_16616,N_12758,N_10340);
or U16617 (N_16617,N_12952,N_14426);
nor U16618 (N_16618,N_14208,N_10965);
or U16619 (N_16619,N_14250,N_14888);
xor U16620 (N_16620,N_10012,N_12694);
or U16621 (N_16621,N_13735,N_12611);
nand U16622 (N_16622,N_13685,N_10625);
and U16623 (N_16623,N_12844,N_13931);
and U16624 (N_16624,N_10441,N_11690);
nor U16625 (N_16625,N_13978,N_12825);
nor U16626 (N_16626,N_11851,N_11477);
and U16627 (N_16627,N_14314,N_11971);
nand U16628 (N_16628,N_13001,N_12386);
nor U16629 (N_16629,N_10019,N_14473);
xnor U16630 (N_16630,N_11465,N_12120);
nor U16631 (N_16631,N_10454,N_12748);
or U16632 (N_16632,N_10029,N_10233);
nand U16633 (N_16633,N_13664,N_14626);
nor U16634 (N_16634,N_11512,N_13802);
or U16635 (N_16635,N_14612,N_12659);
nor U16636 (N_16636,N_11704,N_10921);
or U16637 (N_16637,N_11745,N_11040);
and U16638 (N_16638,N_13750,N_13868);
or U16639 (N_16639,N_14309,N_11182);
nand U16640 (N_16640,N_13680,N_10360);
nand U16641 (N_16641,N_11338,N_14271);
or U16642 (N_16642,N_11853,N_13226);
nor U16643 (N_16643,N_10521,N_14775);
and U16644 (N_16644,N_10382,N_10962);
nand U16645 (N_16645,N_14597,N_12591);
or U16646 (N_16646,N_13111,N_12895);
nor U16647 (N_16647,N_12889,N_10735);
and U16648 (N_16648,N_13934,N_11355);
and U16649 (N_16649,N_13560,N_10911);
nand U16650 (N_16650,N_11592,N_14346);
and U16651 (N_16651,N_14601,N_10851);
nor U16652 (N_16652,N_14830,N_12638);
nand U16653 (N_16653,N_10328,N_10558);
or U16654 (N_16654,N_10526,N_11646);
and U16655 (N_16655,N_13695,N_12888);
and U16656 (N_16656,N_13648,N_13396);
and U16657 (N_16657,N_13089,N_10177);
and U16658 (N_16658,N_13842,N_12693);
or U16659 (N_16659,N_13467,N_11741);
or U16660 (N_16660,N_10083,N_12295);
nand U16661 (N_16661,N_12209,N_13376);
and U16662 (N_16662,N_14102,N_11442);
or U16663 (N_16663,N_13439,N_10571);
or U16664 (N_16664,N_13143,N_13354);
or U16665 (N_16665,N_14989,N_11337);
or U16666 (N_16666,N_11700,N_12163);
nand U16667 (N_16667,N_10798,N_13646);
nor U16668 (N_16668,N_13562,N_10269);
and U16669 (N_16669,N_10800,N_14867);
and U16670 (N_16670,N_14651,N_12240);
xnor U16671 (N_16671,N_10694,N_12115);
nand U16672 (N_16672,N_13102,N_13554);
or U16673 (N_16673,N_12633,N_14244);
xor U16674 (N_16674,N_13718,N_11200);
and U16675 (N_16675,N_11256,N_10691);
xor U16676 (N_16676,N_10878,N_14095);
or U16677 (N_16677,N_13597,N_13696);
nand U16678 (N_16678,N_11720,N_13690);
nand U16679 (N_16679,N_14604,N_13356);
nor U16680 (N_16680,N_13114,N_11786);
nor U16681 (N_16681,N_11695,N_11672);
and U16682 (N_16682,N_14861,N_11289);
or U16683 (N_16683,N_10595,N_12966);
or U16684 (N_16684,N_12727,N_12760);
nor U16685 (N_16685,N_12921,N_12776);
nand U16686 (N_16686,N_12684,N_11284);
and U16687 (N_16687,N_13132,N_11196);
nor U16688 (N_16688,N_14269,N_14941);
nor U16689 (N_16689,N_10693,N_11406);
nor U16690 (N_16690,N_11108,N_11138);
or U16691 (N_16691,N_11880,N_11498);
nand U16692 (N_16692,N_10151,N_11162);
and U16693 (N_16693,N_12929,N_13534);
or U16694 (N_16694,N_13905,N_13100);
nand U16695 (N_16695,N_12664,N_14091);
or U16696 (N_16696,N_13616,N_12051);
or U16697 (N_16697,N_11059,N_11490);
nand U16698 (N_16698,N_12356,N_12865);
xor U16699 (N_16699,N_13587,N_10973);
and U16700 (N_16700,N_14787,N_11359);
or U16701 (N_16701,N_14417,N_11648);
nor U16702 (N_16702,N_11808,N_12718);
nand U16703 (N_16703,N_12118,N_11728);
nand U16704 (N_16704,N_10744,N_12487);
or U16705 (N_16705,N_13161,N_13208);
and U16706 (N_16706,N_11867,N_13984);
nor U16707 (N_16707,N_13943,N_10728);
nand U16708 (N_16708,N_14545,N_12615);
or U16709 (N_16709,N_13300,N_13469);
or U16710 (N_16710,N_12480,N_10101);
or U16711 (N_16711,N_12212,N_14865);
or U16712 (N_16712,N_12910,N_13327);
or U16713 (N_16713,N_11056,N_11817);
nor U16714 (N_16714,N_11429,N_11213);
nor U16715 (N_16715,N_14929,N_10445);
nand U16716 (N_16716,N_10450,N_10272);
or U16717 (N_16717,N_12262,N_13073);
nor U16718 (N_16718,N_11946,N_13793);
and U16719 (N_16719,N_13896,N_14476);
nor U16720 (N_16720,N_11917,N_11637);
nor U16721 (N_16721,N_11240,N_10655);
and U16722 (N_16722,N_11854,N_12778);
nand U16723 (N_16723,N_10055,N_11141);
nor U16724 (N_16724,N_10477,N_13497);
nor U16725 (N_16725,N_12301,N_11222);
and U16726 (N_16726,N_14494,N_13440);
nor U16727 (N_16727,N_14659,N_11606);
nor U16728 (N_16728,N_11676,N_12518);
nor U16729 (N_16729,N_10038,N_10471);
or U16730 (N_16730,N_14796,N_13079);
and U16731 (N_16731,N_13911,N_12902);
and U16732 (N_16732,N_14003,N_10212);
or U16733 (N_16733,N_12802,N_11124);
and U16734 (N_16734,N_14502,N_14600);
nand U16735 (N_16735,N_13448,N_13694);
nor U16736 (N_16736,N_10044,N_11469);
and U16737 (N_16737,N_10887,N_12019);
nor U16738 (N_16738,N_12939,N_14850);
and U16739 (N_16739,N_13558,N_13734);
or U16740 (N_16740,N_13729,N_12231);
nand U16741 (N_16741,N_14118,N_13498);
or U16742 (N_16742,N_13292,N_13339);
nor U16743 (N_16743,N_13264,N_13240);
nor U16744 (N_16744,N_12622,N_12734);
nand U16745 (N_16745,N_10805,N_14749);
nand U16746 (N_16746,N_14290,N_12674);
nor U16747 (N_16747,N_11649,N_13575);
or U16748 (N_16748,N_11819,N_14860);
nand U16749 (N_16749,N_11753,N_13402);
and U16750 (N_16750,N_11788,N_13166);
or U16751 (N_16751,N_11947,N_12218);
nor U16752 (N_16752,N_12581,N_11642);
or U16753 (N_16753,N_14812,N_10533);
and U16754 (N_16754,N_11408,N_12136);
nor U16755 (N_16755,N_14220,N_13393);
nor U16756 (N_16756,N_14516,N_13567);
and U16757 (N_16757,N_13530,N_12970);
or U16758 (N_16758,N_13152,N_14026);
or U16759 (N_16759,N_13125,N_13236);
or U16760 (N_16760,N_12293,N_10917);
nand U16761 (N_16761,N_13494,N_11374);
nor U16762 (N_16762,N_12080,N_13566);
or U16763 (N_16763,N_11568,N_11553);
nand U16764 (N_16764,N_13758,N_12988);
nor U16765 (N_16765,N_13715,N_13109);
nand U16766 (N_16766,N_14105,N_13088);
or U16767 (N_16767,N_14168,N_14022);
and U16768 (N_16768,N_14769,N_12350);
and U16769 (N_16769,N_13645,N_11944);
nand U16770 (N_16770,N_12056,N_10469);
nand U16771 (N_16771,N_10801,N_12256);
and U16772 (N_16772,N_13899,N_14943);
nor U16773 (N_16773,N_10260,N_14938);
nor U16774 (N_16774,N_13985,N_12497);
nor U16775 (N_16775,N_14915,N_13939);
nor U16776 (N_16776,N_12159,N_13529);
nor U16777 (N_16777,N_12427,N_10374);
and U16778 (N_16778,N_10190,N_13594);
and U16779 (N_16779,N_13773,N_14264);
xor U16780 (N_16780,N_13902,N_11348);
xor U16781 (N_16781,N_11698,N_14164);
nor U16782 (N_16782,N_13424,N_10215);
and U16783 (N_16783,N_10026,N_14258);
or U16784 (N_16784,N_11120,N_10016);
or U16785 (N_16785,N_10652,N_11951);
or U16786 (N_16786,N_14547,N_10459);
nor U16787 (N_16787,N_12756,N_12372);
nor U16788 (N_16788,N_10467,N_12735);
nor U16789 (N_16789,N_11924,N_12123);
or U16790 (N_16790,N_14058,N_10071);
or U16791 (N_16791,N_13158,N_12315);
nand U16792 (N_16792,N_10292,N_12395);
or U16793 (N_16793,N_11175,N_12542);
nand U16794 (N_16794,N_11860,N_11366);
and U16795 (N_16795,N_10095,N_10394);
or U16796 (N_16796,N_10942,N_12221);
nand U16797 (N_16797,N_14501,N_12464);
nand U16798 (N_16798,N_14838,N_11413);
nand U16799 (N_16799,N_13065,N_12398);
nor U16800 (N_16800,N_12614,N_11781);
or U16801 (N_16801,N_12512,N_14633);
and U16802 (N_16802,N_13167,N_10051);
nor U16803 (N_16803,N_14893,N_12449);
nand U16804 (N_16804,N_10396,N_13021);
nand U16805 (N_16805,N_13944,N_14833);
nor U16806 (N_16806,N_14443,N_10171);
and U16807 (N_16807,N_10773,N_10825);
and U16808 (N_16808,N_12675,N_11497);
or U16809 (N_16809,N_10956,N_13107);
nor U16810 (N_16810,N_11234,N_12435);
or U16811 (N_16811,N_11039,N_13080);
xnor U16812 (N_16812,N_11480,N_14742);
or U16813 (N_16813,N_11044,N_14810);
or U16814 (N_16814,N_10063,N_13611);
and U16815 (N_16815,N_13621,N_14740);
and U16816 (N_16816,N_12950,N_14498);
nor U16817 (N_16817,N_14563,N_13108);
nor U16818 (N_16818,N_13239,N_13795);
nor U16819 (N_16819,N_13549,N_10428);
and U16820 (N_16820,N_11400,N_13697);
nand U16821 (N_16821,N_13598,N_10668);
nand U16822 (N_16822,N_13913,N_11679);
nand U16823 (N_16823,N_14191,N_14528);
nor U16824 (N_16824,N_12251,N_11228);
or U16825 (N_16825,N_13007,N_11107);
nor U16826 (N_16826,N_13688,N_14487);
and U16827 (N_16827,N_12322,N_11158);
nand U16828 (N_16828,N_10490,N_11008);
xor U16829 (N_16829,N_10967,N_12807);
and U16830 (N_16830,N_12722,N_13076);
nand U16831 (N_16831,N_11399,N_11418);
nand U16832 (N_16832,N_14916,N_13634);
or U16833 (N_16833,N_13458,N_14727);
nor U16834 (N_16834,N_12723,N_10604);
or U16835 (N_16835,N_11716,N_11802);
nand U16836 (N_16836,N_12438,N_14731);
nor U16837 (N_16837,N_13548,N_13274);
and U16838 (N_16838,N_11428,N_14805);
nand U16839 (N_16839,N_10819,N_12018);
nand U16840 (N_16840,N_12026,N_13288);
and U16841 (N_16841,N_14241,N_10472);
or U16842 (N_16842,N_12493,N_11352);
nand U16843 (N_16843,N_11482,N_10392);
or U16844 (N_16844,N_10033,N_12981);
or U16845 (N_16845,N_11371,N_14788);
and U16846 (N_16846,N_12020,N_14878);
and U16847 (N_16847,N_12146,N_10510);
and U16848 (N_16848,N_12309,N_11765);
nand U16849 (N_16849,N_10503,N_13359);
and U16850 (N_16850,N_14029,N_13019);
or U16851 (N_16851,N_12683,N_13988);
nand U16852 (N_16852,N_14606,N_14000);
nand U16853 (N_16853,N_10991,N_11931);
or U16854 (N_16854,N_12553,N_13188);
nor U16855 (N_16855,N_14039,N_12814);
nor U16856 (N_16856,N_11475,N_10456);
or U16857 (N_16857,N_10666,N_10088);
nand U16858 (N_16858,N_14574,N_12907);
nor U16859 (N_16859,N_10371,N_12380);
nor U16860 (N_16860,N_10280,N_10500);
nand U16861 (N_16861,N_10389,N_12233);
and U16862 (N_16862,N_10789,N_14373);
nand U16863 (N_16863,N_10257,N_11832);
nand U16864 (N_16864,N_12873,N_12456);
or U16865 (N_16865,N_11310,N_11798);
or U16866 (N_16866,N_12306,N_10474);
or U16867 (N_16867,N_12445,N_10935);
or U16868 (N_16868,N_12945,N_12170);
and U16869 (N_16869,N_14097,N_13826);
and U16870 (N_16870,N_10582,N_13395);
and U16871 (N_16871,N_13765,N_11285);
and U16872 (N_16872,N_14588,N_13953);
nor U16873 (N_16873,N_14673,N_12167);
nor U16874 (N_16874,N_11380,N_13791);
nor U16875 (N_16875,N_14189,N_10551);
xnor U16876 (N_16876,N_11806,N_10411);
or U16877 (N_16877,N_12013,N_14166);
or U16878 (N_16878,N_12037,N_14184);
and U16879 (N_16879,N_14218,N_12569);
nand U16880 (N_16880,N_10251,N_10407);
and U16881 (N_16881,N_13929,N_12558);
nor U16882 (N_16882,N_12476,N_13832);
nor U16883 (N_16883,N_12444,N_12754);
or U16884 (N_16884,N_11209,N_13427);
nor U16885 (N_16885,N_10149,N_12925);
or U16886 (N_16886,N_14917,N_11678);
or U16887 (N_16887,N_13035,N_13501);
nor U16888 (N_16888,N_10953,N_13173);
or U16889 (N_16889,N_10197,N_12506);
and U16890 (N_16890,N_11052,N_13874);
and U16891 (N_16891,N_12180,N_14752);
and U16892 (N_16892,N_14919,N_13568);
and U16893 (N_16893,N_10326,N_13861);
nand U16894 (N_16894,N_14579,N_14777);
nand U16895 (N_16895,N_13490,N_14423);
or U16896 (N_16896,N_12867,N_11132);
nor U16897 (N_16897,N_10364,N_11905);
and U16898 (N_16898,N_12904,N_10992);
nor U16899 (N_16899,N_12944,N_10564);
xor U16900 (N_16900,N_14388,N_11926);
nand U16901 (N_16901,N_10317,N_10159);
nor U16902 (N_16902,N_10004,N_11579);
or U16903 (N_16903,N_13450,N_14190);
nand U16904 (N_16904,N_14504,N_12267);
nand U16905 (N_16905,N_10966,N_13716);
or U16906 (N_16906,N_10468,N_10335);
or U16907 (N_16907,N_12685,N_11133);
or U16908 (N_16908,N_13545,N_14800);
nand U16909 (N_16909,N_11703,N_11997);
and U16910 (N_16910,N_11217,N_12244);
nor U16911 (N_16911,N_12431,N_11194);
or U16912 (N_16912,N_13350,N_14720);
nor U16913 (N_16913,N_13086,N_14932);
and U16914 (N_16914,N_12317,N_10605);
nand U16915 (N_16915,N_13858,N_13527);
nor U16916 (N_16916,N_10731,N_12808);
nor U16917 (N_16917,N_14639,N_11279);
or U16918 (N_16918,N_13862,N_13064);
nand U16919 (N_16919,N_12875,N_13502);
and U16920 (N_16920,N_11246,N_11459);
or U16921 (N_16921,N_12687,N_14402);
or U16922 (N_16922,N_13678,N_11391);
or U16923 (N_16923,N_13830,N_12436);
nand U16924 (N_16924,N_10637,N_10086);
xnor U16925 (N_16925,N_12661,N_13782);
nor U16926 (N_16926,N_12086,N_13776);
and U16927 (N_16927,N_11609,N_10187);
and U16928 (N_16928,N_10429,N_12658);
nand U16929 (N_16929,N_12979,N_10736);
nor U16930 (N_16930,N_14142,N_13251);
xnor U16931 (N_16931,N_13332,N_14136);
and U16932 (N_16932,N_14944,N_14175);
or U16933 (N_16933,N_11669,N_13371);
nand U16934 (N_16934,N_13411,N_10081);
or U16935 (N_16935,N_13603,N_10496);
or U16936 (N_16936,N_13736,N_11265);
and U16937 (N_16937,N_13420,N_12993);
or U16938 (N_16938,N_14514,N_12165);
nor U16939 (N_16939,N_13482,N_10091);
or U16940 (N_16940,N_12175,N_13950);
and U16941 (N_16941,N_12406,N_13269);
nor U16942 (N_16942,N_11170,N_10877);
nor U16943 (N_16943,N_12847,N_12666);
or U16944 (N_16944,N_12935,N_13144);
or U16945 (N_16945,N_12660,N_10938);
and U16946 (N_16946,N_10548,N_13969);
nor U16947 (N_16947,N_13151,N_12729);
nand U16948 (N_16948,N_11273,N_12587);
xor U16949 (N_16949,N_13480,N_11630);
nor U16950 (N_16950,N_13700,N_11157);
nor U16951 (N_16951,N_11624,N_11395);
nand U16952 (N_16952,N_11829,N_13027);
and U16953 (N_16953,N_13910,N_10211);
or U16954 (N_16954,N_11768,N_13096);
nand U16955 (N_16955,N_13748,N_14926);
nand U16956 (N_16956,N_12704,N_12275);
nor U16957 (N_16957,N_11250,N_10751);
or U16958 (N_16958,N_11038,N_11771);
or U16959 (N_16959,N_10169,N_10707);
nor U16960 (N_16960,N_10682,N_11852);
nand U16961 (N_16961,N_12600,N_12584);
nand U16962 (N_16962,N_11153,N_10458);
nand U16963 (N_16963,N_10855,N_14268);
nand U16964 (N_16964,N_12762,N_11699);
nor U16965 (N_16965,N_13234,N_13563);
nor U16966 (N_16966,N_10308,N_12822);
nand U16967 (N_16967,N_13518,N_13397);
nor U16968 (N_16968,N_10299,N_13609);
or U16969 (N_16969,N_12098,N_10948);
and U16970 (N_16970,N_11259,N_13351);
or U16971 (N_16971,N_11100,N_12647);
nand U16972 (N_16972,N_12654,N_10118);
nor U16973 (N_16973,N_12636,N_12074);
and U16974 (N_16974,N_13417,N_13827);
nand U16975 (N_16975,N_11833,N_12589);
and U16976 (N_16976,N_13789,N_13836);
and U16977 (N_16977,N_11680,N_13122);
xnor U16978 (N_16978,N_11193,N_10220);
and U16979 (N_16979,N_11754,N_11317);
nor U16980 (N_16980,N_14757,N_10416);
xnor U16981 (N_16981,N_14801,N_14643);
and U16982 (N_16982,N_12289,N_11966);
or U16983 (N_16983,N_10433,N_14328);
or U16984 (N_16984,N_14607,N_12138);
and U16985 (N_16985,N_10593,N_10287);
nand U16986 (N_16986,N_14595,N_12279);
nand U16987 (N_16987,N_12682,N_12551);
or U16988 (N_16988,N_12739,N_12189);
or U16989 (N_16989,N_11830,N_11205);
nor U16990 (N_16990,N_11034,N_10680);
and U16991 (N_16991,N_13324,N_10749);
nor U16992 (N_16992,N_11857,N_12815);
and U16993 (N_16993,N_10082,N_13263);
nor U16994 (N_16994,N_11841,N_14050);
nand U16995 (N_16995,N_12927,N_10238);
nor U16996 (N_16996,N_13244,N_13430);
nand U16997 (N_16997,N_10226,N_14978);
nor U16998 (N_16998,N_13628,N_10990);
nor U16999 (N_16999,N_13200,N_14648);
xor U17000 (N_17000,N_14390,N_13342);
or U17001 (N_17001,N_12879,N_14444);
or U17002 (N_17002,N_13547,N_13596);
and U17003 (N_17003,N_13652,N_12308);
and U17004 (N_17004,N_11874,N_14435);
or U17005 (N_17005,N_14320,N_13451);
nand U17006 (N_17006,N_10975,N_12741);
nor U17007 (N_17007,N_14906,N_11930);
or U17008 (N_17008,N_14960,N_12871);
and U17009 (N_17009,N_14040,N_12595);
and U17010 (N_17010,N_14386,N_14092);
and U17011 (N_17011,N_14910,N_11556);
and U17012 (N_17012,N_13246,N_11293);
nor U17013 (N_17013,N_13903,N_11894);
and U17014 (N_17014,N_12023,N_14471);
or U17015 (N_17015,N_13869,N_10797);
nor U17016 (N_17016,N_14682,N_10386);
nand U17017 (N_17017,N_10516,N_13369);
nand U17018 (N_17018,N_14818,N_14345);
and U17019 (N_17019,N_11544,N_10351);
nor U17020 (N_17020,N_13137,N_13653);
or U17021 (N_17021,N_14277,N_13593);
and U17022 (N_17022,N_12714,N_10585);
and U17023 (N_17023,N_14556,N_10778);
nor U17024 (N_17024,N_13872,N_11473);
or U17025 (N_17025,N_10421,N_13296);
nand U17026 (N_17026,N_13479,N_12237);
nand U17027 (N_17027,N_11872,N_12646);
and U17028 (N_17028,N_13070,N_13650);
nor U17029 (N_17029,N_14395,N_14227);
nand U17030 (N_17030,N_12994,N_10532);
and U17031 (N_17031,N_10514,N_14876);
nor U17032 (N_17032,N_11778,N_14278);
or U17033 (N_17033,N_13709,N_11557);
or U17034 (N_17034,N_10341,N_14109);
and U17035 (N_17035,N_12064,N_11960);
nor U17036 (N_17036,N_10486,N_10356);
nand U17037 (N_17037,N_11134,N_10479);
and U17038 (N_17038,N_14738,N_11171);
or U17039 (N_17039,N_14147,N_14377);
or U17040 (N_17040,N_13816,N_11906);
nor U17041 (N_17041,N_13379,N_12513);
or U17042 (N_17042,N_14440,N_13305);
and U17043 (N_17043,N_11522,N_12346);
nand U17044 (N_17044,N_10602,N_12077);
nand U17045 (N_17045,N_11831,N_13656);
nand U17046 (N_17046,N_10286,N_13900);
nor U17047 (N_17047,N_12926,N_14730);
nor U17048 (N_17048,N_10653,N_13979);
nor U17049 (N_17049,N_13328,N_11738);
or U17050 (N_17050,N_11227,N_14422);
and U17051 (N_17051,N_14043,N_12713);
and U17052 (N_17052,N_14135,N_10378);
nor U17053 (N_17053,N_13537,N_14676);
nand U17054 (N_17054,N_11914,N_14605);
or U17055 (N_17055,N_14432,N_14712);
xnor U17056 (N_17056,N_10309,N_12292);
nand U17057 (N_17057,N_10057,N_14464);
nor U17058 (N_17058,N_14054,N_12457);
nor U17059 (N_17059,N_10628,N_11689);
or U17060 (N_17060,N_11450,N_13662);
xnor U17061 (N_17061,N_14967,N_14327);
nand U17062 (N_17062,N_10417,N_14647);
or U17063 (N_17063,N_11376,N_10422);
and U17064 (N_17064,N_14856,N_10568);
or U17065 (N_17065,N_12909,N_11379);
and U17066 (N_17066,N_11834,N_13967);
xor U17067 (N_17067,N_11491,N_11402);
nor U17068 (N_17068,N_12763,N_10096);
and U17069 (N_17069,N_10592,N_12991);
and U17070 (N_17070,N_14034,N_10094);
or U17071 (N_17071,N_13124,N_14824);
nor U17072 (N_17072,N_12725,N_10160);
or U17073 (N_17073,N_14994,N_12737);
nor U17074 (N_17074,N_12696,N_10888);
or U17075 (N_17075,N_14090,N_12899);
and U17076 (N_17076,N_13972,N_12676);
or U17077 (N_17077,N_11779,N_10512);
nor U17078 (N_17078,N_11394,N_14100);
or U17079 (N_17079,N_13705,N_11244);
xor U17080 (N_17080,N_12473,N_10162);
and U17081 (N_17081,N_14866,N_13390);
nor U17082 (N_17082,N_11042,N_10865);
and U17083 (N_17083,N_10318,N_14704);
or U17084 (N_17084,N_11572,N_12239);
and U17085 (N_17085,N_12184,N_12408);
nand U17086 (N_17086,N_14909,N_13719);
nor U17087 (N_17087,N_10932,N_10861);
nor U17088 (N_17088,N_10368,N_14535);
or U17089 (N_17089,N_13258,N_14668);
nor U17090 (N_17090,N_13590,N_14429);
nor U17091 (N_17091,N_10273,N_11268);
and U17092 (N_17092,N_11309,N_13313);
xnor U17093 (N_17093,N_13787,N_10919);
or U17094 (N_17094,N_14044,N_13871);
and U17095 (N_17095,N_14505,N_11195);
nand U17096 (N_17096,N_10536,N_11022);
and U17097 (N_17097,N_12592,N_14790);
nor U17098 (N_17098,N_12990,N_14566);
xnor U17099 (N_17099,N_12689,N_13745);
nor U17100 (N_17100,N_12580,N_10365);
nor U17101 (N_17101,N_11577,N_11541);
nor U17102 (N_17102,N_10964,N_10854);
or U17103 (N_17103,N_14260,N_12204);
and U17104 (N_17104,N_14703,N_12818);
nor U17105 (N_17105,N_14846,N_12223);
nor U17106 (N_17106,N_14699,N_11890);
nor U17107 (N_17107,N_13599,N_14371);
nor U17108 (N_17108,N_12893,N_11436);
and U17109 (N_17109,N_10696,N_11346);
nor U17110 (N_17110,N_13020,N_13042);
or U17111 (N_17111,N_13746,N_13833);
or U17112 (N_17112,N_10105,N_12073);
nor U17113 (N_17113,N_13539,N_13878);
nor U17114 (N_17114,N_12977,N_13801);
or U17115 (N_17115,N_10660,N_11341);
and U17116 (N_17116,N_13473,N_12565);
and U17117 (N_17117,N_11000,N_12183);
nor U17118 (N_17118,N_11083,N_12353);
nand U17119 (N_17119,N_14933,N_13210);
nand U17120 (N_17120,N_10950,N_14186);
and U17121 (N_17121,N_14384,N_12836);
or U17122 (N_17122,N_10567,N_14242);
nand U17123 (N_17123,N_11036,N_10850);
and U17124 (N_17124,N_13487,N_13779);
nand U17125 (N_17125,N_13044,N_10876);
nand U17126 (N_17126,N_14094,N_11451);
nor U17127 (N_17127,N_13809,N_13341);
nor U17128 (N_17128,N_13739,N_12626);
nand U17129 (N_17129,N_11628,N_11382);
nor U17130 (N_17130,N_13622,N_13807);
or U17131 (N_17131,N_11484,N_11333);
and U17132 (N_17132,N_11242,N_11487);
nor U17133 (N_17133,N_12606,N_14642);
or U17134 (N_17134,N_14325,N_13289);
nand U17135 (N_17135,N_11559,N_13708);
nor U17136 (N_17136,N_13580,N_13229);
nand U17137 (N_17137,N_10434,N_12471);
or U17138 (N_17138,N_14364,N_12370);
nor U17139 (N_17139,N_10853,N_10915);
or U17140 (N_17140,N_14404,N_14073);
nand U17141 (N_17141,N_12501,N_11598);
nand U17142 (N_17142,N_13066,N_13462);
and U17143 (N_17143,N_12413,N_12125);
or U17144 (N_17144,N_10039,N_10316);
nor U17145 (N_17145,N_13400,N_14646);
nor U17146 (N_17146,N_11981,N_12804);
or U17147 (N_17147,N_12439,N_12855);
nand U17148 (N_17148,N_13693,N_14491);
nand U17149 (N_17149,N_12478,N_13428);
nand U17150 (N_17150,N_14045,N_11396);
and U17151 (N_17151,N_12806,N_12583);
and U17152 (N_17152,N_14084,N_12290);
nor U17153 (N_17153,N_12467,N_10420);
nor U17154 (N_17154,N_10945,N_12156);
or U17155 (N_17155,N_12488,N_14047);
or U17156 (N_17156,N_13682,N_13572);
and U17157 (N_17157,N_10763,N_11147);
and U17158 (N_17158,N_13050,N_12276);
nand U17159 (N_17159,N_14488,N_13606);
nor U17160 (N_17160,N_13394,N_13880);
nor U17161 (N_17161,N_14561,N_12318);
nor U17162 (N_17162,N_14782,N_14717);
nor U17163 (N_17163,N_12532,N_13806);
nand U17164 (N_17164,N_14970,N_12151);
nor U17165 (N_17165,N_14288,N_11313);
nand U17166 (N_17166,N_12671,N_14137);
and U17167 (N_17167,N_12520,N_11105);
nand U17168 (N_17168,N_11099,N_10895);
and U17169 (N_17169,N_10894,N_12618);
nor U17170 (N_17170,N_10366,N_10621);
nand U17171 (N_17171,N_12716,N_11608);
and U17172 (N_17172,N_12084,N_11028);
or U17173 (N_17173,N_14352,N_11590);
xnor U17174 (N_17174,N_11180,N_10202);
xnor U17175 (N_17175,N_12517,N_13014);
and U17176 (N_17176,N_12548,N_13129);
nor U17177 (N_17177,N_13207,N_11759);
nand U17178 (N_17178,N_13203,N_10077);
nor U17179 (N_17179,N_12753,N_12331);
and U17180 (N_17180,N_13243,N_13493);
or U17181 (N_17181,N_10267,N_14930);
nor U17182 (N_17182,N_14401,N_14420);
nor U17183 (N_17183,N_12044,N_10645);
nand U17184 (N_17184,N_12537,N_10864);
nand U17185 (N_17185,N_10092,N_14724);
nor U17186 (N_17186,N_10509,N_10709);
or U17187 (N_17187,N_14624,N_11295);
nand U17188 (N_17188,N_14129,N_10816);
nor U17189 (N_17189,N_14360,N_14581);
xnor U17190 (N_17190,N_12708,N_12258);
nor U17191 (N_17191,N_10681,N_13459);
nor U17192 (N_17192,N_13153,N_11957);
nand U17193 (N_17193,N_12039,N_12593);
nor U17194 (N_17194,N_11633,N_14552);
or U17195 (N_17195,N_10610,N_11186);
or U17196 (N_17196,N_10836,N_14194);
and U17197 (N_17197,N_10554,N_12434);
or U17198 (N_17198,N_14076,N_10803);
nor U17199 (N_17199,N_12031,N_11278);
nand U17200 (N_17200,N_13955,N_10034);
and U17201 (N_17201,N_11508,N_11912);
nor U17202 (N_17202,N_10480,N_10629);
and U17203 (N_17203,N_14520,N_14188);
nor U17204 (N_17204,N_12916,N_14549);
nand U17205 (N_17205,N_11320,N_14789);
nor U17206 (N_17206,N_11146,N_14101);
nor U17207 (N_17207,N_14018,N_14374);
and U17208 (N_17208,N_10792,N_13131);
and U17209 (N_17209,N_13279,N_13205);
xnor U17210 (N_17210,N_14766,N_14570);
nand U17211 (N_17211,N_13040,N_11775);
nand U17212 (N_17212,N_12181,N_12035);
and U17213 (N_17213,N_12155,N_14365);
and U17214 (N_17214,N_10167,N_13605);
or U17215 (N_17215,N_13326,N_12405);
or U17216 (N_17216,N_11435,N_10978);
nand U17217 (N_17217,N_14653,N_12964);
and U17218 (N_17218,N_10017,N_11865);
and U17219 (N_17219,N_14454,N_11423);
and U17220 (N_17220,N_11670,N_14680);
and U17221 (N_17221,N_10362,N_10241);
nand U17222 (N_17222,N_10404,N_10104);
and U17223 (N_17223,N_11281,N_10968);
nor U17224 (N_17224,N_13576,N_12854);
or U17225 (N_17225,N_12141,N_14702);
nor U17226 (N_17226,N_10384,N_11530);
or U17227 (N_17227,N_14323,N_14669);
nor U17228 (N_17228,N_10793,N_11550);
and U17229 (N_17229,N_10128,N_14983);
nor U17230 (N_17230,N_10373,N_14781);
or U17231 (N_17231,N_12976,N_13583);
xor U17232 (N_17232,N_14236,N_14466);
nand U17233 (N_17233,N_14706,N_12957);
and U17234 (N_17234,N_12458,N_14144);
and U17235 (N_17235,N_14425,N_12509);
xnor U17236 (N_17236,N_11610,N_12420);
nor U17237 (N_17237,N_10001,N_11814);
xnor U17238 (N_17238,N_14042,N_13147);
and U17239 (N_17239,N_13762,N_14667);
and U17240 (N_17240,N_12680,N_12579);
nor U17241 (N_17241,N_12038,N_14477);
nor U17242 (N_17242,N_12777,N_13961);
or U17243 (N_17243,N_14160,N_13447);
nand U17244 (N_17244,N_12097,N_13839);
nor U17245 (N_17245,N_13533,N_14908);
or U17246 (N_17246,N_11114,N_12145);
nor U17247 (N_17247,N_13365,N_13983);
nor U17248 (N_17248,N_13182,N_10410);
nor U17249 (N_17249,N_10357,N_10908);
nand U17250 (N_17250,N_10882,N_10569);
and U17251 (N_17251,N_11445,N_10700);
and U17252 (N_17252,N_10544,N_11277);
or U17253 (N_17253,N_11654,N_11879);
xor U17254 (N_17254,N_11387,N_10988);
and U17255 (N_17255,N_13966,N_10058);
and U17256 (N_17256,N_10769,N_13989);
nand U17257 (N_17257,N_11013,N_13803);
and U17258 (N_17258,N_10358,N_14859);
nand U17259 (N_17259,N_10213,N_11474);
nand U17260 (N_17260,N_11620,N_11002);
nand U17261 (N_17261,N_13492,N_14666);
and U17262 (N_17262,N_12224,N_14107);
nor U17263 (N_17263,N_10121,N_14900);
or U17264 (N_17264,N_10880,N_13759);
nand U17265 (N_17265,N_13749,N_14696);
nand U17266 (N_17266,N_14924,N_11229);
nand U17267 (N_17267,N_11587,N_14210);
nor U17268 (N_17268,N_11725,N_13286);
nand U17269 (N_17269,N_12460,N_11710);
nor U17270 (N_17270,N_13980,N_12712);
nand U17271 (N_17271,N_12811,N_12749);
nand U17272 (N_17272,N_10343,N_10284);
or U17273 (N_17273,N_12556,N_10163);
nand U17274 (N_17274,N_11691,N_11236);
nor U17275 (N_17275,N_12229,N_10833);
and U17276 (N_17276,N_12432,N_12072);
nor U17277 (N_17277,N_13625,N_13509);
nand U17278 (N_17278,N_10607,N_10985);
and U17279 (N_17279,N_13160,N_14507);
nand U17280 (N_17280,N_10310,N_11187);
nor U17281 (N_17281,N_14055,N_13194);
and U17282 (N_17282,N_10253,N_10658);
and U17283 (N_17283,N_14981,N_12048);
nand U17284 (N_17284,N_10354,N_12605);
or U17285 (N_17285,N_10713,N_14206);
and U17286 (N_17286,N_14729,N_13581);
nand U17287 (N_17287,N_12284,N_14139);
nor U17288 (N_17288,N_12287,N_14223);
or U17289 (N_17289,N_12842,N_12631);
nand U17290 (N_17290,N_10221,N_12217);
nand U17291 (N_17291,N_12227,N_13982);
or U17292 (N_17292,N_14891,N_10626);
and U17293 (N_17293,N_10960,N_13507);
or U17294 (N_17294,N_13683,N_10575);
nor U17295 (N_17295,N_14664,N_11719);
or U17296 (N_17296,N_12091,N_11007);
nand U17297 (N_17297,N_13280,N_11693);
and U17298 (N_17298,N_12005,N_14613);
nor U17299 (N_17299,N_10910,N_14780);
and U17300 (N_17300,N_14254,N_13517);
nand U17301 (N_17301,N_11342,N_13755);
or U17302 (N_17302,N_14247,N_13426);
or U17303 (N_17303,N_12111,N_13658);
and U17304 (N_17304,N_11943,N_13238);
nand U17305 (N_17305,N_13556,N_13360);
or U17306 (N_17306,N_10304,N_10047);
and U17307 (N_17307,N_14411,N_14071);
nor U17308 (N_17308,N_13812,N_11001);
and U17309 (N_17309,N_11024,N_10856);
and U17310 (N_17310,N_12931,N_11254);
or U17311 (N_17311,N_12533,N_10164);
and U17312 (N_17312,N_10242,N_10236);
or U17313 (N_17313,N_14725,N_12383);
or U17314 (N_17314,N_13081,N_11032);
or U17315 (N_17315,N_11589,N_10639);
and U17316 (N_17316,N_12378,N_11144);
and U17317 (N_17317,N_14424,N_12627);
nor U17318 (N_17318,N_10157,N_14256);
and U17319 (N_17319,N_12549,N_14334);
and U17320 (N_17320,N_12757,N_14538);
and U17321 (N_17321,N_11622,N_10748);
or U17322 (N_17322,N_12800,N_14515);
and U17323 (N_17323,N_10191,N_14751);
or U17324 (N_17324,N_11658,N_12376);
and U17325 (N_17325,N_13601,N_12479);
xnor U17326 (N_17326,N_11950,N_11793);
nor U17327 (N_17327,N_11838,N_10084);
or U17328 (N_17328,N_14154,N_13382);
nor U17329 (N_17329,N_10804,N_13155);
nor U17330 (N_17330,N_12874,N_11983);
nand U17331 (N_17331,N_13053,N_12607);
or U17332 (N_17332,N_13227,N_14127);
nand U17333 (N_17333,N_11815,N_11467);
nor U17334 (N_17334,N_12747,N_13897);
nand U17335 (N_17335,N_11791,N_14655);
and U17336 (N_17336,N_13348,N_13867);
and U17337 (N_17337,N_13453,N_13457);
and U17338 (N_17338,N_14901,N_14469);
nand U17339 (N_17339,N_11463,N_11792);
or U17340 (N_17340,N_13882,N_13644);
or U17341 (N_17341,N_12357,N_13629);
nand U17342 (N_17342,N_11750,N_10446);
or U17343 (N_17343,N_11385,N_10616);
or U17344 (N_17344,N_13029,N_13466);
and U17345 (N_17345,N_13637,N_14192);
or U17346 (N_17346,N_13248,N_10755);
nand U17347 (N_17347,N_12453,N_10161);
nor U17348 (N_17348,N_11862,N_12839);
nor U17349 (N_17349,N_11881,N_12169);
and U17350 (N_17350,N_13443,N_10881);
nor U17351 (N_17351,N_10845,N_14914);
and U17352 (N_17352,N_14169,N_14436);
or U17353 (N_17353,N_12052,N_13840);
and U17354 (N_17354,N_10296,N_11638);
xnor U17355 (N_17355,N_14339,N_11112);
and U17356 (N_17356,N_10245,N_11166);
nor U17357 (N_17357,N_14778,N_13510);
and U17358 (N_17358,N_10035,N_14760);
nand U17359 (N_17359,N_12362,N_11177);
nand U17360 (N_17360,N_12419,N_14852);
and U17361 (N_17361,N_13220,N_12381);
or U17362 (N_17362,N_10313,N_11448);
nand U17363 (N_17363,N_11325,N_10858);
and U17364 (N_17364,N_11305,N_13800);
nor U17365 (N_17365,N_13295,N_12872);
or U17366 (N_17366,N_12657,N_11510);
and U17367 (N_17367,N_12932,N_12066);
nand U17368 (N_17368,N_11941,N_10705);
or U17369 (N_17369,N_10116,N_13848);
nor U17370 (N_17370,N_12514,N_10791);
or U17371 (N_17371,N_10065,N_11797);
nand U17372 (N_17372,N_12025,N_11631);
nor U17373 (N_17373,N_11762,N_12651);
or U17374 (N_17374,N_13148,N_10432);
nor U17375 (N_17375,N_10875,N_14336);
nand U17376 (N_17376,N_12841,N_11188);
nor U17377 (N_17377,N_12379,N_12554);
or U17378 (N_17378,N_13679,N_12266);
nand U17379 (N_17379,N_12008,N_14577);
and U17380 (N_17380,N_12236,N_12995);
nand U17381 (N_17381,N_10812,N_11017);
or U17382 (N_17382,N_10024,N_12883);
or U17383 (N_17383,N_14614,N_14064);
and U17384 (N_17384,N_10906,N_12996);
or U17385 (N_17385,N_12254,N_10664);
and U17386 (N_17386,N_11197,N_13831);
and U17387 (N_17387,N_10064,N_12027);
or U17388 (N_17388,N_10724,N_12602);
and U17389 (N_17389,N_14447,N_13470);
or U17390 (N_17390,N_13864,N_11316);
xor U17391 (N_17391,N_12575,N_12343);
nand U17392 (N_17392,N_11801,N_11420);
xnor U17393 (N_17393,N_12363,N_10535);
nand U17394 (N_17394,N_12890,N_10470);
and U17395 (N_17395,N_11231,N_10000);
nor U17396 (N_17396,N_12324,N_10636);
nand U17397 (N_17397,N_12483,N_11368);
nor U17398 (N_17398,N_10559,N_10869);
and U17399 (N_17399,N_11045,N_13586);
nor U17400 (N_17400,N_11238,N_13145);
nand U17401 (N_17401,N_14398,N_12521);
nor U17402 (N_17402,N_10155,N_13627);
or U17403 (N_17403,N_11258,N_10689);
and U17404 (N_17404,N_11178,N_13410);
nand U17405 (N_17405,N_10449,N_13588);
and U17406 (N_17406,N_13060,N_13577);
and U17407 (N_17407,N_10726,N_10442);
and U17408 (N_17408,N_14656,N_13643);
or U17409 (N_17409,N_11495,N_12901);
and U17410 (N_17410,N_10586,N_13478);
nor U17411 (N_17411,N_12486,N_12570);
nand U17412 (N_17412,N_13859,N_12157);
nor U17413 (N_17413,N_13636,N_11057);
or U17414 (N_17414,N_11539,N_10941);
nor U17415 (N_17415,N_14586,N_13093);
and U17416 (N_17416,N_10596,N_14126);
xnor U17417 (N_17417,N_11723,N_11332);
or U17418 (N_17418,N_13171,N_10957);
nand U17419 (N_17419,N_14726,N_14609);
nor U17420 (N_17420,N_10452,N_12604);
or U17421 (N_17421,N_11653,N_10327);
nand U17422 (N_17422,N_14178,N_13938);
nand U17423 (N_17423,N_11129,N_10334);
nand U17424 (N_17424,N_10274,N_12154);
and U17425 (N_17425,N_11601,N_14214);
and U17426 (N_17426,N_13895,N_10712);
nor U17427 (N_17427,N_14472,N_11067);
and U17428 (N_17428,N_13157,N_11504);
nor U17429 (N_17429,N_11650,N_10430);
and U17430 (N_17430,N_11126,N_12720);
nor U17431 (N_17431,N_10898,N_14170);
nor U17432 (N_17432,N_12628,N_13760);
nand U17433 (N_17433,N_11661,N_14855);
nor U17434 (N_17434,N_12455,N_13337);
nand U17435 (N_17435,N_12923,N_13055);
nor U17436 (N_17436,N_12230,N_11987);
or U17437 (N_17437,N_13037,N_11548);
nor U17438 (N_17438,N_13522,N_14693);
nor U17439 (N_17439,N_11516,N_10874);
and U17440 (N_17440,N_14593,N_12069);
or U17441 (N_17441,N_12699,N_11726);
nand U17442 (N_17442,N_12504,N_10381);
nor U17443 (N_17443,N_14235,N_11612);
nor U17444 (N_17444,N_11192,N_13651);
nor U17445 (N_17445,N_14450,N_12620);
nand U17446 (N_17446,N_11585,N_10183);
nor U17447 (N_17447,N_14847,N_14691);
nor U17448 (N_17448,N_13378,N_11683);
or U17449 (N_17449,N_14053,N_14185);
nor U17450 (N_17450,N_13707,N_13689);
and U17451 (N_17451,N_14416,N_13271);
or U17452 (N_17452,N_12971,N_10025);
nand U17453 (N_17453,N_13814,N_13163);
or U17454 (N_17454,N_12375,N_11870);
nand U17455 (N_17455,N_12955,N_14332);
nand U17456 (N_17456,N_11261,N_10920);
nand U17457 (N_17457,N_13098,N_14733);
nor U17458 (N_17458,N_13928,N_12686);
or U17459 (N_17459,N_11527,N_12354);
and U17460 (N_17460,N_11327,N_12327);
and U17461 (N_17461,N_13216,N_12459);
nand U17462 (N_17462,N_11933,N_11460);
and U17463 (N_17463,N_14275,N_10560);
nor U17464 (N_17464,N_10355,N_13655);
nor U17465 (N_17465,N_10641,N_11746);
or U17466 (N_17466,N_12108,N_12185);
nor U17467 (N_17467,N_14849,N_12003);
nand U17468 (N_17468,N_13965,N_10283);
nor U17469 (N_17469,N_11297,N_14340);
nor U17470 (N_17470,N_12869,N_12796);
and U17471 (N_17471,N_13865,N_10246);
nand U17472 (N_17472,N_12228,N_10574);
or U17473 (N_17473,N_14995,N_14057);
or U17474 (N_17474,N_11203,N_13130);
and U17475 (N_17475,N_10588,N_13935);
nor U17476 (N_17476,N_11179,N_14391);
nand U17477 (N_17477,N_13681,N_11027);
nand U17478 (N_17478,N_14383,N_11929);
nand U17479 (N_17479,N_10056,N_13211);
or U17480 (N_17480,N_14759,N_11080);
or U17481 (N_17481,N_12715,N_11081);
and U17482 (N_17482,N_11794,N_14959);
and U17483 (N_17483,N_13565,N_14739);
nand U17484 (N_17484,N_14230,N_13526);
and U17485 (N_17485,N_12801,N_10609);
and U17486 (N_17486,N_10147,N_13030);
or U17487 (N_17487,N_10403,N_14690);
nand U17488 (N_17488,N_10438,N_12792);
nand U17489 (N_17489,N_11004,N_13892);
and U17490 (N_17490,N_14937,N_13975);
nor U17491 (N_17491,N_10041,N_11431);
nor U17492 (N_17492,N_11288,N_13671);
or U17493 (N_17493,N_11336,N_14641);
or U17494 (N_17494,N_12070,N_14310);
nor U17495 (N_17495,N_10933,N_11542);
nand U17496 (N_17496,N_12519,N_14329);
nor U17497 (N_17497,N_14544,N_12525);
or U17498 (N_17498,N_10153,N_13881);
nand U17499 (N_17499,N_14857,N_14565);
and U17500 (N_17500,N_13721,N_12896);
or U17501 (N_17501,N_14975,N_11278);
nand U17502 (N_17502,N_12332,N_12279);
or U17503 (N_17503,N_12229,N_11653);
nand U17504 (N_17504,N_14562,N_12347);
or U17505 (N_17505,N_14204,N_13966);
or U17506 (N_17506,N_13193,N_12960);
and U17507 (N_17507,N_12557,N_12224);
nor U17508 (N_17508,N_12270,N_12933);
nand U17509 (N_17509,N_11346,N_11318);
nand U17510 (N_17510,N_14594,N_11188);
and U17511 (N_17511,N_13517,N_11225);
nor U17512 (N_17512,N_10598,N_12734);
and U17513 (N_17513,N_10559,N_10501);
or U17514 (N_17514,N_14969,N_12697);
nand U17515 (N_17515,N_11784,N_11059);
or U17516 (N_17516,N_14760,N_11618);
nand U17517 (N_17517,N_14067,N_12927);
nand U17518 (N_17518,N_12020,N_12186);
nand U17519 (N_17519,N_13003,N_12153);
nand U17520 (N_17520,N_11357,N_13267);
or U17521 (N_17521,N_13277,N_10807);
nor U17522 (N_17522,N_10547,N_10792);
xnor U17523 (N_17523,N_11935,N_11124);
or U17524 (N_17524,N_14190,N_10609);
nand U17525 (N_17525,N_12212,N_14390);
or U17526 (N_17526,N_13875,N_14948);
or U17527 (N_17527,N_14709,N_10766);
or U17528 (N_17528,N_10705,N_14154);
nor U17529 (N_17529,N_13703,N_10882);
or U17530 (N_17530,N_12964,N_13893);
and U17531 (N_17531,N_14354,N_11219);
or U17532 (N_17532,N_14840,N_13229);
nand U17533 (N_17533,N_10969,N_10418);
and U17534 (N_17534,N_12839,N_12058);
xnor U17535 (N_17535,N_13394,N_11334);
nand U17536 (N_17536,N_11463,N_12423);
or U17537 (N_17537,N_10223,N_12419);
or U17538 (N_17538,N_14525,N_13890);
nand U17539 (N_17539,N_10415,N_14419);
nand U17540 (N_17540,N_10817,N_10749);
nor U17541 (N_17541,N_13489,N_14408);
nand U17542 (N_17542,N_10940,N_11514);
or U17543 (N_17543,N_11213,N_12386);
nand U17544 (N_17544,N_12773,N_14268);
nor U17545 (N_17545,N_11815,N_10563);
nor U17546 (N_17546,N_14017,N_11805);
nand U17547 (N_17547,N_13964,N_14967);
nor U17548 (N_17548,N_12703,N_11546);
nor U17549 (N_17549,N_13782,N_12405);
or U17550 (N_17550,N_12508,N_11894);
xnor U17551 (N_17551,N_11236,N_13917);
nand U17552 (N_17552,N_10691,N_12612);
and U17553 (N_17553,N_14300,N_13626);
nor U17554 (N_17554,N_11186,N_11860);
xor U17555 (N_17555,N_11369,N_12625);
nor U17556 (N_17556,N_11741,N_12480);
and U17557 (N_17557,N_11772,N_14831);
xor U17558 (N_17558,N_13197,N_10083);
or U17559 (N_17559,N_10270,N_11620);
nand U17560 (N_17560,N_14450,N_10219);
nor U17561 (N_17561,N_14721,N_12189);
and U17562 (N_17562,N_14293,N_12114);
and U17563 (N_17563,N_12478,N_12213);
nand U17564 (N_17564,N_12811,N_14881);
nor U17565 (N_17565,N_12496,N_11718);
or U17566 (N_17566,N_10830,N_12160);
nand U17567 (N_17567,N_10152,N_10316);
or U17568 (N_17568,N_14949,N_12661);
nor U17569 (N_17569,N_12305,N_13863);
or U17570 (N_17570,N_10052,N_14863);
nand U17571 (N_17571,N_10526,N_13191);
or U17572 (N_17572,N_12876,N_13258);
nand U17573 (N_17573,N_13169,N_14541);
or U17574 (N_17574,N_11584,N_14466);
and U17575 (N_17575,N_11214,N_12775);
xor U17576 (N_17576,N_11139,N_11475);
or U17577 (N_17577,N_11196,N_13069);
xor U17578 (N_17578,N_12968,N_12638);
or U17579 (N_17579,N_11506,N_11424);
or U17580 (N_17580,N_12217,N_10902);
or U17581 (N_17581,N_12226,N_13696);
or U17582 (N_17582,N_14757,N_14529);
and U17583 (N_17583,N_13891,N_12376);
and U17584 (N_17584,N_13842,N_11577);
and U17585 (N_17585,N_11114,N_14312);
nor U17586 (N_17586,N_14542,N_12022);
or U17587 (N_17587,N_14246,N_11829);
nor U17588 (N_17588,N_10539,N_13151);
nand U17589 (N_17589,N_14433,N_13838);
and U17590 (N_17590,N_12992,N_14559);
and U17591 (N_17591,N_14790,N_13179);
nand U17592 (N_17592,N_14005,N_12530);
nand U17593 (N_17593,N_10958,N_13589);
or U17594 (N_17594,N_12764,N_12978);
nor U17595 (N_17595,N_11106,N_13839);
and U17596 (N_17596,N_12095,N_13340);
nand U17597 (N_17597,N_13825,N_12239);
and U17598 (N_17598,N_13119,N_13390);
or U17599 (N_17599,N_10328,N_10845);
nand U17600 (N_17600,N_12579,N_14528);
and U17601 (N_17601,N_11981,N_13469);
and U17602 (N_17602,N_12433,N_14666);
nand U17603 (N_17603,N_10585,N_11748);
nor U17604 (N_17604,N_13499,N_11778);
nor U17605 (N_17605,N_12539,N_14157);
nor U17606 (N_17606,N_11265,N_11995);
or U17607 (N_17607,N_10453,N_11448);
and U17608 (N_17608,N_14445,N_14815);
xor U17609 (N_17609,N_11455,N_12208);
nor U17610 (N_17610,N_12421,N_12729);
and U17611 (N_17611,N_13915,N_13787);
nand U17612 (N_17612,N_11321,N_13563);
nand U17613 (N_17613,N_13831,N_14449);
nand U17614 (N_17614,N_11180,N_12734);
nand U17615 (N_17615,N_14497,N_10421);
nand U17616 (N_17616,N_13891,N_12093);
nor U17617 (N_17617,N_13905,N_10323);
or U17618 (N_17618,N_10206,N_10640);
or U17619 (N_17619,N_12678,N_14945);
nand U17620 (N_17620,N_14717,N_11252);
nand U17621 (N_17621,N_13816,N_12679);
nor U17622 (N_17622,N_14230,N_11771);
or U17623 (N_17623,N_12998,N_12250);
and U17624 (N_17624,N_14538,N_12683);
nand U17625 (N_17625,N_11127,N_12828);
or U17626 (N_17626,N_12010,N_14197);
or U17627 (N_17627,N_13046,N_10151);
xnor U17628 (N_17628,N_11648,N_14661);
nor U17629 (N_17629,N_10964,N_10779);
nand U17630 (N_17630,N_11731,N_13903);
nand U17631 (N_17631,N_14467,N_13277);
and U17632 (N_17632,N_14913,N_11545);
nor U17633 (N_17633,N_11879,N_11968);
or U17634 (N_17634,N_14367,N_10791);
nand U17635 (N_17635,N_14463,N_11442);
nor U17636 (N_17636,N_13359,N_14240);
or U17637 (N_17637,N_13805,N_12374);
nand U17638 (N_17638,N_14297,N_12412);
nor U17639 (N_17639,N_13323,N_11023);
and U17640 (N_17640,N_11076,N_10732);
and U17641 (N_17641,N_14865,N_10053);
or U17642 (N_17642,N_11298,N_13859);
xnor U17643 (N_17643,N_11585,N_13140);
nor U17644 (N_17644,N_10107,N_12296);
xnor U17645 (N_17645,N_11248,N_10397);
nand U17646 (N_17646,N_13678,N_12533);
and U17647 (N_17647,N_13723,N_14563);
and U17648 (N_17648,N_12230,N_13915);
nand U17649 (N_17649,N_11586,N_10328);
nand U17650 (N_17650,N_12563,N_11773);
xnor U17651 (N_17651,N_11915,N_13256);
and U17652 (N_17652,N_11406,N_13492);
and U17653 (N_17653,N_11221,N_14673);
nor U17654 (N_17654,N_10697,N_10864);
or U17655 (N_17655,N_13521,N_13096);
nand U17656 (N_17656,N_12915,N_11512);
nor U17657 (N_17657,N_12507,N_12878);
nor U17658 (N_17658,N_13200,N_14663);
nor U17659 (N_17659,N_10296,N_12508);
nand U17660 (N_17660,N_13551,N_13908);
or U17661 (N_17661,N_12011,N_12837);
or U17662 (N_17662,N_12857,N_10198);
xor U17663 (N_17663,N_11138,N_12713);
or U17664 (N_17664,N_14751,N_14244);
and U17665 (N_17665,N_14882,N_10604);
nor U17666 (N_17666,N_10197,N_13612);
nor U17667 (N_17667,N_14519,N_10584);
nand U17668 (N_17668,N_13416,N_11400);
and U17669 (N_17669,N_10789,N_11337);
nor U17670 (N_17670,N_12705,N_14136);
and U17671 (N_17671,N_14553,N_13046);
nand U17672 (N_17672,N_11087,N_11361);
and U17673 (N_17673,N_12917,N_10359);
and U17674 (N_17674,N_12497,N_13755);
or U17675 (N_17675,N_11843,N_12290);
nor U17676 (N_17676,N_14830,N_13381);
nor U17677 (N_17677,N_13569,N_12590);
and U17678 (N_17678,N_14295,N_11463);
nand U17679 (N_17679,N_13484,N_11624);
and U17680 (N_17680,N_12992,N_11159);
nand U17681 (N_17681,N_13773,N_11318);
or U17682 (N_17682,N_10656,N_13747);
or U17683 (N_17683,N_12934,N_12992);
and U17684 (N_17684,N_11152,N_10490);
and U17685 (N_17685,N_10622,N_11403);
or U17686 (N_17686,N_12159,N_10458);
or U17687 (N_17687,N_10054,N_11836);
nor U17688 (N_17688,N_12044,N_14304);
xnor U17689 (N_17689,N_11334,N_13903);
nor U17690 (N_17690,N_12808,N_10504);
or U17691 (N_17691,N_13252,N_11878);
or U17692 (N_17692,N_13127,N_10709);
and U17693 (N_17693,N_14685,N_10009);
nand U17694 (N_17694,N_11672,N_13013);
nor U17695 (N_17695,N_13969,N_14631);
nand U17696 (N_17696,N_13908,N_10665);
nor U17697 (N_17697,N_12049,N_10476);
nand U17698 (N_17698,N_13929,N_14102);
or U17699 (N_17699,N_13232,N_11932);
and U17700 (N_17700,N_14784,N_11970);
and U17701 (N_17701,N_12057,N_10162);
and U17702 (N_17702,N_11317,N_11138);
nand U17703 (N_17703,N_14446,N_14413);
and U17704 (N_17704,N_10800,N_14946);
nor U17705 (N_17705,N_10046,N_14804);
nor U17706 (N_17706,N_12002,N_12866);
nand U17707 (N_17707,N_14437,N_14294);
nor U17708 (N_17708,N_10439,N_12572);
nand U17709 (N_17709,N_13253,N_14227);
nor U17710 (N_17710,N_12938,N_14503);
nor U17711 (N_17711,N_12590,N_13209);
nand U17712 (N_17712,N_14513,N_12073);
nand U17713 (N_17713,N_11445,N_10872);
or U17714 (N_17714,N_14467,N_12252);
and U17715 (N_17715,N_14899,N_12177);
or U17716 (N_17716,N_12392,N_12287);
or U17717 (N_17717,N_10220,N_14650);
and U17718 (N_17718,N_12469,N_13910);
and U17719 (N_17719,N_14183,N_14282);
nand U17720 (N_17720,N_11102,N_14074);
nor U17721 (N_17721,N_12136,N_13497);
nand U17722 (N_17722,N_13032,N_12822);
nor U17723 (N_17723,N_13801,N_12455);
nor U17724 (N_17724,N_10108,N_13669);
nand U17725 (N_17725,N_14202,N_14071);
and U17726 (N_17726,N_13949,N_12496);
nand U17727 (N_17727,N_12086,N_11406);
and U17728 (N_17728,N_12799,N_14259);
and U17729 (N_17729,N_12224,N_13028);
nor U17730 (N_17730,N_11378,N_12353);
nor U17731 (N_17731,N_12463,N_14674);
and U17732 (N_17732,N_12503,N_12786);
or U17733 (N_17733,N_14857,N_11083);
nand U17734 (N_17734,N_10704,N_11477);
and U17735 (N_17735,N_13061,N_14392);
nor U17736 (N_17736,N_12004,N_11626);
xor U17737 (N_17737,N_14137,N_10897);
nand U17738 (N_17738,N_10707,N_10359);
nand U17739 (N_17739,N_11943,N_14564);
nor U17740 (N_17740,N_12309,N_12325);
nor U17741 (N_17741,N_13775,N_14059);
nor U17742 (N_17742,N_13892,N_12782);
nand U17743 (N_17743,N_13542,N_14602);
and U17744 (N_17744,N_14885,N_14633);
or U17745 (N_17745,N_11375,N_13298);
nand U17746 (N_17746,N_12387,N_11920);
or U17747 (N_17747,N_13635,N_12533);
nor U17748 (N_17748,N_11098,N_12016);
and U17749 (N_17749,N_14605,N_10431);
nor U17750 (N_17750,N_11706,N_10754);
nor U17751 (N_17751,N_13404,N_13007);
nand U17752 (N_17752,N_10008,N_10910);
nand U17753 (N_17753,N_10731,N_12796);
or U17754 (N_17754,N_13287,N_12974);
xor U17755 (N_17755,N_10377,N_13898);
and U17756 (N_17756,N_14162,N_10652);
nor U17757 (N_17757,N_11277,N_12587);
and U17758 (N_17758,N_11406,N_12758);
or U17759 (N_17759,N_13177,N_13491);
nand U17760 (N_17760,N_14562,N_14908);
or U17761 (N_17761,N_14061,N_12727);
nor U17762 (N_17762,N_12179,N_12707);
nand U17763 (N_17763,N_14171,N_12512);
nor U17764 (N_17764,N_14738,N_14474);
and U17765 (N_17765,N_11734,N_12527);
and U17766 (N_17766,N_13755,N_14297);
or U17767 (N_17767,N_12871,N_11396);
nand U17768 (N_17768,N_14499,N_14564);
or U17769 (N_17769,N_11383,N_13163);
nand U17770 (N_17770,N_11095,N_14879);
or U17771 (N_17771,N_11176,N_12930);
or U17772 (N_17772,N_12415,N_11219);
nor U17773 (N_17773,N_12157,N_14192);
nor U17774 (N_17774,N_11771,N_10842);
nor U17775 (N_17775,N_11240,N_10051);
nand U17776 (N_17776,N_11734,N_11278);
nand U17777 (N_17777,N_14176,N_14083);
and U17778 (N_17778,N_13452,N_11468);
nand U17779 (N_17779,N_12275,N_12429);
nor U17780 (N_17780,N_13917,N_11192);
nand U17781 (N_17781,N_14624,N_11080);
or U17782 (N_17782,N_11402,N_10394);
nor U17783 (N_17783,N_12654,N_10516);
or U17784 (N_17784,N_10120,N_14758);
nand U17785 (N_17785,N_12459,N_11024);
and U17786 (N_17786,N_13615,N_14601);
or U17787 (N_17787,N_10833,N_12525);
nor U17788 (N_17788,N_11027,N_13162);
or U17789 (N_17789,N_12079,N_12766);
nand U17790 (N_17790,N_14745,N_12544);
or U17791 (N_17791,N_12921,N_12265);
xnor U17792 (N_17792,N_12269,N_10864);
nand U17793 (N_17793,N_11638,N_10791);
nand U17794 (N_17794,N_13248,N_11563);
nand U17795 (N_17795,N_10708,N_13097);
or U17796 (N_17796,N_11073,N_10351);
nor U17797 (N_17797,N_14627,N_12215);
or U17798 (N_17798,N_13498,N_11191);
or U17799 (N_17799,N_12921,N_13988);
and U17800 (N_17800,N_12028,N_12711);
nor U17801 (N_17801,N_10104,N_10542);
or U17802 (N_17802,N_12521,N_13995);
and U17803 (N_17803,N_13525,N_14206);
and U17804 (N_17804,N_14960,N_13618);
nor U17805 (N_17805,N_10155,N_12871);
or U17806 (N_17806,N_14854,N_10457);
or U17807 (N_17807,N_11112,N_11027);
nor U17808 (N_17808,N_12311,N_13232);
nor U17809 (N_17809,N_14132,N_10519);
nand U17810 (N_17810,N_14651,N_10797);
and U17811 (N_17811,N_12306,N_14640);
nor U17812 (N_17812,N_14429,N_14510);
nand U17813 (N_17813,N_12399,N_11822);
or U17814 (N_17814,N_13751,N_13270);
nand U17815 (N_17815,N_11560,N_11680);
xnor U17816 (N_17816,N_14753,N_13826);
nor U17817 (N_17817,N_10576,N_13845);
or U17818 (N_17818,N_13280,N_11005);
nand U17819 (N_17819,N_12370,N_12597);
nor U17820 (N_17820,N_10418,N_11383);
nor U17821 (N_17821,N_11906,N_14730);
or U17822 (N_17822,N_14247,N_11924);
nand U17823 (N_17823,N_14636,N_12217);
and U17824 (N_17824,N_11063,N_13610);
or U17825 (N_17825,N_10574,N_11643);
nor U17826 (N_17826,N_13525,N_13487);
and U17827 (N_17827,N_10365,N_14313);
or U17828 (N_17828,N_10420,N_13177);
nor U17829 (N_17829,N_13103,N_13778);
nand U17830 (N_17830,N_10031,N_14255);
or U17831 (N_17831,N_14048,N_11718);
or U17832 (N_17832,N_13281,N_14431);
nand U17833 (N_17833,N_14122,N_12227);
nor U17834 (N_17834,N_10097,N_14726);
nand U17835 (N_17835,N_11427,N_14620);
nor U17836 (N_17836,N_13010,N_10530);
or U17837 (N_17837,N_10056,N_14756);
nor U17838 (N_17838,N_10522,N_11624);
and U17839 (N_17839,N_12778,N_12126);
and U17840 (N_17840,N_12259,N_12620);
nor U17841 (N_17841,N_13934,N_10228);
and U17842 (N_17842,N_13974,N_10017);
nand U17843 (N_17843,N_13389,N_12336);
nor U17844 (N_17844,N_11794,N_12852);
nor U17845 (N_17845,N_11401,N_12923);
and U17846 (N_17846,N_13186,N_10939);
nand U17847 (N_17847,N_11457,N_12794);
nor U17848 (N_17848,N_14667,N_14956);
and U17849 (N_17849,N_12195,N_14997);
nor U17850 (N_17850,N_11871,N_13315);
nand U17851 (N_17851,N_11310,N_11195);
and U17852 (N_17852,N_11982,N_13242);
or U17853 (N_17853,N_14118,N_11839);
and U17854 (N_17854,N_13717,N_10368);
and U17855 (N_17855,N_12872,N_11540);
nor U17856 (N_17856,N_11119,N_10048);
nand U17857 (N_17857,N_10606,N_10907);
and U17858 (N_17858,N_14701,N_12368);
and U17859 (N_17859,N_13166,N_13791);
nand U17860 (N_17860,N_14206,N_10794);
nand U17861 (N_17861,N_12962,N_10456);
nor U17862 (N_17862,N_12259,N_12297);
and U17863 (N_17863,N_11164,N_14853);
nand U17864 (N_17864,N_10839,N_11894);
and U17865 (N_17865,N_13166,N_12612);
and U17866 (N_17866,N_12753,N_14772);
or U17867 (N_17867,N_10300,N_13800);
or U17868 (N_17868,N_12055,N_13268);
and U17869 (N_17869,N_14187,N_12876);
nor U17870 (N_17870,N_10556,N_14374);
nor U17871 (N_17871,N_10535,N_13314);
or U17872 (N_17872,N_10369,N_13855);
nand U17873 (N_17873,N_13602,N_14059);
and U17874 (N_17874,N_12259,N_13933);
and U17875 (N_17875,N_13240,N_13159);
or U17876 (N_17876,N_13550,N_12865);
nand U17877 (N_17877,N_10329,N_10314);
or U17878 (N_17878,N_13006,N_13129);
or U17879 (N_17879,N_11653,N_11019);
nor U17880 (N_17880,N_13861,N_13657);
and U17881 (N_17881,N_13643,N_13903);
nor U17882 (N_17882,N_12635,N_14346);
or U17883 (N_17883,N_14465,N_12908);
nor U17884 (N_17884,N_13406,N_10523);
and U17885 (N_17885,N_14683,N_14288);
nor U17886 (N_17886,N_14061,N_11450);
and U17887 (N_17887,N_14867,N_11696);
and U17888 (N_17888,N_13928,N_13336);
nand U17889 (N_17889,N_12075,N_13084);
nor U17890 (N_17890,N_10183,N_10126);
nand U17891 (N_17891,N_12553,N_10209);
nand U17892 (N_17892,N_13280,N_10320);
or U17893 (N_17893,N_13620,N_10382);
or U17894 (N_17894,N_13277,N_14422);
or U17895 (N_17895,N_10597,N_11399);
and U17896 (N_17896,N_14379,N_12386);
nor U17897 (N_17897,N_11529,N_10777);
nand U17898 (N_17898,N_14742,N_11008);
and U17899 (N_17899,N_10271,N_13310);
nand U17900 (N_17900,N_14232,N_14114);
nand U17901 (N_17901,N_10181,N_12751);
nor U17902 (N_17902,N_11773,N_10101);
or U17903 (N_17903,N_11580,N_13010);
or U17904 (N_17904,N_14095,N_10815);
or U17905 (N_17905,N_13696,N_14864);
or U17906 (N_17906,N_12132,N_11327);
xnor U17907 (N_17907,N_10999,N_11771);
nand U17908 (N_17908,N_11560,N_14463);
and U17909 (N_17909,N_14892,N_14079);
nand U17910 (N_17910,N_12827,N_14183);
or U17911 (N_17911,N_11989,N_11503);
and U17912 (N_17912,N_13046,N_14119);
and U17913 (N_17913,N_14050,N_13355);
and U17914 (N_17914,N_13684,N_12961);
or U17915 (N_17915,N_10125,N_11235);
or U17916 (N_17916,N_10302,N_12306);
nand U17917 (N_17917,N_10592,N_13572);
nor U17918 (N_17918,N_12946,N_11280);
nor U17919 (N_17919,N_14789,N_11067);
nand U17920 (N_17920,N_10293,N_12726);
nor U17921 (N_17921,N_13409,N_12482);
and U17922 (N_17922,N_12302,N_12058);
or U17923 (N_17923,N_13603,N_13061);
nor U17924 (N_17924,N_11226,N_14339);
xor U17925 (N_17925,N_11278,N_12215);
and U17926 (N_17926,N_13451,N_12540);
and U17927 (N_17927,N_12973,N_13921);
nand U17928 (N_17928,N_11355,N_14102);
nor U17929 (N_17929,N_10381,N_10979);
and U17930 (N_17930,N_10215,N_14002);
nor U17931 (N_17931,N_13166,N_14524);
nand U17932 (N_17932,N_13873,N_14503);
nand U17933 (N_17933,N_13834,N_12935);
or U17934 (N_17934,N_14595,N_12249);
xnor U17935 (N_17935,N_13241,N_12562);
nor U17936 (N_17936,N_12376,N_10526);
and U17937 (N_17937,N_14972,N_13189);
and U17938 (N_17938,N_14569,N_13556);
nand U17939 (N_17939,N_11369,N_13049);
or U17940 (N_17940,N_10216,N_10109);
nand U17941 (N_17941,N_14212,N_12332);
nor U17942 (N_17942,N_13474,N_11941);
and U17943 (N_17943,N_11575,N_13403);
nand U17944 (N_17944,N_12083,N_10562);
xnor U17945 (N_17945,N_12804,N_14331);
nand U17946 (N_17946,N_12833,N_12487);
or U17947 (N_17947,N_12644,N_12388);
and U17948 (N_17948,N_13228,N_10713);
or U17949 (N_17949,N_11678,N_10046);
nand U17950 (N_17950,N_12696,N_13986);
or U17951 (N_17951,N_10035,N_12765);
and U17952 (N_17952,N_12557,N_14525);
or U17953 (N_17953,N_10901,N_11203);
or U17954 (N_17954,N_13297,N_14714);
or U17955 (N_17955,N_12020,N_14197);
and U17956 (N_17956,N_12144,N_10306);
or U17957 (N_17957,N_14232,N_10336);
nand U17958 (N_17958,N_13317,N_12497);
or U17959 (N_17959,N_11630,N_12003);
nor U17960 (N_17960,N_14351,N_11650);
and U17961 (N_17961,N_12391,N_11796);
nor U17962 (N_17962,N_12408,N_11344);
nand U17963 (N_17963,N_13815,N_11418);
xor U17964 (N_17964,N_10415,N_12152);
xor U17965 (N_17965,N_14164,N_11882);
and U17966 (N_17966,N_12666,N_10480);
nand U17967 (N_17967,N_11527,N_12552);
and U17968 (N_17968,N_13984,N_10775);
nand U17969 (N_17969,N_14432,N_14939);
or U17970 (N_17970,N_13595,N_13968);
and U17971 (N_17971,N_10759,N_13985);
nand U17972 (N_17972,N_11587,N_11940);
nand U17973 (N_17973,N_10693,N_12087);
nor U17974 (N_17974,N_12795,N_12953);
or U17975 (N_17975,N_14242,N_14785);
or U17976 (N_17976,N_12265,N_12382);
nand U17977 (N_17977,N_14115,N_13198);
nand U17978 (N_17978,N_12192,N_10772);
nand U17979 (N_17979,N_14047,N_11947);
nor U17980 (N_17980,N_14650,N_13553);
or U17981 (N_17981,N_13916,N_14619);
and U17982 (N_17982,N_11833,N_12160);
nand U17983 (N_17983,N_11571,N_10218);
nand U17984 (N_17984,N_14977,N_11839);
or U17985 (N_17985,N_10626,N_14383);
nand U17986 (N_17986,N_12430,N_14300);
nand U17987 (N_17987,N_10402,N_14885);
or U17988 (N_17988,N_12212,N_13741);
or U17989 (N_17989,N_11372,N_11709);
or U17990 (N_17990,N_10234,N_12456);
nor U17991 (N_17991,N_14205,N_10473);
and U17992 (N_17992,N_11859,N_13106);
or U17993 (N_17993,N_14553,N_12554);
nor U17994 (N_17994,N_14190,N_13951);
and U17995 (N_17995,N_10371,N_13683);
nand U17996 (N_17996,N_14031,N_11717);
or U17997 (N_17997,N_13254,N_12428);
nand U17998 (N_17998,N_13313,N_11208);
and U17999 (N_17999,N_11793,N_13336);
and U18000 (N_18000,N_11507,N_12750);
nor U18001 (N_18001,N_13812,N_10549);
or U18002 (N_18002,N_12815,N_14214);
nor U18003 (N_18003,N_13897,N_14204);
nand U18004 (N_18004,N_10495,N_11422);
or U18005 (N_18005,N_13007,N_11366);
nor U18006 (N_18006,N_11668,N_14607);
nor U18007 (N_18007,N_12920,N_11927);
nor U18008 (N_18008,N_12789,N_14563);
nor U18009 (N_18009,N_12637,N_14941);
nand U18010 (N_18010,N_13813,N_11762);
nor U18011 (N_18011,N_12142,N_11532);
or U18012 (N_18012,N_14969,N_10366);
xnor U18013 (N_18013,N_12484,N_13141);
and U18014 (N_18014,N_13735,N_10851);
nor U18015 (N_18015,N_13486,N_13299);
and U18016 (N_18016,N_13842,N_12278);
or U18017 (N_18017,N_10217,N_13616);
nor U18018 (N_18018,N_14072,N_10884);
nor U18019 (N_18019,N_11085,N_12044);
or U18020 (N_18020,N_13798,N_11444);
and U18021 (N_18021,N_10853,N_14445);
nand U18022 (N_18022,N_10960,N_10443);
nand U18023 (N_18023,N_13363,N_10579);
and U18024 (N_18024,N_12339,N_13482);
nor U18025 (N_18025,N_11369,N_13372);
nor U18026 (N_18026,N_13798,N_12762);
and U18027 (N_18027,N_10972,N_13128);
nor U18028 (N_18028,N_10709,N_10988);
nand U18029 (N_18029,N_11640,N_11763);
or U18030 (N_18030,N_11012,N_11522);
and U18031 (N_18031,N_13230,N_14532);
nor U18032 (N_18032,N_10481,N_11225);
nand U18033 (N_18033,N_10714,N_12763);
nand U18034 (N_18034,N_14714,N_10873);
or U18035 (N_18035,N_13079,N_10268);
xor U18036 (N_18036,N_13496,N_13186);
and U18037 (N_18037,N_10476,N_10431);
nor U18038 (N_18038,N_14829,N_10942);
and U18039 (N_18039,N_12464,N_11068);
or U18040 (N_18040,N_14550,N_14978);
xor U18041 (N_18041,N_13129,N_14565);
nand U18042 (N_18042,N_12180,N_13355);
or U18043 (N_18043,N_12816,N_14716);
nand U18044 (N_18044,N_10360,N_14268);
and U18045 (N_18045,N_10385,N_14027);
or U18046 (N_18046,N_10713,N_11256);
and U18047 (N_18047,N_14604,N_13819);
nand U18048 (N_18048,N_14641,N_13500);
nor U18049 (N_18049,N_10236,N_12298);
nor U18050 (N_18050,N_11550,N_13200);
nor U18051 (N_18051,N_13025,N_13486);
or U18052 (N_18052,N_12608,N_14109);
and U18053 (N_18053,N_11552,N_12820);
or U18054 (N_18054,N_14383,N_10282);
nor U18055 (N_18055,N_12426,N_12364);
and U18056 (N_18056,N_12216,N_12303);
or U18057 (N_18057,N_13818,N_10147);
or U18058 (N_18058,N_14381,N_13335);
nand U18059 (N_18059,N_13249,N_10971);
nand U18060 (N_18060,N_14964,N_12349);
and U18061 (N_18061,N_13738,N_12339);
nand U18062 (N_18062,N_10770,N_11489);
and U18063 (N_18063,N_10571,N_10878);
nor U18064 (N_18064,N_10145,N_12099);
or U18065 (N_18065,N_11486,N_14051);
and U18066 (N_18066,N_10658,N_14532);
and U18067 (N_18067,N_11979,N_10290);
or U18068 (N_18068,N_12335,N_11894);
and U18069 (N_18069,N_11205,N_13681);
nor U18070 (N_18070,N_14102,N_11007);
nand U18071 (N_18071,N_12028,N_14797);
and U18072 (N_18072,N_13043,N_10070);
or U18073 (N_18073,N_11330,N_12873);
nor U18074 (N_18074,N_13970,N_11095);
and U18075 (N_18075,N_13469,N_10676);
nand U18076 (N_18076,N_11331,N_11611);
nand U18077 (N_18077,N_10064,N_12880);
or U18078 (N_18078,N_11422,N_14272);
and U18079 (N_18079,N_10030,N_11772);
or U18080 (N_18080,N_14112,N_12210);
and U18081 (N_18081,N_13743,N_10907);
or U18082 (N_18082,N_13285,N_14161);
nor U18083 (N_18083,N_13928,N_10331);
or U18084 (N_18084,N_14002,N_13416);
nor U18085 (N_18085,N_10686,N_12861);
nand U18086 (N_18086,N_13358,N_14631);
nand U18087 (N_18087,N_11726,N_13251);
nand U18088 (N_18088,N_10593,N_11844);
nor U18089 (N_18089,N_11857,N_14518);
or U18090 (N_18090,N_14955,N_12784);
nand U18091 (N_18091,N_12371,N_14426);
or U18092 (N_18092,N_10077,N_14832);
nand U18093 (N_18093,N_11556,N_11928);
or U18094 (N_18094,N_10652,N_11942);
and U18095 (N_18095,N_12395,N_11494);
or U18096 (N_18096,N_14387,N_10246);
nand U18097 (N_18097,N_11801,N_10353);
nand U18098 (N_18098,N_14337,N_11097);
nand U18099 (N_18099,N_12240,N_14423);
nor U18100 (N_18100,N_13748,N_11855);
or U18101 (N_18101,N_13289,N_10382);
and U18102 (N_18102,N_13844,N_12202);
nor U18103 (N_18103,N_12321,N_10752);
nand U18104 (N_18104,N_13690,N_10308);
nor U18105 (N_18105,N_14939,N_11662);
or U18106 (N_18106,N_13868,N_12281);
nor U18107 (N_18107,N_14284,N_10183);
or U18108 (N_18108,N_12534,N_11799);
nand U18109 (N_18109,N_14949,N_11262);
or U18110 (N_18110,N_14536,N_12760);
or U18111 (N_18111,N_10696,N_10560);
nor U18112 (N_18112,N_12749,N_10878);
and U18113 (N_18113,N_14707,N_13906);
and U18114 (N_18114,N_12716,N_11992);
and U18115 (N_18115,N_10129,N_12894);
nor U18116 (N_18116,N_12387,N_12811);
and U18117 (N_18117,N_11572,N_14600);
nand U18118 (N_18118,N_10575,N_13810);
nor U18119 (N_18119,N_12292,N_12109);
nor U18120 (N_18120,N_11963,N_12273);
nand U18121 (N_18121,N_13598,N_11061);
nor U18122 (N_18122,N_11414,N_11202);
nor U18123 (N_18123,N_13867,N_12665);
nand U18124 (N_18124,N_12834,N_14796);
and U18125 (N_18125,N_11992,N_11818);
nor U18126 (N_18126,N_12715,N_10931);
nand U18127 (N_18127,N_13823,N_10081);
or U18128 (N_18128,N_10218,N_13533);
nor U18129 (N_18129,N_11889,N_12624);
nor U18130 (N_18130,N_11573,N_12962);
or U18131 (N_18131,N_10407,N_12416);
or U18132 (N_18132,N_13563,N_13971);
nand U18133 (N_18133,N_13625,N_11027);
and U18134 (N_18134,N_14232,N_10190);
and U18135 (N_18135,N_12663,N_10393);
nor U18136 (N_18136,N_10673,N_10129);
or U18137 (N_18137,N_10345,N_11501);
xor U18138 (N_18138,N_14954,N_14853);
or U18139 (N_18139,N_14595,N_10901);
or U18140 (N_18140,N_11844,N_10727);
nor U18141 (N_18141,N_13169,N_14110);
nand U18142 (N_18142,N_14464,N_14210);
or U18143 (N_18143,N_12378,N_11679);
nand U18144 (N_18144,N_14646,N_13979);
or U18145 (N_18145,N_13320,N_14322);
and U18146 (N_18146,N_11457,N_14228);
and U18147 (N_18147,N_13099,N_13941);
nand U18148 (N_18148,N_12420,N_10938);
and U18149 (N_18149,N_14427,N_11362);
and U18150 (N_18150,N_10733,N_10416);
and U18151 (N_18151,N_13322,N_12555);
nor U18152 (N_18152,N_13723,N_12228);
or U18153 (N_18153,N_10102,N_10778);
or U18154 (N_18154,N_11147,N_14853);
nand U18155 (N_18155,N_13394,N_10347);
or U18156 (N_18156,N_11135,N_14988);
or U18157 (N_18157,N_12034,N_14316);
nor U18158 (N_18158,N_12997,N_12398);
or U18159 (N_18159,N_11793,N_12550);
and U18160 (N_18160,N_10066,N_14633);
nor U18161 (N_18161,N_13072,N_11870);
xor U18162 (N_18162,N_12631,N_10507);
nor U18163 (N_18163,N_10493,N_13736);
or U18164 (N_18164,N_13112,N_14033);
and U18165 (N_18165,N_11042,N_14108);
and U18166 (N_18166,N_12298,N_12102);
nand U18167 (N_18167,N_12551,N_14673);
and U18168 (N_18168,N_11569,N_14844);
or U18169 (N_18169,N_10846,N_12372);
or U18170 (N_18170,N_13345,N_10975);
nor U18171 (N_18171,N_13242,N_13933);
and U18172 (N_18172,N_11397,N_12366);
and U18173 (N_18173,N_14499,N_12062);
and U18174 (N_18174,N_11190,N_11711);
or U18175 (N_18175,N_14410,N_10976);
xnor U18176 (N_18176,N_10378,N_14529);
nor U18177 (N_18177,N_11098,N_11511);
or U18178 (N_18178,N_14706,N_12037);
nor U18179 (N_18179,N_13236,N_14187);
and U18180 (N_18180,N_14170,N_14735);
nor U18181 (N_18181,N_12256,N_10755);
and U18182 (N_18182,N_10412,N_11990);
or U18183 (N_18183,N_13617,N_14913);
and U18184 (N_18184,N_13900,N_13509);
and U18185 (N_18185,N_10608,N_11736);
nor U18186 (N_18186,N_14285,N_11107);
and U18187 (N_18187,N_11511,N_11365);
or U18188 (N_18188,N_10516,N_12913);
nand U18189 (N_18189,N_13007,N_13996);
or U18190 (N_18190,N_10581,N_14393);
or U18191 (N_18191,N_11572,N_11522);
and U18192 (N_18192,N_11720,N_14849);
and U18193 (N_18193,N_10905,N_10634);
nand U18194 (N_18194,N_12303,N_14478);
and U18195 (N_18195,N_12607,N_10936);
and U18196 (N_18196,N_10985,N_13637);
and U18197 (N_18197,N_13965,N_10079);
or U18198 (N_18198,N_10574,N_10293);
or U18199 (N_18199,N_14197,N_10123);
and U18200 (N_18200,N_10466,N_13671);
nand U18201 (N_18201,N_14472,N_10028);
and U18202 (N_18202,N_12022,N_10420);
and U18203 (N_18203,N_11283,N_10542);
nor U18204 (N_18204,N_11478,N_10417);
xor U18205 (N_18205,N_14855,N_11020);
nor U18206 (N_18206,N_10001,N_14409);
nand U18207 (N_18207,N_10833,N_14864);
nor U18208 (N_18208,N_11117,N_13508);
or U18209 (N_18209,N_14857,N_10886);
nand U18210 (N_18210,N_14790,N_14436);
nor U18211 (N_18211,N_11851,N_11769);
or U18212 (N_18212,N_10498,N_11256);
nand U18213 (N_18213,N_14403,N_10099);
xnor U18214 (N_18214,N_10703,N_10237);
or U18215 (N_18215,N_10789,N_14692);
nand U18216 (N_18216,N_11516,N_11217);
nand U18217 (N_18217,N_11824,N_12005);
or U18218 (N_18218,N_12221,N_10856);
nor U18219 (N_18219,N_12085,N_11441);
nor U18220 (N_18220,N_12653,N_11128);
and U18221 (N_18221,N_12916,N_10732);
nand U18222 (N_18222,N_13446,N_12752);
and U18223 (N_18223,N_13710,N_12777);
nor U18224 (N_18224,N_11358,N_10943);
and U18225 (N_18225,N_13423,N_10317);
or U18226 (N_18226,N_12489,N_11835);
or U18227 (N_18227,N_10681,N_12293);
nand U18228 (N_18228,N_11194,N_10844);
nand U18229 (N_18229,N_14037,N_10404);
nor U18230 (N_18230,N_10152,N_12763);
nor U18231 (N_18231,N_13060,N_13598);
or U18232 (N_18232,N_12575,N_13694);
nor U18233 (N_18233,N_12419,N_10062);
or U18234 (N_18234,N_11322,N_14097);
or U18235 (N_18235,N_14931,N_11313);
nor U18236 (N_18236,N_13129,N_12530);
or U18237 (N_18237,N_10345,N_13917);
nand U18238 (N_18238,N_12766,N_14402);
and U18239 (N_18239,N_11535,N_10990);
and U18240 (N_18240,N_11501,N_13810);
xor U18241 (N_18241,N_13207,N_13235);
nand U18242 (N_18242,N_10415,N_12084);
and U18243 (N_18243,N_14080,N_11480);
nor U18244 (N_18244,N_11813,N_13158);
and U18245 (N_18245,N_13622,N_10470);
or U18246 (N_18246,N_10835,N_14501);
nor U18247 (N_18247,N_12724,N_13610);
and U18248 (N_18248,N_13922,N_14319);
nand U18249 (N_18249,N_12880,N_14326);
or U18250 (N_18250,N_12857,N_14432);
and U18251 (N_18251,N_11119,N_13766);
nand U18252 (N_18252,N_14593,N_10935);
and U18253 (N_18253,N_10720,N_12109);
xor U18254 (N_18254,N_14319,N_10427);
and U18255 (N_18255,N_14024,N_12372);
and U18256 (N_18256,N_10237,N_10784);
nor U18257 (N_18257,N_12522,N_14425);
nand U18258 (N_18258,N_12003,N_10188);
or U18259 (N_18259,N_11674,N_11633);
or U18260 (N_18260,N_14444,N_14945);
and U18261 (N_18261,N_12019,N_11694);
nand U18262 (N_18262,N_14338,N_11094);
xnor U18263 (N_18263,N_12804,N_13191);
nand U18264 (N_18264,N_11183,N_10441);
nor U18265 (N_18265,N_13462,N_10856);
and U18266 (N_18266,N_13929,N_11707);
nor U18267 (N_18267,N_14159,N_14937);
or U18268 (N_18268,N_14894,N_14486);
and U18269 (N_18269,N_14481,N_13990);
and U18270 (N_18270,N_11507,N_11833);
nor U18271 (N_18271,N_11581,N_13395);
nand U18272 (N_18272,N_12461,N_11351);
nor U18273 (N_18273,N_13153,N_11804);
nand U18274 (N_18274,N_14773,N_13387);
or U18275 (N_18275,N_10178,N_11180);
nor U18276 (N_18276,N_13071,N_11742);
or U18277 (N_18277,N_12236,N_13329);
or U18278 (N_18278,N_14602,N_12516);
or U18279 (N_18279,N_10377,N_11720);
nor U18280 (N_18280,N_11498,N_11278);
nand U18281 (N_18281,N_14374,N_11497);
and U18282 (N_18282,N_10155,N_14908);
nand U18283 (N_18283,N_11724,N_11308);
nand U18284 (N_18284,N_14771,N_10222);
nand U18285 (N_18285,N_10192,N_12396);
nand U18286 (N_18286,N_11334,N_13206);
nor U18287 (N_18287,N_13716,N_13089);
and U18288 (N_18288,N_11140,N_12311);
nand U18289 (N_18289,N_13241,N_11848);
and U18290 (N_18290,N_11734,N_13874);
nand U18291 (N_18291,N_13014,N_14061);
and U18292 (N_18292,N_10097,N_10648);
nand U18293 (N_18293,N_14666,N_11861);
or U18294 (N_18294,N_11716,N_10672);
nor U18295 (N_18295,N_14713,N_10442);
nor U18296 (N_18296,N_11970,N_13448);
xor U18297 (N_18297,N_12521,N_13143);
and U18298 (N_18298,N_11988,N_10988);
nand U18299 (N_18299,N_10003,N_13944);
nand U18300 (N_18300,N_12826,N_12347);
nor U18301 (N_18301,N_12845,N_13484);
or U18302 (N_18302,N_11629,N_12684);
xnor U18303 (N_18303,N_10202,N_14166);
or U18304 (N_18304,N_14286,N_11379);
or U18305 (N_18305,N_11130,N_12057);
or U18306 (N_18306,N_12454,N_10226);
nor U18307 (N_18307,N_12912,N_13329);
nand U18308 (N_18308,N_13981,N_14386);
or U18309 (N_18309,N_10572,N_12465);
and U18310 (N_18310,N_13997,N_10421);
or U18311 (N_18311,N_10422,N_12880);
nor U18312 (N_18312,N_13248,N_13877);
nand U18313 (N_18313,N_10664,N_10735);
nor U18314 (N_18314,N_12855,N_12402);
or U18315 (N_18315,N_11620,N_11289);
nor U18316 (N_18316,N_14194,N_12875);
nor U18317 (N_18317,N_12226,N_13975);
nand U18318 (N_18318,N_11930,N_13147);
nor U18319 (N_18319,N_10316,N_13438);
nand U18320 (N_18320,N_14526,N_11952);
or U18321 (N_18321,N_14121,N_13565);
or U18322 (N_18322,N_12087,N_13133);
nor U18323 (N_18323,N_12948,N_10493);
nor U18324 (N_18324,N_10899,N_10996);
and U18325 (N_18325,N_12508,N_12251);
nand U18326 (N_18326,N_13044,N_12625);
and U18327 (N_18327,N_14535,N_14942);
nor U18328 (N_18328,N_12304,N_14990);
nand U18329 (N_18329,N_11702,N_12328);
or U18330 (N_18330,N_14840,N_13911);
nand U18331 (N_18331,N_14859,N_14648);
and U18332 (N_18332,N_11749,N_11082);
nand U18333 (N_18333,N_14102,N_12590);
nor U18334 (N_18334,N_13575,N_10280);
or U18335 (N_18335,N_14608,N_12494);
xor U18336 (N_18336,N_14852,N_10917);
nor U18337 (N_18337,N_11219,N_13090);
or U18338 (N_18338,N_12474,N_12182);
nand U18339 (N_18339,N_11252,N_12650);
or U18340 (N_18340,N_11150,N_13653);
and U18341 (N_18341,N_10122,N_10541);
nor U18342 (N_18342,N_11169,N_13677);
and U18343 (N_18343,N_14352,N_12492);
nor U18344 (N_18344,N_11501,N_14288);
and U18345 (N_18345,N_10757,N_13777);
or U18346 (N_18346,N_12035,N_14628);
or U18347 (N_18347,N_14831,N_13939);
or U18348 (N_18348,N_11220,N_11667);
xor U18349 (N_18349,N_11026,N_12522);
or U18350 (N_18350,N_10181,N_10774);
nand U18351 (N_18351,N_14013,N_12055);
nor U18352 (N_18352,N_14161,N_14282);
nor U18353 (N_18353,N_12416,N_14459);
nor U18354 (N_18354,N_12115,N_11589);
or U18355 (N_18355,N_12698,N_10118);
or U18356 (N_18356,N_11676,N_12477);
nor U18357 (N_18357,N_11581,N_12039);
nand U18358 (N_18358,N_13308,N_10883);
or U18359 (N_18359,N_10192,N_10925);
or U18360 (N_18360,N_12549,N_14782);
nor U18361 (N_18361,N_10362,N_13068);
nor U18362 (N_18362,N_13363,N_11477);
nand U18363 (N_18363,N_13925,N_10724);
and U18364 (N_18364,N_10819,N_10426);
nor U18365 (N_18365,N_14762,N_11215);
nor U18366 (N_18366,N_10689,N_11206);
nand U18367 (N_18367,N_10546,N_14633);
nand U18368 (N_18368,N_12638,N_12904);
nand U18369 (N_18369,N_12222,N_14795);
and U18370 (N_18370,N_13702,N_12340);
and U18371 (N_18371,N_14101,N_13757);
nand U18372 (N_18372,N_11711,N_11782);
and U18373 (N_18373,N_14760,N_12318);
and U18374 (N_18374,N_13725,N_14190);
nor U18375 (N_18375,N_13933,N_14312);
or U18376 (N_18376,N_12413,N_13139);
or U18377 (N_18377,N_14574,N_10869);
nand U18378 (N_18378,N_13855,N_13716);
nor U18379 (N_18379,N_14155,N_12683);
and U18380 (N_18380,N_12705,N_10617);
or U18381 (N_18381,N_13551,N_12492);
and U18382 (N_18382,N_10706,N_12010);
and U18383 (N_18383,N_11061,N_14201);
nand U18384 (N_18384,N_14158,N_14024);
and U18385 (N_18385,N_14702,N_13751);
nor U18386 (N_18386,N_14170,N_10306);
or U18387 (N_18387,N_13804,N_12928);
nor U18388 (N_18388,N_13721,N_12659);
nor U18389 (N_18389,N_12369,N_14980);
nor U18390 (N_18390,N_11961,N_11709);
nand U18391 (N_18391,N_14586,N_13121);
or U18392 (N_18392,N_14488,N_11389);
or U18393 (N_18393,N_12543,N_13781);
and U18394 (N_18394,N_14824,N_10821);
nor U18395 (N_18395,N_11310,N_12771);
nand U18396 (N_18396,N_12972,N_10789);
nor U18397 (N_18397,N_12425,N_11329);
or U18398 (N_18398,N_13279,N_10556);
nand U18399 (N_18399,N_14920,N_10191);
nand U18400 (N_18400,N_14052,N_11450);
nand U18401 (N_18401,N_14431,N_14357);
and U18402 (N_18402,N_14799,N_14889);
or U18403 (N_18403,N_12601,N_11285);
nor U18404 (N_18404,N_10550,N_12523);
and U18405 (N_18405,N_13139,N_14158);
and U18406 (N_18406,N_14193,N_12726);
and U18407 (N_18407,N_12324,N_14791);
or U18408 (N_18408,N_11910,N_13236);
and U18409 (N_18409,N_13361,N_10844);
or U18410 (N_18410,N_12039,N_12002);
nand U18411 (N_18411,N_11254,N_11325);
or U18412 (N_18412,N_14991,N_13987);
and U18413 (N_18413,N_11392,N_10446);
nand U18414 (N_18414,N_12946,N_12158);
nor U18415 (N_18415,N_13824,N_14250);
or U18416 (N_18416,N_10769,N_12640);
or U18417 (N_18417,N_14130,N_14378);
nor U18418 (N_18418,N_14327,N_10551);
nor U18419 (N_18419,N_11872,N_11247);
nand U18420 (N_18420,N_11161,N_10615);
nor U18421 (N_18421,N_14433,N_12165);
and U18422 (N_18422,N_14292,N_11472);
or U18423 (N_18423,N_12248,N_13005);
nor U18424 (N_18424,N_12084,N_11338);
nor U18425 (N_18425,N_11947,N_13086);
and U18426 (N_18426,N_12577,N_10010);
and U18427 (N_18427,N_14569,N_12218);
nor U18428 (N_18428,N_12645,N_14168);
nor U18429 (N_18429,N_13662,N_12005);
and U18430 (N_18430,N_12230,N_13071);
xor U18431 (N_18431,N_11824,N_12087);
nand U18432 (N_18432,N_11155,N_10475);
and U18433 (N_18433,N_14746,N_14166);
or U18434 (N_18434,N_10732,N_14687);
nand U18435 (N_18435,N_11171,N_10751);
nor U18436 (N_18436,N_10701,N_11936);
or U18437 (N_18437,N_11111,N_11851);
and U18438 (N_18438,N_13043,N_11950);
nand U18439 (N_18439,N_14242,N_13293);
and U18440 (N_18440,N_14267,N_11487);
nor U18441 (N_18441,N_12426,N_13528);
nand U18442 (N_18442,N_14444,N_11680);
and U18443 (N_18443,N_14042,N_14465);
or U18444 (N_18444,N_10519,N_13791);
nor U18445 (N_18445,N_10204,N_11769);
or U18446 (N_18446,N_10135,N_14164);
or U18447 (N_18447,N_13671,N_10317);
nor U18448 (N_18448,N_14411,N_12317);
and U18449 (N_18449,N_10782,N_14913);
nor U18450 (N_18450,N_10638,N_11751);
or U18451 (N_18451,N_14895,N_10575);
and U18452 (N_18452,N_13180,N_12330);
nor U18453 (N_18453,N_13313,N_12143);
nor U18454 (N_18454,N_10977,N_11453);
and U18455 (N_18455,N_12733,N_11476);
and U18456 (N_18456,N_10665,N_13891);
or U18457 (N_18457,N_13036,N_14803);
nor U18458 (N_18458,N_13096,N_14752);
and U18459 (N_18459,N_11574,N_13081);
or U18460 (N_18460,N_12335,N_14742);
and U18461 (N_18461,N_13497,N_12218);
and U18462 (N_18462,N_14981,N_10644);
and U18463 (N_18463,N_13870,N_14586);
and U18464 (N_18464,N_13113,N_13045);
nand U18465 (N_18465,N_14433,N_14458);
and U18466 (N_18466,N_14056,N_13975);
and U18467 (N_18467,N_12913,N_11800);
or U18468 (N_18468,N_11539,N_13930);
nand U18469 (N_18469,N_12435,N_14847);
nor U18470 (N_18470,N_10173,N_14713);
nor U18471 (N_18471,N_11004,N_14196);
and U18472 (N_18472,N_11250,N_14022);
and U18473 (N_18473,N_13705,N_12990);
nor U18474 (N_18474,N_13711,N_10099);
nor U18475 (N_18475,N_14418,N_12635);
nand U18476 (N_18476,N_13961,N_14905);
or U18477 (N_18477,N_11664,N_14571);
nor U18478 (N_18478,N_13074,N_11276);
and U18479 (N_18479,N_11879,N_14195);
nand U18480 (N_18480,N_13915,N_12174);
nand U18481 (N_18481,N_14368,N_14935);
or U18482 (N_18482,N_10723,N_12072);
and U18483 (N_18483,N_11648,N_13587);
nor U18484 (N_18484,N_13424,N_12344);
nand U18485 (N_18485,N_13423,N_14907);
nand U18486 (N_18486,N_13165,N_11338);
nor U18487 (N_18487,N_13651,N_13841);
or U18488 (N_18488,N_11785,N_14397);
or U18489 (N_18489,N_10227,N_10581);
and U18490 (N_18490,N_14076,N_13980);
nor U18491 (N_18491,N_12657,N_13024);
and U18492 (N_18492,N_12157,N_13031);
or U18493 (N_18493,N_12711,N_12744);
nand U18494 (N_18494,N_12541,N_10287);
or U18495 (N_18495,N_14825,N_10567);
or U18496 (N_18496,N_11792,N_13759);
nand U18497 (N_18497,N_10594,N_12124);
nor U18498 (N_18498,N_11869,N_13072);
nor U18499 (N_18499,N_10610,N_14787);
or U18500 (N_18500,N_10899,N_10002);
nor U18501 (N_18501,N_10295,N_11509);
nand U18502 (N_18502,N_10731,N_10301);
and U18503 (N_18503,N_13155,N_14928);
nand U18504 (N_18504,N_13246,N_14924);
nor U18505 (N_18505,N_12268,N_14159);
or U18506 (N_18506,N_10240,N_14253);
xor U18507 (N_18507,N_10582,N_13294);
nand U18508 (N_18508,N_11010,N_11312);
or U18509 (N_18509,N_13681,N_10703);
nor U18510 (N_18510,N_13492,N_10237);
and U18511 (N_18511,N_13461,N_13438);
or U18512 (N_18512,N_13953,N_11616);
and U18513 (N_18513,N_11806,N_11012);
nand U18514 (N_18514,N_13406,N_12045);
nand U18515 (N_18515,N_12327,N_13992);
nor U18516 (N_18516,N_10887,N_13163);
nor U18517 (N_18517,N_13974,N_11930);
nor U18518 (N_18518,N_13207,N_12076);
or U18519 (N_18519,N_14125,N_12063);
and U18520 (N_18520,N_12870,N_11428);
and U18521 (N_18521,N_13819,N_11566);
nor U18522 (N_18522,N_14421,N_14562);
nand U18523 (N_18523,N_14372,N_13939);
nor U18524 (N_18524,N_13287,N_11882);
or U18525 (N_18525,N_13357,N_13904);
nand U18526 (N_18526,N_12307,N_12691);
nor U18527 (N_18527,N_12907,N_14020);
or U18528 (N_18528,N_13773,N_12899);
xor U18529 (N_18529,N_14902,N_11416);
nor U18530 (N_18530,N_14834,N_11485);
nand U18531 (N_18531,N_14419,N_14856);
nand U18532 (N_18532,N_11477,N_14332);
nand U18533 (N_18533,N_13794,N_12429);
and U18534 (N_18534,N_10833,N_12633);
and U18535 (N_18535,N_10636,N_11727);
nor U18536 (N_18536,N_13331,N_13064);
nor U18537 (N_18537,N_12793,N_11762);
nand U18538 (N_18538,N_10531,N_13750);
nand U18539 (N_18539,N_14670,N_12145);
nand U18540 (N_18540,N_14406,N_13779);
nor U18541 (N_18541,N_12786,N_13018);
or U18542 (N_18542,N_12132,N_13931);
nor U18543 (N_18543,N_13842,N_13185);
and U18544 (N_18544,N_11390,N_13518);
nand U18545 (N_18545,N_14907,N_10002);
nor U18546 (N_18546,N_10875,N_14833);
and U18547 (N_18547,N_11647,N_14300);
or U18548 (N_18548,N_11656,N_10654);
or U18549 (N_18549,N_10124,N_14514);
and U18550 (N_18550,N_11487,N_14158);
nand U18551 (N_18551,N_10089,N_11950);
nor U18552 (N_18552,N_12589,N_11717);
and U18553 (N_18553,N_10517,N_12590);
and U18554 (N_18554,N_12280,N_12905);
and U18555 (N_18555,N_12938,N_10931);
and U18556 (N_18556,N_14711,N_13447);
and U18557 (N_18557,N_11842,N_10948);
or U18558 (N_18558,N_11299,N_10367);
and U18559 (N_18559,N_13081,N_10286);
or U18560 (N_18560,N_11504,N_11502);
nor U18561 (N_18561,N_12854,N_12905);
and U18562 (N_18562,N_14895,N_10500);
nor U18563 (N_18563,N_11326,N_12450);
and U18564 (N_18564,N_14942,N_14168);
nor U18565 (N_18565,N_12117,N_12705);
nor U18566 (N_18566,N_14357,N_11482);
nor U18567 (N_18567,N_10716,N_13327);
or U18568 (N_18568,N_11260,N_10117);
or U18569 (N_18569,N_14084,N_12474);
and U18570 (N_18570,N_12517,N_11843);
nor U18571 (N_18571,N_11917,N_13484);
nand U18572 (N_18572,N_11204,N_11303);
nand U18573 (N_18573,N_13197,N_13938);
and U18574 (N_18574,N_12528,N_11284);
nor U18575 (N_18575,N_14812,N_14264);
or U18576 (N_18576,N_14703,N_10480);
or U18577 (N_18577,N_13734,N_14991);
and U18578 (N_18578,N_13498,N_14058);
nor U18579 (N_18579,N_11447,N_10166);
and U18580 (N_18580,N_14837,N_14412);
or U18581 (N_18581,N_10641,N_13272);
nand U18582 (N_18582,N_10750,N_11495);
and U18583 (N_18583,N_13980,N_10872);
and U18584 (N_18584,N_14600,N_13093);
nor U18585 (N_18585,N_10141,N_10307);
nor U18586 (N_18586,N_11908,N_10855);
nand U18587 (N_18587,N_13020,N_10860);
nor U18588 (N_18588,N_12107,N_13615);
and U18589 (N_18589,N_12088,N_13765);
or U18590 (N_18590,N_12486,N_13446);
nand U18591 (N_18591,N_10295,N_11160);
nand U18592 (N_18592,N_12863,N_10411);
and U18593 (N_18593,N_14840,N_11735);
or U18594 (N_18594,N_11132,N_12090);
or U18595 (N_18595,N_14272,N_13596);
and U18596 (N_18596,N_14365,N_11820);
or U18597 (N_18597,N_10680,N_11165);
xnor U18598 (N_18598,N_11141,N_14621);
and U18599 (N_18599,N_12781,N_10294);
nand U18600 (N_18600,N_13105,N_11039);
and U18601 (N_18601,N_10785,N_11541);
nor U18602 (N_18602,N_14404,N_10085);
and U18603 (N_18603,N_10486,N_11926);
or U18604 (N_18604,N_13021,N_13536);
or U18605 (N_18605,N_14626,N_14262);
nand U18606 (N_18606,N_10064,N_11176);
nor U18607 (N_18607,N_12546,N_13242);
nand U18608 (N_18608,N_12253,N_10055);
and U18609 (N_18609,N_10728,N_14257);
nor U18610 (N_18610,N_13090,N_10528);
or U18611 (N_18611,N_10197,N_14107);
and U18612 (N_18612,N_11176,N_13055);
nand U18613 (N_18613,N_14479,N_11335);
nor U18614 (N_18614,N_13993,N_14817);
xnor U18615 (N_18615,N_14381,N_13053);
nor U18616 (N_18616,N_10309,N_12762);
and U18617 (N_18617,N_10835,N_13230);
and U18618 (N_18618,N_11157,N_12802);
nand U18619 (N_18619,N_14209,N_13430);
and U18620 (N_18620,N_13382,N_12375);
and U18621 (N_18621,N_13282,N_14132);
nor U18622 (N_18622,N_12415,N_13000);
xor U18623 (N_18623,N_13879,N_10034);
or U18624 (N_18624,N_10848,N_10432);
nand U18625 (N_18625,N_11135,N_11625);
nor U18626 (N_18626,N_14828,N_12152);
or U18627 (N_18627,N_10062,N_10700);
or U18628 (N_18628,N_14882,N_14830);
and U18629 (N_18629,N_14299,N_10919);
nor U18630 (N_18630,N_10655,N_12797);
or U18631 (N_18631,N_14340,N_14029);
and U18632 (N_18632,N_10889,N_11908);
nor U18633 (N_18633,N_10126,N_10903);
and U18634 (N_18634,N_12076,N_12209);
and U18635 (N_18635,N_14093,N_10249);
and U18636 (N_18636,N_13846,N_13755);
or U18637 (N_18637,N_11984,N_14688);
nor U18638 (N_18638,N_12024,N_11934);
nor U18639 (N_18639,N_12746,N_12738);
nor U18640 (N_18640,N_14659,N_13913);
nand U18641 (N_18641,N_12879,N_14689);
nand U18642 (N_18642,N_13655,N_12878);
or U18643 (N_18643,N_13673,N_12297);
or U18644 (N_18644,N_13780,N_10120);
and U18645 (N_18645,N_12546,N_11614);
or U18646 (N_18646,N_10863,N_14673);
or U18647 (N_18647,N_13818,N_11183);
nand U18648 (N_18648,N_11670,N_12358);
nor U18649 (N_18649,N_12523,N_10477);
xor U18650 (N_18650,N_12569,N_13606);
nand U18651 (N_18651,N_11566,N_11223);
and U18652 (N_18652,N_14663,N_10827);
nand U18653 (N_18653,N_11298,N_14480);
nand U18654 (N_18654,N_13028,N_14275);
nand U18655 (N_18655,N_12226,N_11812);
and U18656 (N_18656,N_12838,N_13786);
nor U18657 (N_18657,N_11063,N_11390);
nor U18658 (N_18658,N_10247,N_11150);
and U18659 (N_18659,N_11805,N_12998);
and U18660 (N_18660,N_14668,N_12844);
nor U18661 (N_18661,N_14029,N_11467);
or U18662 (N_18662,N_11533,N_10171);
and U18663 (N_18663,N_10781,N_11411);
or U18664 (N_18664,N_10825,N_14606);
nor U18665 (N_18665,N_11853,N_13016);
nor U18666 (N_18666,N_11836,N_14236);
nand U18667 (N_18667,N_13771,N_12261);
or U18668 (N_18668,N_11528,N_14731);
nand U18669 (N_18669,N_13503,N_11508);
and U18670 (N_18670,N_10628,N_10662);
nand U18671 (N_18671,N_10514,N_10010);
nand U18672 (N_18672,N_11266,N_12599);
nor U18673 (N_18673,N_11210,N_13398);
nor U18674 (N_18674,N_12086,N_11954);
nand U18675 (N_18675,N_13711,N_11773);
nand U18676 (N_18676,N_10060,N_12846);
xor U18677 (N_18677,N_13788,N_11379);
nor U18678 (N_18678,N_11450,N_10446);
or U18679 (N_18679,N_10614,N_11691);
nand U18680 (N_18680,N_13298,N_12980);
and U18681 (N_18681,N_14484,N_12693);
and U18682 (N_18682,N_12441,N_14578);
nor U18683 (N_18683,N_10524,N_10463);
or U18684 (N_18684,N_13966,N_13190);
nand U18685 (N_18685,N_12053,N_14825);
or U18686 (N_18686,N_14036,N_10365);
and U18687 (N_18687,N_11187,N_12534);
nor U18688 (N_18688,N_13879,N_11225);
or U18689 (N_18689,N_14735,N_10184);
and U18690 (N_18690,N_13053,N_12080);
nor U18691 (N_18691,N_11044,N_14745);
nor U18692 (N_18692,N_11514,N_13285);
and U18693 (N_18693,N_13387,N_13955);
nor U18694 (N_18694,N_14035,N_10455);
or U18695 (N_18695,N_12162,N_11390);
or U18696 (N_18696,N_12930,N_10244);
and U18697 (N_18697,N_12203,N_13406);
and U18698 (N_18698,N_11570,N_13724);
and U18699 (N_18699,N_13640,N_13531);
nor U18700 (N_18700,N_10817,N_14682);
nand U18701 (N_18701,N_10628,N_10637);
and U18702 (N_18702,N_12651,N_10674);
or U18703 (N_18703,N_13741,N_10497);
or U18704 (N_18704,N_14110,N_10848);
nand U18705 (N_18705,N_10660,N_12828);
or U18706 (N_18706,N_12027,N_10889);
and U18707 (N_18707,N_10934,N_10397);
nand U18708 (N_18708,N_12113,N_12400);
or U18709 (N_18709,N_11655,N_14446);
nand U18710 (N_18710,N_12777,N_12079);
or U18711 (N_18711,N_13309,N_13523);
nor U18712 (N_18712,N_13523,N_10456);
nand U18713 (N_18713,N_10557,N_13998);
nand U18714 (N_18714,N_11362,N_12242);
nor U18715 (N_18715,N_14455,N_11260);
nand U18716 (N_18716,N_10888,N_12040);
and U18717 (N_18717,N_12293,N_11744);
or U18718 (N_18718,N_13312,N_11792);
or U18719 (N_18719,N_11657,N_10439);
xnor U18720 (N_18720,N_12787,N_13605);
nor U18721 (N_18721,N_13763,N_10102);
nor U18722 (N_18722,N_10233,N_14656);
or U18723 (N_18723,N_11884,N_13588);
nand U18724 (N_18724,N_12768,N_12039);
and U18725 (N_18725,N_12915,N_12304);
and U18726 (N_18726,N_10735,N_10736);
nand U18727 (N_18727,N_11422,N_11959);
nor U18728 (N_18728,N_11390,N_12525);
nor U18729 (N_18729,N_12655,N_10815);
and U18730 (N_18730,N_12123,N_12589);
or U18731 (N_18731,N_12582,N_10073);
nor U18732 (N_18732,N_10036,N_13364);
and U18733 (N_18733,N_14252,N_11737);
nor U18734 (N_18734,N_11313,N_11476);
and U18735 (N_18735,N_11073,N_13856);
nor U18736 (N_18736,N_13172,N_10656);
xnor U18737 (N_18737,N_11037,N_14321);
and U18738 (N_18738,N_12469,N_11220);
nor U18739 (N_18739,N_10802,N_12633);
nand U18740 (N_18740,N_12303,N_14193);
nand U18741 (N_18741,N_10907,N_14811);
and U18742 (N_18742,N_13008,N_14878);
nand U18743 (N_18743,N_11021,N_12607);
or U18744 (N_18744,N_14826,N_14891);
and U18745 (N_18745,N_14620,N_13787);
nor U18746 (N_18746,N_11848,N_11794);
or U18747 (N_18747,N_12086,N_12582);
and U18748 (N_18748,N_12565,N_10851);
nand U18749 (N_18749,N_14046,N_11254);
or U18750 (N_18750,N_14074,N_14237);
nand U18751 (N_18751,N_10828,N_10890);
and U18752 (N_18752,N_13395,N_12782);
nand U18753 (N_18753,N_11318,N_12351);
or U18754 (N_18754,N_13041,N_14268);
nor U18755 (N_18755,N_11142,N_13676);
nand U18756 (N_18756,N_12977,N_10578);
nor U18757 (N_18757,N_10767,N_12417);
or U18758 (N_18758,N_14463,N_11237);
nor U18759 (N_18759,N_13814,N_10360);
nand U18760 (N_18760,N_11585,N_11987);
or U18761 (N_18761,N_11603,N_14520);
or U18762 (N_18762,N_13656,N_12697);
nand U18763 (N_18763,N_12870,N_12764);
nor U18764 (N_18764,N_12385,N_12365);
or U18765 (N_18765,N_12033,N_14517);
nand U18766 (N_18766,N_11652,N_12910);
nor U18767 (N_18767,N_14027,N_12507);
nor U18768 (N_18768,N_11757,N_13729);
nand U18769 (N_18769,N_11875,N_10638);
or U18770 (N_18770,N_11560,N_12013);
and U18771 (N_18771,N_12414,N_14109);
nor U18772 (N_18772,N_14682,N_13191);
and U18773 (N_18773,N_13829,N_13168);
xnor U18774 (N_18774,N_13227,N_12424);
or U18775 (N_18775,N_11412,N_11162);
nand U18776 (N_18776,N_14692,N_10514);
nand U18777 (N_18777,N_14751,N_14222);
or U18778 (N_18778,N_11480,N_10939);
or U18779 (N_18779,N_10098,N_12525);
nand U18780 (N_18780,N_11229,N_10885);
nor U18781 (N_18781,N_11465,N_12779);
and U18782 (N_18782,N_11637,N_10183);
and U18783 (N_18783,N_13900,N_14741);
and U18784 (N_18784,N_10029,N_13113);
and U18785 (N_18785,N_14625,N_12929);
nor U18786 (N_18786,N_10484,N_11518);
or U18787 (N_18787,N_10509,N_14852);
xor U18788 (N_18788,N_10629,N_12853);
or U18789 (N_18789,N_13766,N_14137);
and U18790 (N_18790,N_10813,N_11154);
nor U18791 (N_18791,N_14893,N_14260);
nand U18792 (N_18792,N_12797,N_14631);
or U18793 (N_18793,N_13121,N_12269);
nor U18794 (N_18794,N_13692,N_12066);
nand U18795 (N_18795,N_13479,N_12515);
nor U18796 (N_18796,N_12016,N_10440);
or U18797 (N_18797,N_10470,N_13061);
nand U18798 (N_18798,N_14399,N_12782);
and U18799 (N_18799,N_11980,N_12574);
nor U18800 (N_18800,N_11769,N_14464);
and U18801 (N_18801,N_11916,N_14501);
nor U18802 (N_18802,N_12786,N_14040);
nor U18803 (N_18803,N_14996,N_14396);
nand U18804 (N_18804,N_14186,N_14166);
nand U18805 (N_18805,N_11999,N_11150);
or U18806 (N_18806,N_10332,N_14571);
nand U18807 (N_18807,N_12884,N_12221);
or U18808 (N_18808,N_13501,N_12295);
or U18809 (N_18809,N_14871,N_11613);
nand U18810 (N_18810,N_11453,N_10202);
or U18811 (N_18811,N_12396,N_11179);
nand U18812 (N_18812,N_12010,N_10756);
nor U18813 (N_18813,N_13528,N_10951);
nand U18814 (N_18814,N_14914,N_10956);
or U18815 (N_18815,N_12685,N_14379);
nand U18816 (N_18816,N_10944,N_14004);
nand U18817 (N_18817,N_11618,N_10460);
nor U18818 (N_18818,N_11023,N_13316);
xnor U18819 (N_18819,N_12793,N_11116);
or U18820 (N_18820,N_12385,N_12546);
or U18821 (N_18821,N_14746,N_12085);
nand U18822 (N_18822,N_13392,N_12411);
nor U18823 (N_18823,N_13583,N_14667);
xor U18824 (N_18824,N_12817,N_11742);
and U18825 (N_18825,N_13653,N_14615);
and U18826 (N_18826,N_14047,N_13657);
or U18827 (N_18827,N_14209,N_12567);
nand U18828 (N_18828,N_11935,N_14823);
nor U18829 (N_18829,N_12827,N_11636);
nand U18830 (N_18830,N_13266,N_12373);
and U18831 (N_18831,N_13338,N_11864);
nand U18832 (N_18832,N_14527,N_14696);
nor U18833 (N_18833,N_12411,N_12518);
nand U18834 (N_18834,N_13582,N_14011);
nor U18835 (N_18835,N_13383,N_12136);
xor U18836 (N_18836,N_13489,N_12022);
or U18837 (N_18837,N_14285,N_14532);
nor U18838 (N_18838,N_13643,N_14788);
or U18839 (N_18839,N_12218,N_12072);
nor U18840 (N_18840,N_12471,N_11839);
or U18841 (N_18841,N_14710,N_13128);
nand U18842 (N_18842,N_14873,N_13385);
nand U18843 (N_18843,N_13786,N_11885);
nor U18844 (N_18844,N_12786,N_14718);
nand U18845 (N_18845,N_11893,N_12216);
and U18846 (N_18846,N_11463,N_12168);
nand U18847 (N_18847,N_13527,N_14268);
nand U18848 (N_18848,N_10034,N_13875);
and U18849 (N_18849,N_13150,N_14880);
nand U18850 (N_18850,N_13941,N_10171);
nand U18851 (N_18851,N_13596,N_13136);
or U18852 (N_18852,N_13723,N_12702);
and U18853 (N_18853,N_13724,N_12794);
nand U18854 (N_18854,N_14029,N_13036);
nand U18855 (N_18855,N_12775,N_12545);
nor U18856 (N_18856,N_11776,N_12993);
nor U18857 (N_18857,N_12196,N_11027);
and U18858 (N_18858,N_13193,N_10037);
or U18859 (N_18859,N_14620,N_14560);
and U18860 (N_18860,N_12525,N_11373);
and U18861 (N_18861,N_13646,N_14694);
and U18862 (N_18862,N_13801,N_14427);
or U18863 (N_18863,N_10893,N_11240);
or U18864 (N_18864,N_12703,N_11768);
or U18865 (N_18865,N_10273,N_11701);
or U18866 (N_18866,N_10494,N_13522);
nand U18867 (N_18867,N_12202,N_11083);
nor U18868 (N_18868,N_10048,N_12612);
xnor U18869 (N_18869,N_12103,N_13388);
and U18870 (N_18870,N_12094,N_10408);
nor U18871 (N_18871,N_13841,N_14025);
and U18872 (N_18872,N_14040,N_11788);
and U18873 (N_18873,N_11883,N_11423);
or U18874 (N_18874,N_13845,N_13521);
nor U18875 (N_18875,N_12869,N_10269);
nor U18876 (N_18876,N_14761,N_11985);
nor U18877 (N_18877,N_11190,N_11404);
xnor U18878 (N_18878,N_12232,N_13863);
nand U18879 (N_18879,N_12267,N_12271);
nand U18880 (N_18880,N_11939,N_13065);
nor U18881 (N_18881,N_12376,N_11448);
nand U18882 (N_18882,N_10337,N_13515);
nor U18883 (N_18883,N_10268,N_12978);
and U18884 (N_18884,N_11564,N_14629);
nand U18885 (N_18885,N_11689,N_10261);
nor U18886 (N_18886,N_10117,N_10761);
nor U18887 (N_18887,N_14984,N_14104);
nand U18888 (N_18888,N_12741,N_14483);
nor U18889 (N_18889,N_13771,N_11685);
nand U18890 (N_18890,N_11249,N_14012);
or U18891 (N_18891,N_12789,N_14474);
nand U18892 (N_18892,N_14916,N_13626);
or U18893 (N_18893,N_14940,N_11458);
nor U18894 (N_18894,N_11362,N_10896);
and U18895 (N_18895,N_11198,N_12482);
and U18896 (N_18896,N_10276,N_11124);
and U18897 (N_18897,N_14710,N_12516);
or U18898 (N_18898,N_13188,N_13233);
and U18899 (N_18899,N_10921,N_14410);
and U18900 (N_18900,N_13472,N_11960);
nand U18901 (N_18901,N_12586,N_14383);
xnor U18902 (N_18902,N_10420,N_12233);
and U18903 (N_18903,N_12600,N_11214);
or U18904 (N_18904,N_13050,N_12300);
nand U18905 (N_18905,N_12850,N_12378);
nand U18906 (N_18906,N_11342,N_14447);
nor U18907 (N_18907,N_12412,N_11901);
or U18908 (N_18908,N_14678,N_14918);
nor U18909 (N_18909,N_10901,N_11002);
and U18910 (N_18910,N_12517,N_12532);
nor U18911 (N_18911,N_14528,N_14219);
nor U18912 (N_18912,N_13531,N_10225);
nor U18913 (N_18913,N_11292,N_13057);
and U18914 (N_18914,N_14426,N_12298);
and U18915 (N_18915,N_13877,N_14401);
or U18916 (N_18916,N_11246,N_12427);
and U18917 (N_18917,N_10593,N_13728);
nand U18918 (N_18918,N_13089,N_11351);
nand U18919 (N_18919,N_12292,N_11140);
and U18920 (N_18920,N_12621,N_13625);
nand U18921 (N_18921,N_11059,N_13060);
nor U18922 (N_18922,N_12730,N_14542);
nand U18923 (N_18923,N_13462,N_13540);
and U18924 (N_18924,N_13801,N_14071);
nor U18925 (N_18925,N_14115,N_12247);
and U18926 (N_18926,N_11028,N_12657);
nor U18927 (N_18927,N_12889,N_13961);
nand U18928 (N_18928,N_10082,N_12009);
or U18929 (N_18929,N_11148,N_12043);
and U18930 (N_18930,N_10284,N_14259);
nand U18931 (N_18931,N_14788,N_11560);
nor U18932 (N_18932,N_13411,N_11053);
and U18933 (N_18933,N_11301,N_13145);
nor U18934 (N_18934,N_14787,N_12901);
nor U18935 (N_18935,N_13800,N_10350);
nand U18936 (N_18936,N_14658,N_14684);
nand U18937 (N_18937,N_10764,N_12082);
nand U18938 (N_18938,N_14064,N_13861);
nor U18939 (N_18939,N_14630,N_10056);
or U18940 (N_18940,N_12937,N_11862);
nor U18941 (N_18941,N_13021,N_14921);
or U18942 (N_18942,N_14058,N_14522);
nor U18943 (N_18943,N_11091,N_13649);
and U18944 (N_18944,N_14804,N_10321);
and U18945 (N_18945,N_10904,N_13634);
and U18946 (N_18946,N_13400,N_11944);
or U18947 (N_18947,N_12641,N_10063);
and U18948 (N_18948,N_12784,N_11116);
or U18949 (N_18949,N_11255,N_12124);
nor U18950 (N_18950,N_11602,N_13716);
nand U18951 (N_18951,N_12828,N_13814);
and U18952 (N_18952,N_12586,N_14307);
nand U18953 (N_18953,N_12476,N_10730);
nor U18954 (N_18954,N_13534,N_10861);
and U18955 (N_18955,N_13666,N_14634);
nor U18956 (N_18956,N_11422,N_10853);
nor U18957 (N_18957,N_14126,N_10302);
nand U18958 (N_18958,N_12600,N_10564);
nor U18959 (N_18959,N_10206,N_13928);
or U18960 (N_18960,N_10526,N_13939);
nand U18961 (N_18961,N_10818,N_11843);
nor U18962 (N_18962,N_11710,N_13975);
and U18963 (N_18963,N_11317,N_10415);
and U18964 (N_18964,N_10814,N_12372);
or U18965 (N_18965,N_10125,N_10267);
nor U18966 (N_18966,N_12061,N_12610);
nand U18967 (N_18967,N_11147,N_13445);
and U18968 (N_18968,N_11887,N_12967);
or U18969 (N_18969,N_13919,N_11722);
or U18970 (N_18970,N_13070,N_12976);
nand U18971 (N_18971,N_13034,N_14995);
nor U18972 (N_18972,N_10866,N_14507);
nor U18973 (N_18973,N_13550,N_11117);
and U18974 (N_18974,N_10766,N_12853);
or U18975 (N_18975,N_11937,N_11669);
and U18976 (N_18976,N_12442,N_13479);
or U18977 (N_18977,N_13293,N_11882);
nand U18978 (N_18978,N_10920,N_14606);
nand U18979 (N_18979,N_14790,N_10384);
nand U18980 (N_18980,N_12086,N_11475);
and U18981 (N_18981,N_13136,N_11090);
or U18982 (N_18982,N_13568,N_14195);
and U18983 (N_18983,N_14114,N_11658);
or U18984 (N_18984,N_13009,N_13991);
nand U18985 (N_18985,N_12969,N_11514);
nand U18986 (N_18986,N_10547,N_10120);
and U18987 (N_18987,N_14344,N_12449);
nand U18988 (N_18988,N_12841,N_11299);
nor U18989 (N_18989,N_10569,N_12445);
nor U18990 (N_18990,N_12721,N_11804);
nand U18991 (N_18991,N_11040,N_12134);
nand U18992 (N_18992,N_11630,N_13117);
or U18993 (N_18993,N_11295,N_13606);
and U18994 (N_18994,N_11157,N_14568);
nor U18995 (N_18995,N_11758,N_10582);
nor U18996 (N_18996,N_12138,N_11795);
nand U18997 (N_18997,N_13074,N_11301);
or U18998 (N_18998,N_12293,N_13241);
and U18999 (N_18999,N_13516,N_12431);
nand U19000 (N_19000,N_12966,N_10668);
nor U19001 (N_19001,N_13516,N_11812);
and U19002 (N_19002,N_12821,N_10687);
nor U19003 (N_19003,N_10310,N_14615);
nor U19004 (N_19004,N_11349,N_10696);
or U19005 (N_19005,N_14074,N_12997);
or U19006 (N_19006,N_13778,N_13054);
or U19007 (N_19007,N_11822,N_12910);
nor U19008 (N_19008,N_11243,N_14399);
nor U19009 (N_19009,N_11259,N_14727);
nand U19010 (N_19010,N_11026,N_13987);
nor U19011 (N_19011,N_11163,N_11332);
nand U19012 (N_19012,N_11494,N_14049);
and U19013 (N_19013,N_14592,N_11369);
or U19014 (N_19014,N_12932,N_13593);
nand U19015 (N_19015,N_12662,N_12004);
nor U19016 (N_19016,N_13858,N_11206);
nor U19017 (N_19017,N_14128,N_13685);
nand U19018 (N_19018,N_14932,N_13314);
or U19019 (N_19019,N_11288,N_14645);
nor U19020 (N_19020,N_10775,N_12936);
or U19021 (N_19021,N_12113,N_13248);
and U19022 (N_19022,N_11407,N_12866);
nor U19023 (N_19023,N_10381,N_10678);
nand U19024 (N_19024,N_11570,N_10055);
or U19025 (N_19025,N_14913,N_13573);
nand U19026 (N_19026,N_14229,N_10380);
and U19027 (N_19027,N_14044,N_10020);
nand U19028 (N_19028,N_11263,N_11585);
and U19029 (N_19029,N_11203,N_10251);
nand U19030 (N_19030,N_11792,N_12333);
and U19031 (N_19031,N_12304,N_11183);
and U19032 (N_19032,N_11178,N_11508);
nor U19033 (N_19033,N_13321,N_14528);
nand U19034 (N_19034,N_14248,N_12246);
or U19035 (N_19035,N_14401,N_14577);
nor U19036 (N_19036,N_10122,N_11554);
or U19037 (N_19037,N_13733,N_13793);
and U19038 (N_19038,N_12595,N_12577);
nand U19039 (N_19039,N_13582,N_10204);
nand U19040 (N_19040,N_12586,N_13591);
and U19041 (N_19041,N_11000,N_13198);
nor U19042 (N_19042,N_13801,N_14555);
and U19043 (N_19043,N_12025,N_10714);
nand U19044 (N_19044,N_10564,N_11114);
nand U19045 (N_19045,N_12798,N_12025);
nand U19046 (N_19046,N_13363,N_13513);
nand U19047 (N_19047,N_12894,N_11345);
nand U19048 (N_19048,N_13149,N_12944);
or U19049 (N_19049,N_10703,N_12751);
and U19050 (N_19050,N_13623,N_12308);
or U19051 (N_19051,N_12346,N_12019);
nor U19052 (N_19052,N_14988,N_14885);
xor U19053 (N_19053,N_13337,N_11604);
and U19054 (N_19054,N_10803,N_11349);
and U19055 (N_19055,N_13520,N_11422);
and U19056 (N_19056,N_12474,N_12488);
and U19057 (N_19057,N_11740,N_10950);
nand U19058 (N_19058,N_13340,N_10071);
and U19059 (N_19059,N_12479,N_12890);
or U19060 (N_19060,N_11574,N_11705);
nand U19061 (N_19061,N_11703,N_14028);
and U19062 (N_19062,N_11418,N_10164);
nor U19063 (N_19063,N_13176,N_12816);
or U19064 (N_19064,N_13192,N_11969);
and U19065 (N_19065,N_11920,N_14136);
or U19066 (N_19066,N_14742,N_14860);
or U19067 (N_19067,N_10047,N_13498);
nand U19068 (N_19068,N_12147,N_13893);
nor U19069 (N_19069,N_13331,N_14956);
nor U19070 (N_19070,N_10057,N_11904);
nor U19071 (N_19071,N_14775,N_13774);
and U19072 (N_19072,N_14810,N_12150);
and U19073 (N_19073,N_12200,N_13645);
nor U19074 (N_19074,N_11230,N_10794);
nor U19075 (N_19075,N_13070,N_11160);
or U19076 (N_19076,N_12330,N_11753);
nor U19077 (N_19077,N_14804,N_14869);
nor U19078 (N_19078,N_11320,N_11103);
nand U19079 (N_19079,N_13589,N_12554);
and U19080 (N_19080,N_13098,N_13525);
or U19081 (N_19081,N_10893,N_13752);
and U19082 (N_19082,N_11670,N_11944);
nand U19083 (N_19083,N_14367,N_12177);
or U19084 (N_19084,N_11537,N_12951);
nand U19085 (N_19085,N_10172,N_13140);
nand U19086 (N_19086,N_10367,N_14763);
and U19087 (N_19087,N_13394,N_10698);
nand U19088 (N_19088,N_14958,N_12443);
nand U19089 (N_19089,N_10513,N_10010);
and U19090 (N_19090,N_14580,N_14238);
and U19091 (N_19091,N_11560,N_10754);
or U19092 (N_19092,N_14959,N_13013);
nand U19093 (N_19093,N_10584,N_13915);
or U19094 (N_19094,N_11366,N_14115);
nand U19095 (N_19095,N_11855,N_11325);
nor U19096 (N_19096,N_11806,N_12747);
or U19097 (N_19097,N_13550,N_13152);
nor U19098 (N_19098,N_12620,N_13190);
and U19099 (N_19099,N_14475,N_10320);
or U19100 (N_19100,N_14813,N_10365);
and U19101 (N_19101,N_14539,N_11159);
nand U19102 (N_19102,N_11976,N_11009);
nor U19103 (N_19103,N_10490,N_14005);
nor U19104 (N_19104,N_12416,N_10388);
nand U19105 (N_19105,N_10737,N_13276);
and U19106 (N_19106,N_13038,N_11433);
and U19107 (N_19107,N_12404,N_12857);
nand U19108 (N_19108,N_12326,N_10816);
or U19109 (N_19109,N_13620,N_13781);
and U19110 (N_19110,N_12041,N_11038);
nand U19111 (N_19111,N_10476,N_12867);
xor U19112 (N_19112,N_13050,N_10474);
or U19113 (N_19113,N_10380,N_13794);
or U19114 (N_19114,N_11165,N_10323);
and U19115 (N_19115,N_10645,N_10455);
nor U19116 (N_19116,N_13056,N_10265);
nor U19117 (N_19117,N_11979,N_10156);
nor U19118 (N_19118,N_10760,N_12735);
and U19119 (N_19119,N_10278,N_13055);
or U19120 (N_19120,N_14517,N_12899);
and U19121 (N_19121,N_14674,N_10423);
xnor U19122 (N_19122,N_13145,N_11444);
or U19123 (N_19123,N_12392,N_13818);
nand U19124 (N_19124,N_12149,N_11539);
nand U19125 (N_19125,N_11663,N_12061);
nand U19126 (N_19126,N_12656,N_11349);
and U19127 (N_19127,N_11944,N_10653);
nand U19128 (N_19128,N_13386,N_14121);
nand U19129 (N_19129,N_13338,N_12134);
or U19130 (N_19130,N_11101,N_10178);
or U19131 (N_19131,N_12957,N_10533);
and U19132 (N_19132,N_12474,N_14880);
nand U19133 (N_19133,N_12456,N_11381);
and U19134 (N_19134,N_10454,N_12085);
or U19135 (N_19135,N_13063,N_11159);
nor U19136 (N_19136,N_11316,N_13827);
nor U19137 (N_19137,N_14461,N_14822);
and U19138 (N_19138,N_12820,N_11119);
or U19139 (N_19139,N_12592,N_10176);
or U19140 (N_19140,N_10623,N_11573);
and U19141 (N_19141,N_13717,N_13390);
or U19142 (N_19142,N_13923,N_11805);
nand U19143 (N_19143,N_13340,N_13973);
and U19144 (N_19144,N_10694,N_11437);
nor U19145 (N_19145,N_12840,N_10704);
nor U19146 (N_19146,N_12947,N_13005);
and U19147 (N_19147,N_12817,N_11777);
nand U19148 (N_19148,N_10313,N_13592);
nand U19149 (N_19149,N_14580,N_14101);
or U19150 (N_19150,N_11615,N_14840);
nor U19151 (N_19151,N_10007,N_14421);
nand U19152 (N_19152,N_14949,N_10793);
or U19153 (N_19153,N_13116,N_12353);
or U19154 (N_19154,N_12970,N_13504);
and U19155 (N_19155,N_11739,N_11761);
nor U19156 (N_19156,N_14018,N_12329);
and U19157 (N_19157,N_12554,N_14395);
or U19158 (N_19158,N_13222,N_14635);
or U19159 (N_19159,N_13940,N_10107);
nor U19160 (N_19160,N_10058,N_12237);
and U19161 (N_19161,N_13662,N_10195);
nand U19162 (N_19162,N_12479,N_11308);
nand U19163 (N_19163,N_10625,N_13196);
or U19164 (N_19164,N_13508,N_10380);
or U19165 (N_19165,N_12598,N_11442);
and U19166 (N_19166,N_11726,N_13784);
or U19167 (N_19167,N_14059,N_11253);
and U19168 (N_19168,N_10138,N_14336);
nand U19169 (N_19169,N_14356,N_10999);
or U19170 (N_19170,N_10125,N_13086);
or U19171 (N_19171,N_12732,N_11068);
nor U19172 (N_19172,N_11250,N_10290);
and U19173 (N_19173,N_10545,N_12338);
nor U19174 (N_19174,N_14128,N_11503);
and U19175 (N_19175,N_10570,N_11009);
or U19176 (N_19176,N_10530,N_11572);
and U19177 (N_19177,N_10215,N_10227);
nor U19178 (N_19178,N_11227,N_13475);
nor U19179 (N_19179,N_10918,N_13453);
and U19180 (N_19180,N_11709,N_12502);
and U19181 (N_19181,N_11537,N_10816);
and U19182 (N_19182,N_12022,N_11963);
and U19183 (N_19183,N_11174,N_12169);
nor U19184 (N_19184,N_11466,N_14365);
and U19185 (N_19185,N_13102,N_10509);
and U19186 (N_19186,N_10469,N_13646);
nor U19187 (N_19187,N_11916,N_10048);
nand U19188 (N_19188,N_12367,N_12907);
nand U19189 (N_19189,N_13249,N_13405);
nand U19190 (N_19190,N_12146,N_12106);
nand U19191 (N_19191,N_10744,N_13396);
and U19192 (N_19192,N_13991,N_13602);
or U19193 (N_19193,N_11809,N_14959);
nor U19194 (N_19194,N_14134,N_11385);
nor U19195 (N_19195,N_11609,N_12617);
nor U19196 (N_19196,N_11301,N_12918);
nand U19197 (N_19197,N_14878,N_11013);
nor U19198 (N_19198,N_12143,N_14494);
or U19199 (N_19199,N_11012,N_14464);
and U19200 (N_19200,N_11017,N_13439);
and U19201 (N_19201,N_12204,N_12593);
or U19202 (N_19202,N_13756,N_14963);
nand U19203 (N_19203,N_13473,N_10383);
or U19204 (N_19204,N_14860,N_10470);
or U19205 (N_19205,N_12224,N_10001);
or U19206 (N_19206,N_11513,N_12426);
nand U19207 (N_19207,N_11787,N_10648);
or U19208 (N_19208,N_12380,N_12486);
nor U19209 (N_19209,N_13315,N_14590);
nor U19210 (N_19210,N_13279,N_12286);
and U19211 (N_19211,N_14726,N_13389);
nor U19212 (N_19212,N_13322,N_13507);
nor U19213 (N_19213,N_10183,N_12038);
nor U19214 (N_19214,N_11805,N_13515);
nand U19215 (N_19215,N_10210,N_11407);
nor U19216 (N_19216,N_11506,N_10575);
nand U19217 (N_19217,N_12940,N_11709);
nor U19218 (N_19218,N_12078,N_14563);
and U19219 (N_19219,N_13170,N_14700);
nand U19220 (N_19220,N_11887,N_12704);
nor U19221 (N_19221,N_12262,N_13907);
nand U19222 (N_19222,N_13909,N_14936);
and U19223 (N_19223,N_11898,N_12881);
nor U19224 (N_19224,N_14882,N_12444);
nand U19225 (N_19225,N_12206,N_11571);
xnor U19226 (N_19226,N_14136,N_12249);
and U19227 (N_19227,N_10701,N_12372);
and U19228 (N_19228,N_11890,N_13261);
nand U19229 (N_19229,N_13993,N_12131);
nor U19230 (N_19230,N_14161,N_14845);
or U19231 (N_19231,N_14448,N_12635);
or U19232 (N_19232,N_14665,N_11761);
nor U19233 (N_19233,N_12779,N_12297);
nand U19234 (N_19234,N_13777,N_12845);
and U19235 (N_19235,N_12893,N_13123);
and U19236 (N_19236,N_11127,N_12212);
nand U19237 (N_19237,N_13945,N_12466);
and U19238 (N_19238,N_10431,N_11402);
nand U19239 (N_19239,N_12574,N_13839);
xnor U19240 (N_19240,N_13402,N_12399);
nor U19241 (N_19241,N_10851,N_12041);
or U19242 (N_19242,N_14810,N_13367);
and U19243 (N_19243,N_12032,N_10424);
or U19244 (N_19244,N_13838,N_13174);
nor U19245 (N_19245,N_10623,N_13415);
nor U19246 (N_19246,N_10268,N_12046);
and U19247 (N_19247,N_12508,N_14543);
nand U19248 (N_19248,N_11547,N_12128);
nor U19249 (N_19249,N_11521,N_12677);
and U19250 (N_19250,N_11430,N_11977);
nor U19251 (N_19251,N_14660,N_14472);
or U19252 (N_19252,N_12575,N_13413);
and U19253 (N_19253,N_10010,N_12159);
and U19254 (N_19254,N_11279,N_10481);
nor U19255 (N_19255,N_14876,N_13442);
or U19256 (N_19256,N_14244,N_14315);
and U19257 (N_19257,N_14250,N_10271);
nand U19258 (N_19258,N_13175,N_14313);
nor U19259 (N_19259,N_10414,N_12480);
and U19260 (N_19260,N_14224,N_10354);
or U19261 (N_19261,N_11376,N_12225);
nor U19262 (N_19262,N_12598,N_12321);
nand U19263 (N_19263,N_10552,N_10672);
nand U19264 (N_19264,N_13303,N_12247);
nand U19265 (N_19265,N_12964,N_12600);
nor U19266 (N_19266,N_10575,N_14556);
or U19267 (N_19267,N_10910,N_14788);
nand U19268 (N_19268,N_14831,N_13648);
nor U19269 (N_19269,N_11583,N_13723);
nor U19270 (N_19270,N_14907,N_10228);
or U19271 (N_19271,N_11076,N_13347);
or U19272 (N_19272,N_11967,N_12227);
nand U19273 (N_19273,N_11552,N_14729);
nand U19274 (N_19274,N_12262,N_11728);
xor U19275 (N_19275,N_11409,N_13083);
and U19276 (N_19276,N_10080,N_13927);
nor U19277 (N_19277,N_11035,N_13407);
or U19278 (N_19278,N_13508,N_12738);
or U19279 (N_19279,N_14544,N_13572);
nor U19280 (N_19280,N_12560,N_14082);
and U19281 (N_19281,N_12838,N_11438);
or U19282 (N_19282,N_10195,N_14658);
xnor U19283 (N_19283,N_10937,N_13203);
or U19284 (N_19284,N_14896,N_10480);
or U19285 (N_19285,N_14911,N_11659);
nand U19286 (N_19286,N_12441,N_12569);
and U19287 (N_19287,N_13396,N_13148);
and U19288 (N_19288,N_11158,N_11536);
and U19289 (N_19289,N_13232,N_13911);
or U19290 (N_19290,N_13210,N_14204);
nor U19291 (N_19291,N_10687,N_12245);
and U19292 (N_19292,N_13360,N_14830);
nand U19293 (N_19293,N_13993,N_10634);
nand U19294 (N_19294,N_12801,N_11119);
nor U19295 (N_19295,N_10749,N_10672);
nor U19296 (N_19296,N_12353,N_14016);
and U19297 (N_19297,N_11646,N_11002);
or U19298 (N_19298,N_13585,N_10943);
nand U19299 (N_19299,N_14803,N_10171);
nand U19300 (N_19300,N_13024,N_14646);
and U19301 (N_19301,N_14010,N_12972);
xor U19302 (N_19302,N_14357,N_14277);
or U19303 (N_19303,N_14248,N_13839);
nand U19304 (N_19304,N_12457,N_13239);
nor U19305 (N_19305,N_13927,N_12109);
nor U19306 (N_19306,N_12835,N_12259);
nand U19307 (N_19307,N_12663,N_11088);
and U19308 (N_19308,N_11109,N_11728);
or U19309 (N_19309,N_12593,N_14647);
or U19310 (N_19310,N_10245,N_11830);
nand U19311 (N_19311,N_11051,N_12140);
or U19312 (N_19312,N_10659,N_14385);
nand U19313 (N_19313,N_10419,N_11172);
or U19314 (N_19314,N_11563,N_14369);
nor U19315 (N_19315,N_13022,N_14185);
and U19316 (N_19316,N_14054,N_11538);
nor U19317 (N_19317,N_13282,N_14371);
or U19318 (N_19318,N_11869,N_11161);
nand U19319 (N_19319,N_11276,N_14352);
nand U19320 (N_19320,N_11650,N_13837);
nor U19321 (N_19321,N_14419,N_14289);
nand U19322 (N_19322,N_11054,N_13360);
nand U19323 (N_19323,N_14415,N_11861);
nor U19324 (N_19324,N_10744,N_14395);
nor U19325 (N_19325,N_11435,N_12743);
nand U19326 (N_19326,N_14617,N_12260);
and U19327 (N_19327,N_13967,N_11782);
and U19328 (N_19328,N_14552,N_10392);
or U19329 (N_19329,N_13198,N_12856);
nor U19330 (N_19330,N_12555,N_13030);
nor U19331 (N_19331,N_13646,N_13385);
and U19332 (N_19332,N_12744,N_14630);
or U19333 (N_19333,N_10594,N_11515);
and U19334 (N_19334,N_13927,N_13874);
nor U19335 (N_19335,N_14514,N_12134);
nor U19336 (N_19336,N_10545,N_13364);
and U19337 (N_19337,N_13754,N_12539);
and U19338 (N_19338,N_13621,N_11824);
and U19339 (N_19339,N_11674,N_12074);
nand U19340 (N_19340,N_10431,N_10847);
nand U19341 (N_19341,N_12429,N_10184);
or U19342 (N_19342,N_13578,N_13505);
nor U19343 (N_19343,N_14015,N_13323);
nand U19344 (N_19344,N_12118,N_13495);
nand U19345 (N_19345,N_11743,N_11614);
and U19346 (N_19346,N_14561,N_11760);
xnor U19347 (N_19347,N_12766,N_14179);
nor U19348 (N_19348,N_11701,N_11363);
or U19349 (N_19349,N_13692,N_10068);
nand U19350 (N_19350,N_14318,N_14981);
or U19351 (N_19351,N_12051,N_14772);
nand U19352 (N_19352,N_13204,N_13074);
or U19353 (N_19353,N_12687,N_10644);
and U19354 (N_19354,N_13774,N_10871);
and U19355 (N_19355,N_11924,N_10132);
nor U19356 (N_19356,N_12748,N_14351);
nand U19357 (N_19357,N_14428,N_14386);
or U19358 (N_19358,N_11096,N_14435);
or U19359 (N_19359,N_11701,N_12774);
and U19360 (N_19360,N_14093,N_10666);
or U19361 (N_19361,N_13091,N_13979);
nand U19362 (N_19362,N_10135,N_13530);
nand U19363 (N_19363,N_14680,N_10083);
nor U19364 (N_19364,N_12908,N_14282);
or U19365 (N_19365,N_10745,N_10078);
or U19366 (N_19366,N_12173,N_14404);
nand U19367 (N_19367,N_14750,N_14565);
nand U19368 (N_19368,N_10950,N_11450);
nand U19369 (N_19369,N_12133,N_14218);
and U19370 (N_19370,N_14994,N_11869);
nor U19371 (N_19371,N_11568,N_13721);
nand U19372 (N_19372,N_13142,N_14743);
or U19373 (N_19373,N_10972,N_12121);
or U19374 (N_19374,N_14950,N_10523);
nor U19375 (N_19375,N_12513,N_14932);
and U19376 (N_19376,N_10528,N_14354);
nor U19377 (N_19377,N_14649,N_14226);
and U19378 (N_19378,N_14201,N_11832);
nand U19379 (N_19379,N_14336,N_12426);
nand U19380 (N_19380,N_11343,N_12987);
and U19381 (N_19381,N_13415,N_14514);
nor U19382 (N_19382,N_13142,N_13066);
or U19383 (N_19383,N_10968,N_11136);
or U19384 (N_19384,N_13127,N_11454);
or U19385 (N_19385,N_11609,N_13123);
nand U19386 (N_19386,N_11516,N_13053);
and U19387 (N_19387,N_12326,N_10952);
and U19388 (N_19388,N_11000,N_11209);
and U19389 (N_19389,N_13010,N_13395);
nand U19390 (N_19390,N_10453,N_13948);
nor U19391 (N_19391,N_11668,N_11279);
and U19392 (N_19392,N_12859,N_12630);
and U19393 (N_19393,N_13355,N_10855);
or U19394 (N_19394,N_10656,N_13253);
nand U19395 (N_19395,N_10228,N_10532);
xor U19396 (N_19396,N_14699,N_13840);
nor U19397 (N_19397,N_13807,N_14402);
nand U19398 (N_19398,N_14265,N_10535);
nand U19399 (N_19399,N_14715,N_14352);
or U19400 (N_19400,N_12378,N_11888);
and U19401 (N_19401,N_14781,N_12406);
nor U19402 (N_19402,N_14820,N_13947);
nand U19403 (N_19403,N_14691,N_14279);
nand U19404 (N_19404,N_14367,N_11900);
nand U19405 (N_19405,N_10310,N_10076);
and U19406 (N_19406,N_13873,N_10775);
or U19407 (N_19407,N_11429,N_14652);
and U19408 (N_19408,N_13417,N_14776);
or U19409 (N_19409,N_14855,N_14906);
and U19410 (N_19410,N_14039,N_14290);
or U19411 (N_19411,N_10219,N_14212);
nor U19412 (N_19412,N_10220,N_12707);
nand U19413 (N_19413,N_10167,N_12186);
nand U19414 (N_19414,N_11452,N_12229);
nand U19415 (N_19415,N_11404,N_14652);
or U19416 (N_19416,N_14278,N_11104);
xnor U19417 (N_19417,N_10654,N_11328);
or U19418 (N_19418,N_13301,N_14541);
nor U19419 (N_19419,N_11110,N_13766);
and U19420 (N_19420,N_11983,N_10170);
and U19421 (N_19421,N_13820,N_10172);
nand U19422 (N_19422,N_10094,N_10938);
or U19423 (N_19423,N_10940,N_10521);
and U19424 (N_19424,N_10851,N_11708);
nand U19425 (N_19425,N_11973,N_13919);
nor U19426 (N_19426,N_11992,N_14082);
or U19427 (N_19427,N_11223,N_14970);
and U19428 (N_19428,N_13571,N_13797);
or U19429 (N_19429,N_14298,N_11499);
and U19430 (N_19430,N_11810,N_10395);
and U19431 (N_19431,N_14540,N_14432);
nor U19432 (N_19432,N_10941,N_14919);
nand U19433 (N_19433,N_14080,N_14947);
or U19434 (N_19434,N_12314,N_11082);
nor U19435 (N_19435,N_10709,N_14962);
nor U19436 (N_19436,N_12724,N_13195);
nor U19437 (N_19437,N_14616,N_12861);
nor U19438 (N_19438,N_10032,N_12303);
nand U19439 (N_19439,N_12383,N_10495);
or U19440 (N_19440,N_14001,N_11098);
and U19441 (N_19441,N_11615,N_12008);
nand U19442 (N_19442,N_12519,N_14822);
nand U19443 (N_19443,N_10228,N_10119);
nand U19444 (N_19444,N_14876,N_13221);
nand U19445 (N_19445,N_12007,N_10195);
or U19446 (N_19446,N_10871,N_10879);
or U19447 (N_19447,N_10645,N_14473);
and U19448 (N_19448,N_11005,N_10397);
xor U19449 (N_19449,N_11862,N_14787);
and U19450 (N_19450,N_11051,N_13822);
nor U19451 (N_19451,N_12917,N_10930);
nand U19452 (N_19452,N_10109,N_13188);
xnor U19453 (N_19453,N_14238,N_10436);
and U19454 (N_19454,N_12598,N_12914);
xor U19455 (N_19455,N_12032,N_13272);
and U19456 (N_19456,N_12530,N_10010);
or U19457 (N_19457,N_12259,N_11200);
nor U19458 (N_19458,N_10695,N_14375);
nand U19459 (N_19459,N_12712,N_12070);
and U19460 (N_19460,N_13709,N_13823);
and U19461 (N_19461,N_14465,N_14856);
and U19462 (N_19462,N_11312,N_13485);
nand U19463 (N_19463,N_13464,N_14534);
nor U19464 (N_19464,N_13982,N_11131);
xor U19465 (N_19465,N_10231,N_13011);
or U19466 (N_19466,N_14421,N_13614);
or U19467 (N_19467,N_14955,N_10280);
nor U19468 (N_19468,N_11380,N_13743);
and U19469 (N_19469,N_14202,N_11431);
nand U19470 (N_19470,N_13399,N_14228);
nor U19471 (N_19471,N_14719,N_10164);
and U19472 (N_19472,N_13201,N_12088);
or U19473 (N_19473,N_10729,N_13472);
nor U19474 (N_19474,N_11559,N_10204);
or U19475 (N_19475,N_12529,N_14849);
nand U19476 (N_19476,N_13174,N_13113);
nor U19477 (N_19477,N_10419,N_11699);
or U19478 (N_19478,N_12516,N_11205);
and U19479 (N_19479,N_10759,N_11574);
nand U19480 (N_19480,N_13166,N_14416);
nor U19481 (N_19481,N_14899,N_14160);
nand U19482 (N_19482,N_10781,N_10032);
nand U19483 (N_19483,N_12050,N_13816);
or U19484 (N_19484,N_14936,N_12643);
or U19485 (N_19485,N_14955,N_10909);
nand U19486 (N_19486,N_14381,N_11331);
and U19487 (N_19487,N_11081,N_13552);
nor U19488 (N_19488,N_13940,N_10941);
nor U19489 (N_19489,N_13478,N_13847);
nand U19490 (N_19490,N_12149,N_13697);
or U19491 (N_19491,N_11008,N_13935);
nand U19492 (N_19492,N_13629,N_10788);
nand U19493 (N_19493,N_10902,N_14651);
and U19494 (N_19494,N_12323,N_10664);
nand U19495 (N_19495,N_12141,N_10162);
xnor U19496 (N_19496,N_12173,N_13480);
nand U19497 (N_19497,N_10669,N_14029);
nand U19498 (N_19498,N_14551,N_14267);
xnor U19499 (N_19499,N_14416,N_13226);
nand U19500 (N_19500,N_14753,N_10034);
nor U19501 (N_19501,N_11158,N_11173);
or U19502 (N_19502,N_13100,N_14028);
nor U19503 (N_19503,N_14907,N_12112);
and U19504 (N_19504,N_12672,N_13988);
and U19505 (N_19505,N_13734,N_13053);
or U19506 (N_19506,N_12272,N_12458);
nand U19507 (N_19507,N_14777,N_11419);
nor U19508 (N_19508,N_12292,N_11307);
nor U19509 (N_19509,N_14356,N_13083);
nand U19510 (N_19510,N_13244,N_12170);
or U19511 (N_19511,N_12708,N_11960);
and U19512 (N_19512,N_14139,N_13343);
nor U19513 (N_19513,N_14182,N_11572);
and U19514 (N_19514,N_13855,N_12642);
and U19515 (N_19515,N_12750,N_12708);
and U19516 (N_19516,N_13387,N_11941);
nand U19517 (N_19517,N_10118,N_10256);
nand U19518 (N_19518,N_12098,N_12951);
or U19519 (N_19519,N_11293,N_13696);
or U19520 (N_19520,N_11191,N_14252);
nand U19521 (N_19521,N_12340,N_12880);
nor U19522 (N_19522,N_10806,N_10082);
nand U19523 (N_19523,N_11780,N_13423);
nor U19524 (N_19524,N_10516,N_11132);
or U19525 (N_19525,N_10190,N_14140);
nor U19526 (N_19526,N_10012,N_10173);
or U19527 (N_19527,N_11657,N_12505);
nor U19528 (N_19528,N_10716,N_12000);
nand U19529 (N_19529,N_10837,N_14825);
or U19530 (N_19530,N_11603,N_11051);
nand U19531 (N_19531,N_10835,N_14157);
or U19532 (N_19532,N_13212,N_12652);
or U19533 (N_19533,N_10228,N_10441);
nand U19534 (N_19534,N_12033,N_13882);
nand U19535 (N_19535,N_13269,N_13717);
nand U19536 (N_19536,N_12943,N_12275);
nand U19537 (N_19537,N_13492,N_12367);
or U19538 (N_19538,N_14230,N_14644);
nand U19539 (N_19539,N_14581,N_10729);
nor U19540 (N_19540,N_12580,N_10731);
nor U19541 (N_19541,N_14708,N_13417);
or U19542 (N_19542,N_11981,N_12010);
and U19543 (N_19543,N_13916,N_13915);
and U19544 (N_19544,N_12820,N_12242);
nand U19545 (N_19545,N_12532,N_12983);
and U19546 (N_19546,N_10243,N_14464);
nor U19547 (N_19547,N_10274,N_14165);
or U19548 (N_19548,N_14259,N_11366);
nor U19549 (N_19549,N_12173,N_13380);
nand U19550 (N_19550,N_13205,N_14378);
nor U19551 (N_19551,N_11405,N_11778);
nand U19552 (N_19552,N_11667,N_13951);
nand U19553 (N_19553,N_12958,N_11307);
and U19554 (N_19554,N_12882,N_12169);
or U19555 (N_19555,N_10298,N_11600);
nand U19556 (N_19556,N_14096,N_12777);
nand U19557 (N_19557,N_12506,N_11897);
or U19558 (N_19558,N_12602,N_12322);
nor U19559 (N_19559,N_11825,N_10801);
and U19560 (N_19560,N_13112,N_10040);
and U19561 (N_19561,N_12847,N_10551);
and U19562 (N_19562,N_13206,N_12931);
and U19563 (N_19563,N_11782,N_10547);
and U19564 (N_19564,N_14870,N_13274);
or U19565 (N_19565,N_12440,N_14438);
nor U19566 (N_19566,N_14322,N_11781);
and U19567 (N_19567,N_14255,N_10373);
nand U19568 (N_19568,N_10082,N_14647);
nor U19569 (N_19569,N_14185,N_14271);
nand U19570 (N_19570,N_12691,N_13127);
or U19571 (N_19571,N_10479,N_14706);
and U19572 (N_19572,N_12108,N_13405);
nor U19573 (N_19573,N_10612,N_12079);
or U19574 (N_19574,N_14541,N_11351);
and U19575 (N_19575,N_14749,N_12325);
or U19576 (N_19576,N_11951,N_11926);
or U19577 (N_19577,N_12659,N_10872);
or U19578 (N_19578,N_10602,N_12048);
xnor U19579 (N_19579,N_12066,N_11441);
nor U19580 (N_19580,N_14253,N_10728);
nand U19581 (N_19581,N_14564,N_10806);
xor U19582 (N_19582,N_10020,N_10080);
nor U19583 (N_19583,N_11885,N_11556);
nand U19584 (N_19584,N_11327,N_10764);
nand U19585 (N_19585,N_10824,N_11286);
nand U19586 (N_19586,N_14509,N_12276);
nor U19587 (N_19587,N_10664,N_12995);
nand U19588 (N_19588,N_11031,N_10616);
nand U19589 (N_19589,N_13022,N_10220);
nand U19590 (N_19590,N_11600,N_12107);
and U19591 (N_19591,N_12735,N_13478);
nor U19592 (N_19592,N_11471,N_12709);
nand U19593 (N_19593,N_12085,N_13461);
or U19594 (N_19594,N_11709,N_10554);
or U19595 (N_19595,N_12320,N_12975);
nand U19596 (N_19596,N_12731,N_13897);
nand U19597 (N_19597,N_12479,N_12183);
and U19598 (N_19598,N_14676,N_14612);
or U19599 (N_19599,N_13594,N_12704);
nor U19600 (N_19600,N_10461,N_13630);
and U19601 (N_19601,N_14237,N_13313);
nor U19602 (N_19602,N_10372,N_12622);
or U19603 (N_19603,N_14502,N_13305);
nor U19604 (N_19604,N_11783,N_12925);
nor U19605 (N_19605,N_12538,N_11313);
and U19606 (N_19606,N_10529,N_11126);
or U19607 (N_19607,N_10103,N_11641);
and U19608 (N_19608,N_13683,N_10239);
nand U19609 (N_19609,N_14011,N_12683);
or U19610 (N_19610,N_14672,N_12253);
nor U19611 (N_19611,N_11650,N_14459);
xnor U19612 (N_19612,N_10572,N_11283);
nand U19613 (N_19613,N_12212,N_13366);
nand U19614 (N_19614,N_14741,N_11994);
and U19615 (N_19615,N_14166,N_11699);
nor U19616 (N_19616,N_12804,N_10431);
nor U19617 (N_19617,N_14214,N_11953);
and U19618 (N_19618,N_13086,N_10366);
nand U19619 (N_19619,N_13195,N_14205);
nor U19620 (N_19620,N_10519,N_13492);
and U19621 (N_19621,N_14881,N_11664);
nand U19622 (N_19622,N_13040,N_12929);
nand U19623 (N_19623,N_10102,N_13390);
and U19624 (N_19624,N_14169,N_13726);
or U19625 (N_19625,N_11145,N_11147);
nand U19626 (N_19626,N_14882,N_14948);
or U19627 (N_19627,N_13746,N_14419);
nor U19628 (N_19628,N_10000,N_12496);
nand U19629 (N_19629,N_12748,N_10972);
and U19630 (N_19630,N_14268,N_11902);
nor U19631 (N_19631,N_13649,N_10657);
or U19632 (N_19632,N_13387,N_11164);
and U19633 (N_19633,N_14423,N_14371);
or U19634 (N_19634,N_10087,N_10034);
nand U19635 (N_19635,N_13161,N_11146);
nor U19636 (N_19636,N_11707,N_10457);
nor U19637 (N_19637,N_11775,N_11308);
or U19638 (N_19638,N_13084,N_12158);
nand U19639 (N_19639,N_12605,N_12542);
nand U19640 (N_19640,N_11040,N_13351);
nand U19641 (N_19641,N_11454,N_14397);
nor U19642 (N_19642,N_13627,N_13575);
nand U19643 (N_19643,N_12517,N_11002);
nand U19644 (N_19644,N_13774,N_11315);
nor U19645 (N_19645,N_12547,N_13704);
nand U19646 (N_19646,N_13110,N_14281);
or U19647 (N_19647,N_12583,N_14071);
nand U19648 (N_19648,N_13335,N_14785);
xor U19649 (N_19649,N_11549,N_13452);
nand U19650 (N_19650,N_14901,N_13901);
nand U19651 (N_19651,N_11630,N_11316);
nand U19652 (N_19652,N_14889,N_14145);
nor U19653 (N_19653,N_13480,N_13240);
nand U19654 (N_19654,N_13443,N_14796);
nor U19655 (N_19655,N_11126,N_14032);
nor U19656 (N_19656,N_13536,N_11090);
or U19657 (N_19657,N_10544,N_14555);
or U19658 (N_19658,N_10694,N_14957);
and U19659 (N_19659,N_14273,N_13166);
nand U19660 (N_19660,N_13334,N_14254);
nor U19661 (N_19661,N_11559,N_13491);
or U19662 (N_19662,N_14364,N_11004);
nor U19663 (N_19663,N_13003,N_14056);
nand U19664 (N_19664,N_10675,N_14766);
nand U19665 (N_19665,N_14235,N_13738);
nor U19666 (N_19666,N_14641,N_13254);
or U19667 (N_19667,N_12103,N_12800);
or U19668 (N_19668,N_13730,N_10969);
or U19669 (N_19669,N_11391,N_14511);
nand U19670 (N_19670,N_13084,N_10215);
and U19671 (N_19671,N_10241,N_10973);
or U19672 (N_19672,N_14270,N_10207);
and U19673 (N_19673,N_14026,N_13779);
nand U19674 (N_19674,N_13152,N_10676);
or U19675 (N_19675,N_11211,N_10429);
nand U19676 (N_19676,N_10360,N_13681);
or U19677 (N_19677,N_13655,N_13158);
nand U19678 (N_19678,N_11505,N_14479);
nor U19679 (N_19679,N_11370,N_11746);
and U19680 (N_19680,N_11016,N_13975);
and U19681 (N_19681,N_11466,N_13944);
or U19682 (N_19682,N_12443,N_10843);
or U19683 (N_19683,N_13387,N_10886);
nor U19684 (N_19684,N_13077,N_12435);
nor U19685 (N_19685,N_14150,N_13320);
or U19686 (N_19686,N_14979,N_14507);
nand U19687 (N_19687,N_11091,N_14588);
nand U19688 (N_19688,N_13295,N_11716);
xnor U19689 (N_19689,N_11008,N_14498);
and U19690 (N_19690,N_14878,N_14566);
or U19691 (N_19691,N_13656,N_12260);
nor U19692 (N_19692,N_14694,N_11368);
nand U19693 (N_19693,N_14829,N_10078);
nor U19694 (N_19694,N_14296,N_10463);
or U19695 (N_19695,N_13102,N_12509);
nand U19696 (N_19696,N_10473,N_12869);
or U19697 (N_19697,N_14821,N_10280);
nand U19698 (N_19698,N_11300,N_12238);
or U19699 (N_19699,N_10602,N_10961);
nand U19700 (N_19700,N_13697,N_14709);
nand U19701 (N_19701,N_13757,N_14567);
nor U19702 (N_19702,N_14100,N_11289);
nor U19703 (N_19703,N_13391,N_10084);
or U19704 (N_19704,N_12805,N_11301);
nand U19705 (N_19705,N_11623,N_12213);
or U19706 (N_19706,N_13238,N_13924);
nor U19707 (N_19707,N_12390,N_13414);
and U19708 (N_19708,N_11405,N_14472);
or U19709 (N_19709,N_10782,N_13969);
nand U19710 (N_19710,N_11528,N_13345);
and U19711 (N_19711,N_10356,N_14529);
xnor U19712 (N_19712,N_12290,N_10970);
nor U19713 (N_19713,N_14319,N_14145);
nand U19714 (N_19714,N_13654,N_13379);
and U19715 (N_19715,N_12488,N_12085);
or U19716 (N_19716,N_10057,N_10260);
and U19717 (N_19717,N_13998,N_10423);
xnor U19718 (N_19718,N_14506,N_12480);
nand U19719 (N_19719,N_12536,N_12407);
and U19720 (N_19720,N_10177,N_12945);
nor U19721 (N_19721,N_11690,N_10875);
nor U19722 (N_19722,N_11833,N_10618);
and U19723 (N_19723,N_12534,N_12593);
or U19724 (N_19724,N_13333,N_10050);
or U19725 (N_19725,N_11153,N_13494);
and U19726 (N_19726,N_14557,N_11057);
and U19727 (N_19727,N_13561,N_14614);
nor U19728 (N_19728,N_10246,N_11967);
nand U19729 (N_19729,N_12608,N_14181);
and U19730 (N_19730,N_10580,N_12286);
or U19731 (N_19731,N_11709,N_12964);
nor U19732 (N_19732,N_14447,N_14086);
and U19733 (N_19733,N_14771,N_10632);
nor U19734 (N_19734,N_11655,N_12020);
and U19735 (N_19735,N_11283,N_14596);
and U19736 (N_19736,N_13773,N_13068);
nand U19737 (N_19737,N_14481,N_11108);
xnor U19738 (N_19738,N_11789,N_10236);
and U19739 (N_19739,N_12606,N_12833);
and U19740 (N_19740,N_11720,N_13451);
and U19741 (N_19741,N_13957,N_10252);
and U19742 (N_19742,N_11930,N_14430);
or U19743 (N_19743,N_12904,N_12479);
or U19744 (N_19744,N_13020,N_11367);
nor U19745 (N_19745,N_14701,N_14569);
nor U19746 (N_19746,N_13098,N_12576);
or U19747 (N_19747,N_13655,N_11969);
and U19748 (N_19748,N_10661,N_10625);
nand U19749 (N_19749,N_11407,N_11825);
or U19750 (N_19750,N_12109,N_10526);
nand U19751 (N_19751,N_11603,N_10468);
nand U19752 (N_19752,N_11513,N_10615);
nor U19753 (N_19753,N_12974,N_13910);
nor U19754 (N_19754,N_11969,N_10342);
nor U19755 (N_19755,N_10546,N_13970);
and U19756 (N_19756,N_10839,N_13123);
nand U19757 (N_19757,N_14934,N_13839);
nand U19758 (N_19758,N_12569,N_12618);
nand U19759 (N_19759,N_12224,N_12395);
nand U19760 (N_19760,N_11987,N_14284);
xor U19761 (N_19761,N_12701,N_14291);
nand U19762 (N_19762,N_10605,N_10587);
nand U19763 (N_19763,N_14663,N_10476);
nor U19764 (N_19764,N_12896,N_12347);
and U19765 (N_19765,N_14599,N_12406);
or U19766 (N_19766,N_13275,N_12990);
nor U19767 (N_19767,N_10721,N_13320);
or U19768 (N_19768,N_11418,N_13809);
and U19769 (N_19769,N_14784,N_11583);
nor U19770 (N_19770,N_13319,N_11874);
and U19771 (N_19771,N_14756,N_12456);
and U19772 (N_19772,N_14994,N_13566);
and U19773 (N_19773,N_10620,N_10046);
and U19774 (N_19774,N_13474,N_10232);
nor U19775 (N_19775,N_10695,N_10497);
or U19776 (N_19776,N_11354,N_12202);
or U19777 (N_19777,N_14044,N_13041);
or U19778 (N_19778,N_14110,N_13982);
nor U19779 (N_19779,N_12452,N_11676);
or U19780 (N_19780,N_12023,N_10974);
and U19781 (N_19781,N_10530,N_14752);
or U19782 (N_19782,N_14178,N_14698);
nand U19783 (N_19783,N_12915,N_11941);
and U19784 (N_19784,N_11021,N_10232);
and U19785 (N_19785,N_13894,N_14942);
xor U19786 (N_19786,N_13383,N_14430);
nor U19787 (N_19787,N_11610,N_12242);
nand U19788 (N_19788,N_10303,N_13709);
or U19789 (N_19789,N_13879,N_14195);
nor U19790 (N_19790,N_13799,N_10621);
or U19791 (N_19791,N_12829,N_11702);
nor U19792 (N_19792,N_12944,N_11344);
nor U19793 (N_19793,N_13888,N_12151);
and U19794 (N_19794,N_10864,N_14031);
nand U19795 (N_19795,N_11919,N_13539);
nand U19796 (N_19796,N_13548,N_12446);
nand U19797 (N_19797,N_11611,N_11761);
nor U19798 (N_19798,N_12675,N_13483);
nand U19799 (N_19799,N_11684,N_10162);
nor U19800 (N_19800,N_12514,N_14456);
nand U19801 (N_19801,N_14455,N_13633);
or U19802 (N_19802,N_11545,N_11730);
nand U19803 (N_19803,N_10987,N_12514);
nand U19804 (N_19804,N_11404,N_10998);
nand U19805 (N_19805,N_13948,N_10868);
nor U19806 (N_19806,N_13472,N_11346);
nor U19807 (N_19807,N_13154,N_10028);
and U19808 (N_19808,N_12113,N_11812);
nand U19809 (N_19809,N_11468,N_11158);
or U19810 (N_19810,N_14974,N_11946);
and U19811 (N_19811,N_12118,N_14623);
nand U19812 (N_19812,N_13022,N_13608);
and U19813 (N_19813,N_10420,N_14800);
and U19814 (N_19814,N_14179,N_12694);
or U19815 (N_19815,N_14356,N_12178);
and U19816 (N_19816,N_13331,N_13833);
nand U19817 (N_19817,N_14258,N_14947);
and U19818 (N_19818,N_12792,N_10382);
nor U19819 (N_19819,N_10210,N_14882);
nor U19820 (N_19820,N_11046,N_11576);
or U19821 (N_19821,N_12629,N_11231);
nor U19822 (N_19822,N_12874,N_11824);
and U19823 (N_19823,N_11855,N_10473);
and U19824 (N_19824,N_12104,N_13810);
and U19825 (N_19825,N_14556,N_13722);
or U19826 (N_19826,N_14227,N_11796);
nor U19827 (N_19827,N_12521,N_14532);
and U19828 (N_19828,N_14576,N_13849);
nand U19829 (N_19829,N_14603,N_13019);
nor U19830 (N_19830,N_13402,N_10154);
and U19831 (N_19831,N_11796,N_14133);
nand U19832 (N_19832,N_13576,N_14349);
nand U19833 (N_19833,N_10658,N_13026);
and U19834 (N_19834,N_11908,N_13121);
or U19835 (N_19835,N_10138,N_13606);
xor U19836 (N_19836,N_12960,N_10031);
nor U19837 (N_19837,N_14977,N_12081);
nand U19838 (N_19838,N_14038,N_14209);
or U19839 (N_19839,N_14674,N_10913);
and U19840 (N_19840,N_11152,N_13006);
and U19841 (N_19841,N_13950,N_11489);
or U19842 (N_19842,N_10002,N_13715);
nand U19843 (N_19843,N_12648,N_12580);
and U19844 (N_19844,N_10033,N_12869);
and U19845 (N_19845,N_11626,N_10473);
nor U19846 (N_19846,N_14898,N_11863);
nand U19847 (N_19847,N_14218,N_13503);
nor U19848 (N_19848,N_10071,N_14657);
and U19849 (N_19849,N_13478,N_10452);
or U19850 (N_19850,N_13280,N_11780);
or U19851 (N_19851,N_12826,N_11499);
nor U19852 (N_19852,N_10668,N_10713);
nor U19853 (N_19853,N_12737,N_11627);
or U19854 (N_19854,N_11663,N_14606);
nand U19855 (N_19855,N_11967,N_12739);
nor U19856 (N_19856,N_10659,N_13766);
nand U19857 (N_19857,N_12040,N_11191);
nor U19858 (N_19858,N_11712,N_12142);
and U19859 (N_19859,N_11109,N_12993);
nor U19860 (N_19860,N_14160,N_14605);
and U19861 (N_19861,N_11281,N_11621);
or U19862 (N_19862,N_12422,N_11031);
nand U19863 (N_19863,N_14886,N_12447);
or U19864 (N_19864,N_13026,N_11216);
nor U19865 (N_19865,N_10990,N_11714);
nand U19866 (N_19866,N_11115,N_14123);
and U19867 (N_19867,N_12099,N_11231);
nand U19868 (N_19868,N_12692,N_10979);
or U19869 (N_19869,N_12827,N_12645);
or U19870 (N_19870,N_13111,N_10084);
nor U19871 (N_19871,N_12251,N_14557);
nor U19872 (N_19872,N_14384,N_14414);
and U19873 (N_19873,N_14130,N_13418);
and U19874 (N_19874,N_13498,N_14770);
and U19875 (N_19875,N_14492,N_10152);
nand U19876 (N_19876,N_10259,N_14362);
nand U19877 (N_19877,N_13494,N_14090);
or U19878 (N_19878,N_10896,N_14535);
or U19879 (N_19879,N_13112,N_10014);
nand U19880 (N_19880,N_11553,N_12808);
nor U19881 (N_19881,N_14216,N_14861);
nand U19882 (N_19882,N_14084,N_12073);
or U19883 (N_19883,N_14094,N_13741);
or U19884 (N_19884,N_12572,N_14549);
nand U19885 (N_19885,N_13564,N_12003);
and U19886 (N_19886,N_10760,N_14497);
or U19887 (N_19887,N_10009,N_14816);
nor U19888 (N_19888,N_10640,N_10051);
nor U19889 (N_19889,N_12998,N_12696);
nand U19890 (N_19890,N_13092,N_10446);
nor U19891 (N_19891,N_12040,N_10642);
nor U19892 (N_19892,N_13631,N_12324);
nor U19893 (N_19893,N_10142,N_11632);
and U19894 (N_19894,N_14989,N_13927);
and U19895 (N_19895,N_10067,N_11472);
nand U19896 (N_19896,N_11604,N_13773);
or U19897 (N_19897,N_11934,N_12258);
and U19898 (N_19898,N_10902,N_14399);
or U19899 (N_19899,N_12340,N_11307);
and U19900 (N_19900,N_10257,N_14145);
nand U19901 (N_19901,N_13330,N_12117);
or U19902 (N_19902,N_10057,N_12268);
or U19903 (N_19903,N_12888,N_11529);
or U19904 (N_19904,N_10657,N_11683);
nor U19905 (N_19905,N_13588,N_14901);
and U19906 (N_19906,N_12830,N_11961);
and U19907 (N_19907,N_14370,N_14203);
nor U19908 (N_19908,N_14708,N_10513);
and U19909 (N_19909,N_12425,N_12976);
or U19910 (N_19910,N_11640,N_10217);
nand U19911 (N_19911,N_13122,N_14362);
and U19912 (N_19912,N_10485,N_14698);
and U19913 (N_19913,N_14440,N_14830);
xor U19914 (N_19914,N_10957,N_14325);
nand U19915 (N_19915,N_14315,N_14453);
nand U19916 (N_19916,N_14620,N_12377);
nand U19917 (N_19917,N_14322,N_12726);
nand U19918 (N_19918,N_13874,N_10559);
nand U19919 (N_19919,N_10110,N_10263);
and U19920 (N_19920,N_12841,N_14503);
nand U19921 (N_19921,N_14921,N_10007);
nand U19922 (N_19922,N_11417,N_13924);
nor U19923 (N_19923,N_11225,N_13894);
nor U19924 (N_19924,N_13601,N_13003);
and U19925 (N_19925,N_14586,N_11922);
and U19926 (N_19926,N_13012,N_10432);
nor U19927 (N_19927,N_12517,N_11183);
nor U19928 (N_19928,N_10406,N_13599);
nor U19929 (N_19929,N_14116,N_12529);
nor U19930 (N_19930,N_10134,N_11881);
nand U19931 (N_19931,N_13337,N_13982);
nor U19932 (N_19932,N_11882,N_11756);
and U19933 (N_19933,N_12564,N_13895);
nor U19934 (N_19934,N_12824,N_11126);
nand U19935 (N_19935,N_14265,N_12833);
and U19936 (N_19936,N_13553,N_11270);
or U19937 (N_19937,N_11540,N_12909);
nor U19938 (N_19938,N_12251,N_12744);
nor U19939 (N_19939,N_12259,N_10755);
and U19940 (N_19940,N_11854,N_10766);
nor U19941 (N_19941,N_12112,N_13465);
or U19942 (N_19942,N_12632,N_14933);
nor U19943 (N_19943,N_11295,N_12594);
and U19944 (N_19944,N_14680,N_11349);
xnor U19945 (N_19945,N_10051,N_12892);
nor U19946 (N_19946,N_11222,N_14936);
nand U19947 (N_19947,N_12332,N_12117);
and U19948 (N_19948,N_10500,N_10424);
and U19949 (N_19949,N_14185,N_10500);
nor U19950 (N_19950,N_11818,N_14721);
nand U19951 (N_19951,N_12041,N_12433);
or U19952 (N_19952,N_11754,N_11375);
and U19953 (N_19953,N_14146,N_14410);
or U19954 (N_19954,N_13849,N_12604);
or U19955 (N_19955,N_14373,N_10691);
and U19956 (N_19956,N_10589,N_13515);
or U19957 (N_19957,N_13493,N_10930);
nand U19958 (N_19958,N_11936,N_14583);
nor U19959 (N_19959,N_13124,N_10445);
nor U19960 (N_19960,N_13216,N_12904);
nor U19961 (N_19961,N_10699,N_10075);
or U19962 (N_19962,N_11082,N_12996);
and U19963 (N_19963,N_12001,N_14067);
or U19964 (N_19964,N_11184,N_10686);
nand U19965 (N_19965,N_13058,N_12782);
and U19966 (N_19966,N_11543,N_13138);
and U19967 (N_19967,N_13497,N_10488);
or U19968 (N_19968,N_11221,N_11363);
or U19969 (N_19969,N_13189,N_14898);
or U19970 (N_19970,N_14633,N_13710);
nor U19971 (N_19971,N_12847,N_13662);
nor U19972 (N_19972,N_10564,N_14182);
and U19973 (N_19973,N_13634,N_13952);
and U19974 (N_19974,N_14006,N_12851);
nor U19975 (N_19975,N_11384,N_14734);
nor U19976 (N_19976,N_14762,N_10049);
nand U19977 (N_19977,N_12948,N_11235);
xnor U19978 (N_19978,N_10942,N_11975);
nand U19979 (N_19979,N_10457,N_12370);
nor U19980 (N_19980,N_14613,N_13424);
nand U19981 (N_19981,N_12285,N_12303);
and U19982 (N_19982,N_12966,N_12285);
and U19983 (N_19983,N_11815,N_13506);
nand U19984 (N_19984,N_14878,N_11788);
nor U19985 (N_19985,N_12767,N_12155);
and U19986 (N_19986,N_11334,N_12949);
nand U19987 (N_19987,N_14727,N_10054);
or U19988 (N_19988,N_10823,N_14900);
or U19989 (N_19989,N_13787,N_14539);
nor U19990 (N_19990,N_11551,N_14256);
and U19991 (N_19991,N_10163,N_10798);
nand U19992 (N_19992,N_11252,N_12109);
nand U19993 (N_19993,N_11885,N_13683);
nand U19994 (N_19994,N_10032,N_13603);
or U19995 (N_19995,N_14965,N_11517);
or U19996 (N_19996,N_11745,N_14480);
or U19997 (N_19997,N_11946,N_13873);
and U19998 (N_19998,N_13640,N_10571);
nor U19999 (N_19999,N_13121,N_10659);
nor U20000 (N_20000,N_16897,N_16603);
nand U20001 (N_20001,N_19756,N_17754);
nand U20002 (N_20002,N_18946,N_19507);
nor U20003 (N_20003,N_16142,N_15389);
nand U20004 (N_20004,N_15051,N_16321);
nor U20005 (N_20005,N_17458,N_17420);
and U20006 (N_20006,N_19172,N_19808);
and U20007 (N_20007,N_19214,N_17663);
nand U20008 (N_20008,N_18953,N_18990);
nor U20009 (N_20009,N_18680,N_19260);
nand U20010 (N_20010,N_16487,N_18863);
and U20011 (N_20011,N_17189,N_16247);
or U20012 (N_20012,N_16550,N_15178);
nand U20013 (N_20013,N_15638,N_19953);
nor U20014 (N_20014,N_18438,N_17201);
or U20015 (N_20015,N_15843,N_15143);
nor U20016 (N_20016,N_15191,N_18021);
and U20017 (N_20017,N_15575,N_15580);
or U20018 (N_20018,N_18419,N_16010);
and U20019 (N_20019,N_17071,N_16392);
nor U20020 (N_20020,N_16264,N_18724);
or U20021 (N_20021,N_19177,N_17440);
nor U20022 (N_20022,N_17709,N_16628);
nor U20023 (N_20023,N_19150,N_19168);
or U20024 (N_20024,N_15342,N_16663);
nand U20025 (N_20025,N_17771,N_18828);
nor U20026 (N_20026,N_19893,N_18456);
nor U20027 (N_20027,N_17051,N_18660);
and U20028 (N_20028,N_15744,N_19544);
nor U20029 (N_20029,N_17326,N_15637);
and U20030 (N_20030,N_15470,N_15232);
nand U20031 (N_20031,N_16342,N_15493);
and U20032 (N_20032,N_15578,N_15210);
nand U20033 (N_20033,N_17827,N_17788);
and U20034 (N_20034,N_15491,N_15540);
nor U20035 (N_20035,N_15416,N_16528);
and U20036 (N_20036,N_15725,N_17441);
nand U20037 (N_20037,N_16749,N_16648);
nand U20038 (N_20038,N_18499,N_19300);
and U20039 (N_20039,N_15648,N_19023);
nor U20040 (N_20040,N_17453,N_15900);
and U20041 (N_20041,N_18309,N_19415);
or U20042 (N_20042,N_19906,N_16845);
nor U20043 (N_20043,N_16959,N_18855);
nand U20044 (N_20044,N_18501,N_19989);
and U20045 (N_20045,N_17579,N_15642);
and U20046 (N_20046,N_15390,N_17977);
or U20047 (N_20047,N_16598,N_17597);
xnor U20048 (N_20048,N_18218,N_19597);
and U20049 (N_20049,N_18704,N_15698);
and U20050 (N_20050,N_15167,N_18697);
or U20051 (N_20051,N_18511,N_16837);
and U20052 (N_20052,N_19620,N_17344);
or U20053 (N_20053,N_18350,N_16785);
nor U20054 (N_20054,N_19262,N_17630);
nand U20055 (N_20055,N_18577,N_16839);
and U20056 (N_20056,N_18343,N_18269);
nand U20057 (N_20057,N_15741,N_17002);
and U20058 (N_20058,N_18742,N_15186);
nor U20059 (N_20059,N_18100,N_18341);
nor U20060 (N_20060,N_18002,N_16049);
nor U20061 (N_20061,N_17947,N_16522);
nor U20062 (N_20062,N_17199,N_15304);
nand U20063 (N_20063,N_16701,N_18125);
and U20064 (N_20064,N_15706,N_19396);
nand U20065 (N_20065,N_15711,N_15433);
or U20066 (N_20066,N_16163,N_16120);
and U20067 (N_20067,N_18722,N_18398);
nor U20068 (N_20068,N_17048,N_15631);
and U20069 (N_20069,N_19083,N_19664);
nand U20070 (N_20070,N_16606,N_15738);
nand U20071 (N_20071,N_17164,N_16587);
nand U20072 (N_20072,N_19929,N_16104);
nand U20073 (N_20073,N_18214,N_15983);
or U20074 (N_20074,N_19435,N_16003);
or U20075 (N_20075,N_19277,N_16161);
or U20076 (N_20076,N_19385,N_15632);
nor U20077 (N_20077,N_19274,N_17196);
or U20078 (N_20078,N_16995,N_19275);
nand U20079 (N_20079,N_18486,N_17726);
nand U20080 (N_20080,N_18320,N_17803);
nand U20081 (N_20081,N_17262,N_18594);
or U20082 (N_20082,N_15244,N_17938);
or U20083 (N_20083,N_19460,N_19139);
nand U20084 (N_20084,N_15996,N_15779);
nor U20085 (N_20085,N_18330,N_15503);
nand U20086 (N_20086,N_15670,N_16886);
xor U20087 (N_20087,N_18378,N_15130);
nor U20088 (N_20088,N_18851,N_15974);
or U20089 (N_20089,N_15356,N_15168);
nor U20090 (N_20090,N_19542,N_17101);
nor U20091 (N_20091,N_18049,N_15514);
and U20092 (N_20092,N_16307,N_17470);
or U20093 (N_20093,N_15241,N_16882);
nor U20094 (N_20094,N_16495,N_19802);
or U20095 (N_20095,N_15700,N_15078);
nand U20096 (N_20096,N_15736,N_15549);
xor U20097 (N_20097,N_19830,N_18224);
or U20098 (N_20098,N_15915,N_18126);
nand U20099 (N_20099,N_16396,N_16071);
nor U20100 (N_20100,N_18063,N_16733);
nand U20101 (N_20101,N_16740,N_19657);
and U20102 (N_20102,N_16731,N_18618);
nor U20103 (N_20103,N_18060,N_16109);
nand U20104 (N_20104,N_19494,N_16772);
nand U20105 (N_20105,N_19676,N_19822);
nor U20106 (N_20106,N_18010,N_19860);
nand U20107 (N_20107,N_18621,N_18368);
nand U20108 (N_20108,N_18839,N_16437);
and U20109 (N_20109,N_18603,N_15404);
and U20110 (N_20110,N_15234,N_16544);
and U20111 (N_20111,N_19883,N_19112);
nor U20112 (N_20112,N_15350,N_16240);
and U20113 (N_20113,N_16332,N_19091);
or U20114 (N_20114,N_16282,N_15257);
nor U20115 (N_20115,N_17358,N_16931);
and U20116 (N_20116,N_17775,N_18778);
nor U20117 (N_20117,N_18519,N_17211);
or U20118 (N_20118,N_18717,N_19010);
nor U20119 (N_20119,N_18489,N_18171);
and U20120 (N_20120,N_19726,N_16583);
or U20121 (N_20121,N_19717,N_17077);
nand U20122 (N_20122,N_18169,N_18963);
nand U20123 (N_20123,N_17118,N_18335);
nand U20124 (N_20124,N_17452,N_15786);
nor U20125 (N_20125,N_16400,N_18738);
or U20126 (N_20126,N_17316,N_19965);
and U20127 (N_20127,N_15913,N_16516);
nor U20128 (N_20128,N_15068,N_18260);
nand U20129 (N_20129,N_19486,N_18133);
and U20130 (N_20130,N_19047,N_16903);
nand U20131 (N_20131,N_19932,N_17473);
nand U20132 (N_20132,N_16928,N_16842);
and U20133 (N_20133,N_17427,N_17357);
nand U20134 (N_20134,N_16883,N_18688);
and U20135 (N_20135,N_18151,N_17626);
nand U20136 (N_20136,N_17577,N_17650);
and U20137 (N_20137,N_16929,N_18497);
nor U20138 (N_20138,N_15753,N_17949);
nand U20139 (N_20139,N_18732,N_17106);
or U20140 (N_20140,N_17796,N_18612);
nand U20141 (N_20141,N_16916,N_19825);
and U20142 (N_20142,N_16742,N_15227);
and U20143 (N_20143,N_16686,N_17995);
nand U20144 (N_20144,N_19667,N_17621);
and U20145 (N_20145,N_15897,N_18087);
and U20146 (N_20146,N_18634,N_18979);
xor U20147 (N_20147,N_19182,N_15732);
and U20148 (N_20148,N_18366,N_15319);
or U20149 (N_20149,N_15772,N_15238);
nand U20150 (N_20150,N_15408,N_16153);
and U20151 (N_20151,N_16377,N_16677);
nor U20152 (N_20152,N_16967,N_15102);
nor U20153 (N_20153,N_18464,N_18769);
nor U20154 (N_20154,N_16140,N_19692);
and U20155 (N_20155,N_19059,N_18574);
xnor U20156 (N_20156,N_18162,N_15634);
and U20157 (N_20157,N_17059,N_19062);
nand U20158 (N_20158,N_19517,N_18128);
nor U20159 (N_20159,N_16541,N_19472);
nor U20160 (N_20160,N_18431,N_19768);
nor U20161 (N_20161,N_18195,N_19280);
and U20162 (N_20162,N_17423,N_16422);
and U20163 (N_20163,N_16399,N_17957);
or U20164 (N_20164,N_16117,N_16750);
nand U20165 (N_20165,N_18976,N_17982);
and U20166 (N_20166,N_19180,N_17555);
or U20167 (N_20167,N_18835,N_18869);
nand U20168 (N_20168,N_15170,N_15454);
nor U20169 (N_20169,N_15534,N_18292);
and U20170 (N_20170,N_15361,N_19980);
nand U20171 (N_20171,N_17000,N_16933);
nand U20172 (N_20172,N_19608,N_19555);
nand U20173 (N_20173,N_16179,N_15141);
or U20174 (N_20174,N_15086,N_18716);
and U20175 (N_20175,N_16610,N_19035);
nor U20176 (N_20176,N_18054,N_19071);
and U20177 (N_20177,N_18600,N_15349);
nor U20178 (N_20178,N_16474,N_16937);
nor U20179 (N_20179,N_17162,N_17264);
and U20180 (N_20180,N_18757,N_19367);
nor U20181 (N_20181,N_16769,N_15466);
nand U20182 (N_20182,N_19924,N_15376);
or U20183 (N_20183,N_16015,N_18579);
or U20184 (N_20184,N_18071,N_18116);
and U20185 (N_20185,N_19409,N_15230);
or U20186 (N_20186,N_16857,N_19271);
nand U20187 (N_20187,N_19610,N_17697);
and U20188 (N_20188,N_19225,N_19451);
and U20189 (N_20189,N_15297,N_16484);
nor U20190 (N_20190,N_15633,N_17397);
nor U20191 (N_20191,N_17350,N_19038);
nor U20192 (N_20192,N_16310,N_15508);
xor U20193 (N_20193,N_16314,N_15699);
and U20194 (N_20194,N_19871,N_18545);
nand U20195 (N_20195,N_17964,N_17558);
and U20196 (N_20196,N_17412,N_15708);
or U20197 (N_20197,N_15807,N_16434);
nand U20198 (N_20198,N_17055,N_17599);
nor U20199 (N_20199,N_17031,N_17306);
nand U20200 (N_20200,N_16803,N_15197);
and U20201 (N_20201,N_18585,N_16617);
and U20202 (N_20202,N_17123,N_15194);
or U20203 (N_20203,N_18203,N_18194);
nor U20204 (N_20204,N_18476,N_17224);
and U20205 (N_20205,N_15379,N_16981);
nor U20206 (N_20206,N_19380,N_18105);
or U20207 (N_20207,N_19829,N_16111);
nor U20208 (N_20208,N_15762,N_19884);
nor U20209 (N_20209,N_15710,N_15668);
nand U20210 (N_20210,N_17718,N_17335);
and U20211 (N_20211,N_17645,N_15588);
nor U20212 (N_20212,N_18437,N_19581);
nand U20213 (N_20213,N_16851,N_18198);
and U20214 (N_20214,N_17111,N_15767);
nor U20215 (N_20215,N_19081,N_16242);
or U20216 (N_20216,N_15105,N_16246);
or U20217 (N_20217,N_17843,N_15850);
nor U20218 (N_20218,N_16483,N_15008);
xor U20219 (N_20219,N_18432,N_18975);
xnor U20220 (N_20220,N_19371,N_18524);
xor U20221 (N_20221,N_17083,N_15801);
and U20222 (N_20222,N_15485,N_17873);
and U20223 (N_20223,N_19152,N_17741);
nor U20224 (N_20224,N_15997,N_19821);
and U20225 (N_20225,N_18560,N_15198);
or U20226 (N_20226,N_15340,N_17755);
or U20227 (N_20227,N_16124,N_19589);
and U20228 (N_20228,N_19431,N_17837);
nor U20229 (N_20229,N_15478,N_16556);
nor U20230 (N_20230,N_16002,N_15891);
or U20231 (N_20231,N_19552,N_15332);
or U20232 (N_20232,N_18472,N_19588);
and U20233 (N_20233,N_15598,N_17219);
nor U20234 (N_20234,N_16275,N_17328);
and U20235 (N_20235,N_18303,N_19702);
or U20236 (N_20236,N_15559,N_15107);
or U20237 (N_20237,N_17618,N_16013);
nand U20238 (N_20238,N_19328,N_18286);
and U20239 (N_20239,N_19587,N_17756);
nand U20240 (N_20240,N_19240,N_19634);
nor U20241 (N_20241,N_16739,N_18760);
and U20242 (N_20242,N_16129,N_18725);
nand U20243 (N_20243,N_19524,N_19499);
nor U20244 (N_20244,N_18905,N_19575);
and U20245 (N_20245,N_16789,N_17005);
or U20246 (N_20246,N_17041,N_18488);
nand U20247 (N_20247,N_19392,N_15576);
or U20248 (N_20248,N_15098,N_16496);
and U20249 (N_20249,N_18097,N_19921);
nand U20250 (N_20250,N_15993,N_17682);
or U20251 (N_20251,N_17578,N_19852);
nor U20252 (N_20252,N_19327,N_17327);
and U20253 (N_20253,N_19074,N_16871);
nor U20254 (N_20254,N_16917,N_16426);
nor U20255 (N_20255,N_16472,N_17105);
nor U20256 (N_20256,N_16992,N_19548);
nor U20257 (N_20257,N_17035,N_17978);
or U20258 (N_20258,N_19176,N_17792);
nand U20259 (N_20259,N_18627,N_16118);
nor U20260 (N_20260,N_19843,N_17714);
nor U20261 (N_20261,N_17329,N_15391);
xor U20262 (N_20262,N_17776,N_17027);
and U20263 (N_20263,N_18122,N_16691);
or U20264 (N_20264,N_17824,N_17401);
nor U20265 (N_20265,N_18506,N_19188);
or U20266 (N_20266,N_16308,N_18825);
nand U20267 (N_20267,N_17519,N_19429);
xnor U20268 (N_20268,N_18943,N_19167);
or U20269 (N_20269,N_19354,N_16651);
nand U20270 (N_20270,N_15305,N_16343);
or U20271 (N_20271,N_17475,N_17355);
nor U20272 (N_20272,N_17334,N_17180);
or U20273 (N_20273,N_19316,N_15326);
and U20274 (N_20274,N_15461,N_19463);
nor U20275 (N_20275,N_15872,N_17253);
xor U20276 (N_20276,N_16784,N_15554);
nor U20277 (N_20277,N_16056,N_18756);
nor U20278 (N_20278,N_19868,N_18158);
nor U20279 (N_20279,N_18446,N_15645);
or U20280 (N_20280,N_15392,N_16086);
and U20281 (N_20281,N_15075,N_15854);
nor U20282 (N_20282,N_16862,N_19775);
and U20283 (N_20283,N_16113,N_17376);
or U20284 (N_20284,N_17391,N_16561);
nand U20285 (N_20285,N_15650,N_15149);
and U20286 (N_20286,N_16228,N_18340);
nand U20287 (N_20287,N_17930,N_16034);
nand U20288 (N_20288,N_16480,N_17594);
or U20289 (N_20289,N_17916,N_18935);
or U20290 (N_20290,N_16868,N_15932);
and U20291 (N_20291,N_17851,N_19485);
and U20292 (N_20292,N_18790,N_15084);
or U20293 (N_20293,N_15898,N_16055);
nor U20294 (N_20294,N_17553,N_18983);
and U20295 (N_20295,N_19411,N_18344);
nor U20296 (N_20296,N_15007,N_17394);
nor U20297 (N_20297,N_15264,N_18598);
nand U20298 (N_20298,N_19049,N_19962);
nor U20299 (N_20299,N_18361,N_16637);
nor U20300 (N_20300,N_16913,N_19662);
or U20301 (N_20301,N_15047,N_15337);
nand U20302 (N_20302,N_15286,N_15518);
nor U20303 (N_20303,N_16471,N_16213);
and U20304 (N_20304,N_15074,N_19912);
and U20305 (N_20305,N_19405,N_19397);
and U20306 (N_20306,N_16988,N_19204);
and U20307 (N_20307,N_17396,N_19437);
nor U20308 (N_20308,N_16751,N_16183);
nor U20309 (N_20309,N_18865,N_18710);
nand U20310 (N_20310,N_18146,N_18179);
nor U20311 (N_20311,N_16304,N_19244);
and U20312 (N_20312,N_18744,N_19872);
nand U20313 (N_20313,N_15569,N_17156);
and U20314 (N_20314,N_18373,N_16311);
and U20315 (N_20315,N_18741,N_19901);
xnor U20316 (N_20316,N_17258,N_17375);
and U20317 (N_20317,N_19757,N_17217);
and U20318 (N_20318,N_19844,N_18871);
nor U20319 (N_20319,N_17918,N_19941);
nor U20320 (N_20320,N_19294,N_17929);
nand U20321 (N_20321,N_16378,N_17512);
nor U20322 (N_20322,N_19909,N_17611);
or U20323 (N_20323,N_19820,N_19623);
and U20324 (N_20324,N_19386,N_16538);
or U20325 (N_20325,N_15583,N_15247);
xnor U20326 (N_20326,N_16136,N_16622);
nor U20327 (N_20327,N_18653,N_15283);
and U20328 (N_20328,N_15510,N_15240);
or U20329 (N_20329,N_15482,N_16414);
nor U20330 (N_20330,N_17290,N_15406);
and U20331 (N_20331,N_17887,N_16822);
and U20332 (N_20332,N_19340,N_18925);
and U20333 (N_20333,N_17500,N_18005);
nand U20334 (N_20334,N_17249,N_17974);
or U20335 (N_20335,N_15043,N_18401);
and U20336 (N_20336,N_18689,N_16028);
or U20337 (N_20337,N_16402,N_16572);
and U20338 (N_20338,N_17170,N_18245);
and U20339 (N_20339,N_15511,N_16257);
nor U20340 (N_20340,N_17989,N_19341);
nand U20341 (N_20341,N_17951,N_19573);
nor U20342 (N_20342,N_16288,N_16668);
and U20343 (N_20343,N_16514,N_18568);
and U20344 (N_20344,N_19351,N_16948);
nand U20345 (N_20345,N_16515,N_18413);
nor U20346 (N_20346,N_19858,N_19925);
and U20347 (N_20347,N_18708,N_16766);
nand U20348 (N_20348,N_17994,N_18672);
and U20349 (N_20349,N_17923,N_18699);
nor U20350 (N_20350,N_18069,N_15285);
nand U20351 (N_20351,N_18613,N_17361);
nor U20352 (N_20352,N_19407,N_19426);
nor U20353 (N_20353,N_15312,N_15790);
nor U20354 (N_20354,N_15839,N_18348);
nor U20355 (N_20355,N_16719,N_16756);
nand U20356 (N_20356,N_17914,N_19388);
or U20357 (N_20357,N_17119,N_17572);
nand U20358 (N_20358,N_15348,N_18980);
and U20359 (N_20359,N_15678,N_19361);
nor U20360 (N_20360,N_19052,N_18042);
or U20361 (N_20361,N_19556,N_19253);
nand U20362 (N_20362,N_18940,N_16040);
nand U20363 (N_20363,N_19848,N_19652);
nand U20364 (N_20364,N_19632,N_17360);
nand U20365 (N_20365,N_19835,N_17400);
and U20366 (N_20366,N_15154,N_17346);
or U20367 (N_20367,N_17437,N_18727);
or U20368 (N_20368,N_15934,N_15359);
nand U20369 (N_20369,N_15959,N_18065);
or U20370 (N_20370,N_15172,N_18371);
or U20371 (N_20371,N_15436,N_16976);
or U20372 (N_20372,N_18402,N_15893);
xor U20373 (N_20373,N_16027,N_17785);
and U20374 (N_20374,N_19899,N_16687);
and U20375 (N_20375,N_17115,N_17214);
nor U20376 (N_20376,N_16649,N_15048);
xnor U20377 (N_20377,N_15474,N_15750);
nor U20378 (N_20378,N_16440,N_17582);
xor U20379 (N_20379,N_19973,N_15602);
or U20380 (N_20380,N_15834,N_17542);
and U20381 (N_20381,N_15472,N_17725);
nor U20382 (N_20382,N_19491,N_17471);
or U20383 (N_20383,N_15327,N_19880);
nor U20384 (N_20384,N_15338,N_16860);
and U20385 (N_20385,N_17309,N_17819);
nor U20386 (N_20386,N_16009,N_19892);
and U20387 (N_20387,N_18903,N_19576);
and U20388 (N_20388,N_15689,N_18238);
nor U20389 (N_20389,N_16627,N_18450);
nand U20390 (N_20390,N_15134,N_17457);
and U20391 (N_20391,N_19381,N_15017);
or U20392 (N_20392,N_16272,N_15004);
and U20393 (N_20393,N_17465,N_15148);
or U20394 (N_20394,N_15473,N_16069);
nand U20395 (N_20395,N_18426,N_16464);
nand U20396 (N_20396,N_16918,N_15329);
and U20397 (N_20397,N_19583,N_15352);
and U20398 (N_20398,N_19646,N_19521);
nor U20399 (N_20399,N_18314,N_15477);
nand U20400 (N_20400,N_17940,N_17606);
and U20401 (N_20401,N_19519,N_17409);
or U20402 (N_20402,N_17576,N_16588);
nor U20403 (N_20403,N_19151,N_15147);
or U20404 (N_20404,N_17121,N_15421);
and U20405 (N_20405,N_18817,N_18525);
nand U20406 (N_20406,N_16060,N_15014);
or U20407 (N_20407,N_18392,N_16831);
xnor U20408 (N_20408,N_16497,N_17063);
and U20409 (N_20409,N_18258,N_15617);
or U20410 (N_20410,N_15582,N_18018);
or U20411 (N_20411,N_16297,N_18761);
nand U20412 (N_20412,N_16051,N_15907);
nor U20413 (N_20413,N_16671,N_16797);
and U20414 (N_20414,N_15748,N_15541);
nand U20415 (N_20415,N_17596,N_19331);
nor U20416 (N_20416,N_18970,N_17871);
or U20417 (N_20417,N_17865,N_19721);
or U20418 (N_20418,N_17620,N_19522);
or U20419 (N_20419,N_17405,N_18277);
nand U20420 (N_20420,N_19599,N_17907);
nand U20421 (N_20421,N_15789,N_17232);
or U20422 (N_20422,N_19051,N_16956);
nand U20423 (N_20423,N_16276,N_15988);
or U20424 (N_20424,N_19303,N_16841);
nand U20425 (N_20425,N_17556,N_17584);
or U20426 (N_20426,N_15111,N_19114);
nor U20427 (N_20427,N_17469,N_19734);
and U20428 (N_20428,N_18683,N_19914);
and U20429 (N_20429,N_18625,N_17607);
nor U20430 (N_20430,N_15164,N_15727);
xor U20431 (N_20431,N_16290,N_15185);
nor U20432 (N_20432,N_17745,N_16728);
nand U20433 (N_20433,N_17767,N_19896);
or U20434 (N_20434,N_18748,N_17036);
nand U20435 (N_20435,N_17700,N_16589);
or U20436 (N_20436,N_15231,N_18204);
or U20437 (N_20437,N_17210,N_17896);
nand U20438 (N_20438,N_15562,N_18607);
and U20439 (N_20439,N_18590,N_19058);
and U20440 (N_20440,N_19714,N_19678);
and U20441 (N_20441,N_19577,N_15529);
or U20442 (N_20442,N_17138,N_17096);
or U20443 (N_20443,N_16058,N_16607);
or U20444 (N_20444,N_18824,N_19732);
and U20445 (N_20445,N_16936,N_16447);
nor U20446 (N_20446,N_15802,N_18362);
or U20447 (N_20447,N_15384,N_17524);
and U20448 (N_20448,N_18193,N_19286);
and U20449 (N_20449,N_16427,N_16873);
nor U20450 (N_20450,N_19506,N_18385);
nor U20451 (N_20451,N_16714,N_19055);
and U20452 (N_20452,N_16094,N_18507);
nor U20453 (N_20453,N_19054,N_17108);
nand U20454 (N_20454,N_15188,N_19982);
and U20455 (N_20455,N_19990,N_18134);
or U20456 (N_20456,N_19336,N_18675);
nand U20457 (N_20457,N_15968,N_17781);
nand U20458 (N_20458,N_15403,N_19161);
and U20459 (N_20459,N_19638,N_15740);
nor U20460 (N_20460,N_18775,N_18491);
nand U20461 (N_20461,N_15896,N_16176);
and U20462 (N_20462,N_15841,N_19272);
nor U20463 (N_20463,N_15873,N_16676);
or U20464 (N_20464,N_18157,N_15695);
and U20465 (N_20465,N_18570,N_17191);
xor U20466 (N_20466,N_16555,N_17102);
and U20467 (N_20467,N_18875,N_19078);
nor U20468 (N_20468,N_17836,N_18147);
or U20469 (N_20469,N_16734,N_18140);
nand U20470 (N_20470,N_17715,N_17013);
nor U20471 (N_20471,N_19826,N_19801);
nor U20472 (N_20472,N_16317,N_15662);
or U20473 (N_20473,N_16261,N_17383);
and U20474 (N_20474,N_16612,N_18428);
nor U20475 (N_20475,N_16961,N_19812);
and U20476 (N_20476,N_18904,N_19546);
or U20477 (N_20477,N_18958,N_15924);
nand U20478 (N_20478,N_19969,N_16680);
nand U20479 (N_20479,N_16007,N_16367);
nand U20480 (N_20480,N_18592,N_19027);
xor U20481 (N_20481,N_15195,N_19543);
nand U20482 (N_20482,N_15490,N_16542);
and U20483 (N_20483,N_15981,N_18984);
and U20484 (N_20484,N_19276,N_18176);
and U20485 (N_20485,N_19375,N_15183);
xor U20486 (N_20486,N_18891,N_16067);
nor U20487 (N_20487,N_16799,N_19269);
and U20488 (N_20488,N_17812,N_17928);
or U20489 (N_20489,N_19915,N_18800);
nor U20490 (N_20490,N_18439,N_18583);
and U20491 (N_20491,N_17670,N_19366);
and U20492 (N_20492,N_18899,N_17646);
nand U20493 (N_20493,N_15973,N_18495);
nand U20494 (N_20494,N_16014,N_15110);
and U20495 (N_20495,N_17937,N_17615);
nand U20496 (N_20496,N_15721,N_17608);
nand U20497 (N_20497,N_19545,N_15365);
or U20498 (N_20498,N_19838,N_15448);
and U20499 (N_20499,N_18274,N_18681);
or U20500 (N_20500,N_16827,N_18374);
or U20501 (N_20501,N_19750,N_18234);
nor U20502 (N_20502,N_17116,N_16095);
nor U20503 (N_20503,N_17415,N_18663);
or U20504 (N_20504,N_18172,N_19311);
and U20505 (N_20505,N_16667,N_19551);
or U20506 (N_20506,N_19224,N_16459);
and U20507 (N_20507,N_15096,N_17125);
or U20508 (N_20508,N_17192,N_19977);
nand U20509 (N_20509,N_18754,N_18770);
or U20510 (N_20510,N_17049,N_19064);
nand U20511 (N_20511,N_17625,N_19574);
nor U20512 (N_20512,N_18111,N_18780);
nand U20513 (N_20513,N_15165,N_16494);
and U20514 (N_20514,N_17438,N_18043);
or U20515 (N_20515,N_18833,N_15769);
nand U20516 (N_20516,N_16989,N_17961);
nand U20517 (N_20517,N_19534,N_18901);
nand U20518 (N_20518,N_19945,N_18230);
and U20519 (N_20519,N_15808,N_16920);
or U20520 (N_20520,N_16532,N_15702);
nor U20521 (N_20521,N_17392,N_17877);
nor U20522 (N_20522,N_16083,N_15053);
and U20523 (N_20523,N_16964,N_16779);
nand U20524 (N_20524,N_16783,N_18287);
and U20525 (N_20525,N_16455,N_17917);
or U20526 (N_20526,N_19512,N_18608);
nand U20527 (N_20527,N_17787,N_15665);
and U20528 (N_20528,N_16208,N_15547);
nand U20529 (N_20529,N_19170,N_15844);
or U20530 (N_20530,N_18076,N_15171);
or U20531 (N_20531,N_18624,N_18528);
and U20532 (N_20532,N_15956,N_19243);
or U20533 (N_20533,N_17926,N_16294);
or U20534 (N_20534,N_18883,N_15258);
nor U20535 (N_20535,N_17416,N_15771);
or U20536 (N_20536,N_19377,N_15140);
xnor U20537 (N_20537,N_15512,N_19727);
or U20538 (N_20538,N_17288,N_19110);
or U20539 (N_20539,N_15201,N_15880);
nand U20540 (N_20540,N_19967,N_16743);
nand U20541 (N_20541,N_18095,N_17213);
or U20542 (N_20542,N_16670,N_19241);
nand U20543 (N_20543,N_17137,N_17250);
nor U20544 (N_20544,N_19339,N_15169);
nor U20545 (N_20545,N_17411,N_18059);
and U20546 (N_20546,N_18591,N_16465);
or U20547 (N_20547,N_18829,N_15581);
or U20548 (N_20548,N_17474,N_19484);
and U20549 (N_20549,N_18882,N_15813);
or U20550 (N_20550,N_16376,N_18093);
nand U20551 (N_20551,N_16896,N_16444);
or U20552 (N_20552,N_18406,N_18075);
nor U20553 (N_20553,N_19668,N_18150);
and U20554 (N_20554,N_16726,N_18687);
or U20555 (N_20555,N_17076,N_19539);
or U20556 (N_20556,N_16836,N_18611);
or U20557 (N_20557,N_17273,N_16320);
or U20558 (N_20558,N_18206,N_17347);
nand U20559 (N_20559,N_17178,N_18582);
or U20560 (N_20560,N_16692,N_18077);
and U20561 (N_20561,N_18933,N_17808);
nor U20562 (N_20562,N_19227,N_19120);
nand U20563 (N_20563,N_18709,N_18914);
or U20564 (N_20564,N_16500,N_18639);
and U20565 (N_20565,N_19414,N_17658);
or U20566 (N_20566,N_16987,N_16243);
nand U20567 (N_20567,N_15784,N_18165);
and U20568 (N_20568,N_19560,N_16358);
nor U20569 (N_20569,N_19016,N_17738);
or U20570 (N_20570,N_16021,N_16313);
and U20571 (N_20571,N_19119,N_18731);
or U20572 (N_20572,N_19712,N_16650);
nand U20573 (N_20573,N_15469,N_18651);
nor U20574 (N_20574,N_19876,N_19073);
nand U20575 (N_20575,N_16081,N_18235);
nor U20576 (N_20576,N_17567,N_17484);
or U20577 (N_20577,N_15521,N_16795);
or U20578 (N_20578,N_19306,N_19160);
nand U20579 (N_20579,N_17820,N_17153);
and U20580 (N_20580,N_18372,N_15810);
and U20581 (N_20581,N_19309,N_19067);
nand U20582 (N_20582,N_17814,N_17089);
xnor U20583 (N_20583,N_17675,N_16925);
or U20584 (N_20584,N_18587,N_15292);
nor U20585 (N_20585,N_17936,N_18452);
nor U20586 (N_20586,N_19740,N_16020);
nor U20587 (N_20587,N_16599,N_16942);
nand U20588 (N_20588,N_16908,N_19538);
nor U20589 (N_20589,N_15316,N_17311);
nand U20590 (N_20590,N_18539,N_17623);
and U20591 (N_20591,N_15037,N_19895);
nand U20592 (N_20592,N_17188,N_17291);
and U20593 (N_20593,N_19840,N_17695);
nand U20594 (N_20594,N_17113,N_18746);
xnor U20595 (N_20595,N_18866,N_15271);
nand U20596 (N_20596,N_15295,N_15557);
nand U20597 (N_20597,N_16996,N_17157);
or U20598 (N_20598,N_18765,N_15214);
nand U20599 (N_20599,N_17228,N_19935);
or U20600 (N_20600,N_19488,N_15203);
nor U20601 (N_20601,N_16406,N_16488);
or U20602 (N_20602,N_17312,N_19847);
or U20603 (N_20603,N_16468,N_19504);
or U20604 (N_20604,N_17421,N_19614);
nor U20605 (N_20605,N_15310,N_19186);
or U20606 (N_20606,N_19104,N_16539);
or U20607 (N_20607,N_18278,N_16168);
and U20608 (N_20608,N_17149,N_15373);
nor U20609 (N_20609,N_16438,N_19850);
or U20610 (N_20610,N_15943,N_15931);
nand U20611 (N_20611,N_18580,N_19325);
nand U20612 (N_20612,N_17750,N_15108);
nor U20613 (N_20613,N_16157,N_19228);
nor U20614 (N_20614,N_18542,N_18174);
and U20615 (N_20615,N_15002,N_17721);
nand U20616 (N_20616,N_19281,N_19954);
xnor U20617 (N_20617,N_19700,N_18082);
or U20618 (N_20618,N_16821,N_19215);
and U20619 (N_20619,N_17979,N_15381);
and U20620 (N_20620,N_19039,N_16266);
or U20621 (N_20621,N_16190,N_17120);
and U20622 (N_20622,N_16417,N_17744);
nand U20623 (N_20623,N_18072,N_19956);
nand U20624 (N_20624,N_17064,N_16485);
nor U20625 (N_20625,N_18342,N_15429);
xor U20626 (N_20626,N_18447,N_19236);
and U20627 (N_20627,N_17284,N_15858);
and U20628 (N_20628,N_18723,N_16334);
nand U20629 (N_20629,N_18531,N_16180);
and U20630 (N_20630,N_18137,N_19258);
nor U20631 (N_20631,N_15212,N_16865);
nor U20632 (N_20632,N_17557,N_16325);
nand U20633 (N_20633,N_18422,N_17795);
nand U20634 (N_20634,N_19572,N_16684);
nand U20635 (N_20635,N_19856,N_16971);
nand U20636 (N_20636,N_18657,N_17921);
nand U20637 (N_20637,N_18484,N_18148);
nor U20638 (N_20638,N_17122,N_16365);
or U20639 (N_20639,N_19744,N_17791);
and U20640 (N_20640,N_15713,N_15615);
xor U20641 (N_20641,N_19202,N_18783);
xor U20642 (N_20642,N_15398,N_15723);
nand U20643 (N_20643,N_15977,N_19441);
and U20644 (N_20644,N_18752,N_17768);
nand U20645 (N_20645,N_19957,N_17286);
and U20646 (N_20646,N_19044,N_16593);
nand U20647 (N_20647,N_15099,N_18795);
nor U20648 (N_20648,N_18696,N_17580);
nor U20649 (N_20649,N_16127,N_18701);
or U20650 (N_20650,N_18633,N_18616);
or U20651 (N_20651,N_15567,N_15150);
nor U20652 (N_20652,N_17380,N_17699);
or U20653 (N_20653,N_16217,N_16469);
or U20654 (N_20654,N_15380,N_18597);
nor U20655 (N_20655,N_17924,N_15208);
nor U20656 (N_20656,N_17943,N_15895);
nand U20657 (N_20657,N_19767,N_19450);
or U20658 (N_20658,N_19611,N_17410);
or U20659 (N_20659,N_16571,N_18811);
and U20660 (N_20660,N_17777,N_18469);
nor U20661 (N_20661,N_16159,N_16810);
nand U20662 (N_20662,N_19770,N_16944);
and U20663 (N_20663,N_17230,N_15462);
and U20664 (N_20664,N_16939,N_18516);
nand U20665 (N_20665,N_19109,N_15399);
or U20666 (N_20666,N_15430,N_18031);
or U20667 (N_20667,N_15401,N_17573);
nor U20668 (N_20668,N_15225,N_15523);
or U20669 (N_20669,N_17259,N_16847);
nand U20670 (N_20670,N_16181,N_15963);
xor U20671 (N_20671,N_18154,N_15112);
or U20672 (N_20672,N_19434,N_17444);
nor U20673 (N_20673,N_15339,N_15531);
or U20674 (N_20674,N_16771,N_17289);
nand U20675 (N_20675,N_17139,N_16251);
nand U20676 (N_20676,N_19918,N_17988);
and U20677 (N_20677,N_16093,N_18327);
nand U20678 (N_20678,N_18339,N_16116);
nand U20679 (N_20679,N_19473,N_17281);
nor U20680 (N_20680,N_19165,N_17884);
nand U20681 (N_20681,N_19729,N_17046);
nand U20682 (N_20682,N_16619,N_17354);
or U20683 (N_20683,N_17319,N_17374);
nand U20684 (N_20684,N_19057,N_18840);
or U20685 (N_20685,N_16112,N_16046);
nor U20686 (N_20686,N_16745,N_17736);
or U20687 (N_20687,N_17632,N_16371);
nor U20688 (N_20688,N_17406,N_18407);
and U20689 (N_20689,N_18027,N_15418);
nor U20690 (N_20690,N_17664,N_15593);
xor U20691 (N_20691,N_17245,N_16711);
nand U20692 (N_20692,N_19986,N_15862);
or U20693 (N_20693,N_19443,N_19103);
and U20694 (N_20694,N_15826,N_18619);
or U20695 (N_20695,N_15929,N_18022);
nor U20696 (N_20696,N_17132,N_17647);
or U20697 (N_20697,N_19013,N_19670);
nand U20698 (N_20698,N_18670,N_17735);
or U20699 (N_20699,N_16006,N_18107);
and U20700 (N_20700,N_19179,N_17499);
and U20701 (N_20701,N_18512,N_15693);
xor U20702 (N_20702,N_18854,N_15090);
nor U20703 (N_20703,N_19398,N_18255);
or U20704 (N_20704,N_17168,N_19703);
nand U20705 (N_20705,N_15239,N_15829);
or U20706 (N_20706,N_15757,N_19890);
nand U20707 (N_20707,N_17965,N_19417);
nor U20708 (N_20708,N_15883,N_15269);
and U20709 (N_20709,N_15556,N_17028);
or U20710 (N_20710,N_16138,N_19553);
or U20711 (N_20711,N_16941,N_15621);
nand U20712 (N_20712,N_19650,N_16349);
nand U20713 (N_20713,N_19661,N_15005);
or U20714 (N_20714,N_15013,N_15358);
or U20715 (N_20715,N_17780,N_19265);
nor U20716 (N_20716,N_17967,N_18463);
nor U20717 (N_20717,N_17868,N_18112);
nand U20718 (N_20718,N_17838,N_19454);
or U20719 (N_20719,N_15387,N_19242);
or U20720 (N_20720,N_17216,N_19762);
nand U20721 (N_20721,N_16277,N_17753);
and U20722 (N_20722,N_16418,N_18892);
nor U20723 (N_20723,N_15526,N_16854);
and U20724 (N_20724,N_17786,N_15679);
nor U20725 (N_20725,N_15483,N_19549);
nor U20726 (N_20726,N_16501,N_16875);
nand U20727 (N_20727,N_15657,N_19881);
nor U20728 (N_20728,N_15624,N_18536);
and U20729 (N_20729,N_19458,N_18376);
nand U20730 (N_20730,N_18471,N_16145);
nand U20731 (N_20731,N_16540,N_16993);
nand U20732 (N_20732,N_17548,N_15815);
nand U20733 (N_20733,N_16192,N_17793);
nand U20734 (N_20734,N_18190,N_16530);
and U20735 (N_20735,N_19694,N_19663);
nor U20736 (N_20736,N_16023,N_17235);
nor U20737 (N_20737,N_17860,N_18604);
and U20738 (N_20738,N_17094,N_16134);
or U20739 (N_20739,N_18123,N_19296);
and U20740 (N_20740,N_17370,N_19533);
or U20741 (N_20741,N_15734,N_17151);
or U20742 (N_20742,N_17001,N_16629);
nor U20743 (N_20743,N_19250,N_17485);
and U20744 (N_20744,N_17686,N_17689);
nor U20745 (N_20745,N_15715,N_16702);
and U20746 (N_20746,N_18142,N_15519);
nand U20747 (N_20747,N_15088,N_17816);
or U20748 (N_20748,N_16765,N_16704);
nand U20749 (N_20749,N_16723,N_19697);
nor U20750 (N_20750,N_16758,N_17082);
xnor U20751 (N_20751,N_19247,N_18009);
and U20752 (N_20752,N_17369,N_16169);
nand U20753 (N_20753,N_16673,N_16802);
nor U20754 (N_20754,N_18168,N_18526);
nor U20755 (N_20755,N_19072,N_16397);
and U20756 (N_20756,N_17809,N_17575);
or U20757 (N_20757,N_19755,N_16082);
or U20758 (N_20758,N_17525,N_15586);
nor U20759 (N_20759,N_16031,N_16826);
and U20760 (N_20760,N_19455,N_15912);
nor U20761 (N_20761,N_18821,N_19823);
nor U20762 (N_20762,N_17985,N_17368);
or U20763 (N_20763,N_17732,N_19446);
nor U20764 (N_20764,N_19642,N_16356);
and U20765 (N_20765,N_15137,N_17941);
or U20766 (N_20766,N_18927,N_16229);
or U20767 (N_20767,N_19068,N_18465);
nand U20768 (N_20768,N_17561,N_17858);
nor U20769 (N_20769,N_15209,N_18739);
and U20770 (N_20770,N_17104,N_15812);
xnor U20771 (N_20771,N_18987,N_16477);
or U20772 (N_20772,N_15821,N_15775);
nor U20773 (N_20773,N_18532,N_15542);
xor U20774 (N_20774,N_18396,N_17110);
nor U20775 (N_20775,N_19862,N_15261);
and U20776 (N_20776,N_15803,N_18552);
and U20777 (N_20777,N_18161,N_17373);
or U20778 (N_20778,N_15032,N_17017);
and U20779 (N_20779,N_18888,N_17913);
and U20780 (N_20780,N_19308,N_18208);
or U20781 (N_20781,N_17660,N_16197);
and U20782 (N_20782,N_17304,N_15160);
and U20783 (N_20783,N_15640,N_19433);
nor U20784 (N_20784,N_17103,N_17414);
nor U20785 (N_20785,N_16700,N_16965);
and U20786 (N_20786,N_19569,N_19395);
nand U20787 (N_20787,N_16158,N_15585);
and U20788 (N_20788,N_19305,N_17212);
nor U20789 (N_20789,N_17086,N_19211);
nand U20790 (N_20790,N_18533,N_18945);
or U20791 (N_20791,N_17806,N_15944);
or U20792 (N_20792,N_15272,N_15960);
and U20793 (N_20793,N_16184,N_17805);
nand U20794 (N_20794,N_17790,N_15654);
and U20795 (N_20795,N_15717,N_18016);
nor U20796 (N_20796,N_15971,N_16080);
or U20797 (N_20797,N_15317,N_19828);
xnor U20798 (N_20798,N_18451,N_16535);
and U20799 (N_20799,N_18061,N_17209);
nor U20800 (N_20800,N_16884,N_15166);
nor U20801 (N_20801,N_16092,N_17953);
or U20802 (N_20802,N_19063,N_17667);
or U20803 (N_20803,N_19839,N_15892);
nor U20804 (N_20804,N_16932,N_15211);
or U20805 (N_20805,N_18306,N_17456);
nor U20806 (N_20806,N_17447,N_16811);
nand U20807 (N_20807,N_19963,N_18614);
nand U20808 (N_20808,N_15372,N_16844);
nand U20809 (N_20809,N_15619,N_17497);
nor U20810 (N_20810,N_17450,N_17842);
or U20811 (N_20811,N_18248,N_16090);
nand U20812 (N_20812,N_15564,N_19806);
nand U20813 (N_20813,N_18220,N_18070);
or U20814 (N_20814,N_16660,N_16703);
nor U20815 (N_20815,N_18403,N_15911);
nor U20816 (N_20816,N_17823,N_18273);
nor U20817 (N_20817,N_16644,N_17815);
nand U20818 (N_20818,N_16905,N_15502);
nand U20819 (N_20819,N_15307,N_18718);
nand U20820 (N_20820,N_16888,N_18623);
or U20821 (N_20821,N_15299,N_16958);
or U20822 (N_20822,N_17716,N_16833);
or U20823 (N_20823,N_16577,N_17155);
nand U20824 (N_20824,N_18279,N_15428);
and U20825 (N_20825,N_16921,N_15354);
nor U20826 (N_20826,N_16248,N_16887);
nand U20827 (N_20827,N_17481,N_15106);
nand U20828 (N_20828,N_18014,N_16131);
or U20829 (N_20829,N_16729,N_16059);
and U20830 (N_20830,N_15036,N_18308);
and U20831 (N_20831,N_18139,N_16352);
nand U20832 (N_20832,N_15532,N_17218);
xnor U20833 (N_20833,N_15480,N_16849);
nand U20834 (N_20834,N_18721,N_15202);
and U20835 (N_20835,N_18543,N_16788);
nand U20836 (N_20836,N_18816,N_18085);
nor U20837 (N_20837,N_19219,N_15607);
nor U20838 (N_20838,N_17413,N_18781);
nand U20839 (N_20839,N_18316,N_17234);
and U20840 (N_20840,N_15536,N_15798);
or U20841 (N_20841,N_19127,N_15995);
nor U20842 (N_20842,N_15504,N_19102);
and U20843 (N_20843,N_19509,N_18885);
and U20844 (N_20844,N_18950,N_16162);
nor U20845 (N_20845,N_16189,N_17900);
or U20846 (N_20846,N_15842,N_16645);
or U20847 (N_20847,N_18196,N_17693);
or U20848 (N_20848,N_15814,N_15745);
or U20849 (N_20849,N_19747,N_18155);
nor U20850 (N_20850,N_17078,N_15363);
or U20851 (N_20851,N_17068,N_15869);
xnor U20852 (N_20852,N_15758,N_19391);
nor U20853 (N_20853,N_16891,N_19659);
nor U20854 (N_20854,N_17766,N_16076);
nand U20855 (N_20855,N_17516,N_17934);
nand U20856 (N_20856,N_16360,N_15041);
or U20857 (N_20857,N_15806,N_17800);
nor U20858 (N_20858,N_18038,N_19394);
or U20859 (N_20859,N_18629,N_19400);
and U20860 (N_20860,N_16102,N_16433);
or U20861 (N_20861,N_19069,N_17303);
or U20862 (N_20862,N_17602,N_19541);
and U20863 (N_20863,N_18572,N_18183);
nor U20864 (N_20864,N_16909,N_16620);
nand U20865 (N_20865,N_16318,N_16204);
and U20866 (N_20866,N_17043,N_16770);
and U20867 (N_20867,N_16281,N_19122);
and U20868 (N_20868,N_16391,N_17378);
xnor U20869 (N_20869,N_19946,N_15252);
nand U20870 (N_20870,N_15737,N_16718);
nand U20871 (N_20871,N_18690,N_19251);
nand U20872 (N_20872,N_16271,N_19837);
nand U20873 (N_20873,N_18805,N_17653);
and U20874 (N_20874,N_19836,N_17074);
and U20875 (N_20875,N_15847,N_19997);
or U20876 (N_20876,N_18584,N_19239);
or U20877 (N_20877,N_19086,N_16840);
nor U20878 (N_20878,N_16220,N_15196);
nor U20879 (N_20879,N_17257,N_17225);
and U20880 (N_20880,N_16721,N_18418);
nor U20881 (N_20881,N_16853,N_16689);
or U20882 (N_20882,N_17047,N_18240);
nand U20883 (N_20883,N_16011,N_15865);
and U20884 (N_20884,N_17761,N_19116);
nor U20885 (N_20885,N_16299,N_17067);
nand U20886 (N_20886,N_15690,N_15226);
or U20887 (N_20887,N_15935,N_16215);
and U20888 (N_20888,N_18423,N_16443);
nand U20889 (N_20889,N_17241,N_18969);
or U20890 (N_20890,N_19516,N_15980);
nor U20891 (N_20891,N_17226,N_16621);
nand U20892 (N_20892,N_19870,N_16019);
nor U20893 (N_20893,N_19807,N_18586);
or U20894 (N_20894,N_16435,N_17956);
nor U20895 (N_20895,N_17605,N_17026);
and U20896 (N_20896,N_18991,N_18601);
and U20897 (N_20897,N_18566,N_18264);
or U20898 (N_20898,N_19252,N_15259);
nand U20899 (N_20899,N_16681,N_17511);
nor U20900 (N_20900,N_15033,N_18007);
xor U20901 (N_20901,N_16753,N_18352);
or U20902 (N_20902,N_17251,N_19748);
and U20903 (N_20903,N_18119,N_19282);
nor U20904 (N_20904,N_19424,N_15603);
nor U20905 (N_20905,N_15347,N_16383);
nor U20906 (N_20906,N_18237,N_16919);
nand U20907 (N_20907,N_18814,N_15902);
nor U20908 (N_20908,N_17672,N_19278);
nor U20909 (N_20909,N_16508,N_16182);
or U20910 (N_20910,N_15597,N_16089);
and U20911 (N_20911,N_18354,N_15411);
and U20912 (N_20912,N_15331,N_19910);
nor U20913 (N_20913,N_16843,N_19480);
nand U20914 (N_20914,N_18886,N_18494);
or U20915 (N_20915,N_17986,N_19230);
and U20916 (N_20916,N_17696,N_16586);
or U20917 (N_20917,N_19233,N_16894);
nor U20918 (N_20918,N_18357,N_18820);
nor U20919 (N_20919,N_16792,N_17431);
or U20920 (N_20920,N_16715,N_19413);
nand U20921 (N_20921,N_19537,N_16462);
or U20922 (N_20922,N_16549,N_17338);
nor U20923 (N_20923,N_17270,N_15357);
nand U20924 (N_20924,N_19644,N_15820);
nor U20925 (N_20925,N_17340,N_15070);
or U20926 (N_20926,N_17287,N_18067);
or U20927 (N_20927,N_19136,N_18384);
nor U20928 (N_20928,N_19312,N_16708);
and U20929 (N_20929,N_17163,N_18858);
and U20930 (N_20930,N_19595,N_18225);
nor U20931 (N_20931,N_15967,N_17980);
nor U20932 (N_20932,N_16348,N_17798);
or U20933 (N_20933,N_15267,N_19908);
nand U20934 (N_20934,N_16335,N_19585);
or U20935 (N_20935,N_18563,N_15494);
nor U20936 (N_20936,N_17222,N_15735);
or U20937 (N_20937,N_16098,N_19690);
and U20938 (N_20938,N_16489,N_15010);
nand U20939 (N_20939,N_17701,N_18911);
nor U20940 (N_20940,N_16174,N_17247);
nor U20941 (N_20941,N_15761,N_15752);
or U20942 (N_20942,N_18051,N_15604);
or U20943 (N_20943,N_16513,N_19192);
nor U20944 (N_20944,N_15687,N_19285);
or U20945 (N_20945,N_15800,N_19978);
nand U20946 (N_20946,N_16968,N_19210);
nand U20947 (N_20947,N_17821,N_16456);
and U20948 (N_20948,N_19612,N_17942);
and U20949 (N_20949,N_18573,N_18909);
nand U20950 (N_20950,N_17782,N_17734);
nor U20951 (N_20951,N_15613,N_19961);
and U20952 (N_20952,N_16171,N_15006);
nand U20953 (N_20953,N_16259,N_18955);
nor U20954 (N_20954,N_17446,N_18907);
and U20955 (N_20955,N_18518,N_16268);
and U20956 (N_20956,N_17057,N_17910);
or U20957 (N_20957,N_19851,N_19601);
or U20958 (N_20958,N_15525,N_18768);
and U20959 (N_20959,N_15298,N_18015);
or U20960 (N_20960,N_19324,N_19001);
nor U20961 (N_20961,N_15774,N_15994);
nor U20962 (N_20962,N_18429,N_18916);
nor U20963 (N_20963,N_16694,N_19679);
or U20964 (N_20964,N_17285,N_15948);
or U20965 (N_20965,N_19362,N_19159);
nor U20966 (N_20966,N_15296,N_18510);
and U20967 (N_20967,N_16274,N_18455);
nand U20968 (N_20968,N_19675,N_19615);
or U20969 (N_20969,N_18822,N_17629);
nor U20970 (N_20970,N_19043,N_17830);
nor U20971 (N_20971,N_16787,N_18728);
nor U20972 (N_20972,N_18921,N_16716);
nand U20973 (N_20973,N_17966,N_18121);
or U20974 (N_20974,N_16167,N_19370);
or U20975 (N_20975,N_19329,N_18241);
and U20976 (N_20976,N_18954,N_16806);
or U20977 (N_20977,N_16133,N_19641);
nor U20978 (N_20978,N_18200,N_18138);
or U20979 (N_20979,N_15894,N_19605);
or U20980 (N_20980,N_18541,N_18939);
nand U20981 (N_20981,N_18453,N_15402);
nand U20982 (N_20982,N_18565,N_16150);
or U20983 (N_20983,N_17293,N_19923);
or U20984 (N_20984,N_19030,N_15199);
nor U20985 (N_20985,N_18135,N_17507);
and U20986 (N_20986,N_18351,N_16223);
nand U20987 (N_20987,N_18114,N_19483);
or U20988 (N_20988,N_15923,N_17829);
nor U20989 (N_20989,N_15066,N_16804);
and U20990 (N_20990,N_16421,N_15496);
nor U20991 (N_20991,N_15778,N_16669);
and U20992 (N_20992,N_18652,N_19390);
or U20993 (N_20993,N_15952,N_17652);
or U20994 (N_20994,N_15965,N_16201);
nor U20995 (N_20995,N_17501,N_16305);
and U20996 (N_20996,N_18223,N_19404);
and U20997 (N_20997,N_19814,N_16085);
nand U20998 (N_20998,N_17968,N_17562);
and U20999 (N_20999,N_17619,N_18635);
and U21000 (N_21000,N_17972,N_19785);
nor U21001 (N_21001,N_17016,N_15658);
nand U21002 (N_21002,N_18250,N_19310);
nand U21003 (N_21003,N_16339,N_18642);
and U21004 (N_21004,N_18050,N_18913);
nor U21005 (N_21005,N_18847,N_19671);
and U21006 (N_21006,N_19350,N_18880);
or U21007 (N_21007,N_17454,N_19259);
and U21008 (N_21008,N_19368,N_18381);
nand U21009 (N_21009,N_18517,N_18771);
nor U21010 (N_21010,N_17540,N_16866);
nand U21011 (N_21011,N_16218,N_17020);
nor U21012 (N_21012,N_16253,N_17757);
or U21013 (N_21013,N_16463,N_19323);
nand U21014 (N_21014,N_16042,N_15260);
nor U21015 (N_21015,N_16614,N_15887);
and U21016 (N_21016,N_18868,N_17702);
or U21017 (N_21017,N_17948,N_17042);
nor U21018 (N_21018,N_19080,N_18941);
or U21019 (N_21019,N_18057,N_15375);
nand U21020 (N_21020,N_15035,N_16173);
and U21021 (N_21021,N_15809,N_16630);
nor U21022 (N_21022,N_17279,N_19547);
or U21023 (N_21023,N_15823,N_16175);
or U21024 (N_21024,N_15138,N_18971);
or U21025 (N_21025,N_17221,N_17384);
nand U21026 (N_21026,N_16946,N_18104);
xnor U21027 (N_21027,N_16760,N_19098);
or U21028 (N_21028,N_18209,N_16962);
nor U21029 (N_21029,N_16835,N_15022);
nor U21030 (N_21030,N_19760,N_18323);
nand U21031 (N_21031,N_19264,N_17893);
nor U21032 (N_21032,N_19903,N_17984);
and U21033 (N_21033,N_17208,N_17707);
and U21034 (N_21034,N_16938,N_18257);
or U21035 (N_21035,N_19944,N_19792);
nand U21036 (N_21036,N_15009,N_18515);
and U21037 (N_21037,N_18040,N_17727);
nor U21038 (N_21038,N_19754,N_15057);
or U21039 (N_21039,N_17451,N_15162);
nand U21040 (N_21040,N_15236,N_19706);
nor U21041 (N_21041,N_18874,N_18391);
xor U21042 (N_21042,N_19777,N_16643);
nand U21043 (N_21043,N_15688,N_17692);
nand U21044 (N_21044,N_15173,N_15233);
or U21045 (N_21045,N_19508,N_15867);
and U21046 (N_21046,N_15499,N_17045);
nand U21047 (N_21047,N_15016,N_17688);
nand U21048 (N_21048,N_18192,N_16453);
and U21049 (N_21049,N_19156,N_16690);
nand U21050 (N_21050,N_17359,N_18304);
nor U21051 (N_21051,N_19031,N_18254);
or U21052 (N_21052,N_18679,N_16774);
or U21053 (N_21053,N_18706,N_18153);
nor U21054 (N_21054,N_19153,N_19568);
and U21055 (N_21055,N_18052,N_15793);
or U21056 (N_21056,N_17428,N_19713);
nand U21057 (N_21057,N_16420,N_19773);
nor U21058 (N_21058,N_15059,N_16125);
or U21059 (N_21059,N_17248,N_18636);
nor U21060 (N_21060,N_19804,N_15223);
nor U21061 (N_21061,N_15038,N_15045);
nand U21062 (N_21062,N_16164,N_18965);
or U21063 (N_21063,N_19117,N_17182);
or U21064 (N_21064,N_17657,N_18897);
or U21065 (N_21065,N_16949,N_18537);
nand U21066 (N_21066,N_16724,N_15612);
nor U21067 (N_21067,N_17314,N_17833);
and U21068 (N_21068,N_15091,N_16449);
nand U21069 (N_21069,N_15135,N_19045);
or U21070 (N_21070,N_17530,N_17295);
and U21071 (N_21071,N_17834,N_18588);
or U21072 (N_21072,N_15724,N_19040);
nor U21073 (N_21073,N_19672,N_17432);
or U21074 (N_21074,N_15939,N_16063);
nor U21075 (N_21075,N_15878,N_19318);
nand U21076 (N_21076,N_15309,N_16737);
and U21077 (N_21077,N_16024,N_19158);
nand U21078 (N_21078,N_15434,N_15262);
and U21079 (N_21079,N_17574,N_19502);
nor U21080 (N_21080,N_15975,N_15205);
or U21081 (N_21081,N_18480,N_15620);
nand U21082 (N_21082,N_16808,N_16725);
nand U21083 (N_21083,N_19853,N_19384);
nor U21084 (N_21084,N_19079,N_17088);
or U21085 (N_21085,N_19154,N_16951);
nor U21086 (N_21086,N_16032,N_18443);
xnor U21087 (N_21087,N_17971,N_15424);
and U21088 (N_21088,N_17100,N_18520);
and U21089 (N_21089,N_16585,N_19827);
and U21090 (N_21090,N_15328,N_16591);
nand U21091 (N_21091,N_19503,N_18482);
nand U21092 (N_21092,N_15760,N_18272);
and U21093 (N_21093,N_17847,N_17872);
nand U21094 (N_21094,N_19682,N_16245);
nand U21095 (N_21095,N_18599,N_19981);
and U21096 (N_21096,N_16518,N_17845);
nor U21097 (N_21097,N_15061,N_18291);
nor U21098 (N_21098,N_15909,N_16001);
and U21099 (N_21099,N_17429,N_18189);
or U21100 (N_21100,N_17857,N_15773);
nor U21101 (N_21101,N_15680,N_15972);
nand U21102 (N_21102,N_16653,N_17198);
nand U21103 (N_21103,N_15431,N_19752);
nand U21104 (N_21104,N_19123,N_19290);
xnor U21105 (N_21105,N_17674,N_15095);
and U21106 (N_21106,N_15610,N_19654);
nand U21107 (N_21107,N_17070,N_15435);
and U21108 (N_21108,N_15290,N_17339);
or U21109 (N_21109,N_15119,N_18175);
nor U21110 (N_21110,N_15733,N_19799);
or U21111 (N_21111,N_15764,N_19774);
or U21112 (N_21112,N_15860,N_16108);
and U21113 (N_21113,N_17598,N_16036);
nand U21114 (N_21114,N_15318,N_19683);
nand U21115 (N_21115,N_18458,N_16776);
nand U21116 (N_21116,N_15343,N_18702);
nand U21117 (N_21117,N_15718,N_16551);
nor U21118 (N_21118,N_16759,N_18427);
nand U21119 (N_21119,N_15749,N_18853);
and U21120 (N_21120,N_19609,N_19619);
and U21121 (N_21121,N_16646,N_16707);
nand U21122 (N_21122,N_15423,N_16486);
nor U21123 (N_21123,N_15533,N_16107);
nor U21124 (N_21124,N_19584,N_19447);
and U21125 (N_21125,N_15840,N_18936);
or U21126 (N_21126,N_16592,N_15184);
and U21127 (N_21127,N_19019,N_15776);
nor U21128 (N_21128,N_19994,N_18233);
nand U21129 (N_21129,N_15371,N_15151);
and U21130 (N_21130,N_19408,N_18186);
nand U21131 (N_21131,N_19053,N_17010);
and U21132 (N_21132,N_17589,N_16519);
nand U21133 (N_21133,N_16608,N_18961);
and U21134 (N_21134,N_15000,N_16512);
nand U21135 (N_21135,N_19111,N_17308);
nor U21136 (N_21136,N_17004,N_17835);
xor U21137 (N_21137,N_16790,N_16966);
and U21138 (N_21138,N_15413,N_19012);
or U21139 (N_21139,N_16374,N_17387);
and U21140 (N_21140,N_15176,N_17310);
and U21141 (N_21141,N_16911,N_16584);
nand U21142 (N_21142,N_16922,N_17635);
nand U21143 (N_21143,N_16580,N_19621);
or U21144 (N_21144,N_17826,N_19759);
nor U21145 (N_21145,N_17442,N_18559);
nor U21146 (N_21146,N_15655,N_18654);
nand U21147 (N_21147,N_15594,N_15447);
and U21148 (N_21148,N_17181,N_19784);
nand U21149 (N_21149,N_17613,N_19976);
nand U21150 (N_21150,N_15664,N_18417);
or U21151 (N_21151,N_19704,N_17018);
and U21152 (N_21152,N_17895,N_18380);
nand U21153 (N_21153,N_16354,N_16017);
or U21154 (N_21154,N_17203,N_17933);
nand U21155 (N_21155,N_19591,N_19163);
nor U21156 (N_21156,N_15833,N_17091);
nand U21157 (N_21157,N_18836,N_17449);
nor U21158 (N_21158,N_16309,N_16997);
or U21159 (N_21159,N_19562,N_18039);
nand U21160 (N_21160,N_17075,N_18977);
nand U21161 (N_21161,N_17764,N_18400);
nand U21162 (N_21162,N_16441,N_17514);
or U21163 (N_21163,N_15906,N_19532);
or U21164 (N_21164,N_19691,N_18364);
nand U21165 (N_21165,N_18753,N_16904);
nor U21166 (N_21166,N_15605,N_18664);
nor U21167 (N_21167,N_18640,N_19200);
nand U21168 (N_21168,N_18645,N_18692);
and U21169 (N_21169,N_19995,N_19778);
xor U21170 (N_21170,N_16830,N_15056);
nand U21171 (N_21171,N_18475,N_18037);
nor U21172 (N_21172,N_16754,N_19907);
and U21173 (N_21173,N_16848,N_19515);
or U21174 (N_21174,N_15315,N_19464);
nand U21175 (N_21175,N_15409,N_16188);
and U21176 (N_21176,N_16381,N_17603);
and U21177 (N_21177,N_17927,N_17973);
nand U21178 (N_21178,N_18008,N_15563);
and U21179 (N_21179,N_15672,N_17643);
or U21180 (N_21180,N_18478,N_17022);
nor U21181 (N_21181,N_15524,N_18412);
nand U21182 (N_21182,N_16387,N_18089);
nand U21183 (N_21183,N_18931,N_18103);
nor U21184 (N_21184,N_19457,N_19926);
and U21185 (N_21185,N_16511,N_18658);
or U21186 (N_21186,N_17894,N_17521);
or U21187 (N_21187,N_16338,N_16688);
or U21188 (N_21188,N_18997,N_17039);
nand U21189 (N_21189,N_17503,N_15830);
nand U21190 (N_21190,N_18715,N_15647);
nor U21191 (N_21191,N_17174,N_18972);
and U21192 (N_21192,N_16088,N_16412);
nor U21193 (N_21193,N_18487,N_18924);
and U21194 (N_21194,N_15982,N_15685);
and U21195 (N_21195,N_17648,N_18295);
or U21196 (N_21196,N_18457,N_17759);
nor U21197 (N_21197,N_16054,N_18558);
and U21198 (N_21198,N_17861,N_16901);
and U21199 (N_21199,N_19403,N_17307);
nor U21200 (N_21200,N_17462,N_19934);
nor U21201 (N_21201,N_16211,N_19026);
nor U21202 (N_21202,N_19326,N_17302);
nand U21203 (N_21203,N_18130,N_15703);
nor U21204 (N_21204,N_15742,N_16341);
nor U21205 (N_21205,N_16221,N_18810);
nor U21206 (N_21206,N_18948,N_17136);
or U21207 (N_21207,N_19772,N_19438);
nand U21208 (N_21208,N_19789,N_15697);
nand U21209 (N_21209,N_16430,N_18239);
and U21210 (N_21210,N_18665,N_16394);
or U21211 (N_21211,N_19217,N_19334);
or U21212 (N_21212,N_16078,N_19048);
nand U21213 (N_21213,N_19291,N_18081);
nand U21214 (N_21214,N_18522,N_17564);
nand U21215 (N_21215,N_18712,N_18890);
and U21216 (N_21216,N_19412,N_15937);
nand U21217 (N_21217,N_19686,N_15622);
and U21218 (N_21218,N_17114,N_19319);
nand U21219 (N_21219,N_18019,N_16675);
or U21220 (N_21220,N_16286,N_18917);
and U21221 (N_21221,N_15368,N_19818);
and U21222 (N_21222,N_19162,N_15280);
nor U21223 (N_21223,N_18684,N_18324);
or U21224 (N_21224,N_15175,N_19731);
and U21225 (N_21225,N_17185,N_15092);
nor U21226 (N_21226,N_18144,N_16527);
nor U21227 (N_21227,N_17752,N_19637);
or U21228 (N_21228,N_15601,N_15804);
and U21229 (N_21229,N_19221,N_16206);
or U21230 (N_21230,N_18850,N_15992);
nor U21231 (N_21231,N_19255,N_18707);
or U21232 (N_21232,N_17704,N_15517);
or U21233 (N_21233,N_17987,N_16390);
or U21234 (N_21234,N_19687,N_17881);
nand U21235 (N_21235,N_18394,N_16798);
xnor U21236 (N_21236,N_16425,N_17490);
nand U21237 (N_21237,N_19942,N_19677);
nand U21238 (N_21238,N_18468,N_17654);
nand U21239 (N_21239,N_15388,N_18503);
and U21240 (N_21240,N_18283,N_19530);
or U21241 (N_21241,N_16284,N_15355);
nor U21242 (N_21242,N_18802,N_15386);
nor U21243 (N_21243,N_15705,N_18889);
or U21244 (N_21244,N_17591,N_16823);
nand U21245 (N_21245,N_15574,N_18647);
nand U21246 (N_21246,N_19175,N_15630);
or U21247 (N_21247,N_18411,N_19579);
nor U21248 (N_21248,N_19523,N_16273);
and U21249 (N_21249,N_19009,N_18408);
and U21250 (N_21250,N_17242,N_15827);
nand U21251 (N_21251,N_17535,N_17142);
nor U21252 (N_21252,N_17038,N_15919);
and U21253 (N_21253,N_17099,N_16809);
nand U21254 (N_21254,N_16570,N_19293);
or U21255 (N_21255,N_15353,N_17638);
and U21256 (N_21256,N_17946,N_15794);
nand U21257 (N_21257,N_18693,N_15817);
nand U21258 (N_21258,N_16216,N_19666);
or U21259 (N_21259,N_18424,N_16154);
nand U21260 (N_21260,N_18349,N_19834);
and U21261 (N_21261,N_15627,N_19492);
and U21262 (N_21262,N_16143,N_18046);
nand U21263 (N_21263,N_16537,N_19470);
and U21264 (N_21264,N_18436,N_16234);
or U21265 (N_21265,N_15270,N_18773);
or U21266 (N_21266,N_19889,N_16442);
and U21267 (N_21267,N_18605,N_15282);
nor U21268 (N_21268,N_17165,N_16568);
and U21269 (N_21269,N_17891,N_15121);
and U21270 (N_21270,N_17642,N_19427);
nor U21271 (N_21271,N_15335,N_19365);
nor U21272 (N_21272,N_15781,N_16146);
nor U21273 (N_21273,N_19449,N_18129);
or U21274 (N_21274,N_18098,N_18275);
and U21275 (N_21275,N_16047,N_17807);
nor U21276 (N_21276,N_15990,N_18529);
nor U21277 (N_21277,N_19187,N_15242);
nand U21278 (N_21278,N_15903,N_17243);
or U21279 (N_21279,N_19000,N_19342);
nor U21280 (N_21280,N_18334,N_16372);
or U21281 (N_21281,N_18667,N_19461);
nand U21282 (N_21282,N_16405,N_17784);
and U21283 (N_21283,N_17506,N_16679);
xor U21284 (N_21284,N_15192,N_16252);
nor U21285 (N_21285,N_16043,N_18908);
nor U21286 (N_21286,N_16732,N_15417);
nand U21287 (N_21287,N_19805,N_19741);
or U21288 (N_21288,N_19453,N_18145);
or U21289 (N_21289,N_17874,N_19145);
or U21290 (N_21290,N_17685,N_19270);
nand U21291 (N_21291,N_15528,N_17087);
nor U21292 (N_21292,N_16050,N_19076);
and U21293 (N_21293,N_17353,N_16177);
nor U21294 (N_21294,N_15344,N_16915);
nor U21295 (N_21295,N_19320,N_16582);
nand U21296 (N_21296,N_16829,N_18159);
and U21297 (N_21297,N_19983,N_18581);
nand U21298 (N_21298,N_16575,N_17662);
nor U21299 (N_21299,N_15692,N_18496);
nand U21300 (N_21300,N_17377,N_15979);
nand U21301 (N_21301,N_18668,N_16214);
or U21302 (N_21302,N_18389,N_17128);
nand U21303 (N_21303,N_18355,N_17301);
nor U21304 (N_21304,N_19347,N_18297);
nand U21305 (N_21305,N_16203,N_17175);
nor U21306 (N_21306,N_15046,N_17831);
nand U21307 (N_21307,N_15487,N_19263);
or U21308 (N_21308,N_19845,N_15479);
nand U21309 (N_21309,N_17878,N_19813);
and U21310 (N_21310,N_19776,N_18102);
nor U21311 (N_21311,N_18096,N_15052);
nand U21312 (N_21312,N_18251,N_17770);
and U21313 (N_21313,N_17095,N_19011);
nand U21314 (N_21314,N_15118,N_18502);
nand U21315 (N_21315,N_15468,N_17822);
and U21316 (N_21316,N_18995,N_15136);
nand U21317 (N_21317,N_15914,N_19719);
nor U21318 (N_21318,N_17193,N_19819);
nor U21319 (N_21319,N_16331,N_17202);
nor U21320 (N_21320,N_15933,N_15544);
or U21321 (N_21321,N_16296,N_18859);
nand U21322 (N_21322,N_19222,N_18567);
nand U21323 (N_21323,N_19146,N_19401);
or U21324 (N_21324,N_18393,N_19195);
or U21325 (N_21325,N_15885,N_16573);
nand U21326 (N_21326,N_18280,N_15663);
and U21327 (N_21327,N_18025,N_17825);
and U21328 (N_21328,N_19066,N_15101);
or U21329 (N_21329,N_19885,N_18986);
nor U21330 (N_21330,N_17362,N_19084);
or U21331 (N_21331,N_17231,N_16730);
and U21332 (N_21332,N_16885,N_19234);
and U21333 (N_21333,N_19498,N_16552);
nand U21334 (N_21334,N_19723,N_19332);
or U21335 (N_21335,N_18325,N_18215);
and U21336 (N_21336,N_17502,N_17052);
or U21337 (N_21337,N_18648,N_17590);
and U21338 (N_21338,N_19194,N_16350);
nor U21339 (N_21339,N_17915,N_18079);
or U21340 (N_21340,N_19094,N_18751);
nand U21341 (N_21341,N_17634,N_16747);
nand U21342 (N_21342,N_17651,N_17436);
nor U21343 (N_21343,N_18363,N_17729);
or U21344 (N_21344,N_17395,N_18792);
nand U21345 (N_21345,N_17604,N_15144);
nand U21346 (N_21346,N_17545,N_16408);
xor U21347 (N_21347,N_16053,N_17852);
nor U21348 (N_21348,N_16543,N_17763);
nor U21349 (N_21349,N_18929,N_17467);
or U21350 (N_21350,N_17024,N_15206);
or U21351 (N_21351,N_17925,N_19439);
and U21352 (N_21352,N_19550,N_19399);
nor U21353 (N_21353,N_16793,N_17817);
nor U21354 (N_21354,N_16115,N_15886);
xnor U21355 (N_21355,N_17543,N_18020);
nor U21356 (N_21356,N_19846,N_17009);
and U21357 (N_21357,N_17708,N_18259);
nor U21358 (N_21358,N_16980,N_18492);
and U21359 (N_21359,N_16517,N_18359);
nor U21360 (N_21360,N_17880,N_18199);
or U21361 (N_21361,N_19904,N_18796);
and U21362 (N_21362,N_15492,N_17526);
nor U21363 (N_21363,N_16357,N_15458);
nand U21364 (N_21364,N_15265,N_16640);
nand U21365 (N_21365,N_17305,N_15268);
nand U21366 (N_21366,N_15816,N_19857);
and U21367 (N_21367,N_15819,N_15157);
nor U21368 (N_21368,N_15694,N_15451);
nor U21369 (N_21369,N_15131,N_15507);
or U21370 (N_21370,N_17135,N_15966);
nor U21371 (N_21371,N_19197,N_18834);
or U21372 (N_21372,N_19736,N_19134);
nand U21373 (N_21373,N_19471,N_16666);
and U21374 (N_21374,N_18041,N_15278);
nand U21375 (N_21375,N_19596,N_17158);
nor U21376 (N_21376,N_18416,N_15720);
or U21377 (N_21377,N_19496,N_19346);
or U21378 (N_21378,N_19101,N_17352);
and U21379 (N_21379,N_15320,N_19410);
nand U21380 (N_21380,N_16879,N_15334);
nor U21381 (N_21381,N_18797,N_15498);
and U21382 (N_21382,N_19505,N_18617);
nand U21383 (N_21383,N_16973,N_16893);
nor U21384 (N_21384,N_17003,N_19373);
nor U21385 (N_21385,N_16232,N_17669);
nor U21386 (N_21386,N_19743,N_19422);
and U21387 (N_21387,N_18508,N_18367);
or U21388 (N_21388,N_15565,N_15346);
nand U21389 (N_21389,N_15497,N_16460);
nor U21390 (N_21390,N_18319,N_17717);
or U21391 (N_21391,N_15908,N_15925);
nor U21392 (N_21392,N_17879,N_15527);
nor U21393 (N_21393,N_15537,N_15832);
nor U21394 (N_21394,N_18178,N_16424);
nand U21395 (N_21395,N_17920,N_15714);
or U21396 (N_21396,N_18293,N_18118);
nor U21397 (N_21397,N_16880,N_18937);
nand U21398 (N_21398,N_18156,N_16429);
nand U21399 (N_21399,N_16139,N_19358);
xor U21400 (N_21400,N_17959,N_18561);
or U21401 (N_21401,N_19948,N_16300);
and U21402 (N_21402,N_17588,N_17532);
nor U21403 (N_21403,N_19475,N_16596);
and U21404 (N_21404,N_15440,N_17053);
nor U21405 (N_21405,N_16475,N_19288);
xor U21406 (N_21406,N_17393,N_16693);
nor U21407 (N_21407,N_15302,N_19720);
or U21408 (N_21408,N_19190,N_18053);
or U21409 (N_21409,N_19379,N_18474);
nor U21410 (N_21410,N_16322,N_15849);
and U21411 (N_21411,N_17568,N_17743);
and U21412 (N_21412,N_19321,N_18564);
or U21413 (N_21413,N_16446,N_15571);
nand U21414 (N_21414,N_16269,N_16870);
nand U21415 (N_21415,N_19226,N_15341);
xnor U21416 (N_21416,N_16389,N_17944);
nand U21417 (N_21417,N_18951,N_19191);
or U21418 (N_21418,N_19796,N_17130);
nand U21419 (N_21419,N_17912,N_16633);
nand U21420 (N_21420,N_15875,N_18074);
nand U21421 (N_21421,N_18160,N_19050);
nor U21422 (N_21422,N_18213,N_16225);
and U21423 (N_21423,N_17866,N_19022);
nand U21424 (N_21424,N_19709,N_19701);
or U21425 (N_21425,N_19658,N_17694);
and U21426 (N_21426,N_17399,N_19432);
and U21427 (N_21427,N_17740,N_16265);
or U21428 (N_21428,N_18873,N_16205);
nand U21429 (N_21429,N_18276,N_19625);
nor U21430 (N_21430,N_19832,N_18271);
and U21431 (N_21431,N_18167,N_19565);
nor U21432 (N_21432,N_15213,N_16330);
nor U21433 (N_21433,N_19133,N_18609);
and U21434 (N_21434,N_17033,N_19971);
nor U21435 (N_21435,N_15759,N_18210);
nor U21436 (N_21436,N_15859,N_19764);
nand U21437 (N_21437,N_15606,N_17124);
and U21438 (N_21438,N_19875,N_18554);
and U21439 (N_21439,N_15686,N_15219);
and U21440 (N_21440,N_18444,N_15190);
and U21441 (N_21441,N_17720,N_15218);
or U21442 (N_21442,N_19298,N_17840);
nor U21443 (N_21443,N_17297,N_19536);
xor U21444 (N_21444,N_15146,N_17783);
nand U21445 (N_21445,N_16558,N_15281);
nand U21446 (N_21446,N_19798,N_15644);
or U21447 (N_21447,N_19301,N_19791);
and U21448 (N_21448,N_17194,N_15716);
or U21449 (N_21449,N_16548,N_16846);
and U21450 (N_21450,N_19528,N_15899);
or U21451 (N_21451,N_15217,N_17282);
xor U21452 (N_21452,N_19629,N_15822);
nand U21453 (N_21453,N_15156,N_18055);
nor U21454 (N_21454,N_17169,N_19113);
and U21455 (N_21455,N_18944,N_17388);
nand U21456 (N_21456,N_19462,N_18962);
and U21457 (N_21457,N_15216,N_15928);
and U21458 (N_21458,N_19289,N_19855);
nor U21459 (N_21459,N_16954,N_18191);
or U21460 (N_21460,N_18000,N_17332);
nand U21461 (N_21461,N_15920,N_16867);
or U21462 (N_21462,N_15378,N_18530);
nand U21463 (N_21463,N_19867,N_16632);
or U21464 (N_21464,N_15855,N_16258);
nand U21465 (N_21465,N_15449,N_18949);
nand U21466 (N_21466,N_18099,N_18934);
nand U21467 (N_21467,N_16008,N_15551);
xnor U21468 (N_21468,N_15730,N_19021);
nand U21469 (N_21469,N_18628,N_15215);
and U21470 (N_21470,N_15124,N_19070);
and U21471 (N_21471,N_15584,N_17908);
nand U21472 (N_21472,N_16604,N_17460);
and U21473 (N_21473,N_18719,N_15555);
nand U21474 (N_21474,N_19105,N_17492);
nor U21475 (N_21475,N_16481,N_16554);
nor U21476 (N_21476,N_17518,N_18301);
nand U21477 (N_21477,N_17906,N_17236);
nor U21478 (N_21478,N_17363,N_16505);
nor U21479 (N_21479,N_16735,N_18894);
and U21480 (N_21480,N_16100,N_16103);
nand U21481 (N_21481,N_18013,N_15568);
or U21482 (N_21482,N_15746,N_17939);
xnor U21483 (N_21483,N_15599,N_16955);
nor U21484 (N_21484,N_15221,N_15069);
or U21485 (N_21485,N_19142,N_17498);
or U21486 (N_21486,N_16553,N_16741);
nor U21487 (N_21487,N_18981,N_19419);
or U21488 (N_21488,N_16978,N_16963);
xnor U21489 (N_21489,N_19886,N_19769);
or U21490 (N_21490,N_16950,N_16567);
nand U21491 (N_21491,N_17592,N_18006);
xor U21492 (N_21492,N_19763,N_19927);
nor U21493 (N_21493,N_17522,N_17523);
or U21494 (N_21494,N_16461,N_16566);
or U21495 (N_21495,N_19559,N_15229);
and U21496 (N_21496,N_19115,N_18310);
nand U21497 (N_21497,N_19531,N_15246);
or U21498 (N_21498,N_17398,N_19639);
nand U21499 (N_21499,N_17478,N_19235);
nand U21500 (N_21500,N_18047,N_18782);
nor U21501 (N_21501,N_19209,N_19869);
or U21502 (N_21502,N_16696,N_17570);
or U21503 (N_21503,N_18353,N_18848);
nand U21504 (N_21504,N_15550,N_17640);
nor U21505 (N_21505,N_17911,N_18818);
nand U21506 (N_21506,N_16470,N_16746);
nor U21507 (N_21507,N_18788,N_16569);
or U21508 (N_21508,N_16306,N_18467);
nand U21509 (N_21509,N_17200,N_15395);
nand U21510 (N_21510,N_16744,N_16039);
nand U21511 (N_21511,N_19497,N_16353);
nand U21512 (N_21512,N_15818,N_19815);
and U21513 (N_21513,N_16812,N_19273);
nor U21514 (N_21514,N_16200,N_18842);
nor U21515 (N_21515,N_18294,N_16407);
and U21516 (N_21516,N_17183,N_17909);
or U21517 (N_21517,N_15838,N_15311);
or U21518 (N_21518,N_18387,N_17356);
xor U21519 (N_21519,N_18184,N_17975);
nor U21520 (N_21520,N_16351,N_19322);
nor U21521 (N_21521,N_18966,N_16524);
nor U21522 (N_21522,N_15366,N_15174);
and U21523 (N_21523,N_19627,N_15026);
and U21524 (N_21524,N_19874,N_18454);
nor U21525 (N_21525,N_19459,N_15628);
and U21526 (N_21526,N_19501,N_15661);
or U21527 (N_21527,N_17488,N_19722);
nor U21528 (N_21528,N_18108,N_16052);
nand U21529 (N_21529,N_15021,N_15614);
nand U21530 (N_21530,N_15274,N_15942);
and U21531 (N_21531,N_15595,N_18555);
and U21532 (N_21532,N_16256,N_19685);
or U21533 (N_21533,N_17612,N_15600);
and U21534 (N_21534,N_15731,N_19647);
or U21535 (N_21535,N_16565,N_19108);
and U21536 (N_21536,N_15093,N_18036);
and U21537 (N_21537,N_15020,N_17846);
and U21538 (N_21538,N_18226,N_19096);
xor U21539 (N_21539,N_19279,N_19947);
or U21540 (N_21540,N_16226,N_15787);
nor U21541 (N_21541,N_19699,N_18550);
nor U21542 (N_21542,N_18767,N_18920);
or U21543 (N_21543,N_15625,N_17848);
or U21544 (N_21544,N_19993,N_18092);
nor U21545 (N_21545,N_15064,N_16999);
or U21546 (N_21546,N_16755,N_18333);
and U21547 (N_21547,N_16316,N_18289);
nor U21548 (N_21548,N_18222,N_15028);
nand U21549 (N_21549,N_18445,N_16613);
nor U21550 (N_21550,N_15250,N_18221);
nor U21551 (N_21551,N_19041,N_19529);
or U21552 (N_21552,N_19888,N_15825);
and U21553 (N_21553,N_15123,N_16210);
nand U21554 (N_21554,N_15998,N_19865);
and U21555 (N_21555,N_18989,N_18677);
nor U21556 (N_21556,N_15279,N_15729);
nor U21557 (N_21557,N_17167,N_17197);
nor U21558 (N_21558,N_15945,N_19626);
nand U21559 (N_21559,N_19527,N_15949);
nand U21560 (N_21560,N_15374,N_16280);
nand U21561 (N_21561,N_19352,N_16035);
nand U21562 (N_21562,N_17811,N_19456);
or U21563 (N_21563,N_15535,N_19337);
and U21564 (N_21564,N_17922,N_19220);
nor U21565 (N_21565,N_16858,N_17520);
or U21566 (N_21566,N_16574,N_16626);
or U21567 (N_21567,N_16907,N_15445);
nor U21568 (N_21568,N_16209,N_15142);
or U21569 (N_21569,N_16025,N_18315);
nand U21570 (N_21570,N_19710,N_16717);
or U21571 (N_21571,N_17671,N_15486);
and U21572 (N_21572,N_18466,N_18772);
and U21573 (N_21573,N_17614,N_18044);
nand U21574 (N_21574,N_17876,N_16368);
or U21575 (N_21575,N_18544,N_16504);
nor U21576 (N_21576,N_16641,N_15362);
or U21577 (N_21577,N_15888,N_17544);
nor U21578 (N_21578,N_16778,N_15050);
nor U21579 (N_21579,N_17056,N_17862);
or U21580 (N_21580,N_18838,N_17509);
and U21581 (N_21581,N_17513,N_18726);
nand U21582 (N_21582,N_18026,N_17144);
nand U21583 (N_21583,N_18211,N_17244);
nor U21584 (N_21584,N_17844,N_18505);
nand U21585 (N_21585,N_15611,N_17261);
and U21586 (N_21586,N_15566,N_18329);
nor U21587 (N_21587,N_19189,N_17560);
or U21588 (N_21588,N_18317,N_18789);
nor U21589 (N_21589,N_16121,N_18678);
nor U21590 (N_21590,N_17616,N_17993);
and U21591 (N_21591,N_18844,N_16403);
and U21592 (N_21592,N_18180,N_16128);
and U21593 (N_21593,N_17935,N_19121);
and U21594 (N_21594,N_16074,N_16506);
nor U21595 (N_21595,N_16972,N_15683);
and U21596 (N_21596,N_16523,N_16947);
or U21597 (N_21597,N_16380,N_16560);
xor U21598 (N_21598,N_18246,N_15405);
and U21599 (N_21599,N_19428,N_15986);
nor U21600 (N_21600,N_16635,N_16818);
or U21601 (N_21601,N_15659,N_15158);
nor U21602 (N_21602,N_15520,N_17037);
and U21603 (N_21603,N_16590,N_19897);
nor U21604 (N_21604,N_19025,N_15522);
nor U21605 (N_21605,N_15616,N_18448);
nand U21606 (N_21606,N_18132,N_19014);
and U21607 (N_21607,N_17668,N_15385);
nor U21608 (N_21608,N_18864,N_18305);
nor U21609 (N_21609,N_15785,N_15127);
nand U21610 (N_21610,N_15921,N_17366);
and U21611 (N_21611,N_19788,N_16110);
and U21612 (N_21612,N_16782,N_15765);
nor U21613 (N_21613,N_19132,N_17903);
nand U21614 (N_21614,N_17379,N_19089);
nand U21615 (N_21615,N_16289,N_19248);
or U21616 (N_21616,N_15044,N_17538);
or U21617 (N_21617,N_15674,N_16178);
or U21618 (N_21618,N_19998,N_15220);
nand U21619 (N_21619,N_18994,N_16148);
nand U21620 (N_21620,N_15836,N_16658);
nand U21621 (N_21621,N_18923,N_17422);
and U21622 (N_21622,N_17143,N_17976);
and U21623 (N_21623,N_18837,N_16752);
and U21624 (N_21624,N_15085,N_19445);
or U21625 (N_21625,N_16084,N_18803);
nand U21626 (N_21626,N_17870,N_18106);
or U21627 (N_21627,N_16536,N_18012);
and U21628 (N_21628,N_18017,N_19824);
and U21629 (N_21629,N_18749,N_19421);
nor U21630 (N_21630,N_19173,N_19905);
nor U21631 (N_21631,N_18084,N_19229);
nor U21632 (N_21632,N_18806,N_16576);
nor U21633 (N_21633,N_19758,N_15369);
nor U21634 (N_21634,N_16852,N_15425);
nor U21635 (N_21635,N_17600,N_16450);
or U21636 (N_21636,N_15407,N_17300);
nor U21637 (N_21637,N_15780,N_16333);
nor U21638 (N_21638,N_16970,N_17583);
nand U21639 (N_21639,N_18252,N_17254);
or U21640 (N_21640,N_19602,N_15450);
nand U21641 (N_21641,N_19029,N_19746);
nor U21642 (N_21642,N_18120,N_15453);
and U21643 (N_21643,N_17998,N_19425);
or U21644 (N_21644,N_16813,N_16863);
or U21645 (N_21645,N_19353,N_15955);
and U21646 (N_21646,N_17885,N_19742);
nor U21647 (N_21647,N_17841,N_17190);
and U21648 (N_21648,N_18370,N_19873);
or U21649 (N_21649,N_17510,N_17869);
and U21650 (N_21650,N_17832,N_18094);
or U21651 (N_21651,N_19841,N_15475);
nor U21652 (N_21652,N_19936,N_15961);
and U21653 (N_21653,N_17931,N_16016);
or U21654 (N_21654,N_16123,N_16324);
nor U21655 (N_21655,N_19930,N_15080);
or U21656 (N_21656,N_15065,N_17875);
or U21657 (N_21657,N_19564,N_15011);
or U21658 (N_21658,N_16065,N_17093);
nand U21659 (N_21659,N_15755,N_15293);
or U21660 (N_21660,N_16895,N_15177);
nand U21661 (N_21661,N_16250,N_15133);
or U21662 (N_21662,N_18143,N_15377);
nand U21663 (N_21663,N_16087,N_15936);
or U21664 (N_21664,N_18763,N_18930);
or U21665 (N_21665,N_15248,N_17537);
nand U21666 (N_21666,N_16699,N_16319);
and U21667 (N_21667,N_15207,N_19126);
or U21668 (N_21668,N_16636,N_16927);
nand U21669 (N_21669,N_17691,N_15861);
and U21670 (N_21670,N_19295,N_15104);
or U21671 (N_21671,N_18181,N_17011);
or U21672 (N_21672,N_17706,N_18569);
nand U21673 (N_21673,N_19302,N_19689);
nand U21674 (N_21674,N_15027,N_17641);
and U21675 (N_21675,N_16710,N_16639);
nand U21676 (N_21676,N_18553,N_16820);
and U21677 (N_21677,N_16890,N_16156);
or U21678 (N_21678,N_15501,N_19698);
and U21679 (N_21679,N_17547,N_16355);
and U21680 (N_21680,N_19212,N_16106);
and U21681 (N_21681,N_18777,N_16364);
xor U21682 (N_21682,N_16479,N_18030);
nor U21683 (N_21683,N_17742,N_18300);
nand U21684 (N_21684,N_16361,N_19877);
nand U21685 (N_21685,N_17897,N_16363);
nand U21686 (N_21686,N_17496,N_17040);
xor U21687 (N_21687,N_19075,N_16238);
nand U21688 (N_21688,N_15852,N_18902);
and U21689 (N_21689,N_17007,N_17769);
and U21690 (N_21690,N_19749,N_16685);
or U21691 (N_21691,N_16149,N_15441);
nor U21692 (N_21692,N_17147,N_15351);
or U21693 (N_21693,N_15739,N_18843);
and U21694 (N_21694,N_16856,N_19141);
nand U21695 (N_21695,N_15756,N_17733);
nand U21696 (N_21696,N_18386,N_18960);
and U21697 (N_21697,N_19975,N_18470);
nand U21698 (N_21698,N_16791,N_19693);
nor U21699 (N_21699,N_19649,N_17109);
nand U21700 (N_21700,N_16207,N_16132);
nor U21701 (N_21701,N_18857,N_16073);
nand U21702 (N_21702,N_15682,N_17550);
nor U21703 (N_21703,N_15303,N_15538);
nor U21704 (N_21704,N_18922,N_16777);
nand U21705 (N_21705,N_15857,N_15848);
nand U21706 (N_21706,N_16712,N_16825);
nand U21707 (N_21707,N_15696,N_15179);
and U21708 (N_21708,N_19442,N_18779);
or U21709 (N_21709,N_19842,N_19166);
nor U21710 (N_21710,N_17546,N_17318);
nor U21711 (N_21711,N_18024,N_16695);
nand U21712 (N_21712,N_15251,N_16395);
or U21713 (N_21713,N_17867,N_15712);
and U21714 (N_21714,N_18703,N_18758);
and U21715 (N_21715,N_17849,N_17256);
nor U21716 (N_21716,N_17853,N_15189);
nor U21717 (N_21717,N_16924,N_16388);
nor U21718 (N_21718,N_18737,N_15639);
and U21719 (N_21719,N_19125,N_17177);
and U21720 (N_21720,N_18345,N_15060);
nand U21721 (N_21721,N_19849,N_18360);
nand U21722 (N_21722,N_17801,N_19087);
nor U21723 (N_21723,N_17684,N_16413);
and U21724 (N_21724,N_15969,N_16327);
nor U21725 (N_21725,N_18872,N_18088);
and U21726 (N_21726,N_17439,N_18244);
nor U21727 (N_21727,N_18477,N_16359);
or U21728 (N_21728,N_18713,N_16068);
and U21729 (N_21729,N_19106,N_16638);
and U21730 (N_21730,N_15420,N_17636);
nand U21731 (N_21731,N_15684,N_15412);
and U21732 (N_21732,N_18091,N_18028);
nor U21733 (N_21733,N_16375,N_18068);
and U21734 (N_21734,N_15957,N_17904);
or U21735 (N_21735,N_17533,N_17673);
and U21736 (N_21736,N_15889,N_17491);
nand U21737 (N_21737,N_17991,N_18124);
or U21738 (N_21738,N_18649,N_15187);
nor U21739 (N_21739,N_19135,N_17204);
nor U21740 (N_21740,N_17610,N_18733);
or U21741 (N_21741,N_19761,N_19185);
or U21742 (N_21742,N_18898,N_18674);
nor U21743 (N_21743,N_18942,N_19960);
and U21744 (N_21744,N_17126,N_17159);
nor U21745 (N_21745,N_16012,N_17751);
nand U21746 (N_21746,N_18655,N_17888);
and U21747 (N_21747,N_19984,N_17705);
nor U21748 (N_21748,N_15139,N_19213);
or U21749 (N_21749,N_16876,N_17072);
or U21750 (N_21750,N_17161,N_16160);
nor U21751 (N_21751,N_16423,N_18974);
or U21752 (N_21752,N_19430,N_16267);
or U21753 (N_21753,N_15155,N_17892);
nor U21754 (N_21754,N_17269,N_19715);
nor U21755 (N_21755,N_16362,N_19416);
nor U21756 (N_21756,N_17655,N_15129);
nand U21757 (N_21757,N_18896,N_19919);
nand U21758 (N_21758,N_17639,N_19964);
nand U21759 (N_21759,N_16431,N_16625);
nor U21760 (N_21760,N_19979,N_18745);
nor U21761 (N_21761,N_15783,N_17531);
xor U21762 (N_21762,N_19554,N_18117);
nand U21763 (N_21763,N_18691,N_17719);
nand U21764 (N_21764,N_16312,N_18390);
or U21765 (N_21765,N_19198,N_17298);
or U21766 (N_21766,N_18576,N_19138);
nand U21767 (N_21767,N_19004,N_16889);
and U21768 (N_21768,N_18557,N_19174);
nand U21769 (N_21769,N_16503,N_17030);
nand U21770 (N_21770,N_15941,N_18115);
or U21771 (N_21771,N_15182,N_15255);
and U21772 (N_21772,N_18409,N_18596);
nor U21773 (N_21773,N_19338,N_19093);
nand U21774 (N_21774,N_17066,N_19970);
nor U21775 (N_21775,N_15200,N_19383);
nand U21776 (N_21776,N_17566,N_17593);
nor U21777 (N_21777,N_18086,N_18033);
nand U21778 (N_21778,N_15012,N_18912);
nand U21779 (N_21779,N_17549,N_17186);
nor U21780 (N_21780,N_17275,N_19561);
and U21781 (N_21781,N_17385,N_17187);
and U21782 (N_21782,N_15922,N_16285);
and U21783 (N_21783,N_16912,N_19782);
and U21784 (N_21784,N_18332,N_16235);
and U21785 (N_21785,N_16609,N_17324);
nand U21786 (N_21786,N_18449,N_19854);
nor U21787 (N_21787,N_16507,N_17958);
nand U21788 (N_21788,N_19307,N_19085);
and U21789 (N_21789,N_16534,N_18534);
nor U21790 (N_21790,N_17097,N_15276);
or U21791 (N_21791,N_18538,N_15291);
and U21792 (N_21792,N_15322,N_17633);
nand U21793 (N_21793,N_19913,N_18626);
xor U21794 (N_21794,N_18229,N_16727);
nor U21795 (N_21795,N_19024,N_16796);
xnor U21796 (N_21796,N_17960,N_15442);
nand U21797 (N_21797,N_17445,N_17098);
nor U21798 (N_21798,N_18887,N_17802);
xor U21799 (N_21799,N_17730,N_15763);
nor U21800 (N_21800,N_18685,N_16683);
nand U21801 (N_21801,N_17828,N_17710);
nor U21802 (N_21802,N_17505,N_18801);
or U21803 (N_21803,N_19745,N_15999);
xor U21804 (N_21804,N_17148,N_15947);
nor U21805 (N_21805,N_16262,N_16337);
nand U21806 (N_21806,N_15904,N_15797);
and U21807 (N_21807,N_18967,N_18110);
or U21808 (N_21808,N_17062,N_16152);
or U21809 (N_21809,N_19603,N_18549);
nand U21810 (N_21810,N_19476,N_19952);
and U21811 (N_21811,N_17969,N_15592);
and U21812 (N_21812,N_16490,N_19781);
or U21813 (N_21813,N_15543,N_19095);
nor U21814 (N_21814,N_19007,N_18268);
or U21815 (N_21815,N_18282,N_19500);
and U21816 (N_21816,N_19440,N_19665);
nand U21817 (N_21817,N_19232,N_15796);
or U21818 (N_21818,N_15870,N_17749);
nand U21819 (N_21819,N_18231,N_19645);
nor U21820 (N_21820,N_16292,N_18915);
xnor U21821 (N_21821,N_18236,N_17854);
nor U21822 (N_21822,N_18593,N_17722);
or U21823 (N_21823,N_19389,N_15677);
and U21824 (N_21824,N_15868,N_15438);
and U21825 (N_21825,N_15467,N_16096);
nand U21826 (N_21826,N_16473,N_19444);
nand U21827 (N_21827,N_19779,N_15991);
nand U21828 (N_21828,N_17983,N_17160);
nor U21829 (N_21829,N_19959,N_16077);
and U21830 (N_21830,N_19635,N_17434);
nand U21831 (N_21831,N_18819,N_15573);
nand U21832 (N_21832,N_19061,N_15039);
nor U21833 (N_21833,N_18787,N_17342);
nor U21834 (N_21834,N_18575,N_17364);
nand U21835 (N_21835,N_15596,N_16119);
nor U21836 (N_21836,N_18485,N_16279);
and U21837 (N_21837,N_19879,N_15505);
nand U21838 (N_21838,N_15643,N_15863);
or U21839 (N_21839,N_18900,N_17084);
and U21840 (N_21840,N_17569,N_17932);
or U21841 (N_21841,N_16061,N_17758);
or U21842 (N_21842,N_16975,N_15333);
and U21843 (N_21843,N_16373,N_19359);
nand U21844 (N_21844,N_17390,N_15835);
nor U21845 (N_21845,N_15077,N_19931);
nand U21846 (N_21846,N_16892,N_19033);
nor U21847 (N_21847,N_19448,N_19231);
nor U21848 (N_21848,N_18336,N_16230);
nand U21849 (N_21849,N_15927,N_16347);
or U21850 (N_21850,N_19436,N_17855);
or U21851 (N_21851,N_16415,N_17215);
xor U21852 (N_21852,N_16382,N_15460);
nand U21853 (N_21853,N_19958,N_15132);
or U21854 (N_21854,N_17515,N_19372);
nor U21855 (N_21855,N_19716,N_18959);
nand U21856 (N_21856,N_16698,N_15415);
and U21857 (N_21857,N_17586,N_15964);
nor U21858 (N_21858,N_17999,N_19474);
or U21859 (N_21859,N_18832,N_16198);
or U21860 (N_21860,N_16509,N_16545);
and U21861 (N_21861,N_19143,N_19100);
or U21862 (N_21862,N_17296,N_19940);
nor U21863 (N_21863,N_17240,N_16263);
nor U21864 (N_21864,N_18267,N_15308);
nand U21865 (N_21865,N_18382,N_17008);
nand U21866 (N_21866,N_19199,N_19493);
nor U21867 (N_21867,N_17713,N_19630);
or U21868 (N_21868,N_18521,N_18109);
nand U21869 (N_21869,N_19730,N_18307);
or U21870 (N_21870,N_19028,N_19034);
nand U21871 (N_21871,N_19171,N_15609);
nand U21872 (N_21872,N_15097,N_19831);
nor U21873 (N_21873,N_17207,N_18846);
nand U21874 (N_21874,N_18056,N_18589);
or U21875 (N_21875,N_17069,N_16869);
and U21876 (N_21876,N_19809,N_15579);
or U21877 (N_21877,N_18711,N_16326);
nor U21878 (N_21878,N_19786,N_19343);
nor U21879 (N_21879,N_16531,N_17320);
or U21880 (N_21880,N_18188,N_18388);
nand U21881 (N_21881,N_18996,N_16037);
nand U21882 (N_21882,N_16005,N_16878);
or U21883 (N_21883,N_18755,N_17624);
and U21884 (N_21884,N_17061,N_16910);
or U21885 (N_21885,N_16521,N_17021);
nor U21886 (N_21886,N_19518,N_18729);
nand U21887 (N_21887,N_18546,N_16398);
or U21888 (N_21888,N_19863,N_19696);
and U21889 (N_21889,N_16155,N_19238);
or U21890 (N_21890,N_16563,N_16786);
nor U21891 (N_21891,N_19201,N_16329);
nand U21892 (N_21892,N_18253,N_19790);
nor U21893 (N_21893,N_19911,N_19144);
nand U21894 (N_21894,N_18281,N_19557);
nand U21895 (N_21895,N_17476,N_15890);
or U21896 (N_21896,N_19206,N_15515);
nor U21897 (N_21897,N_18003,N_16768);
and U21898 (N_21898,N_18982,N_16850);
nor U21899 (N_21899,N_19535,N_15951);
nand U21900 (N_21900,N_19737,N_16340);
or U21901 (N_21901,N_16022,N_19708);
nor U21902 (N_21902,N_15128,N_15456);
and U21903 (N_21903,N_16800,N_17246);
or U21904 (N_21904,N_17278,N_17294);
xnor U21905 (N_21905,N_15653,N_17425);
and U21906 (N_21906,N_19937,N_19283);
or U21907 (N_21907,N_18548,N_19344);
nand U21908 (N_21908,N_15666,N_19600);
or U21909 (N_21909,N_19284,N_19184);
and U21910 (N_21910,N_18786,N_15874);
nor U21911 (N_21911,N_19902,N_17644);
and U21912 (N_21912,N_18131,N_16499);
or U21913 (N_21913,N_18498,N_15646);
or U21914 (N_21914,N_17622,N_16881);
or U21915 (N_21915,N_17963,N_15125);
or U21916 (N_21916,N_19592,N_17233);
or U21917 (N_21917,N_15076,N_16366);
and U21918 (N_21918,N_19008,N_19042);
nor U21919 (N_21919,N_18032,N_17085);
and U21920 (N_21920,N_19018,N_19525);
nor U21921 (N_21921,N_18435,N_19423);
nor U21922 (N_21922,N_15463,N_16458);
or U21923 (N_21923,N_19735,N_15031);
and U21924 (N_21924,N_18669,N_15081);
nor U21925 (N_21925,N_19287,N_18441);
or U21926 (N_21926,N_18313,N_19292);
or U21927 (N_21927,N_17945,N_15722);
or U21928 (N_21928,N_17883,N_15488);
and U21929 (N_21929,N_18483,N_16079);
nand U21930 (N_21930,N_16902,N_19733);
nor U21931 (N_21931,N_16713,N_17274);
nor U21932 (N_21932,N_19479,N_17483);
or U21933 (N_21933,N_17595,N_19951);
and U21934 (N_21934,N_15228,N_16943);
or U21935 (N_21935,N_17534,N_16624);
and U21936 (N_21936,N_18242,N_16030);
nand U21937 (N_21937,N_15626,N_16260);
and U21938 (N_21938,N_17773,N_18893);
and U21939 (N_21939,N_17864,N_19939);
nand U21940 (N_21940,N_19586,N_17617);
nand U21941 (N_21941,N_18878,N_19705);
or U21942 (N_21942,N_16709,N_16662);
or U21943 (N_21943,N_17280,N_18249);
nand U21944 (N_21944,N_15879,N_16763);
or U21945 (N_21945,N_16945,N_17141);
nor U21946 (N_21946,N_19859,N_15083);
nand U21947 (N_21947,N_16815,N_17739);
and U21948 (N_21948,N_16227,N_19891);
nand U21949 (N_21949,N_19469,N_18720);
and U21950 (N_21950,N_15805,N_18610);
or U21951 (N_21951,N_19155,N_16529);
nand U21952 (N_21952,N_16057,N_17487);
nand U21953 (N_21953,N_15926,N_18867);
xnor U21954 (N_21954,N_16977,N_16602);
nor U21955 (N_21955,N_19183,N_19943);
and U21956 (N_21956,N_15019,N_18433);
nand U21957 (N_21957,N_19866,N_19015);
nand U21958 (N_21958,N_18998,N_16934);
or U21959 (N_21959,N_18414,N_18202);
nand U21960 (N_21960,N_15481,N_16191);
nand U21961 (N_21961,N_17536,N_17044);
and U21962 (N_21962,N_17665,N_16482);
and U21963 (N_21963,N_16722,N_16807);
and U21964 (N_21964,N_16436,N_19653);
nor U21965 (N_21965,N_16998,N_15089);
and U21966 (N_21966,N_17090,N_19580);
nand U21967 (N_21967,N_18090,N_17601);
nand U21968 (N_21968,N_16705,N_19261);
or U21969 (N_21969,N_15509,N_19355);
xnor U21970 (N_21970,N_19046,N_15589);
and U21971 (N_21971,N_18694,N_15560);
nand U21972 (N_21972,N_17372,N_17681);
or U21973 (N_21973,N_15364,N_18556);
nand U21974 (N_21974,N_16283,N_15530);
and U21975 (N_21975,N_18700,N_15799);
and U21976 (N_21976,N_17315,N_16493);
or U21977 (N_21977,N_19137,N_18369);
nor U21978 (N_21978,N_17348,N_19216);
or U21979 (N_21979,N_18999,N_19800);
nand U21980 (N_21980,N_16126,N_15728);
or U21981 (N_21981,N_15115,N_16478);
or U21982 (N_21982,N_17737,N_16315);
nor U21983 (N_21983,N_18219,N_17571);
and U21984 (N_21984,N_16099,N_16451);
nor U21985 (N_21985,N_16605,N_16072);
or U21986 (N_21986,N_15954,N_15590);
and U21987 (N_21987,N_18322,N_19208);
and U21988 (N_21988,N_16224,N_16344);
or U21989 (N_21989,N_17265,N_18747);
nor U21990 (N_21990,N_15042,N_16990);
and U21991 (N_21991,N_15224,N_19887);
nor U21992 (N_21992,N_17992,N_18807);
or U21993 (N_21993,N_16757,N_18823);
nand U21994 (N_21994,N_18207,N_16445);
and U21995 (N_21995,N_15881,N_18058);
nor U21996 (N_21996,N_16091,N_19624);
and U21997 (N_21997,N_15180,N_19966);
and U21998 (N_21998,N_18785,N_17336);
or U21999 (N_21999,N_17195,N_15901);
and U22000 (N_22000,N_15457,N_18827);
nor U22001 (N_22001,N_16559,N_17404);
nor U22002 (N_22002,N_16926,N_17779);
nand U22003 (N_22003,N_18262,N_18630);
nand U22004 (N_22004,N_15465,N_15055);
and U22005 (N_22005,N_15109,N_17266);
or U22006 (N_22006,N_16564,N_18346);
nor U22007 (N_22007,N_16656,N_19738);
and U22008 (N_22008,N_17760,N_17140);
nand U22009 (N_22009,N_15782,N_15452);
or U22010 (N_22010,N_17728,N_15651);
nor U22011 (N_22011,N_17117,N_16122);
and U22012 (N_22012,N_16816,N_19203);
nand U22013 (N_22013,N_18073,N_19315);
nor U22014 (N_22014,N_17656,N_15884);
or U22015 (N_22015,N_15117,N_17724);
and U22016 (N_22016,N_19566,N_15410);
and U22017 (N_22017,N_17133,N_17276);
nor U22018 (N_22018,N_15253,N_18632);
or U22019 (N_22019,N_16004,N_15768);
or U22020 (N_22020,N_15962,N_17418);
nand U22021 (N_22021,N_17179,N_17283);
nand U22022 (N_22022,N_15336,N_15120);
and U22023 (N_22023,N_19674,N_15426);
and U22024 (N_22024,N_19766,N_18849);
nor U22025 (N_22025,N_16328,N_17529);
or U22026 (N_22026,N_19739,N_19593);
or U22027 (N_22027,N_18992,N_17171);
nand U22028 (N_22028,N_16254,N_18101);
nor U22029 (N_22029,N_18620,N_18029);
nand U22030 (N_22030,N_19254,N_16278);
and U22031 (N_22031,N_19017,N_17443);
or U22032 (N_22032,N_15546,N_17381);
nand U22033 (N_22033,N_16655,N_16466);
nor U22034 (N_22034,N_17112,N_17631);
nor U22035 (N_22035,N_19363,N_16985);
nor U22036 (N_22036,N_17029,N_17459);
xor U22037 (N_22037,N_15301,N_16923);
nand U22038 (N_22038,N_15561,N_19467);
and U22039 (N_22039,N_18425,N_15067);
nand U22040 (N_22040,N_17252,N_17263);
nand U22041 (N_22041,N_16323,N_17486);
nand U22042 (N_22042,N_16533,N_17661);
nor U22043 (N_22043,N_15245,N_17389);
nand U22044 (N_22044,N_19036,N_19477);
or U22045 (N_22045,N_18671,N_15791);
and U22046 (N_22046,N_19816,N_17585);
and U22047 (N_22047,N_17919,N_18637);
or U22048 (N_22048,N_19267,N_17480);
nor U22049 (N_22049,N_18606,N_16578);
xnor U22050 (N_22050,N_18656,N_16066);
or U22051 (N_22051,N_18926,N_18430);
nand U22052 (N_22052,N_18527,N_15193);
or U22053 (N_22053,N_15553,N_15153);
and U22054 (N_22054,N_16983,N_18216);
and U22055 (N_22055,N_17019,N_18662);
or U22056 (N_22056,N_19218,N_18397);
and U22057 (N_22057,N_16960,N_16270);
or U22058 (N_22058,N_16736,N_18290);
xor U22059 (N_22059,N_18578,N_18296);
nand U22060 (N_22060,N_17006,N_15649);
and U22061 (N_22061,N_18187,N_15984);
nand U22062 (N_22062,N_17433,N_16767);
or U22063 (N_22063,N_17268,N_16141);
nand U22064 (N_22064,N_19803,N_16151);
nor U22065 (N_22065,N_19974,N_16295);
nand U22066 (N_22066,N_17712,N_16611);
nand U22067 (N_22067,N_16991,N_18284);
xnor U22068 (N_22068,N_15444,N_18299);
nor U22069 (N_22069,N_16476,N_15751);
nand U22070 (N_22070,N_15676,N_17092);
nor U22071 (N_22071,N_19771,N_17173);
or U22072 (N_22072,N_18734,N_19582);
nor U22073 (N_22073,N_17495,N_17587);
nand U22074 (N_22074,N_17060,N_16510);
nor U22075 (N_22075,N_18978,N_19878);
xor U22076 (N_22076,N_16195,N_17890);
and U22077 (N_22077,N_17996,N_17954);
nand U22078 (N_22078,N_16239,N_15587);
nand U22079 (N_22079,N_16064,N_18420);
and U22080 (N_22080,N_17317,N_18650);
nor U22081 (N_22081,N_15432,N_16872);
or U22082 (N_22082,N_15837,N_15414);
nand U22083 (N_22083,N_19020,N_15024);
and U22084 (N_22084,N_16298,N_15094);
nor U22085 (N_22085,N_19618,N_18035);
and U22086 (N_22086,N_17856,N_18736);
nand U22087 (N_22087,N_17472,N_16805);
nand U22088 (N_22088,N_19988,N_19787);
or U22089 (N_22089,N_16386,N_17058);
or U22090 (N_22090,N_18879,N_16249);
xnor U22091 (N_22091,N_16952,N_17508);
and U22092 (N_22092,N_16597,N_19207);
nand U22093 (N_22093,N_17345,N_19797);
or U22094 (N_22094,N_18973,N_16864);
and U22095 (N_22095,N_17970,N_17239);
nor U22096 (N_22096,N_17172,N_16775);
nor U22097 (N_22097,N_16859,N_15287);
or U22098 (N_22098,N_18809,N_16345);
and U22099 (N_22099,N_15953,N_17050);
and U22100 (N_22100,N_16762,N_15079);
nand U22101 (N_22101,N_19922,N_16219);
or U22102 (N_22102,N_15570,N_16979);
nand U22103 (N_22103,N_15489,N_15222);
and U22104 (N_22104,N_16130,N_18523);
or U22105 (N_22105,N_15845,N_19382);
nand U22106 (N_22106,N_18876,N_15058);
nand U22107 (N_22107,N_16940,N_16801);
and U22108 (N_22108,N_16581,N_19060);
or U22109 (N_22109,N_19617,N_19526);
and U22110 (N_22110,N_16231,N_17417);
nand U22111 (N_22111,N_18932,N_19563);
or U22112 (N_22112,N_15394,N_18862);
nor U22113 (N_22113,N_18205,N_15360);
and U22114 (N_22114,N_15321,N_15294);
nor U22115 (N_22115,N_15726,N_16634);
nand U22116 (N_22116,N_17489,N_15660);
and U22117 (N_22117,N_16764,N_17676);
xor U22118 (N_22118,N_19468,N_18938);
nand U22119 (N_22119,N_19402,N_17711);
or U22120 (N_22120,N_16385,N_18804);
and U22121 (N_22121,N_15382,N_17371);
or U22122 (N_22122,N_16914,N_15851);
or U22123 (N_22123,N_15396,N_16018);
or U22124 (N_22124,N_16661,N_16654);
or U22125 (N_22125,N_15701,N_16401);
nor U22126 (N_22126,N_19648,N_19140);
or U22127 (N_22127,N_17683,N_15905);
nand U22128 (N_22128,N_19056,N_18442);
and U22129 (N_22129,N_16819,N_18504);
nand U22130 (N_22130,N_16233,N_19357);
nor U22131 (N_22131,N_15306,N_17981);
nand U22132 (N_22132,N_17255,N_16144);
nor U22133 (N_22133,N_16773,N_15446);
or U22134 (N_22134,N_15770,N_18243);
and U22135 (N_22135,N_17223,N_16241);
or U22136 (N_22136,N_16994,N_16172);
nand U22137 (N_22137,N_16631,N_19917);
and U22138 (N_22138,N_19987,N_19999);
nor U22139 (N_22139,N_18856,N_19418);
or U22140 (N_22140,N_16974,N_19753);
or U22141 (N_22141,N_17581,N_17778);
and U22142 (N_22142,N_17330,N_18947);
and U22143 (N_22143,N_19992,N_18698);
nor U22144 (N_22144,N_15495,N_17527);
or U22145 (N_22145,N_16491,N_18957);
nor U22146 (N_22146,N_17466,N_15795);
nor U22147 (N_22147,N_17839,N_15871);
nor U22148 (N_22148,N_15370,N_18358);
nand U22149 (N_22149,N_16657,N_19249);
nor U22150 (N_22150,N_19604,N_19811);
or U22151 (N_22151,N_16346,N_19420);
nor U22152 (N_22152,N_17905,N_17997);
nand U22153 (N_22153,N_19631,N_18919);
nor U22154 (N_22154,N_19178,N_19695);
nor U22155 (N_22155,N_18004,N_15766);
or U22156 (N_22156,N_19333,N_15671);
nor U22157 (N_22157,N_17762,N_19349);
and U22158 (N_22158,N_16678,N_18676);
nor U22159 (N_22159,N_17145,N_17166);
or U22160 (N_22160,N_18127,N_19237);
and U22161 (N_22161,N_15256,N_16170);
or U22162 (N_22162,N_18326,N_17794);
and U22163 (N_22163,N_16070,N_16244);
nor U22164 (N_22164,N_19920,N_16953);
and U22165 (N_22165,N_16814,N_16874);
nor U22166 (N_22166,N_16369,N_19950);
nor U22167 (N_22167,N_19149,N_17952);
nor U22168 (N_22168,N_18023,N_17333);
and U22169 (N_22169,N_15015,N_19510);
nor U22170 (N_22170,N_18638,N_19780);
nand U22171 (N_22171,N_16672,N_16410);
nor U22172 (N_22172,N_16114,N_19037);
and U22173 (N_22173,N_15152,N_15163);
and U22174 (N_22174,N_18985,N_15985);
and U22175 (N_22175,N_15709,N_18149);
and U22176 (N_22176,N_16202,N_15181);
or U22177 (N_22177,N_18182,N_19360);
xor U22178 (N_22178,N_16834,N_17080);
nand U22179 (N_22179,N_15500,N_17237);
nand U22180 (N_22180,N_15548,N_18730);
or U22181 (N_22181,N_19304,N_17419);
nand U22182 (N_22182,N_16502,N_15754);
or U22183 (N_22183,N_16303,N_15071);
or U22184 (N_22184,N_17747,N_15623);
or U22185 (N_22185,N_19489,N_16044);
nor U22186 (N_22186,N_19540,N_18212);
nor U22187 (N_22187,N_18815,N_19164);
nand U22188 (N_22188,N_19567,N_19465);
and U22189 (N_22189,N_16147,N_18379);
nor U22190 (N_22190,N_15484,N_17746);
and U22191 (N_22191,N_19406,N_15987);
and U22192 (N_22192,N_17229,N_15704);
nor U22193 (N_22193,N_19606,N_16291);
and U22194 (N_22194,N_18141,N_16498);
nand U22195 (N_22195,N_18798,N_15864);
xor U22196 (N_22196,N_16526,N_18682);
nand U22197 (N_22197,N_18170,N_16982);
or U22198 (N_22198,N_18232,N_15950);
or U22199 (N_22199,N_16525,N_18509);
or U22200 (N_22200,N_17479,N_18547);
and U22201 (N_22201,N_17731,N_15707);
or U22202 (N_22202,N_18113,N_17271);
nand U22203 (N_22203,N_17267,N_18774);
nand U22204 (N_22204,N_18177,N_18197);
or U22205 (N_22205,N_17539,N_17448);
and U22206 (N_22206,N_17703,N_15459);
or U22207 (N_22207,N_18852,N_19669);
and U22208 (N_22208,N_16199,N_16557);
and U22209 (N_22209,N_18440,N_15455);
and U22210 (N_22210,N_16832,N_16237);
nor U22211 (N_22211,N_17677,N_17528);
and U22212 (N_22212,N_15018,N_19558);
nand U22213 (N_22213,N_18631,N_17184);
nand U22214 (N_22214,N_18861,N_16045);
nor U22215 (N_22215,N_19688,N_15652);
and U22216 (N_22216,N_15263,N_19317);
nand U22217 (N_22217,N_19128,N_15669);
xor U22218 (N_22218,N_17666,N_16105);
and U22219 (N_22219,N_17818,N_17382);
nor U22220 (N_22220,N_19002,N_18166);
and U22221 (N_22221,N_15437,N_15288);
and U22222 (N_22222,N_18318,N_16838);
or U22223 (N_22223,N_15439,N_19157);
nor U22224 (N_22224,N_19006,N_19482);
and U22225 (N_22225,N_15811,N_17698);
xor U22226 (N_22226,N_17073,N_16618);
and U22227 (N_22227,N_18928,N_15397);
nand U22228 (N_22228,N_16137,N_18462);
and U22229 (N_22229,N_15114,N_18377);
nand U22230 (N_22230,N_17386,N_15572);
nor U22231 (N_22231,N_18064,N_16194);
and U22232 (N_22232,N_19616,N_19728);
or U22233 (N_22233,N_18695,N_15249);
and U22234 (N_22234,N_18686,N_17107);
nor U22235 (N_22235,N_16682,N_16594);
nor U22236 (N_22236,N_15636,N_15082);
nand U22237 (N_22237,N_16600,N_18136);
and U22238 (N_22238,N_15917,N_18331);
or U22239 (N_22239,N_15300,N_15675);
and U22240 (N_22240,N_18493,N_16665);
and U22241 (N_22241,N_18481,N_17687);
nor U22242 (N_22242,N_16935,N_18735);
nor U22243 (N_22243,N_18034,N_16986);
or U22244 (N_22244,N_19817,N_17863);
or U22245 (N_22245,N_16547,N_17402);
nand U22246 (N_22246,N_17146,N_17477);
nor U22247 (N_22247,N_17206,N_18740);
nand U22248 (N_22248,N_16761,N_17220);
and U22249 (N_22249,N_17609,N_17351);
or U22250 (N_22250,N_19613,N_16135);
nor U22251 (N_22251,N_16706,N_19256);
xor U22252 (N_22252,N_18791,N_15656);
nand U22253 (N_22253,N_15427,N_16674);
nand U22254 (N_22254,N_19131,N_19594);
or U22255 (N_22255,N_19724,N_16379);
nand U22256 (N_22256,N_19949,N_16562);
nand U22257 (N_22257,N_15747,N_17408);
and U22258 (N_22258,N_19193,N_17955);
or U22259 (N_22259,N_18395,N_19928);
nand U22260 (N_22260,N_18311,N_19972);
and U22261 (N_22261,N_17129,N_18643);
xor U22262 (N_22262,N_18870,N_18078);
and U22263 (N_22263,N_16404,N_19005);
nand U22264 (N_22264,N_18918,N_19099);
or U22265 (N_22265,N_19707,N_15145);
or U22266 (N_22266,N_16236,N_17554);
xnor U22267 (N_22267,N_19268,N_19673);
nand U22268 (N_22268,N_15506,N_15558);
nor U22269 (N_22269,N_16452,N_18845);
and U22270 (N_22270,N_17886,N_18001);
nand U22271 (N_22271,N_15916,N_18813);
nand U22272 (N_22272,N_15023,N_15476);
and U22273 (N_22273,N_18288,N_15235);
nor U22274 (N_22274,N_15673,N_19513);
nor U22275 (N_22275,N_17899,N_17325);
and U22276 (N_22276,N_18666,N_16454);
and U22277 (N_22277,N_17299,N_18540);
nand U22278 (N_22278,N_15618,N_17797);
and U22279 (N_22279,N_15464,N_19633);
nand U22280 (N_22280,N_16855,N_15777);
and U22281 (N_22281,N_15254,N_18884);
nand U22282 (N_22282,N_17407,N_16041);
nor U22283 (N_22283,N_17430,N_19097);
nand U22284 (N_22284,N_15719,N_18993);
nor U22285 (N_22285,N_19810,N_17322);
or U22286 (N_22286,N_19718,N_19147);
and U22287 (N_22287,N_18227,N_15513);
and U22288 (N_22288,N_19299,N_18659);
nor U22289 (N_22289,N_15126,N_15788);
or U22290 (N_22290,N_15910,N_18163);
or U22291 (N_22291,N_18910,N_18644);
or U22292 (N_22292,N_16616,N_17321);
and U22293 (N_22293,N_19900,N_16409);
or U22294 (N_22294,N_17901,N_19490);
or U22295 (N_22295,N_16411,N_15345);
xnor U22296 (N_22296,N_17482,N_15393);
nand U22297 (N_22297,N_19955,N_16898);
nor U22298 (N_22298,N_18338,N_15063);
nor U22299 (N_22299,N_16186,N_19345);
or U22300 (N_22300,N_18759,N_16075);
or U22301 (N_22301,N_19393,N_15204);
nor U22302 (N_22302,N_19369,N_16393);
nand U22303 (N_22303,N_17493,N_18860);
and U22304 (N_22304,N_16457,N_18270);
or U22305 (N_22305,N_19607,N_18646);
nand U22306 (N_22306,N_17628,N_18247);
or U22307 (N_22307,N_18337,N_18228);
nor U22308 (N_22308,N_16097,N_19376);
and U22309 (N_22309,N_17850,N_15641);
or U22310 (N_22310,N_19520,N_18405);
and U22311 (N_22311,N_18830,N_17054);
nor U22312 (N_22312,N_16492,N_18328);
nor U22313 (N_22313,N_17313,N_15122);
and U22314 (N_22314,N_17552,N_19680);
nor U22315 (N_22315,N_15667,N_19894);
nor U22316 (N_22316,N_17205,N_16969);
nand U22317 (N_22317,N_15243,N_17565);
nand U22318 (N_22318,N_16026,N_18571);
and U22319 (N_22319,N_16419,N_16652);
nand U22320 (N_22320,N_16601,N_17065);
nand U22321 (N_22321,N_17341,N_16748);
nand U22322 (N_22322,N_18906,N_18964);
or U22323 (N_22323,N_19684,N_15876);
nor U22324 (N_22324,N_19452,N_15552);
nand U22325 (N_22325,N_19118,N_18831);
or U22326 (N_22326,N_15087,N_17659);
or U22327 (N_22327,N_17015,N_15970);
nand U22328 (N_22328,N_19495,N_19124);
nor U22329 (N_22329,N_18766,N_19938);
or U22330 (N_22330,N_17541,N_18201);
and U22331 (N_22331,N_18459,N_19129);
nand U22332 (N_22332,N_19590,N_19223);
nor U22333 (N_22333,N_18460,N_19374);
nor U22334 (N_22334,N_15313,N_16293);
nand U22335 (N_22335,N_19313,N_17152);
nand U22336 (N_22336,N_17559,N_19257);
nor U22337 (N_22337,N_17343,N_15930);
or U22338 (N_22338,N_19314,N_18595);
nand U22339 (N_22339,N_15989,N_16467);
or U22340 (N_22340,N_19330,N_18812);
nand U22341 (N_22341,N_17723,N_16595);
and U22342 (N_22342,N_16623,N_16642);
xor U22343 (N_22343,N_19833,N_15025);
nand U22344 (N_22344,N_18705,N_18164);
nor U22345 (N_22345,N_18045,N_17079);
nor U22346 (N_22346,N_17227,N_15273);
xor U22347 (N_22347,N_18826,N_17748);
or U22348 (N_22348,N_19246,N_17950);
nand U22349 (N_22349,N_18673,N_17551);
and U22350 (N_22350,N_16647,N_18066);
nor U22351 (N_22351,N_15635,N_15743);
nand U22352 (N_22352,N_16615,N_15323);
nor U22353 (N_22353,N_17464,N_19088);
or U22354 (N_22354,N_18622,N_17504);
nand U22355 (N_22355,N_19571,N_18321);
or U22356 (N_22356,N_15940,N_17154);
or U22357 (N_22357,N_17679,N_19478);
nand U22358 (N_22358,N_15792,N_19643);
or U22359 (N_22359,N_17023,N_16416);
nor U22360 (N_22360,N_19466,N_17455);
nor U22361 (N_22361,N_17678,N_19783);
or U22362 (N_22362,N_15030,N_17563);
nand U22363 (N_22363,N_19032,N_19297);
and U22364 (N_22364,N_16166,N_15100);
and U22365 (N_22365,N_15072,N_19481);
and U22366 (N_22366,N_18881,N_15681);
and U22367 (N_22367,N_18266,N_18461);
nand U22368 (N_22368,N_16520,N_16062);
nand U22369 (N_22369,N_19622,N_15116);
or U22370 (N_22370,N_18365,N_17238);
nor U22371 (N_22371,N_15275,N_17902);
nor U22372 (N_22372,N_18173,N_18808);
nor U22373 (N_22373,N_17690,N_15103);
or U22374 (N_22374,N_18661,N_19065);
nor U22375 (N_22375,N_16906,N_18312);
nor U22376 (N_22376,N_19181,N_16930);
nor U22377 (N_22377,N_18968,N_17813);
and U22378 (N_22378,N_19196,N_15400);
and U22379 (N_22379,N_16817,N_19130);
or U22380 (N_22380,N_16000,N_19655);
or U22381 (N_22381,N_18615,N_17323);
nor U22382 (N_22382,N_18952,N_18500);
nand U22383 (N_22383,N_19795,N_16029);
nor U22384 (N_22384,N_19681,N_18080);
nand U22385 (N_22385,N_18776,N_17014);
nor U22386 (N_22386,N_16899,N_17127);
and U22387 (N_22387,N_16370,N_19711);
nand U22388 (N_22388,N_18062,N_16101);
nor U22389 (N_22389,N_17081,N_18265);
or U22390 (N_22390,N_15289,N_17468);
and U22391 (N_22391,N_16861,N_15237);
nand U22392 (N_22392,N_17882,N_16187);
or U22393 (N_22393,N_15471,N_18551);
nor U22394 (N_22394,N_15029,N_18762);
nor U22395 (N_22395,N_16781,N_18263);
and U22396 (N_22396,N_16212,N_15054);
or U22397 (N_22397,N_19107,N_16697);
nand U22398 (N_22398,N_17337,N_17424);
nand U22399 (N_22399,N_17772,N_16448);
nand U22400 (N_22400,N_18404,N_17134);
and U22401 (N_22401,N_18298,N_15325);
and U22402 (N_22402,N_19092,N_16546);
nor U22403 (N_22403,N_17292,N_19356);
nor U22404 (N_22404,N_15419,N_16780);
or U22405 (N_22405,N_19487,N_17426);
and U22406 (N_22406,N_18421,N_17898);
nor U22407 (N_22407,N_16048,N_16301);
xnor U22408 (N_22408,N_19077,N_19660);
nand U22409 (N_22409,N_17176,N_15866);
nand U22410 (N_22410,N_19205,N_19514);
or U22411 (N_22411,N_16664,N_15049);
nand U22412 (N_22412,N_15577,N_19082);
and U22413 (N_22413,N_16984,N_16038);
nor U22414 (N_22414,N_16877,N_15856);
or U22415 (N_22415,N_17627,N_17649);
and U22416 (N_22416,N_15976,N_18347);
nand U22417 (N_22417,N_17331,N_17789);
nand U22418 (N_22418,N_15539,N_16196);
nor U22419 (N_22419,N_18799,N_17277);
and U22420 (N_22420,N_17272,N_18841);
nor U22421 (N_22421,N_16439,N_15591);
nand U22422 (N_22422,N_15001,N_19794);
and U22423 (N_22423,N_17859,N_17962);
nand U22424 (N_22424,N_15422,N_16193);
nor U22425 (N_22425,N_16185,N_18877);
and U22426 (N_22426,N_17810,N_15161);
nor U22427 (N_22427,N_19628,N_17435);
nand U22428 (N_22428,N_18356,N_15938);
nor U22429 (N_22429,N_18956,N_15691);
nor U22430 (N_22430,N_16165,N_18011);
nor U22431 (N_22431,N_15978,N_16794);
nand U22432 (N_22432,N_16579,N_19335);
or U22433 (N_22433,N_16432,N_17461);
nor U22434 (N_22434,N_18479,N_15062);
and U22435 (N_22435,N_18764,N_16428);
and U22436 (N_22436,N_19636,N_15324);
nand U22437 (N_22437,N_19882,N_18793);
and U22438 (N_22438,N_19898,N_16302);
nor U22439 (N_22439,N_17150,N_18399);
or U22440 (N_22440,N_18083,N_15383);
xor U22441 (N_22441,N_19933,N_19348);
nor U22442 (N_22442,N_18048,N_15831);
nand U22443 (N_22443,N_15367,N_19245);
nand U22444 (N_22444,N_16824,N_16222);
or U22445 (N_22445,N_18750,N_17025);
nand U22446 (N_22446,N_19148,N_18410);
xor U22447 (N_22447,N_18743,N_18261);
and U22448 (N_22448,N_17680,N_18217);
nand U22449 (N_22449,N_19793,N_18988);
nand U22450 (N_22450,N_15330,N_17637);
xnor U22451 (N_22451,N_15608,N_17260);
nor U22452 (N_22452,N_19985,N_18285);
nand U22453 (N_22453,N_19003,N_15828);
nand U22454 (N_22454,N_19765,N_19578);
xnor U22455 (N_22455,N_16957,N_18152);
nor U22456 (N_22456,N_18302,N_17804);
and U22457 (N_22457,N_15443,N_15159);
nor U22458 (N_22458,N_19751,N_19656);
nor U22459 (N_22459,N_17131,N_18383);
and U22460 (N_22460,N_15946,N_15918);
or U22461 (N_22461,N_16659,N_16738);
or U22462 (N_22462,N_15882,N_18490);
or U22463 (N_22463,N_16287,N_19266);
xnor U22464 (N_22464,N_19861,N_15040);
or U22465 (N_22465,N_19378,N_18256);
and U22466 (N_22466,N_18434,N_18794);
and U22467 (N_22467,N_19364,N_19090);
or U22468 (N_22468,N_18535,N_15629);
and U22469 (N_22469,N_15314,N_17494);
and U22470 (N_22470,N_15853,N_18513);
nand U22471 (N_22471,N_17990,N_17349);
and U22472 (N_22472,N_15003,N_18375);
and U22473 (N_22473,N_19598,N_18602);
and U22474 (N_22474,N_18895,N_15266);
and U22475 (N_22475,N_15877,N_18473);
nor U22476 (N_22476,N_17765,N_19968);
and U22477 (N_22477,N_16828,N_18185);
and U22478 (N_22478,N_19651,N_19640);
or U22479 (N_22479,N_16255,N_17367);
nand U22480 (N_22480,N_15277,N_15516);
and U22481 (N_22481,N_17517,N_19864);
nand U22482 (N_22482,N_15073,N_17774);
nor U22483 (N_22483,N_18514,N_17403);
or U22484 (N_22484,N_16900,N_16336);
or U22485 (N_22485,N_19916,N_17032);
and U22486 (N_22486,N_17034,N_15284);
nand U22487 (N_22487,N_19570,N_17463);
nor U22488 (N_22488,N_19387,N_15958);
nor U22489 (N_22489,N_17799,N_15113);
and U22490 (N_22490,N_17889,N_19725);
nor U22491 (N_22491,N_16384,N_15824);
or U22492 (N_22492,N_19991,N_18641);
nor U22493 (N_22493,N_18714,N_15846);
nor U22494 (N_22494,N_15545,N_19996);
xor U22495 (N_22495,N_15034,N_17365);
xnor U22496 (N_22496,N_18562,N_16033);
nor U22497 (N_22497,N_18784,N_16720);
nand U22498 (N_22498,N_18415,N_17012);
nor U22499 (N_22499,N_19511,N_19169);
nand U22500 (N_22500,N_18710,N_19915);
nor U22501 (N_22501,N_15115,N_18946);
or U22502 (N_22502,N_15634,N_18503);
or U22503 (N_22503,N_15220,N_19180);
nand U22504 (N_22504,N_16476,N_17045);
nor U22505 (N_22505,N_18784,N_16781);
nor U22506 (N_22506,N_15093,N_18026);
xnor U22507 (N_22507,N_18539,N_16222);
nand U22508 (N_22508,N_17328,N_17098);
nand U22509 (N_22509,N_17606,N_18906);
nor U22510 (N_22510,N_19138,N_19222);
nand U22511 (N_22511,N_16932,N_17944);
or U22512 (N_22512,N_15897,N_17753);
nor U22513 (N_22513,N_17245,N_16461);
or U22514 (N_22514,N_19440,N_15814);
and U22515 (N_22515,N_19450,N_17712);
and U22516 (N_22516,N_18453,N_15372);
and U22517 (N_22517,N_18327,N_16176);
nor U22518 (N_22518,N_19081,N_19702);
nor U22519 (N_22519,N_18211,N_16343);
nor U22520 (N_22520,N_18030,N_17387);
and U22521 (N_22521,N_17306,N_18626);
and U22522 (N_22522,N_16749,N_15974);
nor U22523 (N_22523,N_17679,N_17911);
and U22524 (N_22524,N_18121,N_15600);
and U22525 (N_22525,N_18440,N_17060);
nor U22526 (N_22526,N_15705,N_19136);
nor U22527 (N_22527,N_15873,N_18232);
nor U22528 (N_22528,N_15537,N_19188);
or U22529 (N_22529,N_19360,N_18078);
nand U22530 (N_22530,N_17228,N_18113);
nand U22531 (N_22531,N_16257,N_16123);
and U22532 (N_22532,N_16867,N_19946);
or U22533 (N_22533,N_18167,N_15831);
nand U22534 (N_22534,N_16736,N_17815);
and U22535 (N_22535,N_19436,N_16937);
nor U22536 (N_22536,N_18138,N_18733);
nand U22537 (N_22537,N_18671,N_15786);
and U22538 (N_22538,N_16182,N_19483);
nand U22539 (N_22539,N_15953,N_19720);
and U22540 (N_22540,N_17272,N_18342);
nand U22541 (N_22541,N_19758,N_18325);
nand U22542 (N_22542,N_17065,N_16503);
and U22543 (N_22543,N_17277,N_15045);
xnor U22544 (N_22544,N_18714,N_18172);
and U22545 (N_22545,N_16984,N_19865);
nor U22546 (N_22546,N_18063,N_18256);
nand U22547 (N_22547,N_16278,N_16286);
and U22548 (N_22548,N_19798,N_17244);
nor U22549 (N_22549,N_17645,N_15421);
and U22550 (N_22550,N_19684,N_19715);
or U22551 (N_22551,N_17020,N_18943);
nand U22552 (N_22552,N_17083,N_19547);
nor U22553 (N_22553,N_19180,N_15441);
nand U22554 (N_22554,N_15329,N_15670);
nor U22555 (N_22555,N_19167,N_19807);
nand U22556 (N_22556,N_19478,N_18255);
and U22557 (N_22557,N_18563,N_16404);
or U22558 (N_22558,N_17693,N_16656);
nor U22559 (N_22559,N_16274,N_15374);
nand U22560 (N_22560,N_15344,N_15016);
or U22561 (N_22561,N_19642,N_18795);
or U22562 (N_22562,N_16062,N_17859);
and U22563 (N_22563,N_18821,N_19039);
or U22564 (N_22564,N_18860,N_15351);
or U22565 (N_22565,N_18417,N_19136);
nand U22566 (N_22566,N_19266,N_15288);
and U22567 (N_22567,N_15359,N_16785);
and U22568 (N_22568,N_16153,N_16980);
nand U22569 (N_22569,N_17615,N_18688);
or U22570 (N_22570,N_19455,N_16903);
or U22571 (N_22571,N_17517,N_19288);
and U22572 (N_22572,N_17659,N_18618);
or U22573 (N_22573,N_15375,N_17919);
nor U22574 (N_22574,N_17507,N_16751);
or U22575 (N_22575,N_17266,N_19826);
and U22576 (N_22576,N_15104,N_19508);
and U22577 (N_22577,N_19603,N_16144);
nand U22578 (N_22578,N_15080,N_16735);
or U22579 (N_22579,N_18912,N_18051);
nand U22580 (N_22580,N_15578,N_18983);
or U22581 (N_22581,N_18573,N_17022);
nand U22582 (N_22582,N_15457,N_17288);
nand U22583 (N_22583,N_16282,N_19429);
or U22584 (N_22584,N_16891,N_16657);
nor U22585 (N_22585,N_19222,N_18379);
nor U22586 (N_22586,N_15482,N_15891);
nand U22587 (N_22587,N_17946,N_17789);
and U22588 (N_22588,N_17000,N_16632);
and U22589 (N_22589,N_15583,N_17545);
nand U22590 (N_22590,N_17625,N_19787);
or U22591 (N_22591,N_17424,N_17369);
and U22592 (N_22592,N_17107,N_17222);
nand U22593 (N_22593,N_18895,N_15356);
or U22594 (N_22594,N_16802,N_18749);
nand U22595 (N_22595,N_19891,N_18970);
or U22596 (N_22596,N_16621,N_17081);
nor U22597 (N_22597,N_16609,N_19858);
and U22598 (N_22598,N_17264,N_17060);
and U22599 (N_22599,N_17946,N_17040);
and U22600 (N_22600,N_16613,N_15199);
nor U22601 (N_22601,N_16701,N_16214);
nand U22602 (N_22602,N_18490,N_17287);
nor U22603 (N_22603,N_16545,N_15125);
nor U22604 (N_22604,N_17255,N_16497);
xor U22605 (N_22605,N_16334,N_18811);
nand U22606 (N_22606,N_15997,N_15273);
or U22607 (N_22607,N_17667,N_17353);
nand U22608 (N_22608,N_18279,N_19781);
nand U22609 (N_22609,N_18039,N_16664);
and U22610 (N_22610,N_15903,N_16756);
nor U22611 (N_22611,N_15876,N_17254);
nor U22612 (N_22612,N_18195,N_16165);
or U22613 (N_22613,N_15339,N_15169);
or U22614 (N_22614,N_19212,N_19340);
and U22615 (N_22615,N_18389,N_18677);
and U22616 (N_22616,N_18035,N_19267);
and U22617 (N_22617,N_18737,N_15893);
or U22618 (N_22618,N_16879,N_17552);
nor U22619 (N_22619,N_19575,N_19456);
nand U22620 (N_22620,N_19531,N_19164);
nor U22621 (N_22621,N_19117,N_18268);
nand U22622 (N_22622,N_17502,N_17172);
nand U22623 (N_22623,N_16516,N_18500);
nor U22624 (N_22624,N_19254,N_19277);
and U22625 (N_22625,N_15415,N_17147);
and U22626 (N_22626,N_17693,N_15992);
or U22627 (N_22627,N_17588,N_15803);
or U22628 (N_22628,N_19722,N_19076);
and U22629 (N_22629,N_18967,N_18350);
nand U22630 (N_22630,N_16014,N_17196);
nand U22631 (N_22631,N_17573,N_15629);
or U22632 (N_22632,N_17818,N_18890);
nand U22633 (N_22633,N_18482,N_18826);
nor U22634 (N_22634,N_15115,N_18980);
and U22635 (N_22635,N_18729,N_16892);
or U22636 (N_22636,N_19904,N_18062);
nor U22637 (N_22637,N_18637,N_15858);
nand U22638 (N_22638,N_15445,N_19434);
or U22639 (N_22639,N_19382,N_19502);
and U22640 (N_22640,N_19188,N_17506);
nand U22641 (N_22641,N_17608,N_17994);
and U22642 (N_22642,N_16314,N_19059);
xor U22643 (N_22643,N_15785,N_17386);
and U22644 (N_22644,N_16223,N_17075);
nor U22645 (N_22645,N_16201,N_17418);
or U22646 (N_22646,N_19810,N_19149);
and U22647 (N_22647,N_17451,N_18447);
nand U22648 (N_22648,N_19433,N_16524);
and U22649 (N_22649,N_15772,N_19632);
or U22650 (N_22650,N_15031,N_19546);
and U22651 (N_22651,N_17203,N_17790);
and U22652 (N_22652,N_16128,N_17852);
nor U22653 (N_22653,N_18827,N_18169);
nand U22654 (N_22654,N_19249,N_17647);
nand U22655 (N_22655,N_15025,N_19869);
or U22656 (N_22656,N_17855,N_16755);
and U22657 (N_22657,N_17097,N_19209);
nor U22658 (N_22658,N_17462,N_17154);
and U22659 (N_22659,N_15348,N_18747);
or U22660 (N_22660,N_15031,N_18204);
nand U22661 (N_22661,N_18467,N_16564);
and U22662 (N_22662,N_18651,N_17406);
nand U22663 (N_22663,N_19386,N_15631);
and U22664 (N_22664,N_15625,N_18017);
nand U22665 (N_22665,N_15053,N_15277);
or U22666 (N_22666,N_17260,N_15929);
or U22667 (N_22667,N_15924,N_15285);
or U22668 (N_22668,N_16591,N_17299);
nand U22669 (N_22669,N_15405,N_16392);
xor U22670 (N_22670,N_16216,N_17772);
nand U22671 (N_22671,N_15040,N_17808);
nand U22672 (N_22672,N_17297,N_16701);
nand U22673 (N_22673,N_19491,N_19881);
and U22674 (N_22674,N_16704,N_18156);
and U22675 (N_22675,N_18013,N_15006);
nor U22676 (N_22676,N_16005,N_15712);
nand U22677 (N_22677,N_16823,N_17859);
and U22678 (N_22678,N_17538,N_18059);
nor U22679 (N_22679,N_15207,N_16328);
and U22680 (N_22680,N_16096,N_19839);
and U22681 (N_22681,N_16110,N_16980);
nor U22682 (N_22682,N_16431,N_18094);
and U22683 (N_22683,N_18524,N_15428);
and U22684 (N_22684,N_19993,N_19974);
xnor U22685 (N_22685,N_15390,N_16226);
and U22686 (N_22686,N_17724,N_16697);
or U22687 (N_22687,N_19944,N_15882);
nand U22688 (N_22688,N_15420,N_19405);
nand U22689 (N_22689,N_18470,N_15202);
nand U22690 (N_22690,N_18212,N_16945);
nor U22691 (N_22691,N_17279,N_18828);
or U22692 (N_22692,N_17153,N_19447);
or U22693 (N_22693,N_18469,N_15676);
nand U22694 (N_22694,N_17669,N_17280);
or U22695 (N_22695,N_18075,N_17762);
nor U22696 (N_22696,N_15078,N_19828);
nor U22697 (N_22697,N_15018,N_16131);
nand U22698 (N_22698,N_17741,N_17558);
nand U22699 (N_22699,N_18615,N_17237);
or U22700 (N_22700,N_18766,N_15570);
and U22701 (N_22701,N_17924,N_18885);
nor U22702 (N_22702,N_16965,N_16130);
nor U22703 (N_22703,N_17067,N_16306);
nand U22704 (N_22704,N_19841,N_19899);
nor U22705 (N_22705,N_18717,N_17344);
and U22706 (N_22706,N_19294,N_17663);
or U22707 (N_22707,N_18849,N_16426);
or U22708 (N_22708,N_18839,N_17430);
nand U22709 (N_22709,N_19849,N_19018);
or U22710 (N_22710,N_18761,N_16011);
or U22711 (N_22711,N_19143,N_16339);
nor U22712 (N_22712,N_18923,N_17559);
nor U22713 (N_22713,N_16678,N_16996);
and U22714 (N_22714,N_17774,N_18779);
or U22715 (N_22715,N_18147,N_19182);
nor U22716 (N_22716,N_15115,N_15890);
and U22717 (N_22717,N_17957,N_18898);
and U22718 (N_22718,N_16437,N_15460);
or U22719 (N_22719,N_15204,N_18240);
or U22720 (N_22720,N_16542,N_19653);
nand U22721 (N_22721,N_18016,N_19919);
or U22722 (N_22722,N_16222,N_18301);
and U22723 (N_22723,N_19419,N_16868);
nor U22724 (N_22724,N_18080,N_16117);
nand U22725 (N_22725,N_19471,N_18483);
and U22726 (N_22726,N_16120,N_15742);
or U22727 (N_22727,N_19414,N_19687);
or U22728 (N_22728,N_17799,N_15073);
and U22729 (N_22729,N_15382,N_15189);
nand U22730 (N_22730,N_19801,N_18861);
or U22731 (N_22731,N_18157,N_19481);
nand U22732 (N_22732,N_16262,N_19992);
nor U22733 (N_22733,N_15578,N_17074);
or U22734 (N_22734,N_19561,N_16686);
and U22735 (N_22735,N_19774,N_16456);
xnor U22736 (N_22736,N_18801,N_17093);
nor U22737 (N_22737,N_15348,N_19765);
and U22738 (N_22738,N_17330,N_18004);
nor U22739 (N_22739,N_19435,N_17664);
nand U22740 (N_22740,N_18479,N_17470);
xnor U22741 (N_22741,N_17593,N_16276);
nand U22742 (N_22742,N_16992,N_18154);
nor U22743 (N_22743,N_17064,N_18951);
nand U22744 (N_22744,N_19848,N_16376);
and U22745 (N_22745,N_16575,N_16460);
nand U22746 (N_22746,N_19031,N_17375);
nand U22747 (N_22747,N_17312,N_18383);
or U22748 (N_22748,N_19176,N_18326);
and U22749 (N_22749,N_19343,N_19248);
nand U22750 (N_22750,N_19140,N_17928);
or U22751 (N_22751,N_16957,N_17212);
or U22752 (N_22752,N_17654,N_17538);
nor U22753 (N_22753,N_18515,N_19053);
or U22754 (N_22754,N_16096,N_19924);
nor U22755 (N_22755,N_16474,N_15517);
nor U22756 (N_22756,N_17774,N_15263);
and U22757 (N_22757,N_15124,N_19642);
nand U22758 (N_22758,N_15404,N_15207);
and U22759 (N_22759,N_15684,N_17850);
or U22760 (N_22760,N_18606,N_18943);
nand U22761 (N_22761,N_19565,N_19439);
or U22762 (N_22762,N_19536,N_17967);
and U22763 (N_22763,N_16493,N_15330);
or U22764 (N_22764,N_16296,N_18134);
and U22765 (N_22765,N_17596,N_17464);
or U22766 (N_22766,N_16519,N_16089);
or U22767 (N_22767,N_19469,N_17536);
and U22768 (N_22768,N_17366,N_19729);
and U22769 (N_22769,N_18022,N_17480);
nor U22770 (N_22770,N_18256,N_17925);
or U22771 (N_22771,N_16543,N_19278);
or U22772 (N_22772,N_18211,N_15172);
or U22773 (N_22773,N_18905,N_19612);
or U22774 (N_22774,N_15745,N_16818);
or U22775 (N_22775,N_19087,N_18966);
or U22776 (N_22776,N_17014,N_17968);
nand U22777 (N_22777,N_15054,N_16416);
nor U22778 (N_22778,N_16661,N_16515);
nor U22779 (N_22779,N_18263,N_17743);
nand U22780 (N_22780,N_18227,N_17013);
nand U22781 (N_22781,N_19542,N_17462);
nor U22782 (N_22782,N_19669,N_16513);
or U22783 (N_22783,N_18955,N_17906);
or U22784 (N_22784,N_19281,N_16419);
and U22785 (N_22785,N_15904,N_16713);
and U22786 (N_22786,N_15118,N_17233);
nor U22787 (N_22787,N_15128,N_19950);
and U22788 (N_22788,N_17324,N_15163);
and U22789 (N_22789,N_17648,N_17762);
nor U22790 (N_22790,N_18864,N_19066);
nor U22791 (N_22791,N_15467,N_16300);
nor U22792 (N_22792,N_19845,N_15687);
nor U22793 (N_22793,N_16325,N_16961);
nor U22794 (N_22794,N_16824,N_19798);
and U22795 (N_22795,N_16456,N_17085);
and U22796 (N_22796,N_15137,N_17345);
and U22797 (N_22797,N_19249,N_18937);
xor U22798 (N_22798,N_15013,N_17729);
and U22799 (N_22799,N_15411,N_15877);
and U22800 (N_22800,N_19257,N_18570);
nand U22801 (N_22801,N_15735,N_18557);
and U22802 (N_22802,N_15862,N_17850);
or U22803 (N_22803,N_19714,N_18447);
nor U22804 (N_22804,N_18657,N_19015);
and U22805 (N_22805,N_15133,N_17350);
nor U22806 (N_22806,N_19602,N_16404);
and U22807 (N_22807,N_15814,N_17140);
and U22808 (N_22808,N_17906,N_15261);
nand U22809 (N_22809,N_17814,N_18610);
or U22810 (N_22810,N_16388,N_15277);
or U22811 (N_22811,N_19933,N_17323);
or U22812 (N_22812,N_15453,N_17460);
and U22813 (N_22813,N_16876,N_18346);
and U22814 (N_22814,N_18645,N_15224);
nor U22815 (N_22815,N_17055,N_16227);
or U22816 (N_22816,N_19581,N_15882);
and U22817 (N_22817,N_19705,N_19904);
nor U22818 (N_22818,N_15853,N_15202);
or U22819 (N_22819,N_16852,N_19265);
nand U22820 (N_22820,N_19424,N_15880);
nand U22821 (N_22821,N_15484,N_19274);
and U22822 (N_22822,N_18864,N_17747);
nor U22823 (N_22823,N_17603,N_19564);
nor U22824 (N_22824,N_15761,N_16820);
and U22825 (N_22825,N_18594,N_16926);
or U22826 (N_22826,N_19456,N_16126);
nand U22827 (N_22827,N_18446,N_16468);
or U22828 (N_22828,N_18538,N_16473);
nor U22829 (N_22829,N_17461,N_19035);
and U22830 (N_22830,N_16602,N_18189);
nand U22831 (N_22831,N_18580,N_18927);
nand U22832 (N_22832,N_18529,N_17117);
nor U22833 (N_22833,N_18051,N_15703);
nand U22834 (N_22834,N_16637,N_16427);
or U22835 (N_22835,N_18311,N_16275);
or U22836 (N_22836,N_18320,N_15784);
nand U22837 (N_22837,N_17460,N_18876);
nor U22838 (N_22838,N_15887,N_17867);
nand U22839 (N_22839,N_19390,N_17258);
and U22840 (N_22840,N_15621,N_17977);
or U22841 (N_22841,N_19845,N_19489);
and U22842 (N_22842,N_16803,N_18101);
nand U22843 (N_22843,N_17393,N_18679);
or U22844 (N_22844,N_19790,N_15665);
or U22845 (N_22845,N_18087,N_17280);
or U22846 (N_22846,N_17351,N_19408);
or U22847 (N_22847,N_15063,N_18566);
or U22848 (N_22848,N_17204,N_19173);
nand U22849 (N_22849,N_18308,N_18325);
or U22850 (N_22850,N_19727,N_17846);
nor U22851 (N_22851,N_17153,N_15482);
xnor U22852 (N_22852,N_18560,N_18739);
nor U22853 (N_22853,N_17401,N_16494);
or U22854 (N_22854,N_19862,N_16700);
or U22855 (N_22855,N_18724,N_19593);
and U22856 (N_22856,N_16240,N_16669);
nor U22857 (N_22857,N_19915,N_18841);
or U22858 (N_22858,N_17229,N_18027);
or U22859 (N_22859,N_19720,N_18290);
nor U22860 (N_22860,N_15412,N_16921);
nor U22861 (N_22861,N_16846,N_15168);
nand U22862 (N_22862,N_17864,N_15844);
nand U22863 (N_22863,N_18647,N_16563);
or U22864 (N_22864,N_18383,N_19060);
or U22865 (N_22865,N_15122,N_17273);
or U22866 (N_22866,N_18535,N_16230);
or U22867 (N_22867,N_15071,N_17318);
and U22868 (N_22868,N_16924,N_16870);
or U22869 (N_22869,N_17550,N_18362);
nand U22870 (N_22870,N_18199,N_17688);
or U22871 (N_22871,N_16304,N_18086);
or U22872 (N_22872,N_17649,N_19304);
nor U22873 (N_22873,N_15240,N_16867);
nand U22874 (N_22874,N_19590,N_19229);
nor U22875 (N_22875,N_17290,N_18398);
or U22876 (N_22876,N_19179,N_17097);
nand U22877 (N_22877,N_19798,N_19410);
and U22878 (N_22878,N_16381,N_15899);
and U22879 (N_22879,N_17510,N_18242);
nand U22880 (N_22880,N_19661,N_19980);
and U22881 (N_22881,N_17317,N_19584);
nand U22882 (N_22882,N_19215,N_19775);
and U22883 (N_22883,N_19549,N_19660);
and U22884 (N_22884,N_16405,N_17444);
or U22885 (N_22885,N_18044,N_17708);
and U22886 (N_22886,N_19372,N_16095);
xor U22887 (N_22887,N_18942,N_15160);
or U22888 (N_22888,N_17403,N_18399);
and U22889 (N_22889,N_15513,N_17619);
or U22890 (N_22890,N_16622,N_19662);
nor U22891 (N_22891,N_17678,N_17275);
nor U22892 (N_22892,N_19385,N_19233);
or U22893 (N_22893,N_18052,N_16667);
nor U22894 (N_22894,N_19298,N_17021);
and U22895 (N_22895,N_15484,N_17139);
and U22896 (N_22896,N_18927,N_16703);
or U22897 (N_22897,N_16779,N_15423);
and U22898 (N_22898,N_16779,N_19932);
or U22899 (N_22899,N_17946,N_18220);
nor U22900 (N_22900,N_18997,N_18377);
or U22901 (N_22901,N_15555,N_19371);
and U22902 (N_22902,N_15687,N_17177);
nor U22903 (N_22903,N_15319,N_19456);
nand U22904 (N_22904,N_19744,N_16943);
or U22905 (N_22905,N_15584,N_16917);
or U22906 (N_22906,N_19127,N_16407);
or U22907 (N_22907,N_15214,N_19556);
and U22908 (N_22908,N_17086,N_17965);
or U22909 (N_22909,N_19037,N_17390);
and U22910 (N_22910,N_18049,N_16601);
nor U22911 (N_22911,N_16421,N_15337);
or U22912 (N_22912,N_16116,N_16618);
nor U22913 (N_22913,N_19555,N_16933);
nor U22914 (N_22914,N_15352,N_18472);
nand U22915 (N_22915,N_15202,N_16208);
nand U22916 (N_22916,N_16787,N_15578);
nand U22917 (N_22917,N_18449,N_17190);
or U22918 (N_22918,N_19979,N_19348);
nand U22919 (N_22919,N_16836,N_16756);
nor U22920 (N_22920,N_16433,N_15962);
and U22921 (N_22921,N_19967,N_17518);
nor U22922 (N_22922,N_17061,N_18725);
nand U22923 (N_22923,N_19603,N_15667);
nor U22924 (N_22924,N_18359,N_18567);
or U22925 (N_22925,N_19610,N_19703);
and U22926 (N_22926,N_16039,N_17219);
or U22927 (N_22927,N_15555,N_19440);
and U22928 (N_22928,N_15193,N_19991);
nand U22929 (N_22929,N_19078,N_19055);
and U22930 (N_22930,N_17682,N_19302);
and U22931 (N_22931,N_19599,N_15051);
nor U22932 (N_22932,N_15999,N_15182);
or U22933 (N_22933,N_15030,N_19719);
xnor U22934 (N_22934,N_17598,N_16068);
or U22935 (N_22935,N_15469,N_15633);
and U22936 (N_22936,N_17756,N_15427);
nand U22937 (N_22937,N_19903,N_18563);
or U22938 (N_22938,N_16323,N_15939);
and U22939 (N_22939,N_19275,N_15915);
xor U22940 (N_22940,N_18770,N_15052);
or U22941 (N_22941,N_16186,N_15636);
nor U22942 (N_22942,N_16484,N_15036);
nor U22943 (N_22943,N_16319,N_19086);
nand U22944 (N_22944,N_18653,N_17670);
nor U22945 (N_22945,N_19022,N_15815);
nor U22946 (N_22946,N_15992,N_18322);
and U22947 (N_22947,N_18188,N_17264);
nand U22948 (N_22948,N_18373,N_16988);
nand U22949 (N_22949,N_18793,N_16662);
xnor U22950 (N_22950,N_18629,N_15747);
nor U22951 (N_22951,N_17906,N_19625);
and U22952 (N_22952,N_18424,N_15031);
nor U22953 (N_22953,N_16805,N_18371);
nand U22954 (N_22954,N_16976,N_15163);
or U22955 (N_22955,N_16838,N_17771);
nor U22956 (N_22956,N_16040,N_16685);
nor U22957 (N_22957,N_15989,N_15271);
nor U22958 (N_22958,N_18059,N_17078);
and U22959 (N_22959,N_18953,N_19901);
and U22960 (N_22960,N_19890,N_17513);
or U22961 (N_22961,N_19643,N_18826);
or U22962 (N_22962,N_19398,N_19827);
xor U22963 (N_22963,N_19784,N_17450);
and U22964 (N_22964,N_16340,N_15565);
and U22965 (N_22965,N_17107,N_19215);
and U22966 (N_22966,N_18181,N_18969);
nor U22967 (N_22967,N_19615,N_15924);
or U22968 (N_22968,N_16994,N_16463);
and U22969 (N_22969,N_18474,N_16414);
nand U22970 (N_22970,N_19335,N_19122);
and U22971 (N_22971,N_17715,N_15602);
nor U22972 (N_22972,N_15963,N_19463);
or U22973 (N_22973,N_16594,N_17017);
or U22974 (N_22974,N_17735,N_18652);
and U22975 (N_22975,N_19041,N_19149);
nand U22976 (N_22976,N_16532,N_17120);
or U22977 (N_22977,N_19595,N_19771);
nand U22978 (N_22978,N_16062,N_17351);
or U22979 (N_22979,N_18305,N_17462);
nand U22980 (N_22980,N_15652,N_16638);
nand U22981 (N_22981,N_18746,N_17092);
nand U22982 (N_22982,N_16113,N_18773);
and U22983 (N_22983,N_15896,N_18445);
nand U22984 (N_22984,N_15777,N_17998);
nor U22985 (N_22985,N_19247,N_18107);
or U22986 (N_22986,N_18394,N_18946);
nand U22987 (N_22987,N_19808,N_18815);
and U22988 (N_22988,N_16001,N_18426);
nor U22989 (N_22989,N_19958,N_15006);
and U22990 (N_22990,N_15445,N_18259);
nand U22991 (N_22991,N_16569,N_19522);
nand U22992 (N_22992,N_16543,N_16569);
nor U22993 (N_22993,N_15768,N_19442);
xor U22994 (N_22994,N_19222,N_17675);
and U22995 (N_22995,N_19480,N_18458);
nor U22996 (N_22996,N_19150,N_17217);
and U22997 (N_22997,N_15622,N_19302);
or U22998 (N_22998,N_19297,N_15595);
nor U22999 (N_22999,N_18889,N_16929);
and U23000 (N_23000,N_18974,N_18411);
nand U23001 (N_23001,N_18250,N_17790);
nor U23002 (N_23002,N_15149,N_19931);
and U23003 (N_23003,N_15125,N_15827);
and U23004 (N_23004,N_15532,N_19974);
or U23005 (N_23005,N_18514,N_15715);
nand U23006 (N_23006,N_16933,N_18741);
nor U23007 (N_23007,N_17764,N_15280);
nand U23008 (N_23008,N_15183,N_16086);
nor U23009 (N_23009,N_17177,N_19827);
or U23010 (N_23010,N_15958,N_18222);
and U23011 (N_23011,N_16150,N_16522);
nand U23012 (N_23012,N_15169,N_19365);
nand U23013 (N_23013,N_15794,N_15209);
nor U23014 (N_23014,N_16117,N_17533);
or U23015 (N_23015,N_17017,N_18777);
nand U23016 (N_23016,N_17674,N_17775);
nand U23017 (N_23017,N_16856,N_19815);
or U23018 (N_23018,N_15860,N_18556);
nand U23019 (N_23019,N_16631,N_17611);
nor U23020 (N_23020,N_18278,N_18391);
or U23021 (N_23021,N_16541,N_15879);
and U23022 (N_23022,N_19056,N_19941);
nor U23023 (N_23023,N_18611,N_19309);
nor U23024 (N_23024,N_19053,N_17664);
and U23025 (N_23025,N_17981,N_19088);
and U23026 (N_23026,N_16051,N_17542);
nor U23027 (N_23027,N_16233,N_18914);
nor U23028 (N_23028,N_19009,N_15291);
nand U23029 (N_23029,N_18225,N_15891);
nand U23030 (N_23030,N_16452,N_19105);
or U23031 (N_23031,N_19675,N_17515);
nor U23032 (N_23032,N_18407,N_18095);
or U23033 (N_23033,N_16866,N_16331);
nor U23034 (N_23034,N_15462,N_17272);
or U23035 (N_23035,N_17587,N_15670);
or U23036 (N_23036,N_15739,N_19273);
nor U23037 (N_23037,N_19742,N_18387);
or U23038 (N_23038,N_18778,N_17654);
nor U23039 (N_23039,N_16115,N_15753);
nor U23040 (N_23040,N_17244,N_15707);
nor U23041 (N_23041,N_19019,N_16537);
nor U23042 (N_23042,N_17289,N_19527);
and U23043 (N_23043,N_19717,N_15602);
nand U23044 (N_23044,N_16808,N_18672);
and U23045 (N_23045,N_15530,N_17828);
nand U23046 (N_23046,N_19185,N_19953);
nor U23047 (N_23047,N_18343,N_18835);
or U23048 (N_23048,N_17576,N_18783);
nand U23049 (N_23049,N_17162,N_17231);
or U23050 (N_23050,N_19110,N_16614);
or U23051 (N_23051,N_18737,N_19195);
nor U23052 (N_23052,N_19247,N_15298);
nor U23053 (N_23053,N_18337,N_16035);
and U23054 (N_23054,N_15267,N_15665);
and U23055 (N_23055,N_16780,N_18401);
and U23056 (N_23056,N_18961,N_18817);
and U23057 (N_23057,N_16635,N_17712);
nand U23058 (N_23058,N_17388,N_17254);
nand U23059 (N_23059,N_15333,N_16409);
nand U23060 (N_23060,N_16446,N_18132);
nand U23061 (N_23061,N_15592,N_18274);
and U23062 (N_23062,N_19581,N_19092);
nand U23063 (N_23063,N_15240,N_16654);
nand U23064 (N_23064,N_15308,N_16660);
nor U23065 (N_23065,N_18668,N_15277);
nor U23066 (N_23066,N_19425,N_18497);
and U23067 (N_23067,N_17677,N_16439);
and U23068 (N_23068,N_15148,N_16778);
or U23069 (N_23069,N_16057,N_15611);
xnor U23070 (N_23070,N_17334,N_15181);
and U23071 (N_23071,N_19132,N_17534);
or U23072 (N_23072,N_17601,N_17804);
nand U23073 (N_23073,N_15262,N_19328);
or U23074 (N_23074,N_17571,N_15585);
nand U23075 (N_23075,N_15606,N_17816);
or U23076 (N_23076,N_17774,N_17211);
nand U23077 (N_23077,N_16765,N_19874);
nand U23078 (N_23078,N_19772,N_16634);
or U23079 (N_23079,N_19696,N_15884);
and U23080 (N_23080,N_17306,N_17879);
nor U23081 (N_23081,N_17407,N_15010);
or U23082 (N_23082,N_19230,N_19567);
nor U23083 (N_23083,N_19089,N_16538);
or U23084 (N_23084,N_18997,N_19381);
or U23085 (N_23085,N_15340,N_18857);
nand U23086 (N_23086,N_16419,N_16508);
nor U23087 (N_23087,N_15205,N_18669);
and U23088 (N_23088,N_18321,N_19052);
or U23089 (N_23089,N_15296,N_16704);
and U23090 (N_23090,N_17056,N_18710);
and U23091 (N_23091,N_15719,N_15532);
or U23092 (N_23092,N_15922,N_18110);
and U23093 (N_23093,N_18975,N_18948);
nand U23094 (N_23094,N_16783,N_16029);
or U23095 (N_23095,N_18905,N_19232);
nand U23096 (N_23096,N_19774,N_18829);
or U23097 (N_23097,N_17234,N_15530);
and U23098 (N_23098,N_16444,N_17766);
or U23099 (N_23099,N_16439,N_17570);
nand U23100 (N_23100,N_18544,N_15102);
nand U23101 (N_23101,N_15587,N_17500);
or U23102 (N_23102,N_16282,N_16698);
nor U23103 (N_23103,N_17181,N_16980);
and U23104 (N_23104,N_15460,N_15040);
or U23105 (N_23105,N_19749,N_18614);
and U23106 (N_23106,N_17232,N_15370);
nand U23107 (N_23107,N_17527,N_15615);
and U23108 (N_23108,N_16333,N_17305);
or U23109 (N_23109,N_18484,N_17515);
nand U23110 (N_23110,N_16215,N_15899);
and U23111 (N_23111,N_17455,N_16831);
or U23112 (N_23112,N_17168,N_19798);
nand U23113 (N_23113,N_17463,N_17775);
nor U23114 (N_23114,N_17838,N_15968);
nand U23115 (N_23115,N_16593,N_16603);
nor U23116 (N_23116,N_15289,N_18119);
and U23117 (N_23117,N_15916,N_15085);
and U23118 (N_23118,N_15396,N_18073);
nor U23119 (N_23119,N_19305,N_18099);
and U23120 (N_23120,N_16762,N_15073);
and U23121 (N_23121,N_19553,N_19716);
nand U23122 (N_23122,N_19585,N_16422);
nor U23123 (N_23123,N_19935,N_17488);
nor U23124 (N_23124,N_17790,N_16685);
nand U23125 (N_23125,N_17182,N_18797);
nor U23126 (N_23126,N_19683,N_15445);
and U23127 (N_23127,N_19060,N_17751);
nor U23128 (N_23128,N_17143,N_16438);
or U23129 (N_23129,N_19435,N_19427);
nor U23130 (N_23130,N_16834,N_17868);
nor U23131 (N_23131,N_17675,N_16036);
or U23132 (N_23132,N_16067,N_17946);
nor U23133 (N_23133,N_17851,N_15106);
nor U23134 (N_23134,N_17773,N_15087);
and U23135 (N_23135,N_16127,N_16260);
or U23136 (N_23136,N_16042,N_15470);
nor U23137 (N_23137,N_16887,N_19766);
and U23138 (N_23138,N_18363,N_17004);
nand U23139 (N_23139,N_15424,N_18492);
nor U23140 (N_23140,N_16975,N_15122);
and U23141 (N_23141,N_15301,N_18647);
and U23142 (N_23142,N_18352,N_18554);
nor U23143 (N_23143,N_19234,N_16971);
nor U23144 (N_23144,N_16962,N_15300);
and U23145 (N_23145,N_18481,N_19437);
nor U23146 (N_23146,N_18120,N_18959);
or U23147 (N_23147,N_15982,N_16260);
nand U23148 (N_23148,N_19463,N_15334);
nor U23149 (N_23149,N_18508,N_15861);
or U23150 (N_23150,N_16073,N_16294);
or U23151 (N_23151,N_17493,N_15223);
or U23152 (N_23152,N_15199,N_16686);
and U23153 (N_23153,N_18521,N_18577);
nor U23154 (N_23154,N_18143,N_16998);
nand U23155 (N_23155,N_17547,N_17765);
nand U23156 (N_23156,N_17717,N_16461);
or U23157 (N_23157,N_18190,N_17853);
or U23158 (N_23158,N_19443,N_18662);
nor U23159 (N_23159,N_16774,N_17153);
nor U23160 (N_23160,N_19120,N_16390);
and U23161 (N_23161,N_19265,N_16696);
nand U23162 (N_23162,N_19249,N_15201);
nor U23163 (N_23163,N_17574,N_16324);
nand U23164 (N_23164,N_16540,N_18609);
and U23165 (N_23165,N_16163,N_15809);
nor U23166 (N_23166,N_16186,N_15546);
or U23167 (N_23167,N_17519,N_15114);
nand U23168 (N_23168,N_17921,N_19556);
and U23169 (N_23169,N_15549,N_19657);
or U23170 (N_23170,N_16179,N_16510);
or U23171 (N_23171,N_17673,N_17496);
and U23172 (N_23172,N_16291,N_18092);
and U23173 (N_23173,N_18132,N_15644);
nand U23174 (N_23174,N_15039,N_15416);
nor U23175 (N_23175,N_17748,N_18431);
and U23176 (N_23176,N_15959,N_19170);
nor U23177 (N_23177,N_16528,N_15154);
xor U23178 (N_23178,N_19281,N_16750);
and U23179 (N_23179,N_17268,N_16377);
nand U23180 (N_23180,N_19271,N_16842);
or U23181 (N_23181,N_18205,N_15689);
and U23182 (N_23182,N_19441,N_18567);
nand U23183 (N_23183,N_19973,N_17713);
or U23184 (N_23184,N_18396,N_19487);
or U23185 (N_23185,N_19357,N_19382);
and U23186 (N_23186,N_16165,N_18932);
nor U23187 (N_23187,N_19472,N_15937);
nor U23188 (N_23188,N_15276,N_17175);
nand U23189 (N_23189,N_19930,N_19966);
and U23190 (N_23190,N_17326,N_15428);
nor U23191 (N_23191,N_18751,N_18526);
nor U23192 (N_23192,N_15352,N_15368);
or U23193 (N_23193,N_16857,N_19774);
or U23194 (N_23194,N_18183,N_17217);
or U23195 (N_23195,N_18753,N_16985);
nand U23196 (N_23196,N_17371,N_16476);
nand U23197 (N_23197,N_17183,N_17814);
xnor U23198 (N_23198,N_19695,N_15871);
nand U23199 (N_23199,N_15120,N_15077);
or U23200 (N_23200,N_16966,N_17447);
and U23201 (N_23201,N_18437,N_15081);
and U23202 (N_23202,N_17849,N_16406);
or U23203 (N_23203,N_18280,N_19552);
nand U23204 (N_23204,N_19102,N_16393);
nor U23205 (N_23205,N_16659,N_17202);
nor U23206 (N_23206,N_16958,N_18084);
and U23207 (N_23207,N_17148,N_15120);
and U23208 (N_23208,N_15729,N_16315);
and U23209 (N_23209,N_18916,N_19093);
and U23210 (N_23210,N_17956,N_18555);
nand U23211 (N_23211,N_18516,N_16493);
or U23212 (N_23212,N_17457,N_16866);
and U23213 (N_23213,N_17735,N_18039);
nor U23214 (N_23214,N_19391,N_15137);
or U23215 (N_23215,N_16824,N_15956);
or U23216 (N_23216,N_17743,N_19289);
and U23217 (N_23217,N_16049,N_19484);
or U23218 (N_23218,N_15249,N_18382);
and U23219 (N_23219,N_17443,N_15709);
or U23220 (N_23220,N_15539,N_17042);
nor U23221 (N_23221,N_19829,N_15650);
nor U23222 (N_23222,N_17412,N_19908);
and U23223 (N_23223,N_17639,N_15882);
and U23224 (N_23224,N_18797,N_16873);
and U23225 (N_23225,N_16351,N_16218);
or U23226 (N_23226,N_19720,N_18251);
or U23227 (N_23227,N_15469,N_19137);
nand U23228 (N_23228,N_18449,N_18685);
and U23229 (N_23229,N_17195,N_15869);
nor U23230 (N_23230,N_19569,N_18573);
nor U23231 (N_23231,N_16285,N_18155);
or U23232 (N_23232,N_16179,N_19850);
nand U23233 (N_23233,N_19570,N_15191);
and U23234 (N_23234,N_15664,N_17637);
nor U23235 (N_23235,N_17581,N_18279);
nand U23236 (N_23236,N_16880,N_17054);
nand U23237 (N_23237,N_18228,N_15770);
or U23238 (N_23238,N_16140,N_16484);
or U23239 (N_23239,N_17442,N_17739);
nor U23240 (N_23240,N_18332,N_17401);
nor U23241 (N_23241,N_19503,N_18755);
nand U23242 (N_23242,N_15616,N_18951);
and U23243 (N_23243,N_15492,N_16168);
nand U23244 (N_23244,N_17873,N_17345);
nor U23245 (N_23245,N_17940,N_18707);
or U23246 (N_23246,N_17829,N_18997);
or U23247 (N_23247,N_18954,N_16712);
and U23248 (N_23248,N_15271,N_17669);
nand U23249 (N_23249,N_16589,N_18404);
nor U23250 (N_23250,N_17038,N_17879);
or U23251 (N_23251,N_17641,N_15805);
nand U23252 (N_23252,N_18128,N_19795);
nand U23253 (N_23253,N_19176,N_16357);
and U23254 (N_23254,N_18194,N_15460);
nand U23255 (N_23255,N_18895,N_16980);
nor U23256 (N_23256,N_17921,N_16593);
and U23257 (N_23257,N_15560,N_18434);
nor U23258 (N_23258,N_18388,N_19471);
xor U23259 (N_23259,N_18960,N_19894);
and U23260 (N_23260,N_16374,N_15836);
and U23261 (N_23261,N_18934,N_15549);
nand U23262 (N_23262,N_19078,N_18354);
and U23263 (N_23263,N_19503,N_18828);
or U23264 (N_23264,N_18201,N_19093);
nand U23265 (N_23265,N_18636,N_18133);
or U23266 (N_23266,N_18921,N_16458);
and U23267 (N_23267,N_15693,N_15032);
nor U23268 (N_23268,N_15625,N_16040);
or U23269 (N_23269,N_15514,N_18849);
and U23270 (N_23270,N_19716,N_18282);
and U23271 (N_23271,N_19034,N_15699);
nor U23272 (N_23272,N_17668,N_15427);
xor U23273 (N_23273,N_18088,N_19859);
and U23274 (N_23274,N_17269,N_17300);
nand U23275 (N_23275,N_15267,N_16894);
xnor U23276 (N_23276,N_16363,N_15280);
and U23277 (N_23277,N_18713,N_15140);
nand U23278 (N_23278,N_19092,N_16433);
or U23279 (N_23279,N_19084,N_19385);
or U23280 (N_23280,N_19412,N_18475);
and U23281 (N_23281,N_18149,N_18926);
xor U23282 (N_23282,N_17007,N_16591);
or U23283 (N_23283,N_16867,N_18480);
nand U23284 (N_23284,N_19035,N_16683);
or U23285 (N_23285,N_16652,N_18617);
and U23286 (N_23286,N_16238,N_19612);
and U23287 (N_23287,N_16901,N_15541);
xnor U23288 (N_23288,N_18407,N_19655);
nand U23289 (N_23289,N_17570,N_17630);
or U23290 (N_23290,N_15643,N_17227);
nor U23291 (N_23291,N_17921,N_15227);
nor U23292 (N_23292,N_15366,N_17848);
nor U23293 (N_23293,N_15254,N_19232);
or U23294 (N_23294,N_18297,N_16255);
nand U23295 (N_23295,N_17806,N_17819);
or U23296 (N_23296,N_19734,N_16149);
nor U23297 (N_23297,N_18777,N_19990);
nand U23298 (N_23298,N_16780,N_18154);
nor U23299 (N_23299,N_17135,N_15528);
nand U23300 (N_23300,N_15293,N_17505);
and U23301 (N_23301,N_19119,N_16339);
and U23302 (N_23302,N_18818,N_17662);
or U23303 (N_23303,N_17598,N_19822);
nand U23304 (N_23304,N_16628,N_15168);
nand U23305 (N_23305,N_15021,N_17768);
nand U23306 (N_23306,N_17283,N_19233);
nor U23307 (N_23307,N_16461,N_17628);
and U23308 (N_23308,N_17506,N_17513);
nor U23309 (N_23309,N_15635,N_16347);
or U23310 (N_23310,N_16875,N_17843);
nand U23311 (N_23311,N_18383,N_19734);
nor U23312 (N_23312,N_18860,N_17266);
and U23313 (N_23313,N_19786,N_19873);
or U23314 (N_23314,N_15852,N_15979);
nand U23315 (N_23315,N_16205,N_19686);
nand U23316 (N_23316,N_17615,N_16735);
or U23317 (N_23317,N_18660,N_16093);
nand U23318 (N_23318,N_18753,N_19208);
nor U23319 (N_23319,N_17404,N_17029);
xnor U23320 (N_23320,N_19562,N_18096);
and U23321 (N_23321,N_17597,N_15676);
and U23322 (N_23322,N_18314,N_15350);
or U23323 (N_23323,N_15392,N_15886);
nand U23324 (N_23324,N_15681,N_17329);
or U23325 (N_23325,N_17249,N_16048);
nand U23326 (N_23326,N_17633,N_17505);
and U23327 (N_23327,N_17812,N_16583);
or U23328 (N_23328,N_16633,N_18839);
and U23329 (N_23329,N_18349,N_15705);
nor U23330 (N_23330,N_16808,N_17022);
nand U23331 (N_23331,N_19726,N_16895);
xor U23332 (N_23332,N_16144,N_18605);
nand U23333 (N_23333,N_18223,N_18375);
and U23334 (N_23334,N_16576,N_16114);
or U23335 (N_23335,N_18213,N_17261);
or U23336 (N_23336,N_16867,N_16850);
and U23337 (N_23337,N_18730,N_19127);
and U23338 (N_23338,N_19280,N_17936);
and U23339 (N_23339,N_17050,N_18131);
nor U23340 (N_23340,N_16490,N_17636);
or U23341 (N_23341,N_17004,N_16667);
xor U23342 (N_23342,N_19289,N_16681);
nand U23343 (N_23343,N_15254,N_17478);
nand U23344 (N_23344,N_18430,N_15364);
nand U23345 (N_23345,N_17954,N_19759);
nor U23346 (N_23346,N_17533,N_19536);
and U23347 (N_23347,N_19088,N_17286);
and U23348 (N_23348,N_18760,N_17051);
and U23349 (N_23349,N_17875,N_17514);
or U23350 (N_23350,N_16766,N_18965);
nor U23351 (N_23351,N_15133,N_19205);
and U23352 (N_23352,N_17924,N_17560);
or U23353 (N_23353,N_15432,N_17979);
and U23354 (N_23354,N_18260,N_17581);
and U23355 (N_23355,N_15593,N_18170);
nor U23356 (N_23356,N_17824,N_19003);
or U23357 (N_23357,N_19349,N_16566);
or U23358 (N_23358,N_16243,N_17740);
and U23359 (N_23359,N_16387,N_17175);
nor U23360 (N_23360,N_16473,N_18069);
or U23361 (N_23361,N_19264,N_18703);
and U23362 (N_23362,N_18712,N_15183);
nor U23363 (N_23363,N_16201,N_17781);
nand U23364 (N_23364,N_18993,N_15272);
nand U23365 (N_23365,N_18514,N_17637);
and U23366 (N_23366,N_17150,N_16666);
nand U23367 (N_23367,N_15778,N_19232);
and U23368 (N_23368,N_18068,N_16078);
nor U23369 (N_23369,N_15015,N_18397);
or U23370 (N_23370,N_16452,N_18327);
and U23371 (N_23371,N_15320,N_16693);
nand U23372 (N_23372,N_18028,N_19748);
and U23373 (N_23373,N_16992,N_16324);
nor U23374 (N_23374,N_18181,N_18252);
and U23375 (N_23375,N_17840,N_18106);
nor U23376 (N_23376,N_15985,N_17911);
nand U23377 (N_23377,N_19576,N_19381);
or U23378 (N_23378,N_16656,N_15662);
nor U23379 (N_23379,N_17590,N_16671);
nand U23380 (N_23380,N_16501,N_19218);
nor U23381 (N_23381,N_15863,N_19527);
nor U23382 (N_23382,N_15007,N_16777);
nor U23383 (N_23383,N_15178,N_18470);
nand U23384 (N_23384,N_15419,N_19719);
nand U23385 (N_23385,N_17386,N_16603);
nand U23386 (N_23386,N_15851,N_16844);
nand U23387 (N_23387,N_18719,N_17920);
nor U23388 (N_23388,N_19835,N_17149);
nand U23389 (N_23389,N_19778,N_18055);
and U23390 (N_23390,N_17101,N_15260);
or U23391 (N_23391,N_16630,N_18128);
or U23392 (N_23392,N_19856,N_19356);
or U23393 (N_23393,N_16415,N_18359);
nor U23394 (N_23394,N_15341,N_18265);
nand U23395 (N_23395,N_17633,N_15472);
and U23396 (N_23396,N_17564,N_19067);
and U23397 (N_23397,N_18732,N_17375);
nand U23398 (N_23398,N_17011,N_19795);
nor U23399 (N_23399,N_18640,N_15708);
nand U23400 (N_23400,N_18132,N_17063);
and U23401 (N_23401,N_19830,N_17523);
nor U23402 (N_23402,N_15139,N_15791);
nor U23403 (N_23403,N_16071,N_15674);
nor U23404 (N_23404,N_16224,N_17479);
nand U23405 (N_23405,N_18638,N_15902);
or U23406 (N_23406,N_17055,N_18113);
and U23407 (N_23407,N_18256,N_17685);
nand U23408 (N_23408,N_18757,N_16086);
nand U23409 (N_23409,N_15620,N_19061);
nor U23410 (N_23410,N_19510,N_17695);
nand U23411 (N_23411,N_15233,N_16875);
nand U23412 (N_23412,N_17771,N_15721);
nand U23413 (N_23413,N_17659,N_17919);
and U23414 (N_23414,N_17910,N_19353);
or U23415 (N_23415,N_15630,N_16452);
nor U23416 (N_23416,N_19867,N_17993);
and U23417 (N_23417,N_17028,N_16563);
nand U23418 (N_23418,N_18373,N_15593);
and U23419 (N_23419,N_17514,N_18835);
or U23420 (N_23420,N_17879,N_15377);
nand U23421 (N_23421,N_16078,N_15772);
nand U23422 (N_23422,N_18426,N_16802);
nand U23423 (N_23423,N_15949,N_15007);
or U23424 (N_23424,N_18993,N_16708);
nor U23425 (N_23425,N_16201,N_15740);
or U23426 (N_23426,N_15282,N_19968);
and U23427 (N_23427,N_19979,N_15629);
nand U23428 (N_23428,N_16808,N_18116);
or U23429 (N_23429,N_15633,N_15767);
and U23430 (N_23430,N_19027,N_16359);
nor U23431 (N_23431,N_18497,N_17566);
nand U23432 (N_23432,N_16263,N_18495);
and U23433 (N_23433,N_17053,N_19883);
and U23434 (N_23434,N_18590,N_17891);
and U23435 (N_23435,N_16560,N_19687);
nor U23436 (N_23436,N_19679,N_17382);
and U23437 (N_23437,N_18350,N_19408);
and U23438 (N_23438,N_17235,N_17244);
nor U23439 (N_23439,N_17762,N_19923);
nand U23440 (N_23440,N_18339,N_17961);
nor U23441 (N_23441,N_19729,N_19537);
or U23442 (N_23442,N_18953,N_18879);
nor U23443 (N_23443,N_19158,N_17706);
nor U23444 (N_23444,N_17487,N_16507);
nor U23445 (N_23445,N_16914,N_16749);
nand U23446 (N_23446,N_19072,N_18284);
nor U23447 (N_23447,N_15421,N_18121);
and U23448 (N_23448,N_19682,N_19486);
or U23449 (N_23449,N_16056,N_18525);
nand U23450 (N_23450,N_18485,N_18347);
or U23451 (N_23451,N_18310,N_16451);
nand U23452 (N_23452,N_17439,N_17097);
and U23453 (N_23453,N_18268,N_15563);
nand U23454 (N_23454,N_17385,N_17360);
or U23455 (N_23455,N_17297,N_17543);
nor U23456 (N_23456,N_16087,N_16193);
and U23457 (N_23457,N_18799,N_19881);
and U23458 (N_23458,N_18077,N_17732);
xor U23459 (N_23459,N_15314,N_17002);
or U23460 (N_23460,N_17897,N_18446);
or U23461 (N_23461,N_16742,N_17108);
nor U23462 (N_23462,N_17286,N_18470);
nor U23463 (N_23463,N_15501,N_16958);
or U23464 (N_23464,N_16801,N_18408);
or U23465 (N_23465,N_16753,N_15128);
or U23466 (N_23466,N_19661,N_19471);
nor U23467 (N_23467,N_15292,N_16264);
and U23468 (N_23468,N_17983,N_19474);
and U23469 (N_23469,N_15078,N_15115);
and U23470 (N_23470,N_15014,N_19738);
or U23471 (N_23471,N_19153,N_19268);
nand U23472 (N_23472,N_19171,N_18382);
or U23473 (N_23473,N_18817,N_16760);
nor U23474 (N_23474,N_19211,N_15634);
or U23475 (N_23475,N_18310,N_18377);
nor U23476 (N_23476,N_15288,N_15147);
or U23477 (N_23477,N_16139,N_15293);
nor U23478 (N_23478,N_16472,N_17439);
nand U23479 (N_23479,N_16752,N_17410);
nand U23480 (N_23480,N_17069,N_19358);
nand U23481 (N_23481,N_19174,N_17594);
nor U23482 (N_23482,N_17284,N_15454);
nor U23483 (N_23483,N_15994,N_15692);
and U23484 (N_23484,N_15417,N_15963);
or U23485 (N_23485,N_18251,N_17202);
nor U23486 (N_23486,N_17817,N_18316);
and U23487 (N_23487,N_19533,N_15982);
or U23488 (N_23488,N_19451,N_18913);
nor U23489 (N_23489,N_16627,N_17591);
or U23490 (N_23490,N_15454,N_19007);
and U23491 (N_23491,N_16421,N_16872);
or U23492 (N_23492,N_15907,N_15563);
or U23493 (N_23493,N_19225,N_15082);
and U23494 (N_23494,N_19374,N_15340);
and U23495 (N_23495,N_17778,N_17166);
and U23496 (N_23496,N_18512,N_19404);
or U23497 (N_23497,N_19037,N_15577);
nand U23498 (N_23498,N_19345,N_18705);
and U23499 (N_23499,N_17127,N_17760);
nor U23500 (N_23500,N_19874,N_16398);
or U23501 (N_23501,N_15859,N_16474);
or U23502 (N_23502,N_18075,N_16087);
and U23503 (N_23503,N_15721,N_16594);
and U23504 (N_23504,N_17232,N_17493);
nand U23505 (N_23505,N_18661,N_19589);
nor U23506 (N_23506,N_15814,N_15784);
or U23507 (N_23507,N_18500,N_18424);
nor U23508 (N_23508,N_15463,N_18046);
xor U23509 (N_23509,N_15931,N_18413);
or U23510 (N_23510,N_15392,N_19849);
nor U23511 (N_23511,N_18154,N_19603);
nor U23512 (N_23512,N_19031,N_17999);
or U23513 (N_23513,N_16781,N_19043);
nand U23514 (N_23514,N_16802,N_15120);
and U23515 (N_23515,N_19047,N_16762);
nand U23516 (N_23516,N_15688,N_16047);
nor U23517 (N_23517,N_16734,N_19394);
nand U23518 (N_23518,N_17201,N_15740);
nor U23519 (N_23519,N_18937,N_19086);
xor U23520 (N_23520,N_15544,N_18496);
nand U23521 (N_23521,N_15353,N_19649);
nor U23522 (N_23522,N_15375,N_18457);
nor U23523 (N_23523,N_18341,N_16996);
and U23524 (N_23524,N_17467,N_15313);
or U23525 (N_23525,N_19183,N_18794);
nand U23526 (N_23526,N_17503,N_15533);
or U23527 (N_23527,N_16837,N_16527);
or U23528 (N_23528,N_16201,N_18244);
nand U23529 (N_23529,N_19019,N_18983);
and U23530 (N_23530,N_16808,N_15470);
or U23531 (N_23531,N_16142,N_18124);
and U23532 (N_23532,N_16208,N_16235);
or U23533 (N_23533,N_15075,N_16197);
and U23534 (N_23534,N_18947,N_18418);
nand U23535 (N_23535,N_15594,N_19650);
nand U23536 (N_23536,N_18280,N_19248);
nor U23537 (N_23537,N_17409,N_16015);
nor U23538 (N_23538,N_17869,N_18929);
nand U23539 (N_23539,N_16079,N_18384);
nand U23540 (N_23540,N_17815,N_18666);
and U23541 (N_23541,N_18939,N_18413);
nand U23542 (N_23542,N_16500,N_19684);
or U23543 (N_23543,N_15569,N_16834);
and U23544 (N_23544,N_17480,N_19116);
and U23545 (N_23545,N_15550,N_16137);
nor U23546 (N_23546,N_18845,N_15094);
nor U23547 (N_23547,N_17520,N_18507);
nor U23548 (N_23548,N_18163,N_18213);
nor U23549 (N_23549,N_17427,N_17289);
nor U23550 (N_23550,N_19688,N_15076);
or U23551 (N_23551,N_18217,N_15642);
nand U23552 (N_23552,N_15623,N_16344);
nand U23553 (N_23553,N_16823,N_15689);
or U23554 (N_23554,N_15695,N_17885);
and U23555 (N_23555,N_18611,N_19017);
or U23556 (N_23556,N_16995,N_17726);
and U23557 (N_23557,N_19313,N_17984);
nand U23558 (N_23558,N_19389,N_17019);
nor U23559 (N_23559,N_16110,N_19167);
and U23560 (N_23560,N_15324,N_16400);
nor U23561 (N_23561,N_17495,N_15149);
nand U23562 (N_23562,N_18788,N_18330);
nand U23563 (N_23563,N_19807,N_18514);
nand U23564 (N_23564,N_18227,N_16975);
and U23565 (N_23565,N_19814,N_15743);
or U23566 (N_23566,N_18697,N_15515);
or U23567 (N_23567,N_19413,N_16300);
nand U23568 (N_23568,N_18700,N_16396);
nor U23569 (N_23569,N_19240,N_18024);
nand U23570 (N_23570,N_18138,N_19618);
and U23571 (N_23571,N_16200,N_15447);
nor U23572 (N_23572,N_15686,N_16829);
nor U23573 (N_23573,N_19502,N_19838);
or U23574 (N_23574,N_17263,N_18735);
nand U23575 (N_23575,N_16974,N_16309);
nand U23576 (N_23576,N_16732,N_15446);
nor U23577 (N_23577,N_15203,N_17053);
or U23578 (N_23578,N_16241,N_15524);
or U23579 (N_23579,N_16771,N_18615);
nor U23580 (N_23580,N_17091,N_16279);
nand U23581 (N_23581,N_16205,N_17045);
and U23582 (N_23582,N_15839,N_15251);
or U23583 (N_23583,N_18478,N_15965);
and U23584 (N_23584,N_18795,N_18643);
and U23585 (N_23585,N_17187,N_18572);
or U23586 (N_23586,N_15781,N_19779);
and U23587 (N_23587,N_19030,N_18238);
and U23588 (N_23588,N_16825,N_16219);
nand U23589 (N_23589,N_18450,N_17390);
or U23590 (N_23590,N_15451,N_19950);
nor U23591 (N_23591,N_17908,N_18276);
and U23592 (N_23592,N_16832,N_16770);
nor U23593 (N_23593,N_16571,N_17926);
or U23594 (N_23594,N_15844,N_17966);
nand U23595 (N_23595,N_18174,N_19661);
and U23596 (N_23596,N_15872,N_15952);
xnor U23597 (N_23597,N_18183,N_15389);
nor U23598 (N_23598,N_16927,N_15388);
and U23599 (N_23599,N_18948,N_19356);
or U23600 (N_23600,N_19054,N_16949);
or U23601 (N_23601,N_18185,N_17892);
nand U23602 (N_23602,N_18622,N_16170);
nand U23603 (N_23603,N_16703,N_16675);
nor U23604 (N_23604,N_19130,N_16961);
or U23605 (N_23605,N_18493,N_16957);
and U23606 (N_23606,N_19662,N_16201);
nand U23607 (N_23607,N_19297,N_17718);
nand U23608 (N_23608,N_16072,N_15377);
nor U23609 (N_23609,N_18465,N_18955);
or U23610 (N_23610,N_18814,N_17826);
nor U23611 (N_23611,N_17723,N_19623);
or U23612 (N_23612,N_17920,N_18995);
and U23613 (N_23613,N_18016,N_16446);
and U23614 (N_23614,N_17127,N_19120);
nor U23615 (N_23615,N_19406,N_15521);
nor U23616 (N_23616,N_18661,N_15911);
and U23617 (N_23617,N_18272,N_18682);
or U23618 (N_23618,N_17108,N_18351);
and U23619 (N_23619,N_17073,N_19851);
nor U23620 (N_23620,N_16025,N_19136);
or U23621 (N_23621,N_17891,N_19744);
nor U23622 (N_23622,N_15887,N_18645);
or U23623 (N_23623,N_19778,N_18494);
and U23624 (N_23624,N_18175,N_17369);
nand U23625 (N_23625,N_19528,N_19380);
nor U23626 (N_23626,N_17818,N_15099);
nand U23627 (N_23627,N_16069,N_16494);
and U23628 (N_23628,N_19188,N_16336);
nand U23629 (N_23629,N_19229,N_19360);
or U23630 (N_23630,N_16235,N_18499);
and U23631 (N_23631,N_16149,N_17443);
xor U23632 (N_23632,N_18481,N_16164);
or U23633 (N_23633,N_18021,N_16679);
nand U23634 (N_23634,N_19949,N_18726);
and U23635 (N_23635,N_19716,N_17779);
nor U23636 (N_23636,N_16610,N_19644);
and U23637 (N_23637,N_17605,N_17166);
xor U23638 (N_23638,N_15819,N_19199);
nor U23639 (N_23639,N_18637,N_18295);
or U23640 (N_23640,N_18967,N_17931);
and U23641 (N_23641,N_17173,N_17899);
nand U23642 (N_23642,N_16709,N_16795);
and U23643 (N_23643,N_19355,N_15794);
nand U23644 (N_23644,N_16802,N_15197);
or U23645 (N_23645,N_17189,N_17692);
nor U23646 (N_23646,N_15045,N_18627);
xor U23647 (N_23647,N_15803,N_16599);
and U23648 (N_23648,N_18178,N_17002);
nor U23649 (N_23649,N_16368,N_19440);
xor U23650 (N_23650,N_16910,N_18347);
or U23651 (N_23651,N_16968,N_18579);
and U23652 (N_23652,N_17258,N_15465);
nor U23653 (N_23653,N_16467,N_18828);
nand U23654 (N_23654,N_19332,N_19121);
and U23655 (N_23655,N_18112,N_15326);
nor U23656 (N_23656,N_17624,N_16353);
and U23657 (N_23657,N_19545,N_19831);
nor U23658 (N_23658,N_18180,N_17609);
nand U23659 (N_23659,N_18052,N_17676);
and U23660 (N_23660,N_16552,N_16219);
nand U23661 (N_23661,N_16646,N_17761);
nand U23662 (N_23662,N_18837,N_17264);
or U23663 (N_23663,N_17611,N_15767);
or U23664 (N_23664,N_18102,N_17608);
or U23665 (N_23665,N_17015,N_16496);
or U23666 (N_23666,N_16989,N_17741);
nor U23667 (N_23667,N_18327,N_18539);
or U23668 (N_23668,N_17197,N_16773);
nor U23669 (N_23669,N_18852,N_17593);
nand U23670 (N_23670,N_18904,N_15757);
and U23671 (N_23671,N_15708,N_16053);
nand U23672 (N_23672,N_15122,N_15154);
nand U23673 (N_23673,N_17836,N_18009);
nor U23674 (N_23674,N_18243,N_17404);
or U23675 (N_23675,N_15998,N_16811);
or U23676 (N_23676,N_19229,N_18933);
or U23677 (N_23677,N_18422,N_16514);
or U23678 (N_23678,N_15633,N_17243);
nor U23679 (N_23679,N_18097,N_19398);
or U23680 (N_23680,N_18429,N_16000);
nand U23681 (N_23681,N_19271,N_16359);
or U23682 (N_23682,N_19058,N_17507);
or U23683 (N_23683,N_16878,N_19236);
nor U23684 (N_23684,N_19503,N_16612);
nand U23685 (N_23685,N_16839,N_17916);
or U23686 (N_23686,N_15610,N_15541);
nand U23687 (N_23687,N_18710,N_16607);
nor U23688 (N_23688,N_18941,N_16604);
nand U23689 (N_23689,N_18911,N_19572);
nor U23690 (N_23690,N_19734,N_15048);
or U23691 (N_23691,N_19859,N_17279);
and U23692 (N_23692,N_19065,N_16892);
or U23693 (N_23693,N_18814,N_17141);
or U23694 (N_23694,N_18918,N_16752);
nor U23695 (N_23695,N_16045,N_16290);
xnor U23696 (N_23696,N_15774,N_15649);
or U23697 (N_23697,N_16390,N_17925);
nand U23698 (N_23698,N_15578,N_19191);
and U23699 (N_23699,N_18138,N_18910);
and U23700 (N_23700,N_19204,N_18336);
or U23701 (N_23701,N_17547,N_17661);
and U23702 (N_23702,N_17645,N_16765);
and U23703 (N_23703,N_18350,N_15433);
nand U23704 (N_23704,N_18937,N_19727);
and U23705 (N_23705,N_16122,N_19251);
nand U23706 (N_23706,N_19230,N_16142);
nand U23707 (N_23707,N_17444,N_18298);
nor U23708 (N_23708,N_19486,N_18520);
or U23709 (N_23709,N_17989,N_16167);
xor U23710 (N_23710,N_19107,N_18124);
nand U23711 (N_23711,N_17403,N_15382);
nor U23712 (N_23712,N_16823,N_15797);
nor U23713 (N_23713,N_15154,N_19473);
nand U23714 (N_23714,N_19692,N_15024);
or U23715 (N_23715,N_17120,N_15276);
and U23716 (N_23716,N_17970,N_19209);
nor U23717 (N_23717,N_17870,N_16895);
nand U23718 (N_23718,N_15058,N_18388);
nor U23719 (N_23719,N_16403,N_17547);
or U23720 (N_23720,N_18697,N_19329);
nor U23721 (N_23721,N_16710,N_17466);
nor U23722 (N_23722,N_17619,N_18654);
or U23723 (N_23723,N_19279,N_19131);
nand U23724 (N_23724,N_18375,N_15479);
xnor U23725 (N_23725,N_19918,N_15088);
nor U23726 (N_23726,N_15548,N_15206);
or U23727 (N_23727,N_18654,N_19703);
or U23728 (N_23728,N_17526,N_18920);
nand U23729 (N_23729,N_18118,N_16996);
nor U23730 (N_23730,N_18338,N_18111);
nand U23731 (N_23731,N_15283,N_17540);
nand U23732 (N_23732,N_15607,N_15966);
or U23733 (N_23733,N_16298,N_15377);
or U23734 (N_23734,N_18774,N_17323);
and U23735 (N_23735,N_15890,N_16060);
and U23736 (N_23736,N_18585,N_19019);
or U23737 (N_23737,N_17188,N_18963);
and U23738 (N_23738,N_17151,N_15086);
and U23739 (N_23739,N_17803,N_17717);
nor U23740 (N_23740,N_17434,N_16703);
nor U23741 (N_23741,N_16921,N_18636);
or U23742 (N_23742,N_19821,N_16778);
nor U23743 (N_23743,N_18898,N_19266);
and U23744 (N_23744,N_19882,N_15993);
xnor U23745 (N_23745,N_18573,N_19310);
and U23746 (N_23746,N_15536,N_15260);
nand U23747 (N_23747,N_18379,N_19335);
nor U23748 (N_23748,N_15575,N_19350);
nand U23749 (N_23749,N_15251,N_17428);
and U23750 (N_23750,N_17315,N_18762);
nor U23751 (N_23751,N_18495,N_16453);
nand U23752 (N_23752,N_17832,N_15048);
and U23753 (N_23753,N_16434,N_17343);
or U23754 (N_23754,N_16981,N_17673);
nand U23755 (N_23755,N_19194,N_15999);
nor U23756 (N_23756,N_17159,N_17350);
or U23757 (N_23757,N_15162,N_19238);
and U23758 (N_23758,N_15280,N_17853);
nand U23759 (N_23759,N_17750,N_17580);
xnor U23760 (N_23760,N_17203,N_19893);
nor U23761 (N_23761,N_18973,N_17586);
nand U23762 (N_23762,N_16423,N_19459);
and U23763 (N_23763,N_18563,N_15548);
and U23764 (N_23764,N_17987,N_19878);
nand U23765 (N_23765,N_19617,N_18569);
nor U23766 (N_23766,N_16299,N_18322);
or U23767 (N_23767,N_17413,N_15554);
nand U23768 (N_23768,N_15571,N_15614);
nand U23769 (N_23769,N_15130,N_15849);
nand U23770 (N_23770,N_18088,N_19456);
nand U23771 (N_23771,N_19019,N_15877);
xnor U23772 (N_23772,N_16373,N_15493);
and U23773 (N_23773,N_15187,N_18778);
or U23774 (N_23774,N_17402,N_15633);
nand U23775 (N_23775,N_15887,N_19129);
or U23776 (N_23776,N_18852,N_16528);
nand U23777 (N_23777,N_18629,N_19050);
or U23778 (N_23778,N_19782,N_17532);
nor U23779 (N_23779,N_19407,N_15305);
and U23780 (N_23780,N_18028,N_15489);
xor U23781 (N_23781,N_17844,N_17674);
or U23782 (N_23782,N_19765,N_16101);
or U23783 (N_23783,N_18472,N_16657);
and U23784 (N_23784,N_18815,N_16493);
nand U23785 (N_23785,N_15598,N_17846);
and U23786 (N_23786,N_17346,N_18894);
or U23787 (N_23787,N_19081,N_19646);
nand U23788 (N_23788,N_15580,N_19167);
and U23789 (N_23789,N_17933,N_16991);
and U23790 (N_23790,N_15051,N_15822);
or U23791 (N_23791,N_17423,N_16777);
and U23792 (N_23792,N_16774,N_17834);
nor U23793 (N_23793,N_16044,N_18149);
or U23794 (N_23794,N_17759,N_17493);
or U23795 (N_23795,N_19294,N_16116);
nand U23796 (N_23796,N_15465,N_19007);
and U23797 (N_23797,N_17322,N_17116);
nor U23798 (N_23798,N_19903,N_17482);
nor U23799 (N_23799,N_19599,N_15382);
nand U23800 (N_23800,N_15881,N_19290);
nor U23801 (N_23801,N_16849,N_15697);
or U23802 (N_23802,N_17752,N_15801);
nor U23803 (N_23803,N_18304,N_19355);
nand U23804 (N_23804,N_18793,N_19046);
or U23805 (N_23805,N_16066,N_15723);
nand U23806 (N_23806,N_15327,N_18368);
nand U23807 (N_23807,N_15019,N_16548);
and U23808 (N_23808,N_16574,N_15844);
and U23809 (N_23809,N_15230,N_15914);
and U23810 (N_23810,N_19733,N_16776);
or U23811 (N_23811,N_17076,N_15455);
and U23812 (N_23812,N_15700,N_19159);
nand U23813 (N_23813,N_16710,N_18068);
nand U23814 (N_23814,N_16614,N_15738);
nand U23815 (N_23815,N_17613,N_19760);
nor U23816 (N_23816,N_19082,N_18177);
nor U23817 (N_23817,N_16728,N_16727);
or U23818 (N_23818,N_16243,N_18079);
nor U23819 (N_23819,N_18616,N_19680);
xnor U23820 (N_23820,N_19326,N_15351);
or U23821 (N_23821,N_19264,N_15284);
nor U23822 (N_23822,N_17193,N_15971);
nor U23823 (N_23823,N_18789,N_19356);
and U23824 (N_23824,N_17179,N_17499);
nor U23825 (N_23825,N_15077,N_15358);
and U23826 (N_23826,N_18049,N_16249);
nand U23827 (N_23827,N_18777,N_18214);
nand U23828 (N_23828,N_15577,N_16567);
or U23829 (N_23829,N_17849,N_17090);
nor U23830 (N_23830,N_18602,N_19300);
and U23831 (N_23831,N_18988,N_18626);
or U23832 (N_23832,N_19116,N_18879);
nor U23833 (N_23833,N_15159,N_15232);
nand U23834 (N_23834,N_17992,N_15218);
nand U23835 (N_23835,N_15523,N_19625);
nand U23836 (N_23836,N_19997,N_16757);
nor U23837 (N_23837,N_17975,N_16367);
or U23838 (N_23838,N_17487,N_18375);
and U23839 (N_23839,N_16439,N_19425);
nor U23840 (N_23840,N_16146,N_19242);
or U23841 (N_23841,N_17501,N_16812);
nor U23842 (N_23842,N_15528,N_16923);
nor U23843 (N_23843,N_18961,N_19431);
or U23844 (N_23844,N_19784,N_18999);
nand U23845 (N_23845,N_17999,N_15597);
and U23846 (N_23846,N_17696,N_18433);
nand U23847 (N_23847,N_15167,N_15983);
or U23848 (N_23848,N_19033,N_18752);
or U23849 (N_23849,N_17359,N_16223);
nor U23850 (N_23850,N_17090,N_19479);
or U23851 (N_23851,N_16720,N_16627);
nand U23852 (N_23852,N_19014,N_16923);
nor U23853 (N_23853,N_15295,N_17582);
nand U23854 (N_23854,N_18770,N_17804);
nand U23855 (N_23855,N_15281,N_19829);
or U23856 (N_23856,N_17081,N_19427);
nand U23857 (N_23857,N_19150,N_19708);
nor U23858 (N_23858,N_19089,N_16155);
nor U23859 (N_23859,N_17463,N_16288);
nand U23860 (N_23860,N_16647,N_17222);
nand U23861 (N_23861,N_19789,N_15283);
nor U23862 (N_23862,N_15875,N_17239);
or U23863 (N_23863,N_18677,N_17024);
or U23864 (N_23864,N_15256,N_19444);
nor U23865 (N_23865,N_17513,N_15223);
and U23866 (N_23866,N_16743,N_15020);
nor U23867 (N_23867,N_17039,N_17711);
nor U23868 (N_23868,N_18012,N_16482);
and U23869 (N_23869,N_15264,N_15246);
or U23870 (N_23870,N_19440,N_15997);
nand U23871 (N_23871,N_17196,N_15520);
nor U23872 (N_23872,N_17245,N_15505);
nor U23873 (N_23873,N_15989,N_15808);
nand U23874 (N_23874,N_15972,N_16415);
nand U23875 (N_23875,N_19568,N_15790);
nor U23876 (N_23876,N_16230,N_18114);
and U23877 (N_23877,N_19670,N_16772);
xor U23878 (N_23878,N_19113,N_18103);
nand U23879 (N_23879,N_15247,N_19590);
and U23880 (N_23880,N_15306,N_17019);
and U23881 (N_23881,N_18805,N_16171);
nor U23882 (N_23882,N_18069,N_16237);
or U23883 (N_23883,N_17111,N_17174);
and U23884 (N_23884,N_19938,N_18442);
nor U23885 (N_23885,N_16152,N_18470);
or U23886 (N_23886,N_18727,N_16722);
and U23887 (N_23887,N_17562,N_18588);
or U23888 (N_23888,N_18857,N_19490);
or U23889 (N_23889,N_15161,N_18805);
or U23890 (N_23890,N_16585,N_16614);
nand U23891 (N_23891,N_15419,N_16329);
nor U23892 (N_23892,N_16391,N_19471);
and U23893 (N_23893,N_19638,N_16479);
and U23894 (N_23894,N_15416,N_19987);
nor U23895 (N_23895,N_18343,N_19201);
nand U23896 (N_23896,N_16716,N_17931);
or U23897 (N_23897,N_18608,N_18929);
nand U23898 (N_23898,N_17672,N_17552);
or U23899 (N_23899,N_16297,N_19159);
and U23900 (N_23900,N_18284,N_17607);
and U23901 (N_23901,N_17571,N_17840);
and U23902 (N_23902,N_17287,N_15090);
or U23903 (N_23903,N_16854,N_16335);
nand U23904 (N_23904,N_15318,N_19881);
nand U23905 (N_23905,N_19257,N_17758);
nand U23906 (N_23906,N_19695,N_18685);
nand U23907 (N_23907,N_16702,N_17685);
or U23908 (N_23908,N_17997,N_17251);
nand U23909 (N_23909,N_18977,N_18213);
nor U23910 (N_23910,N_17945,N_16874);
nor U23911 (N_23911,N_17972,N_17725);
and U23912 (N_23912,N_19288,N_16143);
nor U23913 (N_23913,N_15439,N_17163);
and U23914 (N_23914,N_19569,N_16600);
or U23915 (N_23915,N_18296,N_17532);
or U23916 (N_23916,N_15122,N_19334);
nand U23917 (N_23917,N_19247,N_19795);
or U23918 (N_23918,N_16239,N_18531);
or U23919 (N_23919,N_15704,N_19915);
and U23920 (N_23920,N_16539,N_19254);
nor U23921 (N_23921,N_18769,N_19750);
nand U23922 (N_23922,N_17640,N_18168);
nor U23923 (N_23923,N_19796,N_15906);
or U23924 (N_23924,N_16936,N_19139);
or U23925 (N_23925,N_16211,N_15592);
or U23926 (N_23926,N_17756,N_16863);
nor U23927 (N_23927,N_15610,N_16513);
or U23928 (N_23928,N_16800,N_19177);
and U23929 (N_23929,N_19339,N_17134);
or U23930 (N_23930,N_15369,N_16309);
and U23931 (N_23931,N_16542,N_15749);
or U23932 (N_23932,N_15341,N_19193);
nor U23933 (N_23933,N_18621,N_17967);
or U23934 (N_23934,N_17540,N_15910);
nor U23935 (N_23935,N_17593,N_16008);
nand U23936 (N_23936,N_16431,N_19196);
nor U23937 (N_23937,N_19816,N_18387);
and U23938 (N_23938,N_19390,N_19412);
and U23939 (N_23939,N_15484,N_15652);
nand U23940 (N_23940,N_18358,N_16329);
and U23941 (N_23941,N_19802,N_19410);
nor U23942 (N_23942,N_17281,N_19483);
or U23943 (N_23943,N_16115,N_18797);
nand U23944 (N_23944,N_18130,N_16875);
or U23945 (N_23945,N_15939,N_16165);
and U23946 (N_23946,N_19924,N_15952);
and U23947 (N_23947,N_16610,N_16067);
nand U23948 (N_23948,N_17397,N_18058);
nand U23949 (N_23949,N_15631,N_17798);
nor U23950 (N_23950,N_16399,N_17826);
nor U23951 (N_23951,N_19263,N_16941);
and U23952 (N_23952,N_16939,N_16615);
and U23953 (N_23953,N_16569,N_18243);
and U23954 (N_23954,N_19049,N_15371);
and U23955 (N_23955,N_15047,N_15255);
or U23956 (N_23956,N_19038,N_15351);
nand U23957 (N_23957,N_17642,N_15368);
or U23958 (N_23958,N_17515,N_19883);
nor U23959 (N_23959,N_19650,N_15663);
nand U23960 (N_23960,N_16689,N_16045);
and U23961 (N_23961,N_17463,N_15122);
and U23962 (N_23962,N_18894,N_19941);
or U23963 (N_23963,N_19177,N_18826);
and U23964 (N_23964,N_15789,N_17486);
nor U23965 (N_23965,N_15186,N_17181);
nand U23966 (N_23966,N_17183,N_18084);
nor U23967 (N_23967,N_18015,N_19230);
nor U23968 (N_23968,N_17578,N_17210);
nor U23969 (N_23969,N_18258,N_16514);
nand U23970 (N_23970,N_18896,N_17269);
nand U23971 (N_23971,N_18943,N_15736);
or U23972 (N_23972,N_18758,N_18448);
or U23973 (N_23973,N_17243,N_15161);
or U23974 (N_23974,N_17793,N_19212);
nand U23975 (N_23975,N_18344,N_18006);
and U23976 (N_23976,N_16549,N_17266);
and U23977 (N_23977,N_17828,N_15429);
and U23978 (N_23978,N_17156,N_16637);
and U23979 (N_23979,N_16534,N_17841);
nand U23980 (N_23980,N_18002,N_17625);
and U23981 (N_23981,N_19318,N_16923);
and U23982 (N_23982,N_18122,N_19291);
nor U23983 (N_23983,N_17325,N_15710);
and U23984 (N_23984,N_18021,N_17882);
nand U23985 (N_23985,N_15498,N_15367);
nand U23986 (N_23986,N_17447,N_19408);
and U23987 (N_23987,N_16785,N_15347);
nor U23988 (N_23988,N_15848,N_19246);
xor U23989 (N_23989,N_17237,N_16206);
or U23990 (N_23990,N_16434,N_17732);
nor U23991 (N_23991,N_15475,N_17430);
nand U23992 (N_23992,N_18746,N_17321);
nor U23993 (N_23993,N_15741,N_19492);
or U23994 (N_23994,N_17305,N_15594);
and U23995 (N_23995,N_16672,N_18002);
and U23996 (N_23996,N_16906,N_17069);
nor U23997 (N_23997,N_16614,N_16183);
and U23998 (N_23998,N_16808,N_17129);
xnor U23999 (N_23999,N_17007,N_17743);
and U24000 (N_24000,N_15382,N_17240);
and U24001 (N_24001,N_17150,N_16453);
and U24002 (N_24002,N_18264,N_15032);
or U24003 (N_24003,N_19867,N_17648);
and U24004 (N_24004,N_17973,N_15243);
and U24005 (N_24005,N_19950,N_15339);
xnor U24006 (N_24006,N_17294,N_15723);
and U24007 (N_24007,N_17549,N_17863);
nand U24008 (N_24008,N_18393,N_19728);
nor U24009 (N_24009,N_18717,N_15900);
and U24010 (N_24010,N_16484,N_16556);
or U24011 (N_24011,N_15141,N_19028);
and U24012 (N_24012,N_15750,N_17572);
and U24013 (N_24013,N_17298,N_18735);
nand U24014 (N_24014,N_17787,N_17269);
and U24015 (N_24015,N_15127,N_19524);
and U24016 (N_24016,N_19682,N_16337);
and U24017 (N_24017,N_18612,N_16815);
nor U24018 (N_24018,N_15794,N_16684);
or U24019 (N_24019,N_19388,N_19612);
and U24020 (N_24020,N_15678,N_19510);
nand U24021 (N_24021,N_18226,N_17021);
nor U24022 (N_24022,N_17295,N_15657);
or U24023 (N_24023,N_19979,N_18756);
nor U24024 (N_24024,N_19149,N_19280);
nor U24025 (N_24025,N_18696,N_19954);
nor U24026 (N_24026,N_19561,N_15098);
nand U24027 (N_24027,N_18386,N_17010);
nor U24028 (N_24028,N_15010,N_17972);
nor U24029 (N_24029,N_19169,N_18868);
or U24030 (N_24030,N_16176,N_15703);
and U24031 (N_24031,N_18371,N_18565);
xnor U24032 (N_24032,N_15242,N_18644);
or U24033 (N_24033,N_19610,N_18659);
nand U24034 (N_24034,N_16313,N_18514);
nor U24035 (N_24035,N_17976,N_16588);
nand U24036 (N_24036,N_17701,N_16373);
or U24037 (N_24037,N_16290,N_17783);
nor U24038 (N_24038,N_19667,N_19166);
nand U24039 (N_24039,N_16981,N_18438);
or U24040 (N_24040,N_19086,N_16621);
and U24041 (N_24041,N_18152,N_17689);
nand U24042 (N_24042,N_19841,N_16188);
or U24043 (N_24043,N_15237,N_19929);
or U24044 (N_24044,N_16705,N_17217);
or U24045 (N_24045,N_19237,N_15217);
nand U24046 (N_24046,N_17954,N_18248);
and U24047 (N_24047,N_19053,N_18434);
and U24048 (N_24048,N_17771,N_18832);
or U24049 (N_24049,N_16736,N_15141);
and U24050 (N_24050,N_17465,N_18818);
nand U24051 (N_24051,N_16825,N_15546);
or U24052 (N_24052,N_18080,N_19847);
and U24053 (N_24053,N_17577,N_16514);
xor U24054 (N_24054,N_19618,N_18023);
nor U24055 (N_24055,N_15379,N_17568);
nand U24056 (N_24056,N_19930,N_15608);
and U24057 (N_24057,N_17765,N_16904);
or U24058 (N_24058,N_19777,N_19318);
xnor U24059 (N_24059,N_18943,N_17775);
nand U24060 (N_24060,N_17567,N_16522);
xnor U24061 (N_24061,N_18265,N_15108);
or U24062 (N_24062,N_17517,N_16200);
nor U24063 (N_24063,N_18866,N_18182);
nand U24064 (N_24064,N_15680,N_18148);
and U24065 (N_24065,N_19452,N_15370);
nor U24066 (N_24066,N_16516,N_18766);
nand U24067 (N_24067,N_16398,N_19226);
or U24068 (N_24068,N_18015,N_19524);
and U24069 (N_24069,N_18314,N_18155);
or U24070 (N_24070,N_16331,N_17297);
or U24071 (N_24071,N_18229,N_19280);
or U24072 (N_24072,N_19647,N_17524);
nor U24073 (N_24073,N_19190,N_15272);
or U24074 (N_24074,N_18234,N_17890);
nor U24075 (N_24075,N_15849,N_19002);
and U24076 (N_24076,N_19655,N_18534);
nor U24077 (N_24077,N_18426,N_18851);
or U24078 (N_24078,N_19021,N_19993);
or U24079 (N_24079,N_17449,N_19013);
and U24080 (N_24080,N_15205,N_19454);
and U24081 (N_24081,N_18558,N_17556);
nand U24082 (N_24082,N_19819,N_18226);
nor U24083 (N_24083,N_16606,N_15450);
and U24084 (N_24084,N_15025,N_16785);
or U24085 (N_24085,N_19176,N_16868);
nand U24086 (N_24086,N_15067,N_15251);
and U24087 (N_24087,N_18180,N_16490);
nor U24088 (N_24088,N_18495,N_18530);
nand U24089 (N_24089,N_15713,N_17022);
nor U24090 (N_24090,N_19573,N_15200);
xor U24091 (N_24091,N_15284,N_17579);
nand U24092 (N_24092,N_16421,N_19991);
nand U24093 (N_24093,N_16316,N_17879);
nand U24094 (N_24094,N_17915,N_18286);
and U24095 (N_24095,N_17664,N_17162);
or U24096 (N_24096,N_15290,N_19032);
or U24097 (N_24097,N_18763,N_16056);
and U24098 (N_24098,N_16782,N_16812);
nor U24099 (N_24099,N_19055,N_19012);
nand U24100 (N_24100,N_16669,N_18798);
nand U24101 (N_24101,N_19924,N_18666);
or U24102 (N_24102,N_18733,N_19913);
and U24103 (N_24103,N_18049,N_19356);
or U24104 (N_24104,N_17299,N_19764);
nor U24105 (N_24105,N_16738,N_19877);
nand U24106 (N_24106,N_15029,N_15748);
or U24107 (N_24107,N_15276,N_16086);
nor U24108 (N_24108,N_19128,N_15726);
and U24109 (N_24109,N_16135,N_15096);
and U24110 (N_24110,N_17076,N_15153);
nand U24111 (N_24111,N_18208,N_18498);
nor U24112 (N_24112,N_17147,N_16735);
nor U24113 (N_24113,N_15264,N_19295);
or U24114 (N_24114,N_18567,N_16017);
nor U24115 (N_24115,N_19277,N_16640);
nand U24116 (N_24116,N_17889,N_15588);
nand U24117 (N_24117,N_15902,N_16093);
and U24118 (N_24118,N_17108,N_16679);
or U24119 (N_24119,N_17040,N_19755);
xor U24120 (N_24120,N_17270,N_15740);
nand U24121 (N_24121,N_17182,N_17885);
xor U24122 (N_24122,N_19868,N_19386);
and U24123 (N_24123,N_19308,N_19666);
nor U24124 (N_24124,N_17342,N_17278);
nand U24125 (N_24125,N_17778,N_17069);
or U24126 (N_24126,N_19375,N_16182);
and U24127 (N_24127,N_19686,N_16321);
nand U24128 (N_24128,N_18501,N_17943);
nor U24129 (N_24129,N_15352,N_16586);
or U24130 (N_24130,N_16371,N_19741);
xnor U24131 (N_24131,N_18016,N_19133);
nand U24132 (N_24132,N_15071,N_15214);
or U24133 (N_24133,N_17788,N_16616);
or U24134 (N_24134,N_18779,N_19588);
nand U24135 (N_24135,N_17877,N_15837);
nor U24136 (N_24136,N_18987,N_19550);
nand U24137 (N_24137,N_18731,N_15557);
and U24138 (N_24138,N_17213,N_17621);
nor U24139 (N_24139,N_18612,N_16019);
nor U24140 (N_24140,N_16241,N_19716);
or U24141 (N_24141,N_15734,N_19791);
and U24142 (N_24142,N_18527,N_18793);
nand U24143 (N_24143,N_19952,N_18479);
nand U24144 (N_24144,N_16178,N_15290);
nand U24145 (N_24145,N_16838,N_15133);
and U24146 (N_24146,N_16513,N_19887);
or U24147 (N_24147,N_15869,N_16788);
nand U24148 (N_24148,N_18951,N_16403);
nand U24149 (N_24149,N_16463,N_15014);
nor U24150 (N_24150,N_16893,N_16787);
and U24151 (N_24151,N_15181,N_19499);
nor U24152 (N_24152,N_15863,N_15026);
nand U24153 (N_24153,N_18886,N_18726);
nand U24154 (N_24154,N_16681,N_17221);
nor U24155 (N_24155,N_15547,N_17493);
or U24156 (N_24156,N_15766,N_17131);
xnor U24157 (N_24157,N_16178,N_16206);
nor U24158 (N_24158,N_15828,N_15972);
or U24159 (N_24159,N_17801,N_19419);
nor U24160 (N_24160,N_15002,N_19902);
and U24161 (N_24161,N_18733,N_16542);
or U24162 (N_24162,N_18414,N_18894);
or U24163 (N_24163,N_17996,N_17667);
nor U24164 (N_24164,N_16289,N_17465);
and U24165 (N_24165,N_17865,N_19890);
and U24166 (N_24166,N_15705,N_19063);
and U24167 (N_24167,N_18669,N_15040);
nand U24168 (N_24168,N_18961,N_18065);
nand U24169 (N_24169,N_16345,N_19087);
nor U24170 (N_24170,N_18637,N_15670);
nor U24171 (N_24171,N_19271,N_18407);
and U24172 (N_24172,N_17178,N_18952);
nand U24173 (N_24173,N_18749,N_18864);
nand U24174 (N_24174,N_18644,N_15969);
or U24175 (N_24175,N_17896,N_17307);
or U24176 (N_24176,N_19597,N_15579);
nor U24177 (N_24177,N_19521,N_15047);
nor U24178 (N_24178,N_16870,N_19119);
and U24179 (N_24179,N_17336,N_18643);
and U24180 (N_24180,N_16278,N_18259);
or U24181 (N_24181,N_16172,N_19437);
and U24182 (N_24182,N_19985,N_15188);
and U24183 (N_24183,N_17710,N_19847);
nand U24184 (N_24184,N_16402,N_19654);
and U24185 (N_24185,N_17014,N_17294);
and U24186 (N_24186,N_19571,N_18479);
nand U24187 (N_24187,N_18728,N_17559);
nor U24188 (N_24188,N_15235,N_16442);
nor U24189 (N_24189,N_17339,N_16708);
and U24190 (N_24190,N_16556,N_15358);
and U24191 (N_24191,N_18482,N_16196);
nand U24192 (N_24192,N_15164,N_16539);
nor U24193 (N_24193,N_17734,N_17135);
nand U24194 (N_24194,N_17200,N_19918);
or U24195 (N_24195,N_19779,N_17101);
and U24196 (N_24196,N_15555,N_18529);
nor U24197 (N_24197,N_19562,N_18923);
nor U24198 (N_24198,N_19721,N_16546);
nand U24199 (N_24199,N_18110,N_15025);
or U24200 (N_24200,N_16497,N_15523);
nand U24201 (N_24201,N_19715,N_17461);
or U24202 (N_24202,N_15764,N_18935);
nand U24203 (N_24203,N_17056,N_17075);
or U24204 (N_24204,N_16987,N_18620);
or U24205 (N_24205,N_19488,N_17878);
or U24206 (N_24206,N_17061,N_15591);
or U24207 (N_24207,N_16664,N_16845);
or U24208 (N_24208,N_15123,N_17925);
nor U24209 (N_24209,N_15938,N_19158);
nor U24210 (N_24210,N_19620,N_18527);
and U24211 (N_24211,N_19474,N_17280);
nor U24212 (N_24212,N_15736,N_16749);
and U24213 (N_24213,N_15533,N_18688);
xor U24214 (N_24214,N_15561,N_17604);
and U24215 (N_24215,N_17155,N_16390);
nor U24216 (N_24216,N_16046,N_19069);
nand U24217 (N_24217,N_19460,N_15905);
nand U24218 (N_24218,N_17460,N_16945);
nand U24219 (N_24219,N_17590,N_16634);
or U24220 (N_24220,N_18770,N_17430);
or U24221 (N_24221,N_17828,N_18422);
nor U24222 (N_24222,N_16706,N_16078);
nor U24223 (N_24223,N_19209,N_16071);
and U24224 (N_24224,N_18661,N_17288);
nor U24225 (N_24225,N_17199,N_17999);
nor U24226 (N_24226,N_16520,N_16394);
or U24227 (N_24227,N_17011,N_15352);
nor U24228 (N_24228,N_16201,N_17531);
and U24229 (N_24229,N_15363,N_17189);
and U24230 (N_24230,N_17755,N_17248);
and U24231 (N_24231,N_16560,N_15816);
nand U24232 (N_24232,N_15345,N_18856);
or U24233 (N_24233,N_16752,N_16577);
nor U24234 (N_24234,N_15402,N_17708);
and U24235 (N_24235,N_17710,N_19486);
nand U24236 (N_24236,N_19508,N_16402);
nor U24237 (N_24237,N_18582,N_16350);
nand U24238 (N_24238,N_15993,N_15178);
or U24239 (N_24239,N_18560,N_16641);
nand U24240 (N_24240,N_16408,N_19574);
or U24241 (N_24241,N_15891,N_19911);
or U24242 (N_24242,N_16926,N_16958);
or U24243 (N_24243,N_17522,N_18025);
nor U24244 (N_24244,N_18892,N_18845);
and U24245 (N_24245,N_15643,N_16990);
nand U24246 (N_24246,N_16146,N_19071);
and U24247 (N_24247,N_15229,N_16359);
or U24248 (N_24248,N_18209,N_15954);
and U24249 (N_24249,N_19148,N_18348);
or U24250 (N_24250,N_18380,N_19641);
nand U24251 (N_24251,N_16520,N_18771);
nand U24252 (N_24252,N_17412,N_15820);
nor U24253 (N_24253,N_16837,N_19703);
nand U24254 (N_24254,N_17633,N_19080);
nor U24255 (N_24255,N_18217,N_18070);
nand U24256 (N_24256,N_19328,N_15379);
nand U24257 (N_24257,N_16334,N_19398);
or U24258 (N_24258,N_19681,N_19846);
nand U24259 (N_24259,N_19102,N_15877);
and U24260 (N_24260,N_19989,N_16008);
or U24261 (N_24261,N_15510,N_17262);
nor U24262 (N_24262,N_18089,N_16373);
nor U24263 (N_24263,N_19741,N_15698);
nand U24264 (N_24264,N_19021,N_18515);
and U24265 (N_24265,N_17779,N_17093);
nand U24266 (N_24266,N_16898,N_19122);
or U24267 (N_24267,N_17560,N_16172);
and U24268 (N_24268,N_17071,N_17032);
nor U24269 (N_24269,N_19338,N_18292);
and U24270 (N_24270,N_17403,N_19750);
nor U24271 (N_24271,N_19443,N_17776);
nand U24272 (N_24272,N_16204,N_19948);
nand U24273 (N_24273,N_19582,N_18668);
and U24274 (N_24274,N_16761,N_16627);
nand U24275 (N_24275,N_17382,N_16518);
nand U24276 (N_24276,N_15036,N_15458);
nand U24277 (N_24277,N_16939,N_18913);
nand U24278 (N_24278,N_15689,N_19393);
nor U24279 (N_24279,N_19235,N_15932);
and U24280 (N_24280,N_16915,N_15451);
nand U24281 (N_24281,N_18537,N_15315);
nand U24282 (N_24282,N_17894,N_15461);
or U24283 (N_24283,N_17761,N_18305);
nor U24284 (N_24284,N_16801,N_17368);
and U24285 (N_24285,N_16820,N_16832);
and U24286 (N_24286,N_16646,N_16492);
nor U24287 (N_24287,N_19006,N_15081);
nor U24288 (N_24288,N_19172,N_18558);
nor U24289 (N_24289,N_16893,N_17263);
nor U24290 (N_24290,N_17764,N_18513);
nand U24291 (N_24291,N_16727,N_18156);
nor U24292 (N_24292,N_15860,N_16865);
and U24293 (N_24293,N_15567,N_19637);
and U24294 (N_24294,N_19418,N_18976);
or U24295 (N_24295,N_18657,N_18270);
and U24296 (N_24296,N_16025,N_18481);
nor U24297 (N_24297,N_19922,N_15963);
and U24298 (N_24298,N_18662,N_15642);
xnor U24299 (N_24299,N_18397,N_19703);
nor U24300 (N_24300,N_19802,N_19829);
nor U24301 (N_24301,N_16566,N_18682);
nor U24302 (N_24302,N_16027,N_18081);
and U24303 (N_24303,N_16186,N_17035);
nand U24304 (N_24304,N_16830,N_19496);
nand U24305 (N_24305,N_17387,N_17590);
or U24306 (N_24306,N_16218,N_19532);
or U24307 (N_24307,N_15086,N_18096);
nand U24308 (N_24308,N_16736,N_19007);
and U24309 (N_24309,N_16610,N_15231);
nor U24310 (N_24310,N_15563,N_16724);
nor U24311 (N_24311,N_16148,N_17629);
and U24312 (N_24312,N_17939,N_18248);
or U24313 (N_24313,N_15908,N_16864);
and U24314 (N_24314,N_18905,N_18283);
and U24315 (N_24315,N_19200,N_15690);
and U24316 (N_24316,N_15203,N_19528);
nor U24317 (N_24317,N_18511,N_18311);
and U24318 (N_24318,N_17756,N_17400);
or U24319 (N_24319,N_17984,N_15701);
and U24320 (N_24320,N_18312,N_19322);
nand U24321 (N_24321,N_18706,N_16913);
nor U24322 (N_24322,N_16727,N_15541);
and U24323 (N_24323,N_16554,N_19088);
nand U24324 (N_24324,N_18911,N_17190);
or U24325 (N_24325,N_16373,N_15055);
nand U24326 (N_24326,N_17824,N_18167);
nor U24327 (N_24327,N_16893,N_19210);
and U24328 (N_24328,N_18559,N_19697);
and U24329 (N_24329,N_19804,N_19728);
xor U24330 (N_24330,N_15503,N_17548);
or U24331 (N_24331,N_15889,N_18367);
or U24332 (N_24332,N_19529,N_17700);
or U24333 (N_24333,N_19677,N_16555);
and U24334 (N_24334,N_15160,N_16784);
or U24335 (N_24335,N_16978,N_17018);
or U24336 (N_24336,N_18508,N_19682);
and U24337 (N_24337,N_16702,N_17577);
nor U24338 (N_24338,N_18480,N_19636);
and U24339 (N_24339,N_18037,N_17832);
or U24340 (N_24340,N_17028,N_15721);
nor U24341 (N_24341,N_17421,N_19262);
nor U24342 (N_24342,N_17310,N_15177);
nor U24343 (N_24343,N_16723,N_17369);
nor U24344 (N_24344,N_16801,N_17126);
nand U24345 (N_24345,N_15752,N_16865);
and U24346 (N_24346,N_17664,N_15671);
and U24347 (N_24347,N_15539,N_18672);
or U24348 (N_24348,N_15076,N_19098);
and U24349 (N_24349,N_19131,N_18918);
xnor U24350 (N_24350,N_18176,N_18406);
nor U24351 (N_24351,N_17203,N_18419);
or U24352 (N_24352,N_15164,N_19959);
nand U24353 (N_24353,N_17367,N_15681);
or U24354 (N_24354,N_17658,N_19794);
and U24355 (N_24355,N_16330,N_18385);
nand U24356 (N_24356,N_17698,N_17239);
or U24357 (N_24357,N_17924,N_19128);
or U24358 (N_24358,N_17405,N_18259);
nor U24359 (N_24359,N_18604,N_16842);
and U24360 (N_24360,N_19232,N_19851);
nand U24361 (N_24361,N_16270,N_19008);
nand U24362 (N_24362,N_15751,N_18651);
nor U24363 (N_24363,N_15280,N_18614);
and U24364 (N_24364,N_15311,N_17012);
nand U24365 (N_24365,N_18376,N_15737);
or U24366 (N_24366,N_19080,N_16168);
and U24367 (N_24367,N_15048,N_19304);
nand U24368 (N_24368,N_17559,N_17958);
and U24369 (N_24369,N_18783,N_18733);
and U24370 (N_24370,N_17229,N_15065);
and U24371 (N_24371,N_16022,N_15627);
or U24372 (N_24372,N_18537,N_17410);
and U24373 (N_24373,N_16560,N_15452);
nor U24374 (N_24374,N_18881,N_15676);
and U24375 (N_24375,N_16187,N_18930);
and U24376 (N_24376,N_19250,N_15867);
nor U24377 (N_24377,N_17591,N_15418);
nor U24378 (N_24378,N_18854,N_15000);
or U24379 (N_24379,N_18310,N_16839);
and U24380 (N_24380,N_18887,N_19230);
nand U24381 (N_24381,N_19352,N_18006);
or U24382 (N_24382,N_15846,N_18501);
nor U24383 (N_24383,N_16561,N_18638);
and U24384 (N_24384,N_16581,N_15519);
and U24385 (N_24385,N_15860,N_15132);
nor U24386 (N_24386,N_18719,N_17087);
nor U24387 (N_24387,N_19245,N_16115);
nand U24388 (N_24388,N_17549,N_19496);
nor U24389 (N_24389,N_18807,N_17188);
and U24390 (N_24390,N_15785,N_17493);
and U24391 (N_24391,N_16925,N_15873);
nand U24392 (N_24392,N_19768,N_17678);
nor U24393 (N_24393,N_19923,N_19396);
and U24394 (N_24394,N_15777,N_19009);
nor U24395 (N_24395,N_16478,N_18372);
or U24396 (N_24396,N_16053,N_17451);
nor U24397 (N_24397,N_19647,N_17714);
and U24398 (N_24398,N_16375,N_17400);
and U24399 (N_24399,N_15699,N_15741);
or U24400 (N_24400,N_17072,N_15785);
nand U24401 (N_24401,N_15468,N_18199);
or U24402 (N_24402,N_19656,N_15875);
and U24403 (N_24403,N_18538,N_15413);
nand U24404 (N_24404,N_16041,N_15026);
or U24405 (N_24405,N_18316,N_18425);
or U24406 (N_24406,N_19087,N_15025);
or U24407 (N_24407,N_15774,N_16329);
and U24408 (N_24408,N_19062,N_15995);
nor U24409 (N_24409,N_18880,N_15654);
nor U24410 (N_24410,N_19786,N_19981);
and U24411 (N_24411,N_16022,N_15179);
xor U24412 (N_24412,N_18734,N_15632);
or U24413 (N_24413,N_18567,N_18069);
or U24414 (N_24414,N_19011,N_18527);
and U24415 (N_24415,N_18345,N_15769);
nor U24416 (N_24416,N_19275,N_17012);
nor U24417 (N_24417,N_17468,N_15733);
and U24418 (N_24418,N_19222,N_17772);
nor U24419 (N_24419,N_16545,N_18255);
nand U24420 (N_24420,N_17914,N_17715);
xor U24421 (N_24421,N_17531,N_18729);
nand U24422 (N_24422,N_16605,N_19404);
or U24423 (N_24423,N_17600,N_17313);
nand U24424 (N_24424,N_15348,N_19710);
and U24425 (N_24425,N_18255,N_18615);
nand U24426 (N_24426,N_18944,N_18275);
and U24427 (N_24427,N_17402,N_19811);
or U24428 (N_24428,N_19769,N_17098);
and U24429 (N_24429,N_18774,N_15476);
and U24430 (N_24430,N_16973,N_16691);
or U24431 (N_24431,N_19173,N_18719);
and U24432 (N_24432,N_18795,N_17278);
nand U24433 (N_24433,N_19933,N_19816);
nand U24434 (N_24434,N_18406,N_19833);
and U24435 (N_24435,N_19372,N_19555);
and U24436 (N_24436,N_18282,N_17039);
and U24437 (N_24437,N_19143,N_19189);
or U24438 (N_24438,N_18299,N_15059);
and U24439 (N_24439,N_15493,N_18885);
nand U24440 (N_24440,N_15595,N_18374);
or U24441 (N_24441,N_19328,N_16274);
nor U24442 (N_24442,N_15347,N_18529);
xnor U24443 (N_24443,N_15128,N_16534);
nor U24444 (N_24444,N_17629,N_15397);
or U24445 (N_24445,N_15014,N_16483);
and U24446 (N_24446,N_17583,N_19428);
nor U24447 (N_24447,N_17942,N_19938);
nor U24448 (N_24448,N_19159,N_18379);
or U24449 (N_24449,N_15176,N_19185);
nand U24450 (N_24450,N_19248,N_16031);
nor U24451 (N_24451,N_19372,N_19947);
nor U24452 (N_24452,N_19747,N_17377);
xnor U24453 (N_24453,N_18665,N_19803);
or U24454 (N_24454,N_18426,N_15484);
nor U24455 (N_24455,N_19541,N_18773);
or U24456 (N_24456,N_18440,N_17988);
or U24457 (N_24457,N_17895,N_19768);
and U24458 (N_24458,N_16461,N_17361);
nand U24459 (N_24459,N_15696,N_15926);
nand U24460 (N_24460,N_18310,N_15261);
nor U24461 (N_24461,N_18488,N_19021);
or U24462 (N_24462,N_16727,N_18922);
or U24463 (N_24463,N_18027,N_19534);
xnor U24464 (N_24464,N_17020,N_17225);
or U24465 (N_24465,N_17233,N_19880);
nor U24466 (N_24466,N_15936,N_15945);
or U24467 (N_24467,N_18096,N_15061);
and U24468 (N_24468,N_15604,N_15109);
or U24469 (N_24469,N_19792,N_17926);
nor U24470 (N_24470,N_18879,N_18878);
nand U24471 (N_24471,N_18656,N_19120);
xor U24472 (N_24472,N_17244,N_15420);
or U24473 (N_24473,N_17113,N_17607);
and U24474 (N_24474,N_16693,N_19873);
nand U24475 (N_24475,N_19394,N_18743);
nor U24476 (N_24476,N_18313,N_17455);
nor U24477 (N_24477,N_16946,N_18190);
and U24478 (N_24478,N_17226,N_18784);
xor U24479 (N_24479,N_17169,N_16026);
nor U24480 (N_24480,N_15483,N_19892);
nor U24481 (N_24481,N_16713,N_18950);
or U24482 (N_24482,N_18729,N_17895);
and U24483 (N_24483,N_16953,N_18778);
nand U24484 (N_24484,N_18909,N_19613);
or U24485 (N_24485,N_18263,N_17104);
nand U24486 (N_24486,N_15372,N_16943);
nand U24487 (N_24487,N_18374,N_17631);
xnor U24488 (N_24488,N_19780,N_15355);
and U24489 (N_24489,N_19724,N_15440);
and U24490 (N_24490,N_19560,N_17703);
or U24491 (N_24491,N_15322,N_18339);
nor U24492 (N_24492,N_19720,N_19510);
nor U24493 (N_24493,N_17229,N_16637);
and U24494 (N_24494,N_15962,N_17707);
nand U24495 (N_24495,N_16613,N_15849);
nor U24496 (N_24496,N_16900,N_16553);
nor U24497 (N_24497,N_18295,N_19557);
nand U24498 (N_24498,N_19565,N_15435);
nand U24499 (N_24499,N_16621,N_16743);
nor U24500 (N_24500,N_19179,N_18347);
or U24501 (N_24501,N_16815,N_18119);
or U24502 (N_24502,N_16291,N_16732);
nand U24503 (N_24503,N_17814,N_19037);
and U24504 (N_24504,N_15781,N_17965);
nor U24505 (N_24505,N_15715,N_16080);
nand U24506 (N_24506,N_18419,N_15547);
or U24507 (N_24507,N_17177,N_17534);
and U24508 (N_24508,N_15266,N_16509);
nor U24509 (N_24509,N_16351,N_17342);
or U24510 (N_24510,N_17700,N_18937);
or U24511 (N_24511,N_18983,N_19144);
xor U24512 (N_24512,N_19224,N_17802);
xor U24513 (N_24513,N_18012,N_16458);
or U24514 (N_24514,N_15612,N_15548);
and U24515 (N_24515,N_15596,N_15841);
nand U24516 (N_24516,N_15390,N_15833);
nand U24517 (N_24517,N_18754,N_19564);
nor U24518 (N_24518,N_17894,N_19181);
nor U24519 (N_24519,N_15524,N_15627);
and U24520 (N_24520,N_18312,N_16729);
nand U24521 (N_24521,N_19178,N_17250);
nor U24522 (N_24522,N_18327,N_15869);
or U24523 (N_24523,N_15878,N_15776);
nand U24524 (N_24524,N_19573,N_16863);
nor U24525 (N_24525,N_16203,N_19633);
or U24526 (N_24526,N_17689,N_16703);
or U24527 (N_24527,N_19457,N_16631);
and U24528 (N_24528,N_17783,N_19837);
nand U24529 (N_24529,N_19958,N_17944);
and U24530 (N_24530,N_17097,N_16460);
nand U24531 (N_24531,N_19954,N_19114);
and U24532 (N_24532,N_18357,N_16639);
nand U24533 (N_24533,N_17994,N_15874);
or U24534 (N_24534,N_16417,N_19990);
nor U24535 (N_24535,N_16246,N_15247);
nand U24536 (N_24536,N_16151,N_15267);
nand U24537 (N_24537,N_17841,N_19199);
and U24538 (N_24538,N_18654,N_19180);
and U24539 (N_24539,N_19515,N_18103);
nand U24540 (N_24540,N_18224,N_17261);
and U24541 (N_24541,N_18215,N_18598);
and U24542 (N_24542,N_17275,N_17571);
or U24543 (N_24543,N_18848,N_18405);
nand U24544 (N_24544,N_17344,N_15505);
nand U24545 (N_24545,N_17711,N_16161);
nand U24546 (N_24546,N_16001,N_16470);
nand U24547 (N_24547,N_16572,N_19852);
nand U24548 (N_24548,N_15176,N_17604);
or U24549 (N_24549,N_17938,N_18232);
nand U24550 (N_24550,N_15701,N_16407);
nand U24551 (N_24551,N_17620,N_15956);
nor U24552 (N_24552,N_18401,N_18685);
or U24553 (N_24553,N_15962,N_19174);
and U24554 (N_24554,N_18931,N_16573);
nor U24555 (N_24555,N_16160,N_18917);
or U24556 (N_24556,N_19491,N_15897);
and U24557 (N_24557,N_16389,N_16073);
and U24558 (N_24558,N_15129,N_16729);
nor U24559 (N_24559,N_19222,N_18301);
nand U24560 (N_24560,N_16866,N_17539);
or U24561 (N_24561,N_19711,N_19809);
nand U24562 (N_24562,N_15624,N_19430);
or U24563 (N_24563,N_18860,N_17938);
nand U24564 (N_24564,N_18742,N_18257);
and U24565 (N_24565,N_19117,N_19532);
and U24566 (N_24566,N_16389,N_15217);
and U24567 (N_24567,N_18768,N_17385);
and U24568 (N_24568,N_16689,N_17535);
nand U24569 (N_24569,N_17217,N_18404);
nor U24570 (N_24570,N_19966,N_18368);
nand U24571 (N_24571,N_16263,N_19022);
nor U24572 (N_24572,N_19483,N_17243);
nor U24573 (N_24573,N_18894,N_15384);
or U24574 (N_24574,N_16195,N_19960);
or U24575 (N_24575,N_16665,N_15773);
or U24576 (N_24576,N_17471,N_16068);
and U24577 (N_24577,N_15024,N_18595);
nor U24578 (N_24578,N_15067,N_17496);
nor U24579 (N_24579,N_16700,N_15770);
and U24580 (N_24580,N_15158,N_15178);
and U24581 (N_24581,N_15267,N_17424);
nand U24582 (N_24582,N_17124,N_15814);
nand U24583 (N_24583,N_19136,N_15479);
nand U24584 (N_24584,N_16473,N_19588);
nor U24585 (N_24585,N_15012,N_18389);
and U24586 (N_24586,N_17336,N_18851);
nor U24587 (N_24587,N_19848,N_18076);
xnor U24588 (N_24588,N_19875,N_19721);
nor U24589 (N_24589,N_18304,N_18848);
and U24590 (N_24590,N_18958,N_16074);
and U24591 (N_24591,N_16578,N_15744);
and U24592 (N_24592,N_15107,N_15055);
or U24593 (N_24593,N_16194,N_15317);
or U24594 (N_24594,N_19513,N_15909);
and U24595 (N_24595,N_16904,N_18748);
or U24596 (N_24596,N_18159,N_18324);
nand U24597 (N_24597,N_16266,N_15639);
nor U24598 (N_24598,N_17224,N_15542);
nor U24599 (N_24599,N_19082,N_19936);
and U24600 (N_24600,N_19443,N_16667);
or U24601 (N_24601,N_18948,N_17181);
nor U24602 (N_24602,N_18472,N_17401);
and U24603 (N_24603,N_19942,N_19003);
and U24604 (N_24604,N_16784,N_17888);
and U24605 (N_24605,N_19916,N_19676);
and U24606 (N_24606,N_19716,N_17817);
or U24607 (N_24607,N_15538,N_16155);
nor U24608 (N_24608,N_18309,N_16759);
nand U24609 (N_24609,N_16601,N_19192);
or U24610 (N_24610,N_17319,N_18476);
and U24611 (N_24611,N_16976,N_18358);
or U24612 (N_24612,N_16160,N_17033);
or U24613 (N_24613,N_15302,N_15255);
nand U24614 (N_24614,N_18256,N_16053);
and U24615 (N_24615,N_17982,N_18623);
and U24616 (N_24616,N_15584,N_19682);
nor U24617 (N_24617,N_15596,N_16667);
nor U24618 (N_24618,N_17489,N_19266);
or U24619 (N_24619,N_17328,N_17334);
nand U24620 (N_24620,N_16523,N_15669);
or U24621 (N_24621,N_18395,N_19090);
nand U24622 (N_24622,N_16386,N_16392);
nand U24623 (N_24623,N_19059,N_17054);
nand U24624 (N_24624,N_17453,N_19725);
nand U24625 (N_24625,N_18384,N_18428);
and U24626 (N_24626,N_19489,N_15400);
nor U24627 (N_24627,N_17576,N_15868);
nor U24628 (N_24628,N_15977,N_15139);
nand U24629 (N_24629,N_16775,N_18342);
nor U24630 (N_24630,N_19276,N_16595);
nand U24631 (N_24631,N_18035,N_19586);
and U24632 (N_24632,N_19094,N_17504);
and U24633 (N_24633,N_16172,N_16045);
and U24634 (N_24634,N_16729,N_15857);
nand U24635 (N_24635,N_17858,N_18770);
nor U24636 (N_24636,N_15230,N_17687);
or U24637 (N_24637,N_18409,N_19112);
or U24638 (N_24638,N_16668,N_17090);
or U24639 (N_24639,N_15401,N_16121);
and U24640 (N_24640,N_15943,N_16737);
nor U24641 (N_24641,N_17695,N_16787);
nor U24642 (N_24642,N_15088,N_19909);
nor U24643 (N_24643,N_15644,N_19605);
or U24644 (N_24644,N_19491,N_16182);
nand U24645 (N_24645,N_19669,N_16913);
nand U24646 (N_24646,N_18733,N_16838);
or U24647 (N_24647,N_18525,N_17026);
or U24648 (N_24648,N_18403,N_16564);
or U24649 (N_24649,N_19431,N_19042);
nor U24650 (N_24650,N_19413,N_16690);
or U24651 (N_24651,N_16698,N_15730);
nor U24652 (N_24652,N_18158,N_19764);
and U24653 (N_24653,N_17719,N_19887);
nor U24654 (N_24654,N_19822,N_18046);
and U24655 (N_24655,N_19969,N_17144);
and U24656 (N_24656,N_15390,N_17789);
and U24657 (N_24657,N_19866,N_18301);
or U24658 (N_24658,N_19164,N_17207);
and U24659 (N_24659,N_17951,N_16887);
or U24660 (N_24660,N_17202,N_19339);
and U24661 (N_24661,N_16953,N_18347);
nand U24662 (N_24662,N_15539,N_19906);
nand U24663 (N_24663,N_18295,N_18125);
nand U24664 (N_24664,N_15383,N_17161);
or U24665 (N_24665,N_19300,N_16627);
or U24666 (N_24666,N_17560,N_16577);
nand U24667 (N_24667,N_19845,N_18664);
nor U24668 (N_24668,N_15569,N_18805);
and U24669 (N_24669,N_16119,N_18828);
and U24670 (N_24670,N_17579,N_18798);
nor U24671 (N_24671,N_15274,N_18100);
and U24672 (N_24672,N_16774,N_17714);
nand U24673 (N_24673,N_19043,N_15488);
and U24674 (N_24674,N_17098,N_16652);
nand U24675 (N_24675,N_15302,N_15292);
and U24676 (N_24676,N_15439,N_15396);
nand U24677 (N_24677,N_15908,N_17251);
and U24678 (N_24678,N_17456,N_16992);
nor U24679 (N_24679,N_16060,N_17785);
nand U24680 (N_24680,N_16714,N_15830);
nand U24681 (N_24681,N_17780,N_18383);
xor U24682 (N_24682,N_15933,N_17333);
or U24683 (N_24683,N_17787,N_16912);
or U24684 (N_24684,N_16126,N_18682);
and U24685 (N_24685,N_15407,N_17096);
nand U24686 (N_24686,N_15871,N_18845);
nand U24687 (N_24687,N_19930,N_15088);
nor U24688 (N_24688,N_19255,N_15017);
nand U24689 (N_24689,N_15975,N_18198);
nand U24690 (N_24690,N_16994,N_17128);
or U24691 (N_24691,N_16218,N_19088);
nor U24692 (N_24692,N_15488,N_17150);
and U24693 (N_24693,N_17944,N_17873);
nor U24694 (N_24694,N_15744,N_18981);
and U24695 (N_24695,N_15997,N_17928);
xnor U24696 (N_24696,N_18167,N_17093);
nand U24697 (N_24697,N_19953,N_15245);
and U24698 (N_24698,N_18019,N_16514);
nand U24699 (N_24699,N_17250,N_16875);
and U24700 (N_24700,N_18508,N_15447);
or U24701 (N_24701,N_18656,N_16100);
and U24702 (N_24702,N_18024,N_16204);
nand U24703 (N_24703,N_19836,N_15764);
nor U24704 (N_24704,N_16062,N_17986);
nor U24705 (N_24705,N_15340,N_16571);
and U24706 (N_24706,N_19948,N_19580);
nor U24707 (N_24707,N_15372,N_19136);
nand U24708 (N_24708,N_17184,N_19553);
nand U24709 (N_24709,N_16580,N_15917);
nor U24710 (N_24710,N_15758,N_17089);
and U24711 (N_24711,N_19637,N_18386);
and U24712 (N_24712,N_16127,N_18455);
xnor U24713 (N_24713,N_19185,N_19740);
nor U24714 (N_24714,N_19009,N_15898);
or U24715 (N_24715,N_15170,N_16163);
nor U24716 (N_24716,N_15696,N_19220);
and U24717 (N_24717,N_17280,N_19043);
nand U24718 (N_24718,N_19871,N_19821);
nand U24719 (N_24719,N_19627,N_17236);
nor U24720 (N_24720,N_15423,N_16665);
or U24721 (N_24721,N_15189,N_17593);
and U24722 (N_24722,N_15377,N_18213);
nand U24723 (N_24723,N_17247,N_19393);
nand U24724 (N_24724,N_18649,N_18826);
or U24725 (N_24725,N_18506,N_18027);
and U24726 (N_24726,N_17983,N_18522);
and U24727 (N_24727,N_19893,N_19235);
or U24728 (N_24728,N_17942,N_15098);
nand U24729 (N_24729,N_15653,N_19696);
nand U24730 (N_24730,N_19438,N_18719);
and U24731 (N_24731,N_16241,N_15231);
nand U24732 (N_24732,N_18268,N_17151);
nand U24733 (N_24733,N_16698,N_17754);
and U24734 (N_24734,N_16414,N_16016);
or U24735 (N_24735,N_17403,N_19344);
nor U24736 (N_24736,N_19966,N_19673);
nand U24737 (N_24737,N_16129,N_17612);
and U24738 (N_24738,N_19078,N_19225);
nor U24739 (N_24739,N_16815,N_17220);
and U24740 (N_24740,N_15628,N_15822);
and U24741 (N_24741,N_19104,N_17324);
xor U24742 (N_24742,N_17605,N_17899);
nor U24743 (N_24743,N_18055,N_19574);
or U24744 (N_24744,N_17083,N_16247);
nor U24745 (N_24745,N_19128,N_18533);
and U24746 (N_24746,N_18511,N_19249);
or U24747 (N_24747,N_18846,N_16365);
and U24748 (N_24748,N_16880,N_15045);
nand U24749 (N_24749,N_15617,N_18059);
or U24750 (N_24750,N_17367,N_18856);
xor U24751 (N_24751,N_16076,N_19623);
or U24752 (N_24752,N_16636,N_15969);
and U24753 (N_24753,N_19358,N_16776);
nor U24754 (N_24754,N_18371,N_19124);
nand U24755 (N_24755,N_19208,N_17302);
and U24756 (N_24756,N_18109,N_16330);
or U24757 (N_24757,N_17135,N_19487);
or U24758 (N_24758,N_18248,N_18852);
and U24759 (N_24759,N_19643,N_19193);
or U24760 (N_24760,N_19792,N_15042);
or U24761 (N_24761,N_18420,N_18666);
and U24762 (N_24762,N_15788,N_18438);
or U24763 (N_24763,N_17196,N_15042);
nor U24764 (N_24764,N_15499,N_18899);
or U24765 (N_24765,N_19001,N_16474);
or U24766 (N_24766,N_19124,N_18953);
and U24767 (N_24767,N_15580,N_19716);
xnor U24768 (N_24768,N_19858,N_19572);
nand U24769 (N_24769,N_16387,N_15513);
or U24770 (N_24770,N_16355,N_19794);
nor U24771 (N_24771,N_17474,N_15211);
nor U24772 (N_24772,N_17537,N_19584);
and U24773 (N_24773,N_18774,N_16137);
nor U24774 (N_24774,N_16506,N_19492);
or U24775 (N_24775,N_19956,N_19974);
and U24776 (N_24776,N_17498,N_19812);
and U24777 (N_24777,N_19331,N_18259);
nor U24778 (N_24778,N_19529,N_15787);
and U24779 (N_24779,N_18635,N_15220);
nor U24780 (N_24780,N_18753,N_17908);
and U24781 (N_24781,N_18627,N_19074);
xnor U24782 (N_24782,N_16945,N_19028);
nor U24783 (N_24783,N_19512,N_16129);
nand U24784 (N_24784,N_16223,N_15877);
nand U24785 (N_24785,N_15128,N_17423);
nand U24786 (N_24786,N_17313,N_19232);
and U24787 (N_24787,N_16712,N_19524);
nor U24788 (N_24788,N_15449,N_17510);
and U24789 (N_24789,N_17490,N_15186);
nor U24790 (N_24790,N_17065,N_16456);
nand U24791 (N_24791,N_18847,N_15641);
or U24792 (N_24792,N_18558,N_19087);
and U24793 (N_24793,N_19874,N_16505);
or U24794 (N_24794,N_18977,N_15792);
and U24795 (N_24795,N_18186,N_17083);
nand U24796 (N_24796,N_19298,N_19078);
nand U24797 (N_24797,N_19651,N_18620);
or U24798 (N_24798,N_15714,N_15602);
or U24799 (N_24799,N_19414,N_18717);
or U24800 (N_24800,N_18197,N_19501);
nor U24801 (N_24801,N_18124,N_19420);
nand U24802 (N_24802,N_16707,N_16208);
nor U24803 (N_24803,N_17701,N_17562);
or U24804 (N_24804,N_17795,N_19413);
nor U24805 (N_24805,N_17198,N_16122);
nor U24806 (N_24806,N_16063,N_17841);
nand U24807 (N_24807,N_19476,N_17031);
or U24808 (N_24808,N_16414,N_18503);
and U24809 (N_24809,N_19627,N_15845);
nand U24810 (N_24810,N_17447,N_15640);
nor U24811 (N_24811,N_18676,N_18129);
and U24812 (N_24812,N_15524,N_18812);
nand U24813 (N_24813,N_18481,N_18272);
nor U24814 (N_24814,N_19954,N_18387);
nor U24815 (N_24815,N_15061,N_17752);
or U24816 (N_24816,N_17406,N_17409);
nor U24817 (N_24817,N_16942,N_16068);
nor U24818 (N_24818,N_17774,N_16225);
and U24819 (N_24819,N_15181,N_18086);
nor U24820 (N_24820,N_19563,N_16991);
or U24821 (N_24821,N_16083,N_18089);
and U24822 (N_24822,N_19183,N_19463);
nand U24823 (N_24823,N_17331,N_19961);
nand U24824 (N_24824,N_18395,N_16851);
nor U24825 (N_24825,N_16005,N_15128);
and U24826 (N_24826,N_18894,N_17577);
or U24827 (N_24827,N_16451,N_17693);
and U24828 (N_24828,N_19873,N_15246);
nor U24829 (N_24829,N_15539,N_17251);
nand U24830 (N_24830,N_15819,N_19784);
or U24831 (N_24831,N_17617,N_19653);
nand U24832 (N_24832,N_15249,N_18631);
or U24833 (N_24833,N_19618,N_16230);
nor U24834 (N_24834,N_17316,N_17319);
nand U24835 (N_24835,N_18893,N_16496);
nand U24836 (N_24836,N_16590,N_19755);
nand U24837 (N_24837,N_17832,N_19575);
and U24838 (N_24838,N_16921,N_15148);
nand U24839 (N_24839,N_16748,N_15739);
and U24840 (N_24840,N_18523,N_17379);
or U24841 (N_24841,N_15748,N_18404);
or U24842 (N_24842,N_17713,N_17105);
nor U24843 (N_24843,N_15523,N_15333);
and U24844 (N_24844,N_17496,N_18059);
nor U24845 (N_24845,N_17192,N_18435);
or U24846 (N_24846,N_16728,N_15979);
or U24847 (N_24847,N_15778,N_19367);
or U24848 (N_24848,N_18440,N_17240);
and U24849 (N_24849,N_19848,N_16472);
or U24850 (N_24850,N_15092,N_15799);
nand U24851 (N_24851,N_16748,N_16761);
or U24852 (N_24852,N_18083,N_18488);
nor U24853 (N_24853,N_16242,N_16515);
nor U24854 (N_24854,N_18922,N_18993);
nand U24855 (N_24855,N_18785,N_18776);
nor U24856 (N_24856,N_19532,N_17184);
or U24857 (N_24857,N_19847,N_18410);
or U24858 (N_24858,N_15412,N_16130);
and U24859 (N_24859,N_18505,N_19512);
and U24860 (N_24860,N_18301,N_18198);
and U24861 (N_24861,N_16482,N_18151);
nor U24862 (N_24862,N_17390,N_17261);
or U24863 (N_24863,N_16324,N_15072);
or U24864 (N_24864,N_17814,N_16454);
or U24865 (N_24865,N_17636,N_19857);
and U24866 (N_24866,N_17743,N_17045);
nor U24867 (N_24867,N_15135,N_18744);
nand U24868 (N_24868,N_17000,N_16467);
and U24869 (N_24869,N_18433,N_15384);
and U24870 (N_24870,N_15279,N_18131);
nor U24871 (N_24871,N_18332,N_19485);
nor U24872 (N_24872,N_15147,N_17841);
or U24873 (N_24873,N_17181,N_16001);
nand U24874 (N_24874,N_17119,N_16802);
and U24875 (N_24875,N_19124,N_15271);
or U24876 (N_24876,N_17814,N_15121);
nor U24877 (N_24877,N_15191,N_19299);
and U24878 (N_24878,N_18592,N_15688);
or U24879 (N_24879,N_18333,N_15652);
or U24880 (N_24880,N_17364,N_17051);
nor U24881 (N_24881,N_16862,N_15009);
and U24882 (N_24882,N_15036,N_17213);
or U24883 (N_24883,N_15363,N_17435);
nor U24884 (N_24884,N_15318,N_19168);
nor U24885 (N_24885,N_17823,N_16618);
and U24886 (N_24886,N_15928,N_19591);
nand U24887 (N_24887,N_17826,N_17213);
or U24888 (N_24888,N_15606,N_19435);
nor U24889 (N_24889,N_16212,N_15350);
nor U24890 (N_24890,N_19545,N_19272);
nor U24891 (N_24891,N_19899,N_19716);
nor U24892 (N_24892,N_19962,N_19121);
xnor U24893 (N_24893,N_15839,N_17107);
nor U24894 (N_24894,N_18966,N_18575);
or U24895 (N_24895,N_17260,N_18593);
xor U24896 (N_24896,N_18082,N_19070);
and U24897 (N_24897,N_17391,N_16544);
nand U24898 (N_24898,N_16141,N_17298);
or U24899 (N_24899,N_17261,N_15328);
nor U24900 (N_24900,N_15950,N_19406);
or U24901 (N_24901,N_17472,N_19230);
nand U24902 (N_24902,N_17538,N_19481);
nand U24903 (N_24903,N_15086,N_17117);
or U24904 (N_24904,N_16484,N_16539);
nor U24905 (N_24905,N_19513,N_19550);
nand U24906 (N_24906,N_17604,N_15985);
nor U24907 (N_24907,N_16112,N_16599);
or U24908 (N_24908,N_17916,N_18639);
nand U24909 (N_24909,N_16237,N_19095);
and U24910 (N_24910,N_19064,N_16879);
and U24911 (N_24911,N_15782,N_18409);
nor U24912 (N_24912,N_15650,N_19225);
nand U24913 (N_24913,N_15070,N_16901);
xnor U24914 (N_24914,N_18092,N_17272);
nor U24915 (N_24915,N_16860,N_16794);
or U24916 (N_24916,N_15116,N_19157);
or U24917 (N_24917,N_19442,N_19480);
or U24918 (N_24918,N_15198,N_15974);
or U24919 (N_24919,N_17843,N_16489);
or U24920 (N_24920,N_19823,N_18047);
and U24921 (N_24921,N_17998,N_17564);
and U24922 (N_24922,N_18329,N_15702);
nand U24923 (N_24923,N_16031,N_15519);
and U24924 (N_24924,N_17697,N_16204);
nand U24925 (N_24925,N_19362,N_16280);
and U24926 (N_24926,N_19887,N_18864);
nand U24927 (N_24927,N_15666,N_17195);
xor U24928 (N_24928,N_18864,N_16435);
or U24929 (N_24929,N_15085,N_19491);
nor U24930 (N_24930,N_15243,N_16330);
or U24931 (N_24931,N_16253,N_15118);
and U24932 (N_24932,N_16932,N_18853);
and U24933 (N_24933,N_16213,N_16455);
nand U24934 (N_24934,N_16763,N_15409);
and U24935 (N_24935,N_17183,N_19421);
and U24936 (N_24936,N_17044,N_19299);
or U24937 (N_24937,N_15234,N_17225);
nand U24938 (N_24938,N_16764,N_18931);
and U24939 (N_24939,N_17888,N_15887);
and U24940 (N_24940,N_18126,N_15438);
or U24941 (N_24941,N_15504,N_15620);
xnor U24942 (N_24942,N_18237,N_18881);
nor U24943 (N_24943,N_17213,N_18135);
nand U24944 (N_24944,N_19736,N_18606);
nor U24945 (N_24945,N_17510,N_18943);
nor U24946 (N_24946,N_16605,N_19702);
or U24947 (N_24947,N_16804,N_19275);
and U24948 (N_24948,N_15954,N_19525);
nand U24949 (N_24949,N_16187,N_15912);
and U24950 (N_24950,N_19652,N_18544);
nor U24951 (N_24951,N_16693,N_15358);
and U24952 (N_24952,N_18559,N_17146);
or U24953 (N_24953,N_16999,N_17709);
or U24954 (N_24954,N_18616,N_19603);
nor U24955 (N_24955,N_17586,N_16713);
and U24956 (N_24956,N_15895,N_19674);
and U24957 (N_24957,N_19310,N_19430);
and U24958 (N_24958,N_17313,N_18117);
nor U24959 (N_24959,N_15383,N_17955);
nor U24960 (N_24960,N_16950,N_15042);
nand U24961 (N_24961,N_16617,N_19317);
nand U24962 (N_24962,N_15058,N_16986);
or U24963 (N_24963,N_18573,N_17620);
and U24964 (N_24964,N_15132,N_17671);
and U24965 (N_24965,N_17978,N_18181);
nand U24966 (N_24966,N_18197,N_16510);
and U24967 (N_24967,N_18914,N_17888);
or U24968 (N_24968,N_17121,N_17348);
or U24969 (N_24969,N_16491,N_19452);
and U24970 (N_24970,N_15732,N_17378);
and U24971 (N_24971,N_17191,N_15760);
nand U24972 (N_24972,N_19181,N_18942);
and U24973 (N_24973,N_15178,N_17214);
nor U24974 (N_24974,N_15863,N_15231);
and U24975 (N_24975,N_18934,N_17629);
and U24976 (N_24976,N_16479,N_19880);
nor U24977 (N_24977,N_17974,N_16925);
nand U24978 (N_24978,N_18442,N_18221);
nand U24979 (N_24979,N_17516,N_18560);
nand U24980 (N_24980,N_18116,N_17655);
nor U24981 (N_24981,N_15899,N_17104);
nand U24982 (N_24982,N_15476,N_15550);
and U24983 (N_24983,N_16815,N_17194);
or U24984 (N_24984,N_19406,N_18533);
or U24985 (N_24985,N_15095,N_16734);
nor U24986 (N_24986,N_16710,N_18896);
nand U24987 (N_24987,N_19687,N_17373);
and U24988 (N_24988,N_15121,N_17955);
or U24989 (N_24989,N_15061,N_17551);
or U24990 (N_24990,N_19382,N_18484);
nor U24991 (N_24991,N_18589,N_16922);
nand U24992 (N_24992,N_15022,N_17909);
and U24993 (N_24993,N_15086,N_19826);
xor U24994 (N_24994,N_16926,N_18373);
and U24995 (N_24995,N_16493,N_17943);
and U24996 (N_24996,N_16046,N_18195);
nand U24997 (N_24997,N_19835,N_18403);
nand U24998 (N_24998,N_19820,N_18929);
nand U24999 (N_24999,N_17921,N_18812);
and UO_0 (O_0,N_24490,N_20964);
nand UO_1 (O_1,N_24110,N_23718);
nand UO_2 (O_2,N_24882,N_23640);
and UO_3 (O_3,N_23984,N_23288);
nand UO_4 (O_4,N_21931,N_21684);
nor UO_5 (O_5,N_23180,N_24706);
nand UO_6 (O_6,N_22722,N_23780);
nor UO_7 (O_7,N_21746,N_22659);
nand UO_8 (O_8,N_20838,N_22434);
or UO_9 (O_9,N_23281,N_23460);
and UO_10 (O_10,N_22804,N_20966);
or UO_11 (O_11,N_24446,N_24371);
nand UO_12 (O_12,N_20733,N_22065);
nand UO_13 (O_13,N_21258,N_24941);
nand UO_14 (O_14,N_20318,N_20083);
or UO_15 (O_15,N_21210,N_22921);
and UO_16 (O_16,N_21159,N_20165);
or UO_17 (O_17,N_21731,N_21094);
nand UO_18 (O_18,N_20128,N_21079);
and UO_19 (O_19,N_24937,N_24125);
or UO_20 (O_20,N_20059,N_21398);
nor UO_21 (O_21,N_23435,N_23500);
nor UO_22 (O_22,N_22574,N_24903);
nor UO_23 (O_23,N_22932,N_21471);
nor UO_24 (O_24,N_21757,N_23765);
and UO_25 (O_25,N_23998,N_23709);
and UO_26 (O_26,N_21744,N_20276);
nand UO_27 (O_27,N_22358,N_24392);
nand UO_28 (O_28,N_22644,N_20492);
nor UO_29 (O_29,N_22918,N_20396);
nand UO_30 (O_30,N_21327,N_20946);
and UO_31 (O_31,N_22144,N_21638);
nor UO_32 (O_32,N_21752,N_22159);
and UO_33 (O_33,N_24845,N_21206);
and UO_34 (O_34,N_20412,N_20445);
and UO_35 (O_35,N_20817,N_22118);
and UO_36 (O_36,N_20006,N_22108);
xor UO_37 (O_37,N_20973,N_24766);
nand UO_38 (O_38,N_22189,N_22666);
or UO_39 (O_39,N_21216,N_23600);
nand UO_40 (O_40,N_23262,N_24993);
and UO_41 (O_41,N_20827,N_24409);
or UO_42 (O_42,N_20545,N_21552);
nand UO_43 (O_43,N_22606,N_22853);
nand UO_44 (O_44,N_22436,N_22753);
nand UO_45 (O_45,N_22775,N_21445);
or UO_46 (O_46,N_20155,N_23991);
or UO_47 (O_47,N_22825,N_23205);
or UO_48 (O_48,N_21771,N_21228);
and UO_49 (O_49,N_22640,N_23565);
and UO_50 (O_50,N_22662,N_22878);
or UO_51 (O_51,N_21201,N_23093);
or UO_52 (O_52,N_24948,N_20609);
nor UO_53 (O_53,N_24359,N_20661);
nand UO_54 (O_54,N_24986,N_20452);
nor UO_55 (O_55,N_21676,N_21839);
nor UO_56 (O_56,N_24553,N_20259);
and UO_57 (O_57,N_20951,N_23446);
nor UO_58 (O_58,N_21918,N_21399);
nor UO_59 (O_59,N_23508,N_21468);
or UO_60 (O_60,N_22516,N_21437);
nand UO_61 (O_61,N_21775,N_24761);
nand UO_62 (O_62,N_21707,N_23261);
or UO_63 (O_63,N_21174,N_20715);
or UO_64 (O_64,N_23485,N_23767);
nor UO_65 (O_65,N_21614,N_23029);
and UO_66 (O_66,N_21902,N_24032);
or UO_67 (O_67,N_24156,N_23252);
nor UO_68 (O_68,N_21211,N_22546);
nor UO_69 (O_69,N_20922,N_21974);
and UO_70 (O_70,N_23422,N_23987);
nand UO_71 (O_71,N_21263,N_22768);
or UO_72 (O_72,N_21161,N_24978);
nor UO_73 (O_73,N_22355,N_23358);
nand UO_74 (O_74,N_20927,N_24206);
nand UO_75 (O_75,N_24456,N_20408);
nor UO_76 (O_76,N_22415,N_23650);
and UO_77 (O_77,N_23363,N_21591);
and UO_78 (O_78,N_20269,N_22622);
nor UO_79 (O_79,N_23339,N_23254);
nand UO_80 (O_80,N_23213,N_23246);
and UO_81 (O_81,N_24234,N_23057);
or UO_82 (O_82,N_20806,N_23831);
or UO_83 (O_83,N_23175,N_21182);
or UO_84 (O_84,N_22255,N_24000);
nor UO_85 (O_85,N_22981,N_20509);
nor UO_86 (O_86,N_22519,N_20892);
nand UO_87 (O_87,N_23668,N_24135);
or UO_88 (O_88,N_21240,N_21451);
nand UO_89 (O_89,N_22506,N_24150);
nand UO_90 (O_90,N_22429,N_20608);
and UO_91 (O_91,N_22154,N_20461);
and UO_92 (O_92,N_24900,N_22368);
or UO_93 (O_93,N_21932,N_20521);
or UO_94 (O_94,N_21589,N_22010);
or UO_95 (O_95,N_24265,N_24231);
nand UO_96 (O_96,N_21338,N_24038);
and UO_97 (O_97,N_21654,N_20582);
nand UO_98 (O_98,N_24057,N_24830);
xnor UO_99 (O_99,N_21652,N_23675);
or UO_100 (O_100,N_20907,N_23226);
nand UO_101 (O_101,N_24537,N_24756);
or UO_102 (O_102,N_20302,N_24893);
and UO_103 (O_103,N_23577,N_22289);
or UO_104 (O_104,N_23691,N_23857);
and UO_105 (O_105,N_22317,N_22861);
nor UO_106 (O_106,N_23316,N_21186);
nand UO_107 (O_107,N_23391,N_24436);
nor UO_108 (O_108,N_20558,N_21950);
or UO_109 (O_109,N_20022,N_20961);
nand UO_110 (O_110,N_21660,N_23575);
nor UO_111 (O_111,N_21212,N_20679);
and UO_112 (O_112,N_21926,N_22504);
xnor UO_113 (O_113,N_24638,N_23834);
nor UO_114 (O_114,N_21070,N_21016);
xor UO_115 (O_115,N_20390,N_20926);
and UO_116 (O_116,N_24827,N_21307);
nand UO_117 (O_117,N_22969,N_22297);
or UO_118 (O_118,N_23352,N_23992);
nand UO_119 (O_119,N_22402,N_21925);
or UO_120 (O_120,N_20983,N_23805);
or UO_121 (O_121,N_23777,N_20754);
nand UO_122 (O_122,N_21082,N_23340);
and UO_123 (O_123,N_23940,N_21848);
nor UO_124 (O_124,N_20482,N_23383);
nor UO_125 (O_125,N_24533,N_21028);
or UO_126 (O_126,N_23404,N_21975);
nand UO_127 (O_127,N_22174,N_21215);
nor UO_128 (O_128,N_21528,N_24612);
xnor UO_129 (O_129,N_24095,N_21237);
nand UO_130 (O_130,N_22898,N_24796);
and UO_131 (O_131,N_24107,N_20965);
nand UO_132 (O_132,N_20583,N_23152);
xnor UO_133 (O_133,N_20316,N_21455);
and UO_134 (O_134,N_21345,N_23617);
and UO_135 (O_135,N_20264,N_20912);
xnor UO_136 (O_136,N_24445,N_21716);
and UO_137 (O_137,N_20695,N_20606);
nand UO_138 (O_138,N_20779,N_22551);
nand UO_139 (O_139,N_24179,N_21321);
and UO_140 (O_140,N_24485,N_22095);
nor UO_141 (O_141,N_22196,N_20923);
and UO_142 (O_142,N_23364,N_21012);
nor UO_143 (O_143,N_20291,N_20982);
or UO_144 (O_144,N_24825,N_20321);
or UO_145 (O_145,N_24417,N_24259);
nor UO_146 (O_146,N_22889,N_21244);
nor UO_147 (O_147,N_23696,N_22613);
nor UO_148 (O_148,N_23637,N_23924);
xnor UO_149 (O_149,N_23366,N_22202);
and UO_150 (O_150,N_20124,N_24894);
nand UO_151 (O_151,N_24718,N_22812);
nand UO_152 (O_152,N_20065,N_21875);
nor UO_153 (O_153,N_22617,N_20080);
nor UO_154 (O_154,N_20954,N_21639);
nor UO_155 (O_155,N_23414,N_22066);
or UO_156 (O_156,N_22822,N_23452);
or UO_157 (O_157,N_20389,N_23193);
nand UO_158 (O_158,N_20010,N_24593);
or UO_159 (O_159,N_22034,N_22470);
nand UO_160 (O_160,N_24588,N_22512);
nor UO_161 (O_161,N_24868,N_24608);
nor UO_162 (O_162,N_22782,N_23525);
nand UO_163 (O_163,N_24737,N_20672);
nor UO_164 (O_164,N_22684,N_23351);
nand UO_165 (O_165,N_21196,N_20913);
nand UO_166 (O_166,N_22230,N_22928);
nor UO_167 (O_167,N_22605,N_24073);
nand UO_168 (O_168,N_21063,N_21050);
nor UO_169 (O_169,N_22949,N_22961);
or UO_170 (O_170,N_21293,N_20601);
and UO_171 (O_171,N_23545,N_24580);
nor UO_172 (O_172,N_24838,N_23131);
or UO_173 (O_173,N_23549,N_24357);
nand UO_174 (O_174,N_24369,N_20114);
nand UO_175 (O_175,N_24366,N_23573);
or UO_176 (O_176,N_21694,N_22685);
or UO_177 (O_177,N_23682,N_22441);
nor UO_178 (O_178,N_22811,N_20930);
nor UO_179 (O_179,N_24988,N_22858);
nor UO_180 (O_180,N_24382,N_20924);
or UO_181 (O_181,N_24616,N_23529);
nand UO_182 (O_182,N_22176,N_24952);
nand UO_183 (O_183,N_22002,N_22270);
and UO_184 (O_184,N_21463,N_23304);
or UO_185 (O_185,N_22972,N_21904);
and UO_186 (O_186,N_20981,N_23027);
and UO_187 (O_187,N_20807,N_20953);
or UO_188 (O_188,N_21381,N_20737);
nor UO_189 (O_189,N_24972,N_20447);
nor UO_190 (O_190,N_22403,N_24667);
or UO_191 (O_191,N_20021,N_21722);
or UO_192 (O_192,N_21609,N_22071);
nand UO_193 (O_193,N_24386,N_24270);
nand UO_194 (O_194,N_22448,N_20699);
or UO_195 (O_195,N_21369,N_20014);
and UO_196 (O_196,N_22269,N_23438);
nor UO_197 (O_197,N_20100,N_20222);
or UO_198 (O_198,N_22696,N_22778);
nand UO_199 (O_199,N_20796,N_21986);
nor UO_200 (O_200,N_21059,N_20749);
and UO_201 (O_201,N_24657,N_24944);
or UO_202 (O_202,N_23056,N_20064);
nand UO_203 (O_203,N_21596,N_23865);
or UO_204 (O_204,N_20168,N_22978);
nor UO_205 (O_205,N_24636,N_21563);
or UO_206 (O_206,N_20840,N_24603);
nand UO_207 (O_207,N_21426,N_21120);
nand UO_208 (O_208,N_22654,N_22423);
xor UO_209 (O_209,N_22757,N_24431);
nand UO_210 (O_210,N_21852,N_20500);
nand UO_211 (O_211,N_24690,N_20283);
or UO_212 (O_212,N_22761,N_20795);
or UO_213 (O_213,N_21302,N_24904);
nor UO_214 (O_214,N_24506,N_24115);
nor UO_215 (O_215,N_21826,N_24330);
xnor UO_216 (O_216,N_23506,N_24679);
or UO_217 (O_217,N_23025,N_22234);
nor UO_218 (O_218,N_21319,N_21601);
nand UO_219 (O_219,N_22367,N_22924);
nor UO_220 (O_220,N_23970,N_21264);
or UO_221 (O_221,N_22123,N_23719);
nor UO_222 (O_222,N_22838,N_24124);
or UO_223 (O_223,N_21308,N_22560);
or UO_224 (O_224,N_22916,N_21077);
and UO_225 (O_225,N_24644,N_21666);
xnor UO_226 (O_226,N_20477,N_20287);
or UO_227 (O_227,N_23367,N_22345);
or UO_228 (O_228,N_23277,N_22321);
and UO_229 (O_229,N_24814,N_24731);
or UO_230 (O_230,N_23004,N_24130);
nor UO_231 (O_231,N_24983,N_22061);
and UO_232 (O_232,N_21149,N_21485);
nand UO_233 (O_233,N_20329,N_22211);
nor UO_234 (O_234,N_21243,N_23976);
or UO_235 (O_235,N_20734,N_20868);
and UO_236 (O_236,N_21667,N_21089);
nor UO_237 (O_237,N_22814,N_22287);
and UO_238 (O_238,N_22523,N_24284);
or UO_239 (O_239,N_24987,N_21655);
nand UO_240 (O_240,N_23921,N_20599);
nor UO_241 (O_241,N_22507,N_23464);
or UO_242 (O_242,N_24572,N_21780);
or UO_243 (O_243,N_23168,N_22735);
nand UO_244 (O_244,N_23278,N_22618);
or UO_245 (O_245,N_21583,N_22561);
and UO_246 (O_246,N_24397,N_21505);
or UO_247 (O_247,N_20766,N_20569);
and UO_248 (O_248,N_20540,N_20888);
and UO_249 (O_249,N_20675,N_21928);
and UO_250 (O_250,N_24458,N_24406);
nor UO_251 (O_251,N_24450,N_24811);
xor UO_252 (O_252,N_24077,N_21701);
or UO_253 (O_253,N_20593,N_24540);
and UO_254 (O_254,N_21980,N_23893);
nand UO_255 (O_255,N_22087,N_21976);
nand UO_256 (O_256,N_21085,N_24262);
nand UO_257 (O_257,N_23566,N_24875);
or UO_258 (O_258,N_24689,N_21661);
nand UO_259 (O_259,N_21984,N_24797);
nor UO_260 (O_260,N_22779,N_22306);
nor UO_261 (O_261,N_20422,N_20642);
or UO_262 (O_262,N_22678,N_24426);
nor UO_263 (O_263,N_24619,N_22182);
and UO_264 (O_264,N_23387,N_23729);
or UO_265 (O_265,N_20471,N_23109);
and UO_266 (O_266,N_20822,N_24907);
nand UO_267 (O_267,N_23178,N_21127);
or UO_268 (O_268,N_23299,N_23249);
and UO_269 (O_269,N_20305,N_24685);
and UO_270 (O_270,N_22938,N_23877);
nand UO_271 (O_271,N_24724,N_22937);
nand UO_272 (O_272,N_21170,N_22337);
or UO_273 (O_273,N_23049,N_23182);
or UO_274 (O_274,N_23771,N_23171);
nor UO_275 (O_275,N_23898,N_24097);
and UO_276 (O_276,N_22510,N_20296);
and UO_277 (O_277,N_20811,N_21372);
or UO_278 (O_278,N_24951,N_22899);
nor UO_279 (O_279,N_23842,N_23909);
and UO_280 (O_280,N_21409,N_23018);
and UO_281 (O_281,N_24622,N_22271);
nand UO_282 (O_282,N_21656,N_24563);
nand UO_283 (O_283,N_21927,N_24524);
or UO_284 (O_284,N_23815,N_24999);
nor UO_285 (O_285,N_23328,N_24854);
or UO_286 (O_286,N_20539,N_21823);
nor UO_287 (O_287,N_24692,N_23701);
and UO_288 (O_288,N_22895,N_23220);
and UO_289 (O_289,N_23493,N_22794);
nand UO_290 (O_290,N_23198,N_24696);
nand UO_291 (O_291,N_22464,N_22375);
and UO_292 (O_292,N_23875,N_24017);
nand UO_293 (O_293,N_24379,N_21286);
nand UO_294 (O_294,N_24361,N_22826);
nor UO_295 (O_295,N_20220,N_22480);
or UO_296 (O_296,N_21136,N_22896);
and UO_297 (O_297,N_21121,N_23658);
or UO_298 (O_298,N_21953,N_20654);
or UO_299 (O_299,N_24314,N_22704);
or UO_300 (O_300,N_24149,N_23016);
nor UO_301 (O_301,N_21693,N_21817);
nor UO_302 (O_302,N_23953,N_22428);
nand UO_303 (O_303,N_21122,N_24264);
nor UO_304 (O_304,N_20156,N_20074);
nand UO_305 (O_305,N_20327,N_23326);
and UO_306 (O_306,N_23135,N_22763);
nor UO_307 (O_307,N_23546,N_20476);
and UO_308 (O_308,N_20903,N_21886);
xnor UO_309 (O_309,N_22840,N_22747);
nand UO_310 (O_310,N_21856,N_22278);
or UO_311 (O_311,N_22503,N_24628);
and UO_312 (O_312,N_21424,N_21330);
nand UO_313 (O_313,N_22832,N_22450);
nor UO_314 (O_314,N_20058,N_22968);
nor UO_315 (O_315,N_20328,N_23775);
xor UO_316 (O_316,N_24278,N_23944);
and UO_317 (O_317,N_22310,N_22904);
nand UO_318 (O_318,N_23344,N_23216);
nand UO_319 (O_319,N_24243,N_22378);
and UO_320 (O_320,N_21725,N_24216);
or UO_321 (O_321,N_22730,N_20381);
or UO_322 (O_322,N_22101,N_21756);
nor UO_323 (O_323,N_23643,N_24958);
and UO_324 (O_324,N_22384,N_20303);
or UO_325 (O_325,N_23279,N_20893);
and UO_326 (O_326,N_24633,N_20752);
nand UO_327 (O_327,N_20219,N_20067);
and UO_328 (O_328,N_21720,N_23132);
xor UO_329 (O_329,N_22260,N_23950);
and UO_330 (O_330,N_23149,N_20768);
nor UO_331 (O_331,N_23601,N_22212);
or UO_332 (O_332,N_20194,N_22455);
xor UO_333 (O_333,N_20257,N_23702);
or UO_334 (O_334,N_21246,N_20292);
nor UO_335 (O_335,N_22712,N_22107);
nand UO_336 (O_336,N_20849,N_21483);
nor UO_337 (O_337,N_20392,N_24920);
or UO_338 (O_338,N_24559,N_20132);
nand UO_339 (O_339,N_22973,N_21699);
nand UO_340 (O_340,N_21824,N_22802);
nor UO_341 (O_341,N_24404,N_23878);
nand UO_342 (O_342,N_22721,N_24650);
nand UO_343 (O_343,N_23794,N_22307);
or UO_344 (O_344,N_23388,N_24926);
nor UO_345 (O_345,N_24437,N_21232);
xor UO_346 (O_346,N_21099,N_20306);
nor UO_347 (O_347,N_23502,N_22097);
nand UO_348 (O_348,N_23562,N_24851);
and UO_349 (O_349,N_21200,N_21313);
nor UO_350 (O_350,N_22357,N_20967);
nand UO_351 (O_351,N_20762,N_23954);
nand UO_352 (O_352,N_23870,N_23750);
or UO_353 (O_353,N_21000,N_22449);
nand UO_354 (O_354,N_23726,N_20998);
and UO_355 (O_355,N_24050,N_22670);
or UO_356 (O_356,N_22369,N_24185);
and UO_357 (O_357,N_21727,N_21758);
or UO_358 (O_358,N_24162,N_23542);
nor UO_359 (O_359,N_22746,N_23849);
nor UO_360 (O_360,N_22251,N_23440);
nor UO_361 (O_361,N_20794,N_24452);
or UO_362 (O_362,N_20190,N_22079);
nor UO_363 (O_363,N_22575,N_21815);
or UO_364 (O_364,N_20159,N_23959);
and UO_365 (O_365,N_23167,N_24080);
xnor UO_366 (O_366,N_22620,N_24775);
and UO_367 (O_367,N_22572,N_22282);
nor UO_368 (O_368,N_20855,N_23732);
nor UO_369 (O_369,N_23022,N_23443);
nor UO_370 (O_370,N_20110,N_21167);
or UO_371 (O_371,N_20170,N_22243);
and UO_372 (O_372,N_23517,N_21858);
and UO_373 (O_373,N_20720,N_20936);
nor UO_374 (O_374,N_23509,N_22513);
nor UO_375 (O_375,N_20107,N_20378);
and UO_376 (O_376,N_23163,N_22217);
nand UO_377 (O_377,N_22195,N_21990);
nand UO_378 (O_378,N_23059,N_22266);
or UO_379 (O_379,N_20862,N_21557);
or UO_380 (O_380,N_24841,N_22559);
nand UO_381 (O_381,N_21594,N_24784);
nand UO_382 (O_382,N_22914,N_24850);
nor UO_383 (O_383,N_24837,N_21977);
nor UO_384 (O_384,N_23519,N_24783);
and UO_385 (O_385,N_24739,N_21585);
nand UO_386 (O_386,N_23189,N_23406);
and UO_387 (O_387,N_20487,N_23720);
and UO_388 (O_388,N_24554,N_23431);
nand UO_389 (O_389,N_20181,N_21968);
nor UO_390 (O_390,N_23951,N_20620);
nand UO_391 (O_391,N_23156,N_20959);
or UO_392 (O_392,N_22328,N_21795);
and UO_393 (O_393,N_23782,N_21616);
nor UO_394 (O_394,N_21578,N_22294);
and UO_395 (O_395,N_21712,N_23392);
nor UO_396 (O_396,N_22036,N_23521);
and UO_397 (O_397,N_22229,N_20832);
or UO_398 (O_398,N_21550,N_23830);
xnor UO_399 (O_399,N_24326,N_20527);
or UO_400 (O_400,N_21023,N_20567);
and UO_401 (O_401,N_22518,N_20294);
nor UO_402 (O_402,N_23541,N_23801);
nor UO_403 (O_403,N_20861,N_20773);
and UO_404 (O_404,N_24045,N_20637);
nor UO_405 (O_405,N_24196,N_23080);
or UO_406 (O_406,N_20809,N_24096);
nand UO_407 (O_407,N_22766,N_22447);
nand UO_408 (O_408,N_22634,N_21091);
nor UO_409 (O_409,N_22445,N_23483);
nor UO_410 (O_410,N_22201,N_22153);
and UO_411 (O_411,N_23848,N_24843);
and UO_412 (O_412,N_20829,N_20193);
and UO_413 (O_413,N_21957,N_22422);
and UO_414 (O_414,N_21665,N_20345);
nand UO_415 (O_415,N_24912,N_21456);
nand UO_416 (O_416,N_22485,N_20577);
nand UO_417 (O_417,N_24448,N_21715);
nor UO_418 (O_418,N_21208,N_24961);
nor UO_419 (O_419,N_20858,N_23808);
or UO_420 (O_420,N_22024,N_20728);
or UO_421 (O_421,N_20008,N_20383);
nor UO_422 (O_422,N_22726,N_24488);
or UO_423 (O_423,N_24394,N_24982);
nor UO_424 (O_424,N_22293,N_20522);
and UO_425 (O_425,N_24024,N_20910);
nor UO_426 (O_426,N_20211,N_23348);
nand UO_427 (O_427,N_22602,N_21462);
or UO_428 (O_428,N_21385,N_20857);
and UO_429 (O_429,N_21179,N_20919);
and UO_430 (O_430,N_23218,N_24304);
and UO_431 (O_431,N_21311,N_23065);
nor UO_432 (O_432,N_23335,N_20813);
nand UO_433 (O_433,N_22073,N_23532);
nand UO_434 (O_434,N_20628,N_20721);
nor UO_435 (O_435,N_23449,N_21873);
nor UO_436 (O_436,N_23456,N_23539);
and UO_437 (O_437,N_20744,N_20043);
nor UO_438 (O_438,N_23302,N_21621);
nand UO_439 (O_439,N_24001,N_22709);
and UO_440 (O_440,N_21611,N_23883);
or UO_441 (O_441,N_24892,N_23162);
or UO_442 (O_442,N_23570,N_21157);
nor UO_443 (O_443,N_24886,N_22515);
nand UO_444 (O_444,N_23096,N_20799);
nand UO_445 (O_445,N_24871,N_24496);
nor UO_446 (O_446,N_24584,N_20034);
nor UO_447 (O_447,N_23749,N_22815);
xor UO_448 (O_448,N_21116,N_21628);
or UO_449 (O_449,N_22451,N_20578);
or UO_450 (O_450,N_24697,N_24810);
and UO_451 (O_451,N_21105,N_20130);
or UO_452 (O_452,N_24313,N_23122);
nor UO_453 (O_453,N_24911,N_23874);
and UO_454 (O_454,N_24175,N_24530);
and UO_455 (O_455,N_22134,N_24344);
nor UO_456 (O_456,N_21491,N_23257);
nor UO_457 (O_457,N_23212,N_22483);
or UO_458 (O_458,N_24672,N_20505);
and UO_459 (O_459,N_20340,N_22929);
or UO_460 (O_460,N_20202,N_20409);
xnor UO_461 (O_461,N_20828,N_22163);
and UO_462 (O_462,N_21499,N_23086);
nand UO_463 (O_463,N_21561,N_20191);
and UO_464 (O_464,N_24316,N_20039);
and UO_465 (O_465,N_23294,N_21640);
and UO_466 (O_466,N_21914,N_23999);
nor UO_467 (O_467,N_21484,N_21316);
or UO_468 (O_468,N_24155,N_23863);
and UO_469 (O_469,N_23614,N_20576);
or UO_470 (O_470,N_24088,N_21791);
xnor UO_471 (O_471,N_20691,N_23264);
or UO_472 (O_472,N_23856,N_24031);
nand UO_473 (O_473,N_21364,N_20723);
and UO_474 (O_474,N_23219,N_23918);
nor UO_475 (O_475,N_23173,N_23929);
nand UO_476 (O_476,N_20719,N_20393);
nor UO_477 (O_477,N_24544,N_24643);
nor UO_478 (O_478,N_23239,N_20437);
nand UO_479 (O_479,N_23873,N_21446);
nor UO_480 (O_480,N_21870,N_23561);
or UO_481 (O_481,N_21617,N_22089);
xor UO_482 (O_482,N_24505,N_24807);
nand UO_483 (O_483,N_21419,N_21115);
nor UO_484 (O_484,N_21230,N_21774);
nand UO_485 (O_485,N_24538,N_22740);
or UO_486 (O_486,N_21188,N_21650);
and UO_487 (O_487,N_22256,N_21075);
nand UO_488 (O_488,N_24592,N_24507);
nor UO_489 (O_489,N_24469,N_20013);
and UO_490 (O_490,N_21022,N_20091);
xnor UO_491 (O_491,N_20639,N_20777);
nor UO_492 (O_492,N_20253,N_21129);
or UO_493 (O_493,N_24755,N_22372);
or UO_494 (O_494,N_24678,N_20572);
and UO_495 (O_495,N_24717,N_22554);
nand UO_496 (O_496,N_24831,N_20357);
nor UO_497 (O_497,N_23832,N_22194);
or UO_498 (O_498,N_23957,N_20032);
nand UO_499 (O_499,N_24883,N_23926);
or UO_500 (O_500,N_23273,N_21348);
or UO_501 (O_501,N_20410,N_24430);
nand UO_502 (O_502,N_20182,N_24773);
nor UO_503 (O_503,N_21314,N_24033);
or UO_504 (O_504,N_23073,N_22109);
nand UO_505 (O_505,N_21921,N_20183);
nor UO_506 (O_506,N_22016,N_23628);
nand UO_507 (O_507,N_20689,N_21588);
and UO_508 (O_508,N_24627,N_21812);
nor UO_509 (O_509,N_23333,N_20687);
or UO_510 (O_510,N_24415,N_24372);
or UO_511 (O_511,N_22824,N_24116);
nand UO_512 (O_512,N_24671,N_23705);
or UO_513 (O_513,N_20493,N_20945);
nand UO_514 (O_514,N_22942,N_20872);
nand UO_515 (O_515,N_22276,N_24688);
and UO_516 (O_516,N_21155,N_24880);
and UO_517 (O_517,N_22412,N_22151);
nor UO_518 (O_518,N_21466,N_21525);
or UO_519 (O_519,N_23781,N_21982);
xnor UO_520 (O_520,N_21154,N_20075);
nor UO_521 (O_521,N_24774,N_20564);
and UO_522 (O_522,N_21592,N_22093);
or UO_523 (O_523,N_23111,N_21140);
or UO_524 (O_524,N_21490,N_23853);
nand UO_525 (O_525,N_24310,N_20650);
or UO_526 (O_526,N_21397,N_21416);
nor UO_527 (O_527,N_21641,N_23776);
xnor UO_528 (O_528,N_24929,N_22754);
nand UO_529 (O_529,N_21458,N_22253);
nor UO_530 (O_530,N_23956,N_20125);
nor UO_531 (O_531,N_21229,N_21770);
nand UO_532 (O_532,N_24898,N_20876);
or UO_533 (O_533,N_24018,N_20142);
xnor UO_534 (O_534,N_24932,N_23112);
and UO_535 (O_535,N_20942,N_24659);
nand UO_536 (O_536,N_20245,N_20789);
or UO_537 (O_537,N_21259,N_22386);
or UO_538 (O_538,N_23136,N_24081);
nand UO_539 (O_539,N_20076,N_24931);
nor UO_540 (O_540,N_23590,N_24617);
or UO_541 (O_541,N_20023,N_20985);
nor UO_542 (O_542,N_21645,N_20897);
xor UO_543 (O_543,N_20950,N_24562);
or UO_544 (O_544,N_22494,N_20821);
and UO_545 (O_545,N_22490,N_22508);
nor UO_546 (O_546,N_22931,N_21929);
and UO_547 (O_547,N_22579,N_22492);
and UO_548 (O_548,N_22370,N_20248);
nor UO_549 (O_549,N_21504,N_23434);
and UO_550 (O_550,N_24029,N_21498);
nor UO_551 (O_551,N_21710,N_24647);
or UO_552 (O_552,N_22244,N_24188);
and UO_553 (O_553,N_21547,N_23901);
xor UO_554 (O_554,N_23448,N_23116);
nor UO_555 (O_555,N_20490,N_22698);
nor UO_556 (O_556,N_22582,N_20753);
or UO_557 (O_557,N_20460,N_22841);
nand UO_558 (O_558,N_22162,N_22742);
nor UO_559 (O_559,N_20271,N_24566);
nor UO_560 (O_560,N_21124,N_21622);
nand UO_561 (O_561,N_22362,N_20596);
nand UO_562 (O_562,N_20463,N_22103);
nand UO_563 (O_563,N_23522,N_22142);
nor UO_564 (O_564,N_23169,N_21909);
and UO_565 (O_565,N_21708,N_20755);
nand UO_566 (O_566,N_22703,N_20956);
nor UO_567 (O_567,N_20604,N_21801);
or UO_568 (O_568,N_24235,N_21544);
and UO_569 (O_569,N_22420,N_21938);
nor UO_570 (O_570,N_22708,N_21788);
or UO_571 (O_571,N_21003,N_20592);
and UO_572 (O_572,N_23552,N_24703);
and UO_573 (O_573,N_23074,N_20388);
and UO_574 (O_574,N_22444,N_22267);
and UO_575 (O_575,N_21787,N_21646);
nor UO_576 (O_576,N_23747,N_24373);
nor UO_577 (O_577,N_22584,N_20638);
nor UO_578 (O_578,N_20207,N_20002);
nor UO_579 (O_579,N_24292,N_23044);
nand UO_580 (O_580,N_22477,N_24856);
or UO_581 (O_581,N_23948,N_23418);
and UO_582 (O_582,N_21959,N_23917);
nor UO_583 (O_583,N_24826,N_24614);
nor UO_584 (O_584,N_24639,N_20534);
nand UO_585 (O_585,N_21021,N_23664);
and UO_586 (O_586,N_23688,N_23572);
nor UO_587 (O_587,N_23607,N_24347);
or UO_588 (O_588,N_21804,N_21970);
and UO_589 (O_589,N_21342,N_23360);
nor UO_590 (O_590,N_21749,N_23994);
nor UO_591 (O_591,N_22971,N_21074);
and UO_592 (O_592,N_24860,N_21139);
nor UO_593 (O_593,N_24582,N_20629);
nor UO_594 (O_594,N_22406,N_24497);
or UO_595 (O_595,N_20096,N_21719);
and UO_596 (O_596,N_22501,N_23740);
xor UO_597 (O_597,N_24075,N_20859);
nor UO_598 (O_598,N_24339,N_23906);
nor UO_599 (O_599,N_24645,N_21090);
nor UO_600 (O_600,N_23370,N_23120);
or UO_601 (O_601,N_21797,N_23420);
or UO_602 (O_602,N_24381,N_22901);
or UO_603 (O_603,N_20311,N_20200);
or UO_604 (O_604,N_22992,N_21303);
nor UO_605 (O_605,N_23076,N_23911);
or UO_606 (O_606,N_23574,N_22130);
or UO_607 (O_607,N_24279,N_21422);
nor UO_608 (O_608,N_20844,N_21796);
nor UO_609 (O_609,N_20020,N_20761);
and UO_610 (O_610,N_22424,N_21438);
and UO_611 (O_611,N_22221,N_24611);
and UO_612 (O_612,N_24401,N_22498);
nor UO_613 (O_613,N_23647,N_24888);
and UO_614 (O_614,N_24771,N_21998);
or UO_615 (O_615,N_23158,N_23200);
and UO_616 (O_616,N_24061,N_20150);
or UO_617 (O_617,N_24172,N_24213);
nand UO_618 (O_618,N_20727,N_24176);
nor UO_619 (O_619,N_23454,N_21011);
or UO_620 (O_620,N_22393,N_21741);
and UO_621 (O_621,N_21930,N_23098);
nor UO_622 (O_622,N_23685,N_24652);
or UO_623 (O_623,N_21072,N_22945);
nand UO_624 (O_624,N_24848,N_22304);
or UO_625 (O_625,N_23206,N_23773);
nor UO_626 (O_626,N_21577,N_23265);
and UO_627 (O_627,N_24656,N_20237);
nand UO_628 (O_628,N_21613,N_23784);
or UO_629 (O_629,N_23300,N_23210);
or UO_630 (O_630,N_22788,N_22553);
nand UO_631 (O_631,N_24317,N_24010);
or UO_632 (O_632,N_20891,N_20785);
nand UO_633 (O_633,N_20914,N_22725);
nor UO_634 (O_634,N_24121,N_24670);
nand UO_635 (O_635,N_24294,N_21768);
and UO_636 (O_636,N_20431,N_24597);
nand UO_637 (O_637,N_23678,N_20580);
nand UO_638 (O_638,N_22785,N_22299);
and UO_639 (O_639,N_22541,N_21207);
nand UO_640 (O_640,N_22012,N_22674);
nor UO_641 (O_641,N_22600,N_20515);
nand UO_642 (O_642,N_20421,N_20173);
or UO_643 (O_643,N_21049,N_20512);
nand UO_644 (O_644,N_21647,N_21305);
nor UO_645 (O_645,N_23822,N_22146);
nor UO_646 (O_646,N_22543,N_20680);
and UO_647 (O_647,N_21256,N_23341);
nor UO_648 (O_648,N_23982,N_24577);
and UO_649 (O_649,N_21060,N_20201);
or UO_650 (O_650,N_21695,N_23321);
or UO_651 (O_651,N_20147,N_23155);
or UO_652 (O_652,N_23134,N_23034);
nand UO_653 (O_653,N_23672,N_24040);
or UO_654 (O_654,N_22866,N_21217);
nand UO_655 (O_655,N_24427,N_21729);
nand UO_656 (O_656,N_21546,N_23318);
nand UO_657 (O_657,N_24526,N_21737);
nand UO_658 (O_658,N_24816,N_20420);
nor UO_659 (O_659,N_24682,N_21353);
or UO_660 (O_660,N_23230,N_23094);
or UO_661 (O_661,N_23324,N_22873);
and UO_662 (O_662,N_24391,N_20788);
nor UO_663 (O_663,N_21387,N_24661);
xnor UO_664 (O_664,N_23141,N_20517);
and UO_665 (O_665,N_22114,N_24862);
nand UO_666 (O_666,N_20456,N_24859);
or UO_667 (O_667,N_20295,N_24187);
nor UO_668 (O_668,N_20700,N_22625);
or UO_669 (O_669,N_22636,N_20122);
nand UO_670 (O_670,N_22392,N_21663);
nor UO_671 (O_671,N_22366,N_23920);
nand UO_672 (O_672,N_21162,N_21067);
and UO_673 (O_673,N_20631,N_20688);
nand UO_674 (O_674,N_22091,N_24570);
or UO_675 (O_675,N_22183,N_20833);
nand UO_676 (O_676,N_23413,N_20198);
or UO_677 (O_677,N_22259,N_23932);
nor UO_678 (O_678,N_23645,N_23490);
xor UO_679 (O_679,N_21908,N_24324);
nor UO_680 (O_680,N_20106,N_21281);
nor UO_681 (O_681,N_21199,N_21555);
nor UO_682 (O_682,N_22209,N_23543);
xor UO_683 (O_683,N_23569,N_20771);
and UO_684 (O_684,N_20491,N_23484);
nor UO_685 (O_685,N_20049,N_21711);
and UO_686 (O_686,N_24762,N_21829);
nor UO_687 (O_687,N_21123,N_21160);
nor UO_688 (O_688,N_21678,N_20387);
or UO_689 (O_689,N_24668,N_20474);
nand UO_690 (O_690,N_22165,N_22975);
and UO_691 (O_691,N_23088,N_22350);
and UO_692 (O_692,N_21501,N_20450);
nor UO_693 (O_693,N_24863,N_21709);
nand UO_694 (O_694,N_20233,N_24380);
or UO_695 (O_695,N_22522,N_23965);
and UO_696 (O_696,N_24090,N_23481);
and UO_697 (O_697,N_22784,N_20144);
or UO_698 (O_698,N_20879,N_24305);
and UO_699 (O_699,N_23563,N_21052);
nor UO_700 (O_700,N_21825,N_21517);
xor UO_701 (O_701,N_24290,N_23587);
or UO_702 (O_702,N_22935,N_20187);
and UO_703 (O_703,N_22122,N_23635);
nor UO_704 (O_704,N_20341,N_20864);
nor UO_705 (O_705,N_22064,N_23028);
nor UO_706 (O_706,N_24519,N_24076);
and UO_707 (O_707,N_21093,N_23133);
nor UO_708 (O_708,N_20591,N_24306);
nor UO_709 (O_709,N_20089,N_20671);
and UO_710 (O_710,N_20589,N_21636);
nand UO_711 (O_711,N_23735,N_21562);
or UO_712 (O_712,N_22573,N_24020);
and UO_713 (O_713,N_24475,N_23661);
and UO_714 (O_714,N_22847,N_24145);
nand UO_715 (O_715,N_23746,N_24337);
or UO_716 (O_716,N_20775,N_20030);
and UO_717 (O_717,N_24895,N_24794);
and UO_718 (O_718,N_23296,N_22489);
nor UO_719 (O_719,N_23276,N_23745);
xor UO_720 (O_720,N_23269,N_21745);
and UO_721 (O_721,N_24189,N_24683);
and UO_722 (O_722,N_20231,N_22987);
nand UO_723 (O_723,N_24399,N_21776);
or UO_724 (O_724,N_23401,N_23774);
nor UO_725 (O_725,N_23390,N_23106);
and UO_726 (O_726,N_24642,N_20653);
or UO_727 (O_727,N_22771,N_20145);
and UO_728 (O_728,N_22440,N_23217);
and UO_729 (O_729,N_21283,N_22343);
and UO_730 (O_730,N_21602,N_21026);
nor UO_731 (O_731,N_20652,N_21278);
or UO_732 (O_732,N_23833,N_20146);
and UO_733 (O_733,N_21042,N_24151);
and UO_734 (O_734,N_21470,N_20630);
nand UO_735 (O_735,N_24801,N_22245);
nand UO_736 (O_736,N_20725,N_22713);
nand UO_737 (O_737,N_20898,N_20038);
and UO_738 (O_738,N_23902,N_22020);
nand UO_739 (O_739,N_24281,N_23931);
or UO_740 (O_740,N_22475,N_24098);
or UO_741 (O_741,N_24864,N_24037);
nor UO_742 (O_742,N_24268,N_20293);
nand UO_743 (O_743,N_24515,N_23751);
or UO_744 (O_744,N_21763,N_21511);
nand UO_745 (O_745,N_24494,N_21861);
nor UO_746 (O_746,N_21840,N_23648);
or UO_747 (O_747,N_20590,N_24174);
or UO_748 (O_748,N_22707,N_20299);
and UO_749 (O_749,N_22538,N_21610);
or UO_750 (O_750,N_21867,N_20717);
nand UO_751 (O_751,N_22032,N_20070);
and UO_752 (O_752,N_24955,N_20810);
nor UO_753 (O_753,N_20226,N_22765);
nor UO_754 (O_754,N_22115,N_23380);
or UO_755 (O_755,N_24821,N_22342);
nor UO_756 (O_756,N_22139,N_22926);
or UO_757 (O_757,N_23763,N_22571);
nor UO_758 (O_758,N_22875,N_24028);
nand UO_759 (O_759,N_21697,N_23433);
nor UO_760 (O_760,N_22152,N_20495);
xor UO_761 (O_761,N_21857,N_23896);
and UO_762 (O_762,N_21881,N_23686);
nor UO_763 (O_763,N_23934,N_22528);
nor UO_764 (O_764,N_24787,N_20585);
or UO_765 (O_765,N_24011,N_22021);
nand UO_766 (O_766,N_20473,N_24936);
and UO_767 (O_767,N_21062,N_21152);
nor UO_768 (O_768,N_22925,N_22789);
and UO_769 (O_769,N_20339,N_24414);
or UO_770 (O_770,N_21005,N_22124);
or UO_771 (O_771,N_24122,N_23235);
nor UO_772 (O_772,N_21282,N_20322);
or UO_773 (O_773,N_23530,N_22829);
or UO_774 (O_774,N_20344,N_21623);
nand UO_775 (O_775,N_24778,N_24803);
nor UO_776 (O_776,N_22246,N_24873);
or UO_777 (O_777,N_20722,N_20649);
and UO_778 (O_778,N_22806,N_21037);
and UO_779 (O_779,N_24541,N_23009);
nor UO_780 (O_780,N_22565,N_21047);
xnor UO_781 (O_781,N_23290,N_23819);
nand UO_782 (O_782,N_22453,N_20915);
nor UO_783 (O_783,N_22580,N_20875);
xnor UO_784 (O_784,N_22970,N_22381);
or UO_785 (O_785,N_22208,N_24068);
and UO_786 (O_786,N_24992,N_23892);
and UO_787 (O_787,N_21428,N_23512);
or UO_788 (O_788,N_24959,N_24829);
xor UO_789 (O_789,N_23538,N_20882);
nor UO_790 (O_790,N_23963,N_22192);
nor UO_791 (O_791,N_22380,N_23285);
and UO_792 (O_792,N_20665,N_23854);
nand UO_793 (O_793,N_22550,N_21371);
nand UO_794 (O_794,N_24093,N_21556);
or UO_795 (O_795,N_20488,N_21095);
nand UO_796 (O_796,N_21910,N_21431);
nor UO_797 (O_797,N_22249,N_24486);
nor UO_798 (O_798,N_21607,N_21352);
nand UO_799 (O_799,N_24743,N_23199);
and UO_800 (O_800,N_23221,N_23503);
nor UO_801 (O_801,N_21429,N_23609);
or UO_802 (O_802,N_23710,N_20575);
nand UO_803 (O_803,N_23184,N_20900);
nand UO_804 (O_804,N_22474,N_22974);
nor UO_805 (O_805,N_21488,N_20192);
nand UO_806 (O_806,N_24333,N_23524);
nand UO_807 (O_807,N_22643,N_20499);
nand UO_808 (O_808,N_21254,N_21325);
and UO_809 (O_809,N_23639,N_20149);
nand UO_810 (O_810,N_20109,N_24780);
and UO_811 (O_811,N_22791,N_20741);
or UO_812 (O_812,N_21117,N_20033);
and UO_813 (O_813,N_23303,N_20932);
or UO_814 (O_814,N_23342,N_23396);
nand UO_815 (O_815,N_24767,N_21535);
and UO_816 (O_816,N_22462,N_22312);
nand UO_817 (O_817,N_22922,N_24210);
or UO_818 (O_818,N_23047,N_23764);
or UO_819 (O_819,N_23862,N_20468);
nand UO_820 (O_820,N_24199,N_21537);
nand UO_821 (O_821,N_20469,N_23013);
nand UO_822 (O_822,N_21400,N_23376);
and UO_823 (O_823,N_22220,N_20823);
nand UO_824 (O_824,N_22479,N_21618);
and UO_825 (O_825,N_21298,N_24327);
or UO_826 (O_826,N_21326,N_20818);
nand UO_827 (O_827,N_22049,N_20479);
and UO_828 (O_828,N_20426,N_22689);
nor UO_829 (O_829,N_22223,N_20116);
and UO_830 (O_830,N_23003,N_21495);
xnor UO_831 (O_831,N_21312,N_20791);
nor UO_832 (O_832,N_24979,N_23827);
or UO_833 (O_833,N_23222,N_24990);
or UO_834 (O_834,N_21883,N_21777);
or UO_835 (O_835,N_22277,N_24207);
and UO_836 (O_836,N_20433,N_22595);
nor UO_837 (O_837,N_22564,N_20834);
nand UO_838 (O_838,N_24833,N_24709);
or UO_839 (O_839,N_21531,N_20407);
nand UO_840 (O_840,N_20581,N_20673);
nor UO_841 (O_841,N_22692,N_24008);
or UO_842 (O_842,N_20172,N_24177);
nor UO_843 (O_843,N_23128,N_22069);
or UO_844 (O_844,N_22953,N_22072);
and UO_845 (O_845,N_21169,N_21584);
or UO_846 (O_846,N_23855,N_24605);
nand UO_847 (O_847,N_20320,N_23791);
nor UO_848 (O_848,N_23807,N_22481);
and UO_849 (O_849,N_21334,N_23424);
nor UO_850 (O_850,N_20355,N_23505);
nand UO_851 (O_851,N_23298,N_22476);
and UO_852 (O_852,N_24131,N_23817);
nand UO_853 (O_853,N_22288,N_21767);
nor UO_854 (O_854,N_21444,N_22263);
nor UO_855 (O_855,N_22446,N_20758);
nor UO_856 (O_856,N_20310,N_20475);
nand UO_857 (O_857,N_22473,N_20851);
nor UO_858 (O_858,N_23280,N_23499);
or UO_859 (O_859,N_21222,N_21860);
nor UO_860 (O_860,N_23669,N_21390);
and UO_861 (O_861,N_21479,N_21057);
or UO_862 (O_862,N_24089,N_22701);
or UO_863 (O_863,N_22774,N_21033);
and UO_864 (O_864,N_21534,N_24750);
nor UO_865 (O_865,N_22389,N_24658);
nor UO_866 (O_866,N_20958,N_22919);
and UO_867 (O_867,N_20353,N_23263);
nand UO_868 (O_868,N_21078,N_24209);
and UO_869 (O_869,N_20356,N_24291);
nor UO_870 (O_870,N_21713,N_20203);
or UO_871 (O_871,N_23641,N_24167);
and UO_872 (O_872,N_23707,N_21043);
nand UO_873 (O_873,N_23103,N_20360);
nand UO_874 (O_874,N_24217,N_22604);
nand UO_875 (O_875,N_22354,N_20209);
nand UO_876 (O_876,N_23736,N_24143);
nand UO_877 (O_877,N_21635,N_22723);
nor UO_878 (O_878,N_20169,N_20137);
and UO_879 (O_879,N_24791,N_24004);
and UO_880 (O_880,N_22950,N_23608);
nor UO_881 (O_881,N_21176,N_20770);
xor UO_882 (O_882,N_22917,N_21669);
and UO_883 (O_883,N_22131,N_23554);
or UO_884 (O_884,N_21172,N_23325);
nor UO_885 (O_885,N_20373,N_21102);
or UO_886 (O_886,N_22976,N_23084);
or UO_887 (O_887,N_20645,N_22817);
and UO_888 (O_888,N_24922,N_22442);
or UO_889 (O_889,N_20786,N_24699);
nand UO_890 (O_890,N_24569,N_20802);
nand UO_891 (O_891,N_22727,N_23191);
and UO_892 (O_892,N_23186,N_21750);
nor UO_893 (O_893,N_21017,N_22593);
and UO_894 (O_894,N_21907,N_21295);
nor UO_895 (O_895,N_22887,N_21066);
nor UO_896 (O_896,N_20977,N_22557);
and UO_897 (O_897,N_24511,N_20764);
nand UO_898 (O_898,N_21036,N_22807);
nand UO_899 (O_899,N_20525,N_20312);
and UO_900 (O_900,N_22776,N_24869);
nand UO_901 (O_901,N_24367,N_24030);
and UO_902 (O_902,N_24484,N_24462);
nor UO_903 (O_903,N_20175,N_21171);
xor UO_904 (O_904,N_20750,N_21375);
or UO_905 (O_905,N_22621,N_21204);
or UO_906 (O_906,N_20315,N_23620);
nand UO_907 (O_907,N_22116,N_23194);
nor UO_908 (O_908,N_23450,N_23869);
or UO_909 (O_909,N_24201,N_24419);
nor UO_910 (O_910,N_20781,N_22009);
or UO_911 (O_911,N_24967,N_23979);
nor UO_912 (O_912,N_21356,N_22164);
or UO_913 (O_913,N_23204,N_23211);
nor UO_914 (O_914,N_23284,N_20297);
nor UO_915 (O_915,N_22236,N_23501);
or UO_916 (O_916,N_22491,N_21778);
nor UO_917 (O_917,N_20994,N_24763);
or UO_918 (O_918,N_24092,N_23757);
nor UO_919 (O_919,N_21262,N_21519);
nand UO_920 (O_920,N_21435,N_24285);
nand UO_921 (O_921,N_24499,N_22333);
or UO_922 (O_922,N_22262,N_20656);
nor UO_923 (O_923,N_22849,N_20889);
or UO_924 (O_924,N_22371,N_21605);
nor UO_925 (O_925,N_23087,N_22452);
and UO_926 (O_926,N_20757,N_20745);
or UO_927 (O_927,N_22298,N_21551);
or UO_928 (O_928,N_23779,N_20459);
or UO_929 (O_929,N_22081,N_24153);
nand UO_930 (O_930,N_23126,N_20979);
or UO_931 (O_931,N_22356,N_22694);
nor UO_932 (O_932,N_23489,N_22085);
nor UO_933 (O_933,N_21866,N_21800);
and UO_934 (O_934,N_20793,N_23876);
or UO_935 (O_935,N_22347,N_24318);
nand UO_936 (O_936,N_21747,N_24891);
or UO_937 (O_937,N_21692,N_22225);
and UO_938 (O_938,N_24144,N_20826);
nor UO_939 (O_939,N_20554,N_22856);
nor UO_940 (O_940,N_20934,N_20708);
nor UO_941 (O_941,N_24832,N_21978);
or UO_942 (O_942,N_22404,N_23904);
or UO_943 (O_943,N_22843,N_21138);
or UO_944 (O_944,N_20657,N_23868);
nor UO_945 (O_945,N_20997,N_20854);
nand UO_946 (O_946,N_20729,N_22111);
or UO_947 (O_947,N_24120,N_23208);
and UO_948 (O_948,N_24019,N_23301);
and UO_949 (O_949,N_21383,N_24621);
or UO_950 (O_950,N_24277,N_22170);
nor UO_951 (O_951,N_22456,N_22998);
nor UO_952 (O_952,N_22567,N_21792);
nand UO_953 (O_953,N_21404,N_22257);
or UO_954 (O_954,N_24924,N_20029);
nand UO_955 (O_955,N_21408,N_24710);
nor UO_956 (O_956,N_24915,N_21343);
or UO_957 (O_957,N_24909,N_24857);
and UO_958 (O_958,N_20366,N_22186);
and UO_959 (O_959,N_21472,N_20041);
and UO_960 (O_960,N_20284,N_23922);
and UO_961 (O_961,N_21682,N_20587);
or UO_962 (O_962,N_21425,N_21620);
and UO_963 (O_963,N_20503,N_23283);
nor UO_964 (O_964,N_24648,N_22214);
nand UO_965 (O_965,N_24694,N_21252);
xor UO_966 (O_966,N_23410,N_21738);
nor UO_967 (O_967,N_20713,N_24950);
and UO_968 (O_968,N_24522,N_20921);
nand UO_969 (O_969,N_24275,N_22029);
or UO_970 (O_970,N_20135,N_20423);
nand UO_971 (O_971,N_20238,N_24348);
nor UO_972 (O_972,N_24989,N_21361);
and UO_973 (O_973,N_22648,N_24820);
nand UO_974 (O_974,N_23914,N_21106);
and UO_975 (O_975,N_21192,N_22461);
or UO_976 (O_976,N_21933,N_20863);
and UO_977 (O_977,N_24133,N_24996);
nand UO_978 (O_978,N_24191,N_24631);
or UO_979 (O_979,N_23947,N_20677);
or UO_980 (O_980,N_24844,N_24640);
nor UO_981 (O_981,N_24684,N_22206);
xor UO_982 (O_982,N_20223,N_21734);
nor UO_983 (O_983,N_21339,N_22318);
and UO_984 (O_984,N_24890,N_20304);
and UO_985 (O_985,N_23268,N_23196);
and UO_986 (O_986,N_21759,N_24940);
or UO_987 (O_987,N_23997,N_20280);
nand UO_988 (O_988,N_21703,N_22880);
nand UO_989 (O_989,N_21934,N_24094);
or UO_990 (O_990,N_21261,N_24374);
nor UO_991 (O_991,N_23967,N_24815);
nand UO_992 (O_992,N_22008,N_20166);
nand UO_993 (O_993,N_21098,N_20415);
nand UO_994 (O_994,N_24808,N_20279);
nor UO_995 (O_995,N_21841,N_24148);
or UO_996 (O_996,N_21513,N_21449);
nand UO_997 (O_997,N_23083,N_20404);
and UO_998 (O_998,N_21285,N_24355);
xor UO_999 (O_999,N_21001,N_22545);
nor UO_1000 (O_1000,N_21581,N_21936);
or UO_1001 (O_1001,N_21963,N_24273);
or UO_1002 (O_1002,N_22999,N_20735);
and UO_1003 (O_1003,N_23240,N_24514);
nand UO_1004 (O_1004,N_22910,N_24768);
nand UO_1005 (O_1005,N_24681,N_22043);
and UO_1006 (O_1006,N_22891,N_24965);
nand UO_1007 (O_1007,N_24211,N_21053);
and UO_1008 (O_1008,N_23295,N_20562);
nor UO_1009 (O_1009,N_22982,N_24568);
nand UO_1010 (O_1010,N_22272,N_22933);
nor UO_1011 (O_1011,N_23627,N_20848);
nand UO_1012 (O_1012,N_23835,N_23759);
and UO_1013 (O_1013,N_20739,N_20372);
nor UO_1014 (O_1014,N_21507,N_24653);
nand UO_1015 (O_1015,N_22156,N_20704);
nand UO_1016 (O_1016,N_22664,N_20079);
and UO_1017 (O_1017,N_24233,N_22993);
or UO_1018 (O_1018,N_23250,N_21943);
and UO_1019 (O_1019,N_23271,N_22022);
or UO_1020 (O_1020,N_20714,N_23814);
nand UO_1021 (O_1021,N_20676,N_24014);
or UO_1022 (O_1022,N_24835,N_23527);
nand UO_1023 (O_1023,N_20548,N_22117);
nand UO_1024 (O_1024,N_24067,N_20004);
nand UO_1025 (O_1025,N_23728,N_22374);
nand UO_1026 (O_1026,N_21634,N_22138);
nor UO_1027 (O_1027,N_21835,N_24804);
or UO_1028 (O_1028,N_24457,N_21276);
nand UO_1029 (O_1029,N_24471,N_21855);
nand UO_1030 (O_1030,N_20718,N_24585);
xor UO_1031 (O_1031,N_20805,N_23913);
or UO_1032 (O_1032,N_23373,N_23715);
or UO_1033 (O_1033,N_21146,N_21224);
nor UO_1034 (O_1034,N_21392,N_21143);
or UO_1035 (O_1035,N_21659,N_20325);
and UO_1036 (O_1036,N_23568,N_21671);
or UO_1037 (O_1037,N_23398,N_21582);
nand UO_1038 (O_1038,N_22502,N_22752);
nand UO_1039 (O_1039,N_23330,N_22859);
nand UO_1040 (O_1040,N_21046,N_21350);
and UO_1041 (O_1041,N_22943,N_23308);
and UO_1042 (O_1042,N_21896,N_24637);
and UO_1043 (O_1043,N_20016,N_22338);
and UO_1044 (O_1044,N_21198,N_23806);
nor UO_1045 (O_1045,N_23385,N_24776);
nand UO_1046 (O_1046,N_24698,N_24970);
nand UO_1047 (O_1047,N_22870,N_24288);
or UO_1048 (O_1048,N_24980,N_22607);
or UO_1049 (O_1049,N_24106,N_20017);
nor UO_1050 (O_1050,N_22418,N_23514);
nor UO_1051 (O_1051,N_21674,N_22530);
and UO_1052 (O_1052,N_20380,N_21813);
nor UO_1053 (O_1053,N_23972,N_22860);
and UO_1054 (O_1054,N_23988,N_24253);
or UO_1055 (O_1055,N_20523,N_22329);
nand UO_1056 (O_1056,N_23192,N_24919);
and UO_1057 (O_1057,N_21142,N_20313);
nand UO_1058 (O_1058,N_21002,N_21493);
nor UO_1059 (O_1059,N_21845,N_23014);
nor UO_1060 (O_1060,N_21443,N_23354);
and UO_1061 (O_1061,N_23531,N_22332);
or UO_1062 (O_1062,N_22578,N_24525);
nor UO_1063 (O_1063,N_22598,N_20281);
and UO_1064 (O_1064,N_21790,N_23095);
nand UO_1065 (O_1065,N_21629,N_21065);
nor UO_1066 (O_1066,N_21341,N_24879);
and UO_1067 (O_1067,N_23470,N_23037);
or UO_1068 (O_1068,N_23144,N_23595);
nand UO_1069 (O_1069,N_22877,N_20991);
nand UO_1070 (O_1070,N_24197,N_21015);
or UO_1071 (O_1071,N_21101,N_23462);
and UO_1072 (O_1072,N_23105,N_22984);
and UO_1073 (O_1073,N_22786,N_23622);
and UO_1074 (O_1074,N_22397,N_20260);
and UO_1075 (O_1075,N_22027,N_22181);
nand UO_1076 (O_1076,N_21689,N_24132);
and UO_1077 (O_1077,N_24536,N_23006);
nand UO_1078 (O_1078,N_22110,N_22511);
and UO_1079 (O_1079,N_22790,N_23516);
or UO_1080 (O_1080,N_22762,N_20268);
and UO_1081 (O_1081,N_24781,N_20547);
nor UO_1082 (O_1082,N_20663,N_22524);
or UO_1083 (O_1083,N_24400,N_20842);
nand UO_1084 (O_1084,N_22232,N_21844);
nand UO_1085 (O_1085,N_24015,N_23187);
or UO_1086 (O_1086,N_23867,N_24748);
nand UO_1087 (O_1087,N_20035,N_21854);
and UO_1088 (O_1088,N_24403,N_24215);
and UO_1089 (O_1089,N_24725,N_23060);
nand UO_1090 (O_1090,N_22017,N_24842);
nor UO_1091 (O_1091,N_22376,N_21205);
and UO_1092 (O_1092,N_20262,N_23311);
nand UO_1093 (O_1093,N_24205,N_21233);
nand UO_1094 (O_1094,N_20438,N_22426);
nor UO_1095 (O_1095,N_24365,N_24735);
and UO_1096 (O_1096,N_24438,N_20068);
or UO_1097 (O_1097,N_23309,N_24727);
nand UO_1098 (O_1098,N_20536,N_20298);
nand UO_1099 (O_1099,N_20835,N_21755);
and UO_1100 (O_1100,N_24377,N_22172);
and UO_1101 (O_1101,N_20171,N_21332);
nor UO_1102 (O_1102,N_23772,N_21294);
nand UO_1103 (O_1103,N_23792,N_23166);
nand UO_1104 (O_1104,N_23345,N_21527);
nor UO_1105 (O_1105,N_23334,N_24509);
nor UO_1106 (O_1106,N_22222,N_21785);
nor UO_1107 (O_1107,N_22140,N_20635);
or UO_1108 (O_1108,N_23305,N_22330);
or UO_1109 (O_1109,N_20189,N_22652);
nor UO_1110 (O_1110,N_22728,N_20678);
or UO_1111 (O_1111,N_23306,N_21580);
nand UO_1112 (O_1112,N_24323,N_23942);
or UO_1113 (O_1113,N_24202,N_20972);
nand UO_1114 (O_1114,N_20414,N_23588);
and UO_1115 (O_1115,N_20746,N_23670);
and UO_1116 (O_1116,N_24977,N_22190);
nor UO_1117 (O_1117,N_23594,N_20494);
nor UO_1118 (O_1118,N_24049,N_20740);
or UO_1119 (O_1119,N_23559,N_22218);
and UO_1120 (O_1120,N_21723,N_21850);
or UO_1121 (O_1121,N_23317,N_23864);
or UO_1122 (O_1122,N_20546,N_20158);
nor UO_1123 (O_1123,N_23046,N_20055);
nand UO_1124 (O_1124,N_21355,N_20767);
and UO_1125 (O_1125,N_24332,N_23621);
nor UO_1126 (O_1126,N_21554,N_20706);
nand UO_1127 (O_1127,N_21164,N_20636);
nor UO_1128 (O_1128,N_22309,N_20097);
nor UO_1129 (O_1129,N_23458,N_24732);
and UO_1130 (O_1130,N_22886,N_21366);
xnor UO_1131 (O_1131,N_23933,N_21702);
nand UO_1132 (O_1132,N_23445,N_21236);
nor UO_1133 (O_1133,N_21292,N_20342);
nand UO_1134 (O_1134,N_24312,N_20444);
and UO_1135 (O_1135,N_21735,N_22809);
nor UO_1136 (O_1136,N_23312,N_21242);
nand UO_1137 (O_1137,N_20975,N_21643);
xnor UO_1138 (O_1138,N_23253,N_24342);
or UO_1139 (O_1139,N_22800,N_21794);
nand UO_1140 (O_1140,N_23137,N_22359);
and UO_1141 (O_1141,N_21742,N_22136);
or UO_1142 (O_1142,N_23712,N_23741);
nor UO_1143 (O_1143,N_22649,N_23584);
and UO_1144 (O_1144,N_24171,N_20570);
or UO_1145 (O_1145,N_24897,N_24646);
and UO_1146 (O_1146,N_23473,N_22388);
and UO_1147 (O_1147,N_20533,N_23015);
and UO_1148 (O_1148,N_24261,N_22979);
nand UO_1149 (O_1149,N_24047,N_22417);
and UO_1150 (O_1150,N_22905,N_22001);
and UO_1151 (O_1151,N_20748,N_20772);
nor UO_1152 (O_1152,N_24058,N_23520);
and UO_1153 (O_1153,N_22795,N_21271);
nand UO_1154 (O_1154,N_24402,N_23889);
and UO_1155 (O_1155,N_22588,N_22876);
nor UO_1156 (O_1156,N_21949,N_22525);
or UO_1157 (O_1157,N_21346,N_22000);
and UO_1158 (O_1158,N_23544,N_22373);
nand UO_1159 (O_1159,N_20099,N_23752);
and UO_1160 (O_1160,N_23130,N_22421);
nand UO_1161 (O_1161,N_21384,N_22749);
nand UO_1162 (O_1162,N_20968,N_21799);
or UO_1163 (O_1163,N_23616,N_22798);
nor UO_1164 (O_1164,N_23660,N_20057);
nor UO_1165 (O_1165,N_22088,N_23361);
nor UO_1166 (O_1166,N_24474,N_20947);
and UO_1167 (O_1167,N_22792,N_21828);
or UO_1168 (O_1168,N_20376,N_24480);
and UO_1169 (O_1169,N_24772,N_24629);
nor UO_1170 (O_1170,N_20736,N_24303);
and UO_1171 (O_1171,N_24280,N_24676);
nor UO_1172 (O_1172,N_20069,N_22497);
and UO_1173 (O_1173,N_20153,N_23119);
or UO_1174 (O_1174,N_23125,N_24429);
and UO_1175 (O_1175,N_24928,N_20104);
xnor UO_1176 (O_1176,N_23455,N_22760);
nor UO_1177 (O_1177,N_22058,N_20906);
nor UO_1178 (O_1178,N_24885,N_21113);
nor UO_1179 (O_1179,N_23760,N_21112);
nor UO_1180 (O_1180,N_20197,N_21822);
xor UO_1181 (O_1181,N_20073,N_24074);
or UO_1182 (O_1182,N_24453,N_23708);
nor UO_1183 (O_1183,N_23082,N_23267);
or UO_1184 (O_1184,N_22046,N_24296);
nor UO_1185 (O_1185,N_22292,N_21624);
and UO_1186 (O_1186,N_24203,N_21418);
and UO_1187 (O_1187,N_23646,N_22055);
and UO_1188 (O_1188,N_24126,N_21148);
nand UO_1189 (O_1189,N_21901,N_22514);
xnor UO_1190 (O_1190,N_23259,N_24322);
nand UO_1191 (O_1191,N_20229,N_22233);
nor UO_1192 (O_1192,N_23560,N_24052);
and UO_1193 (O_1193,N_22601,N_21954);
and UO_1194 (O_1194,N_20571,N_22767);
or UO_1195 (O_1195,N_24204,N_23229);
or UO_1196 (O_1196,N_22352,N_22745);
and UO_1197 (O_1197,N_23021,N_20955);
nor UO_1198 (O_1198,N_23494,N_24424);
nand UO_1199 (O_1199,N_22274,N_20506);
nor UO_1200 (O_1200,N_22671,N_21476);
nor UO_1201 (O_1201,N_23846,N_21524);
or UO_1202 (O_1202,N_24276,N_22053);
nand UO_1203 (O_1203,N_21454,N_22149);
nand UO_1204 (O_1204,N_23859,N_23513);
or UO_1205 (O_1205,N_22351,N_21724);
nand UO_1206 (O_1206,N_23337,N_24165);
and UO_1207 (O_1207,N_24118,N_20952);
nand UO_1208 (O_1208,N_23706,N_24169);
and UO_1209 (O_1209,N_23185,N_20877);
and UO_1210 (O_1210,N_24016,N_24104);
and UO_1211 (O_1211,N_22056,N_24245);
or UO_1212 (O_1212,N_20267,N_24384);
nor UO_1213 (O_1213,N_20710,N_23251);
and UO_1214 (O_1214,N_22900,N_24740);
or UO_1215 (O_1215,N_24673,N_20508);
nor UO_1216 (O_1216,N_20542,N_21051);
nand UO_1217 (O_1217,N_20301,N_20454);
and UO_1218 (O_1218,N_24460,N_23722);
nor UO_1219 (O_1219,N_22327,N_24055);
or UO_1220 (O_1220,N_21987,N_24501);
or UO_1221 (O_1221,N_20240,N_20108);
nor UO_1222 (O_1222,N_20228,N_21367);
and UO_1223 (O_1223,N_22672,N_21141);
nand UO_1224 (O_1224,N_24158,N_22537);
nand UO_1225 (O_1225,N_22361,N_24790);
and UO_1226 (O_1226,N_20690,N_20681);
nor UO_1227 (O_1227,N_21819,N_21919);
or UO_1228 (O_1228,N_21502,N_22614);
or UO_1229 (O_1229,N_20513,N_22769);
nor UO_1230 (O_1230,N_20485,N_21842);
or UO_1231 (O_1231,N_20703,N_24529);
nand UO_1232 (O_1232,N_23786,N_22408);
nor UO_1233 (O_1233,N_20782,N_22731);
nor UO_1234 (O_1234,N_21009,N_24720);
or UO_1235 (O_1235,N_23556,N_22063);
nor UO_1236 (O_1236,N_22031,N_22273);
nor UO_1237 (O_1237,N_24146,N_21830);
nand UO_1238 (O_1238,N_20394,N_22316);
nor UO_1239 (O_1239,N_21518,N_24985);
or UO_1240 (O_1240,N_21753,N_23195);
nand UO_1241 (O_1241,N_20019,N_22341);
or UO_1242 (O_1242,N_23800,N_24241);
and UO_1243 (O_1243,N_21195,N_23910);
and UO_1244 (O_1244,N_21573,N_23866);
or UO_1245 (O_1245,N_20163,N_20519);
nand UO_1246 (O_1246,N_20308,N_23816);
nor UO_1247 (O_1247,N_21940,N_21441);
or UO_1248 (O_1248,N_20751,N_24232);
nand UO_1249 (O_1249,N_23381,N_20330);
and UO_1250 (O_1250,N_23721,N_20127);
or UO_1251 (O_1251,N_23550,N_23700);
or UO_1252 (O_1252,N_22834,N_22038);
nor UO_1253 (O_1253,N_24244,N_21128);
nor UO_1254 (O_1254,N_21389,N_20453);
nor UO_1255 (O_1255,N_22732,N_24013);
or UO_1256 (O_1256,N_20094,N_23993);
and UO_1257 (O_1257,N_24700,N_22591);
and UO_1258 (O_1258,N_23459,N_21299);
or UO_1259 (O_1259,N_21657,N_21955);
nor UO_1260 (O_1260,N_20176,N_20693);
nor UO_1261 (O_1261,N_21523,N_24345);
or UO_1262 (O_1262,N_20309,N_22720);
nor UO_1263 (O_1263,N_22363,N_23402);
nand UO_1264 (O_1264,N_21202,N_20218);
nor UO_1265 (O_1265,N_20277,N_22655);
xor UO_1266 (O_1266,N_23463,N_21898);
xnor UO_1267 (O_1267,N_20416,N_23960);
nor UO_1268 (O_1268,N_23511,N_21478);
and UO_1269 (O_1269,N_21993,N_23030);
or UO_1270 (O_1270,N_20999,N_23012);
nand UO_1271 (O_1271,N_21604,N_21590);
nor UO_1272 (O_1272,N_23659,N_23908);
nand UO_1273 (O_1273,N_24470,N_23895);
nor UO_1274 (O_1274,N_20362,N_21880);
or UO_1275 (O_1275,N_22141,N_22188);
xnor UO_1276 (O_1276,N_21994,N_20624);
and UO_1277 (O_1277,N_20894,N_22028);
nand UO_1278 (O_1278,N_20402,N_21784);
nand UO_1279 (O_1279,N_23036,N_24398);
or UO_1280 (O_1280,N_20425,N_20532);
and UO_1281 (O_1281,N_23041,N_23310);
nor UO_1282 (O_1282,N_21370,N_22801);
and UO_1283 (O_1283,N_21553,N_22995);
and UO_1284 (O_1284,N_21816,N_23894);
nand UO_1285 (O_1285,N_22075,N_21945);
and UO_1286 (O_1286,N_24039,N_24908);
and UO_1287 (O_1287,N_21110,N_20451);
xnor UO_1288 (O_1288,N_21071,N_24493);
nand UO_1289 (O_1289,N_24721,N_24482);
and UO_1290 (O_1290,N_23197,N_22353);
nand UO_1291 (O_1291,N_23558,N_23486);
nor UO_1292 (O_1292,N_24421,N_24129);
or UO_1293 (O_1293,N_21598,N_23108);
and UO_1294 (O_1294,N_20996,N_22772);
and UO_1295 (O_1295,N_20151,N_22239);
nor UO_1296 (O_1296,N_22216,N_24137);
or UO_1297 (O_1297,N_24351,N_23619);
and UO_1298 (O_1298,N_22881,N_22626);
and UO_1299 (O_1299,N_23723,N_23075);
or UO_1300 (O_1300,N_23591,N_21087);
nor UO_1301 (O_1301,N_22592,N_23079);
nor UO_1302 (O_1302,N_22305,N_20258);
or UO_1303 (O_1303,N_23880,N_24625);
nor UO_1304 (O_1304,N_24164,N_21436);
nand UO_1305 (O_1305,N_20559,N_23407);
nor UO_1306 (O_1306,N_23078,N_21615);
and UO_1307 (O_1307,N_22642,N_22836);
and UO_1308 (O_1308,N_22203,N_22099);
nand UO_1309 (O_1309,N_22780,N_20800);
and UO_1310 (O_1310,N_21183,N_21863);
nand UO_1311 (O_1311,N_22952,N_20027);
and UO_1312 (O_1312,N_21672,N_24906);
and UO_1313 (O_1313,N_23881,N_23471);
xnor UO_1314 (O_1314,N_21275,N_20442);
nor UO_1315 (O_1315,N_22590,N_20160);
or UO_1316 (O_1316,N_23287,N_21916);
and UO_1317 (O_1317,N_22951,N_23938);
nor UO_1318 (O_1318,N_24389,N_24100);
nand UO_1319 (O_1319,N_23177,N_23007);
or UO_1320 (O_1320,N_23840,N_22119);
or UO_1321 (O_1321,N_24353,N_22160);
nor UO_1322 (O_1322,N_24412,N_22147);
nor UO_1323 (O_1323,N_24995,N_21134);
and UO_1324 (O_1324,N_24109,N_20904);
nand UO_1325 (O_1325,N_24613,N_22912);
nand UO_1326 (O_1326,N_23734,N_21625);
nor UO_1327 (O_1327,N_23649,N_24396);
nand UO_1328 (O_1328,N_20658,N_24422);
nand UO_1329 (O_1329,N_21890,N_24302);
and UO_1330 (O_1330,N_23331,N_22665);
nor UO_1331 (O_1331,N_21039,N_21423);
nor UO_1332 (O_1332,N_22054,N_22835);
nand UO_1333 (O_1333,N_20152,N_22258);
or UO_1334 (O_1334,N_22646,N_24733);
nor UO_1335 (O_1335,N_22661,N_23844);
nand UO_1336 (O_1336,N_23002,N_21714);
or UO_1337 (O_1337,N_20349,N_21064);
and UO_1338 (O_1338,N_21869,N_21433);
nor UO_1339 (O_1339,N_23142,N_21721);
and UO_1340 (O_1340,N_24719,N_23825);
or UO_1341 (O_1341,N_23753,N_24749);
nand UO_1342 (O_1342,N_21530,N_24889);
or UO_1343 (O_1343,N_21427,N_23291);
or UO_1344 (O_1344,N_20467,N_22520);
or UO_1345 (O_1345,N_22882,N_23426);
and UO_1346 (O_1346,N_21956,N_24086);
or UO_1347 (O_1347,N_20115,N_24329);
nor UO_1348 (O_1348,N_20920,N_20648);
and UO_1349 (O_1349,N_23769,N_20529);
or UO_1350 (O_1350,N_22733,N_21539);
and UO_1351 (O_1351,N_23416,N_22991);
and UO_1352 (O_1352,N_21274,N_22983);
xnor UO_1353 (O_1353,N_20045,N_21705);
and UO_1354 (O_1354,N_23968,N_21675);
nand UO_1355 (O_1355,N_22125,N_21846);
nand UO_1356 (O_1356,N_20931,N_23761);
nand UO_1357 (O_1357,N_21489,N_20666);
or UO_1358 (O_1358,N_21453,N_24053);
nor UO_1359 (O_1359,N_21220,N_22777);
nand UO_1360 (O_1360,N_22430,N_21608);
nand UO_1361 (O_1361,N_23441,N_24935);
or UO_1362 (O_1362,N_24663,N_23841);
or UO_1363 (O_1363,N_21996,N_20561);
and UO_1364 (O_1364,N_22803,N_23069);
nor UO_1365 (O_1365,N_24461,N_22076);
nor UO_1366 (O_1366,N_20816,N_22011);
or UO_1367 (O_1367,N_24407,N_22965);
and UO_1368 (O_1368,N_23923,N_24192);
and UO_1369 (O_1369,N_21567,N_24105);
nand UO_1370 (O_1370,N_21853,N_22177);
nand UO_1371 (O_1371,N_22677,N_21935);
nand UO_1372 (O_1372,N_23523,N_21849);
nor UO_1373 (O_1373,N_23852,N_23357);
nand UO_1374 (O_1374,N_24575,N_24119);
and UO_1375 (O_1375,N_24934,N_24250);
or UO_1376 (O_1376,N_23955,N_22923);
xor UO_1377 (O_1377,N_23000,N_22499);
and UO_1378 (O_1378,N_23847,N_24887);
nor UO_1379 (O_1379,N_22484,N_24836);
nand UO_1380 (O_1380,N_23665,N_20319);
or UO_1381 (O_1381,N_24527,N_24021);
and UO_1382 (O_1382,N_23689,N_23170);
or UO_1383 (O_1383,N_22997,N_24655);
nand UO_1384 (O_1384,N_22334,N_22128);
nand UO_1385 (O_1385,N_20780,N_23117);
nor UO_1386 (O_1386,N_20379,N_22311);
or UO_1387 (O_1387,N_24777,N_20988);
nor UO_1388 (O_1388,N_23802,N_22629);
nor UO_1389 (O_1389,N_24586,N_20441);
nor UO_1390 (O_1390,N_21832,N_23072);
nand UO_1391 (O_1391,N_22377,N_23989);
nor UO_1392 (O_1392,N_24666,N_22533);
nand UO_1393 (O_1393,N_23971,N_24680);
and UO_1394 (O_1394,N_21700,N_24368);
nand UO_1395 (O_1395,N_20148,N_21482);
or UO_1396 (O_1396,N_20911,N_21061);
nand UO_1397 (O_1397,N_24746,N_22067);
and UO_1398 (O_1398,N_23397,N_20364);
or UO_1399 (O_1399,N_21642,N_23332);
and UO_1400 (O_1400,N_22691,N_21069);
nor UO_1401 (O_1401,N_23624,N_20970);
nor UO_1402 (O_1402,N_21434,N_21762);
nor UO_1403 (O_1403,N_24954,N_23555);
and UO_1404 (O_1404,N_22175,N_21912);
or UO_1405 (O_1405,N_21718,N_23209);
nand UO_1406 (O_1406,N_23038,N_24849);
nand UO_1407 (O_1407,N_21575,N_23551);
and UO_1408 (O_1408,N_22207,N_24757);
nand UO_1409 (O_1409,N_24227,N_23515);
or UO_1410 (O_1410,N_20496,N_24548);
nand UO_1411 (O_1411,N_23201,N_23224);
or UO_1412 (O_1412,N_20031,N_24847);
and UO_1413 (O_1413,N_23739,N_22549);
and UO_1414 (O_1414,N_23161,N_21473);
nand UO_1415 (O_1415,N_21177,N_20516);
nor UO_1416 (O_1416,N_22816,N_22724);
nand UO_1417 (O_1417,N_20261,N_20787);
and UO_1418 (O_1418,N_21378,N_21421);
and UO_1419 (O_1419,N_22050,N_24043);
or UO_1420 (O_1420,N_20256,N_20448);
nand UO_1421 (O_1421,N_22133,N_20929);
or UO_1422 (O_1422,N_20938,N_22086);
and UO_1423 (O_1423,N_21040,N_24555);
nor UO_1424 (O_1424,N_24609,N_23930);
nor UO_1425 (O_1425,N_23714,N_21969);
xor UO_1426 (O_1426,N_22717,N_21328);
and UO_1427 (O_1427,N_24128,N_20391);
nand UO_1428 (O_1428,N_23024,N_21736);
or UO_1429 (O_1429,N_20644,N_23202);
or UO_1430 (O_1430,N_24321,N_22113);
or UO_1431 (O_1431,N_21871,N_21549);
nor UO_1432 (O_1432,N_20969,N_21008);
nand UO_1433 (O_1433,N_23783,N_22906);
and UO_1434 (O_1434,N_24114,N_24994);
or UO_1435 (O_1435,N_22228,N_24247);
nor UO_1436 (O_1436,N_24451,N_21430);
nand UO_1437 (O_1437,N_22734,N_22635);
or UO_1438 (O_1438,N_24997,N_20543);
nor UO_1439 (O_1439,N_23408,N_23183);
nand UO_1440 (O_1440,N_24949,N_23068);
or UO_1441 (O_1441,N_21268,N_20323);
nand UO_1442 (O_1442,N_24005,N_24183);
and UO_1443 (O_1443,N_24905,N_24649);
or UO_1444 (O_1444,N_21512,N_24464);
or UO_1445 (O_1445,N_22532,N_21786);
nor UO_1446 (O_1446,N_24552,N_20174);
nor UO_1447 (O_1447,N_20674,N_22893);
or UO_1448 (O_1448,N_24269,N_23737);
and UO_1449 (O_1449,N_20368,N_24601);
nand UO_1450 (O_1450,N_20742,N_21191);
nor UO_1451 (O_1451,N_21782,N_20873);
nand UO_1452 (O_1452,N_20881,N_23386);
and UO_1453 (O_1453,N_21789,N_24238);
nor UO_1454 (O_1454,N_24942,N_22023);
nor UO_1455 (O_1455,N_24338,N_21255);
or UO_1456 (O_1456,N_22637,N_22729);
and UO_1457 (O_1457,N_23327,N_24716);
or UO_1458 (O_1458,N_21803,N_20123);
and UO_1459 (O_1459,N_24465,N_21481);
nor UO_1460 (O_1460,N_21895,N_22624);
and UO_1461 (O_1461,N_24714,N_24226);
or UO_1462 (O_1462,N_21500,N_20082);
nand UO_1463 (O_1463,N_23207,N_24331);
or UO_1464 (O_1464,N_21333,N_23100);
or UO_1465 (O_1465,N_22862,N_24606);
nand UO_1466 (O_1466,N_22030,N_21447);
nor UO_1467 (O_1467,N_22562,N_24925);
nor UO_1468 (O_1468,N_21915,N_21733);
nor UO_1469 (O_1469,N_23838,N_21538);
nand UO_1470 (O_1470,N_24362,N_23077);
and UO_1471 (O_1471,N_20603,N_23743);
and UO_1472 (O_1472,N_24441,N_21991);
nor UO_1473 (O_1473,N_20307,N_24308);
or UO_1474 (O_1474,N_24839,N_22478);
xor UO_1475 (O_1475,N_23063,N_24660);
and UO_1476 (O_1476,N_24747,N_24263);
or UO_1477 (O_1477,N_23986,N_23888);
nand UO_1478 (O_1478,N_20524,N_22963);
and UO_1479 (O_1479,N_21906,N_21386);
and UO_1480 (O_1480,N_23430,N_23663);
or UO_1481 (O_1481,N_22948,N_24223);
and UO_1482 (O_1482,N_22185,N_22959);
or UO_1483 (O_1483,N_20634,N_24933);
and UO_1484 (O_1484,N_24534,N_23860);
nor UO_1485 (O_1485,N_20347,N_22821);
or UO_1486 (O_1486,N_24375,N_24590);
nor UO_1487 (O_1487,N_24558,N_23051);
and UO_1488 (O_1488,N_21357,N_20895);
nand UO_1489 (O_1489,N_24025,N_20119);
nand UO_1490 (O_1490,N_23576,N_23343);
nand UO_1491 (O_1491,N_20588,N_21765);
and UO_1492 (O_1492,N_23071,N_22346);
and UO_1493 (O_1493,N_20278,N_23476);
nor UO_1494 (O_1494,N_22083,N_20597);
nor UO_1495 (O_1495,N_21696,N_23785);
and UO_1496 (O_1496,N_23272,N_22435);
nor UO_1497 (O_1497,N_24782,N_21360);
nor UO_1498 (O_1498,N_24071,N_20384);
nor UO_1499 (O_1499,N_24405,N_23255);
nor UO_1500 (O_1500,N_21187,N_24354);
nand UO_1501 (O_1501,N_21092,N_22398);
nand UO_1502 (O_1502,N_22121,N_23961);
or UO_1503 (O_1503,N_24007,N_23405);
nand UO_1504 (O_1504,N_23322,N_24009);
and UO_1505 (O_1505,N_20759,N_20255);
or UO_1506 (O_1506,N_21288,N_23845);
or UO_1507 (O_1507,N_21266,N_24325);
xor UO_1508 (O_1508,N_20121,N_22300);
nor UO_1509 (O_1509,N_21772,N_20557);
or UO_1510 (O_1510,N_20180,N_23157);
nand UO_1511 (O_1511,N_24502,N_21301);
nand UO_1512 (O_1512,N_21648,N_21888);
or UO_1513 (O_1513,N_22885,N_24282);
nand UO_1514 (O_1514,N_20288,N_21868);
nor UO_1515 (O_1515,N_22884,N_22955);
nor UO_1516 (O_1516,N_23962,N_22157);
and UO_1517 (O_1517,N_22739,N_22409);
nand UO_1518 (O_1518,N_20335,N_22823);
xnor UO_1519 (O_1519,N_23293,N_22197);
and UO_1520 (O_1520,N_23666,N_20026);
and UO_1521 (O_1521,N_20037,N_23223);
or UO_1522 (O_1522,N_21651,N_20655);
and UO_1523 (O_1523,N_20282,N_20711);
nand UO_1524 (O_1524,N_24500,N_20732);
and UO_1525 (O_1525,N_20024,N_21317);
nor UO_1526 (O_1526,N_23676,N_22526);
or UO_1527 (O_1527,N_21323,N_22797);
and UO_1528 (O_1528,N_24817,N_24166);
nor UO_1529 (O_1529,N_23797,N_22638);
or UO_1530 (O_1530,N_22947,N_21586);
nand UO_1531 (O_1531,N_22639,N_21876);
xor UO_1532 (O_1532,N_21603,N_22459);
and UO_1533 (O_1533,N_20054,N_22360);
nand UO_1534 (O_1534,N_23941,N_20865);
nand UO_1535 (O_1535,N_21247,N_24819);
and UO_1536 (O_1536,N_23153,N_21899);
nor UO_1537 (O_1537,N_24439,N_21764);
or UO_1538 (O_1538,N_24726,N_24271);
and UO_1539 (O_1539,N_21245,N_22344);
and UO_1540 (O_1540,N_24256,N_24587);
or UO_1541 (O_1541,N_20136,N_24872);
and UO_1542 (O_1542,N_20617,N_21658);
and UO_1543 (O_1543,N_24669,N_20535);
and UO_1544 (O_1544,N_23526,N_23315);
and UO_1545 (O_1545,N_24610,N_22405);
nand UO_1546 (O_1546,N_22096,N_22750);
and UO_1547 (O_1547,N_24806,N_22966);
nand UO_1548 (O_1548,N_21465,N_23102);
and UO_1549 (O_1549,N_22281,N_24565);
nor UO_1550 (O_1550,N_22084,N_21893);
nand UO_1551 (O_1551,N_20528,N_23035);
nand UO_1552 (O_1552,N_22770,N_20244);
nor UO_1553 (O_1553,N_22419,N_20326);
and UO_1554 (O_1554,N_22379,N_20670);
nand UO_1555 (O_1555,N_24301,N_22710);
and UO_1556 (O_1556,N_20941,N_24630);
nor UO_1557 (O_1557,N_24770,N_24200);
nand UO_1558 (O_1558,N_24023,N_23091);
and UO_1559 (O_1559,N_22509,N_22705);
and UO_1560 (O_1560,N_21670,N_22148);
or UO_1561 (O_1561,N_20531,N_24963);
or UO_1562 (O_1562,N_22132,N_24939);
nand UO_1563 (O_1563,N_22395,N_21748);
or UO_1564 (O_1564,N_23039,N_23081);
nor UO_1565 (O_1565,N_22813,N_22566);
or UO_1566 (O_1566,N_21686,N_23905);
or UO_1567 (O_1567,N_21133,N_22015);
and UO_1568 (O_1568,N_22986,N_22908);
nor UO_1569 (O_1569,N_20611,N_21779);
or UO_1570 (O_1570,N_22427,N_24913);
or UO_1571 (O_1571,N_20986,N_21100);
or UO_1572 (O_1572,N_20696,N_23884);
nand UO_1573 (O_1573,N_23799,N_23181);
nand UO_1574 (O_1574,N_21536,N_23491);
nand UO_1575 (O_1575,N_20465,N_23674);
nor UO_1576 (O_1576,N_21595,N_23928);
or UO_1577 (O_1577,N_24957,N_22180);
or UO_1578 (O_1578,N_22868,N_23258);
nor UO_1579 (O_1579,N_21942,N_24378);
nand UO_1580 (O_1580,N_22505,N_22314);
or UO_1581 (O_1581,N_20348,N_21532);
nor UO_1582 (O_1582,N_23174,N_24799);
or UO_1583 (O_1583,N_20382,N_23820);
or UO_1584 (O_1584,N_21961,N_22126);
nand UO_1585 (O_1585,N_22848,N_23475);
nor UO_1586 (O_1586,N_20235,N_20618);
nor UO_1587 (O_1587,N_20660,N_20847);
nor UO_1588 (O_1588,N_22616,N_22433);
nand UO_1589 (O_1589,N_21971,N_21337);
and UO_1590 (O_1590,N_22989,N_24127);
or UO_1591 (O_1591,N_21214,N_24420);
nand UO_1592 (O_1592,N_22669,N_23451);
or UO_1593 (O_1593,N_24334,N_24968);
or UO_1594 (O_1594,N_20337,N_24641);
or UO_1595 (O_1595,N_23468,N_20214);
nor UO_1596 (O_1596,N_21027,N_20105);
nor UO_1597 (O_1597,N_24691,N_24194);
nand UO_1598 (O_1598,N_22787,N_21807);
and UO_1599 (O_1599,N_21209,N_21683);
nand UO_1600 (O_1600,N_23419,N_23630);
nand UO_1601 (O_1601,N_23583,N_21529);
or UO_1602 (O_1602,N_20856,N_23085);
and UO_1603 (O_1603,N_22548,N_22322);
nand UO_1604 (O_1604,N_21181,N_20664);
nand UO_1605 (O_1605,N_21010,N_21474);
and UO_1606 (O_1606,N_21088,N_24674);
or UO_1607 (O_1607,N_22326,N_22268);
nand UO_1608 (O_1608,N_21924,N_24181);
nor UO_1609 (O_1609,N_24340,N_20113);
nor UO_1610 (O_1610,N_24620,N_23338);
and UO_1611 (O_1611,N_23375,N_21704);
or UO_1612 (O_1612,N_24410,N_23651);
or UO_1613 (O_1613,N_22425,N_23336);
nor UO_1614 (O_1614,N_24923,N_20090);
nor UO_1615 (O_1615,N_24360,N_20908);
nand UO_1616 (O_1616,N_20274,N_20709);
nor UO_1617 (O_1617,N_21793,N_24248);
or UO_1618 (O_1618,N_23673,N_20483);
and UO_1619 (O_1619,N_20619,N_24416);
nor UO_1620 (O_1620,N_21304,N_20399);
or UO_1621 (O_1621,N_23818,N_23121);
nand UO_1622 (O_1622,N_20808,N_22911);
or UO_1623 (O_1623,N_21685,N_21175);
and UO_1624 (O_1624,N_20289,N_22700);
or UO_1625 (O_1625,N_22077,N_20984);
nor UO_1626 (O_1626,N_20901,N_20333);
and UO_1627 (O_1627,N_20213,N_21080);
nand UO_1628 (O_1628,N_22400,N_23604);
or UO_1629 (O_1629,N_22319,N_21439);
nand UO_1630 (O_1630,N_24447,N_24433);
or UO_1631 (O_1631,N_24186,N_24517);
nand UO_1632 (O_1632,N_20978,N_20625);
nand UO_1633 (O_1633,N_21865,N_24249);
nand UO_1634 (O_1634,N_23861,N_22714);
nor UO_1635 (O_1635,N_20612,N_21810);
nand UO_1636 (O_1636,N_21213,N_22173);
nor UO_1637 (O_1637,N_22082,N_23919);
or UO_1638 (O_1638,N_20555,N_20085);
and UO_1639 (O_1639,N_23436,N_20435);
or UO_1640 (O_1640,N_23005,N_20177);
and UO_1641 (O_1641,N_23282,N_20697);
nand UO_1642 (O_1642,N_21564,N_23821);
and UO_1643 (O_1643,N_20501,N_20072);
or UO_1644 (O_1644,N_22302,N_23242);
nor UO_1645 (O_1645,N_20948,N_21937);
or UO_1646 (O_1646,N_24221,N_20239);
nor UO_1647 (O_1647,N_23055,N_24476);
or UO_1648 (O_1648,N_22224,N_24240);
and UO_1649 (O_1649,N_24686,N_24286);
and UO_1650 (O_1650,N_22291,N_22555);
nand UO_1651 (O_1651,N_22890,N_24159);
and UO_1652 (O_1652,N_23796,N_20470);
nand UO_1653 (O_1653,N_23061,N_20398);
nor UO_1654 (O_1654,N_24618,N_22044);
nand UO_1655 (O_1655,N_23828,N_24960);
nor UO_1656 (O_1656,N_20831,N_20011);
and UO_1657 (O_1657,N_22248,N_21126);
nand UO_1658 (O_1658,N_24598,N_21668);
xor UO_1659 (O_1659,N_21834,N_24564);
and UO_1660 (O_1660,N_22647,N_21225);
nand UO_1661 (O_1661,N_22619,N_23680);
and UO_1662 (O_1662,N_21410,N_20884);
and UO_1663 (O_1663,N_21269,N_20643);
or UO_1664 (O_1664,N_22443,N_22569);
nand UO_1665 (O_1665,N_24254,N_22007);
and UO_1666 (O_1666,N_24229,N_23534);
nor UO_1667 (O_1667,N_23897,N_20210);
or UO_1668 (O_1668,N_21560,N_20909);
nand UO_1669 (O_1669,N_21239,N_20705);
and UO_1670 (O_1670,N_21706,N_23234);
nand UO_1671 (O_1671,N_20458,N_24444);
and UO_1672 (O_1672,N_21178,N_20896);
or UO_1673 (O_1673,N_20429,N_24341);
nor UO_1674 (O_1674,N_23969,N_22237);
and UO_1675 (O_1675,N_22855,N_20265);
nor UO_1676 (O_1676,N_23936,N_20595);
nand UO_1677 (O_1677,N_24581,N_20087);
or UO_1678 (O_1678,N_23592,N_20731);
or UO_1679 (O_1679,N_22718,N_20899);
and UO_1680 (O_1680,N_22888,N_20610);
nor UO_1681 (O_1681,N_21981,N_20263);
nand UO_1682 (O_1682,N_23790,N_23695);
or UO_1683 (O_1683,N_23618,N_21831);
or UO_1684 (O_1684,N_22581,N_24463);
nand UO_1685 (O_1685,N_20088,N_20825);
nor UO_1686 (O_1686,N_22869,N_22401);
nor UO_1687 (O_1687,N_24393,N_21728);
nand UO_1688 (O_1688,N_24547,N_20566);
nand UO_1689 (O_1689,N_22323,N_23347);
nand UO_1690 (O_1690,N_20397,N_24753);
nand UO_1691 (O_1691,N_20351,N_21287);
or UO_1692 (O_1692,N_23974,N_22576);
and UO_1693 (O_1693,N_20427,N_24498);
nor UO_1694 (O_1694,N_21234,N_21626);
and UO_1695 (O_1695,N_24051,N_22178);
or UO_1696 (O_1696,N_21503,N_23237);
or UO_1697 (O_1697,N_21802,N_21475);
nor UO_1698 (O_1698,N_22226,N_20853);
nor UO_1699 (O_1699,N_21235,N_23939);
nand UO_1700 (O_1700,N_23798,N_20995);
and UO_1701 (O_1701,N_21249,N_21494);
nand UO_1702 (O_1702,N_23008,N_23472);
and UO_1703 (O_1703,N_23232,N_23020);
and UO_1704 (O_1704,N_24881,N_22184);
nand UO_1705 (O_1705,N_20056,N_23598);
nor UO_1706 (O_1706,N_24865,N_21962);
and UO_1707 (O_1707,N_22285,N_24662);
and UO_1708 (O_1708,N_20667,N_22265);
or UO_1709 (O_1709,N_21058,N_20331);
nand UO_1710 (O_1710,N_21632,N_22250);
and UO_1711 (O_1711,N_21144,N_24056);
or UO_1712 (O_1712,N_22168,N_23165);
nand UO_1713 (O_1713,N_23518,N_24634);
nor UO_1714 (O_1714,N_21158,N_23758);
nor UO_1715 (O_1715,N_21811,N_21698);
nor UO_1716 (O_1716,N_24532,N_21238);
nand UO_1717 (O_1717,N_21218,N_21989);
nor UO_1718 (O_1718,N_23872,N_22894);
nor UO_1719 (O_1719,N_22850,N_24741);
and UO_1720 (O_1720,N_23394,N_21018);
or UO_1721 (O_1721,N_23457,N_20641);
xor UO_1722 (O_1722,N_24752,N_20905);
nor UO_1723 (O_1723,N_24535,N_22437);
nand UO_1724 (O_1724,N_22879,N_24760);
xor UO_1725 (O_1725,N_22399,N_23140);
and UO_1726 (O_1726,N_21958,N_23176);
or UO_1727 (O_1727,N_24504,N_23248);
nand UO_1728 (O_1728,N_24195,N_24917);
or UO_1729 (O_1729,N_24635,N_24026);
nand UO_1730 (O_1730,N_20987,N_21396);
and UO_1731 (O_1731,N_23699,N_21664);
and UO_1732 (O_1732,N_22737,N_24736);
nand UO_1733 (O_1733,N_21032,N_21260);
nor UO_1734 (O_1734,N_22074,N_24701);
nand UO_1735 (O_1735,N_21349,N_20098);
nand UO_1736 (O_1736,N_20272,N_20205);
or UO_1737 (O_1737,N_23245,N_22958);
and UO_1738 (O_1738,N_20184,N_23603);
nand UO_1739 (O_1739,N_23429,N_22458);
or UO_1740 (O_1740,N_21995,N_23478);
nand UO_1741 (O_1741,N_24712,N_22577);
or UO_1742 (O_1742,N_23042,N_21903);
nand UO_1743 (O_1743,N_23742,N_22527);
nand UO_1744 (O_1744,N_24870,N_20092);
xor UO_1745 (O_1745,N_22764,N_24626);
xor UO_1746 (O_1746,N_21467,N_22365);
nand UO_1747 (O_1747,N_23858,N_24154);
nor UO_1748 (O_1748,N_20251,N_24971);
and UO_1749 (O_1749,N_24975,N_22939);
and UO_1750 (O_1750,N_23693,N_24489);
or UO_1751 (O_1751,N_24274,N_21574);
nand UO_1752 (O_1752,N_24079,N_22198);
nand UO_1753 (O_1753,N_22563,N_20686);
and UO_1754 (O_1754,N_20324,N_21291);
or UO_1755 (O_1755,N_20063,N_22542);
or UO_1756 (O_1756,N_23427,N_24411);
nand UO_1757 (O_1757,N_23656,N_23439);
nand UO_1758 (O_1758,N_21231,N_22846);
or UO_1759 (O_1759,N_20756,N_20712);
nand UO_1760 (O_1760,N_21569,N_23589);
nor UO_1761 (O_1761,N_20111,N_23488);
or UO_1762 (O_1762,N_22135,N_22934);
or UO_1763 (O_1763,N_22104,N_22241);
or UO_1764 (O_1764,N_21034,N_21272);
nand UO_1765 (O_1765,N_22988,N_24521);
nor UO_1766 (O_1766,N_21024,N_23717);
nand UO_1767 (O_1767,N_24855,N_22587);
nand UO_1768 (O_1768,N_21805,N_20526);
and UO_1769 (O_1769,N_23793,N_24503);
and UO_1770 (O_1770,N_21194,N_22106);
or UO_1771 (O_1771,N_24163,N_22413);
or UO_1772 (O_1772,N_24170,N_22005);
or UO_1773 (O_1773,N_23172,N_24054);
and UO_1774 (O_1774,N_22871,N_21545);
nor UO_1775 (O_1775,N_23307,N_20738);
nand UO_1776 (O_1776,N_21754,N_24468);
or UO_1777 (O_1777,N_20497,N_24812);
or UO_1778 (O_1778,N_20216,N_23687);
nand UO_1779 (O_1779,N_23423,N_20439);
or UO_1780 (O_1780,N_23129,N_21377);
nor UO_1781 (O_1781,N_22738,N_21309);
nand UO_1782 (O_1782,N_22094,N_20133);
and UO_1783 (O_1783,N_20208,N_20359);
or UO_1784 (O_1784,N_22668,N_21168);
or UO_1785 (O_1785,N_20971,N_20424);
nand UO_1786 (O_1786,N_23731,N_21516);
and UO_1787 (O_1787,N_24902,N_22068);
or UO_1788 (O_1788,N_22695,N_21362);
and UO_1789 (O_1789,N_21884,N_22035);
nand UO_1790 (O_1790,N_20867,N_23355);
nor UO_1791 (O_1791,N_20204,N_23243);
or UO_1792 (O_1792,N_21081,N_24099);
nand UO_1793 (O_1793,N_22864,N_24173);
nand UO_1794 (O_1794,N_22903,N_21690);
nand UO_1795 (O_1795,N_21732,N_24180);
and UO_1796 (O_1796,N_20866,N_21923);
nand UO_1797 (O_1797,N_20830,N_22092);
nand UO_1798 (O_1798,N_23147,N_22439);
or UO_1799 (O_1799,N_24161,N_24408);
and UO_1800 (O_1800,N_22432,N_23912);
or UO_1801 (O_1801,N_20052,N_20797);
xnor UO_1802 (O_1802,N_21960,N_23466);
and UO_1803 (O_1803,N_22155,N_24713);
nor UO_1804 (O_1804,N_24190,N_20798);
nor UO_1805 (O_1805,N_21997,N_22004);
nand UO_1806 (O_1806,N_23787,N_21223);
nor UO_1807 (O_1807,N_21597,N_23738);
and UO_1808 (O_1808,N_23836,N_23730);
xor UO_1809 (O_1809,N_24943,N_20221);
or UO_1810 (O_1810,N_24311,N_24758);
and UO_1811 (O_1811,N_20317,N_20621);
nor UO_1812 (O_1812,N_21320,N_21911);
xnor UO_1813 (O_1813,N_22632,N_23615);
nand UO_1814 (O_1814,N_24309,N_22810);
or UO_1815 (O_1815,N_23190,N_22040);
and UO_1816 (O_1816,N_23597,N_21251);
nand UO_1817 (O_1817,N_24237,N_20401);
or UO_1818 (O_1818,N_20078,N_20270);
nor UO_1819 (O_1819,N_21315,N_24152);
nor UO_1820 (O_1820,N_20484,N_21568);
or UO_1821 (O_1821,N_22090,N_20841);
nor UO_1822 (O_1822,N_20586,N_24065);
xor UO_1823 (O_1823,N_23727,N_23593);
or UO_1824 (O_1824,N_20081,N_20066);
and UO_1825 (O_1825,N_22865,N_22517);
nor UO_1826 (O_1826,N_22589,N_24876);
and UO_1827 (O_1827,N_21917,N_21406);
nand UO_1828 (O_1828,N_22957,N_24576);
and UO_1829 (O_1829,N_23139,N_20937);
nand UO_1830 (O_1830,N_20047,N_22496);
nand UO_1831 (O_1831,N_22633,N_22045);
or UO_1832 (O_1832,N_23681,N_22098);
nor UO_1833 (O_1833,N_22552,N_20234);
or UO_1834 (O_1834,N_22396,N_23981);
and UO_1835 (O_1835,N_20336,N_21730);
nand UO_1836 (O_1836,N_23935,N_24823);
nor UO_1837 (O_1837,N_24370,N_20480);
nor UO_1838 (O_1838,N_21297,N_22711);
and UO_1839 (O_1839,N_23118,N_24283);
and UO_1840 (O_1840,N_22471,N_22596);
and UO_1841 (O_1841,N_23713,N_22238);
or UO_1842 (O_1842,N_20682,N_20990);
or UO_1843 (O_1843,N_20940,N_20455);
nor UO_1844 (O_1844,N_22466,N_24693);
or UO_1845 (O_1845,N_22630,N_21948);
xnor UO_1846 (O_1846,N_20186,N_21119);
or UO_1847 (O_1847,N_23150,N_20236);
nor UO_1848 (O_1848,N_22927,N_24734);
nand UO_1849 (O_1849,N_22827,N_23368);
nand UO_1850 (O_1850,N_21783,N_24022);
nand UO_1851 (O_1851,N_23596,N_21351);
nand UO_1852 (O_1852,N_23937,N_23725);
xnor UO_1853 (O_1853,N_23415,N_20724);
and UO_1854 (O_1854,N_21380,N_20837);
and UO_1855 (O_1855,N_23417,N_20743);
nor UO_1856 (O_1856,N_20553,N_20626);
or UO_1857 (O_1857,N_23605,N_20574);
and UO_1858 (O_1858,N_24012,N_22681);
xor UO_1859 (O_1859,N_20511,N_22006);
and UO_1860 (O_1860,N_22594,N_24769);
and UO_1861 (O_1861,N_20685,N_21432);
or UO_1862 (O_1862,N_20552,N_20869);
nor UO_1863 (O_1863,N_20584,N_24036);
nand UO_1864 (O_1864,N_21920,N_21452);
nor UO_1865 (O_1865,N_21515,N_23477);
and UO_1866 (O_1866,N_22867,N_22187);
and UO_1867 (O_1867,N_23553,N_24542);
and UO_1868 (O_1868,N_23667,N_20623);
or UO_1869 (O_1869,N_23350,N_20647);
nor UO_1870 (O_1870,N_24138,N_21673);
nand UO_1871 (O_1871,N_22556,N_23652);
nor UO_1872 (O_1872,N_23683,N_21114);
xor UO_1873 (O_1873,N_21677,N_22469);
nand UO_1874 (O_1874,N_22793,N_21118);
nor UO_1875 (O_1875,N_21681,N_24550);
or UO_1876 (O_1876,N_23582,N_24878);
and UO_1877 (O_1877,N_21533,N_22026);
and UO_1878 (O_1878,N_23540,N_20403);
nand UO_1879 (O_1879,N_22495,N_22872);
and UO_1880 (O_1880,N_23001,N_24224);
nand UO_1881 (O_1881,N_23054,N_20928);
or UO_1882 (O_1882,N_22313,N_23421);
or UO_1883 (O_1883,N_21402,N_24914);
nor UO_1884 (O_1884,N_24664,N_24139);
and UO_1885 (O_1885,N_21593,N_21111);
or UO_1886 (O_1886,N_24938,N_23602);
nand UO_1887 (O_1887,N_20018,N_21892);
nand UO_1888 (O_1888,N_22410,N_21833);
or UO_1889 (O_1889,N_23498,N_21459);
or UO_1890 (O_1890,N_23154,N_20845);
nand UO_1891 (O_1891,N_22568,N_23890);
nand UO_1892 (O_1892,N_24387,N_22570);
and UO_1893 (O_1893,N_24003,N_22463);
nor UO_1894 (O_1894,N_23444,N_20206);
xnor UO_1895 (O_1895,N_21227,N_20243);
or UO_1896 (O_1896,N_22706,N_24953);
or UO_1897 (O_1897,N_24583,N_21631);
or UO_1898 (O_1898,N_21864,N_23851);
nand UO_1899 (O_1899,N_21109,N_21013);
nor UO_1900 (O_1900,N_24571,N_22715);
nand UO_1901 (O_1901,N_20051,N_22874);
and UO_1902 (O_1902,N_20790,N_21038);
and UO_1903 (O_1903,N_20371,N_20520);
nor UO_1904 (O_1904,N_24267,N_24675);
xnor UO_1905 (O_1905,N_20071,N_22295);
nand UO_1906 (O_1906,N_21464,N_20549);
or UO_1907 (O_1907,N_21460,N_20195);
and UO_1908 (O_1908,N_20411,N_21156);
nor UO_1909 (O_1909,N_21030,N_22839);
or UO_1910 (O_1910,N_22531,N_21130);
and UO_1911 (O_1911,N_23275,N_23425);
nor UO_1912 (O_1912,N_20338,N_22773);
nand UO_1913 (O_1913,N_22586,N_22070);
nand UO_1914 (O_1914,N_21872,N_23032);
nand UO_1915 (O_1915,N_21487,N_21680);
nand UO_1916 (O_1916,N_23755,N_21769);
and UO_1917 (O_1917,N_24764,N_20273);
xor UO_1918 (O_1918,N_24822,N_21185);
or UO_1919 (O_1919,N_20242,N_23958);
and UO_1920 (O_1920,N_22037,N_21163);
nand UO_1921 (O_1921,N_23353,N_21329);
nand UO_1922 (O_1922,N_20046,N_23123);
nand UO_1923 (O_1923,N_22382,N_22191);
nor UO_1924 (O_1924,N_21221,N_21006);
nor UO_1925 (O_1925,N_22653,N_21497);
or UO_1926 (O_1926,N_20602,N_23045);
xnor UO_1927 (O_1927,N_24006,N_24069);
and UO_1928 (O_1928,N_24046,N_22414);
or UO_1929 (O_1929,N_20960,N_23803);
nor UO_1930 (O_1930,N_24840,N_23885);
nand UO_1931 (O_1931,N_21600,N_24385);
nor UO_1932 (O_1932,N_23679,N_23145);
or UO_1933 (O_1933,N_22060,N_21798);
or UO_1934 (O_1934,N_24567,N_21165);
and UO_1935 (O_1935,N_22454,N_23778);
and UO_1936 (O_1936,N_22468,N_20185);
nand UO_1937 (O_1937,N_23362,N_23062);
nand UO_1938 (O_1938,N_23504,N_21988);
and UO_1939 (O_1939,N_21612,N_24824);
nor UO_1940 (O_1940,N_24083,N_21900);
and UO_1941 (O_1941,N_24193,N_20730);
and UO_1942 (O_1942,N_22783,N_24297);
or UO_1943 (O_1943,N_24208,N_21627);
or UO_1944 (O_1944,N_20361,N_24454);
xor UO_1945 (O_1945,N_21151,N_22946);
or UO_1946 (O_1946,N_22039,N_20974);
nand UO_1947 (O_1947,N_21566,N_21104);
or UO_1948 (O_1948,N_21411,N_24556);
or UO_1949 (O_1949,N_23995,N_24251);
nand UO_1950 (O_1950,N_20933,N_24910);
and UO_1951 (O_1951,N_22603,N_23633);
nand UO_1952 (O_1952,N_20846,N_20769);
or UO_1953 (O_1953,N_23610,N_24228);
or UO_1954 (O_1954,N_22080,N_21096);
and UO_1955 (O_1955,N_22854,N_22100);
nand UO_1956 (O_1956,N_23048,N_23850);
or UO_1957 (O_1957,N_22597,N_20246);
nor UO_1958 (O_1958,N_20141,N_20544);
or UO_1959 (O_1959,N_21131,N_24874);
or UO_1960 (O_1960,N_21496,N_20385);
nor UO_1961 (O_1961,N_20763,N_22690);
nand UO_1962 (O_1962,N_23403,N_20157);
or UO_1963 (O_1963,N_20963,N_20627);
and UO_1964 (O_1964,N_21691,N_20434);
and UO_1965 (O_1965,N_20760,N_21891);
nand UO_1966 (O_1966,N_20917,N_24707);
nand UO_1967 (O_1967,N_23437,N_20765);
nor UO_1968 (O_1968,N_23606,N_20358);
or UO_1969 (O_1969,N_21939,N_23033);
and UO_1970 (O_1970,N_22892,N_21619);
and UO_1971 (O_1971,N_20598,N_24328);
nor UO_1972 (O_1972,N_21324,N_22679);
nand UO_1973 (O_1973,N_22716,N_24423);
and UO_1974 (O_1974,N_22907,N_22663);
or UO_1975 (O_1975,N_21818,N_22199);
nor UO_1976 (O_1976,N_22416,N_23766);
or UO_1977 (O_1977,N_20095,N_21885);
or UO_1978 (O_1978,N_23684,N_22808);
nand UO_1979 (O_1979,N_21250,N_24852);
or UO_1980 (O_1980,N_22482,N_20568);
or UO_1981 (O_1981,N_21097,N_21241);
xnor UO_1982 (O_1982,N_24861,N_22844);
nand UO_1983 (O_1983,N_23585,N_22254);
or UO_1984 (O_1984,N_21572,N_24956);
or UO_1985 (O_1985,N_20698,N_20776);
and UO_1986 (O_1986,N_24574,N_22667);
nand UO_1987 (O_1987,N_22697,N_21843);
and UO_1988 (O_1988,N_24289,N_23692);
and UO_1989 (O_1989,N_20102,N_22286);
or UO_1990 (O_1990,N_23040,N_23655);
nor UO_1991 (O_1991,N_21055,N_22985);
and UO_1992 (O_1992,N_22493,N_23966);
and UO_1993 (O_1993,N_20413,N_20086);
nand UO_1994 (O_1994,N_20820,N_22544);
and UO_1995 (O_1995,N_22631,N_23949);
or UO_1996 (O_1996,N_23891,N_22819);
or UO_1997 (O_1997,N_22460,N_20053);
and UO_1998 (O_1998,N_20814,N_20131);
nand UO_1999 (O_1999,N_23703,N_23813);
nor UO_2000 (O_2000,N_20783,N_21576);
and UO_2001 (O_2001,N_21821,N_22242);
and UO_2002 (O_2002,N_20252,N_21894);
nand UO_2003 (O_2003,N_20918,N_21964);
and UO_2004 (O_2004,N_21558,N_23400);
nand UO_2005 (O_2005,N_22599,N_20883);
and UO_2006 (O_2006,N_24899,N_21766);
nand UO_2007 (O_2007,N_23138,N_23548);
or UO_2008 (O_2008,N_20212,N_24449);
nand UO_2009 (O_2009,N_22743,N_23159);
nor UO_2010 (O_2010,N_24478,N_21045);
and UO_2011 (O_2011,N_21054,N_20870);
or UO_2012 (O_2012,N_20126,N_20363);
nand UO_2013 (O_2013,N_23578,N_23943);
or UO_2014 (O_2014,N_20139,N_20935);
or UO_2015 (O_2015,N_23754,N_22394);
nor UO_2016 (O_2016,N_21820,N_22686);
nand UO_2017 (O_2017,N_20778,N_21717);
nand UO_2018 (O_2018,N_22673,N_24140);
and UO_2019 (O_2019,N_21809,N_20890);
nand UO_2020 (O_2020,N_23653,N_21760);
nor UO_2021 (O_2021,N_20254,N_20430);
and UO_2022 (O_2022,N_21420,N_24350);
and UO_2023 (O_2023,N_20980,N_23359);
nor UO_2024 (O_2024,N_24546,N_24467);
nand UO_2025 (O_2025,N_20887,N_21965);
nor UO_2026 (O_2026,N_24969,N_21025);
and UO_2027 (O_2027,N_23770,N_23748);
nor UO_2028 (O_2028,N_21571,N_24358);
and UO_2029 (O_2029,N_24549,N_20939);
nor UO_2030 (O_2030,N_24523,N_21379);
nand UO_2031 (O_2031,N_24578,N_20615);
nand UO_2032 (O_2032,N_23657,N_21521);
and UO_2033 (O_2033,N_21296,N_20613);
nor UO_2034 (O_2034,N_21007,N_21405);
and UO_2035 (O_2035,N_23266,N_24336);
nor UO_2036 (O_2036,N_24677,N_20188);
and UO_2037 (O_2037,N_22897,N_22264);
nor UO_2038 (O_2038,N_24723,N_22842);
or UO_2039 (O_2039,N_21184,N_22431);
nand UO_2040 (O_2040,N_22219,N_20614);
nor UO_2041 (O_2041,N_20250,N_24070);
or UO_2042 (O_2042,N_23031,N_20129);
or UO_2043 (O_2043,N_20354,N_21412);
and UO_2044 (O_2044,N_22558,N_22828);
or UO_2045 (O_2045,N_21150,N_22820);
nand UO_2046 (O_2046,N_22013,N_22051);
or UO_2047 (O_2047,N_24084,N_20616);
nor UO_2048 (O_2048,N_22996,N_24722);
and UO_2049 (O_2049,N_24218,N_20048);
nand UO_2050 (O_2050,N_23978,N_21506);
and UO_2051 (O_2051,N_22320,N_22411);
or UO_2052 (O_2052,N_24813,N_21662);
nand UO_2053 (O_2053,N_20812,N_21897);
and UO_2054 (O_2054,N_20565,N_22583);
or UO_2055 (O_2055,N_24182,N_23238);
or UO_2056 (O_2056,N_22349,N_20025);
and UO_2057 (O_2057,N_22756,N_24087);
nor UO_2058 (O_2058,N_23756,N_24945);
nor UO_2059 (O_2059,N_20992,N_24442);
nor UO_2060 (O_2060,N_22167,N_21457);
or UO_2061 (O_2061,N_21193,N_24113);
and UO_2062 (O_2062,N_23698,N_21827);
nor UO_2063 (O_2063,N_20462,N_21401);
nor UO_2064 (O_2064,N_20350,N_22383);
or UO_2065 (O_2065,N_20406,N_24136);
nor UO_2066 (O_2066,N_24383,N_24946);
and UO_2067 (O_2067,N_21882,N_20944);
and UO_2068 (O_2068,N_21394,N_24573);
nor UO_2069 (O_2069,N_22143,N_20976);
and UO_2070 (O_2070,N_20419,N_24828);
nand UO_2071 (O_2071,N_21086,N_20684);
or UO_2072 (O_2072,N_22171,N_22615);
xnor UO_2073 (O_2073,N_24513,N_22179);
or UO_2074 (O_2074,N_24596,N_24560);
or UO_2075 (O_2075,N_23964,N_20062);
nand UO_2076 (O_2076,N_22936,N_20632);
and UO_2077 (O_2077,N_23127,N_22465);
and UO_2078 (O_2078,N_22102,N_20486);
or UO_2079 (O_2079,N_20370,N_22676);
and UO_2080 (O_2080,N_23533,N_24495);
and UO_2081 (O_2081,N_21508,N_23289);
nor UO_2082 (O_2082,N_24413,N_23762);
nand UO_2083 (O_2083,N_21318,N_24225);
and UO_2084 (O_2084,N_23810,N_24623);
and UO_2085 (O_2085,N_22127,N_22852);
and UO_2086 (O_2086,N_23557,N_21973);
and UO_2087 (O_2087,N_24299,N_23399);
nand UO_2088 (O_2088,N_24315,N_21137);
nand UO_2089 (O_2089,N_21056,N_24711);
or UO_2090 (O_2090,N_23023,N_20537);
nand UO_2091 (O_2091,N_21847,N_24921);
or UO_2092 (O_2092,N_21041,N_24376);
or UO_2093 (O_2093,N_22324,N_20481);
nand UO_2094 (O_2094,N_20852,N_24751);
nor UO_2095 (O_2095,N_23824,N_22301);
nand UO_2096 (O_2096,N_24027,N_23089);
nand UO_2097 (O_2097,N_22340,N_23671);
nand UO_2098 (O_2098,N_20916,N_23384);
nor UO_2099 (O_2099,N_20077,N_23480);
nand UO_2100 (O_2100,N_22231,N_22657);
nand UO_2101 (O_2101,N_20418,N_22909);
or UO_2102 (O_2102,N_21197,N_24059);
and UO_2103 (O_2103,N_24044,N_22741);
and UO_2104 (O_2104,N_23927,N_20120);
nor UO_2105 (O_2105,N_23983,N_22215);
xor UO_2106 (O_2106,N_21189,N_22487);
nand UO_2107 (O_2107,N_23101,N_23996);
and UO_2108 (O_2108,N_22486,N_20377);
or UO_2109 (O_2109,N_22980,N_22748);
or UO_2110 (O_2110,N_21522,N_22944);
and UO_2111 (O_2111,N_24157,N_22252);
nand UO_2112 (O_2112,N_22296,N_24356);
and UO_2113 (O_2113,N_22940,N_20633);
or UO_2114 (O_2114,N_24319,N_24108);
nor UO_2115 (O_2115,N_21344,N_24877);
nand UO_2116 (O_2116,N_21999,N_22385);
nor UO_2117 (O_2117,N_22857,N_24035);
nor UO_2118 (O_2118,N_24082,N_24528);
or UO_2119 (O_2119,N_24178,N_21363);
nand UO_2120 (O_2120,N_20824,N_20957);
nand UO_2121 (O_2121,N_20874,N_20005);
and UO_2122 (O_2122,N_21944,N_21407);
and UO_2123 (O_2123,N_23623,N_21773);
xnor UO_2124 (O_2124,N_22833,N_20836);
or UO_2125 (O_2125,N_23811,N_24300);
or UO_2126 (O_2126,N_23662,N_20784);
nor UO_2127 (O_2127,N_24792,N_24042);
and UO_2128 (O_2128,N_24335,N_22521);
nor UO_2129 (O_2129,N_21941,N_23975);
or UO_2130 (O_2130,N_21440,N_24434);
nor UO_2131 (O_2131,N_21851,N_21972);
nor UO_2132 (O_2132,N_20550,N_22609);
and UO_2133 (O_2133,N_22883,N_21469);
and UO_2134 (O_2134,N_22650,N_24466);
or UO_2135 (O_2135,N_21359,N_20215);
and UO_2136 (O_2136,N_23945,N_24604);
and UO_2137 (O_2137,N_24624,N_20084);
xnor UO_2138 (O_2138,N_24901,N_23432);
nand UO_2139 (O_2139,N_24272,N_21391);
xor UO_2140 (O_2140,N_24543,N_23537);
and UO_2141 (O_2141,N_23442,N_23638);
nand UO_2142 (O_2142,N_20607,N_23907);
and UO_2143 (O_2143,N_20560,N_21048);
or UO_2144 (O_2144,N_22348,N_21688);
and UO_2145 (O_2145,N_20464,N_20989);
nor UO_2146 (O_2146,N_24520,N_23492);
nor UO_2147 (O_2147,N_24425,N_22112);
nor UO_2148 (O_2148,N_24072,N_23164);
or UO_2149 (O_2149,N_21284,N_24102);
nor UO_2150 (O_2150,N_21644,N_20285);
and UO_2151 (O_2151,N_23411,N_23110);
or UO_2152 (O_2152,N_24060,N_24085);
and UO_2153 (O_2153,N_22488,N_23017);
and UO_2154 (O_2154,N_20662,N_24160);
nand UO_2155 (O_2155,N_21461,N_23453);
nand UO_2156 (O_2156,N_20694,N_24966);
or UO_2157 (O_2157,N_24349,N_21265);
or UO_2158 (O_2158,N_21153,N_20101);
nor UO_2159 (O_2159,N_20036,N_22641);
nand UO_2160 (O_2160,N_21922,N_23612);
nand UO_2161 (O_2161,N_20925,N_24557);
and UO_2162 (O_2162,N_20154,N_20541);
and UO_2163 (O_2163,N_20000,N_22041);
or UO_2164 (O_2164,N_22247,N_24222);
and UO_2165 (O_2165,N_21219,N_24395);
nor UO_2166 (O_2166,N_23052,N_21280);
or UO_2167 (O_2167,N_22325,N_20247);
nand UO_2168 (O_2168,N_20028,N_22680);
nor UO_2169 (O_2169,N_20179,N_24858);
nor UO_2170 (O_2170,N_21946,N_21306);
or UO_2171 (O_2171,N_23372,N_24343);
nand UO_2172 (O_2172,N_24759,N_24363);
nand UO_2173 (O_2173,N_20507,N_24704);
or UO_2174 (O_2174,N_20646,N_21029);
nand UO_2175 (O_2175,N_23837,N_24962);
and UO_2176 (O_2176,N_22585,N_22275);
nand UO_2177 (O_2177,N_20885,N_21031);
nand UO_2178 (O_2178,N_24607,N_21520);
and UO_2179 (O_2179,N_20850,N_20943);
nand UO_2180 (O_2180,N_24508,N_20375);
or UO_2181 (O_2181,N_24390,N_22682);
and UO_2182 (O_2182,N_20140,N_21300);
and UO_2183 (O_2183,N_23789,N_22042);
xor UO_2184 (O_2184,N_20003,N_24483);
or UO_2185 (O_2185,N_24599,N_23292);
and UO_2186 (O_2186,N_21761,N_23378);
nand UO_2187 (O_2187,N_22335,N_21132);
nand UO_2188 (O_2188,N_21543,N_20290);
or UO_2189 (O_2189,N_24805,N_23482);
and UO_2190 (O_2190,N_21382,N_20286);
nor UO_2191 (O_2191,N_23829,N_22003);
nor UO_2192 (O_2192,N_24479,N_24428);
and UO_2193 (O_2193,N_20530,N_22660);
nand UO_2194 (O_2194,N_24352,N_20405);
nor UO_2195 (O_2195,N_23393,N_24062);
nor UO_2196 (O_2196,N_22954,N_23887);
and UO_2197 (O_2197,N_24255,N_21743);
or UO_2198 (O_2198,N_22213,N_23711);
nand UO_2199 (O_2199,N_23903,N_24551);
or UO_2200 (O_2200,N_24112,N_23214);
or UO_2201 (O_2201,N_21395,N_22120);
or UO_2202 (O_2202,N_23510,N_20774);
or UO_2203 (O_2203,N_21633,N_21068);
nor UO_2204 (O_2204,N_23146,N_22204);
nor UO_2205 (O_2205,N_24786,N_23704);
nor UO_2206 (O_2206,N_22751,N_23314);
nor UO_2207 (O_2207,N_24487,N_21739);
nand UO_2208 (O_2208,N_22845,N_24346);
and UO_2209 (O_2209,N_24600,N_21966);
nor UO_2210 (O_2210,N_22227,N_22018);
or UO_2211 (O_2211,N_24459,N_24595);
and UO_2212 (O_2212,N_21510,N_23346);
or UO_2213 (O_2213,N_22014,N_21450);
or UO_2214 (O_2214,N_21322,N_22799);
nor UO_2215 (O_2215,N_21814,N_22902);
or UO_2216 (O_2216,N_20346,N_20518);
nand UO_2217 (O_2217,N_21368,N_22137);
and UO_2218 (O_2218,N_23203,N_24516);
and UO_2219 (O_2219,N_24705,N_23636);
or UO_2220 (O_2220,N_22755,N_23879);
and UO_2221 (O_2221,N_22052,N_23389);
and UO_2222 (O_2222,N_22364,N_23795);
and UO_2223 (O_2223,N_23886,N_22736);
or UO_2224 (O_2224,N_20334,N_21952);
and UO_2225 (O_2225,N_20040,N_23233);
nor UO_2226 (O_2226,N_23690,N_21913);
or UO_2227 (O_2227,N_20266,N_24745);
and UO_2228 (O_2228,N_24212,N_23313);
nand UO_2229 (O_2229,N_22391,N_22059);
or UO_2230 (O_2230,N_21290,N_20275);
and UO_2231 (O_2231,N_20217,N_23179);
and UO_2232 (O_2232,N_21542,N_24134);
and UO_2233 (O_2233,N_20902,N_24930);
nor UO_2234 (O_2234,N_24991,N_21859);
or UO_2235 (O_2235,N_24579,N_23724);
or UO_2236 (O_2236,N_22960,N_23043);
nand UO_2237 (O_2237,N_23487,N_21335);
or UO_2238 (O_2238,N_21336,N_23365);
and UO_2239 (O_2239,N_20622,N_24111);
and UO_2240 (O_2240,N_23064,N_23274);
and UO_2241 (O_2241,N_23227,N_24632);
nor UO_2242 (O_2242,N_21166,N_23899);
nand UO_2243 (O_2243,N_20804,N_20514);
nand UO_2244 (O_2244,N_20241,N_22744);
nor UO_2245 (O_2245,N_20498,N_21726);
and UO_2246 (O_2246,N_23356,N_21442);
and UO_2247 (O_2247,N_23474,N_22913);
and UO_2248 (O_2248,N_24665,N_24765);
nor UO_2249 (O_2249,N_21887,N_23058);
nand UO_2250 (O_2250,N_20042,N_24435);
nand UO_2251 (O_2251,N_23382,N_23629);
or UO_2252 (O_2252,N_24214,N_21838);
or UO_2253 (O_2253,N_21526,N_20012);
or UO_2254 (O_2254,N_21376,N_24473);
or UO_2255 (O_2255,N_24219,N_24117);
and UO_2256 (O_2256,N_23634,N_21862);
or UO_2257 (O_2257,N_21267,N_24246);
and UO_2258 (O_2258,N_20225,N_24947);
and UO_2259 (O_2259,N_20489,N_22390);
nor UO_2260 (O_2260,N_21751,N_22457);
or UO_2261 (O_2261,N_20600,N_24440);
and UO_2262 (O_2262,N_21879,N_21565);
or UO_2263 (O_2263,N_20819,N_20466);
and UO_2264 (O_2264,N_23228,N_20199);
or UO_2265 (O_2265,N_23286,N_23547);
nand UO_2266 (O_2266,N_21393,N_23626);
nor UO_2267 (O_2267,N_24101,N_20232);
and UO_2268 (O_2268,N_24063,N_21548);
nand UO_2269 (O_2269,N_23244,N_23104);
and UO_2270 (O_2270,N_21147,N_20502);
nand UO_2271 (O_2271,N_20683,N_21653);
and UO_2272 (O_2272,N_22687,N_22500);
and UO_2273 (O_2273,N_22627,N_21340);
nand UO_2274 (O_2274,N_23236,N_24964);
nor UO_2275 (O_2275,N_22438,N_20716);
or UO_2276 (O_2276,N_24884,N_24048);
nor UO_2277 (O_2277,N_22930,N_23580);
nor UO_2278 (O_2278,N_23148,N_22407);
or UO_2279 (O_2279,N_23241,N_20449);
xor UO_2280 (O_2280,N_21083,N_21509);
or UO_2281 (O_2281,N_23428,N_23507);
nand UO_2282 (O_2282,N_21107,N_24545);
nand UO_2283 (O_2283,N_20472,N_24744);
or UO_2284 (O_2284,N_22261,N_24730);
and UO_2285 (O_2285,N_23090,N_20162);
or UO_2286 (O_2286,N_23843,N_22057);
nand UO_2287 (O_2287,N_22467,N_20093);
nor UO_2288 (O_2288,N_21203,N_21606);
and UO_2289 (O_2289,N_24491,N_23215);
nor UO_2290 (O_2290,N_20369,N_20440);
or UO_2291 (O_2291,N_23642,N_24729);
or UO_2292 (O_2292,N_22990,N_23323);
nor UO_2293 (O_2293,N_24239,N_20417);
or UO_2294 (O_2294,N_23768,N_21014);
nand UO_2295 (O_2295,N_23826,N_21492);
nor UO_2296 (O_2296,N_22280,N_22105);
or UO_2297 (O_2297,N_20061,N_23379);
nor UO_2298 (O_2298,N_20747,N_23564);
and UO_2299 (O_2299,N_21388,N_23297);
nand UO_2300 (O_2300,N_22628,N_21806);
and UO_2301 (O_2301,N_21253,N_24066);
nand UO_2302 (O_2302,N_24184,N_22210);
and UO_2303 (O_2303,N_20196,N_22303);
nor UO_2304 (O_2304,N_24654,N_24976);
nor UO_2305 (O_2305,N_22290,N_20669);
nor UO_2306 (O_2306,N_23371,N_20551);
or UO_2307 (O_2307,N_22331,N_22336);
and UO_2308 (O_2308,N_24258,N_24531);
and UO_2309 (O_2309,N_23329,N_22656);
nand UO_2310 (O_2310,N_20594,N_20300);
and UO_2311 (O_2311,N_23374,N_23900);
nor UO_2312 (O_2312,N_21947,N_23812);
nor UO_2313 (O_2313,N_20510,N_22129);
and UO_2314 (O_2314,N_23611,N_21637);
or UO_2315 (O_2315,N_21579,N_22161);
and UO_2316 (O_2316,N_22977,N_23019);
or UO_2317 (O_2317,N_22941,N_22915);
nor UO_2318 (O_2318,N_20878,N_24809);
nor UO_2319 (O_2319,N_21279,N_23599);
or UO_2320 (O_2320,N_23092,N_24236);
nor UO_2321 (O_2321,N_24364,N_20103);
or UO_2322 (O_2322,N_24754,N_20659);
and UO_2323 (O_2323,N_20880,N_24147);
nor UO_2324 (O_2324,N_22956,N_24853);
nor UO_2325 (O_2325,N_21331,N_24779);
nand UO_2326 (O_2326,N_20949,N_21277);
nand UO_2327 (O_2327,N_24866,N_24981);
or UO_2328 (O_2328,N_23973,N_24798);
and UO_2329 (O_2329,N_22019,N_23697);
nand UO_2330 (O_2330,N_24916,N_24287);
nor UO_2331 (O_2331,N_21951,N_24728);
or UO_2332 (O_2332,N_24539,N_23990);
nand UO_2333 (O_2333,N_24472,N_21837);
nor UO_2334 (O_2334,N_22688,N_20792);
nor UO_2335 (O_2335,N_24418,N_20143);
nand UO_2336 (O_2336,N_24230,N_22805);
nor UO_2337 (O_2337,N_23567,N_22962);
nand UO_2338 (O_2338,N_23677,N_21145);
nor UO_2339 (O_2339,N_23952,N_20044);
and UO_2340 (O_2340,N_21514,N_20668);
nand UO_2341 (O_2341,N_24788,N_23412);
nor UO_2342 (O_2342,N_22193,N_24198);
nor UO_2343 (O_2343,N_24443,N_23871);
or UO_2344 (O_2344,N_24293,N_20224);
nand UO_2345 (O_2345,N_22699,N_22831);
nor UO_2346 (O_2346,N_21477,N_24789);
or UO_2347 (O_2347,N_23579,N_23496);
nor UO_2348 (O_2348,N_20230,N_20227);
or UO_2349 (O_2349,N_20436,N_24591);
nand UO_2350 (O_2350,N_22693,N_20860);
and UO_2351 (O_2351,N_20400,N_24695);
nand UO_2352 (O_2352,N_23107,N_21985);
or UO_2353 (O_2353,N_23369,N_20428);
nor UO_2354 (O_2354,N_21983,N_21373);
or UO_2355 (O_2355,N_23067,N_21180);
nor UO_2356 (O_2356,N_22200,N_24708);
and UO_2357 (O_2357,N_20640,N_24795);
nand UO_2358 (O_2358,N_24091,N_24123);
or UO_2359 (O_2359,N_23977,N_24260);
nor UO_2360 (O_2360,N_23461,N_24702);
nand UO_2361 (O_2361,N_21781,N_20692);
and UO_2362 (O_2362,N_23447,N_20060);
and UO_2363 (O_2363,N_22315,N_22818);
nor UO_2364 (O_2364,N_21740,N_24974);
nand UO_2365 (O_2365,N_24034,N_23010);
nand UO_2366 (O_2366,N_21414,N_20395);
nor UO_2367 (O_2367,N_23050,N_22837);
and UO_2368 (O_2368,N_22994,N_23644);
nor UO_2369 (O_2369,N_24510,N_21599);
and UO_2370 (O_2370,N_21480,N_21687);
nor UO_2371 (O_2371,N_23026,N_23882);
nand UO_2372 (O_2372,N_24220,N_20432);
nor UO_2373 (O_2373,N_24738,N_20556);
and UO_2374 (O_2374,N_22166,N_21035);
or UO_2375 (O_2375,N_24432,N_20138);
xor UO_2376 (O_2376,N_24834,N_20386);
nand UO_2377 (O_2377,N_22702,N_20651);
nor UO_2378 (O_2378,N_22759,N_24793);
and UO_2379 (O_2379,N_24615,N_23625);
nand UO_2380 (O_2380,N_20702,N_21374);
or UO_2381 (O_2381,N_21226,N_21486);
nor UO_2382 (O_2382,N_22658,N_24252);
or UO_2383 (O_2383,N_21190,N_23915);
or UO_2384 (O_2384,N_21354,N_20478);
nand UO_2385 (O_2385,N_23124,N_23916);
or UO_2386 (O_2386,N_24103,N_23946);
xor UO_2387 (O_2387,N_23631,N_23097);
nand UO_2388 (O_2388,N_20801,N_24927);
and UO_2389 (O_2389,N_22387,N_23613);
or UO_2390 (O_2390,N_21358,N_22539);
xor UO_2391 (O_2391,N_20117,N_21413);
nand UO_2392 (O_2392,N_23256,N_24307);
and UO_2393 (O_2393,N_22078,N_23467);
and UO_2394 (O_2394,N_24257,N_20443);
or UO_2395 (O_2395,N_24298,N_20365);
nand UO_2396 (O_2396,N_23011,N_20707);
and UO_2397 (O_2397,N_23744,N_21347);
and UO_2398 (O_2398,N_21103,N_23823);
or UO_2399 (O_2399,N_22796,N_24295);
nor UO_2400 (O_2400,N_23247,N_23495);
and UO_2401 (O_2401,N_20167,N_24918);
nor UO_2402 (O_2402,N_22529,N_22547);
or UO_2403 (O_2403,N_21905,N_21415);
nor UO_2404 (O_2404,N_23349,N_24973);
and UO_2405 (O_2405,N_20001,N_22920);
nor UO_2406 (O_2406,N_24687,N_24481);
and UO_2407 (O_2407,N_21073,N_21310);
xor UO_2408 (O_2408,N_23188,N_21248);
nand UO_2409 (O_2409,N_21084,N_24589);
and UO_2410 (O_2410,N_21679,N_24998);
and UO_2411 (O_2411,N_24561,N_24602);
or UO_2412 (O_2412,N_23115,N_22283);
and UO_2413 (O_2413,N_22540,N_22150);
nor UO_2414 (O_2414,N_23632,N_24078);
or UO_2415 (O_2415,N_23536,N_20962);
nor UO_2416 (O_2416,N_23143,N_23654);
or UO_2417 (O_2417,N_23469,N_20374);
and UO_2418 (O_2418,N_23985,N_23535);
or UO_2419 (O_2419,N_24141,N_23716);
and UO_2420 (O_2420,N_20314,N_20332);
and UO_2421 (O_2421,N_23980,N_23804);
nand UO_2422 (O_2422,N_21878,N_24785);
nand UO_2423 (O_2423,N_23733,N_24002);
or UO_2424 (O_2424,N_22830,N_23151);
or UO_2425 (O_2425,N_23270,N_20573);
or UO_2426 (O_2426,N_21044,N_22284);
and UO_2427 (O_2427,N_24388,N_22339);
or UO_2428 (O_2428,N_21874,N_20563);
nor UO_2429 (O_2429,N_20701,N_23099);
nand UO_2430 (O_2430,N_24242,N_23925);
nor UO_2431 (O_2431,N_20367,N_24041);
nand UO_2432 (O_2432,N_24320,N_22536);
nor UO_2433 (O_2433,N_20815,N_24518);
xor UO_2434 (O_2434,N_22534,N_22535);
nor UO_2435 (O_2435,N_20803,N_20161);
nor UO_2436 (O_2436,N_23839,N_22169);
nand UO_2437 (O_2437,N_21125,N_20118);
and UO_2438 (O_2438,N_21403,N_21270);
nor UO_2439 (O_2439,N_22472,N_20007);
nand UO_2440 (O_2440,N_24594,N_20343);
and UO_2441 (O_2441,N_20579,N_21076);
nand UO_2442 (O_2442,N_22235,N_22781);
nand UO_2443 (O_2443,N_21570,N_21020);
or UO_2444 (O_2444,N_22610,N_21019);
nand UO_2445 (O_2445,N_23586,N_21448);
or UO_2446 (O_2446,N_23320,N_22683);
nor UO_2447 (O_2447,N_21257,N_22967);
xnor UO_2448 (O_2448,N_23395,N_20164);
and UO_2449 (O_2449,N_23066,N_22205);
nor UO_2450 (O_2450,N_24477,N_22851);
and UO_2451 (O_2451,N_22158,N_22062);
nand UO_2452 (O_2452,N_21836,N_21365);
and UO_2453 (O_2453,N_20050,N_24142);
nor UO_2454 (O_2454,N_20504,N_23225);
nand UO_2455 (O_2455,N_21108,N_24168);
xor UO_2456 (O_2456,N_21967,N_22675);
nand UO_2457 (O_2457,N_22047,N_23113);
and UO_2458 (O_2458,N_23788,N_22645);
and UO_2459 (O_2459,N_20009,N_23694);
nor UO_2460 (O_2460,N_20993,N_21289);
nor UO_2461 (O_2461,N_20839,N_24512);
nand UO_2462 (O_2462,N_20538,N_23571);
and UO_2463 (O_2463,N_23581,N_20605);
or UO_2464 (O_2464,N_23528,N_21649);
or UO_2465 (O_2465,N_22719,N_24800);
nor UO_2466 (O_2466,N_22612,N_21587);
or UO_2467 (O_2467,N_21173,N_22651);
and UO_2468 (O_2468,N_24455,N_20726);
or UO_2469 (O_2469,N_24984,N_21541);
or UO_2470 (O_2470,N_24818,N_21877);
and UO_2471 (O_2471,N_23260,N_23231);
and UO_2472 (O_2472,N_24266,N_24742);
nor UO_2473 (O_2473,N_23497,N_21559);
nand UO_2474 (O_2474,N_23053,N_20134);
nor UO_2475 (O_2475,N_21889,N_24846);
or UO_2476 (O_2476,N_23160,N_20015);
or UO_2477 (O_2477,N_23479,N_20446);
or UO_2478 (O_2478,N_21630,N_21004);
nor UO_2479 (O_2479,N_23114,N_21808);
or UO_2480 (O_2480,N_24064,N_20457);
xor UO_2481 (O_2481,N_22145,N_20843);
or UO_2482 (O_2482,N_21417,N_23465);
nand UO_2483 (O_2483,N_20352,N_24492);
nor UO_2484 (O_2484,N_22048,N_20886);
and UO_2485 (O_2485,N_22025,N_24802);
nand UO_2486 (O_2486,N_24651,N_24896);
nand UO_2487 (O_2487,N_22308,N_22623);
and UO_2488 (O_2488,N_23409,N_21273);
nor UO_2489 (O_2489,N_24867,N_23070);
xor UO_2490 (O_2490,N_22608,N_22758);
and UO_2491 (O_2491,N_22964,N_21992);
nand UO_2492 (O_2492,N_23809,N_21979);
or UO_2493 (O_2493,N_22279,N_22863);
or UO_2494 (O_2494,N_24715,N_21135);
and UO_2495 (O_2495,N_21540,N_20178);
nand UO_2496 (O_2496,N_20249,N_22240);
or UO_2497 (O_2497,N_20871,N_22611);
and UO_2498 (O_2498,N_22033,N_23377);
nand UO_2499 (O_2499,N_23319,N_20112);
or UO_2500 (O_2500,N_24373,N_21162);
or UO_2501 (O_2501,N_20403,N_21668);
xnor UO_2502 (O_2502,N_22971,N_20190);
and UO_2503 (O_2503,N_23770,N_23481);
and UO_2504 (O_2504,N_24477,N_20766);
nand UO_2505 (O_2505,N_21615,N_24081);
nand UO_2506 (O_2506,N_23113,N_24255);
or UO_2507 (O_2507,N_20819,N_21267);
or UO_2508 (O_2508,N_22943,N_24629);
or UO_2509 (O_2509,N_23891,N_22058);
or UO_2510 (O_2510,N_23163,N_20054);
nor UO_2511 (O_2511,N_24622,N_23748);
nor UO_2512 (O_2512,N_22498,N_22171);
nor UO_2513 (O_2513,N_21898,N_20392);
or UO_2514 (O_2514,N_21657,N_24284);
nand UO_2515 (O_2515,N_22999,N_22462);
or UO_2516 (O_2516,N_21432,N_23920);
or UO_2517 (O_2517,N_21773,N_20683);
nand UO_2518 (O_2518,N_23812,N_24313);
or UO_2519 (O_2519,N_22962,N_21962);
nor UO_2520 (O_2520,N_23007,N_22582);
or UO_2521 (O_2521,N_24736,N_23169);
nand UO_2522 (O_2522,N_21165,N_24618);
nor UO_2523 (O_2523,N_21528,N_21385);
or UO_2524 (O_2524,N_24175,N_24469);
or UO_2525 (O_2525,N_23885,N_20797);
nor UO_2526 (O_2526,N_24389,N_20940);
nor UO_2527 (O_2527,N_20204,N_24163);
or UO_2528 (O_2528,N_21112,N_23133);
or UO_2529 (O_2529,N_24010,N_22245);
nand UO_2530 (O_2530,N_23333,N_20853);
and UO_2531 (O_2531,N_24608,N_20973);
and UO_2532 (O_2532,N_20041,N_23983);
xor UO_2533 (O_2533,N_20755,N_20857);
or UO_2534 (O_2534,N_23931,N_21227);
nand UO_2535 (O_2535,N_22421,N_23118);
nor UO_2536 (O_2536,N_21802,N_23397);
nor UO_2537 (O_2537,N_21246,N_22312);
or UO_2538 (O_2538,N_23356,N_23370);
or UO_2539 (O_2539,N_22003,N_23474);
xor UO_2540 (O_2540,N_24831,N_22193);
or UO_2541 (O_2541,N_23829,N_21452);
nand UO_2542 (O_2542,N_24297,N_23432);
and UO_2543 (O_2543,N_24645,N_22094);
nor UO_2544 (O_2544,N_23595,N_22055);
nand UO_2545 (O_2545,N_21604,N_20724);
nor UO_2546 (O_2546,N_22802,N_21283);
nor UO_2547 (O_2547,N_24630,N_24301);
nand UO_2548 (O_2548,N_21152,N_22881);
and UO_2549 (O_2549,N_22672,N_23321);
or UO_2550 (O_2550,N_21523,N_22921);
or UO_2551 (O_2551,N_20906,N_21340);
nand UO_2552 (O_2552,N_20066,N_23049);
nand UO_2553 (O_2553,N_22304,N_23922);
and UO_2554 (O_2554,N_24000,N_20978);
nor UO_2555 (O_2555,N_21792,N_23171);
and UO_2556 (O_2556,N_24771,N_23114);
nand UO_2557 (O_2557,N_20761,N_20237);
and UO_2558 (O_2558,N_21442,N_23520);
nand UO_2559 (O_2559,N_22502,N_22148);
or UO_2560 (O_2560,N_24920,N_21324);
nand UO_2561 (O_2561,N_24897,N_24614);
and UO_2562 (O_2562,N_21044,N_22392);
and UO_2563 (O_2563,N_23158,N_22386);
xnor UO_2564 (O_2564,N_21795,N_24165);
or UO_2565 (O_2565,N_22344,N_22264);
nand UO_2566 (O_2566,N_24450,N_22591);
nand UO_2567 (O_2567,N_21483,N_20698);
nor UO_2568 (O_2568,N_20421,N_23079);
and UO_2569 (O_2569,N_24661,N_21726);
and UO_2570 (O_2570,N_20662,N_24716);
xnor UO_2571 (O_2571,N_23696,N_22908);
nand UO_2572 (O_2572,N_22284,N_22842);
nor UO_2573 (O_2573,N_24184,N_22907);
nor UO_2574 (O_2574,N_20091,N_23251);
nor UO_2575 (O_2575,N_24860,N_22480);
nor UO_2576 (O_2576,N_22102,N_22322);
and UO_2577 (O_2577,N_20847,N_20720);
and UO_2578 (O_2578,N_23186,N_21039);
nor UO_2579 (O_2579,N_21690,N_21083);
or UO_2580 (O_2580,N_24967,N_22702);
nor UO_2581 (O_2581,N_23685,N_20317);
nor UO_2582 (O_2582,N_20302,N_22938);
and UO_2583 (O_2583,N_21865,N_23642);
nor UO_2584 (O_2584,N_23389,N_24580);
nand UO_2585 (O_2585,N_22295,N_20906);
nor UO_2586 (O_2586,N_21071,N_23849);
or UO_2587 (O_2587,N_24540,N_24770);
nor UO_2588 (O_2588,N_22615,N_22807);
nand UO_2589 (O_2589,N_21093,N_24998);
nand UO_2590 (O_2590,N_22828,N_20056);
nor UO_2591 (O_2591,N_24092,N_20984);
nand UO_2592 (O_2592,N_21044,N_24244);
and UO_2593 (O_2593,N_24324,N_24588);
nor UO_2594 (O_2594,N_23829,N_21643);
nor UO_2595 (O_2595,N_22313,N_23014);
nor UO_2596 (O_2596,N_20483,N_24312);
nor UO_2597 (O_2597,N_20398,N_21138);
and UO_2598 (O_2598,N_22335,N_24843);
nor UO_2599 (O_2599,N_24556,N_20784);
or UO_2600 (O_2600,N_24418,N_24132);
nand UO_2601 (O_2601,N_20680,N_24420);
or UO_2602 (O_2602,N_24985,N_21506);
or UO_2603 (O_2603,N_21801,N_24652);
nand UO_2604 (O_2604,N_22148,N_22261);
nor UO_2605 (O_2605,N_23636,N_22350);
or UO_2606 (O_2606,N_23799,N_23972);
nand UO_2607 (O_2607,N_23254,N_22584);
or UO_2608 (O_2608,N_22006,N_20350);
nand UO_2609 (O_2609,N_22350,N_23821);
or UO_2610 (O_2610,N_20717,N_22467);
and UO_2611 (O_2611,N_24242,N_23143);
nor UO_2612 (O_2612,N_20880,N_21220);
nand UO_2613 (O_2613,N_20993,N_21489);
nand UO_2614 (O_2614,N_22662,N_23289);
nand UO_2615 (O_2615,N_20208,N_22178);
and UO_2616 (O_2616,N_22288,N_23460);
and UO_2617 (O_2617,N_22215,N_23047);
and UO_2618 (O_2618,N_21714,N_24283);
nand UO_2619 (O_2619,N_23860,N_20042);
nor UO_2620 (O_2620,N_24429,N_22100);
or UO_2621 (O_2621,N_24766,N_24857);
or UO_2622 (O_2622,N_23167,N_21365);
or UO_2623 (O_2623,N_23122,N_23830);
nand UO_2624 (O_2624,N_22594,N_20525);
nand UO_2625 (O_2625,N_20849,N_24454);
and UO_2626 (O_2626,N_22005,N_24663);
nor UO_2627 (O_2627,N_22427,N_23403);
or UO_2628 (O_2628,N_20366,N_22933);
nand UO_2629 (O_2629,N_23163,N_22963);
nand UO_2630 (O_2630,N_22512,N_24608);
or UO_2631 (O_2631,N_23397,N_23339);
nand UO_2632 (O_2632,N_24207,N_23959);
nand UO_2633 (O_2633,N_24943,N_24869);
nand UO_2634 (O_2634,N_23193,N_22836);
nand UO_2635 (O_2635,N_22272,N_24365);
nor UO_2636 (O_2636,N_20104,N_23538);
nand UO_2637 (O_2637,N_22788,N_21030);
or UO_2638 (O_2638,N_23827,N_24652);
and UO_2639 (O_2639,N_21704,N_22496);
nand UO_2640 (O_2640,N_22067,N_21139);
nand UO_2641 (O_2641,N_23811,N_21223);
and UO_2642 (O_2642,N_24165,N_22373);
nand UO_2643 (O_2643,N_22070,N_23894);
or UO_2644 (O_2644,N_22963,N_21911);
xnor UO_2645 (O_2645,N_23303,N_20998);
nor UO_2646 (O_2646,N_22449,N_22623);
and UO_2647 (O_2647,N_22935,N_22367);
nand UO_2648 (O_2648,N_20330,N_21557);
nor UO_2649 (O_2649,N_24698,N_24636);
nand UO_2650 (O_2650,N_23371,N_24100);
or UO_2651 (O_2651,N_24514,N_23687);
nand UO_2652 (O_2652,N_20916,N_22551);
nor UO_2653 (O_2653,N_23809,N_24566);
or UO_2654 (O_2654,N_23387,N_21667);
and UO_2655 (O_2655,N_24725,N_24683);
and UO_2656 (O_2656,N_21415,N_21159);
xor UO_2657 (O_2657,N_23702,N_24490);
or UO_2658 (O_2658,N_20465,N_23065);
or UO_2659 (O_2659,N_22923,N_22715);
or UO_2660 (O_2660,N_22615,N_21958);
nor UO_2661 (O_2661,N_24579,N_21258);
and UO_2662 (O_2662,N_22675,N_23812);
and UO_2663 (O_2663,N_23192,N_22952);
nand UO_2664 (O_2664,N_22263,N_20128);
and UO_2665 (O_2665,N_21002,N_24163);
nand UO_2666 (O_2666,N_23136,N_21062);
and UO_2667 (O_2667,N_21450,N_22692);
or UO_2668 (O_2668,N_21668,N_24735);
nor UO_2669 (O_2669,N_21023,N_23471);
xor UO_2670 (O_2670,N_24911,N_24631);
or UO_2671 (O_2671,N_21620,N_23070);
or UO_2672 (O_2672,N_23801,N_20259);
nor UO_2673 (O_2673,N_21945,N_20666);
and UO_2674 (O_2674,N_23497,N_24325);
or UO_2675 (O_2675,N_24368,N_24363);
nand UO_2676 (O_2676,N_24362,N_22491);
or UO_2677 (O_2677,N_24190,N_22233);
nor UO_2678 (O_2678,N_22682,N_21423);
and UO_2679 (O_2679,N_20240,N_21609);
or UO_2680 (O_2680,N_21486,N_22374);
and UO_2681 (O_2681,N_20148,N_24312);
nand UO_2682 (O_2682,N_24054,N_21180);
or UO_2683 (O_2683,N_23370,N_20345);
nor UO_2684 (O_2684,N_24857,N_23309);
or UO_2685 (O_2685,N_21899,N_20252);
nor UO_2686 (O_2686,N_21162,N_23780);
and UO_2687 (O_2687,N_22887,N_23148);
xnor UO_2688 (O_2688,N_23163,N_24347);
nor UO_2689 (O_2689,N_21194,N_22870);
nand UO_2690 (O_2690,N_20396,N_23963);
nand UO_2691 (O_2691,N_23602,N_24436);
nand UO_2692 (O_2692,N_20147,N_22921);
and UO_2693 (O_2693,N_21655,N_21519);
nand UO_2694 (O_2694,N_24501,N_21750);
or UO_2695 (O_2695,N_22445,N_20076);
nor UO_2696 (O_2696,N_20745,N_23874);
or UO_2697 (O_2697,N_23477,N_21068);
nor UO_2698 (O_2698,N_22962,N_21609);
nand UO_2699 (O_2699,N_20003,N_22917);
or UO_2700 (O_2700,N_21115,N_20155);
xnor UO_2701 (O_2701,N_21397,N_23856);
nor UO_2702 (O_2702,N_21017,N_23087);
or UO_2703 (O_2703,N_21780,N_20901);
xnor UO_2704 (O_2704,N_20954,N_24355);
nor UO_2705 (O_2705,N_22389,N_20774);
nand UO_2706 (O_2706,N_20132,N_23137);
nor UO_2707 (O_2707,N_24834,N_22413);
nor UO_2708 (O_2708,N_23187,N_22220);
nand UO_2709 (O_2709,N_20917,N_20769);
nor UO_2710 (O_2710,N_20972,N_22345);
and UO_2711 (O_2711,N_20078,N_23277);
or UO_2712 (O_2712,N_24519,N_21535);
xnor UO_2713 (O_2713,N_20633,N_21677);
and UO_2714 (O_2714,N_20404,N_22252);
or UO_2715 (O_2715,N_24547,N_22023);
nor UO_2716 (O_2716,N_23508,N_23002);
and UO_2717 (O_2717,N_20776,N_21448);
or UO_2718 (O_2718,N_22337,N_23169);
nand UO_2719 (O_2719,N_24475,N_24363);
nor UO_2720 (O_2720,N_20337,N_23374);
nor UO_2721 (O_2721,N_23829,N_21077);
nand UO_2722 (O_2722,N_22350,N_24762);
and UO_2723 (O_2723,N_21334,N_22894);
nor UO_2724 (O_2724,N_23455,N_20196);
or UO_2725 (O_2725,N_24847,N_22261);
or UO_2726 (O_2726,N_20635,N_24026);
nand UO_2727 (O_2727,N_23678,N_22743);
and UO_2728 (O_2728,N_22340,N_20864);
and UO_2729 (O_2729,N_22094,N_21547);
and UO_2730 (O_2730,N_22718,N_20487);
nand UO_2731 (O_2731,N_24511,N_20648);
or UO_2732 (O_2732,N_20797,N_23394);
nor UO_2733 (O_2733,N_21139,N_21987);
or UO_2734 (O_2734,N_21992,N_21596);
or UO_2735 (O_2735,N_22449,N_20219);
nand UO_2736 (O_2736,N_22434,N_24797);
nor UO_2737 (O_2737,N_21069,N_23795);
or UO_2738 (O_2738,N_22763,N_21167);
nor UO_2739 (O_2739,N_23606,N_22895);
nand UO_2740 (O_2740,N_21116,N_20189);
or UO_2741 (O_2741,N_23290,N_20198);
and UO_2742 (O_2742,N_22674,N_23416);
nor UO_2743 (O_2743,N_24510,N_23115);
xnor UO_2744 (O_2744,N_21983,N_22155);
nand UO_2745 (O_2745,N_24907,N_20160);
and UO_2746 (O_2746,N_20571,N_22686);
nor UO_2747 (O_2747,N_22837,N_21238);
or UO_2748 (O_2748,N_24090,N_23887);
nor UO_2749 (O_2749,N_23154,N_23248);
nand UO_2750 (O_2750,N_20650,N_22757);
nand UO_2751 (O_2751,N_20079,N_24175);
or UO_2752 (O_2752,N_24467,N_23596);
nand UO_2753 (O_2753,N_21365,N_20743);
nand UO_2754 (O_2754,N_21426,N_21948);
and UO_2755 (O_2755,N_24470,N_24399);
xnor UO_2756 (O_2756,N_20343,N_22803);
nor UO_2757 (O_2757,N_21566,N_24401);
or UO_2758 (O_2758,N_23485,N_21717);
or UO_2759 (O_2759,N_21138,N_23059);
and UO_2760 (O_2760,N_20576,N_23426);
or UO_2761 (O_2761,N_24765,N_21759);
nand UO_2762 (O_2762,N_24697,N_20561);
or UO_2763 (O_2763,N_22145,N_22153);
and UO_2764 (O_2764,N_22798,N_22953);
nor UO_2765 (O_2765,N_21966,N_21821);
nor UO_2766 (O_2766,N_20519,N_20375);
and UO_2767 (O_2767,N_22063,N_20562);
nor UO_2768 (O_2768,N_23690,N_22407);
nand UO_2769 (O_2769,N_24501,N_21357);
xnor UO_2770 (O_2770,N_23796,N_24785);
or UO_2771 (O_2771,N_21661,N_23718);
and UO_2772 (O_2772,N_23476,N_20155);
nand UO_2773 (O_2773,N_21883,N_20660);
or UO_2774 (O_2774,N_20443,N_21147);
and UO_2775 (O_2775,N_22497,N_21358);
nor UO_2776 (O_2776,N_20049,N_24344);
nor UO_2777 (O_2777,N_23972,N_23099);
nand UO_2778 (O_2778,N_20858,N_22179);
and UO_2779 (O_2779,N_22459,N_22163);
nand UO_2780 (O_2780,N_23312,N_22475);
nor UO_2781 (O_2781,N_21445,N_23995);
nand UO_2782 (O_2782,N_21849,N_22579);
and UO_2783 (O_2783,N_24606,N_23789);
xor UO_2784 (O_2784,N_23719,N_22161);
nand UO_2785 (O_2785,N_20379,N_20626);
or UO_2786 (O_2786,N_24163,N_23386);
or UO_2787 (O_2787,N_21003,N_23913);
and UO_2788 (O_2788,N_21961,N_24974);
and UO_2789 (O_2789,N_22793,N_24126);
or UO_2790 (O_2790,N_21291,N_24368);
nand UO_2791 (O_2791,N_21921,N_20093);
nor UO_2792 (O_2792,N_24418,N_24592);
nand UO_2793 (O_2793,N_24641,N_22250);
nor UO_2794 (O_2794,N_20545,N_24449);
nor UO_2795 (O_2795,N_21477,N_24263);
nand UO_2796 (O_2796,N_22147,N_20305);
and UO_2797 (O_2797,N_20655,N_20427);
nand UO_2798 (O_2798,N_22639,N_21576);
or UO_2799 (O_2799,N_24680,N_23147);
or UO_2800 (O_2800,N_21499,N_24069);
and UO_2801 (O_2801,N_24564,N_22025);
nor UO_2802 (O_2802,N_24411,N_23203);
nor UO_2803 (O_2803,N_22344,N_21011);
nand UO_2804 (O_2804,N_21532,N_22288);
or UO_2805 (O_2805,N_24964,N_24533);
nand UO_2806 (O_2806,N_20042,N_23616);
nor UO_2807 (O_2807,N_22394,N_20378);
nand UO_2808 (O_2808,N_21503,N_22430);
nor UO_2809 (O_2809,N_21943,N_22364);
nand UO_2810 (O_2810,N_22749,N_20711);
and UO_2811 (O_2811,N_22275,N_20371);
xor UO_2812 (O_2812,N_21693,N_23370);
nand UO_2813 (O_2813,N_22078,N_23659);
nor UO_2814 (O_2814,N_24998,N_24775);
and UO_2815 (O_2815,N_21335,N_23882);
nor UO_2816 (O_2816,N_23263,N_24016);
and UO_2817 (O_2817,N_22834,N_23436);
or UO_2818 (O_2818,N_23361,N_24536);
and UO_2819 (O_2819,N_20681,N_21592);
nor UO_2820 (O_2820,N_24514,N_21346);
nor UO_2821 (O_2821,N_22581,N_20776);
or UO_2822 (O_2822,N_21291,N_24793);
and UO_2823 (O_2823,N_20353,N_22114);
nand UO_2824 (O_2824,N_23696,N_23384);
or UO_2825 (O_2825,N_24318,N_22630);
and UO_2826 (O_2826,N_21338,N_20174);
nor UO_2827 (O_2827,N_23273,N_21464);
nor UO_2828 (O_2828,N_24324,N_21957);
nand UO_2829 (O_2829,N_24146,N_21751);
or UO_2830 (O_2830,N_20376,N_22767);
nor UO_2831 (O_2831,N_24080,N_21488);
or UO_2832 (O_2832,N_23346,N_24518);
nor UO_2833 (O_2833,N_22320,N_23549);
nor UO_2834 (O_2834,N_20757,N_22726);
nor UO_2835 (O_2835,N_23405,N_20367);
or UO_2836 (O_2836,N_24461,N_23987);
or UO_2837 (O_2837,N_22357,N_22092);
nand UO_2838 (O_2838,N_20089,N_23711);
or UO_2839 (O_2839,N_24860,N_23093);
and UO_2840 (O_2840,N_21596,N_23525);
nor UO_2841 (O_2841,N_22272,N_24194);
and UO_2842 (O_2842,N_20942,N_24961);
and UO_2843 (O_2843,N_21704,N_22949);
nand UO_2844 (O_2844,N_22364,N_24648);
nor UO_2845 (O_2845,N_23082,N_24322);
and UO_2846 (O_2846,N_20928,N_24511);
nand UO_2847 (O_2847,N_21770,N_22527);
and UO_2848 (O_2848,N_20016,N_20642);
nand UO_2849 (O_2849,N_23652,N_22165);
and UO_2850 (O_2850,N_20848,N_22124);
and UO_2851 (O_2851,N_23897,N_21516);
nor UO_2852 (O_2852,N_24860,N_23982);
nand UO_2853 (O_2853,N_22153,N_20732);
and UO_2854 (O_2854,N_23466,N_24486);
and UO_2855 (O_2855,N_22487,N_22068);
or UO_2856 (O_2856,N_20047,N_24444);
nor UO_2857 (O_2857,N_20567,N_24517);
nor UO_2858 (O_2858,N_22305,N_21962);
nor UO_2859 (O_2859,N_24180,N_20819);
or UO_2860 (O_2860,N_23357,N_23475);
nand UO_2861 (O_2861,N_24929,N_23802);
and UO_2862 (O_2862,N_24065,N_20716);
nand UO_2863 (O_2863,N_20126,N_20346);
nor UO_2864 (O_2864,N_22935,N_23500);
nor UO_2865 (O_2865,N_21432,N_20748);
xor UO_2866 (O_2866,N_20897,N_24150);
nor UO_2867 (O_2867,N_20662,N_24748);
nand UO_2868 (O_2868,N_20516,N_24779);
or UO_2869 (O_2869,N_20465,N_22574);
and UO_2870 (O_2870,N_23527,N_23832);
and UO_2871 (O_2871,N_23663,N_24527);
nor UO_2872 (O_2872,N_20907,N_21824);
xor UO_2873 (O_2873,N_20485,N_24918);
and UO_2874 (O_2874,N_20550,N_22370);
and UO_2875 (O_2875,N_23463,N_22483);
xor UO_2876 (O_2876,N_21688,N_21352);
nand UO_2877 (O_2877,N_24347,N_23448);
and UO_2878 (O_2878,N_22348,N_20567);
and UO_2879 (O_2879,N_20092,N_22741);
nor UO_2880 (O_2880,N_24905,N_21329);
nor UO_2881 (O_2881,N_22594,N_23503);
xnor UO_2882 (O_2882,N_23563,N_23635);
nor UO_2883 (O_2883,N_23985,N_24512);
nand UO_2884 (O_2884,N_24075,N_22709);
and UO_2885 (O_2885,N_22674,N_21490);
or UO_2886 (O_2886,N_21122,N_24203);
nand UO_2887 (O_2887,N_22858,N_20412);
and UO_2888 (O_2888,N_22640,N_24440);
or UO_2889 (O_2889,N_20133,N_24684);
nand UO_2890 (O_2890,N_20375,N_23541);
nor UO_2891 (O_2891,N_21411,N_21799);
nor UO_2892 (O_2892,N_20501,N_23240);
or UO_2893 (O_2893,N_23703,N_20992);
or UO_2894 (O_2894,N_23080,N_20833);
or UO_2895 (O_2895,N_24000,N_23454);
nor UO_2896 (O_2896,N_23029,N_24817);
nand UO_2897 (O_2897,N_24792,N_23647);
or UO_2898 (O_2898,N_23356,N_21117);
nor UO_2899 (O_2899,N_24599,N_20852);
nand UO_2900 (O_2900,N_23572,N_24193);
nor UO_2901 (O_2901,N_21624,N_21683);
nor UO_2902 (O_2902,N_23504,N_20257);
or UO_2903 (O_2903,N_21718,N_21552);
and UO_2904 (O_2904,N_20881,N_22742);
or UO_2905 (O_2905,N_23841,N_20711);
and UO_2906 (O_2906,N_21271,N_23161);
and UO_2907 (O_2907,N_22798,N_22786);
or UO_2908 (O_2908,N_20883,N_22658);
and UO_2909 (O_2909,N_20910,N_24215);
or UO_2910 (O_2910,N_23105,N_20099);
nand UO_2911 (O_2911,N_24874,N_21404);
and UO_2912 (O_2912,N_22841,N_21549);
or UO_2913 (O_2913,N_23623,N_23222);
and UO_2914 (O_2914,N_21948,N_23213);
or UO_2915 (O_2915,N_20959,N_22411);
nor UO_2916 (O_2916,N_20089,N_22339);
and UO_2917 (O_2917,N_21060,N_21047);
or UO_2918 (O_2918,N_23365,N_21133);
nor UO_2919 (O_2919,N_22655,N_24233);
nand UO_2920 (O_2920,N_21503,N_21925);
or UO_2921 (O_2921,N_20256,N_24180);
or UO_2922 (O_2922,N_24689,N_23809);
nor UO_2923 (O_2923,N_23382,N_23418);
nor UO_2924 (O_2924,N_24957,N_23721);
nor UO_2925 (O_2925,N_22907,N_24031);
nor UO_2926 (O_2926,N_20840,N_20926);
nand UO_2927 (O_2927,N_21066,N_23131);
and UO_2928 (O_2928,N_20097,N_24785);
nand UO_2929 (O_2929,N_21143,N_20972);
nand UO_2930 (O_2930,N_24118,N_22175);
and UO_2931 (O_2931,N_20633,N_20395);
and UO_2932 (O_2932,N_20523,N_22208);
and UO_2933 (O_2933,N_22244,N_22271);
or UO_2934 (O_2934,N_22622,N_24154);
and UO_2935 (O_2935,N_23123,N_24933);
and UO_2936 (O_2936,N_22915,N_24652);
nand UO_2937 (O_2937,N_24967,N_23325);
nand UO_2938 (O_2938,N_20649,N_20378);
and UO_2939 (O_2939,N_21907,N_23203);
or UO_2940 (O_2940,N_20092,N_20264);
or UO_2941 (O_2941,N_21837,N_21276);
nor UO_2942 (O_2942,N_24263,N_21874);
and UO_2943 (O_2943,N_21893,N_20300);
and UO_2944 (O_2944,N_21184,N_24047);
or UO_2945 (O_2945,N_22230,N_21962);
nor UO_2946 (O_2946,N_20823,N_20118);
and UO_2947 (O_2947,N_24784,N_21788);
nand UO_2948 (O_2948,N_22956,N_21420);
and UO_2949 (O_2949,N_21788,N_23383);
or UO_2950 (O_2950,N_22213,N_22506);
nor UO_2951 (O_2951,N_20411,N_22835);
or UO_2952 (O_2952,N_20902,N_23584);
or UO_2953 (O_2953,N_21996,N_21141);
nor UO_2954 (O_2954,N_21338,N_22891);
nor UO_2955 (O_2955,N_21252,N_21268);
nor UO_2956 (O_2956,N_23598,N_23323);
and UO_2957 (O_2957,N_23848,N_22443);
or UO_2958 (O_2958,N_24715,N_22432);
nand UO_2959 (O_2959,N_21676,N_21354);
and UO_2960 (O_2960,N_23234,N_20890);
nand UO_2961 (O_2961,N_20647,N_21624);
or UO_2962 (O_2962,N_20577,N_24512);
nor UO_2963 (O_2963,N_24993,N_24209);
nor UO_2964 (O_2964,N_24958,N_24218);
nor UO_2965 (O_2965,N_24462,N_24216);
and UO_2966 (O_2966,N_21508,N_22119);
nand UO_2967 (O_2967,N_22042,N_20848);
nor UO_2968 (O_2968,N_20625,N_20263);
or UO_2969 (O_2969,N_23858,N_20954);
nand UO_2970 (O_2970,N_24303,N_20831);
nand UO_2971 (O_2971,N_24579,N_23929);
nor UO_2972 (O_2972,N_20320,N_21805);
nand UO_2973 (O_2973,N_21461,N_23091);
or UO_2974 (O_2974,N_20088,N_21332);
nand UO_2975 (O_2975,N_21888,N_22310);
and UO_2976 (O_2976,N_20527,N_21116);
nor UO_2977 (O_2977,N_22186,N_22455);
nor UO_2978 (O_2978,N_21681,N_22005);
and UO_2979 (O_2979,N_21314,N_20230);
or UO_2980 (O_2980,N_21983,N_23444);
nand UO_2981 (O_2981,N_21520,N_22236);
or UO_2982 (O_2982,N_23817,N_20296);
nor UO_2983 (O_2983,N_22862,N_23587);
nor UO_2984 (O_2984,N_22141,N_21482);
and UO_2985 (O_2985,N_21158,N_20065);
nand UO_2986 (O_2986,N_20545,N_20780);
nand UO_2987 (O_2987,N_20172,N_21041);
nor UO_2988 (O_2988,N_22646,N_22591);
nor UO_2989 (O_2989,N_24255,N_22160);
nand UO_2990 (O_2990,N_22597,N_22843);
nor UO_2991 (O_2991,N_24689,N_21696);
nor UO_2992 (O_2992,N_20868,N_20195);
nor UO_2993 (O_2993,N_24493,N_21175);
nand UO_2994 (O_2994,N_23183,N_22749);
or UO_2995 (O_2995,N_22441,N_23346);
and UO_2996 (O_2996,N_22171,N_20843);
and UO_2997 (O_2997,N_20037,N_20239);
or UO_2998 (O_2998,N_21054,N_21795);
nor UO_2999 (O_2999,N_20072,N_22737);
endmodule