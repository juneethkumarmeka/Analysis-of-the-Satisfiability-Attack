module basic_2500_25000_3000_8_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1141,In_2460);
nand U1 (N_1,In_1093,In_575);
nor U2 (N_2,In_1107,In_797);
or U3 (N_3,In_541,In_4);
xnor U4 (N_4,In_2334,In_1285);
nor U5 (N_5,In_2445,In_66);
and U6 (N_6,In_1371,In_1822);
nor U7 (N_7,In_565,In_1769);
nor U8 (N_8,In_266,In_519);
or U9 (N_9,In_453,In_2236);
nand U10 (N_10,In_544,In_919);
or U11 (N_11,In_1132,In_631);
nor U12 (N_12,In_480,In_2486);
nor U13 (N_13,In_786,In_621);
and U14 (N_14,In_2181,In_2462);
or U15 (N_15,In_1852,In_1147);
and U16 (N_16,In_2169,In_1097);
nand U17 (N_17,In_1414,In_2069);
and U18 (N_18,In_1581,In_2484);
or U19 (N_19,In_1816,In_433);
nand U20 (N_20,In_1508,In_1880);
and U21 (N_21,In_1191,In_1441);
or U22 (N_22,In_1905,In_1194);
or U23 (N_23,In_1864,In_496);
nor U24 (N_24,In_1545,In_1682);
nor U25 (N_25,In_304,In_1683);
xnor U26 (N_26,In_1134,In_2367);
and U27 (N_27,In_2386,In_1224);
and U28 (N_28,In_398,In_721);
nand U29 (N_29,In_1247,In_883);
xnor U30 (N_30,In_2320,In_975);
nor U31 (N_31,In_1321,In_1150);
and U32 (N_32,In_185,In_1961);
xor U33 (N_33,In_1201,In_2120);
and U34 (N_34,In_657,In_133);
nand U35 (N_35,In_8,In_684);
and U36 (N_36,In_1832,In_1317);
and U37 (N_37,In_638,In_1050);
and U38 (N_38,In_1466,In_2318);
or U39 (N_39,In_2332,In_973);
and U40 (N_40,In_2251,In_481);
nand U41 (N_41,In_1989,In_1451);
nor U42 (N_42,In_2263,In_978);
and U43 (N_43,In_417,In_220);
nand U44 (N_44,In_92,In_193);
and U45 (N_45,In_2047,In_1155);
and U46 (N_46,In_1084,In_929);
or U47 (N_47,In_1969,In_853);
nand U48 (N_48,In_1206,In_998);
nand U49 (N_49,In_891,In_1916);
and U50 (N_50,In_600,In_188);
nor U51 (N_51,In_892,In_1018);
or U52 (N_52,In_1073,In_831);
xor U53 (N_53,In_1721,In_1300);
xor U54 (N_54,In_1697,In_1533);
nor U55 (N_55,In_1437,In_2117);
xor U56 (N_56,In_202,In_869);
nor U57 (N_57,In_1921,In_2452);
or U58 (N_58,In_1372,In_1177);
or U59 (N_59,In_830,In_297);
and U60 (N_60,In_817,In_1641);
nand U61 (N_61,In_767,In_400);
and U62 (N_62,In_347,In_1216);
nor U63 (N_63,In_2275,In_1282);
nand U64 (N_64,In_1516,In_597);
nor U65 (N_65,In_312,In_1014);
nand U66 (N_66,In_834,In_2267);
or U67 (N_67,In_844,In_1502);
nand U68 (N_68,In_695,In_2076);
or U69 (N_69,In_840,In_2158);
and U70 (N_70,In_2284,In_1395);
or U71 (N_71,In_261,In_1814);
nor U72 (N_72,In_1311,In_611);
nand U73 (N_73,In_812,In_1857);
xor U74 (N_74,In_293,In_149);
nor U75 (N_75,In_619,In_582);
nand U76 (N_76,In_1181,In_635);
xor U77 (N_77,In_1917,In_1529);
xor U78 (N_78,In_518,In_1657);
nand U79 (N_79,In_2326,In_2212);
nor U80 (N_80,In_332,In_1075);
nor U81 (N_81,In_1166,In_663);
nor U82 (N_82,In_2388,In_1910);
nand U83 (N_83,In_2115,In_2430);
nand U84 (N_84,In_2382,In_1861);
nor U85 (N_85,In_86,In_445);
nand U86 (N_86,In_160,In_172);
nor U87 (N_87,In_52,In_1557);
xor U88 (N_88,In_1526,In_1101);
nand U89 (N_89,In_2059,In_1066);
xor U90 (N_90,In_1031,In_706);
and U91 (N_91,In_1779,In_1784);
and U92 (N_92,In_1119,In_2232);
and U93 (N_93,In_1870,In_738);
nand U94 (N_94,In_1777,In_615);
or U95 (N_95,In_2258,In_241);
or U96 (N_96,In_311,In_879);
and U97 (N_97,In_406,In_2277);
nand U98 (N_98,In_1500,In_557);
and U99 (N_99,In_1251,In_948);
nand U100 (N_100,In_1030,In_1479);
nand U101 (N_101,In_321,In_119);
nor U102 (N_102,In_934,In_677);
nor U103 (N_103,In_1047,In_871);
and U104 (N_104,In_2434,In_1692);
xnor U105 (N_105,In_1994,In_1045);
xnor U106 (N_106,In_1358,In_803);
xor U107 (N_107,In_932,In_302);
nand U108 (N_108,In_2215,In_906);
and U109 (N_109,In_1923,In_1320);
nor U110 (N_110,In_191,In_2003);
xor U111 (N_111,In_2216,In_753);
xnor U112 (N_112,In_1696,In_789);
nor U113 (N_113,In_1123,In_171);
nand U114 (N_114,In_2057,In_654);
nand U115 (N_115,In_1106,In_2202);
nor U116 (N_116,In_1405,In_378);
nand U117 (N_117,In_1912,In_2444);
nor U118 (N_118,In_1408,In_670);
or U119 (N_119,In_130,In_2105);
nand U120 (N_120,In_1620,In_1716);
nor U121 (N_121,In_128,In_151);
or U122 (N_122,In_144,In_2393);
and U123 (N_123,In_1310,In_751);
and U124 (N_124,In_2193,In_1749);
or U125 (N_125,In_1801,In_605);
or U126 (N_126,In_1977,In_970);
and U127 (N_127,In_959,In_1077);
nor U128 (N_128,In_874,In_5);
xnor U129 (N_129,In_1867,In_2234);
nor U130 (N_130,In_181,In_1443);
or U131 (N_131,In_1681,In_2276);
xor U132 (N_132,In_1088,In_554);
xor U133 (N_133,In_1950,In_1274);
nor U134 (N_134,In_2458,In_1722);
nand U135 (N_135,In_2361,In_105);
nor U136 (N_136,In_1347,In_1660);
or U137 (N_137,In_2199,In_2294);
or U138 (N_138,In_2219,In_377);
nand U139 (N_139,In_32,In_1636);
or U140 (N_140,In_336,In_1809);
xor U141 (N_141,In_546,In_1256);
and U142 (N_142,In_2228,In_1403);
and U143 (N_143,In_1313,In_1780);
nand U144 (N_144,In_2079,In_2470);
nor U145 (N_145,In_758,In_584);
nor U146 (N_146,In_447,In_1860);
or U147 (N_147,In_1829,In_432);
and U148 (N_148,In_1118,In_419);
or U149 (N_149,In_68,In_1143);
nor U150 (N_150,In_1853,In_1968);
xnor U151 (N_151,In_1307,In_776);
and U152 (N_152,In_1028,In_1293);
or U153 (N_153,In_2131,In_2259);
or U154 (N_154,In_1919,In_2133);
and U155 (N_155,In_1599,In_2422);
or U156 (N_156,In_1691,In_2487);
nand U157 (N_157,In_2005,In_442);
nand U158 (N_158,In_647,In_1148);
nand U159 (N_159,In_2307,In_839);
nand U160 (N_160,In_774,In_2438);
nand U161 (N_161,In_153,In_972);
nand U162 (N_162,In_325,In_858);
or U163 (N_163,In_87,In_1944);
nor U164 (N_164,In_1512,In_2078);
nor U165 (N_165,In_381,In_250);
nand U166 (N_166,In_538,In_1505);
nand U167 (N_167,In_1808,In_1163);
nand U168 (N_168,In_1487,In_1035);
or U169 (N_169,In_334,In_612);
nand U170 (N_170,In_1607,In_324);
xor U171 (N_171,In_561,In_411);
nor U172 (N_172,In_2315,In_1671);
nand U173 (N_173,In_1621,In_529);
nor U174 (N_174,In_2223,In_995);
nor U175 (N_175,In_1810,In_748);
nand U176 (N_176,In_372,In_731);
nor U177 (N_177,In_507,In_762);
nor U178 (N_178,In_1708,In_2072);
or U179 (N_179,In_806,In_2190);
and U180 (N_180,In_796,In_484);
nor U181 (N_181,In_1773,In_1005);
nand U182 (N_182,In_1121,In_1334);
and U183 (N_183,In_2132,In_1985);
and U184 (N_184,In_1039,In_2139);
and U185 (N_185,In_268,In_2111);
and U186 (N_186,In_1850,In_1684);
nor U187 (N_187,In_2449,In_1930);
xor U188 (N_188,In_787,In_1903);
or U189 (N_189,In_364,In_1333);
and U190 (N_190,In_2207,In_2420);
or U191 (N_191,In_209,In_1764);
and U192 (N_192,In_1575,In_1878);
nand U193 (N_193,In_1927,In_2421);
and U194 (N_194,In_1459,In_2163);
and U195 (N_195,In_848,In_1315);
and U196 (N_196,In_989,In_1794);
or U197 (N_197,In_410,In_864);
or U198 (N_198,In_1149,In_264);
nor U199 (N_199,In_1913,In_1344);
xor U200 (N_200,In_520,In_1244);
nand U201 (N_201,In_2476,In_1125);
nor U202 (N_202,In_24,In_1133);
nand U203 (N_203,In_1411,In_1995);
and U204 (N_204,In_438,In_2363);
nand U205 (N_205,In_111,In_140);
nand U206 (N_206,In_2289,In_1021);
nand U207 (N_207,In_1770,In_687);
and U208 (N_208,In_843,In_1048);
or U209 (N_209,In_894,In_716);
or U210 (N_210,In_2092,In_627);
nor U211 (N_211,In_2292,In_1704);
nand U212 (N_212,In_623,In_389);
nand U213 (N_213,In_2376,In_614);
and U214 (N_214,In_986,In_965);
or U215 (N_215,In_613,In_1436);
nor U216 (N_216,In_847,In_1258);
nor U217 (N_217,In_388,In_788);
or U218 (N_218,In_2056,In_2210);
or U219 (N_219,In_11,In_963);
or U220 (N_220,In_1531,In_522);
xnor U221 (N_221,In_218,In_903);
or U222 (N_222,In_2359,In_54);
xnor U223 (N_223,In_1876,In_1378);
xor U224 (N_224,In_1953,In_1496);
xnor U225 (N_225,In_504,In_1335);
nor U226 (N_226,In_1171,In_977);
nor U227 (N_227,In_656,In_1992);
or U228 (N_228,In_6,In_1527);
and U229 (N_229,In_1362,In_2031);
nor U230 (N_230,In_644,In_2142);
or U231 (N_231,In_12,In_1643);
and U232 (N_232,In_307,In_2391);
nor U233 (N_233,In_350,In_120);
nor U234 (N_234,In_1830,In_1693);
xor U235 (N_235,In_808,In_490);
or U236 (N_236,In_2039,In_2340);
nor U237 (N_237,In_44,In_472);
or U238 (N_238,In_1834,In_882);
or U239 (N_239,In_158,In_1338);
or U240 (N_240,In_254,In_1615);
nand U241 (N_241,In_2002,In_435);
xor U242 (N_242,In_732,In_397);
and U243 (N_243,In_733,In_503);
or U244 (N_244,In_837,In_711);
nor U245 (N_245,In_327,In_1237);
nand U246 (N_246,In_65,In_370);
nor U247 (N_247,In_76,In_434);
and U248 (N_248,In_809,In_828);
xnor U249 (N_249,In_567,In_2036);
nor U250 (N_250,In_1614,In_1227);
and U251 (N_251,In_374,In_1042);
or U252 (N_252,In_1598,In_1115);
nand U253 (N_253,In_375,In_1129);
nand U254 (N_254,In_1986,In_2218);
nand U255 (N_255,In_2197,In_1036);
nand U256 (N_256,In_221,In_99);
or U257 (N_257,In_845,In_662);
nand U258 (N_258,In_1493,In_2488);
or U259 (N_259,In_1080,In_884);
nand U260 (N_260,In_1550,In_431);
or U261 (N_261,In_50,In_1145);
and U262 (N_262,In_1564,In_899);
nand U263 (N_263,In_1752,In_1078);
xor U264 (N_264,In_441,In_1477);
or U265 (N_265,In_1397,In_1924);
xnor U266 (N_266,In_1276,In_826);
or U267 (N_267,In_1561,In_1655);
nor U268 (N_268,In_1204,In_1745);
or U269 (N_269,In_1863,In_259);
nand U270 (N_270,In_835,In_147);
nor U271 (N_271,In_110,In_921);
nand U272 (N_272,In_1972,In_2186);
xnor U273 (N_273,In_590,In_1714);
or U274 (N_274,In_1698,In_1732);
or U275 (N_275,In_127,In_2113);
xor U276 (N_276,In_1492,In_1346);
nor U277 (N_277,In_90,In_1538);
nor U278 (N_278,In_1025,In_2203);
nor U279 (N_279,In_1065,In_1758);
nand U280 (N_280,In_1182,In_1580);
and U281 (N_281,In_1336,In_1393);
or U282 (N_282,In_1278,In_2125);
nor U283 (N_283,In_10,In_1109);
nor U284 (N_284,In_2364,In_1694);
or U285 (N_285,In_2052,In_1634);
nand U286 (N_286,In_1907,In_1011);
xor U287 (N_287,In_1006,In_1517);
or U288 (N_288,In_138,In_1153);
nor U289 (N_289,In_2074,In_1914);
or U290 (N_290,In_1983,In_560);
nor U291 (N_291,In_960,In_881);
and U292 (N_292,In_2129,In_2135);
nand U293 (N_293,In_669,In_1639);
or U294 (N_294,In_2295,In_1677);
nand U295 (N_295,In_1843,In_2008);
nor U296 (N_296,In_2040,In_904);
or U297 (N_297,In_428,In_857);
or U298 (N_298,In_274,In_326);
or U299 (N_299,In_498,In_1076);
and U300 (N_300,In_653,In_269);
nor U301 (N_301,In_2349,In_829);
xnor U302 (N_302,In_703,In_1043);
nor U303 (N_303,In_1130,In_705);
or U304 (N_304,In_2362,In_1246);
nand U305 (N_305,In_2335,In_1624);
or U306 (N_306,In_2415,In_280);
nand U307 (N_307,In_1528,In_512);
and U308 (N_308,In_1685,In_329);
or U309 (N_309,In_2402,In_2328);
or U310 (N_310,In_2245,In_2269);
or U311 (N_311,In_1128,In_2184);
and U312 (N_312,In_1546,In_1720);
nor U313 (N_313,In_562,In_1622);
and U314 (N_314,In_2222,In_1236);
nor U315 (N_315,In_107,In_2384);
nor U316 (N_316,In_271,In_887);
xor U317 (N_317,In_992,In_1603);
or U318 (N_318,In_1859,In_1602);
and U319 (N_319,In_1175,In_984);
nor U320 (N_320,In_2073,In_942);
and U321 (N_321,In_1438,In_1595);
and U322 (N_322,In_1690,In_198);
xor U323 (N_323,In_543,In_523);
nand U324 (N_324,In_2042,In_1753);
nor U325 (N_325,In_211,In_2370);
or U326 (N_326,In_1284,In_466);
nor U327 (N_327,In_1209,In_730);
or U328 (N_328,In_159,In_1458);
and U329 (N_329,In_1900,In_230);
or U330 (N_330,In_1015,In_27);
and U331 (N_331,In_58,In_33);
xor U332 (N_332,In_1197,In_207);
and U333 (N_333,In_2427,In_527);
nor U334 (N_334,In_2271,In_102);
nor U335 (N_335,In_1488,In_1768);
and U336 (N_336,In_2435,In_1566);
nor U337 (N_337,In_1288,In_524);
xnor U338 (N_338,In_675,In_1886);
and U339 (N_339,In_9,In_1444);
and U340 (N_340,In_2217,In_1172);
or U341 (N_341,In_2439,In_2351);
and U342 (N_342,In_1824,In_176);
nor U343 (N_343,In_2225,In_1183);
nor U344 (N_344,In_1707,In_632);
nor U345 (N_345,In_1819,In_403);
and U346 (N_346,In_2165,In_1356);
nand U347 (N_347,In_2145,In_2424);
nand U348 (N_348,In_248,In_2397);
nor U349 (N_349,In_1180,In_777);
and U350 (N_350,In_219,In_573);
nor U351 (N_351,In_1427,In_448);
or U352 (N_352,In_1584,In_579);
nor U353 (N_353,In_2241,In_1261);
nor U354 (N_354,In_2214,In_1044);
or U355 (N_355,In_45,In_1243);
and U356 (N_356,In_616,In_1594);
nor U357 (N_357,In_486,In_604);
xnor U358 (N_358,In_455,In_1741);
or U359 (N_359,In_1901,In_1740);
nand U360 (N_360,In_1932,In_1999);
nand U361 (N_361,In_2020,In_2099);
nand U362 (N_362,In_810,In_1203);
or U363 (N_363,In_1,In_1793);
nor U364 (N_364,In_1471,In_1851);
or U365 (N_365,In_2230,In_2206);
and U366 (N_366,In_1349,In_310);
and U367 (N_367,In_862,In_69);
and U368 (N_368,In_72,In_578);
nor U369 (N_369,In_1926,In_1855);
or U370 (N_370,In_2301,In_1152);
nand U371 (N_371,In_2012,In_1790);
xnor U372 (N_372,In_689,In_569);
nor U373 (N_373,In_1124,In_1888);
or U374 (N_374,In_164,In_1316);
nor U375 (N_375,In_2119,In_933);
or U376 (N_376,In_399,In_1612);
nor U377 (N_377,In_1717,In_821);
xnor U378 (N_378,In_36,In_500);
nor U379 (N_379,In_1482,In_51);
xor U380 (N_380,In_229,In_1522);
xor U381 (N_381,In_1398,In_1198);
and U382 (N_382,In_2387,In_224);
or U383 (N_383,In_1448,In_234);
nor U384 (N_384,In_626,In_2455);
or U385 (N_385,In_1723,In_359);
nand U386 (N_386,In_938,In_426);
or U387 (N_387,In_1895,In_2338);
nor U388 (N_388,In_2242,In_768);
xnor U389 (N_389,In_540,In_1421);
nor U390 (N_390,In_896,In_80);
nor U391 (N_391,In_1844,In_1290);
nor U392 (N_392,In_1823,In_595);
nand U393 (N_393,In_2287,In_780);
nor U394 (N_394,In_1877,In_83);
or U395 (N_395,In_2423,In_1450);
or U396 (N_396,In_603,In_1331);
nand U397 (N_397,In_852,In_2088);
or U398 (N_398,In_1733,In_1611);
nor U399 (N_399,In_1007,In_1215);
nor U400 (N_400,In_1475,In_2446);
nand U401 (N_401,In_690,In_79);
or U402 (N_402,In_1235,In_449);
or U403 (N_403,In_673,In_439);
nor U404 (N_404,In_1280,In_1387);
nand U405 (N_405,In_2268,In_1009);
nor U406 (N_406,In_1573,In_210);
nor U407 (N_407,In_485,In_1666);
nand U408 (N_408,In_1756,In_637);
and U409 (N_409,In_1483,In_233);
or U410 (N_410,In_113,In_1956);
nand U411 (N_411,In_2454,In_1719);
or U412 (N_412,In_303,In_1559);
or U413 (N_413,In_2237,In_2380);
xor U414 (N_414,In_1783,In_1884);
nand U415 (N_415,In_1805,In_239);
or U416 (N_416,In_813,In_2442);
nor U417 (N_417,In_1640,In_784);
nand U418 (N_418,In_1178,In_328);
nor U419 (N_419,In_1254,In_517);
nand U420 (N_420,In_2265,In_949);
and U421 (N_421,In_1565,In_1645);
nand U422 (N_422,In_206,In_165);
nor U423 (N_423,In_888,In_1225);
and U424 (N_424,In_2379,In_1069);
nand U425 (N_425,In_1551,In_2086);
nor U426 (N_426,In_201,In_1579);
nor U427 (N_427,In_1665,In_947);
xor U428 (N_428,In_2306,In_1757);
and U429 (N_429,In_2481,In_1105);
nand U430 (N_430,In_976,In_982);
or U431 (N_431,In_1510,In_2483);
nor U432 (N_432,In_727,In_134);
or U433 (N_433,In_1457,In_953);
and U434 (N_434,In_1114,In_1485);
nand U435 (N_435,In_2479,In_1476);
nor U436 (N_436,In_686,In_1626);
nand U437 (N_437,In_2182,In_1951);
nand U438 (N_438,In_444,In_1499);
or U439 (N_439,In_1739,In_383);
xnor U440 (N_440,In_1102,In_1918);
nand U441 (N_441,In_1778,In_539);
nand U442 (N_442,In_2112,In_698);
and U443 (N_443,In_1200,In_1491);
nand U444 (N_444,In_1990,In_2024);
or U445 (N_445,In_2467,In_2026);
nor U446 (N_446,In_1894,In_1020);
nor U447 (N_447,In_2409,In_396);
nor U448 (N_448,In_674,In_408);
nor U449 (N_449,In_1937,In_999);
or U450 (N_450,In_1613,In_495);
and U451 (N_451,In_1882,In_1815);
nand U452 (N_452,In_118,In_2180);
nor U453 (N_453,In_1214,In_723);
nor U454 (N_454,In_296,In_2175);
or U455 (N_455,In_384,In_1373);
nand U456 (N_456,In_73,In_231);
and U457 (N_457,In_2231,In_436);
nand U458 (N_458,In_424,In_1041);
nand U459 (N_459,In_1792,In_1226);
nand U460 (N_460,In_1842,In_534);
or U461 (N_461,In_1319,In_2121);
and U462 (N_462,In_2095,In_1710);
and U463 (N_463,In_924,In_643);
xnor U464 (N_464,In_1137,In_2122);
nand U465 (N_465,In_474,In_1339);
or U466 (N_466,In_1889,In_1872);
nor U467 (N_467,In_2143,In_2308);
or U468 (N_468,In_2248,In_2336);
nor U469 (N_469,In_1649,In_1978);
or U470 (N_470,In_772,In_1954);
nor U471 (N_471,In_1418,In_1323);
and U472 (N_472,In_925,In_1841);
and U473 (N_473,In_1552,In_2281);
or U474 (N_474,In_2313,In_415);
and U475 (N_475,In_166,In_2344);
nand U476 (N_476,In_273,In_2100);
nor U477 (N_477,In_376,In_15);
or U478 (N_478,In_818,In_1211);
nand U479 (N_479,In_2495,In_779);
and U480 (N_480,In_850,In_2432);
and U481 (N_481,In_1068,In_1836);
nand U482 (N_482,In_1355,In_1383);
nand U483 (N_483,In_1473,In_680);
nor U484 (N_484,In_97,In_2262);
and U485 (N_485,In_1623,In_1498);
nand U486 (N_486,In_1117,In_648);
nand U487 (N_487,In_1578,In_2450);
and U488 (N_488,In_91,In_890);
nor U489 (N_489,In_671,In_2342);
or U490 (N_490,In_747,In_1588);
nor U491 (N_491,In_798,In_1385);
and U492 (N_492,In_290,In_1345);
nor U493 (N_493,In_2085,In_773);
nand U494 (N_494,In_494,In_1099);
nand U495 (N_495,In_822,In_2102);
or U496 (N_496,In_340,In_2065);
and U497 (N_497,In_263,In_2164);
nand U498 (N_498,In_1348,In_1965);
and U499 (N_499,In_170,In_257);
and U500 (N_500,In_1802,In_2372);
nor U501 (N_501,In_458,In_1273);
and U502 (N_502,In_2224,In_2461);
nor U503 (N_503,In_2323,In_710);
and U504 (N_504,In_593,In_2309);
and U505 (N_505,In_2192,In_1675);
nor U506 (N_506,In_591,In_2116);
nand U507 (N_507,In_1763,In_2463);
or U508 (N_508,In_104,In_926);
nand U509 (N_509,In_2201,In_694);
nand U510 (N_510,In_2451,In_2080);
or U511 (N_511,In_2136,In_1091);
xor U512 (N_512,In_2285,In_1154);
nor U513 (N_513,In_1825,In_479);
nand U514 (N_514,In_40,In_1388);
and U515 (N_515,In_1868,In_2290);
nor U516 (N_516,In_2166,In_470);
nand U517 (N_517,In_1052,In_2282);
or U518 (N_518,In_386,In_345);
nand U519 (N_519,In_1266,In_824);
xor U520 (N_520,In_736,In_1363);
or U521 (N_521,In_62,In_291);
nand U522 (N_522,In_719,In_1416);
and U523 (N_523,In_1727,In_1269);
nand U524 (N_524,In_962,In_2188);
nor U525 (N_525,In_1013,In_1017);
or U526 (N_526,In_2447,In_969);
nor U527 (N_527,In_742,In_1071);
and U528 (N_528,In_550,In_525);
and U529 (N_529,In_566,In_1332);
or U530 (N_530,In_761,In_936);
and U531 (N_531,In_279,In_1731);
xnor U532 (N_532,In_2110,In_1547);
or U533 (N_533,In_1667,In_2107);
xor U534 (N_534,In_749,In_1596);
nand U535 (N_535,In_2489,In_815);
nor U536 (N_536,In_1104,In_175);
nand U537 (N_537,In_782,In_2260);
nor U538 (N_538,In_407,In_849);
nor U539 (N_539,In_1548,In_1949);
nand U540 (N_540,In_1556,In_2345);
nor U541 (N_541,In_1424,In_287);
nor U542 (N_542,In_352,In_443);
and U543 (N_543,In_1661,In_868);
or U544 (N_544,In_1555,In_1299);
nand U545 (N_545,In_1159,In_391);
and U546 (N_546,In_1328,In_1838);
nor U547 (N_547,In_1688,In_851);
nand U548 (N_548,In_1997,In_260);
nor U549 (N_549,In_1432,In_88);
or U550 (N_550,In_288,In_1151);
nand U551 (N_551,In_775,In_870);
nand U552 (N_552,In_1952,In_2254);
nand U553 (N_553,In_1560,In_183);
nand U554 (N_554,In_401,In_577);
or U555 (N_555,In_1804,In_82);
xnor U556 (N_556,In_1002,In_395);
and U557 (N_557,In_1070,In_2325);
nor U558 (N_558,In_744,In_1798);
xor U559 (N_559,In_2302,In_1662);
and U560 (N_560,In_988,In_795);
and U561 (N_561,In_387,In_1423);
nor U562 (N_562,In_2399,In_1037);
nor U563 (N_563,In_1447,In_2288);
nor U564 (N_564,In_2303,In_2090);
xnor U565 (N_565,In_136,In_1360);
or U566 (N_566,In_954,In_1384);
xnor U567 (N_567,In_583,In_123);
nor U568 (N_568,In_380,In_900);
nor U569 (N_569,In_2272,In_57);
nand U570 (N_570,In_2235,In_2478);
nand U571 (N_571,In_2279,In_267);
and U572 (N_572,In_1748,In_2353);
nor U573 (N_573,In_1541,In_2398);
nand U574 (N_574,In_572,In_2273);
nor U575 (N_575,In_665,In_820);
and U576 (N_576,In_754,In_2494);
nor U577 (N_577,In_1652,In_510);
and U578 (N_578,In_1590,In_2050);
xnor U579 (N_579,In_2063,In_634);
nor U580 (N_580,In_964,In_60);
nand U581 (N_581,In_1286,In_2091);
or U582 (N_582,In_549,In_316);
xor U583 (N_583,In_412,In_1135);
nor U584 (N_584,In_179,In_1250);
and U585 (N_585,In_704,In_668);
and U586 (N_586,In_807,In_1314);
nand U587 (N_587,In_429,In_836);
nor U588 (N_588,In_1245,In_1298);
nor U589 (N_589,In_109,In_2060);
nand U590 (N_590,In_67,In_2466);
nand U591 (N_591,In_1605,In_1729);
xnor U592 (N_592,In_1539,In_1330);
or U593 (N_593,In_927,In_1521);
nor U594 (N_594,In_1160,In_169);
nand U595 (N_595,In_2441,In_679);
xnor U596 (N_596,In_1821,In_2352);
nor U597 (N_597,In_766,In_305);
xor U598 (N_598,In_141,In_366);
nand U599 (N_599,In_2298,In_1157);
and U600 (N_600,In_649,In_265);
nor U601 (N_601,In_1765,In_1908);
xor U602 (N_602,In_235,In_935);
or U603 (N_603,In_1343,In_1389);
or U604 (N_604,In_276,In_740);
and U605 (N_605,In_2493,In_2305);
and U606 (N_606,In_979,In_875);
and U607 (N_607,In_124,In_56);
nor U608 (N_608,In_2155,In_846);
nand U609 (N_609,In_1653,In_178);
nor U610 (N_610,In_84,In_2053);
nand U611 (N_611,In_2173,In_2067);
nor U612 (N_612,In_955,In_96);
or U613 (N_613,In_951,In_2213);
nor U614 (N_614,In_1629,In_94);
nor U615 (N_615,In_588,In_2436);
or U616 (N_616,In_2373,In_1567);
or U617 (N_617,In_1279,In_1987);
and U618 (N_618,In_245,In_2);
nand U619 (N_619,In_190,In_1647);
nand U620 (N_620,In_363,In_1023);
and U621 (N_621,In_2071,In_1220);
nor U622 (N_622,In_1518,In_1947);
nand U623 (N_623,In_755,In_683);
nor U624 (N_624,In_46,In_162);
nand U625 (N_625,In_2239,In_283);
or U626 (N_626,In_1658,In_945);
nor U627 (N_627,In_1813,In_157);
or U628 (N_628,In_2319,In_2474);
or U629 (N_629,In_2001,In_791);
nor U630 (N_630,In_369,In_790);
xor U631 (N_631,In_2106,In_912);
nand U632 (N_632,In_95,In_404);
or U633 (N_633,In_2428,In_101);
nand U634 (N_634,In_14,In_1396);
or U635 (N_635,In_2459,In_1938);
xnor U636 (N_636,In_2138,In_1353);
or U637 (N_637,In_2000,In_536);
or U638 (N_638,In_1656,In_1267);
nand U639 (N_639,In_473,In_353);
xor U640 (N_640,In_2425,In_696);
nand U641 (N_641,In_708,In_532);
and U642 (N_642,In_2149,In_342);
and U643 (N_643,In_1301,In_462);
nand U644 (N_644,In_620,In_664);
nor U645 (N_645,In_1608,In_1000);
and U646 (N_646,In_651,In_1369);
nand U647 (N_647,In_351,In_1663);
nand U648 (N_648,In_1484,In_240);
nor U649 (N_649,In_2278,In_349);
nor U650 (N_650,In_2198,In_1379);
or U651 (N_651,In_1352,In_1775);
and U652 (N_652,In_692,In_2126);
nor U653 (N_653,In_1571,In_1957);
and U654 (N_654,In_156,In_1817);
and U655 (N_655,In_701,In_1127);
or U656 (N_656,In_1295,In_1359);
or U657 (N_657,In_242,In_1828);
and U658 (N_658,In_939,In_2286);
nand U659 (N_659,In_385,In_196);
and U660 (N_660,In_1260,In_2167);
nor U661 (N_661,In_922,In_1158);
or U662 (N_662,In_535,In_901);
xor U663 (N_663,In_2153,In_1094);
or U664 (N_664,In_322,In_1399);
nand U665 (N_665,In_1231,In_1188);
nand U666 (N_666,In_528,In_1839);
nand U667 (N_667,In_1616,In_393);
nor U668 (N_668,In_576,In_2310);
xor U669 (N_669,In_639,In_1059);
nor U670 (N_670,In_355,In_1281);
or U671 (N_671,In_317,In_1929);
nor U672 (N_672,In_460,In_1701);
nor U673 (N_673,In_1664,In_1292);
nand U674 (N_674,In_2497,In_2061);
or U675 (N_675,In_1169,In_1193);
xnor U676 (N_676,In_707,In_1381);
nor U677 (N_677,In_475,In_854);
nor U678 (N_678,In_915,In_2150);
nor U679 (N_679,In_477,In_137);
and U680 (N_680,In_2498,In_1846);
or U681 (N_681,In_1219,In_2485);
or U682 (N_682,In_1390,In_2070);
nor U683 (N_683,In_917,In_771);
or U684 (N_684,In_1920,In_610);
nand U685 (N_685,In_1646,In_476);
nand U686 (N_686,In_770,In_139);
and U687 (N_687,In_493,In_1087);
and U688 (N_688,In_941,In_599);
or U689 (N_689,In_100,In_2041);
nand U690 (N_690,In_1980,In_2027);
or U691 (N_691,In_1012,In_2331);
or U692 (N_692,In_1772,In_114);
nand U693 (N_693,In_750,In_1144);
nor U694 (N_694,In_301,In_1650);
xnor U695 (N_695,In_2366,In_1858);
nor U696 (N_696,In_1164,In_931);
nor U697 (N_697,In_1435,In_2097);
or U698 (N_698,In_1103,In_1079);
and U699 (N_699,In_1303,In_1271);
xnor U700 (N_700,In_1326,In_1807);
nand U701 (N_701,In_1361,In_63);
and U702 (N_702,In_1234,In_2037);
and U703 (N_703,In_2233,In_70);
nor U704 (N_704,In_1974,In_2337);
and U705 (N_705,In_1948,In_186);
and U706 (N_706,In_2087,In_197);
or U707 (N_707,In_1187,In_2141);
and U708 (N_708,In_1670,In_1811);
and U709 (N_709,In_1189,In_468);
nand U710 (N_710,In_1519,In_1883);
xor U711 (N_711,In_1536,In_1549);
nor U712 (N_712,In_1112,In_129);
and U713 (N_713,In_1966,In_1543);
nand U714 (N_714,In_29,In_1287);
nor U715 (N_715,In_2032,In_28);
or U716 (N_716,In_173,In_1507);
or U717 (N_717,In_38,In_2009);
nand U718 (N_718,In_2414,In_618);
nor U719 (N_719,In_47,In_390);
nand U720 (N_720,In_1309,In_878);
nor U721 (N_721,In_827,In_908);
nor U722 (N_722,In_2183,In_1933);
nand U723 (N_723,In_1981,In_285);
nor U724 (N_724,In_200,In_2118);
xnor U725 (N_725,In_2297,In_35);
or U726 (N_726,In_452,In_49);
xnor U727 (N_727,In_1167,In_804);
and U728 (N_728,In_421,In_379);
or U729 (N_729,In_559,In_420);
and U730 (N_730,In_189,In_658);
or U731 (N_731,In_1341,In_819);
nand U732 (N_732,In_1464,In_2226);
and U733 (N_733,In_2229,In_1840);
nor U734 (N_734,In_2051,In_1709);
xnor U735 (N_735,In_215,In_108);
or U736 (N_736,In_1871,In_34);
nor U737 (N_737,In_1376,In_7);
nand U738 (N_738,In_1506,In_1486);
and U739 (N_739,In_2179,In_1468);
and U740 (N_740,In_232,In_526);
nand U741 (N_741,In_885,In_1940);
or U742 (N_742,In_1744,In_743);
nor U743 (N_743,In_469,In_243);
nor U744 (N_744,In_1058,In_682);
or U745 (N_745,In_1420,In_2270);
nand U746 (N_746,In_2374,In_769);
xor U747 (N_747,In_1909,In_1742);
and U748 (N_748,In_1873,In_1406);
nand U749 (N_749,In_1737,In_1060);
nand U750 (N_750,In_1382,In_1632);
nor U751 (N_751,In_568,In_685);
nor U752 (N_752,In_2300,In_23);
xor U753 (N_753,In_1122,In_895);
nand U754 (N_754,In_1016,In_278);
nand U755 (N_755,In_1513,In_1055);
nor U756 (N_756,In_2392,In_1881);
nor U757 (N_757,In_861,In_734);
nand U758 (N_758,In_841,In_580);
and U759 (N_759,In_636,In_2400);
nand U760 (N_760,In_228,In_1374);
xnor U761 (N_761,In_1849,In_205);
xnor U762 (N_762,In_783,In_548);
and U763 (N_763,In_2033,In_1803);
and U764 (N_764,In_2490,In_227);
nor U765 (N_765,In_697,In_1754);
nor U766 (N_766,In_1263,In_2014);
or U767 (N_767,In_726,In_1221);
or U768 (N_768,In_2411,In_2205);
or U769 (N_769,In_1192,In_1092);
or U770 (N_770,In_348,In_655);
or U771 (N_771,In_451,In_131);
and U772 (N_772,In_1195,In_607);
nand U773 (N_773,In_725,In_461);
xnor U774 (N_774,In_499,In_1785);
or U775 (N_775,In_2081,In_30);
or U776 (N_776,In_1096,In_1165);
and U777 (N_777,In_1364,In_360);
nor U778 (N_778,In_997,In_2068);
and U779 (N_779,In_2346,In_1576);
nor U780 (N_780,In_1257,In_2377);
nand U781 (N_781,In_1988,In_1264);
or U782 (N_782,In_1265,In_2256);
nor U783 (N_783,In_966,In_1086);
nand U784 (N_784,In_1022,In_1501);
or U785 (N_785,In_645,In_574);
or U786 (N_786,In_1365,In_1056);
or U787 (N_787,In_2159,In_1774);
nor U788 (N_788,In_77,In_2160);
xor U789 (N_789,In_2006,In_609);
nor U790 (N_790,In_1038,In_42);
nand U791 (N_791,In_2381,In_249);
nand U792 (N_792,In_223,In_1472);
xnor U793 (N_793,In_1213,In_1642);
and U794 (N_794,In_855,In_1680);
xnor U795 (N_795,In_2389,In_2348);
xnor U796 (N_796,In_2369,In_1587);
nor U797 (N_797,In_2378,In_1202);
nand U798 (N_798,In_78,In_323);
or U799 (N_799,In_358,In_1146);
or U800 (N_800,In_2124,In_1329);
or U801 (N_801,In_1687,In_2401);
and U802 (N_802,In_2176,In_2062);
or U803 (N_803,In_1161,In_1941);
nand U804 (N_804,In_1439,In_161);
nor U805 (N_805,In_907,In_1495);
nand U806 (N_806,In_1689,In_1312);
and U807 (N_807,In_553,In_2187);
xnor U808 (N_808,In_1845,In_298);
nor U809 (N_809,In_1064,In_1606);
or U810 (N_810,In_2048,In_222);
nor U811 (N_811,In_1676,In_1730);
nand U812 (N_812,In_833,In_1480);
and U813 (N_813,In_1703,In_2101);
or U814 (N_814,In_286,In_1572);
nand U815 (N_815,In_1604,In_859);
or U816 (N_816,In_1003,In_2443);
nor U817 (N_817,In_967,In_971);
nor U818 (N_818,In_1786,In_457);
or U819 (N_819,In_2429,In_1781);
and U820 (N_820,In_1176,In_1497);
or U821 (N_821,In_1268,In_944);
nand U822 (N_822,In_1991,In_2299);
nor U823 (N_823,In_272,In_482);
or U824 (N_824,In_22,In_1074);
or U825 (N_825,In_1367,In_1542);
nand U826 (N_826,In_125,In_2200);
or U827 (N_827,In_1205,In_2456);
nand U828 (N_828,In_2220,In_910);
nand U829 (N_829,In_1277,In_2482);
and U830 (N_830,In_1019,In_722);
nor U831 (N_831,In_987,In_983);
or U832 (N_832,In_2440,In_1297);
nand U833 (N_833,In_1638,In_1111);
nor U834 (N_834,In_1034,In_1524);
nor U835 (N_835,In_1755,In_1568);
nand U836 (N_836,In_25,In_2496);
and U837 (N_837,In_1711,In_437);
or U838 (N_838,In_533,In_2419);
or U839 (N_839,In_1404,In_956);
or U840 (N_840,In_1249,In_1401);
nand U841 (N_841,In_1899,In_1442);
and U842 (N_842,In_1318,In_2480);
or U843 (N_843,In_1619,In_2171);
or U844 (N_844,In_423,In_180);
or U845 (N_845,In_1410,In_2317);
or U846 (N_846,In_1095,In_1138);
nand U847 (N_847,In_61,In_1591);
nor U848 (N_848,In_1090,In_1712);
nand U849 (N_849,In_212,In_1366);
nand U850 (N_850,In_508,In_1509);
or U851 (N_851,In_292,In_1848);
and U852 (N_852,In_1449,In_41);
nor U853 (N_853,In_1718,In_1915);
or U854 (N_854,In_1460,In_551);
and U855 (N_855,In_1600,In_1375);
nor U856 (N_856,In_920,In_511);
xor U857 (N_857,In_402,In_2055);
and U858 (N_858,In_75,In_1583);
xor U859 (N_859,In_89,In_1162);
nor U860 (N_860,In_1702,In_2208);
and U861 (N_861,In_1001,In_150);
nand U862 (N_862,In_320,In_1465);
nand U863 (N_863,In_394,In_1417);
or U864 (N_864,In_2343,In_940);
or U865 (N_865,In_530,In_624);
or U866 (N_866,In_253,In_294);
nand U867 (N_867,In_1008,In_1156);
xnor U868 (N_868,In_1305,In_217);
and U869 (N_869,In_1445,In_1750);
nor U870 (N_870,In_1218,In_1040);
nor U871 (N_871,In_1898,In_1998);
and U872 (N_872,In_515,In_709);
nand U873 (N_873,In_74,In_1467);
nand U874 (N_874,In_284,In_509);
nand U875 (N_875,In_361,In_1976);
or U876 (N_876,In_1456,In_18);
and U877 (N_877,In_1207,In_880);
xor U878 (N_878,In_1939,In_886);
or U879 (N_879,In_902,In_1585);
or U880 (N_880,In_31,In_2178);
nand U881 (N_881,In_1272,In_571);
nand U882 (N_882,In_244,In_339);
nand U883 (N_883,In_865,In_1946);
and U884 (N_884,In_720,In_660);
or U885 (N_885,In_1142,In_1654);
xor U886 (N_886,In_246,In_208);
or U887 (N_887,In_1659,In_1223);
nor U888 (N_888,In_633,In_1893);
and U889 (N_889,In_1648,In_1503);
and U890 (N_890,In_1462,In_1577);
nor U891 (N_891,In_2127,In_581);
or U892 (N_892,In_225,In_531);
nand U893 (N_893,In_867,In_1936);
nand U894 (N_894,In_601,In_625);
nand U895 (N_895,In_1057,In_856);
nor U896 (N_896,In_802,In_1061);
or U897 (N_897,In_1186,In_2104);
or U898 (N_898,In_1942,In_2082);
nor U899 (N_899,In_641,In_2390);
or U900 (N_900,In_693,In_1170);
nand U901 (N_901,In_367,In_425);
nand U902 (N_902,In_996,In_1217);
nor U903 (N_903,In_1979,In_1054);
nand U904 (N_904,In_2010,In_2358);
nand U905 (N_905,In_2437,In_1520);
nand U906 (N_906,In_187,In_2238);
nor U907 (N_907,In_371,In_606);
nand U908 (N_908,In_2274,In_2375);
nand U909 (N_909,In_914,In_2148);
or U910 (N_910,In_691,In_2185);
and U911 (N_911,In_2023,In_1252);
and U912 (N_912,In_2261,In_2096);
or U913 (N_913,In_2015,In_778);
xnor U914 (N_914,In_2355,In_1422);
or U915 (N_915,In_122,In_1725);
nor U916 (N_916,In_2280,In_702);
nand U917 (N_917,In_1532,In_2296);
and U918 (N_918,In_2410,In_893);
or U919 (N_919,In_1199,In_1380);
nor U920 (N_920,In_2431,In_594);
nor U921 (N_921,In_1453,In_338);
or U922 (N_922,In_1562,In_1955);
or U923 (N_923,In_1004,In_897);
xnor U924 (N_924,In_558,In_446);
or U925 (N_925,In_666,In_514);
or U926 (N_926,In_365,In_2108);
or U927 (N_927,In_2330,In_1751);
nand U928 (N_928,In_492,In_2350);
or U929 (N_929,In_1699,In_1993);
or U930 (N_930,In_1735,In_2064);
or U931 (N_931,In_55,In_373);
nand U932 (N_932,In_800,In_19);
and U933 (N_933,In_2211,In_1906);
and U934 (N_934,In_1592,In_2038);
or U935 (N_935,In_1053,In_309);
and U936 (N_936,In_1228,In_1869);
or U937 (N_937,In_1357,In_1574);
nor U938 (N_938,In_1796,In_622);
and U939 (N_939,In_981,In_713);
xnor U940 (N_940,In_759,In_923);
and U941 (N_941,In_681,In_667);
xnor U942 (N_942,In_1469,In_916);
nor U943 (N_943,In_2283,In_1351);
nor U944 (N_944,In_1100,In_2151);
and U945 (N_945,In_295,In_642);
and U946 (N_946,In_418,In_1570);
and U947 (N_947,In_64,In_1478);
and U948 (N_948,In_2371,In_343);
nand U949 (N_949,In_652,In_0);
or U950 (N_950,In_2084,In_2011);
nand U951 (N_951,In_1027,In_1185);
nand U952 (N_952,In_2354,In_1324);
or U953 (N_953,In_860,In_346);
nor U954 (N_954,In_1960,In_756);
and U955 (N_955,In_1874,In_1738);
nor U956 (N_956,In_1419,In_255);
nand U957 (N_957,In_1325,In_1116);
and U958 (N_958,In_331,In_2089);
and U959 (N_959,In_1222,In_1540);
nor U960 (N_960,In_745,In_184);
or U961 (N_961,In_1072,In_414);
and U962 (N_962,In_2314,In_735);
nor U963 (N_963,In_177,In_1700);
and U964 (N_964,In_2034,In_1259);
nor U965 (N_965,In_1782,In_1651);
and U966 (N_966,In_2134,In_700);
and U967 (N_967,In_2007,In_1812);
xnor U968 (N_968,In_135,In_39);
nand U969 (N_969,In_974,In_1601);
nand U970 (N_970,In_1085,In_1504);
nand U971 (N_971,In_1628,In_2029);
nor U972 (N_972,In_563,In_450);
xor U973 (N_973,In_1558,In_1120);
or U974 (N_974,In_547,In_2356);
nand U975 (N_975,In_1232,In_1455);
and U976 (N_976,In_2468,In_1922);
nor U977 (N_977,In_587,In_2492);
and U978 (N_978,In_1024,In_985);
nor U979 (N_979,In_281,In_2250);
nor U980 (N_980,In_2195,In_337);
nor U981 (N_981,In_1470,In_1296);
or U982 (N_982,In_825,In_1776);
or U983 (N_983,In_2417,In_832);
nor U984 (N_984,In_1208,In_1430);
nand U985 (N_985,In_37,In_2161);
nand U986 (N_986,In_1627,In_640);
and U987 (N_987,In_678,In_2019);
nor U988 (N_988,In_2469,In_2499);
or U989 (N_989,In_112,In_2473);
or U990 (N_990,In_465,In_728);
nor U991 (N_991,In_2368,In_1970);
nor U992 (N_992,In_994,In_1625);
nand U993 (N_993,In_1386,In_1108);
nand U994 (N_994,In_1306,In_764);
or U995 (N_995,In_2004,In_1586);
and U996 (N_996,In_335,In_1928);
and U997 (N_997,In_1514,In_214);
or U998 (N_998,In_2266,In_545);
nand U999 (N_999,In_2196,In_2028);
and U1000 (N_1000,In_823,In_2018);
nand U1001 (N_1001,In_2103,In_2146);
and U1002 (N_1002,In_318,In_2017);
and U1003 (N_1003,In_1791,In_928);
nand U1004 (N_1004,In_1168,In_1026);
xor U1005 (N_1005,In_555,In_877);
nand U1006 (N_1006,In_2049,In_2357);
and U1007 (N_1007,In_521,In_2426);
and U1008 (N_1008,In_1762,In_1377);
nand U1009 (N_1009,In_1062,In_2054);
nand U1010 (N_1010,In_1715,In_1402);
nand U1011 (N_1011,In_1806,In_1582);
and U1012 (N_1012,In_672,In_154);
nor U1013 (N_1013,In_199,In_1554);
nand U1014 (N_1014,In_1046,In_2471);
and U1015 (N_1015,In_1820,In_1461);
nor U1016 (N_1016,In_2170,In_103);
nor U1017 (N_1017,In_1270,In_2046);
nand U1018 (N_1018,In_1523,In_2311);
and U1019 (N_1019,In_516,In_506);
nand U1020 (N_1020,In_362,In_1081);
or U1021 (N_1021,In_556,In_238);
or U1022 (N_1022,In_1891,In_2177);
or U1023 (N_1023,In_1865,In_873);
nand U1024 (N_1024,In_729,In_911);
nand U1025 (N_1025,In_943,In_1637);
nor U1026 (N_1026,In_21,In_1747);
or U1027 (N_1027,In_1973,In_1262);
or U1028 (N_1028,In_2416,In_204);
nand U1029 (N_1029,In_1854,In_785);
or U1030 (N_1030,In_889,In_483);
or U1031 (N_1031,In_1706,In_1407);
xnor U1032 (N_1032,In_715,In_1233);
or U1033 (N_1033,In_1644,In_1728);
nand U1034 (N_1034,In_2168,In_203);
and U1035 (N_1035,In_1440,In_1771);
nor U1036 (N_1036,In_497,In_991);
or U1037 (N_1037,In_2109,In_801);
and U1038 (N_1038,In_1354,In_564);
or U1039 (N_1039,In_2066,In_1734);
and U1040 (N_1040,In_2383,In_1010);
nor U1041 (N_1041,In_592,In_2321);
or U1042 (N_1042,In_454,In_2123);
nand U1043 (N_1043,In_1975,In_1412);
nand U1044 (N_1044,In_478,In_1534);
and U1045 (N_1045,In_1425,In_2030);
nand U1046 (N_1046,In_456,In_1673);
nor U1047 (N_1047,In_630,In_282);
nand U1048 (N_1048,In_876,In_2403);
nor U1049 (N_1049,In_3,In_168);
nand U1050 (N_1050,In_471,In_463);
or U1051 (N_1051,In_1489,In_148);
or U1052 (N_1052,In_1897,In_1963);
nor U1053 (N_1053,In_1190,In_2137);
or U1054 (N_1054,In_699,In_13);
and U1055 (N_1055,In_752,In_1713);
and U1056 (N_1056,In_2035,In_1569);
or U1057 (N_1057,In_2246,In_354);
or U1058 (N_1058,In_2433,In_712);
or U1059 (N_1059,In_430,In_628);
xnor U1060 (N_1060,In_1433,In_1255);
nand U1061 (N_1061,In_236,In_814);
and U1062 (N_1062,In_344,In_2406);
nor U1063 (N_1063,In_1866,In_1537);
nor U1064 (N_1064,In_319,In_1327);
or U1065 (N_1065,In_863,In_1686);
and U1066 (N_1066,In_737,In_1481);
or U1067 (N_1067,In_289,In_1337);
and U1068 (N_1068,In_2209,In_1248);
nor U1069 (N_1069,In_1241,In_1179);
nor U1070 (N_1070,In_617,In_1835);
nand U1071 (N_1071,In_1051,In_816);
nand U1072 (N_1072,In_659,In_2404);
nor U1073 (N_1073,In_487,In_1589);
nor U1074 (N_1074,In_299,In_1240);
and U1075 (N_1075,In_341,In_1082);
and U1076 (N_1076,In_1618,In_1945);
or U1077 (N_1077,In_792,In_1818);
or U1078 (N_1078,In_2347,In_1544);
or U1079 (N_1079,In_958,In_650);
xnor U1080 (N_1080,In_1833,In_143);
nand U1081 (N_1081,In_1887,In_513);
nand U1082 (N_1082,In_2407,In_2043);
nand U1083 (N_1083,In_993,In_1931);
nand U1084 (N_1084,In_314,In_1173);
nand U1085 (N_1085,In_2477,In_1943);
nor U1086 (N_1086,In_2396,In_1609);
xor U1087 (N_1087,In_2128,In_48);
xor U1088 (N_1088,In_1230,In_1964);
nor U1089 (N_1089,In_2152,In_1563);
and U1090 (N_1090,In_629,In_1630);
and U1091 (N_1091,In_1089,In_1067);
xnor U1092 (N_1092,In_2329,In_121);
or U1093 (N_1093,In_20,In_2240);
xnor U1094 (N_1094,In_489,In_2412);
xnor U1095 (N_1095,In_676,In_258);
xnor U1096 (N_1096,In_1847,In_1672);
or U1097 (N_1097,In_277,In_1695);
and U1098 (N_1098,In_1110,In_2418);
and U1099 (N_1099,In_93,In_2475);
nor U1100 (N_1100,In_300,In_81);
nand U1101 (N_1101,In_427,In_2385);
and U1102 (N_1102,In_2156,In_1892);
nand U1103 (N_1103,In_1431,In_1392);
nand U1104 (N_1104,In_2247,In_781);
nor U1105 (N_1105,In_1925,In_1746);
nand U1106 (N_1106,In_1322,In_866);
and U1107 (N_1107,In_1787,In_1113);
xor U1108 (N_1108,In_2394,In_1827);
nand U1109 (N_1109,In_1934,In_1856);
nand U1110 (N_1110,In_1885,In_2324);
nor U1111 (N_1111,In_2058,In_1239);
nand U1112 (N_1112,In_589,In_382);
and U1113 (N_1113,In_930,In_1862);
nand U1114 (N_1114,In_237,In_1674);
nand U1115 (N_1115,In_757,In_1617);
nor U1116 (N_1116,In_1736,In_1446);
and U1117 (N_1117,In_1238,In_1032);
nor U1118 (N_1118,In_357,In_126);
nor U1119 (N_1119,In_392,In_1400);
nand U1120 (N_1120,In_1875,In_1962);
or U1121 (N_1121,In_505,In_132);
nand U1122 (N_1122,In_2093,In_1904);
nor U1123 (N_1123,In_333,In_1294);
nand U1124 (N_1124,In_2204,In_43);
and U1125 (N_1125,In_646,In_2172);
or U1126 (N_1126,In_142,In_182);
xor U1127 (N_1127,In_2395,In_262);
nand U1128 (N_1128,In_256,In_2083);
nor U1129 (N_1129,In_1669,In_811);
and U1130 (N_1130,In_952,In_2264);
and U1131 (N_1131,In_1098,In_688);
xnor U1132 (N_1132,In_1350,In_416);
nand U1133 (N_1133,In_1610,In_1724);
nand U1134 (N_1134,In_98,In_502);
nand U1135 (N_1135,In_1049,In_2140);
nand U1136 (N_1136,In_1971,In_1063);
nand U1137 (N_1137,In_1131,In_1631);
or U1138 (N_1138,In_174,In_1454);
and U1139 (N_1139,In_585,In_1283);
and U1140 (N_1140,In_1253,In_608);
and U1141 (N_1141,In_422,In_405);
nor U1142 (N_1142,In_872,In_501);
or U1143 (N_1143,In_724,In_2147);
and U1144 (N_1144,In_226,In_2013);
and U1145 (N_1145,In_1413,In_2341);
nor U1146 (N_1146,In_16,In_2221);
nor U1147 (N_1147,In_2257,In_842);
nand U1148 (N_1148,In_937,In_59);
and U1149 (N_1149,In_1535,In_765);
nor U1150 (N_1150,In_718,In_1474);
or U1151 (N_1151,In_1530,In_2457);
nand U1152 (N_1152,In_85,In_1429);
and U1153 (N_1153,In_1743,In_2448);
nand U1154 (N_1154,In_1984,In_2157);
nor U1155 (N_1155,In_71,In_1959);
nor U1156 (N_1156,In_918,In_2130);
or U1157 (N_1157,In_17,In_537);
and U1158 (N_1158,In_586,In_763);
or U1159 (N_1159,In_2025,In_192);
or U1160 (N_1160,In_2408,In_2465);
and U1161 (N_1161,In_1242,In_2189);
nor U1162 (N_1162,In_1635,In_194);
nand U1163 (N_1163,In_1308,In_1766);
or U1164 (N_1164,In_356,In_2016);
and U1165 (N_1165,In_308,In_488);
and U1166 (N_1166,In_145,In_1800);
or U1167 (N_1167,In_957,In_2472);
or U1168 (N_1168,In_146,In_275);
nand U1169 (N_1169,In_1788,In_898);
and U1170 (N_1170,In_661,In_1196);
and U1171 (N_1171,In_909,In_1415);
or U1172 (N_1172,In_1342,In_1289);
nand U1173 (N_1173,In_216,In_1136);
and U1174 (N_1174,In_1434,In_252);
or U1175 (N_1175,In_2162,In_2044);
or U1176 (N_1176,In_53,In_1831);
and U1177 (N_1177,In_1679,In_990);
nand U1178 (N_1178,In_1879,In_1525);
nor U1179 (N_1179,In_2098,In_961);
or U1180 (N_1180,In_2094,In_714);
nor U1181 (N_1181,In_1515,In_247);
and U1182 (N_1182,In_794,In_805);
nor U1183 (N_1183,In_306,In_1391);
and U1184 (N_1184,In_760,In_1890);
nand U1185 (N_1185,In_1996,In_2333);
xnor U1186 (N_1186,In_1304,In_1767);
or U1187 (N_1187,In_1409,In_195);
and U1188 (N_1188,In_2194,In_1597);
nor U1189 (N_1189,In_1668,In_1463);
and U1190 (N_1190,In_2327,In_2255);
nor U1191 (N_1191,In_2243,In_1902);
and U1192 (N_1192,In_1368,In_1982);
nand U1193 (N_1193,In_2464,In_552);
or U1194 (N_1194,In_1761,In_313);
nor U1195 (N_1195,In_2339,In_1760);
nor U1196 (N_1196,In_467,In_2405);
or U1197 (N_1197,In_2293,In_838);
and U1198 (N_1198,In_946,In_2227);
and U1199 (N_1199,In_116,In_1126);
nand U1200 (N_1200,In_1229,In_2491);
nand U1201 (N_1201,In_793,In_602);
nor U1202 (N_1202,In_1759,In_1553);
or U1203 (N_1203,In_1184,In_26);
or U1204 (N_1204,In_1958,In_542);
nand U1205 (N_1205,In_1896,In_2316);
and U1206 (N_1206,In_2249,In_464);
or U1207 (N_1207,In_1212,In_1029);
and U1208 (N_1208,In_570,In_1083);
nand U1209 (N_1209,In_1394,In_2322);
nand U1210 (N_1210,In_1033,In_1967);
and U1211 (N_1211,In_980,In_913);
or U1212 (N_1212,In_2075,In_2312);
nand U1213 (N_1213,In_1210,In_968);
nor U1214 (N_1214,In_1494,In_1174);
nor U1215 (N_1215,In_491,In_1726);
nand U1216 (N_1216,In_2174,In_1789);
nor U1217 (N_1217,In_459,In_1370);
or U1218 (N_1218,In_741,In_739);
nor U1219 (N_1219,In_413,In_2252);
nor U1220 (N_1220,In_905,In_1911);
xor U1221 (N_1221,In_1705,In_746);
nand U1222 (N_1222,In_2191,In_1511);
or U1223 (N_1223,In_1340,In_152);
nor U1224 (N_1224,In_2022,In_598);
nand U1225 (N_1225,In_1275,In_1139);
nand U1226 (N_1226,In_1302,In_1593);
nor U1227 (N_1227,In_2453,In_1490);
or U1228 (N_1228,In_2077,In_2304);
xnor U1229 (N_1229,In_1797,In_409);
and U1230 (N_1230,In_1291,In_1633);
or U1231 (N_1231,In_2045,In_1452);
or U1232 (N_1232,In_167,In_799);
nor U1233 (N_1233,In_117,In_1837);
xnor U1234 (N_1234,In_270,In_1678);
nand U1235 (N_1235,In_596,In_1426);
or U1236 (N_1236,In_330,In_2291);
xnor U1237 (N_1237,In_1428,In_368);
xnor U1238 (N_1238,In_717,In_2114);
nor U1239 (N_1239,In_2360,In_2154);
xnor U1240 (N_1240,In_213,In_950);
or U1241 (N_1241,In_2413,In_1935);
or U1242 (N_1242,In_1799,In_163);
and U1243 (N_1243,In_1140,In_251);
nand U1244 (N_1244,In_2144,In_2244);
xor U1245 (N_1245,In_115,In_1826);
and U1246 (N_1246,In_315,In_1795);
or U1247 (N_1247,In_440,In_155);
or U1248 (N_1248,In_2021,In_106);
xnor U1249 (N_1249,In_2365,In_2253);
and U1250 (N_1250,In_1071,In_2202);
and U1251 (N_1251,In_1984,In_1228);
or U1252 (N_1252,In_1100,In_22);
and U1253 (N_1253,In_2451,In_2171);
nand U1254 (N_1254,In_2263,In_1613);
nor U1255 (N_1255,In_1455,In_127);
and U1256 (N_1256,In_304,In_1079);
and U1257 (N_1257,In_43,In_322);
nand U1258 (N_1258,In_1526,In_164);
and U1259 (N_1259,In_878,In_1107);
and U1260 (N_1260,In_1642,In_2281);
nor U1261 (N_1261,In_1632,In_1840);
nand U1262 (N_1262,In_777,In_1793);
and U1263 (N_1263,In_1131,In_1199);
or U1264 (N_1264,In_2369,In_2499);
and U1265 (N_1265,In_1720,In_1330);
nor U1266 (N_1266,In_1850,In_213);
nor U1267 (N_1267,In_1963,In_1294);
nor U1268 (N_1268,In_426,In_2);
nand U1269 (N_1269,In_1994,In_2011);
nand U1270 (N_1270,In_146,In_1684);
and U1271 (N_1271,In_390,In_2370);
xnor U1272 (N_1272,In_1307,In_2185);
xor U1273 (N_1273,In_1062,In_880);
or U1274 (N_1274,In_2200,In_1499);
nor U1275 (N_1275,In_1464,In_2427);
nor U1276 (N_1276,In_564,In_533);
or U1277 (N_1277,In_1629,In_1798);
nand U1278 (N_1278,In_2122,In_768);
nor U1279 (N_1279,In_1567,In_714);
nor U1280 (N_1280,In_1028,In_1294);
nor U1281 (N_1281,In_563,In_954);
nor U1282 (N_1282,In_153,In_1311);
and U1283 (N_1283,In_158,In_1340);
or U1284 (N_1284,In_1322,In_1856);
nor U1285 (N_1285,In_2096,In_1475);
nand U1286 (N_1286,In_2344,In_128);
or U1287 (N_1287,In_1253,In_242);
nor U1288 (N_1288,In_2478,In_2255);
nand U1289 (N_1289,In_2131,In_376);
or U1290 (N_1290,In_589,In_669);
and U1291 (N_1291,In_2331,In_1520);
nand U1292 (N_1292,In_1403,In_946);
xnor U1293 (N_1293,In_1805,In_1517);
or U1294 (N_1294,In_607,In_847);
or U1295 (N_1295,In_2092,In_2096);
nor U1296 (N_1296,In_537,In_1235);
xnor U1297 (N_1297,In_2235,In_134);
and U1298 (N_1298,In_2381,In_2365);
and U1299 (N_1299,In_2247,In_2245);
and U1300 (N_1300,In_1912,In_2425);
or U1301 (N_1301,In_491,In_1937);
nand U1302 (N_1302,In_2221,In_1699);
and U1303 (N_1303,In_534,In_1483);
or U1304 (N_1304,In_1971,In_2337);
nor U1305 (N_1305,In_2256,In_517);
nand U1306 (N_1306,In_2209,In_2270);
and U1307 (N_1307,In_2072,In_522);
nor U1308 (N_1308,In_60,In_827);
nand U1309 (N_1309,In_966,In_724);
nor U1310 (N_1310,In_1186,In_1085);
nand U1311 (N_1311,In_91,In_2003);
nand U1312 (N_1312,In_417,In_403);
and U1313 (N_1313,In_2469,In_1635);
xnor U1314 (N_1314,In_1362,In_66);
and U1315 (N_1315,In_1434,In_279);
xnor U1316 (N_1316,In_11,In_748);
or U1317 (N_1317,In_1560,In_1260);
xnor U1318 (N_1318,In_1259,In_1562);
and U1319 (N_1319,In_176,In_2181);
nor U1320 (N_1320,In_751,In_1435);
nand U1321 (N_1321,In_1750,In_145);
and U1322 (N_1322,In_2459,In_2111);
xor U1323 (N_1323,In_2139,In_2224);
nand U1324 (N_1324,In_1204,In_1028);
and U1325 (N_1325,In_824,In_766);
and U1326 (N_1326,In_251,In_1189);
or U1327 (N_1327,In_2236,In_1929);
nand U1328 (N_1328,In_1489,In_1945);
or U1329 (N_1329,In_455,In_1086);
and U1330 (N_1330,In_2272,In_1685);
or U1331 (N_1331,In_2225,In_287);
nor U1332 (N_1332,In_2009,In_1386);
or U1333 (N_1333,In_1446,In_566);
nand U1334 (N_1334,In_1893,In_874);
nand U1335 (N_1335,In_501,In_1541);
or U1336 (N_1336,In_958,In_1448);
nor U1337 (N_1337,In_700,In_1757);
xnor U1338 (N_1338,In_374,In_858);
nand U1339 (N_1339,In_365,In_958);
or U1340 (N_1340,In_2133,In_1498);
or U1341 (N_1341,In_418,In_782);
or U1342 (N_1342,In_259,In_2214);
nand U1343 (N_1343,In_1857,In_1553);
or U1344 (N_1344,In_1663,In_1495);
or U1345 (N_1345,In_2139,In_153);
and U1346 (N_1346,In_884,In_1806);
and U1347 (N_1347,In_1720,In_1883);
nor U1348 (N_1348,In_1726,In_1842);
and U1349 (N_1349,In_2426,In_1159);
xor U1350 (N_1350,In_848,In_67);
nor U1351 (N_1351,In_424,In_1105);
nor U1352 (N_1352,In_1028,In_1447);
or U1353 (N_1353,In_2448,In_209);
nor U1354 (N_1354,In_84,In_2384);
and U1355 (N_1355,In_976,In_1325);
nand U1356 (N_1356,In_1242,In_98);
and U1357 (N_1357,In_2167,In_2060);
nor U1358 (N_1358,In_1054,In_342);
nor U1359 (N_1359,In_430,In_2200);
and U1360 (N_1360,In_2436,In_1942);
nand U1361 (N_1361,In_1948,In_1952);
nor U1362 (N_1362,In_1594,In_1608);
and U1363 (N_1363,In_2147,In_92);
nand U1364 (N_1364,In_1085,In_979);
and U1365 (N_1365,In_558,In_443);
xor U1366 (N_1366,In_862,In_2260);
or U1367 (N_1367,In_101,In_1494);
or U1368 (N_1368,In_1256,In_2277);
nand U1369 (N_1369,In_2268,In_2214);
nand U1370 (N_1370,In_906,In_2496);
and U1371 (N_1371,In_198,In_901);
or U1372 (N_1372,In_2049,In_519);
and U1373 (N_1373,In_2136,In_608);
nand U1374 (N_1374,In_1695,In_1462);
and U1375 (N_1375,In_1664,In_507);
nor U1376 (N_1376,In_2343,In_2297);
nor U1377 (N_1377,In_2140,In_579);
and U1378 (N_1378,In_1171,In_587);
and U1379 (N_1379,In_764,In_714);
xor U1380 (N_1380,In_921,In_56);
or U1381 (N_1381,In_1193,In_325);
or U1382 (N_1382,In_10,In_1715);
nand U1383 (N_1383,In_1594,In_740);
or U1384 (N_1384,In_1847,In_1917);
xnor U1385 (N_1385,In_1554,In_131);
nand U1386 (N_1386,In_1735,In_608);
nand U1387 (N_1387,In_2209,In_1387);
nand U1388 (N_1388,In_908,In_1980);
nor U1389 (N_1389,In_2465,In_950);
or U1390 (N_1390,In_2131,In_132);
or U1391 (N_1391,In_1123,In_1440);
and U1392 (N_1392,In_342,In_1555);
nor U1393 (N_1393,In_1046,In_1429);
and U1394 (N_1394,In_2196,In_1248);
and U1395 (N_1395,In_1833,In_483);
nor U1396 (N_1396,In_1619,In_2248);
and U1397 (N_1397,In_1804,In_1552);
and U1398 (N_1398,In_507,In_1589);
nor U1399 (N_1399,In_1813,In_575);
or U1400 (N_1400,In_2143,In_97);
and U1401 (N_1401,In_2322,In_2132);
nand U1402 (N_1402,In_489,In_1586);
xnor U1403 (N_1403,In_339,In_873);
xnor U1404 (N_1404,In_1885,In_786);
nand U1405 (N_1405,In_1518,In_76);
and U1406 (N_1406,In_1389,In_54);
nand U1407 (N_1407,In_2320,In_1998);
or U1408 (N_1408,In_496,In_2462);
nand U1409 (N_1409,In_47,In_1449);
or U1410 (N_1410,In_327,In_972);
nor U1411 (N_1411,In_260,In_1375);
nand U1412 (N_1412,In_2487,In_726);
nor U1413 (N_1413,In_841,In_340);
or U1414 (N_1414,In_455,In_2148);
or U1415 (N_1415,In_2144,In_299);
or U1416 (N_1416,In_2424,In_858);
nor U1417 (N_1417,In_812,In_1355);
or U1418 (N_1418,In_50,In_370);
or U1419 (N_1419,In_2,In_1729);
xor U1420 (N_1420,In_330,In_378);
and U1421 (N_1421,In_1051,In_311);
and U1422 (N_1422,In_1120,In_1891);
and U1423 (N_1423,In_2205,In_1870);
nand U1424 (N_1424,In_927,In_2245);
or U1425 (N_1425,In_1666,In_444);
nor U1426 (N_1426,In_1357,In_2070);
nor U1427 (N_1427,In_1093,In_1095);
xor U1428 (N_1428,In_702,In_206);
nand U1429 (N_1429,In_1986,In_836);
nor U1430 (N_1430,In_1935,In_614);
nand U1431 (N_1431,In_397,In_1257);
and U1432 (N_1432,In_541,In_1431);
nor U1433 (N_1433,In_1744,In_1815);
nand U1434 (N_1434,In_599,In_342);
or U1435 (N_1435,In_12,In_1135);
and U1436 (N_1436,In_1565,In_72);
nor U1437 (N_1437,In_268,In_1600);
nand U1438 (N_1438,In_1201,In_2399);
or U1439 (N_1439,In_2046,In_459);
and U1440 (N_1440,In_2286,In_2418);
nor U1441 (N_1441,In_328,In_1899);
and U1442 (N_1442,In_1692,In_2304);
and U1443 (N_1443,In_2118,In_2414);
nand U1444 (N_1444,In_1347,In_811);
and U1445 (N_1445,In_964,In_798);
xor U1446 (N_1446,In_2424,In_335);
and U1447 (N_1447,In_1066,In_151);
nor U1448 (N_1448,In_69,In_1518);
and U1449 (N_1449,In_152,In_2473);
nor U1450 (N_1450,In_1292,In_666);
or U1451 (N_1451,In_2156,In_2388);
nand U1452 (N_1452,In_888,In_697);
nor U1453 (N_1453,In_1609,In_682);
or U1454 (N_1454,In_229,In_1382);
or U1455 (N_1455,In_59,In_1960);
xor U1456 (N_1456,In_54,In_1676);
or U1457 (N_1457,In_1165,In_1701);
nor U1458 (N_1458,In_1447,In_1938);
and U1459 (N_1459,In_2394,In_1188);
or U1460 (N_1460,In_2060,In_1083);
nor U1461 (N_1461,In_7,In_1125);
xnor U1462 (N_1462,In_569,In_986);
nor U1463 (N_1463,In_1846,In_2451);
nand U1464 (N_1464,In_1534,In_1491);
and U1465 (N_1465,In_997,In_693);
and U1466 (N_1466,In_653,In_775);
xor U1467 (N_1467,In_1304,In_2101);
nand U1468 (N_1468,In_2092,In_132);
and U1469 (N_1469,In_2438,In_1710);
nand U1470 (N_1470,In_59,In_742);
xor U1471 (N_1471,In_1143,In_266);
or U1472 (N_1472,In_686,In_2437);
nand U1473 (N_1473,In_90,In_2233);
xor U1474 (N_1474,In_285,In_1076);
nand U1475 (N_1475,In_1215,In_1467);
nor U1476 (N_1476,In_352,In_1420);
and U1477 (N_1477,In_548,In_2413);
or U1478 (N_1478,In_146,In_1925);
or U1479 (N_1479,In_1449,In_2222);
nor U1480 (N_1480,In_486,In_155);
nand U1481 (N_1481,In_358,In_1428);
or U1482 (N_1482,In_133,In_1552);
xor U1483 (N_1483,In_362,In_100);
and U1484 (N_1484,In_942,In_710);
nor U1485 (N_1485,In_382,In_1680);
or U1486 (N_1486,In_744,In_2013);
xor U1487 (N_1487,In_404,In_384);
nor U1488 (N_1488,In_589,In_1953);
nor U1489 (N_1489,In_242,In_256);
and U1490 (N_1490,In_1791,In_2238);
or U1491 (N_1491,In_1892,In_104);
or U1492 (N_1492,In_1616,In_140);
and U1493 (N_1493,In_19,In_1343);
or U1494 (N_1494,In_1005,In_563);
nor U1495 (N_1495,In_1929,In_140);
nand U1496 (N_1496,In_2089,In_81);
nor U1497 (N_1497,In_932,In_1098);
and U1498 (N_1498,In_540,In_630);
and U1499 (N_1499,In_2037,In_1962);
and U1500 (N_1500,In_226,In_2353);
nor U1501 (N_1501,In_825,In_946);
and U1502 (N_1502,In_2013,In_1556);
nand U1503 (N_1503,In_1753,In_2343);
xnor U1504 (N_1504,In_2027,In_2498);
or U1505 (N_1505,In_1748,In_1808);
nor U1506 (N_1506,In_1941,In_95);
nand U1507 (N_1507,In_1631,In_1946);
and U1508 (N_1508,In_868,In_2360);
nor U1509 (N_1509,In_1015,In_1309);
nand U1510 (N_1510,In_1551,In_1968);
or U1511 (N_1511,In_88,In_367);
and U1512 (N_1512,In_1706,In_1380);
or U1513 (N_1513,In_2352,In_1930);
or U1514 (N_1514,In_2017,In_1550);
nor U1515 (N_1515,In_2051,In_196);
nand U1516 (N_1516,In_2002,In_1015);
nor U1517 (N_1517,In_1068,In_683);
or U1518 (N_1518,In_2029,In_293);
or U1519 (N_1519,In_2357,In_685);
and U1520 (N_1520,In_636,In_702);
and U1521 (N_1521,In_1086,In_633);
nand U1522 (N_1522,In_38,In_2337);
nand U1523 (N_1523,In_101,In_2312);
and U1524 (N_1524,In_288,In_1255);
xor U1525 (N_1525,In_664,In_1422);
or U1526 (N_1526,In_1290,In_1187);
nand U1527 (N_1527,In_515,In_1191);
nor U1528 (N_1528,In_2076,In_2360);
and U1529 (N_1529,In_793,In_1829);
and U1530 (N_1530,In_333,In_1238);
nand U1531 (N_1531,In_1146,In_1413);
nand U1532 (N_1532,In_1527,In_1949);
xnor U1533 (N_1533,In_949,In_221);
and U1534 (N_1534,In_2444,In_896);
nor U1535 (N_1535,In_2039,In_594);
and U1536 (N_1536,In_1935,In_748);
nor U1537 (N_1537,In_2194,In_2223);
or U1538 (N_1538,In_1037,In_1961);
nor U1539 (N_1539,In_2076,In_2250);
nand U1540 (N_1540,In_1305,In_67);
xor U1541 (N_1541,In_514,In_2287);
and U1542 (N_1542,In_1032,In_2141);
or U1543 (N_1543,In_1350,In_470);
nor U1544 (N_1544,In_1757,In_1443);
or U1545 (N_1545,In_161,In_2224);
nand U1546 (N_1546,In_1747,In_628);
xnor U1547 (N_1547,In_2477,In_1035);
and U1548 (N_1548,In_2314,In_1374);
nor U1549 (N_1549,In_94,In_2117);
nor U1550 (N_1550,In_144,In_1249);
nand U1551 (N_1551,In_1252,In_1274);
nor U1552 (N_1552,In_772,In_462);
xor U1553 (N_1553,In_1701,In_1247);
and U1554 (N_1554,In_99,In_1910);
nand U1555 (N_1555,In_1166,In_2021);
and U1556 (N_1556,In_1181,In_885);
nor U1557 (N_1557,In_737,In_459);
nor U1558 (N_1558,In_1255,In_1968);
nor U1559 (N_1559,In_2379,In_1648);
and U1560 (N_1560,In_900,In_2442);
nand U1561 (N_1561,In_1928,In_1886);
and U1562 (N_1562,In_539,In_1414);
nor U1563 (N_1563,In_2126,In_1675);
nor U1564 (N_1564,In_2360,In_721);
nor U1565 (N_1565,In_1926,In_1628);
nand U1566 (N_1566,In_2441,In_1789);
and U1567 (N_1567,In_1480,In_226);
nor U1568 (N_1568,In_2220,In_28);
nand U1569 (N_1569,In_1212,In_1652);
and U1570 (N_1570,In_401,In_1570);
and U1571 (N_1571,In_1493,In_2196);
nor U1572 (N_1572,In_1620,In_1253);
nor U1573 (N_1573,In_660,In_581);
nand U1574 (N_1574,In_2309,In_1917);
or U1575 (N_1575,In_1708,In_1484);
nand U1576 (N_1576,In_1718,In_1607);
and U1577 (N_1577,In_1681,In_1044);
nor U1578 (N_1578,In_1325,In_1358);
and U1579 (N_1579,In_661,In_683);
and U1580 (N_1580,In_813,In_102);
nor U1581 (N_1581,In_1122,In_1603);
and U1582 (N_1582,In_1984,In_1581);
nand U1583 (N_1583,In_886,In_2284);
nand U1584 (N_1584,In_647,In_1440);
or U1585 (N_1585,In_1221,In_584);
or U1586 (N_1586,In_590,In_1590);
xnor U1587 (N_1587,In_1251,In_916);
nand U1588 (N_1588,In_2465,In_87);
nand U1589 (N_1589,In_536,In_69);
or U1590 (N_1590,In_2222,In_510);
nor U1591 (N_1591,In_2377,In_2192);
nand U1592 (N_1592,In_2173,In_64);
or U1593 (N_1593,In_1780,In_2238);
and U1594 (N_1594,In_787,In_2165);
and U1595 (N_1595,In_1273,In_737);
nor U1596 (N_1596,In_291,In_2316);
nor U1597 (N_1597,In_2014,In_1806);
and U1598 (N_1598,In_701,In_1538);
nand U1599 (N_1599,In_71,In_793);
nor U1600 (N_1600,In_1047,In_430);
or U1601 (N_1601,In_1350,In_84);
nor U1602 (N_1602,In_1335,In_364);
or U1603 (N_1603,In_1747,In_20);
nand U1604 (N_1604,In_2480,In_2476);
or U1605 (N_1605,In_1170,In_1394);
nand U1606 (N_1606,In_2489,In_881);
nor U1607 (N_1607,In_2182,In_213);
nor U1608 (N_1608,In_1434,In_941);
nand U1609 (N_1609,In_637,In_1298);
nand U1610 (N_1610,In_1346,In_282);
nor U1611 (N_1611,In_1200,In_1255);
xnor U1612 (N_1612,In_2100,In_899);
xor U1613 (N_1613,In_779,In_2290);
nor U1614 (N_1614,In_1667,In_1688);
and U1615 (N_1615,In_323,In_2021);
and U1616 (N_1616,In_2119,In_645);
nand U1617 (N_1617,In_860,In_2125);
nand U1618 (N_1618,In_1820,In_1778);
nand U1619 (N_1619,In_1329,In_1933);
or U1620 (N_1620,In_1002,In_1230);
nor U1621 (N_1621,In_2356,In_250);
nor U1622 (N_1622,In_627,In_2482);
or U1623 (N_1623,In_865,In_1952);
and U1624 (N_1624,In_53,In_1556);
or U1625 (N_1625,In_150,In_2181);
or U1626 (N_1626,In_1473,In_987);
nand U1627 (N_1627,In_640,In_198);
nand U1628 (N_1628,In_2235,In_1985);
nor U1629 (N_1629,In_1812,In_1533);
and U1630 (N_1630,In_1507,In_931);
and U1631 (N_1631,In_1884,In_1059);
nand U1632 (N_1632,In_2440,In_1703);
or U1633 (N_1633,In_2,In_88);
and U1634 (N_1634,In_2071,In_189);
nor U1635 (N_1635,In_829,In_247);
and U1636 (N_1636,In_1945,In_1214);
nor U1637 (N_1637,In_2106,In_330);
xnor U1638 (N_1638,In_1412,In_2060);
nand U1639 (N_1639,In_2136,In_885);
nand U1640 (N_1640,In_1751,In_670);
or U1641 (N_1641,In_849,In_1086);
or U1642 (N_1642,In_2272,In_571);
and U1643 (N_1643,In_2246,In_1594);
and U1644 (N_1644,In_1817,In_1461);
xor U1645 (N_1645,In_2277,In_891);
and U1646 (N_1646,In_1368,In_2000);
xor U1647 (N_1647,In_698,In_1359);
nor U1648 (N_1648,In_2406,In_2213);
and U1649 (N_1649,In_2406,In_1723);
and U1650 (N_1650,In_1279,In_2440);
nor U1651 (N_1651,In_2297,In_526);
nor U1652 (N_1652,In_68,In_565);
nand U1653 (N_1653,In_2178,In_2226);
nor U1654 (N_1654,In_302,In_2364);
or U1655 (N_1655,In_389,In_1976);
nand U1656 (N_1656,In_2376,In_1761);
and U1657 (N_1657,In_460,In_983);
nor U1658 (N_1658,In_1552,In_1982);
nand U1659 (N_1659,In_626,In_1568);
or U1660 (N_1660,In_851,In_1628);
nand U1661 (N_1661,In_2277,In_922);
nand U1662 (N_1662,In_440,In_1363);
or U1663 (N_1663,In_1867,In_1152);
nand U1664 (N_1664,In_1104,In_1936);
or U1665 (N_1665,In_1511,In_734);
nand U1666 (N_1666,In_1339,In_2076);
nor U1667 (N_1667,In_2320,In_658);
nor U1668 (N_1668,In_1644,In_2104);
and U1669 (N_1669,In_1018,In_1500);
and U1670 (N_1670,In_650,In_1362);
or U1671 (N_1671,In_1346,In_397);
nor U1672 (N_1672,In_1210,In_398);
nor U1673 (N_1673,In_1343,In_1926);
nor U1674 (N_1674,In_2040,In_1487);
nand U1675 (N_1675,In_2008,In_2146);
and U1676 (N_1676,In_414,In_2482);
or U1677 (N_1677,In_1972,In_800);
nor U1678 (N_1678,In_693,In_1189);
or U1679 (N_1679,In_1996,In_1090);
or U1680 (N_1680,In_1580,In_2101);
nand U1681 (N_1681,In_956,In_1907);
nor U1682 (N_1682,In_1100,In_1107);
nand U1683 (N_1683,In_398,In_708);
and U1684 (N_1684,In_2259,In_1009);
and U1685 (N_1685,In_1779,In_871);
xnor U1686 (N_1686,In_2210,In_1216);
nor U1687 (N_1687,In_1082,In_65);
and U1688 (N_1688,In_1653,In_470);
or U1689 (N_1689,In_1566,In_2215);
xnor U1690 (N_1690,In_648,In_350);
nor U1691 (N_1691,In_442,In_1524);
and U1692 (N_1692,In_2298,In_2204);
nand U1693 (N_1693,In_303,In_1930);
and U1694 (N_1694,In_2274,In_853);
or U1695 (N_1695,In_1263,In_2125);
or U1696 (N_1696,In_1573,In_716);
nand U1697 (N_1697,In_654,In_1133);
and U1698 (N_1698,In_133,In_698);
xnor U1699 (N_1699,In_814,In_1072);
or U1700 (N_1700,In_1003,In_678);
nor U1701 (N_1701,In_2336,In_607);
and U1702 (N_1702,In_1127,In_218);
nor U1703 (N_1703,In_1135,In_604);
nand U1704 (N_1704,In_1898,In_214);
nand U1705 (N_1705,In_1459,In_2087);
nor U1706 (N_1706,In_2058,In_906);
nor U1707 (N_1707,In_415,In_1715);
nor U1708 (N_1708,In_1716,In_810);
nor U1709 (N_1709,In_1718,In_607);
nor U1710 (N_1710,In_231,In_988);
or U1711 (N_1711,In_1023,In_445);
nor U1712 (N_1712,In_245,In_1455);
and U1713 (N_1713,In_1007,In_1038);
nand U1714 (N_1714,In_1714,In_1439);
nor U1715 (N_1715,In_1999,In_618);
nor U1716 (N_1716,In_388,In_1913);
and U1717 (N_1717,In_127,In_1640);
or U1718 (N_1718,In_2059,In_1567);
nor U1719 (N_1719,In_1790,In_431);
nand U1720 (N_1720,In_1272,In_593);
xor U1721 (N_1721,In_787,In_76);
nor U1722 (N_1722,In_1380,In_1999);
nand U1723 (N_1723,In_1624,In_1450);
and U1724 (N_1724,In_1671,In_2128);
or U1725 (N_1725,In_2085,In_2049);
and U1726 (N_1726,In_2493,In_829);
xnor U1727 (N_1727,In_915,In_2396);
xnor U1728 (N_1728,In_2082,In_1083);
and U1729 (N_1729,In_1084,In_1263);
nand U1730 (N_1730,In_7,In_478);
or U1731 (N_1731,In_1931,In_2065);
and U1732 (N_1732,In_73,In_1095);
nand U1733 (N_1733,In_440,In_2448);
nor U1734 (N_1734,In_2088,In_1142);
and U1735 (N_1735,In_2011,In_1684);
and U1736 (N_1736,In_1238,In_1693);
or U1737 (N_1737,In_968,In_805);
and U1738 (N_1738,In_616,In_1829);
nor U1739 (N_1739,In_1170,In_21);
or U1740 (N_1740,In_1988,In_1035);
nor U1741 (N_1741,In_1063,In_1992);
nor U1742 (N_1742,In_1927,In_2094);
and U1743 (N_1743,In_516,In_2040);
nand U1744 (N_1744,In_2052,In_424);
nor U1745 (N_1745,In_2252,In_97);
nor U1746 (N_1746,In_794,In_8);
nand U1747 (N_1747,In_2371,In_2309);
nand U1748 (N_1748,In_2377,In_243);
or U1749 (N_1749,In_193,In_2370);
nand U1750 (N_1750,In_1213,In_43);
or U1751 (N_1751,In_950,In_159);
or U1752 (N_1752,In_1077,In_1845);
or U1753 (N_1753,In_863,In_68);
nor U1754 (N_1754,In_1121,In_754);
or U1755 (N_1755,In_605,In_2161);
nor U1756 (N_1756,In_861,In_2280);
nor U1757 (N_1757,In_2335,In_1788);
or U1758 (N_1758,In_1716,In_1018);
or U1759 (N_1759,In_384,In_245);
nor U1760 (N_1760,In_1150,In_1630);
xnor U1761 (N_1761,In_675,In_125);
or U1762 (N_1762,In_1923,In_2472);
xor U1763 (N_1763,In_1540,In_625);
nor U1764 (N_1764,In_384,In_840);
nand U1765 (N_1765,In_1418,In_2030);
and U1766 (N_1766,In_1695,In_105);
and U1767 (N_1767,In_2008,In_1263);
and U1768 (N_1768,In_584,In_689);
nor U1769 (N_1769,In_628,In_2417);
nand U1770 (N_1770,In_1415,In_632);
nor U1771 (N_1771,In_759,In_1037);
and U1772 (N_1772,In_61,In_2404);
or U1773 (N_1773,In_1830,In_1314);
or U1774 (N_1774,In_2104,In_1001);
and U1775 (N_1775,In_483,In_1085);
nor U1776 (N_1776,In_336,In_70);
xnor U1777 (N_1777,In_2043,In_2317);
nand U1778 (N_1778,In_572,In_537);
xor U1779 (N_1779,In_2497,In_2041);
xnor U1780 (N_1780,In_1328,In_2051);
and U1781 (N_1781,In_508,In_2014);
nand U1782 (N_1782,In_2249,In_1398);
xnor U1783 (N_1783,In_845,In_1008);
nor U1784 (N_1784,In_1337,In_2415);
nor U1785 (N_1785,In_654,In_1888);
nand U1786 (N_1786,In_197,In_2364);
or U1787 (N_1787,In_1004,In_469);
and U1788 (N_1788,In_1784,In_706);
nor U1789 (N_1789,In_410,In_1539);
nand U1790 (N_1790,In_218,In_1013);
or U1791 (N_1791,In_8,In_1034);
and U1792 (N_1792,In_1068,In_1708);
or U1793 (N_1793,In_2254,In_2057);
nand U1794 (N_1794,In_1695,In_506);
nand U1795 (N_1795,In_1880,In_1643);
and U1796 (N_1796,In_1687,In_1427);
or U1797 (N_1797,In_1601,In_737);
and U1798 (N_1798,In_1288,In_1072);
nand U1799 (N_1799,In_2228,In_636);
nand U1800 (N_1800,In_48,In_1955);
nand U1801 (N_1801,In_1677,In_1171);
nand U1802 (N_1802,In_463,In_2161);
nand U1803 (N_1803,In_793,In_1384);
xnor U1804 (N_1804,In_1606,In_196);
nand U1805 (N_1805,In_1435,In_217);
xor U1806 (N_1806,In_1652,In_714);
nor U1807 (N_1807,In_747,In_1644);
or U1808 (N_1808,In_2089,In_885);
or U1809 (N_1809,In_628,In_1141);
nor U1810 (N_1810,In_1953,In_386);
nor U1811 (N_1811,In_1531,In_1228);
nand U1812 (N_1812,In_892,In_1986);
nor U1813 (N_1813,In_2345,In_1149);
and U1814 (N_1814,In_903,In_1171);
or U1815 (N_1815,In_1660,In_593);
or U1816 (N_1816,In_1456,In_2478);
nor U1817 (N_1817,In_2280,In_271);
or U1818 (N_1818,In_1040,In_1089);
xnor U1819 (N_1819,In_1627,In_1497);
nand U1820 (N_1820,In_1818,In_1565);
nand U1821 (N_1821,In_759,In_10);
nand U1822 (N_1822,In_1010,In_2327);
or U1823 (N_1823,In_1087,In_359);
nor U1824 (N_1824,In_1145,In_1651);
nor U1825 (N_1825,In_936,In_2065);
nor U1826 (N_1826,In_2139,In_302);
and U1827 (N_1827,In_271,In_1760);
and U1828 (N_1828,In_1718,In_493);
nand U1829 (N_1829,In_2407,In_1787);
or U1830 (N_1830,In_220,In_2145);
and U1831 (N_1831,In_2131,In_661);
and U1832 (N_1832,In_969,In_846);
and U1833 (N_1833,In_1168,In_795);
nor U1834 (N_1834,In_1791,In_657);
nor U1835 (N_1835,In_1274,In_2482);
nand U1836 (N_1836,In_2004,In_2402);
or U1837 (N_1837,In_2315,In_1306);
nor U1838 (N_1838,In_1608,In_1784);
nand U1839 (N_1839,In_366,In_1937);
xor U1840 (N_1840,In_2358,In_1052);
and U1841 (N_1841,In_955,In_479);
xnor U1842 (N_1842,In_1636,In_1664);
or U1843 (N_1843,In_1247,In_2378);
nand U1844 (N_1844,In_2413,In_1019);
nor U1845 (N_1845,In_875,In_70);
and U1846 (N_1846,In_526,In_716);
xor U1847 (N_1847,In_42,In_1060);
nor U1848 (N_1848,In_1041,In_668);
nor U1849 (N_1849,In_430,In_668);
and U1850 (N_1850,In_2005,In_809);
nand U1851 (N_1851,In_359,In_1808);
nor U1852 (N_1852,In_368,In_826);
nand U1853 (N_1853,In_606,In_2330);
xor U1854 (N_1854,In_2191,In_1240);
nor U1855 (N_1855,In_1451,In_110);
or U1856 (N_1856,In_569,In_100);
xnor U1857 (N_1857,In_104,In_653);
or U1858 (N_1858,In_218,In_588);
and U1859 (N_1859,In_1683,In_1583);
nor U1860 (N_1860,In_2226,In_1989);
or U1861 (N_1861,In_117,In_664);
or U1862 (N_1862,In_1629,In_2043);
or U1863 (N_1863,In_1588,In_520);
xnor U1864 (N_1864,In_424,In_2055);
and U1865 (N_1865,In_2081,In_1708);
nor U1866 (N_1866,In_12,In_1572);
and U1867 (N_1867,In_170,In_1722);
or U1868 (N_1868,In_905,In_1953);
nor U1869 (N_1869,In_2101,In_2355);
nor U1870 (N_1870,In_2176,In_1049);
and U1871 (N_1871,In_389,In_107);
nand U1872 (N_1872,In_1851,In_1026);
and U1873 (N_1873,In_559,In_2350);
or U1874 (N_1874,In_1652,In_564);
or U1875 (N_1875,In_363,In_2082);
or U1876 (N_1876,In_1009,In_24);
nor U1877 (N_1877,In_536,In_2238);
and U1878 (N_1878,In_2499,In_1111);
or U1879 (N_1879,In_2438,In_386);
and U1880 (N_1880,In_2136,In_914);
or U1881 (N_1881,In_1282,In_70);
and U1882 (N_1882,In_372,In_2223);
and U1883 (N_1883,In_2390,In_293);
nand U1884 (N_1884,In_1712,In_2058);
nand U1885 (N_1885,In_735,In_406);
and U1886 (N_1886,In_1343,In_1732);
nor U1887 (N_1887,In_952,In_2363);
nor U1888 (N_1888,In_2390,In_1341);
and U1889 (N_1889,In_917,In_1925);
or U1890 (N_1890,In_282,In_424);
and U1891 (N_1891,In_1510,In_2143);
nor U1892 (N_1892,In_738,In_2025);
nand U1893 (N_1893,In_811,In_1148);
or U1894 (N_1894,In_1740,In_2095);
nor U1895 (N_1895,In_1175,In_1161);
and U1896 (N_1896,In_485,In_124);
nand U1897 (N_1897,In_189,In_2120);
xor U1898 (N_1898,In_919,In_2377);
or U1899 (N_1899,In_2173,In_335);
nand U1900 (N_1900,In_1338,In_133);
nand U1901 (N_1901,In_2112,In_1351);
and U1902 (N_1902,In_929,In_546);
nand U1903 (N_1903,In_2069,In_1068);
nand U1904 (N_1904,In_2229,In_2171);
or U1905 (N_1905,In_1764,In_21);
and U1906 (N_1906,In_2102,In_616);
nand U1907 (N_1907,In_1717,In_2285);
or U1908 (N_1908,In_1673,In_1731);
nand U1909 (N_1909,In_1791,In_490);
or U1910 (N_1910,In_86,In_1194);
nand U1911 (N_1911,In_252,In_275);
or U1912 (N_1912,In_1928,In_738);
nand U1913 (N_1913,In_1400,In_1455);
or U1914 (N_1914,In_617,In_1771);
or U1915 (N_1915,In_560,In_416);
or U1916 (N_1916,In_1979,In_1005);
nand U1917 (N_1917,In_153,In_898);
nor U1918 (N_1918,In_1952,In_1564);
nand U1919 (N_1919,In_472,In_2323);
nor U1920 (N_1920,In_23,In_685);
or U1921 (N_1921,In_2220,In_1469);
or U1922 (N_1922,In_154,In_252);
and U1923 (N_1923,In_1140,In_2310);
nor U1924 (N_1924,In_1623,In_277);
or U1925 (N_1925,In_532,In_895);
xor U1926 (N_1926,In_802,In_560);
nor U1927 (N_1927,In_2384,In_376);
nand U1928 (N_1928,In_1606,In_872);
and U1929 (N_1929,In_172,In_1225);
or U1930 (N_1930,In_951,In_1607);
and U1931 (N_1931,In_1350,In_732);
or U1932 (N_1932,In_1248,In_1209);
nand U1933 (N_1933,In_470,In_1384);
nand U1934 (N_1934,In_776,In_1459);
or U1935 (N_1935,In_2365,In_911);
or U1936 (N_1936,In_557,In_160);
or U1937 (N_1937,In_1307,In_1159);
nor U1938 (N_1938,In_1342,In_1409);
and U1939 (N_1939,In_2155,In_2454);
nor U1940 (N_1940,In_2079,In_577);
or U1941 (N_1941,In_1421,In_2028);
nand U1942 (N_1942,In_2454,In_2004);
nor U1943 (N_1943,In_991,In_1100);
and U1944 (N_1944,In_61,In_2119);
and U1945 (N_1945,In_1665,In_1441);
and U1946 (N_1946,In_2083,In_1626);
nand U1947 (N_1947,In_1542,In_1442);
and U1948 (N_1948,In_352,In_1325);
or U1949 (N_1949,In_2320,In_287);
or U1950 (N_1950,In_1368,In_2171);
or U1951 (N_1951,In_874,In_1969);
xnor U1952 (N_1952,In_616,In_711);
nor U1953 (N_1953,In_1684,In_1459);
xnor U1954 (N_1954,In_2397,In_495);
or U1955 (N_1955,In_1549,In_1259);
and U1956 (N_1956,In_77,In_1824);
nand U1957 (N_1957,In_883,In_1912);
or U1958 (N_1958,In_1313,In_924);
xnor U1959 (N_1959,In_587,In_718);
or U1960 (N_1960,In_582,In_1251);
nand U1961 (N_1961,In_1142,In_671);
and U1962 (N_1962,In_162,In_1779);
nor U1963 (N_1963,In_5,In_1209);
nand U1964 (N_1964,In_2193,In_737);
nand U1965 (N_1965,In_505,In_1036);
or U1966 (N_1966,In_576,In_7);
nand U1967 (N_1967,In_83,In_2225);
xnor U1968 (N_1968,In_492,In_1845);
and U1969 (N_1969,In_84,In_989);
nor U1970 (N_1970,In_2422,In_1394);
nand U1971 (N_1971,In_2408,In_1684);
or U1972 (N_1972,In_512,In_873);
nor U1973 (N_1973,In_415,In_912);
nand U1974 (N_1974,In_1158,In_1416);
and U1975 (N_1975,In_139,In_595);
nand U1976 (N_1976,In_36,In_1668);
nand U1977 (N_1977,In_724,In_1690);
and U1978 (N_1978,In_194,In_1479);
nor U1979 (N_1979,In_1404,In_1108);
or U1980 (N_1980,In_2077,In_646);
nor U1981 (N_1981,In_108,In_615);
xor U1982 (N_1982,In_765,In_776);
xnor U1983 (N_1983,In_982,In_146);
or U1984 (N_1984,In_562,In_405);
nor U1985 (N_1985,In_1355,In_1);
and U1986 (N_1986,In_1626,In_1404);
xnor U1987 (N_1987,In_1617,In_1353);
and U1988 (N_1988,In_1674,In_2095);
and U1989 (N_1989,In_182,In_1144);
nand U1990 (N_1990,In_2206,In_2485);
nand U1991 (N_1991,In_202,In_178);
or U1992 (N_1992,In_2146,In_406);
and U1993 (N_1993,In_4,In_2007);
and U1994 (N_1994,In_810,In_1277);
nor U1995 (N_1995,In_2072,In_145);
or U1996 (N_1996,In_1515,In_965);
nand U1997 (N_1997,In_1724,In_976);
nor U1998 (N_1998,In_2084,In_1571);
or U1999 (N_1999,In_652,In_110);
and U2000 (N_2000,In_343,In_2384);
or U2001 (N_2001,In_2222,In_1975);
nand U2002 (N_2002,In_1394,In_1035);
nor U2003 (N_2003,In_1895,In_1270);
or U2004 (N_2004,In_67,In_2381);
or U2005 (N_2005,In_548,In_1932);
or U2006 (N_2006,In_2213,In_2400);
or U2007 (N_2007,In_2177,In_1218);
nor U2008 (N_2008,In_872,In_555);
xnor U2009 (N_2009,In_982,In_1521);
and U2010 (N_2010,In_1890,In_1902);
and U2011 (N_2011,In_340,In_330);
nor U2012 (N_2012,In_292,In_1094);
and U2013 (N_2013,In_2235,In_2107);
nand U2014 (N_2014,In_2172,In_120);
nor U2015 (N_2015,In_2176,In_949);
nand U2016 (N_2016,In_1572,In_1478);
xnor U2017 (N_2017,In_2447,In_1572);
or U2018 (N_2018,In_2442,In_252);
and U2019 (N_2019,In_1429,In_2452);
or U2020 (N_2020,In_2444,In_1394);
and U2021 (N_2021,In_1865,In_687);
nand U2022 (N_2022,In_1288,In_1841);
nand U2023 (N_2023,In_66,In_15);
and U2024 (N_2024,In_1607,In_174);
nand U2025 (N_2025,In_808,In_1049);
or U2026 (N_2026,In_792,In_105);
nand U2027 (N_2027,In_958,In_435);
or U2028 (N_2028,In_1318,In_55);
nand U2029 (N_2029,In_1855,In_1249);
or U2030 (N_2030,In_2159,In_671);
and U2031 (N_2031,In_2031,In_1528);
and U2032 (N_2032,In_1582,In_1536);
nand U2033 (N_2033,In_565,In_892);
nand U2034 (N_2034,In_1723,In_1459);
and U2035 (N_2035,In_1643,In_1035);
and U2036 (N_2036,In_1071,In_1718);
nand U2037 (N_2037,In_1616,In_2266);
nand U2038 (N_2038,In_94,In_1526);
nor U2039 (N_2039,In_240,In_1467);
and U2040 (N_2040,In_2391,In_1990);
nand U2041 (N_2041,In_710,In_320);
nand U2042 (N_2042,In_1063,In_1995);
nor U2043 (N_2043,In_885,In_1087);
or U2044 (N_2044,In_1259,In_1493);
or U2045 (N_2045,In_1253,In_1536);
nand U2046 (N_2046,In_97,In_144);
and U2047 (N_2047,In_1858,In_905);
and U2048 (N_2048,In_2145,In_323);
nand U2049 (N_2049,In_589,In_1464);
or U2050 (N_2050,In_1906,In_298);
nand U2051 (N_2051,In_141,In_2360);
or U2052 (N_2052,In_376,In_579);
and U2053 (N_2053,In_406,In_958);
xor U2054 (N_2054,In_1858,In_1267);
and U2055 (N_2055,In_275,In_1058);
nand U2056 (N_2056,In_2051,In_2295);
or U2057 (N_2057,In_1456,In_876);
and U2058 (N_2058,In_784,In_1747);
nor U2059 (N_2059,In_769,In_2194);
nor U2060 (N_2060,In_1685,In_560);
nor U2061 (N_2061,In_627,In_2433);
and U2062 (N_2062,In_80,In_145);
nor U2063 (N_2063,In_626,In_1637);
nor U2064 (N_2064,In_2165,In_658);
and U2065 (N_2065,In_1650,In_1214);
nor U2066 (N_2066,In_1181,In_2195);
nor U2067 (N_2067,In_996,In_637);
nor U2068 (N_2068,In_886,In_1685);
or U2069 (N_2069,In_314,In_2410);
xor U2070 (N_2070,In_1805,In_2185);
nor U2071 (N_2071,In_706,In_2010);
and U2072 (N_2072,In_5,In_2492);
and U2073 (N_2073,In_1269,In_2017);
nand U2074 (N_2074,In_1736,In_1162);
xnor U2075 (N_2075,In_638,In_1794);
and U2076 (N_2076,In_1196,In_1615);
or U2077 (N_2077,In_1727,In_1248);
nor U2078 (N_2078,In_1166,In_505);
nor U2079 (N_2079,In_545,In_1352);
nor U2080 (N_2080,In_299,In_1401);
or U2081 (N_2081,In_1883,In_45);
nor U2082 (N_2082,In_1905,In_2465);
nor U2083 (N_2083,In_801,In_2099);
nor U2084 (N_2084,In_1684,In_1141);
or U2085 (N_2085,In_1598,In_382);
nand U2086 (N_2086,In_1215,In_1660);
and U2087 (N_2087,In_75,In_1166);
or U2088 (N_2088,In_998,In_2096);
nand U2089 (N_2089,In_349,In_1226);
nand U2090 (N_2090,In_1836,In_1083);
and U2091 (N_2091,In_1628,In_511);
or U2092 (N_2092,In_1103,In_8);
nor U2093 (N_2093,In_535,In_2214);
and U2094 (N_2094,In_174,In_1349);
nor U2095 (N_2095,In_2000,In_829);
nand U2096 (N_2096,In_1403,In_845);
and U2097 (N_2097,In_1862,In_2023);
nor U2098 (N_2098,In_2380,In_771);
nand U2099 (N_2099,In_1367,In_2235);
nor U2100 (N_2100,In_387,In_2318);
and U2101 (N_2101,In_784,In_2420);
or U2102 (N_2102,In_2456,In_1284);
nand U2103 (N_2103,In_889,In_885);
and U2104 (N_2104,In_373,In_517);
nand U2105 (N_2105,In_704,In_2378);
or U2106 (N_2106,In_1146,In_291);
nor U2107 (N_2107,In_1390,In_1157);
or U2108 (N_2108,In_1289,In_1135);
nand U2109 (N_2109,In_2051,In_1715);
nand U2110 (N_2110,In_1758,In_746);
nor U2111 (N_2111,In_52,In_2078);
nor U2112 (N_2112,In_168,In_955);
nor U2113 (N_2113,In_1186,In_2290);
nor U2114 (N_2114,In_1637,In_1358);
nor U2115 (N_2115,In_341,In_369);
nand U2116 (N_2116,In_1705,In_1001);
nand U2117 (N_2117,In_1692,In_1589);
xor U2118 (N_2118,In_2230,In_1674);
xnor U2119 (N_2119,In_1146,In_742);
nor U2120 (N_2120,In_1072,In_215);
or U2121 (N_2121,In_1906,In_1698);
nor U2122 (N_2122,In_1377,In_1343);
nor U2123 (N_2123,In_1017,In_1003);
or U2124 (N_2124,In_273,In_2331);
nand U2125 (N_2125,In_730,In_694);
xor U2126 (N_2126,In_2187,In_1715);
nor U2127 (N_2127,In_2440,In_466);
nand U2128 (N_2128,In_1879,In_1262);
nand U2129 (N_2129,In_936,In_2051);
and U2130 (N_2130,In_2326,In_504);
or U2131 (N_2131,In_1639,In_2403);
nand U2132 (N_2132,In_1128,In_1118);
nand U2133 (N_2133,In_2236,In_619);
nor U2134 (N_2134,In_466,In_1228);
or U2135 (N_2135,In_932,In_15);
nand U2136 (N_2136,In_1440,In_2257);
and U2137 (N_2137,In_1539,In_2207);
and U2138 (N_2138,In_1170,In_260);
or U2139 (N_2139,In_283,In_710);
nand U2140 (N_2140,In_2310,In_1829);
or U2141 (N_2141,In_1066,In_73);
nor U2142 (N_2142,In_415,In_2420);
nor U2143 (N_2143,In_1061,In_2079);
nand U2144 (N_2144,In_2495,In_1287);
or U2145 (N_2145,In_1548,In_1228);
nor U2146 (N_2146,In_1578,In_2371);
or U2147 (N_2147,In_1081,In_839);
nand U2148 (N_2148,In_1799,In_2075);
nand U2149 (N_2149,In_1423,In_956);
or U2150 (N_2150,In_2069,In_1943);
nand U2151 (N_2151,In_1353,In_1223);
or U2152 (N_2152,In_1481,In_690);
and U2153 (N_2153,In_2039,In_2482);
or U2154 (N_2154,In_475,In_268);
or U2155 (N_2155,In_992,In_818);
and U2156 (N_2156,In_895,In_1984);
nor U2157 (N_2157,In_858,In_420);
and U2158 (N_2158,In_1951,In_2334);
xor U2159 (N_2159,In_1499,In_657);
nand U2160 (N_2160,In_1446,In_1958);
and U2161 (N_2161,In_999,In_509);
and U2162 (N_2162,In_0,In_1495);
xnor U2163 (N_2163,In_1459,In_357);
nor U2164 (N_2164,In_426,In_452);
or U2165 (N_2165,In_893,In_2113);
xnor U2166 (N_2166,In_777,In_326);
xnor U2167 (N_2167,In_2454,In_630);
and U2168 (N_2168,In_1665,In_533);
or U2169 (N_2169,In_574,In_549);
and U2170 (N_2170,In_198,In_2152);
or U2171 (N_2171,In_1830,In_1612);
and U2172 (N_2172,In_923,In_1632);
or U2173 (N_2173,In_1465,In_1585);
nand U2174 (N_2174,In_915,In_281);
or U2175 (N_2175,In_1417,In_2344);
and U2176 (N_2176,In_1538,In_373);
and U2177 (N_2177,In_2290,In_990);
nand U2178 (N_2178,In_1077,In_231);
nand U2179 (N_2179,In_1237,In_1712);
and U2180 (N_2180,In_1751,In_426);
nor U2181 (N_2181,In_1804,In_1756);
or U2182 (N_2182,In_1808,In_51);
nor U2183 (N_2183,In_1368,In_95);
and U2184 (N_2184,In_963,In_1516);
nand U2185 (N_2185,In_1436,In_1972);
nor U2186 (N_2186,In_719,In_1406);
nor U2187 (N_2187,In_1122,In_509);
and U2188 (N_2188,In_1851,In_1315);
xnor U2189 (N_2189,In_1651,In_1585);
or U2190 (N_2190,In_674,In_601);
and U2191 (N_2191,In_1226,In_354);
nand U2192 (N_2192,In_1570,In_1962);
nand U2193 (N_2193,In_1480,In_738);
nor U2194 (N_2194,In_522,In_1310);
nand U2195 (N_2195,In_979,In_1264);
nand U2196 (N_2196,In_402,In_2151);
and U2197 (N_2197,In_1334,In_255);
and U2198 (N_2198,In_847,In_366);
and U2199 (N_2199,In_238,In_638);
or U2200 (N_2200,In_2269,In_912);
xor U2201 (N_2201,In_151,In_1355);
nand U2202 (N_2202,In_703,In_831);
xor U2203 (N_2203,In_783,In_701);
nor U2204 (N_2204,In_168,In_274);
and U2205 (N_2205,In_1972,In_1570);
and U2206 (N_2206,In_90,In_2488);
nor U2207 (N_2207,In_240,In_1478);
xor U2208 (N_2208,In_27,In_45);
xor U2209 (N_2209,In_485,In_642);
and U2210 (N_2210,In_561,In_542);
nor U2211 (N_2211,In_553,In_2053);
nand U2212 (N_2212,In_1242,In_1538);
nand U2213 (N_2213,In_727,In_1864);
and U2214 (N_2214,In_2072,In_176);
nand U2215 (N_2215,In_14,In_276);
or U2216 (N_2216,In_1591,In_1682);
and U2217 (N_2217,In_1938,In_246);
xor U2218 (N_2218,In_1672,In_1343);
or U2219 (N_2219,In_1184,In_1995);
xnor U2220 (N_2220,In_562,In_1503);
nor U2221 (N_2221,In_1164,In_768);
and U2222 (N_2222,In_946,In_172);
nor U2223 (N_2223,In_2258,In_397);
nor U2224 (N_2224,In_1115,In_1385);
nand U2225 (N_2225,In_90,In_662);
and U2226 (N_2226,In_1516,In_1088);
or U2227 (N_2227,In_14,In_1425);
and U2228 (N_2228,In_1577,In_2135);
and U2229 (N_2229,In_1871,In_2241);
and U2230 (N_2230,In_1818,In_0);
nand U2231 (N_2231,In_2284,In_2004);
nand U2232 (N_2232,In_1257,In_1781);
nand U2233 (N_2233,In_1512,In_1689);
or U2234 (N_2234,In_1036,In_1351);
nor U2235 (N_2235,In_161,In_1917);
or U2236 (N_2236,In_951,In_85);
or U2237 (N_2237,In_1514,In_1185);
and U2238 (N_2238,In_82,In_1564);
and U2239 (N_2239,In_2129,In_1530);
nor U2240 (N_2240,In_107,In_2113);
nor U2241 (N_2241,In_6,In_2426);
or U2242 (N_2242,In_1610,In_324);
or U2243 (N_2243,In_506,In_1007);
or U2244 (N_2244,In_2457,In_2191);
nand U2245 (N_2245,In_280,In_761);
nor U2246 (N_2246,In_1530,In_2259);
nor U2247 (N_2247,In_1366,In_2039);
xnor U2248 (N_2248,In_1527,In_2429);
and U2249 (N_2249,In_805,In_208);
and U2250 (N_2250,In_2401,In_1304);
or U2251 (N_2251,In_286,In_1679);
or U2252 (N_2252,In_2237,In_794);
nor U2253 (N_2253,In_1739,In_2349);
xnor U2254 (N_2254,In_688,In_1005);
and U2255 (N_2255,In_1100,In_1774);
nand U2256 (N_2256,In_776,In_1799);
and U2257 (N_2257,In_778,In_1681);
and U2258 (N_2258,In_1111,In_1556);
nor U2259 (N_2259,In_738,In_610);
nor U2260 (N_2260,In_2056,In_1491);
nand U2261 (N_2261,In_1063,In_1685);
or U2262 (N_2262,In_566,In_1008);
nor U2263 (N_2263,In_175,In_720);
or U2264 (N_2264,In_453,In_253);
nor U2265 (N_2265,In_2128,In_1554);
nand U2266 (N_2266,In_1178,In_636);
or U2267 (N_2267,In_2431,In_355);
and U2268 (N_2268,In_153,In_901);
nand U2269 (N_2269,In_604,In_2403);
xor U2270 (N_2270,In_1410,In_555);
xnor U2271 (N_2271,In_1452,In_2492);
nor U2272 (N_2272,In_1293,In_1996);
nand U2273 (N_2273,In_1490,In_1380);
nor U2274 (N_2274,In_959,In_699);
xor U2275 (N_2275,In_274,In_1108);
or U2276 (N_2276,In_1442,In_982);
and U2277 (N_2277,In_1107,In_1771);
or U2278 (N_2278,In_1049,In_2221);
nor U2279 (N_2279,In_1256,In_278);
and U2280 (N_2280,In_1518,In_2292);
and U2281 (N_2281,In_820,In_263);
nand U2282 (N_2282,In_410,In_1293);
or U2283 (N_2283,In_669,In_1373);
or U2284 (N_2284,In_360,In_477);
nor U2285 (N_2285,In_732,In_1158);
nor U2286 (N_2286,In_1674,In_1453);
nand U2287 (N_2287,In_2355,In_1954);
nor U2288 (N_2288,In_603,In_2369);
and U2289 (N_2289,In_2092,In_2043);
nor U2290 (N_2290,In_628,In_2155);
nor U2291 (N_2291,In_575,In_984);
and U2292 (N_2292,In_1403,In_849);
xnor U2293 (N_2293,In_1191,In_1632);
nand U2294 (N_2294,In_1251,In_377);
nand U2295 (N_2295,In_1782,In_499);
nand U2296 (N_2296,In_814,In_1171);
nor U2297 (N_2297,In_1628,In_1313);
and U2298 (N_2298,In_26,In_850);
and U2299 (N_2299,In_1248,In_130);
nand U2300 (N_2300,In_1513,In_1014);
nand U2301 (N_2301,In_1360,In_957);
nor U2302 (N_2302,In_1417,In_1212);
nor U2303 (N_2303,In_306,In_1369);
nand U2304 (N_2304,In_2259,In_642);
and U2305 (N_2305,In_1777,In_1085);
nor U2306 (N_2306,In_585,In_797);
and U2307 (N_2307,In_1496,In_2248);
or U2308 (N_2308,In_1635,In_1390);
and U2309 (N_2309,In_135,In_670);
nand U2310 (N_2310,In_2302,In_915);
and U2311 (N_2311,In_1668,In_519);
nor U2312 (N_2312,In_2045,In_1474);
and U2313 (N_2313,In_1276,In_1348);
nor U2314 (N_2314,In_871,In_1607);
nor U2315 (N_2315,In_386,In_165);
nor U2316 (N_2316,In_274,In_5);
nand U2317 (N_2317,In_174,In_2334);
nand U2318 (N_2318,In_191,In_893);
and U2319 (N_2319,In_1485,In_931);
or U2320 (N_2320,In_621,In_2362);
or U2321 (N_2321,In_338,In_2145);
nand U2322 (N_2322,In_333,In_1680);
nor U2323 (N_2323,In_1517,In_2230);
nand U2324 (N_2324,In_447,In_1282);
and U2325 (N_2325,In_1890,In_1850);
or U2326 (N_2326,In_1628,In_1468);
and U2327 (N_2327,In_758,In_1889);
nand U2328 (N_2328,In_66,In_1845);
nand U2329 (N_2329,In_2139,In_636);
nor U2330 (N_2330,In_1031,In_1528);
nand U2331 (N_2331,In_24,In_53);
and U2332 (N_2332,In_2420,In_1825);
nand U2333 (N_2333,In_209,In_596);
or U2334 (N_2334,In_1286,In_142);
nand U2335 (N_2335,In_1762,In_2360);
xor U2336 (N_2336,In_1231,In_1053);
nand U2337 (N_2337,In_1780,In_379);
nand U2338 (N_2338,In_2095,In_1102);
or U2339 (N_2339,In_2234,In_1837);
or U2340 (N_2340,In_280,In_424);
nand U2341 (N_2341,In_237,In_2164);
nand U2342 (N_2342,In_1125,In_1853);
xor U2343 (N_2343,In_1191,In_2391);
xnor U2344 (N_2344,In_129,In_591);
and U2345 (N_2345,In_2025,In_1267);
nor U2346 (N_2346,In_879,In_1225);
and U2347 (N_2347,In_837,In_1192);
nor U2348 (N_2348,In_401,In_964);
and U2349 (N_2349,In_1487,In_279);
xnor U2350 (N_2350,In_98,In_2046);
nor U2351 (N_2351,In_170,In_1145);
nor U2352 (N_2352,In_2171,In_308);
nor U2353 (N_2353,In_2401,In_828);
or U2354 (N_2354,In_1623,In_50);
xnor U2355 (N_2355,In_1685,In_1642);
and U2356 (N_2356,In_2208,In_546);
nand U2357 (N_2357,In_807,In_203);
and U2358 (N_2358,In_1510,In_265);
and U2359 (N_2359,In_176,In_968);
and U2360 (N_2360,In_775,In_1977);
nor U2361 (N_2361,In_1692,In_1149);
nand U2362 (N_2362,In_262,In_21);
or U2363 (N_2363,In_122,In_1721);
nand U2364 (N_2364,In_2292,In_597);
and U2365 (N_2365,In_196,In_615);
or U2366 (N_2366,In_1894,In_621);
and U2367 (N_2367,In_2268,In_1315);
nand U2368 (N_2368,In_650,In_1070);
nor U2369 (N_2369,In_1263,In_880);
or U2370 (N_2370,In_168,In_84);
or U2371 (N_2371,In_1397,In_151);
and U2372 (N_2372,In_1052,In_620);
or U2373 (N_2373,In_1836,In_691);
xor U2374 (N_2374,In_2166,In_690);
nand U2375 (N_2375,In_1275,In_1772);
or U2376 (N_2376,In_792,In_100);
xnor U2377 (N_2377,In_2060,In_205);
nor U2378 (N_2378,In_1769,In_1691);
or U2379 (N_2379,In_2012,In_1080);
nor U2380 (N_2380,In_858,In_1627);
and U2381 (N_2381,In_1822,In_1900);
nor U2382 (N_2382,In_1225,In_105);
nand U2383 (N_2383,In_1484,In_245);
xnor U2384 (N_2384,In_275,In_1987);
nor U2385 (N_2385,In_2167,In_209);
nor U2386 (N_2386,In_258,In_634);
nor U2387 (N_2387,In_286,In_927);
nor U2388 (N_2388,In_1070,In_1986);
xor U2389 (N_2389,In_885,In_1339);
nor U2390 (N_2390,In_1272,In_8);
and U2391 (N_2391,In_505,In_1429);
and U2392 (N_2392,In_1558,In_287);
and U2393 (N_2393,In_278,In_2192);
nand U2394 (N_2394,In_2295,In_1282);
nand U2395 (N_2395,In_2082,In_551);
or U2396 (N_2396,In_2205,In_441);
nor U2397 (N_2397,In_2380,In_1439);
nand U2398 (N_2398,In_74,In_235);
or U2399 (N_2399,In_1808,In_1902);
xor U2400 (N_2400,In_2400,In_2391);
or U2401 (N_2401,In_1070,In_2097);
nand U2402 (N_2402,In_145,In_611);
nand U2403 (N_2403,In_1776,In_567);
nor U2404 (N_2404,In_2004,In_962);
xnor U2405 (N_2405,In_1209,In_1058);
or U2406 (N_2406,In_2210,In_354);
nor U2407 (N_2407,In_1684,In_720);
xnor U2408 (N_2408,In_1597,In_892);
nor U2409 (N_2409,In_2021,In_411);
nor U2410 (N_2410,In_1969,In_1219);
nand U2411 (N_2411,In_259,In_74);
or U2412 (N_2412,In_95,In_1051);
xor U2413 (N_2413,In_322,In_1534);
nor U2414 (N_2414,In_430,In_1931);
or U2415 (N_2415,In_2216,In_62);
nor U2416 (N_2416,In_2451,In_2069);
nor U2417 (N_2417,In_1893,In_1085);
nor U2418 (N_2418,In_1146,In_1218);
and U2419 (N_2419,In_809,In_1609);
xnor U2420 (N_2420,In_103,In_307);
and U2421 (N_2421,In_293,In_774);
or U2422 (N_2422,In_1863,In_1206);
and U2423 (N_2423,In_215,In_1335);
nor U2424 (N_2424,In_1417,In_2423);
xor U2425 (N_2425,In_1827,In_2380);
and U2426 (N_2426,In_1285,In_312);
or U2427 (N_2427,In_357,In_490);
nand U2428 (N_2428,In_331,In_1788);
nor U2429 (N_2429,In_2366,In_542);
and U2430 (N_2430,In_1844,In_1125);
or U2431 (N_2431,In_1109,In_794);
and U2432 (N_2432,In_1184,In_454);
nand U2433 (N_2433,In_1464,In_141);
nor U2434 (N_2434,In_1422,In_1099);
or U2435 (N_2435,In_882,In_1365);
or U2436 (N_2436,In_749,In_2048);
nor U2437 (N_2437,In_1186,In_1095);
xor U2438 (N_2438,In_2219,In_661);
or U2439 (N_2439,In_741,In_390);
nand U2440 (N_2440,In_1639,In_1637);
or U2441 (N_2441,In_1729,In_51);
nor U2442 (N_2442,In_1199,In_1178);
and U2443 (N_2443,In_256,In_1845);
nand U2444 (N_2444,In_978,In_1264);
and U2445 (N_2445,In_1472,In_1520);
and U2446 (N_2446,In_1481,In_266);
or U2447 (N_2447,In_2042,In_657);
or U2448 (N_2448,In_2156,In_2153);
nor U2449 (N_2449,In_2447,In_288);
or U2450 (N_2450,In_75,In_1578);
nand U2451 (N_2451,In_294,In_1488);
nor U2452 (N_2452,In_1172,In_1542);
or U2453 (N_2453,In_1970,In_472);
or U2454 (N_2454,In_1931,In_697);
nor U2455 (N_2455,In_430,In_2116);
and U2456 (N_2456,In_1575,In_392);
xor U2457 (N_2457,In_504,In_1819);
and U2458 (N_2458,In_1473,In_313);
nor U2459 (N_2459,In_988,In_240);
nor U2460 (N_2460,In_453,In_2238);
and U2461 (N_2461,In_1130,In_2125);
nor U2462 (N_2462,In_1885,In_1957);
nand U2463 (N_2463,In_2113,In_1578);
or U2464 (N_2464,In_1114,In_2067);
nor U2465 (N_2465,In_2274,In_1578);
nor U2466 (N_2466,In_864,In_360);
and U2467 (N_2467,In_1079,In_1715);
or U2468 (N_2468,In_1451,In_1718);
nand U2469 (N_2469,In_814,In_2311);
xnor U2470 (N_2470,In_2235,In_727);
nor U2471 (N_2471,In_989,In_298);
nand U2472 (N_2472,In_1581,In_1169);
nor U2473 (N_2473,In_10,In_1504);
nand U2474 (N_2474,In_119,In_1207);
nor U2475 (N_2475,In_2075,In_931);
nor U2476 (N_2476,In_1661,In_402);
nand U2477 (N_2477,In_1340,In_1245);
and U2478 (N_2478,In_2328,In_1136);
and U2479 (N_2479,In_305,In_923);
and U2480 (N_2480,In_995,In_1177);
and U2481 (N_2481,In_2417,In_2084);
xor U2482 (N_2482,In_2265,In_1211);
or U2483 (N_2483,In_1181,In_2176);
nor U2484 (N_2484,In_1130,In_414);
nand U2485 (N_2485,In_917,In_522);
nand U2486 (N_2486,In_2084,In_1045);
nand U2487 (N_2487,In_973,In_1527);
or U2488 (N_2488,In_325,In_2473);
nor U2489 (N_2489,In_381,In_29);
or U2490 (N_2490,In_1183,In_1207);
nor U2491 (N_2491,In_2024,In_566);
nor U2492 (N_2492,In_913,In_2342);
nand U2493 (N_2493,In_1143,In_501);
and U2494 (N_2494,In_941,In_2087);
nor U2495 (N_2495,In_106,In_262);
and U2496 (N_2496,In_330,In_1102);
and U2497 (N_2497,In_2445,In_1877);
and U2498 (N_2498,In_1036,In_2139);
nand U2499 (N_2499,In_259,In_2248);
and U2500 (N_2500,In_817,In_541);
xnor U2501 (N_2501,In_2025,In_2208);
nand U2502 (N_2502,In_1864,In_286);
and U2503 (N_2503,In_2008,In_26);
xor U2504 (N_2504,In_2331,In_54);
nor U2505 (N_2505,In_1303,In_1149);
and U2506 (N_2506,In_1049,In_1403);
xnor U2507 (N_2507,In_1797,In_2185);
and U2508 (N_2508,In_117,In_2059);
and U2509 (N_2509,In_143,In_1314);
and U2510 (N_2510,In_543,In_462);
nor U2511 (N_2511,In_2203,In_503);
or U2512 (N_2512,In_1618,In_2475);
and U2513 (N_2513,In_6,In_1685);
xnor U2514 (N_2514,In_41,In_1267);
and U2515 (N_2515,In_2097,In_93);
nand U2516 (N_2516,In_1272,In_970);
or U2517 (N_2517,In_1873,In_999);
or U2518 (N_2518,In_1514,In_2176);
nor U2519 (N_2519,In_1918,In_2308);
xor U2520 (N_2520,In_2378,In_1320);
or U2521 (N_2521,In_1636,In_311);
or U2522 (N_2522,In_234,In_945);
nand U2523 (N_2523,In_519,In_979);
nor U2524 (N_2524,In_620,In_2469);
or U2525 (N_2525,In_571,In_2033);
nand U2526 (N_2526,In_382,In_1048);
and U2527 (N_2527,In_617,In_1363);
nor U2528 (N_2528,In_1488,In_1403);
nand U2529 (N_2529,In_835,In_105);
or U2530 (N_2530,In_640,In_2371);
or U2531 (N_2531,In_313,In_779);
or U2532 (N_2532,In_2312,In_369);
or U2533 (N_2533,In_1962,In_1634);
and U2534 (N_2534,In_915,In_2331);
or U2535 (N_2535,In_120,In_458);
nor U2536 (N_2536,In_380,In_1633);
xnor U2537 (N_2537,In_297,In_2010);
nor U2538 (N_2538,In_1631,In_732);
and U2539 (N_2539,In_1344,In_549);
or U2540 (N_2540,In_2244,In_2286);
and U2541 (N_2541,In_380,In_1033);
xor U2542 (N_2542,In_2162,In_1981);
nand U2543 (N_2543,In_208,In_1123);
and U2544 (N_2544,In_2225,In_775);
nor U2545 (N_2545,In_2290,In_2474);
nor U2546 (N_2546,In_2068,In_1201);
and U2547 (N_2547,In_256,In_765);
or U2548 (N_2548,In_2394,In_1042);
or U2549 (N_2549,In_1247,In_739);
and U2550 (N_2550,In_2301,In_2095);
or U2551 (N_2551,In_693,In_1288);
or U2552 (N_2552,In_1589,In_2346);
or U2553 (N_2553,In_637,In_1182);
nor U2554 (N_2554,In_138,In_953);
or U2555 (N_2555,In_128,In_1628);
or U2556 (N_2556,In_57,In_1121);
nor U2557 (N_2557,In_845,In_522);
nand U2558 (N_2558,In_732,In_2418);
or U2559 (N_2559,In_56,In_616);
and U2560 (N_2560,In_1284,In_1161);
and U2561 (N_2561,In_1112,In_60);
or U2562 (N_2562,In_1996,In_1520);
nor U2563 (N_2563,In_749,In_1871);
or U2564 (N_2564,In_402,In_495);
or U2565 (N_2565,In_16,In_2411);
or U2566 (N_2566,In_1076,In_1477);
and U2567 (N_2567,In_1976,In_1352);
xor U2568 (N_2568,In_148,In_726);
or U2569 (N_2569,In_1609,In_2005);
nand U2570 (N_2570,In_2160,In_1473);
or U2571 (N_2571,In_1866,In_762);
or U2572 (N_2572,In_1486,In_62);
and U2573 (N_2573,In_519,In_1923);
xor U2574 (N_2574,In_1159,In_1337);
or U2575 (N_2575,In_428,In_2195);
and U2576 (N_2576,In_493,In_2180);
and U2577 (N_2577,In_482,In_74);
and U2578 (N_2578,In_466,In_1860);
or U2579 (N_2579,In_1660,In_2126);
nand U2580 (N_2580,In_2496,In_241);
nand U2581 (N_2581,In_365,In_2154);
or U2582 (N_2582,In_774,In_519);
nand U2583 (N_2583,In_1110,In_1893);
nor U2584 (N_2584,In_2407,In_2125);
and U2585 (N_2585,In_1544,In_1126);
or U2586 (N_2586,In_1614,In_1125);
nand U2587 (N_2587,In_2169,In_1523);
nor U2588 (N_2588,In_1937,In_124);
nand U2589 (N_2589,In_211,In_1343);
or U2590 (N_2590,In_34,In_358);
nand U2591 (N_2591,In_1502,In_1734);
xor U2592 (N_2592,In_360,In_1272);
nor U2593 (N_2593,In_544,In_1027);
and U2594 (N_2594,In_2099,In_1336);
and U2595 (N_2595,In_393,In_758);
and U2596 (N_2596,In_1532,In_985);
or U2597 (N_2597,In_796,In_1955);
nand U2598 (N_2598,In_2388,In_1649);
nor U2599 (N_2599,In_1427,In_1503);
or U2600 (N_2600,In_916,In_461);
xnor U2601 (N_2601,In_896,In_2208);
or U2602 (N_2602,In_551,In_2399);
xnor U2603 (N_2603,In_1664,In_1269);
and U2604 (N_2604,In_2237,In_1342);
nand U2605 (N_2605,In_464,In_577);
or U2606 (N_2606,In_1774,In_370);
nor U2607 (N_2607,In_1265,In_1353);
nand U2608 (N_2608,In_2374,In_2266);
or U2609 (N_2609,In_1375,In_157);
nor U2610 (N_2610,In_909,In_1892);
and U2611 (N_2611,In_797,In_880);
nor U2612 (N_2612,In_1104,In_1486);
and U2613 (N_2613,In_2415,In_1545);
and U2614 (N_2614,In_2189,In_1804);
and U2615 (N_2615,In_967,In_347);
xnor U2616 (N_2616,In_1490,In_2249);
nor U2617 (N_2617,In_1302,In_1762);
nor U2618 (N_2618,In_101,In_802);
nor U2619 (N_2619,In_1711,In_870);
nand U2620 (N_2620,In_2369,In_1025);
xor U2621 (N_2621,In_1090,In_519);
nand U2622 (N_2622,In_1180,In_833);
and U2623 (N_2623,In_904,In_908);
or U2624 (N_2624,In_747,In_671);
and U2625 (N_2625,In_78,In_972);
or U2626 (N_2626,In_1261,In_868);
nor U2627 (N_2627,In_1222,In_1726);
and U2628 (N_2628,In_393,In_2102);
nand U2629 (N_2629,In_2075,In_1881);
and U2630 (N_2630,In_692,In_504);
nor U2631 (N_2631,In_1922,In_42);
or U2632 (N_2632,In_1578,In_1575);
or U2633 (N_2633,In_1009,In_2431);
nor U2634 (N_2634,In_1564,In_784);
nand U2635 (N_2635,In_1984,In_828);
nor U2636 (N_2636,In_1284,In_1428);
nand U2637 (N_2637,In_1729,In_1988);
and U2638 (N_2638,In_1566,In_2410);
xnor U2639 (N_2639,In_799,In_1700);
or U2640 (N_2640,In_2470,In_2492);
nor U2641 (N_2641,In_1052,In_603);
nand U2642 (N_2642,In_366,In_2442);
and U2643 (N_2643,In_1558,In_1802);
xnor U2644 (N_2644,In_2025,In_889);
nand U2645 (N_2645,In_1702,In_26);
and U2646 (N_2646,In_883,In_107);
or U2647 (N_2647,In_2,In_450);
nor U2648 (N_2648,In_2206,In_146);
nand U2649 (N_2649,In_1492,In_107);
nand U2650 (N_2650,In_623,In_1733);
nand U2651 (N_2651,In_1813,In_185);
nand U2652 (N_2652,In_242,In_1469);
and U2653 (N_2653,In_1484,In_614);
nand U2654 (N_2654,In_1854,In_119);
or U2655 (N_2655,In_1553,In_2442);
nand U2656 (N_2656,In_742,In_76);
xor U2657 (N_2657,In_121,In_2368);
xor U2658 (N_2658,In_33,In_611);
nand U2659 (N_2659,In_2287,In_298);
or U2660 (N_2660,In_1500,In_1899);
nor U2661 (N_2661,In_1787,In_655);
or U2662 (N_2662,In_489,In_984);
nor U2663 (N_2663,In_2058,In_198);
nand U2664 (N_2664,In_1584,In_1471);
nand U2665 (N_2665,In_496,In_1148);
nor U2666 (N_2666,In_1230,In_2239);
nand U2667 (N_2667,In_1749,In_1600);
nor U2668 (N_2668,In_1188,In_1556);
nor U2669 (N_2669,In_686,In_255);
nor U2670 (N_2670,In_87,In_2384);
nor U2671 (N_2671,In_2350,In_2034);
nand U2672 (N_2672,In_328,In_525);
or U2673 (N_2673,In_2307,In_1604);
or U2674 (N_2674,In_18,In_467);
or U2675 (N_2675,In_175,In_1269);
nand U2676 (N_2676,In_1718,In_1433);
nand U2677 (N_2677,In_984,In_1482);
and U2678 (N_2678,In_2124,In_2121);
and U2679 (N_2679,In_22,In_1195);
nor U2680 (N_2680,In_442,In_706);
nor U2681 (N_2681,In_2113,In_2340);
and U2682 (N_2682,In_1424,In_262);
and U2683 (N_2683,In_2437,In_2375);
nand U2684 (N_2684,In_1290,In_249);
and U2685 (N_2685,In_256,In_2132);
and U2686 (N_2686,In_410,In_1957);
and U2687 (N_2687,In_610,In_2341);
or U2688 (N_2688,In_101,In_1556);
and U2689 (N_2689,In_819,In_2419);
nor U2690 (N_2690,In_251,In_981);
and U2691 (N_2691,In_2484,In_902);
xnor U2692 (N_2692,In_2142,In_14);
and U2693 (N_2693,In_2091,In_533);
nand U2694 (N_2694,In_1533,In_289);
and U2695 (N_2695,In_1753,In_1947);
and U2696 (N_2696,In_515,In_306);
and U2697 (N_2697,In_329,In_76);
xnor U2698 (N_2698,In_1524,In_966);
nand U2699 (N_2699,In_368,In_1330);
or U2700 (N_2700,In_2389,In_1789);
nor U2701 (N_2701,In_303,In_1670);
or U2702 (N_2702,In_171,In_2347);
xnor U2703 (N_2703,In_2495,In_517);
nor U2704 (N_2704,In_240,In_251);
nor U2705 (N_2705,In_1937,In_769);
or U2706 (N_2706,In_1721,In_1258);
nor U2707 (N_2707,In_262,In_264);
and U2708 (N_2708,In_147,In_39);
or U2709 (N_2709,In_1205,In_1492);
and U2710 (N_2710,In_1297,In_2487);
and U2711 (N_2711,In_924,In_707);
nand U2712 (N_2712,In_1182,In_1591);
nor U2713 (N_2713,In_588,In_2089);
or U2714 (N_2714,In_1038,In_179);
or U2715 (N_2715,In_1809,In_320);
or U2716 (N_2716,In_909,In_203);
or U2717 (N_2717,In_2411,In_1469);
or U2718 (N_2718,In_1532,In_1517);
nand U2719 (N_2719,In_177,In_557);
nand U2720 (N_2720,In_748,In_412);
nor U2721 (N_2721,In_1805,In_2246);
xnor U2722 (N_2722,In_746,In_493);
or U2723 (N_2723,In_1965,In_714);
or U2724 (N_2724,In_352,In_29);
or U2725 (N_2725,In_737,In_2240);
and U2726 (N_2726,In_733,In_835);
nor U2727 (N_2727,In_1101,In_427);
nand U2728 (N_2728,In_231,In_217);
and U2729 (N_2729,In_2377,In_2117);
and U2730 (N_2730,In_98,In_327);
nand U2731 (N_2731,In_600,In_2481);
nor U2732 (N_2732,In_322,In_1910);
and U2733 (N_2733,In_519,In_1621);
nand U2734 (N_2734,In_1791,In_2000);
nand U2735 (N_2735,In_1823,In_1835);
xnor U2736 (N_2736,In_1663,In_1028);
xnor U2737 (N_2737,In_1043,In_1197);
and U2738 (N_2738,In_742,In_195);
nor U2739 (N_2739,In_703,In_673);
nand U2740 (N_2740,In_2393,In_2223);
nor U2741 (N_2741,In_1792,In_1167);
nand U2742 (N_2742,In_919,In_41);
and U2743 (N_2743,In_59,In_2254);
or U2744 (N_2744,In_178,In_2015);
and U2745 (N_2745,In_641,In_380);
or U2746 (N_2746,In_395,In_1214);
xor U2747 (N_2747,In_1467,In_400);
nand U2748 (N_2748,In_2076,In_813);
xor U2749 (N_2749,In_1227,In_1886);
or U2750 (N_2750,In_811,In_1270);
nand U2751 (N_2751,In_2061,In_1538);
nand U2752 (N_2752,In_1838,In_2442);
or U2753 (N_2753,In_668,In_578);
nand U2754 (N_2754,In_2349,In_1560);
and U2755 (N_2755,In_1637,In_587);
or U2756 (N_2756,In_106,In_1780);
or U2757 (N_2757,In_496,In_1701);
and U2758 (N_2758,In_379,In_850);
and U2759 (N_2759,In_2435,In_1639);
nor U2760 (N_2760,In_2118,In_1353);
nor U2761 (N_2761,In_26,In_1457);
nor U2762 (N_2762,In_954,In_1237);
nand U2763 (N_2763,In_2452,In_2024);
or U2764 (N_2764,In_1353,In_236);
and U2765 (N_2765,In_2363,In_1385);
xor U2766 (N_2766,In_661,In_1345);
nor U2767 (N_2767,In_837,In_1258);
xor U2768 (N_2768,In_1277,In_1459);
and U2769 (N_2769,In_784,In_1946);
nand U2770 (N_2770,In_1776,In_726);
or U2771 (N_2771,In_276,In_1130);
nand U2772 (N_2772,In_1553,In_1082);
nor U2773 (N_2773,In_1214,In_2026);
nor U2774 (N_2774,In_1117,In_2195);
or U2775 (N_2775,In_1645,In_397);
or U2776 (N_2776,In_260,In_1537);
xnor U2777 (N_2777,In_1659,In_2197);
or U2778 (N_2778,In_2213,In_2045);
and U2779 (N_2779,In_1070,In_1601);
nor U2780 (N_2780,In_288,In_902);
or U2781 (N_2781,In_1689,In_10);
and U2782 (N_2782,In_465,In_1744);
or U2783 (N_2783,In_1692,In_800);
or U2784 (N_2784,In_1282,In_1185);
and U2785 (N_2785,In_95,In_753);
nor U2786 (N_2786,In_1947,In_1873);
nor U2787 (N_2787,In_209,In_1387);
or U2788 (N_2788,In_855,In_379);
and U2789 (N_2789,In_1963,In_519);
or U2790 (N_2790,In_39,In_2150);
and U2791 (N_2791,In_1381,In_596);
or U2792 (N_2792,In_1696,In_834);
nor U2793 (N_2793,In_1301,In_143);
xor U2794 (N_2794,In_2244,In_1005);
xnor U2795 (N_2795,In_699,In_1951);
and U2796 (N_2796,In_2213,In_2397);
nor U2797 (N_2797,In_2414,In_1304);
nand U2798 (N_2798,In_1259,In_1383);
or U2799 (N_2799,In_880,In_1765);
and U2800 (N_2800,In_1835,In_949);
nand U2801 (N_2801,In_2074,In_1263);
and U2802 (N_2802,In_1199,In_1546);
xnor U2803 (N_2803,In_2189,In_2065);
or U2804 (N_2804,In_1978,In_1653);
xnor U2805 (N_2805,In_1077,In_201);
nor U2806 (N_2806,In_1077,In_1434);
nand U2807 (N_2807,In_31,In_1999);
nor U2808 (N_2808,In_2214,In_1923);
or U2809 (N_2809,In_1025,In_1345);
nand U2810 (N_2810,In_1831,In_904);
nor U2811 (N_2811,In_1812,In_2195);
nor U2812 (N_2812,In_1178,In_1627);
or U2813 (N_2813,In_1767,In_1004);
xor U2814 (N_2814,In_641,In_2402);
and U2815 (N_2815,In_2397,In_164);
and U2816 (N_2816,In_155,In_2499);
nor U2817 (N_2817,In_987,In_2194);
nor U2818 (N_2818,In_514,In_483);
nor U2819 (N_2819,In_839,In_2419);
and U2820 (N_2820,In_1370,In_585);
and U2821 (N_2821,In_1951,In_1183);
nand U2822 (N_2822,In_277,In_1649);
nor U2823 (N_2823,In_1312,In_1057);
or U2824 (N_2824,In_400,In_1243);
and U2825 (N_2825,In_925,In_2224);
or U2826 (N_2826,In_1409,In_2214);
nand U2827 (N_2827,In_600,In_1379);
nand U2828 (N_2828,In_1163,In_2188);
or U2829 (N_2829,In_1959,In_2181);
nand U2830 (N_2830,In_1680,In_532);
xnor U2831 (N_2831,In_1323,In_1083);
nor U2832 (N_2832,In_2151,In_438);
nand U2833 (N_2833,In_975,In_1073);
or U2834 (N_2834,In_1890,In_1680);
nand U2835 (N_2835,In_961,In_1305);
nor U2836 (N_2836,In_1604,In_321);
or U2837 (N_2837,In_2482,In_458);
nand U2838 (N_2838,In_23,In_246);
or U2839 (N_2839,In_311,In_111);
nand U2840 (N_2840,In_1198,In_2474);
and U2841 (N_2841,In_68,In_138);
nand U2842 (N_2842,In_949,In_1201);
nor U2843 (N_2843,In_2432,In_1779);
nand U2844 (N_2844,In_3,In_2279);
nand U2845 (N_2845,In_1939,In_1029);
and U2846 (N_2846,In_2252,In_29);
nand U2847 (N_2847,In_1359,In_2114);
nor U2848 (N_2848,In_717,In_2187);
nand U2849 (N_2849,In_379,In_236);
nand U2850 (N_2850,In_2387,In_463);
xnor U2851 (N_2851,In_499,In_21);
or U2852 (N_2852,In_2124,In_1434);
nand U2853 (N_2853,In_1545,In_2117);
nand U2854 (N_2854,In_997,In_833);
nor U2855 (N_2855,In_111,In_1069);
or U2856 (N_2856,In_992,In_649);
and U2857 (N_2857,In_2308,In_735);
nor U2858 (N_2858,In_72,In_846);
nand U2859 (N_2859,In_297,In_789);
or U2860 (N_2860,In_40,In_818);
nor U2861 (N_2861,In_2098,In_1664);
or U2862 (N_2862,In_164,In_409);
xor U2863 (N_2863,In_1698,In_1369);
or U2864 (N_2864,In_411,In_2426);
nand U2865 (N_2865,In_2334,In_237);
nor U2866 (N_2866,In_412,In_2080);
nor U2867 (N_2867,In_2155,In_149);
nor U2868 (N_2868,In_1639,In_2013);
nor U2869 (N_2869,In_606,In_803);
or U2870 (N_2870,In_1371,In_1147);
nand U2871 (N_2871,In_1861,In_533);
nand U2872 (N_2872,In_1863,In_1003);
nor U2873 (N_2873,In_1835,In_1336);
and U2874 (N_2874,In_133,In_680);
xnor U2875 (N_2875,In_496,In_1024);
nor U2876 (N_2876,In_1965,In_113);
nand U2877 (N_2877,In_327,In_700);
nand U2878 (N_2878,In_120,In_1647);
nand U2879 (N_2879,In_2012,In_1334);
or U2880 (N_2880,In_2298,In_2461);
or U2881 (N_2881,In_2385,In_1245);
and U2882 (N_2882,In_1479,In_506);
nor U2883 (N_2883,In_1798,In_898);
xnor U2884 (N_2884,In_189,In_2455);
xor U2885 (N_2885,In_2322,In_2342);
nand U2886 (N_2886,In_2334,In_1249);
and U2887 (N_2887,In_2116,In_2470);
or U2888 (N_2888,In_1821,In_1951);
and U2889 (N_2889,In_89,In_1242);
and U2890 (N_2890,In_1223,In_1632);
nand U2891 (N_2891,In_1572,In_1058);
nand U2892 (N_2892,In_1679,In_816);
or U2893 (N_2893,In_1339,In_2250);
nand U2894 (N_2894,In_2282,In_389);
or U2895 (N_2895,In_1344,In_1491);
nor U2896 (N_2896,In_212,In_958);
nand U2897 (N_2897,In_651,In_2295);
or U2898 (N_2898,In_1604,In_1179);
nor U2899 (N_2899,In_976,In_1898);
nor U2900 (N_2900,In_1522,In_2281);
and U2901 (N_2901,In_309,In_2141);
and U2902 (N_2902,In_1624,In_1626);
and U2903 (N_2903,In_649,In_725);
and U2904 (N_2904,In_1751,In_2391);
or U2905 (N_2905,In_869,In_1772);
and U2906 (N_2906,In_1828,In_1320);
nand U2907 (N_2907,In_2369,In_1447);
nand U2908 (N_2908,In_1728,In_1890);
and U2909 (N_2909,In_266,In_549);
or U2910 (N_2910,In_2438,In_2046);
nor U2911 (N_2911,In_707,In_1090);
nor U2912 (N_2912,In_1346,In_1412);
nand U2913 (N_2913,In_2498,In_157);
nor U2914 (N_2914,In_1899,In_906);
nor U2915 (N_2915,In_1268,In_1146);
nor U2916 (N_2916,In_1139,In_2024);
nor U2917 (N_2917,In_768,In_1835);
nand U2918 (N_2918,In_1881,In_1513);
nand U2919 (N_2919,In_6,In_2220);
nor U2920 (N_2920,In_239,In_33);
or U2921 (N_2921,In_302,In_278);
nand U2922 (N_2922,In_649,In_328);
nor U2923 (N_2923,In_1801,In_2204);
and U2924 (N_2924,In_1943,In_280);
xnor U2925 (N_2925,In_1201,In_340);
xnor U2926 (N_2926,In_1780,In_2468);
nand U2927 (N_2927,In_1042,In_2370);
or U2928 (N_2928,In_1772,In_1595);
nand U2929 (N_2929,In_2043,In_1805);
xnor U2930 (N_2930,In_959,In_2381);
nand U2931 (N_2931,In_652,In_2236);
nor U2932 (N_2932,In_1551,In_1485);
or U2933 (N_2933,In_2476,In_1610);
nor U2934 (N_2934,In_227,In_797);
or U2935 (N_2935,In_1922,In_1375);
xnor U2936 (N_2936,In_2472,In_1527);
xor U2937 (N_2937,In_899,In_72);
nand U2938 (N_2938,In_1527,In_605);
or U2939 (N_2939,In_1505,In_277);
or U2940 (N_2940,In_1008,In_1780);
and U2941 (N_2941,In_1698,In_1943);
and U2942 (N_2942,In_674,In_1128);
and U2943 (N_2943,In_216,In_154);
or U2944 (N_2944,In_1294,In_2436);
nor U2945 (N_2945,In_808,In_329);
nor U2946 (N_2946,In_1546,In_875);
nor U2947 (N_2947,In_418,In_1124);
xor U2948 (N_2948,In_2355,In_1493);
and U2949 (N_2949,In_1865,In_1622);
xnor U2950 (N_2950,In_756,In_1025);
and U2951 (N_2951,In_1233,In_1843);
xnor U2952 (N_2952,In_2369,In_709);
and U2953 (N_2953,In_945,In_1741);
xor U2954 (N_2954,In_1598,In_647);
nand U2955 (N_2955,In_606,In_1175);
and U2956 (N_2956,In_2088,In_1008);
nand U2957 (N_2957,In_1084,In_2166);
and U2958 (N_2958,In_2402,In_2248);
nand U2959 (N_2959,In_1236,In_249);
and U2960 (N_2960,In_1857,In_2170);
nor U2961 (N_2961,In_1042,In_2010);
nor U2962 (N_2962,In_2266,In_531);
nand U2963 (N_2963,In_1278,In_2451);
or U2964 (N_2964,In_657,In_798);
or U2965 (N_2965,In_1688,In_2332);
or U2966 (N_2966,In_752,In_884);
or U2967 (N_2967,In_1206,In_145);
xor U2968 (N_2968,In_548,In_2255);
and U2969 (N_2969,In_182,In_199);
nand U2970 (N_2970,In_197,In_987);
nor U2971 (N_2971,In_267,In_731);
nor U2972 (N_2972,In_1522,In_1034);
or U2973 (N_2973,In_767,In_754);
and U2974 (N_2974,In_53,In_665);
nor U2975 (N_2975,In_2313,In_2052);
nor U2976 (N_2976,In_915,In_773);
nand U2977 (N_2977,In_305,In_65);
and U2978 (N_2978,In_355,In_2204);
or U2979 (N_2979,In_463,In_529);
nor U2980 (N_2980,In_242,In_1564);
nor U2981 (N_2981,In_5,In_889);
or U2982 (N_2982,In_189,In_1519);
xnor U2983 (N_2983,In_117,In_2178);
or U2984 (N_2984,In_1900,In_971);
nand U2985 (N_2985,In_830,In_1132);
or U2986 (N_2986,In_473,In_2273);
nor U2987 (N_2987,In_740,In_1206);
and U2988 (N_2988,In_488,In_986);
nor U2989 (N_2989,In_195,In_1227);
and U2990 (N_2990,In_263,In_73);
xor U2991 (N_2991,In_2472,In_2402);
xor U2992 (N_2992,In_2449,In_2366);
nor U2993 (N_2993,In_693,In_1232);
nand U2994 (N_2994,In_1571,In_290);
and U2995 (N_2995,In_2117,In_1098);
nor U2996 (N_2996,In_2108,In_634);
nand U2997 (N_2997,In_904,In_2370);
and U2998 (N_2998,In_1846,In_634);
or U2999 (N_2999,In_1351,In_1372);
nor U3000 (N_3000,In_1880,In_420);
nor U3001 (N_3001,In_719,In_509);
nand U3002 (N_3002,In_1691,In_2165);
nor U3003 (N_3003,In_1857,In_1739);
xnor U3004 (N_3004,In_2301,In_420);
or U3005 (N_3005,In_1676,In_675);
or U3006 (N_3006,In_1358,In_2224);
nor U3007 (N_3007,In_98,In_1939);
and U3008 (N_3008,In_2181,In_2036);
nand U3009 (N_3009,In_2412,In_950);
nand U3010 (N_3010,In_1412,In_1432);
nand U3011 (N_3011,In_1674,In_650);
nand U3012 (N_3012,In_1434,In_2214);
and U3013 (N_3013,In_2188,In_104);
and U3014 (N_3014,In_273,In_1070);
nand U3015 (N_3015,In_651,In_1149);
xor U3016 (N_3016,In_809,In_579);
or U3017 (N_3017,In_832,In_605);
xnor U3018 (N_3018,In_1259,In_834);
nor U3019 (N_3019,In_1447,In_2424);
nor U3020 (N_3020,In_143,In_2063);
and U3021 (N_3021,In_1543,In_914);
xor U3022 (N_3022,In_1389,In_122);
nor U3023 (N_3023,In_2384,In_1512);
and U3024 (N_3024,In_2231,In_1240);
nor U3025 (N_3025,In_763,In_1930);
nor U3026 (N_3026,In_2336,In_2260);
xnor U3027 (N_3027,In_1413,In_765);
or U3028 (N_3028,In_2094,In_1244);
or U3029 (N_3029,In_2010,In_1901);
nor U3030 (N_3030,In_1750,In_2388);
and U3031 (N_3031,In_218,In_365);
nor U3032 (N_3032,In_2163,In_319);
nor U3033 (N_3033,In_2183,In_1458);
xor U3034 (N_3034,In_1017,In_1372);
nand U3035 (N_3035,In_700,In_2040);
nor U3036 (N_3036,In_236,In_1421);
or U3037 (N_3037,In_1984,In_1091);
and U3038 (N_3038,In_1724,In_2221);
xor U3039 (N_3039,In_1649,In_1696);
nor U3040 (N_3040,In_59,In_664);
or U3041 (N_3041,In_708,In_229);
nor U3042 (N_3042,In_2204,In_1052);
or U3043 (N_3043,In_639,In_829);
nor U3044 (N_3044,In_603,In_978);
and U3045 (N_3045,In_139,In_1672);
xnor U3046 (N_3046,In_1799,In_2419);
xor U3047 (N_3047,In_2396,In_1321);
or U3048 (N_3048,In_436,In_1389);
xor U3049 (N_3049,In_1278,In_980);
and U3050 (N_3050,In_589,In_851);
and U3051 (N_3051,In_157,In_2126);
and U3052 (N_3052,In_2232,In_69);
nor U3053 (N_3053,In_440,In_1922);
nor U3054 (N_3054,In_1177,In_1718);
and U3055 (N_3055,In_593,In_621);
and U3056 (N_3056,In_2101,In_406);
nor U3057 (N_3057,In_1217,In_1480);
and U3058 (N_3058,In_1743,In_453);
and U3059 (N_3059,In_1356,In_418);
and U3060 (N_3060,In_1346,In_1755);
nand U3061 (N_3061,In_1943,In_1814);
or U3062 (N_3062,In_171,In_1148);
and U3063 (N_3063,In_2186,In_412);
and U3064 (N_3064,In_28,In_2105);
xor U3065 (N_3065,In_655,In_419);
xnor U3066 (N_3066,In_2106,In_333);
nor U3067 (N_3067,In_955,In_970);
nor U3068 (N_3068,In_206,In_1415);
nand U3069 (N_3069,In_1889,In_1981);
and U3070 (N_3070,In_1541,In_1774);
and U3071 (N_3071,In_2333,In_2287);
and U3072 (N_3072,In_470,In_626);
nand U3073 (N_3073,In_2073,In_2053);
or U3074 (N_3074,In_1832,In_1873);
xnor U3075 (N_3075,In_2142,In_179);
or U3076 (N_3076,In_2458,In_1407);
nand U3077 (N_3077,In_575,In_979);
nor U3078 (N_3078,In_1366,In_1277);
or U3079 (N_3079,In_2060,In_1066);
and U3080 (N_3080,In_388,In_1085);
nand U3081 (N_3081,In_467,In_524);
xor U3082 (N_3082,In_261,In_2340);
xnor U3083 (N_3083,In_977,In_1222);
nor U3084 (N_3084,In_1190,In_2134);
nor U3085 (N_3085,In_282,In_826);
nor U3086 (N_3086,In_1829,In_1784);
nand U3087 (N_3087,In_2413,In_696);
nor U3088 (N_3088,In_497,In_2192);
nor U3089 (N_3089,In_1361,In_698);
or U3090 (N_3090,In_865,In_116);
and U3091 (N_3091,In_2087,In_2017);
or U3092 (N_3092,In_1728,In_1032);
nand U3093 (N_3093,In_1718,In_2333);
nor U3094 (N_3094,In_2313,In_605);
or U3095 (N_3095,In_2258,In_2289);
and U3096 (N_3096,In_153,In_1373);
nand U3097 (N_3097,In_1337,In_303);
and U3098 (N_3098,In_819,In_867);
nand U3099 (N_3099,In_962,In_540);
nand U3100 (N_3100,In_579,In_71);
or U3101 (N_3101,In_1288,In_1582);
nand U3102 (N_3102,In_885,In_1799);
nor U3103 (N_3103,In_1558,In_1770);
nor U3104 (N_3104,In_1988,In_488);
nand U3105 (N_3105,In_2059,In_2074);
or U3106 (N_3106,In_738,In_779);
nand U3107 (N_3107,In_2247,In_395);
xor U3108 (N_3108,In_2120,In_483);
and U3109 (N_3109,In_314,In_587);
xnor U3110 (N_3110,In_976,In_734);
or U3111 (N_3111,In_1550,In_1589);
or U3112 (N_3112,In_1350,In_153);
nand U3113 (N_3113,In_1906,In_516);
nand U3114 (N_3114,In_1072,In_868);
and U3115 (N_3115,In_762,In_1166);
and U3116 (N_3116,In_450,In_1636);
nand U3117 (N_3117,In_1727,In_584);
and U3118 (N_3118,In_300,In_1537);
or U3119 (N_3119,In_202,In_393);
nand U3120 (N_3120,In_844,In_1431);
xor U3121 (N_3121,In_834,In_1889);
nand U3122 (N_3122,In_1839,In_569);
xor U3123 (N_3123,In_1726,In_2);
and U3124 (N_3124,In_1083,In_550);
and U3125 (N_3125,N_2886,N_240);
nand U3126 (N_3126,N_553,N_2947);
nand U3127 (N_3127,N_1850,N_1202);
xor U3128 (N_3128,N_1725,N_1740);
or U3129 (N_3129,N_1532,N_2759);
nand U3130 (N_3130,N_1751,N_1133);
nand U3131 (N_3131,N_2426,N_221);
nor U3132 (N_3132,N_1134,N_206);
or U3133 (N_3133,N_959,N_2789);
or U3134 (N_3134,N_2549,N_1713);
nor U3135 (N_3135,N_474,N_1887);
and U3136 (N_3136,N_3103,N_2192);
nand U3137 (N_3137,N_2744,N_2904);
nand U3138 (N_3138,N_171,N_2634);
xor U3139 (N_3139,N_2331,N_851);
xnor U3140 (N_3140,N_2043,N_1561);
nand U3141 (N_3141,N_1185,N_971);
and U3142 (N_3142,N_2275,N_1307);
or U3143 (N_3143,N_755,N_2738);
and U3144 (N_3144,N_305,N_2638);
or U3145 (N_3145,N_1959,N_312);
nand U3146 (N_3146,N_1719,N_3044);
or U3147 (N_3147,N_583,N_1374);
nor U3148 (N_3148,N_1580,N_30);
and U3149 (N_3149,N_3102,N_2942);
nor U3150 (N_3150,N_1557,N_2501);
and U3151 (N_3151,N_1602,N_1593);
nand U3152 (N_3152,N_820,N_2939);
nor U3153 (N_3153,N_1196,N_2060);
or U3154 (N_3154,N_1223,N_945);
nand U3155 (N_3155,N_192,N_2380);
and U3156 (N_3156,N_1705,N_2495);
and U3157 (N_3157,N_329,N_208);
nor U3158 (N_3158,N_2677,N_2040);
nor U3159 (N_3159,N_1412,N_1228);
and U3160 (N_3160,N_1062,N_2628);
nor U3161 (N_3161,N_379,N_390);
nor U3162 (N_3162,N_1966,N_20);
nor U3163 (N_3163,N_951,N_2340);
and U3164 (N_3164,N_1184,N_2674);
and U3165 (N_3165,N_3005,N_1110);
xor U3166 (N_3166,N_1220,N_3008);
nor U3167 (N_3167,N_380,N_2989);
and U3168 (N_3168,N_1188,N_1954);
nand U3169 (N_3169,N_2037,N_2257);
or U3170 (N_3170,N_67,N_2277);
nand U3171 (N_3171,N_1927,N_1317);
nand U3172 (N_3172,N_1801,N_2418);
or U3173 (N_3173,N_1132,N_1404);
and U3174 (N_3174,N_2899,N_2400);
nor U3175 (N_3175,N_447,N_317);
nand U3176 (N_3176,N_1926,N_2028);
and U3177 (N_3177,N_1457,N_487);
or U3178 (N_3178,N_607,N_2562);
nand U3179 (N_3179,N_2826,N_2035);
and U3180 (N_3180,N_2747,N_2099);
or U3181 (N_3181,N_2221,N_1799);
and U3182 (N_3182,N_1794,N_1967);
xnor U3183 (N_3183,N_187,N_485);
nor U3184 (N_3184,N_2681,N_2154);
nand U3185 (N_3185,N_1230,N_738);
nand U3186 (N_3186,N_2498,N_729);
xnor U3187 (N_3187,N_678,N_1351);
or U3188 (N_3188,N_158,N_1283);
and U3189 (N_3189,N_1796,N_630);
nand U3190 (N_3190,N_1314,N_2843);
and U3191 (N_3191,N_327,N_1089);
nand U3192 (N_3192,N_2551,N_499);
xor U3193 (N_3193,N_2298,N_692);
nand U3194 (N_3194,N_494,N_11);
nand U3195 (N_3195,N_2,N_842);
or U3196 (N_3196,N_773,N_2053);
nand U3197 (N_3197,N_792,N_1902);
xnor U3198 (N_3198,N_3114,N_1426);
nor U3199 (N_3199,N_1911,N_59);
xnor U3200 (N_3200,N_782,N_589);
nand U3201 (N_3201,N_744,N_3006);
and U3202 (N_3202,N_2961,N_525);
nor U3203 (N_3203,N_2813,N_1509);
nand U3204 (N_3204,N_776,N_1588);
and U3205 (N_3205,N_283,N_130);
xor U3206 (N_3206,N_2309,N_817);
or U3207 (N_3207,N_1310,N_2379);
or U3208 (N_3208,N_1732,N_845);
nand U3209 (N_3209,N_2537,N_1256);
nand U3210 (N_3210,N_1393,N_688);
and U3211 (N_3211,N_2541,N_465);
and U3212 (N_3212,N_941,N_2656);
nand U3213 (N_3213,N_716,N_89);
xor U3214 (N_3214,N_2065,N_1689);
and U3215 (N_3215,N_2610,N_2974);
nand U3216 (N_3216,N_1095,N_2991);
nor U3217 (N_3217,N_2440,N_804);
and U3218 (N_3218,N_1271,N_2249);
and U3219 (N_3219,N_1748,N_2621);
nor U3220 (N_3220,N_2609,N_1253);
or U3221 (N_3221,N_1913,N_878);
nor U3222 (N_3222,N_2078,N_2251);
and U3223 (N_3223,N_707,N_1644);
nor U3224 (N_3224,N_1222,N_2336);
and U3225 (N_3225,N_1045,N_1829);
nand U3226 (N_3226,N_2546,N_2887);
or U3227 (N_3227,N_602,N_1108);
nand U3228 (N_3228,N_80,N_1570);
and U3229 (N_3229,N_1147,N_51);
and U3230 (N_3230,N_3077,N_2150);
nand U3231 (N_3231,N_2468,N_40);
and U3232 (N_3232,N_1478,N_970);
or U3233 (N_3233,N_2783,N_2911);
nand U3234 (N_3234,N_2346,N_1493);
and U3235 (N_3235,N_1445,N_1894);
or U3236 (N_3236,N_475,N_1325);
or U3237 (N_3237,N_183,N_469);
and U3238 (N_3238,N_2750,N_1016);
nor U3239 (N_3239,N_1073,N_1336);
and U3240 (N_3240,N_2864,N_1984);
nor U3241 (N_3241,N_423,N_2914);
and U3242 (N_3242,N_2545,N_230);
nor U3243 (N_3243,N_1687,N_3096);
nor U3244 (N_3244,N_1119,N_1060);
and U3245 (N_3245,N_1760,N_1503);
nor U3246 (N_3246,N_1684,N_558);
nor U3247 (N_3247,N_129,N_1093);
or U3248 (N_3248,N_3118,N_1573);
and U3249 (N_3249,N_2419,N_2829);
or U3250 (N_3250,N_1679,N_2872);
or U3251 (N_3251,N_2922,N_1581);
or U3252 (N_3252,N_2413,N_814);
xor U3253 (N_3253,N_2281,N_1653);
and U3254 (N_3254,N_3040,N_2892);
nor U3255 (N_3255,N_1254,N_404);
nor U3256 (N_3256,N_426,N_1433);
and U3257 (N_3257,N_1474,N_1327);
nand U3258 (N_3258,N_764,N_1510);
nor U3259 (N_3259,N_2633,N_2590);
xor U3260 (N_3260,N_1168,N_1259);
xor U3261 (N_3261,N_1475,N_2850);
and U3262 (N_3262,N_1237,N_2692);
and U3263 (N_3263,N_2987,N_1257);
or U3264 (N_3264,N_2721,N_2349);
or U3265 (N_3265,N_1768,N_689);
and U3266 (N_3266,N_219,N_2175);
nor U3267 (N_3267,N_1008,N_174);
and U3268 (N_3268,N_2095,N_900);
and U3269 (N_3269,N_933,N_2569);
or U3270 (N_3270,N_1920,N_2220);
nand U3271 (N_3271,N_2619,N_121);
nor U3272 (N_3272,N_139,N_1523);
nor U3273 (N_3273,N_2671,N_1007);
or U3274 (N_3274,N_1945,N_579);
or U3275 (N_3275,N_2529,N_982);
nand U3276 (N_3276,N_55,N_1847);
xnor U3277 (N_3277,N_1671,N_1377);
nand U3278 (N_3278,N_676,N_1448);
nor U3279 (N_3279,N_1214,N_1813);
and U3280 (N_3280,N_1654,N_977);
nand U3281 (N_3281,N_497,N_1741);
or U3282 (N_3282,N_166,N_3123);
nor U3283 (N_3283,N_747,N_1960);
nor U3284 (N_3284,N_2881,N_615);
nor U3285 (N_3285,N_1178,N_271);
nor U3286 (N_3286,N_813,N_176);
and U3287 (N_3287,N_2780,N_756);
xor U3288 (N_3288,N_983,N_636);
and U3289 (N_3289,N_2019,N_1406);
nor U3290 (N_3290,N_619,N_3056);
and U3291 (N_3291,N_2423,N_521);
nor U3292 (N_3292,N_1494,N_2174);
or U3293 (N_3293,N_2951,N_212);
or U3294 (N_3294,N_1919,N_1239);
nor U3295 (N_3295,N_1519,N_155);
or U3296 (N_3296,N_2354,N_2845);
xor U3297 (N_3297,N_848,N_2201);
or U3298 (N_3298,N_838,N_2494);
nor U3299 (N_3299,N_1826,N_507);
or U3300 (N_3300,N_1549,N_2123);
nor U3301 (N_3301,N_2810,N_2580);
nand U3302 (N_3302,N_1604,N_2685);
xnor U3303 (N_3303,N_2982,N_1331);
nand U3304 (N_3304,N_397,N_260);
nand U3305 (N_3305,N_3117,N_815);
nor U3306 (N_3306,N_2478,N_548);
nor U3307 (N_3307,N_1366,N_1203);
or U3308 (N_3308,N_1368,N_1765);
and U3309 (N_3309,N_458,N_569);
or U3310 (N_3310,N_500,N_1333);
and U3311 (N_3311,N_1096,N_2070);
nand U3312 (N_3312,N_82,N_1703);
and U3313 (N_3313,N_1611,N_277);
and U3314 (N_3314,N_837,N_2970);
nand U3315 (N_3315,N_2771,N_2477);
nor U3316 (N_3316,N_1047,N_291);
or U3317 (N_3317,N_3003,N_87);
or U3318 (N_3318,N_556,N_479);
and U3319 (N_3319,N_1461,N_440);
or U3320 (N_3320,N_114,N_2582);
or U3321 (N_3321,N_879,N_3020);
or U3322 (N_3322,N_1849,N_2552);
or U3323 (N_3323,N_378,N_1638);
nand U3324 (N_3324,N_1169,N_2009);
or U3325 (N_3325,N_1153,N_1018);
xnor U3326 (N_3326,N_143,N_1209);
nor U3327 (N_3327,N_2191,N_2823);
nor U3328 (N_3328,N_177,N_989);
nor U3329 (N_3329,N_38,N_2842);
or U3330 (N_3330,N_1560,N_2695);
or U3331 (N_3331,N_1738,N_109);
or U3332 (N_3332,N_1288,N_2639);
nand U3333 (N_3333,N_517,N_2289);
or U3334 (N_3334,N_2021,N_2000);
xnor U3335 (N_3335,N_1628,N_561);
nor U3336 (N_3336,N_2458,N_3032);
nor U3337 (N_3337,N_2058,N_1213);
nor U3338 (N_3338,N_3112,N_101);
or U3339 (N_3339,N_2788,N_1903);
nor U3340 (N_3340,N_2885,N_2714);
or U3341 (N_3341,N_2001,N_601);
nand U3342 (N_3342,N_659,N_153);
and U3343 (N_3343,N_2466,N_2958);
nand U3344 (N_3344,N_3079,N_1914);
nand U3345 (N_3345,N_2386,N_1662);
or U3346 (N_3346,N_760,N_849);
nor U3347 (N_3347,N_1236,N_1845);
nand U3348 (N_3348,N_2948,N_2840);
nor U3349 (N_3349,N_2875,N_1250);
nor U3350 (N_3350,N_102,N_3013);
or U3351 (N_3351,N_2111,N_918);
or U3352 (N_3352,N_1437,N_2793);
nand U3353 (N_3353,N_1099,N_2055);
nor U3354 (N_3354,N_2712,N_3015);
or U3355 (N_3355,N_314,N_1001);
nor U3356 (N_3356,N_1859,N_944);
nor U3357 (N_3357,N_1962,N_1619);
nor U3358 (N_3358,N_2110,N_339);
or U3359 (N_3359,N_681,N_626);
and U3360 (N_3360,N_1935,N_10);
nor U3361 (N_3361,N_2026,N_753);
or U3362 (N_3362,N_713,N_2225);
and U3363 (N_3363,N_962,N_213);
nor U3364 (N_3364,N_793,N_1241);
xor U3365 (N_3365,N_122,N_1780);
or U3366 (N_3366,N_958,N_1907);
nor U3367 (N_3367,N_1082,N_743);
nor U3368 (N_3368,N_34,N_686);
and U3369 (N_3369,N_2320,N_2637);
nor U3370 (N_3370,N_1371,N_598);
nand U3371 (N_3371,N_1527,N_2965);
nor U3372 (N_3372,N_2461,N_2996);
nor U3373 (N_3373,N_2623,N_1197);
or U3374 (N_3374,N_2764,N_797);
nand U3375 (N_3375,N_286,N_2563);
and U3376 (N_3376,N_980,N_394);
nand U3377 (N_3377,N_2817,N_133);
nand U3378 (N_3378,N_3099,N_229);
and U3379 (N_3379,N_606,N_1301);
or U3380 (N_3380,N_1171,N_2596);
or U3381 (N_3381,N_2069,N_924);
and U3382 (N_3382,N_1886,N_1425);
nor U3383 (N_3383,N_2560,N_1453);
or U3384 (N_3384,N_825,N_1925);
nand U3385 (N_3385,N_1126,N_2263);
nor U3386 (N_3386,N_146,N_2283);
or U3387 (N_3387,N_795,N_2411);
and U3388 (N_3388,N_255,N_974);
or U3389 (N_3389,N_516,N_46);
and U3390 (N_3390,N_2235,N_292);
and U3391 (N_3391,N_2530,N_1234);
and U3392 (N_3392,N_2555,N_893);
nand U3393 (N_3393,N_1391,N_1548);
nor U3394 (N_3394,N_224,N_2393);
or U3395 (N_3395,N_2469,N_700);
nand U3396 (N_3396,N_169,N_735);
or U3397 (N_3397,N_1430,N_310);
or U3398 (N_3398,N_2740,N_2168);
or U3399 (N_3399,N_1338,N_1358);
nand U3400 (N_3400,N_1490,N_103);
nand U3401 (N_3401,N_1405,N_1212);
nand U3402 (N_3402,N_1779,N_1979);
and U3403 (N_3403,N_1855,N_2134);
and U3404 (N_3404,N_720,N_1320);
nor U3405 (N_3405,N_1727,N_459);
and U3406 (N_3406,N_547,N_969);
and U3407 (N_3407,N_3016,N_1943);
and U3408 (N_3408,N_2465,N_1415);
nand U3409 (N_3409,N_2969,N_1612);
or U3410 (N_3410,N_2353,N_2601);
nor U3411 (N_3411,N_1791,N_642);
or U3412 (N_3412,N_1516,N_27);
or U3413 (N_3413,N_1322,N_3035);
nor U3414 (N_3414,N_2972,N_2149);
or U3415 (N_3415,N_1873,N_318);
xor U3416 (N_3416,N_2179,N_2757);
and U3417 (N_3417,N_667,N_766);
and U3418 (N_3418,N_835,N_301);
nor U3419 (N_3419,N_1881,N_2526);
nor U3420 (N_3420,N_58,N_2932);
nor U3421 (N_3421,N_182,N_2857);
and U3422 (N_3422,N_53,N_2247);
nand U3423 (N_3423,N_1485,N_1578);
or U3424 (N_3424,N_2640,N_1879);
nor U3425 (N_3425,N_1315,N_2373);
nor U3426 (N_3426,N_1563,N_2189);
and U3427 (N_3427,N_1266,N_2462);
nor U3428 (N_3428,N_2278,N_1931);
and U3429 (N_3429,N_1942,N_786);
or U3430 (N_3430,N_1141,N_2586);
nor U3431 (N_3431,N_2851,N_2934);
nor U3432 (N_3432,N_603,N_2625);
xor U3433 (N_3433,N_2085,N_2135);
or U3434 (N_3434,N_2983,N_610);
and U3435 (N_3435,N_644,N_2509);
xor U3436 (N_3436,N_2572,N_2330);
nor U3437 (N_3437,N_1111,N_3078);
nand U3438 (N_3438,N_1399,N_178);
nor U3439 (N_3439,N_1674,N_2715);
xnor U3440 (N_3440,N_2884,N_2790);
nand U3441 (N_3441,N_1835,N_1896);
nor U3442 (N_3442,N_874,N_629);
nor U3443 (N_3443,N_2205,N_2758);
or U3444 (N_3444,N_2701,N_737);
nor U3445 (N_3445,N_2532,N_1888);
nor U3446 (N_3446,N_2635,N_2363);
and U3447 (N_3447,N_931,N_1422);
xnor U3448 (N_3448,N_1709,N_2253);
and U3449 (N_3449,N_645,N_2518);
and U3450 (N_3450,N_2956,N_333);
nand U3451 (N_3451,N_2279,N_822);
or U3452 (N_3452,N_967,N_2612);
nand U3453 (N_3453,N_880,N_2866);
and U3454 (N_3454,N_1970,N_1897);
nor U3455 (N_3455,N_1981,N_1973);
or U3456 (N_3456,N_1118,N_867);
nand U3457 (N_3457,N_1484,N_715);
nor U3458 (N_3458,N_1989,N_1782);
and U3459 (N_3459,N_762,N_2038);
or U3460 (N_3460,N_975,N_2870);
xor U3461 (N_3461,N_3104,N_624);
or U3462 (N_3462,N_1949,N_1194);
nand U3463 (N_3463,N_3041,N_1528);
and U3464 (N_3464,N_2211,N_2897);
nor U3465 (N_3465,N_204,N_1483);
nor U3466 (N_3466,N_1758,N_2763);
and U3467 (N_3467,N_2809,N_396);
and U3468 (N_3468,N_1695,N_2093);
nand U3469 (N_3469,N_655,N_1225);
xor U3470 (N_3470,N_1539,N_1058);
nor U3471 (N_3471,N_1722,N_1825);
nor U3472 (N_3472,N_2825,N_2256);
nand U3473 (N_3473,N_1379,N_2500);
or U3474 (N_3474,N_2753,N_966);
and U3475 (N_3475,N_2091,N_2720);
and U3476 (N_3476,N_268,N_308);
and U3477 (N_3477,N_2136,N_2867);
xnor U3478 (N_3478,N_670,N_635);
and U3479 (N_3479,N_1800,N_2709);
and U3480 (N_3480,N_936,N_1023);
nand U3481 (N_3481,N_2482,N_549);
nand U3482 (N_3482,N_1034,N_1071);
nor U3483 (N_3483,N_1027,N_2997);
nand U3484 (N_3484,N_2248,N_2234);
or U3485 (N_3485,N_1786,N_1244);
and U3486 (N_3486,N_2933,N_2307);
nand U3487 (N_3487,N_2077,N_2265);
nor U3488 (N_3488,N_2903,N_462);
nor U3489 (N_3489,N_1515,N_1750);
nor U3490 (N_3490,N_2362,N_1854);
nor U3491 (N_3491,N_690,N_2818);
or U3492 (N_3492,N_572,N_1159);
nor U3493 (N_3493,N_1339,N_2909);
and U3494 (N_3494,N_413,N_251);
or U3495 (N_3495,N_905,N_1451);
xnor U3496 (N_3496,N_2074,N_2003);
nand U3497 (N_3497,N_1831,N_403);
and U3498 (N_3498,N_161,N_2686);
or U3499 (N_3499,N_436,N_641);
and U3500 (N_3500,N_2290,N_662);
nor U3501 (N_3501,N_1871,N_1694);
and U3502 (N_3502,N_2344,N_2873);
and U3503 (N_3503,N_1972,N_1592);
and U3504 (N_3504,N_2990,N_1918);
and U3505 (N_3505,N_1033,N_226);
nand U3506 (N_3506,N_1639,N_1436);
nand U3507 (N_3507,N_2962,N_1499);
nor U3508 (N_3508,N_2244,N_1890);
nand U3509 (N_3509,N_2274,N_576);
or U3510 (N_3510,N_1075,N_803);
and U3511 (N_3511,N_3,N_91);
nand U3512 (N_3512,N_488,N_564);
or U3513 (N_3513,N_2960,N_2350);
nand U3514 (N_3514,N_928,N_1964);
nand U3515 (N_3515,N_1407,N_348);
and U3516 (N_3516,N_1462,N_1867);
and U3517 (N_3517,N_1844,N_142);
and U3518 (N_3518,N_1810,N_1924);
nor U3519 (N_3519,N_858,N_1620);
and U3520 (N_3520,N_1174,N_2605);
or U3521 (N_3521,N_2194,N_3089);
nor U3522 (N_3522,N_528,N_136);
nor U3523 (N_3523,N_726,N_1382);
nand U3524 (N_3524,N_2056,N_906);
nor U3525 (N_3525,N_2728,N_228);
nand U3526 (N_3526,N_1675,N_62);
nor U3527 (N_3527,N_640,N_1504);
nor U3528 (N_3528,N_1305,N_1252);
and U3529 (N_3529,N_2597,N_537);
nor U3530 (N_3530,N_1384,N_2450);
and U3531 (N_3531,N_3070,N_1677);
or U3532 (N_3532,N_1086,N_1577);
or U3533 (N_3533,N_282,N_1010);
or U3534 (N_3534,N_1392,N_1356);
and U3535 (N_3535,N_368,N_3066);
and U3536 (N_3536,N_1100,N_311);
or U3537 (N_3537,N_1376,N_2779);
xnor U3538 (N_3538,N_2856,N_1063);
nor U3539 (N_3539,N_3082,N_2553);
or U3540 (N_3540,N_425,N_1297);
or U3541 (N_3541,N_1658,N_352);
nand U3542 (N_3542,N_1987,N_1357);
nand U3543 (N_3543,N_2854,N_450);
nand U3544 (N_3544,N_2925,N_783);
nor U3545 (N_3545,N_1992,N_2470);
nor U3546 (N_3546,N_2266,N_202);
or U3547 (N_3547,N_2427,N_861);
nor U3548 (N_3548,N_1908,N_1540);
nand U3549 (N_3549,N_54,N_340);
nand U3550 (N_3550,N_994,N_1828);
and U3551 (N_3551,N_1559,N_1556);
or U3552 (N_3552,N_1637,N_2017);
nand U3553 (N_3553,N_1569,N_2160);
nand U3554 (N_3554,N_2971,N_751);
or U3555 (N_3555,N_1041,N_1417);
nor U3556 (N_3556,N_343,N_398);
nand U3557 (N_3557,N_3101,N_859);
nand U3558 (N_3558,N_2337,N_1534);
nand U3559 (N_3559,N_1884,N_1757);
nor U3560 (N_3560,N_631,N_2632);
and U3561 (N_3561,N_847,N_1610);
nor U3562 (N_3562,N_1953,N_2130);
nor U3563 (N_3563,N_2981,N_1541);
or U3564 (N_3564,N_2141,N_1038);
and U3565 (N_3565,N_660,N_2472);
and U3566 (N_3566,N_273,N_677);
and U3567 (N_3567,N_1771,N_470);
nand U3568 (N_3568,N_2358,N_1889);
and U3569 (N_3569,N_388,N_617);
or U3570 (N_3570,N_2007,N_2658);
or U3571 (N_3571,N_2282,N_322);
xnor U3572 (N_3572,N_2062,N_2827);
or U3573 (N_3573,N_2305,N_1745);
and U3574 (N_3574,N_1797,N_596);
xor U3575 (N_3575,N_1956,N_826);
nor U3576 (N_3576,N_342,N_1416);
and U3577 (N_3577,N_3057,N_2539);
or U3578 (N_3578,N_60,N_2163);
nand U3579 (N_3579,N_2143,N_100);
nand U3580 (N_3580,N_976,N_2806);
xnor U3581 (N_3581,N_1024,N_501);
and U3582 (N_3582,N_2893,N_1988);
and U3583 (N_3583,N_1963,N_1127);
or U3584 (N_3584,N_36,N_1818);
xnor U3585 (N_3585,N_2139,N_854);
or U3586 (N_3586,N_2755,N_1112);
nand U3587 (N_3587,N_2202,N_2908);
or U3588 (N_3588,N_2550,N_2369);
xnor U3589 (N_3589,N_527,N_767);
nor U3590 (N_3590,N_2930,N_287);
xnor U3591 (N_3591,N_1892,N_680);
or U3592 (N_3592,N_986,N_1055);
and U3593 (N_3593,N_392,N_42);
or U3594 (N_3594,N_625,N_1530);
xor U3595 (N_3595,N_2812,N_2447);
or U3596 (N_3596,N_2357,N_1245);
nand U3597 (N_3597,N_1231,N_682);
or U3598 (N_3598,N_2067,N_438);
nand U3599 (N_3599,N_802,N_498);
nand U3600 (N_3600,N_2782,N_2242);
and U3601 (N_3601,N_846,N_5);
xnor U3602 (N_3602,N_1621,N_730);
or U3603 (N_3603,N_303,N_2587);
nand U3604 (N_3604,N_1520,N_1455);
nand U3605 (N_3605,N_2381,N_1558);
or U3606 (N_3606,N_324,N_2729);
and U3607 (N_3607,N_3119,N_2226);
nand U3608 (N_3608,N_1562,N_2272);
nand U3609 (N_3609,N_908,N_2215);
and U3610 (N_3610,N_411,N_1840);
and U3611 (N_3611,N_505,N_2464);
nand U3612 (N_3612,N_930,N_123);
nand U3613 (N_3613,N_2853,N_482);
and U3614 (N_3614,N_2161,N_1078);
nand U3615 (N_3615,N_222,N_745);
or U3616 (N_3616,N_248,N_2158);
xor U3617 (N_3617,N_1498,N_214);
nor U3618 (N_3618,N_1158,N_3122);
nand U3619 (N_3619,N_749,N_56);
or U3620 (N_3620,N_2185,N_722);
xnor U3621 (N_3621,N_2296,N_2928);
nor U3622 (N_3622,N_1770,N_913);
and U3623 (N_3623,N_2371,N_464);
nand U3624 (N_3624,N_2408,N_777);
or U3625 (N_3625,N_1006,N_1090);
or U3626 (N_3626,N_2329,N_2120);
and U3627 (N_3627,N_1864,N_2424);
or U3628 (N_3628,N_1037,N_2314);
and U3629 (N_3629,N_964,N_266);
nor U3630 (N_3630,N_1723,N_833);
or U3631 (N_3631,N_1866,N_496);
or U3632 (N_3632,N_927,N_661);
and U3633 (N_3633,N_1706,N_2072);
or U3634 (N_3634,N_876,N_421);
nor U3635 (N_3635,N_1135,N_2535);
nor U3636 (N_3636,N_2071,N_882);
and U3637 (N_3637,N_2444,N_2006);
nand U3638 (N_3638,N_2577,N_536);
or U3639 (N_3639,N_2445,N_3053);
and U3640 (N_3640,N_778,N_359);
nor U3641 (N_3641,N_3060,N_434);
and U3642 (N_3642,N_1057,N_2585);
xnor U3643 (N_3643,N_3109,N_718);
and U3644 (N_3644,N_2651,N_2848);
nor U3645 (N_3645,N_1650,N_1216);
and U3646 (N_3646,N_993,N_250);
and U3647 (N_3647,N_2403,N_2100);
nand U3648 (N_3648,N_1952,N_1772);
xnor U3649 (N_3649,N_2581,N_4);
and U3650 (N_3650,N_3069,N_2548);
nor U3651 (N_3651,N_1454,N_2334);
nor U3652 (N_3652,N_3093,N_2439);
xor U3653 (N_3653,N_3064,N_113);
and U3654 (N_3654,N_1776,N_2504);
xor U3655 (N_3655,N_2250,N_389);
and U3656 (N_3656,N_2271,N_376);
nand U3657 (N_3657,N_509,N_2317);
nor U3658 (N_3658,N_370,N_2820);
or U3659 (N_3659,N_1468,N_774);
nor U3660 (N_3660,N_1156,N_1488);
or U3661 (N_3661,N_2702,N_2162);
or U3662 (N_3662,N_2097,N_1633);
xor U3663 (N_3663,N_665,N_1365);
or U3664 (N_3664,N_2322,N_2173);
nor U3665 (N_3665,N_1264,N_2300);
xnor U3666 (N_3666,N_2308,N_1292);
nand U3667 (N_3667,N_853,N_1120);
xor U3668 (N_3668,N_1575,N_3111);
nor U3669 (N_3669,N_2547,N_1961);
xnor U3670 (N_3670,N_698,N_2404);
xor U3671 (N_3671,N_1420,N_2531);
and U3672 (N_3672,N_1506,N_1550);
and U3673 (N_3673,N_1400,N_2938);
nand U3674 (N_3674,N_761,N_2855);
and U3675 (N_3675,N_1995,N_150);
and U3676 (N_3676,N_2646,N_1716);
nor U3677 (N_3677,N_775,N_2558);
nor U3678 (N_3678,N_1242,N_1247);
or U3679 (N_3679,N_1277,N_801);
and U3680 (N_3680,N_2044,N_181);
nor U3681 (N_3681,N_2033,N_3048);
and U3682 (N_3682,N_2064,N_1587);
nor U3683 (N_3683,N_2394,N_13);
nand U3684 (N_3684,N_2184,N_1162);
nor U3685 (N_3685,N_1505,N_524);
xnor U3686 (N_3686,N_154,N_1734);
nand U3687 (N_3687,N_1603,N_2324);
nor U3688 (N_3688,N_2802,N_2725);
nand U3689 (N_3689,N_1891,N_1274);
and U3690 (N_3690,N_965,N_1092);
or U3691 (N_3691,N_1893,N_1950);
or U3692 (N_3692,N_2953,N_2406);
or U3693 (N_3693,N_1465,N_2238);
and U3694 (N_3694,N_942,N_2260);
or U3695 (N_3695,N_2387,N_2452);
nand U3696 (N_3696,N_895,N_1744);
nand U3697 (N_3697,N_2066,N_294);
or U3698 (N_3698,N_2116,N_407);
nor U3699 (N_3699,N_2112,N_186);
and U3700 (N_3700,N_1281,N_1172);
nand U3701 (N_3701,N_2285,N_2119);
nand U3702 (N_3702,N_480,N_650);
nor U3703 (N_3703,N_2303,N_990);
nand U3704 (N_3704,N_2900,N_1481);
nand U3705 (N_3705,N_1817,N_2280);
or U3706 (N_3706,N_2708,N_1998);
nand U3707 (N_3707,N_1328,N_2929);
nand U3708 (N_3708,N_1806,N_1900);
xnor U3709 (N_3709,N_3054,N_2841);
nand U3710 (N_3710,N_1767,N_1634);
nand U3711 (N_3711,N_1615,N_2047);
xnor U3712 (N_3712,N_2068,N_2483);
nor U3713 (N_3713,N_950,N_2684);
or U3714 (N_3714,N_911,N_3098);
nand U3715 (N_3715,N_2591,N_1629);
nand U3716 (N_3716,N_3074,N_2181);
nor U3717 (N_3717,N_1039,N_163);
or U3718 (N_3718,N_3067,N_3027);
or U3719 (N_3719,N_1401,N_1370);
and U3720 (N_3720,N_2687,N_742);
nand U3721 (N_3721,N_2457,N_2233);
and U3722 (N_3722,N_570,N_1291);
and U3723 (N_3723,N_2034,N_863);
xnor U3724 (N_3724,N_1525,N_47);
or U3725 (N_3725,N_1347,N_95);
or U3726 (N_3726,N_2668,N_220);
xnor U3727 (N_3727,N_193,N_2527);
or U3728 (N_3728,N_560,N_2463);
and U3729 (N_3729,N_2401,N_2528);
or U3730 (N_3730,N_1642,N_739);
and U3731 (N_3731,N_1761,N_2787);
or U3732 (N_3732,N_127,N_2428);
xor U3733 (N_3733,N_1334,N_1646);
nor U3734 (N_3734,N_1431,N_119);
nor U3735 (N_3735,N_912,N_65);
nor U3736 (N_3736,N_227,N_2807);
nand U3737 (N_3737,N_551,N_48);
or U3738 (N_3738,N_2641,N_1067);
nand U3739 (N_3739,N_2901,N_2849);
and U3740 (N_3740,N_1865,N_1711);
nand U3741 (N_3741,N_2325,N_727);
nand U3742 (N_3742,N_1452,N_1480);
nand U3743 (N_3743,N_1990,N_2898);
nand U3744 (N_3744,N_839,N_568);
or U3745 (N_3745,N_2847,N_1852);
xnor U3746 (N_3746,N_1069,N_1502);
nor U3747 (N_3747,N_2385,N_1324);
or U3748 (N_3748,N_1666,N_2598);
nand U3749 (N_3749,N_702,N_798);
nand U3750 (N_3750,N_2888,N_3045);
and U3751 (N_3751,N_2889,N_1300);
or U3752 (N_3752,N_1720,N_1496);
and U3753 (N_3753,N_1189,N_1076);
nand U3754 (N_3754,N_1598,N_1833);
and U3755 (N_3755,N_1441,N_1955);
nand U3756 (N_3756,N_1932,N_3097);
or U3757 (N_3757,N_2032,N_2910);
and U3758 (N_3758,N_2024,N_541);
or U3759 (N_3759,N_543,N_888);
and U3760 (N_3760,N_2018,N_3055);
xor U3761 (N_3761,N_1743,N_2227);
xor U3762 (N_3762,N_2574,N_1795);
or U3763 (N_3763,N_947,N_2650);
nand U3764 (N_3764,N_1584,N_2415);
nand U3765 (N_3765,N_3092,N_2103);
nor U3766 (N_3766,N_2013,N_184);
xnor U3767 (N_3767,N_889,N_1101);
xnor U3768 (N_3768,N_49,N_1286);
and U3769 (N_3769,N_2575,N_1160);
nor U3770 (N_3770,N_391,N_750);
xor U3771 (N_3771,N_2094,N_2844);
xor U3772 (N_3772,N_673,N_1659);
or U3773 (N_3773,N_37,N_1429);
nor U3774 (N_3774,N_1812,N_3038);
nand U3775 (N_3775,N_545,N_600);
xnor U3776 (N_3776,N_1443,N_2487);
and U3777 (N_3777,N_2521,N_2240);
nand U3778 (N_3778,N_2459,N_2467);
nor U3779 (N_3779,N_1608,N_3022);
and U3780 (N_3780,N_409,N_890);
and U3781 (N_3781,N_2435,N_3068);
xnor U3782 (N_3782,N_1996,N_623);
or U3783 (N_3783,N_375,N_1109);
nand U3784 (N_3784,N_138,N_540);
or U3785 (N_3785,N_3019,N_2286);
nor U3786 (N_3786,N_2741,N_215);
nor U3787 (N_3787,N_2743,N_806);
nand U3788 (N_3788,N_909,N_2902);
nand U3789 (N_3789,N_1295,N_594);
and U3790 (N_3790,N_2950,N_1811);
and U3791 (N_3791,N_2378,N_418);
and U3792 (N_3792,N_159,N_1150);
nor U3793 (N_3793,N_1219,N_1514);
nand U3794 (N_3794,N_21,N_529);
and U3795 (N_3795,N_1681,N_2816);
nor U3796 (N_3796,N_1778,N_821);
or U3797 (N_3797,N_2819,N_877);
and U3798 (N_3798,N_2739,N_972);
and U3799 (N_3799,N_2155,N_372);
xor U3800 (N_3800,N_1941,N_571);
nor U3801 (N_3801,N_811,N_476);
xor U3802 (N_3802,N_1427,N_1238);
or U3803 (N_3803,N_2377,N_492);
nor U3804 (N_3804,N_581,N_1249);
nand U3805 (N_3805,N_1383,N_785);
or U3806 (N_3806,N_429,N_2828);
xor U3807 (N_3807,N_628,N_1105);
or U3808 (N_3808,N_1491,N_2396);
nor U3809 (N_3809,N_2036,N_26);
nor U3810 (N_3810,N_3121,N_22);
xor U3811 (N_3811,N_2800,N_2051);
or U3812 (N_3812,N_1036,N_6);
or U3813 (N_3813,N_2441,N_1363);
nor U3814 (N_3814,N_1597,N_2717);
nor U3815 (N_3815,N_1968,N_111);
nor U3816 (N_3816,N_988,N_2088);
or U3817 (N_3817,N_554,N_1535);
and U3818 (N_3818,N_2730,N_367);
or U3819 (N_3819,N_1369,N_1877);
and U3820 (N_3820,N_257,N_2315);
nand U3821 (N_3821,N_984,N_1190);
and U3822 (N_3822,N_97,N_832);
nand U3823 (N_3823,N_1341,N_2824);
and U3824 (N_3824,N_1477,N_52);
nor U3825 (N_3825,N_1129,N_2792);
nor U3826 (N_3826,N_2301,N_1362);
and U3827 (N_3827,N_489,N_1648);
or U3828 (N_3828,N_2493,N_857);
nand U3829 (N_3829,N_1280,N_2984);
nor U3830 (N_3830,N_2705,N_1068);
nor U3831 (N_3831,N_2108,N_943);
or U3832 (N_3832,N_2508,N_2284);
xnor U3833 (N_3833,N_94,N_2104);
nor U3834 (N_3834,N_2049,N_2343);
and U3835 (N_3835,N_66,N_2319);
and U3836 (N_3836,N_580,N_2177);
nor U3837 (N_3837,N_2138,N_1815);
or U3838 (N_3838,N_957,N_265);
nand U3839 (N_3839,N_2607,N_712);
nand U3840 (N_3840,N_297,N_663);
nor U3841 (N_3841,N_417,N_2785);
and U3842 (N_3842,N_337,N_2786);
xnor U3843 (N_3843,N_2421,N_2131);
or U3844 (N_3844,N_1165,N_98);
nor U3845 (N_3845,N_1083,N_463);
and U3846 (N_3846,N_29,N_2506);
nand U3847 (N_3847,N_1669,N_2722);
and U3848 (N_3848,N_2451,N_843);
nand U3849 (N_3849,N_2236,N_2255);
nand U3850 (N_3850,N_613,N_79);
nand U3851 (N_3851,N_1342,N_385);
xnor U3852 (N_3852,N_1054,N_1187);
nand U3853 (N_3853,N_19,N_1762);
or U3854 (N_3854,N_198,N_1177);
nand U3855 (N_3855,N_1388,N_2977);
and U3856 (N_3856,N_2797,N_515);
nand U3857 (N_3857,N_519,N_315);
or U3858 (N_3858,N_1097,N_395);
nor U3859 (N_3859,N_998,N_2342);
and U3860 (N_3860,N_1019,N_2648);
and U3861 (N_3861,N_2258,N_555);
xnor U3862 (N_3862,N_746,N_2678);
or U3863 (N_3863,N_2736,N_2367);
or U3864 (N_3864,N_522,N_355);
nor U3865 (N_3865,N_2252,N_195);
and U3866 (N_3866,N_1789,N_1787);
or U3867 (N_3867,N_439,N_1623);
or U3868 (N_3868,N_2030,N_898);
and U3869 (N_3869,N_32,N_687);
nand U3870 (N_3870,N_855,N_2425);
nand U3871 (N_3871,N_200,N_2664);
and U3872 (N_3872,N_344,N_2967);
or U3873 (N_3873,N_1792,N_1591);
xnor U3874 (N_3874,N_1991,N_2814);
or U3875 (N_3875,N_1590,N_531);
and U3876 (N_3876,N_759,N_1707);
or U3877 (N_3877,N_1318,N_1807);
nand U3878 (N_3878,N_330,N_1839);
nand U3879 (N_3879,N_493,N_2949);
xor U3880 (N_3880,N_647,N_2772);
or U3881 (N_3881,N_2505,N_1094);
or U3882 (N_3882,N_706,N_1868);
nor U3883 (N_3883,N_460,N_955);
nor U3884 (N_3884,N_2896,N_1115);
or U3885 (N_3885,N_1035,N_916);
xor U3886 (N_3886,N_3039,N_247);
and U3887 (N_3887,N_2169,N_696);
nand U3888 (N_3888,N_349,N_875);
or U3889 (N_3889,N_891,N_658);
xnor U3890 (N_3890,N_1031,N_1860);
nor U3891 (N_3891,N_2568,N_2973);
or U3892 (N_3892,N_2799,N_740);
or U3893 (N_3893,N_364,N_149);
or U3894 (N_3894,N_2652,N_871);
nand U3895 (N_3895,N_1564,N_1210);
nand U3896 (N_3896,N_112,N_1572);
and U3897 (N_3897,N_1298,N_520);
xor U3898 (N_3898,N_1284,N_935);
nor U3899 (N_3899,N_2593,N_2653);
nand U3900 (N_3900,N_860,N_1017);
nand U3901 (N_3901,N_1329,N_1715);
or U3902 (N_3902,N_2774,N_2148);
and U3903 (N_3903,N_634,N_1471);
nor U3904 (N_3904,N_345,N_1005);
or U3905 (N_3905,N_1136,N_784);
and U3906 (N_3906,N_840,N_2287);
or U3907 (N_3907,N_165,N_1613);
or U3908 (N_3908,N_559,N_2010);
and U3909 (N_3909,N_584,N_2410);
nand U3910 (N_3910,N_406,N_2776);
nor U3911 (N_3911,N_2723,N_1232);
or U3912 (N_3912,N_1353,N_2698);
or U3913 (N_3913,N_225,N_1827);
xnor U3914 (N_3914,N_1495,N_382);
nor U3915 (N_3915,N_2269,N_2204);
nand U3916 (N_3916,N_2907,N_592);
and U3917 (N_3917,N_1895,N_609);
and U3918 (N_3918,N_3065,N_2891);
and U3919 (N_3919,N_3033,N_2643);
xor U3920 (N_3920,N_1769,N_2361);
nor U3921 (N_3921,N_1670,N_332);
nor U3922 (N_3922,N_1428,N_2304);
nand U3923 (N_3923,N_1201,N_3085);
or U3924 (N_3924,N_262,N_968);
or U3925 (N_3925,N_1858,N_1199);
and U3926 (N_3926,N_2481,N_360);
or U3927 (N_3927,N_2420,N_765);
and U3928 (N_3928,N_1808,N_1282);
and U3929 (N_3929,N_638,N_2335);
or U3930 (N_3930,N_2446,N_1043);
and U3931 (N_3931,N_414,N_824);
or U3932 (N_3932,N_449,N_2022);
or U3933 (N_3933,N_511,N_1565);
and U3934 (N_3934,N_586,N_1790);
or U3935 (N_3935,N_1957,N_2015);
or U3936 (N_3936,N_1166,N_2835);
xnor U3937 (N_3937,N_3000,N_1625);
and U3938 (N_3938,N_461,N_1186);
or U3939 (N_3939,N_2559,N_1651);
and U3940 (N_3940,N_1167,N_2366);
and U3941 (N_3941,N_160,N_126);
and U3942 (N_3942,N_386,N_1128);
nand U3943 (N_3943,N_1985,N_152);
nand U3944 (N_3944,N_979,N_61);
xor U3945 (N_3945,N_194,N_173);
xor U3946 (N_3946,N_2496,N_96);
and U3947 (N_3947,N_2752,N_1710);
or U3948 (N_3948,N_2520,N_2383);
or U3949 (N_3949,N_2975,N_141);
nand U3950 (N_3950,N_2491,N_2654);
and U3951 (N_3951,N_578,N_1102);
nor U3952 (N_3952,N_510,N_1114);
nor U3953 (N_3953,N_1753,N_335);
and U3954 (N_3954,N_191,N_1061);
and U3955 (N_3955,N_2534,N_2600);
nor U3956 (N_3956,N_3018,N_1435);
and U3957 (N_3957,N_3091,N_566);
nand U3958 (N_3958,N_539,N_978);
nand U3959 (N_3959,N_683,N_1712);
or U3960 (N_3960,N_309,N_2196);
or U3961 (N_3961,N_2012,N_627);
and U3962 (N_3962,N_2894,N_1661);
nor U3963 (N_3963,N_2670,N_1726);
or U3964 (N_3964,N_679,N_25);
or U3965 (N_3965,N_2666,N_197);
nor U3966 (N_3966,N_2955,N_168);
nand U3967 (N_3967,N_3058,N_1673);
and U3968 (N_3968,N_1255,N_1117);
and U3969 (N_3969,N_35,N_1756);
and U3970 (N_3970,N_2449,N_2499);
nand U3971 (N_3971,N_2348,N_2206);
nand U3972 (N_3972,N_1217,N_3083);
nand U3973 (N_3973,N_1279,N_1880);
nor U3974 (N_3974,N_719,N_2719);
or U3975 (N_3975,N_218,N_2096);
nand U3976 (N_3976,N_2492,N_196);
nand U3977 (N_3977,N_422,N_1064);
nand U3978 (N_3978,N_86,N_925);
nor U3979 (N_3979,N_1632,N_106);
nor U3980 (N_3980,N_711,N_2436);
nor U3981 (N_3981,N_124,N_1226);
xnor U3982 (N_3982,N_2063,N_614);
or U3983 (N_3983,N_2432,N_1969);
nor U3984 (N_3984,N_1170,N_2261);
nand U3985 (N_3985,N_258,N_1);
and U3986 (N_3986,N_2259,N_503);
nand U3987 (N_3987,N_338,N_205);
nor U3988 (N_3988,N_1874,N_1492);
xnor U3989 (N_3989,N_2838,N_3061);
nand U3990 (N_3990,N_420,N_2490);
and U3991 (N_3991,N_1655,N_1176);
xor U3992 (N_3992,N_472,N_1319);
and U3993 (N_3993,N_334,N_235);
nor U3994 (N_3994,N_1290,N_3086);
nand U3995 (N_3995,N_2197,N_1163);
nor U3996 (N_3996,N_1070,N_590);
nand U3997 (N_3997,N_2422,N_293);
or U3998 (N_3998,N_399,N_563);
xnor U3999 (N_3999,N_68,N_267);
nor U4000 (N_4000,N_2405,N_2270);
nand U4001 (N_4001,N_827,N_2153);
and U4002 (N_4002,N_2375,N_2207);
xor U4003 (N_4003,N_862,N_416);
or U4004 (N_4004,N_2943,N_241);
nand U4005 (N_4005,N_1375,N_2732);
or U4006 (N_4006,N_622,N_2660);
or U4007 (N_4007,N_1688,N_108);
nand U4008 (N_4008,N_2767,N_270);
and U4009 (N_4009,N_1870,N_791);
or U4010 (N_4010,N_2657,N_2756);
xnor U4011 (N_4011,N_1193,N_365);
nand U4012 (N_4012,N_2615,N_3075);
and U4013 (N_4013,N_512,N_83);
and U4014 (N_4014,N_1306,N_3031);
nand U4015 (N_4015,N_808,N_93);
nand U4016 (N_4016,N_940,N_1299);
and U4017 (N_4017,N_2871,N_2124);
or U4018 (N_4018,N_1285,N_1755);
and U4019 (N_4019,N_2102,N_290);
nand U4020 (N_4020,N_2734,N_453);
xor U4021 (N_4021,N_1211,N_923);
and U4022 (N_4022,N_2218,N_1965);
nor U4023 (N_4023,N_823,N_2538);
or U4024 (N_4024,N_44,N_1837);
xnor U4025 (N_4025,N_674,N_1056);
xor U4026 (N_4026,N_1372,N_137);
xor U4027 (N_4027,N_2510,N_2193);
or U4028 (N_4028,N_76,N_358);
xor U4029 (N_4029,N_2372,N_2667);
nor U4030 (N_4030,N_2618,N_1386);
nor U4031 (N_4031,N_1993,N_366);
nand U4032 (N_4032,N_350,N_233);
nor U4033 (N_4033,N_1149,N_664);
nor U4034 (N_4034,N_299,N_2137);
nor U4035 (N_4035,N_2433,N_1905);
nor U4036 (N_4036,N_953,N_2145);
nor U4037 (N_4037,N_2390,N_269);
or U4038 (N_4038,N_1822,N_234);
or U4039 (N_4039,N_1398,N_437);
nor U4040 (N_4040,N_996,N_2479);
nand U4041 (N_4041,N_562,N_1656);
or U4042 (N_4042,N_1081,N_1878);
xnor U4043 (N_4043,N_1272,N_736);
and U4044 (N_4044,N_3106,N_298);
nor U4045 (N_4045,N_1262,N_772);
nand U4046 (N_4046,N_73,N_415);
xnor U4047 (N_4047,N_1180,N_2624);
nand U4048 (N_4048,N_2448,N_574);
nand U4049 (N_4049,N_3094,N_2883);
and U4050 (N_4050,N_346,N_354);
or U4051 (N_4051,N_2046,N_2727);
and U4052 (N_4052,N_1387,N_2246);
nand U4053 (N_4053,N_717,N_705);
xor U4054 (N_4054,N_1668,N_1258);
xor U4055 (N_4055,N_864,N_2703);
or U4056 (N_4056,N_1233,N_1630);
nand U4057 (N_4057,N_2083,N_915);
or U4058 (N_4058,N_1553,N_1270);
nor U4059 (N_4059,N_2706,N_1423);
and U4060 (N_4060,N_1066,N_1104);
or U4061 (N_4061,N_2944,N_2749);
or U4062 (N_4062,N_1737,N_1014);
nand U4063 (N_4063,N_2232,N_2454);
and U4064 (N_4064,N_2834,N_1736);
nand U4065 (N_4065,N_2392,N_2359);
and U4066 (N_4066,N_542,N_3002);
and U4067 (N_4067,N_57,N_323);
and U4068 (N_4068,N_81,N_1148);
and U4069 (N_4069,N_2513,N_714);
nor U4070 (N_4070,N_2926,N_2059);
xnor U4071 (N_4071,N_2127,N_2710);
and U4072 (N_4072,N_467,N_2210);
and U4073 (N_4073,N_2675,N_2642);
nand U4074 (N_4074,N_2713,N_1567);
nand U4075 (N_4075,N_1218,N_3051);
nor U4076 (N_4076,N_236,N_259);
nand U4077 (N_4077,N_1944,N_2952);
nor U4078 (N_4078,N_1616,N_2243);
nor U4079 (N_4079,N_207,N_1335);
and U4080 (N_4080,N_697,N_2474);
nand U4081 (N_4081,N_728,N_1700);
and U4082 (N_4082,N_1635,N_1450);
or U4083 (N_4083,N_232,N_2368);
or U4084 (N_4084,N_997,N_1293);
nand U4085 (N_4085,N_2152,N_1263);
nor U4086 (N_4086,N_281,N_2254);
and U4087 (N_4087,N_1235,N_2761);
nand U4088 (N_4088,N_1785,N_2882);
nor U4089 (N_4089,N_694,N_1976);
nand U4090 (N_4090,N_484,N_1566);
and U4091 (N_4091,N_2777,N_2791);
nor U4092 (N_4092,N_885,N_2014);
nor U4093 (N_4093,N_1004,N_2751);
and U4094 (N_4094,N_1875,N_1313);
xnor U4095 (N_4095,N_2769,N_1440);
nand U4096 (N_4096,N_1543,N_599);
and U4097 (N_4097,N_2986,N_2554);
and U4098 (N_4098,N_2398,N_2874);
and U4099 (N_4099,N_2485,N_1410);
or U4100 (N_4100,N_70,N_1125);
nand U4101 (N_4101,N_2565,N_1594);
and U4102 (N_4102,N_2614,N_1053);
nand U4103 (N_4103,N_2050,N_1554);
or U4104 (N_4104,N_1048,N_1568);
xnor U4105 (N_4105,N_771,N_1012);
and U4106 (N_4106,N_612,N_1733);
nand U4107 (N_4107,N_2118,N_2156);
or U4108 (N_4108,N_1051,N_2663);
nor U4109 (N_4109,N_789,N_671);
or U4110 (N_4110,N_1355,N_175);
xnor U4111 (N_4111,N_1020,N_2318);
nor U4112 (N_4112,N_1507,N_2556);
or U4113 (N_4113,N_1836,N_1522);
nand U4114 (N_4114,N_2339,N_1982);
nor U4115 (N_4115,N_620,N_1746);
nand U4116 (N_4116,N_361,N_110);
and U4117 (N_4117,N_2649,N_3120);
or U4118 (N_4118,N_326,N_2376);
nor U4119 (N_4119,N_1986,N_2693);
nor U4120 (N_4120,N_1143,N_2742);
xnor U4121 (N_4121,N_1842,N_1596);
and U4122 (N_4122,N_780,N_1350);
or U4123 (N_4123,N_1389,N_1862);
nor U4124 (N_4124,N_1721,N_1106);
nand U4125 (N_4125,N_2890,N_2188);
or U4126 (N_4126,N_852,N_2803);
nor U4127 (N_4127,N_2128,N_2599);
and U4128 (N_4128,N_2409,N_1763);
and U4129 (N_4129,N_841,N_502);
nand U4130 (N_4130,N_2918,N_2417);
and U4131 (N_4131,N_3076,N_1605);
or U4132 (N_4132,N_1702,N_296);
nand U4133 (N_4133,N_731,N_960);
nor U4134 (N_4134,N_2567,N_374);
nor U4135 (N_4135,N_2688,N_304);
and U4136 (N_4136,N_316,N_937);
xor U4137 (N_4137,N_704,N_1161);
xnor U4138 (N_4138,N_2523,N_2147);
and U4139 (N_4139,N_455,N_1144);
nor U4140 (N_4140,N_2724,N_2592);
and U4141 (N_4141,N_1195,N_2122);
nand U4142 (N_4142,N_856,N_2121);
nor U4143 (N_4143,N_2726,N_1978);
and U4144 (N_4144,N_1124,N_919);
or U4145 (N_4145,N_2880,N_1489);
and U4146 (N_4146,N_2503,N_2544);
or U4147 (N_4147,N_1343,N_1009);
nand U4148 (N_4148,N_1265,N_2696);
and U4149 (N_4149,N_1434,N_557);
nand U4150 (N_4150,N_140,N_1999);
and U4151 (N_4151,N_2860,N_1497);
nor U4152 (N_4152,N_899,N_2214);
nor U4153 (N_4153,N_2691,N_1824);
nor U4154 (N_4154,N_2267,N_1805);
or U4155 (N_4155,N_884,N_393);
and U4156 (N_4156,N_1901,N_419);
nor U4157 (N_4157,N_1576,N_1802);
or U4158 (N_4158,N_2583,N_1781);
and U4159 (N_4159,N_816,N_870);
and U4160 (N_4160,N_2735,N_652);
or U4161 (N_4161,N_504,N_892);
nand U4162 (N_4162,N_2766,N_685);
xnor U4163 (N_4163,N_1028,N_1974);
and U4164 (N_4164,N_1788,N_272);
and U4165 (N_4165,N_1275,N_1107);
nor U4166 (N_4166,N_2195,N_1221);
nand U4167 (N_4167,N_691,N_306);
nand U4168 (N_4168,N_1348,N_2865);
nand U4169 (N_4169,N_633,N_242);
or U4170 (N_4170,N_1463,N_2988);
nand U4171 (N_4171,N_2821,N_2557);
and U4172 (N_4172,N_1346,N_446);
and U4173 (N_4173,N_567,N_637);
nand U4174 (N_4174,N_2114,N_1164);
xnor U4175 (N_4175,N_2606,N_2748);
and U4176 (N_4176,N_779,N_850);
or U4177 (N_4177,N_3059,N_1137);
and U4178 (N_4178,N_1814,N_1011);
nand U4179 (N_4179,N_2968,N_2837);
nand U4180 (N_4180,N_1044,N_1660);
or U4181 (N_4181,N_1524,N_1856);
or U4182 (N_4182,N_514,N_28);
nand U4183 (N_4183,N_1181,N_2313);
nor U4184 (N_4184,N_2442,N_2183);
nand U4185 (N_4185,N_699,N_2519);
nor U4186 (N_4186,N_1087,N_873);
nor U4187 (N_4187,N_2775,N_3034);
nor U4188 (N_4188,N_934,N_1899);
nor U4189 (N_4189,N_288,N_427);
nor U4190 (N_4190,N_1000,N_1473);
xnor U4191 (N_4191,N_1904,N_263);
or U4192 (N_4192,N_518,N_2927);
nor U4193 (N_4193,N_433,N_125);
or U4194 (N_4194,N_190,N_2576);
or U4195 (N_4195,N_1928,N_2798);
nand U4196 (N_4196,N_1065,N_2073);
and U4197 (N_4197,N_90,N_2517);
nor U4198 (N_4198,N_961,N_956);
and U4199 (N_4199,N_1533,N_216);
or U4200 (N_4200,N_1046,N_1582);
and U4201 (N_4201,N_1122,N_591);
and U4202 (N_4202,N_2164,N_1636);
and U4203 (N_4203,N_1832,N_920);
nor U4204 (N_4204,N_2080,N_320);
nand U4205 (N_4205,N_2781,N_1079);
xor U4206 (N_4206,N_243,N_2570);
and U4207 (N_4207,N_2966,N_995);
nor U4208 (N_4208,N_1983,N_2190);
nand U4209 (N_4209,N_2052,N_2109);
and U4210 (N_4210,N_252,N_921);
nor U4211 (N_4211,N_1940,N_3042);
and U4212 (N_4212,N_78,N_1085);
nand U4213 (N_4213,N_1714,N_2115);
or U4214 (N_4214,N_794,N_651);
xnor U4215 (N_4215,N_1851,N_1759);
and U4216 (N_4216,N_2680,N_1243);
nor U4217 (N_4217,N_1798,N_1287);
nand U4218 (N_4218,N_351,N_1678);
and U4219 (N_4219,N_325,N_1175);
or U4220 (N_4220,N_721,N_963);
and U4221 (N_4221,N_356,N_973);
nor U4222 (N_4222,N_506,N_2345);
and U4223 (N_4223,N_1517,N_981);
nand U4224 (N_4224,N_734,N_3124);
and U4225 (N_4225,N_2276,N_1049);
and U4226 (N_4226,N_2694,N_903);
nand U4227 (N_4227,N_371,N_1312);
and U4228 (N_4228,N_353,N_3080);
nand U4229 (N_4229,N_2846,N_809);
nor U4230 (N_4230,N_217,N_992);
nand U4231 (N_4231,N_145,N_264);
nand U4232 (N_4232,N_2879,N_481);
or U4233 (N_4233,N_3028,N_2002);
or U4234 (N_4234,N_2382,N_1321);
nor U4235 (N_4235,N_538,N_1098);
and U4236 (N_4236,N_1459,N_2092);
nand U4237 (N_4237,N_3021,N_668);
nand U4238 (N_4238,N_2241,N_781);
nand U4239 (N_4239,N_1015,N_1680);
nor U4240 (N_4240,N_1841,N_2912);
nand U4241 (N_4241,N_1113,N_2877);
and U4242 (N_4242,N_2113,N_1340);
and U4243 (N_4243,N_2106,N_2689);
and U4244 (N_4244,N_1747,N_2042);
and U4245 (N_4245,N_2906,N_2480);
nand U4246 (N_4246,N_88,N_2584);
nand U4247 (N_4247,N_491,N_1929);
nor U4248 (N_4248,N_653,N_8);
or U4249 (N_4249,N_869,N_748);
nand U4250 (N_4250,N_1916,N_2976);
nor U4251 (N_4251,N_2937,N_2836);
or U4252 (N_4252,N_2711,N_1848);
or U4253 (N_4253,N_295,N_1072);
and U4254 (N_4254,N_1843,N_1330);
or U4255 (N_4255,N_2126,N_1192);
and U4256 (N_4256,N_2931,N_1446);
or U4257 (N_4257,N_2295,N_917);
nand U4258 (N_4258,N_1820,N_3046);
nor U4259 (N_4259,N_535,N_1131);
and U4260 (N_4260,N_2351,N_1512);
nand U4261 (N_4261,N_3110,N_1975);
and U4262 (N_4262,N_84,N_1542);
or U4263 (N_4263,N_2497,N_932);
or U4264 (N_4264,N_1229,N_1444);
xor U4265 (N_4265,N_2460,N_807);
nor U4266 (N_4266,N_1345,N_231);
nand U4267 (N_4267,N_1883,N_1316);
nor U4268 (N_4268,N_3029,N_3073);
xor U4269 (N_4269,N_1409,N_2733);
or U4270 (N_4270,N_2237,N_868);
nand U4271 (N_4271,N_2081,N_3007);
or U4272 (N_4272,N_1693,N_1729);
nor U4273 (N_4273,N_1042,N_2198);
and U4274 (N_4274,N_575,N_115);
or U4275 (N_4275,N_799,N_2993);
and U4276 (N_4276,N_1885,N_1618);
or U4277 (N_4277,N_2475,N_2655);
nand U4278 (N_4278,N_2076,N_1627);
and U4279 (N_4279,N_457,N_151);
or U4280 (N_4280,N_0,N_12);
and U4281 (N_4281,N_2171,N_2434);
nor U4282 (N_4282,N_2978,N_1140);
nor U4283 (N_4283,N_448,N_2941);
xor U4284 (N_4284,N_2166,N_2443);
nand U4285 (N_4285,N_907,N_530);
nand U4286 (N_4286,N_1397,N_2923);
and U4287 (N_4287,N_1182,N_2594);
or U4288 (N_4288,N_1311,N_656);
and U4289 (N_4289,N_1403,N_2299);
nor U4290 (N_4290,N_1551,N_1418);
xnor U4291 (N_4291,N_1251,N_3011);
or U4292 (N_4292,N_1518,N_1261);
nand U4293 (N_4293,N_2760,N_63);
nor U4294 (N_4294,N_2954,N_2994);
nor U4295 (N_4295,N_2229,N_2617);
nand U4296 (N_4296,N_2878,N_1224);
or U4297 (N_4297,N_256,N_2511);
nand U4298 (N_4298,N_2935,N_1708);
nand U4299 (N_4299,N_2801,N_818);
or U4300 (N_4300,N_1026,N_733);
xor U4301 (N_4301,N_618,N_949);
nand U4302 (N_4302,N_1544,N_2412);
nand U4303 (N_4303,N_2754,N_1304);
nand U4304 (N_4304,N_1951,N_321);
xor U4305 (N_4305,N_1511,N_2999);
nand U4306 (N_4306,N_1672,N_2852);
nor U4307 (N_4307,N_1909,N_402);
or U4308 (N_4308,N_442,N_1191);
and U4309 (N_4309,N_1460,N_223);
nor U4310 (N_4310,N_2029,N_254);
or U4311 (N_4311,N_2484,N_72);
nand U4312 (N_4312,N_2107,N_1373);
nor U4313 (N_4313,N_2985,N_2796);
xnor U4314 (N_4314,N_2402,N_2876);
nor U4315 (N_4315,N_1381,N_2861);
or U4316 (N_4316,N_1846,N_180);
or U4317 (N_4317,N_1438,N_1857);
nor U4318 (N_4318,N_1206,N_210);
and U4319 (N_4319,N_544,N_1663);
or U4320 (N_4320,N_1869,N_2916);
nand U4321 (N_4321,N_1838,N_2486);
nor U4322 (N_4322,N_2957,N_1138);
or U4323 (N_4323,N_1088,N_1724);
nor U4324 (N_4324,N_2588,N_3047);
and U4325 (N_4325,N_2630,N_2522);
or U4326 (N_4326,N_1645,N_1538);
nand U4327 (N_4327,N_3004,N_1464);
nor U4328 (N_4328,N_1643,N_669);
nand U4329 (N_4329,N_883,N_1804);
nand U4330 (N_4330,N_1912,N_1977);
or U4331 (N_4331,N_565,N_1040);
or U4332 (N_4332,N_1472,N_1622);
or U4333 (N_4333,N_1766,N_1606);
nor U4334 (N_4334,N_2917,N_275);
or U4335 (N_4335,N_2023,N_2453);
and U4336 (N_4336,N_3095,N_796);
and U4337 (N_4337,N_1774,N_585);
xor U4338 (N_4338,N_2533,N_701);
nor U4339 (N_4339,N_3113,N_2338);
nand U4340 (N_4340,N_1208,N_1764);
nor U4341 (N_4341,N_2765,N_790);
nor U4342 (N_4342,N_237,N_1354);
nand U4343 (N_4343,N_363,N_526);
and U4344 (N_4344,N_2132,N_1775);
and U4345 (N_4345,N_632,N_473);
or U4346 (N_4346,N_77,N_1686);
nand U4347 (N_4347,N_3107,N_2564);
and U4348 (N_4348,N_2611,N_1816);
nand U4349 (N_4349,N_1728,N_1130);
nand U4350 (N_4350,N_1142,N_341);
and U4351 (N_4351,N_2959,N_834);
nand U4352 (N_4352,N_2516,N_1302);
nand U4353 (N_4353,N_2245,N_2291);
xor U4354 (N_4354,N_1332,N_3090);
nor U4355 (N_4355,N_3088,N_2731);
xnor U4356 (N_4356,N_3043,N_3026);
nor U4357 (N_4357,N_1585,N_593);
nor U4358 (N_4358,N_3100,N_800);
xnor U4359 (N_4359,N_2697,N_2101);
and U4360 (N_4360,N_1501,N_2895);
or U4361 (N_4361,N_2525,N_2665);
nor U4362 (N_4362,N_1624,N_384);
and U4363 (N_4363,N_2020,N_649);
or U4364 (N_4364,N_2025,N_675);
xnor U4365 (N_4365,N_2388,N_162);
and U4366 (N_4366,N_201,N_7);
nor U4367 (N_4367,N_2327,N_2084);
nor U4368 (N_4368,N_107,N_2647);
nor U4369 (N_4369,N_805,N_495);
and U4370 (N_4370,N_2669,N_1599);
nor U4371 (N_4371,N_2230,N_3116);
and U4372 (N_4372,N_1586,N_2716);
or U4373 (N_4373,N_639,N_946);
and U4374 (N_4374,N_1419,N_2645);
and U4375 (N_4375,N_1408,N_1583);
nor U4376 (N_4376,N_3072,N_3036);
and U4377 (N_4377,N_2395,N_1555);
and U4378 (N_4378,N_167,N_2429);
or U4379 (N_4379,N_588,N_144);
nor U4380 (N_4380,N_2946,N_1731);
nand U4381 (N_4381,N_1872,N_313);
and U4382 (N_4382,N_2365,N_1432);
or U4383 (N_4383,N_1917,N_2384);
nor U4384 (N_4384,N_1308,N_1683);
nor U4385 (N_4385,N_2507,N_1273);
and U4386 (N_4386,N_1439,N_1657);
xnor U4387 (N_4387,N_1665,N_131);
or U4388 (N_4388,N_244,N_2374);
nor U4389 (N_4389,N_2041,N_2682);
nor U4390 (N_4390,N_1260,N_1296);
nor U4391 (N_4391,N_1692,N_1294);
or U4392 (N_4392,N_1676,N_508);
or U4393 (N_4393,N_443,N_477);
nand U4394 (N_4394,N_1173,N_1360);
xnor U4395 (N_4395,N_597,N_1773);
nand U4396 (N_4396,N_1183,N_672);
nand U4397 (N_4397,N_1647,N_2089);
nor U4398 (N_4398,N_39,N_2180);
and U4399 (N_4399,N_2016,N_2125);
and U4400 (N_4400,N_2512,N_9);
nand U4401 (N_4401,N_2264,N_684);
or U4402 (N_4402,N_2672,N_1793);
nor U4403 (N_4403,N_2312,N_134);
and U4404 (N_4404,N_15,N_1784);
nand U4405 (N_4405,N_2075,N_2347);
nor U4406 (N_4406,N_752,N_185);
or U4407 (N_4407,N_1749,N_954);
and U4408 (N_4408,N_2919,N_3037);
nor U4409 (N_4409,N_2578,N_2005);
nor U4410 (N_4410,N_276,N_2326);
and U4411 (N_4411,N_18,N_1414);
nor U4412 (N_4412,N_128,N_428);
nor U4413 (N_4413,N_2086,N_1380);
nor U4414 (N_4414,N_2473,N_787);
or U4415 (N_4415,N_2352,N_573);
or U4416 (N_4416,N_3084,N_534);
nand U4417 (N_4417,N_2603,N_2644);
or U4418 (N_4418,N_2208,N_1819);
and U4419 (N_4419,N_894,N_2133);
and U4420 (N_4420,N_3062,N_2913);
nor U4421 (N_4421,N_2833,N_1863);
nor U4422 (N_4422,N_828,N_261);
xnor U4423 (N_4423,N_2832,N_2048);
nor U4424 (N_4424,N_1685,N_999);
nand U4425 (N_4425,N_2629,N_319);
nor U4426 (N_4426,N_2117,N_1103);
nor U4427 (N_4427,N_2316,N_2858);
or U4428 (N_4428,N_1021,N_1155);
nor U4429 (N_4429,N_2936,N_2082);
or U4430 (N_4430,N_64,N_910);
nor U4431 (N_4431,N_1571,N_471);
and U4432 (N_4432,N_284,N_2940);
nor U4433 (N_4433,N_2579,N_2746);
nand U4434 (N_4434,N_646,N_2306);
nand U4435 (N_4435,N_2288,N_1910);
or U4436 (N_4436,N_757,N_1458);
nor U4437 (N_4437,N_1948,N_2231);
or U4438 (N_4438,N_1876,N_2920);
nor U4439 (N_4439,N_1479,N_2341);
nand U4440 (N_4440,N_939,N_1701);
nor U4441 (N_4441,N_147,N_2831);
nor U4442 (N_4442,N_2561,N_148);
nand U4443 (N_4443,N_2328,N_948);
nor U4444 (N_4444,N_2165,N_31);
or U4445 (N_4445,N_758,N_1456);
nor U4446 (N_4446,N_1344,N_1091);
nand U4447 (N_4447,N_2964,N_357);
nor U4448 (N_4448,N_246,N_985);
nand U4449 (N_4449,N_1537,N_2620);
nor U4450 (N_4450,N_2311,N_1080);
nand U4451 (N_4451,N_1667,N_2045);
nand U4452 (N_4452,N_1486,N_2176);
and U4453 (N_4453,N_2602,N_3017);
nor U4454 (N_4454,N_1980,N_886);
and U4455 (N_4455,N_902,N_2294);
nand U4456 (N_4456,N_1385,N_336);
nor U4457 (N_4457,N_132,N_1742);
or U4458 (N_4458,N_2008,N_1718);
and U4459 (N_4459,N_1922,N_1123);
nor U4460 (N_4460,N_170,N_513);
nand U4461 (N_4461,N_926,N_2676);
nor U4462 (N_4462,N_1361,N_2144);
and U4463 (N_4463,N_1367,N_952);
or U4464 (N_4464,N_1303,N_253);
and U4465 (N_4465,N_2573,N_3108);
nor U4466 (N_4466,N_209,N_2488);
and U4467 (N_4467,N_2203,N_456);
nor U4468 (N_4468,N_810,N_2431);
and U4469 (N_4469,N_604,N_2151);
nand U4470 (N_4470,N_2399,N_1032);
nor U4471 (N_4471,N_2784,N_987);
or U4472 (N_4472,N_435,N_85);
nand U4473 (N_4473,N_2839,N_2090);
nor U4474 (N_4474,N_2924,N_400);
nor U4475 (N_4475,N_1003,N_1349);
nor U4476 (N_4476,N_1739,N_2679);
xor U4477 (N_4477,N_468,N_608);
and U4478 (N_4478,N_546,N_490);
nand U4479 (N_4479,N_1077,N_769);
nor U4480 (N_4480,N_105,N_135);
or U4481 (N_4481,N_1609,N_831);
and U4482 (N_4482,N_3024,N_2054);
and U4483 (N_4483,N_1958,N_331);
or U4484 (N_4484,N_1526,N_2170);
nand U4485 (N_4485,N_1574,N_595);
nor U4486 (N_4486,N_3063,N_901);
xnor U4487 (N_4487,N_754,N_2456);
and U4488 (N_4488,N_71,N_328);
and U4489 (N_4489,N_1121,N_2662);
xnor U4490 (N_4490,N_239,N_307);
nand U4491 (N_4491,N_2140,N_381);
nor U4492 (N_4492,N_2200,N_1269);
and U4493 (N_4493,N_552,N_725);
nand U4494 (N_4494,N_92,N_2762);
nand U4495 (N_4495,N_1752,N_2031);
or U4496 (N_4496,N_383,N_703);
xor U4497 (N_4497,N_1652,N_2323);
xnor U4498 (N_4498,N_1268,N_763);
nand U4499 (N_4499,N_2808,N_1600);
nor U4500 (N_4500,N_2768,N_2293);
or U4501 (N_4501,N_2514,N_1531);
nor U4502 (N_4502,N_3014,N_1084);
or U4503 (N_4503,N_1390,N_844);
nor U4504 (N_4504,N_1699,N_387);
nor U4505 (N_4505,N_1205,N_2589);
and U4506 (N_4506,N_120,N_708);
xor U4507 (N_4507,N_1248,N_377);
or U4508 (N_4508,N_432,N_1402);
nand U4509 (N_4509,N_1882,N_45);
xnor U4510 (N_4510,N_1215,N_1467);
or U4511 (N_4511,N_188,N_1470);
nand U4512 (N_4512,N_2219,N_1595);
nor U4513 (N_4513,N_424,N_1207);
and U4514 (N_4514,N_2098,N_830);
nand U4515 (N_4515,N_1552,N_16);
and U4516 (N_4516,N_2437,N_1151);
nand U4517 (N_4517,N_788,N_1240);
nand U4518 (N_4518,N_1309,N_3087);
and U4519 (N_4519,N_2167,N_1735);
nand U4520 (N_4520,N_2566,N_2502);
and U4521 (N_4521,N_2310,N_1536);
or U4522 (N_4522,N_1500,N_1050);
and U4523 (N_4523,N_99,N_3049);
nand U4524 (N_4524,N_1589,N_23);
or U4525 (N_4525,N_1469,N_2364);
or U4526 (N_4526,N_1052,N_451);
nand U4527 (N_4527,N_896,N_2795);
xor U4528 (N_4528,N_2863,N_2011);
or U4529 (N_4529,N_1276,N_648);
xnor U4530 (N_4530,N_1649,N_285);
or U4531 (N_4531,N_1013,N_1267);
xnor U4532 (N_4532,N_2268,N_172);
or U4533 (N_4533,N_1411,N_2992);
nor U4534 (N_4534,N_2262,N_2659);
xnor U4535 (N_4535,N_2661,N_2631);
nand U4536 (N_4536,N_2718,N_2690);
nor U4537 (N_4537,N_2868,N_2471);
and U4538 (N_4538,N_2604,N_1997);
nor U4539 (N_4539,N_2515,N_1898);
or U4540 (N_4540,N_1030,N_2027);
nand U4541 (N_4541,N_1029,N_2216);
xor U4542 (N_4542,N_179,N_2360);
nor U4543 (N_4543,N_2004,N_616);
nor U4544 (N_4544,N_452,N_938);
xnor U4545 (N_4545,N_732,N_1704);
nor U4546 (N_4546,N_2223,N_770);
and U4547 (N_4547,N_2921,N_2157);
nor U4548 (N_4548,N_1521,N_1022);
nand U4549 (N_4549,N_1395,N_2770);
or U4550 (N_4550,N_2273,N_1529);
nand U4551 (N_4551,N_274,N_431);
or U4552 (N_4552,N_2822,N_441);
nor U4553 (N_4553,N_881,N_1915);
nor U4554 (N_4554,N_1754,N_1937);
nor U4555 (N_4555,N_17,N_408);
or U4556 (N_4556,N_2370,N_2859);
or U4557 (N_4557,N_1933,N_1337);
or U4558 (N_4558,N_2704,N_723);
or U4559 (N_4559,N_1002,N_1157);
or U4560 (N_4560,N_532,N_1930);
nand U4561 (N_4561,N_1154,N_104);
nor U4562 (N_4562,N_2571,N_2773);
nor U4563 (N_4563,N_1278,N_2355);
or U4564 (N_4564,N_50,N_2915);
and U4565 (N_4565,N_2980,N_2172);
or U4566 (N_4566,N_2869,N_1146);
nand U4567 (N_4567,N_2778,N_621);
or U4568 (N_4568,N_2489,N_2087);
nor U4569 (N_4569,N_582,N_2626);
or U4570 (N_4570,N_695,N_69);
and U4571 (N_4571,N_2142,N_1198);
or U4572 (N_4572,N_164,N_189);
and U4573 (N_4573,N_211,N_2057);
or U4574 (N_4574,N_1971,N_373);
and U4575 (N_4575,N_2297,N_1640);
or U4576 (N_4576,N_2416,N_245);
or U4577 (N_4577,N_1378,N_1204);
nor U4578 (N_4578,N_2963,N_238);
nand U4579 (N_4579,N_523,N_2224);
or U4580 (N_4580,N_2199,N_3105);
or U4581 (N_4581,N_454,N_1579);
or U4582 (N_4582,N_302,N_369);
nor U4583 (N_4583,N_611,N_278);
xor U4584 (N_4584,N_1326,N_2979);
or U4585 (N_4585,N_3023,N_1547);
nor U4586 (N_4586,N_483,N_741);
xor U4587 (N_4587,N_2407,N_2737);
and U4588 (N_4588,N_1853,N_1424);
nand U4589 (N_4589,N_1777,N_2811);
nand U4590 (N_4590,N_2622,N_2707);
or U4591 (N_4591,N_1690,N_156);
xnor U4592 (N_4592,N_1994,N_991);
and U4593 (N_4593,N_2212,N_1691);
and U4594 (N_4594,N_1938,N_643);
nand U4595 (N_4595,N_2129,N_1626);
and U4596 (N_4596,N_401,N_1449);
and U4597 (N_4597,N_430,N_724);
xnor U4598 (N_4598,N_2061,N_3030);
and U4599 (N_4599,N_2105,N_2187);
nand U4600 (N_4600,N_1783,N_300);
nand U4601 (N_4601,N_2039,N_33);
xor U4602 (N_4602,N_1487,N_1861);
xnor U4603 (N_4603,N_657,N_1641);
xnor U4604 (N_4604,N_829,N_2804);
xnor U4605 (N_4605,N_2391,N_2356);
nor U4606 (N_4606,N_533,N_279);
nand U4607 (N_4607,N_1059,N_587);
nor U4608 (N_4608,N_2414,N_1617);
or U4609 (N_4609,N_1025,N_2536);
nand U4610 (N_4610,N_3025,N_1631);
or U4611 (N_4611,N_75,N_289);
or U4612 (N_4612,N_2182,N_2699);
nor U4613 (N_4613,N_3052,N_3001);
or U4614 (N_4614,N_478,N_3115);
nand U4615 (N_4615,N_2673,N_203);
nor U4616 (N_4616,N_410,N_865);
nor U4617 (N_4617,N_2213,N_2540);
nor U4618 (N_4618,N_550,N_812);
nand U4619 (N_4619,N_2862,N_1682);
or U4620 (N_4620,N_2159,N_3050);
nand U4621 (N_4621,N_412,N_2430);
or U4622 (N_4622,N_2476,N_1352);
or U4623 (N_4623,N_2683,N_904);
xnor U4624 (N_4624,N_2945,N_836);
nand U4625 (N_4625,N_1947,N_2389);
and U4626 (N_4626,N_2178,N_1394);
and U4627 (N_4627,N_1809,N_41);
nor U4628 (N_4628,N_1607,N_1936);
nor U4629 (N_4629,N_1508,N_2333);
and U4630 (N_4630,N_466,N_2146);
nor U4631 (N_4631,N_1664,N_116);
or U4632 (N_4632,N_2222,N_1821);
or U4633 (N_4633,N_1074,N_709);
or U4634 (N_4634,N_3010,N_2905);
and U4635 (N_4635,N_2321,N_819);
nor U4636 (N_4636,N_1830,N_1601);
nor U4637 (N_4637,N_1246,N_2186);
xor U4638 (N_4638,N_577,N_1921);
nor U4639 (N_4639,N_2815,N_872);
and U4640 (N_4640,N_1116,N_1152);
or U4641 (N_4641,N_1696,N_1442);
or U4642 (N_4642,N_1614,N_1513);
and U4643 (N_4643,N_445,N_1227);
or U4644 (N_4644,N_1546,N_280);
and U4645 (N_4645,N_1717,N_117);
nor U4646 (N_4646,N_914,N_1934);
nor U4647 (N_4647,N_2805,N_2627);
or U4648 (N_4648,N_2217,N_1323);
nor U4649 (N_4649,N_2543,N_2524);
nor U4650 (N_4650,N_14,N_605);
or U4651 (N_4651,N_444,N_2995);
and U4652 (N_4652,N_486,N_3012);
nor U4653 (N_4653,N_1421,N_1289);
or U4654 (N_4654,N_710,N_1139);
or U4655 (N_4655,N_1179,N_1939);
and U4656 (N_4656,N_1466,N_2636);
nand U4657 (N_4657,N_2228,N_2830);
xnor U4658 (N_4658,N_768,N_347);
nand U4659 (N_4659,N_2542,N_922);
and U4660 (N_4660,N_2613,N_249);
and U4661 (N_4661,N_2616,N_866);
nand U4662 (N_4662,N_74,N_1482);
or U4663 (N_4663,N_1698,N_1200);
or U4664 (N_4664,N_2397,N_2455);
nand U4665 (N_4665,N_2079,N_1413);
nor U4666 (N_4666,N_2745,N_2595);
and U4667 (N_4667,N_2438,N_1946);
xor U4668 (N_4668,N_1396,N_24);
or U4669 (N_4669,N_654,N_43);
and U4670 (N_4670,N_1476,N_897);
nor U4671 (N_4671,N_2998,N_2332);
nand U4672 (N_4672,N_929,N_1906);
nor U4673 (N_4673,N_2700,N_2209);
nand U4674 (N_4674,N_887,N_693);
nor U4675 (N_4675,N_199,N_1803);
xnor U4676 (N_4676,N_1545,N_3071);
nand U4677 (N_4677,N_2239,N_2292);
and U4678 (N_4678,N_1834,N_1364);
nand U4679 (N_4679,N_2608,N_1145);
nor U4680 (N_4680,N_3081,N_2302);
xor U4681 (N_4681,N_3009,N_405);
xor U4682 (N_4682,N_118,N_362);
or U4683 (N_4683,N_1447,N_1923);
nand U4684 (N_4684,N_2794,N_1730);
nand U4685 (N_4685,N_157,N_1823);
nor U4686 (N_4686,N_1359,N_1697);
nor U4687 (N_4687,N_666,N_1105);
nor U4688 (N_4688,N_2869,N_1044);
xor U4689 (N_4689,N_1222,N_2168);
or U4690 (N_4690,N_252,N_1547);
nor U4691 (N_4691,N_1403,N_2527);
nor U4692 (N_4692,N_2462,N_994);
nor U4693 (N_4693,N_1991,N_2722);
nor U4694 (N_4694,N_231,N_2166);
or U4695 (N_4695,N_2660,N_644);
nand U4696 (N_4696,N_1232,N_2682);
xnor U4697 (N_4697,N_2924,N_731);
nand U4698 (N_4698,N_2484,N_1068);
nor U4699 (N_4699,N_1084,N_3085);
or U4700 (N_4700,N_1997,N_1368);
and U4701 (N_4701,N_731,N_1208);
and U4702 (N_4702,N_1102,N_1050);
nor U4703 (N_4703,N_657,N_1178);
and U4704 (N_4704,N_2228,N_772);
nor U4705 (N_4705,N_2065,N_1671);
nand U4706 (N_4706,N_2215,N_1232);
xnor U4707 (N_4707,N_1773,N_2336);
nand U4708 (N_4708,N_1107,N_1019);
xnor U4709 (N_4709,N_275,N_381);
nand U4710 (N_4710,N_586,N_1270);
and U4711 (N_4711,N_1921,N_1846);
or U4712 (N_4712,N_2698,N_430);
nand U4713 (N_4713,N_1213,N_575);
xor U4714 (N_4714,N_917,N_1152);
and U4715 (N_4715,N_1657,N_461);
nand U4716 (N_4716,N_985,N_1605);
and U4717 (N_4717,N_1049,N_1884);
nand U4718 (N_4718,N_1414,N_410);
nor U4719 (N_4719,N_1788,N_2038);
and U4720 (N_4720,N_1858,N_657);
nand U4721 (N_4721,N_1970,N_1194);
or U4722 (N_4722,N_2085,N_252);
xor U4723 (N_4723,N_1202,N_2205);
and U4724 (N_4724,N_1538,N_2545);
or U4725 (N_4725,N_3085,N_2031);
and U4726 (N_4726,N_1794,N_679);
nand U4727 (N_4727,N_490,N_769);
or U4728 (N_4728,N_1335,N_2538);
nor U4729 (N_4729,N_1402,N_269);
nor U4730 (N_4730,N_382,N_1899);
nor U4731 (N_4731,N_72,N_885);
and U4732 (N_4732,N_3118,N_2957);
nand U4733 (N_4733,N_930,N_1086);
and U4734 (N_4734,N_2044,N_800);
nor U4735 (N_4735,N_2340,N_2354);
and U4736 (N_4736,N_1308,N_2252);
nor U4737 (N_4737,N_1823,N_1059);
nand U4738 (N_4738,N_2795,N_2097);
xnor U4739 (N_4739,N_1004,N_2876);
and U4740 (N_4740,N_287,N_1833);
nand U4741 (N_4741,N_2269,N_80);
xnor U4742 (N_4742,N_1803,N_456);
and U4743 (N_4743,N_550,N_2300);
or U4744 (N_4744,N_200,N_1908);
and U4745 (N_4745,N_2196,N_2633);
nand U4746 (N_4746,N_315,N_2911);
and U4747 (N_4747,N_2037,N_1064);
nor U4748 (N_4748,N_1130,N_1219);
or U4749 (N_4749,N_2581,N_307);
nor U4750 (N_4750,N_2177,N_912);
nand U4751 (N_4751,N_1071,N_2632);
and U4752 (N_4752,N_763,N_1788);
nor U4753 (N_4753,N_1358,N_2425);
and U4754 (N_4754,N_718,N_2087);
nor U4755 (N_4755,N_2545,N_1834);
nor U4756 (N_4756,N_213,N_89);
or U4757 (N_4757,N_1721,N_409);
nor U4758 (N_4758,N_3098,N_2221);
nor U4759 (N_4759,N_896,N_2008);
and U4760 (N_4760,N_494,N_1271);
or U4761 (N_4761,N_140,N_1320);
nor U4762 (N_4762,N_2291,N_113);
nand U4763 (N_4763,N_210,N_476);
and U4764 (N_4764,N_1785,N_2786);
nand U4765 (N_4765,N_2244,N_1668);
nand U4766 (N_4766,N_2993,N_2129);
nand U4767 (N_4767,N_2494,N_2430);
xnor U4768 (N_4768,N_2635,N_2321);
nor U4769 (N_4769,N_1967,N_2425);
nand U4770 (N_4770,N_1992,N_2045);
nor U4771 (N_4771,N_590,N_669);
nand U4772 (N_4772,N_3123,N_1421);
nor U4773 (N_4773,N_1005,N_2137);
or U4774 (N_4774,N_2270,N_153);
nand U4775 (N_4775,N_2075,N_511);
nor U4776 (N_4776,N_1765,N_2162);
or U4777 (N_4777,N_1653,N_946);
nand U4778 (N_4778,N_344,N_957);
nand U4779 (N_4779,N_1133,N_596);
or U4780 (N_4780,N_505,N_1055);
and U4781 (N_4781,N_1409,N_1848);
xor U4782 (N_4782,N_2172,N_152);
nand U4783 (N_4783,N_1200,N_2877);
or U4784 (N_4784,N_2315,N_1394);
nor U4785 (N_4785,N_1500,N_3017);
or U4786 (N_4786,N_189,N_171);
nand U4787 (N_4787,N_1700,N_2374);
nor U4788 (N_4788,N_1775,N_1749);
and U4789 (N_4789,N_2935,N_1396);
or U4790 (N_4790,N_434,N_1255);
nor U4791 (N_4791,N_3022,N_255);
nand U4792 (N_4792,N_2038,N_2146);
or U4793 (N_4793,N_1900,N_537);
nor U4794 (N_4794,N_2880,N_1313);
or U4795 (N_4795,N_1119,N_1398);
and U4796 (N_4796,N_211,N_271);
nand U4797 (N_4797,N_114,N_959);
and U4798 (N_4798,N_225,N_737);
or U4799 (N_4799,N_2476,N_1252);
or U4800 (N_4800,N_2404,N_2296);
nor U4801 (N_4801,N_2836,N_3102);
xnor U4802 (N_4802,N_3034,N_1815);
nor U4803 (N_4803,N_2553,N_1948);
and U4804 (N_4804,N_2637,N_2023);
or U4805 (N_4805,N_1955,N_925);
or U4806 (N_4806,N_621,N_2395);
nand U4807 (N_4807,N_504,N_759);
nor U4808 (N_4808,N_298,N_1298);
and U4809 (N_4809,N_869,N_436);
and U4810 (N_4810,N_2214,N_994);
nand U4811 (N_4811,N_1394,N_2089);
xnor U4812 (N_4812,N_1850,N_766);
nand U4813 (N_4813,N_592,N_2128);
nand U4814 (N_4814,N_1917,N_570);
nand U4815 (N_4815,N_1217,N_1414);
nand U4816 (N_4816,N_8,N_1055);
or U4817 (N_4817,N_848,N_2542);
and U4818 (N_4818,N_470,N_1243);
and U4819 (N_4819,N_2055,N_419);
nand U4820 (N_4820,N_2826,N_2633);
or U4821 (N_4821,N_1172,N_895);
nor U4822 (N_4822,N_2374,N_3084);
nand U4823 (N_4823,N_2837,N_1181);
nor U4824 (N_4824,N_1704,N_734);
or U4825 (N_4825,N_1217,N_2357);
nor U4826 (N_4826,N_177,N_1914);
nand U4827 (N_4827,N_929,N_201);
and U4828 (N_4828,N_623,N_594);
nor U4829 (N_4829,N_2782,N_2792);
xnor U4830 (N_4830,N_2881,N_471);
xnor U4831 (N_4831,N_318,N_1162);
nand U4832 (N_4832,N_2879,N_372);
or U4833 (N_4833,N_2860,N_354);
or U4834 (N_4834,N_86,N_620);
and U4835 (N_4835,N_2136,N_338);
nor U4836 (N_4836,N_1979,N_460);
and U4837 (N_4837,N_116,N_2504);
and U4838 (N_4838,N_528,N_1168);
nand U4839 (N_4839,N_712,N_699);
or U4840 (N_4840,N_1357,N_1027);
or U4841 (N_4841,N_2084,N_276);
nand U4842 (N_4842,N_1718,N_1978);
and U4843 (N_4843,N_2547,N_2743);
or U4844 (N_4844,N_124,N_778);
nand U4845 (N_4845,N_343,N_1565);
and U4846 (N_4846,N_1663,N_742);
nor U4847 (N_4847,N_638,N_2946);
nand U4848 (N_4848,N_1036,N_1369);
nor U4849 (N_4849,N_2175,N_1726);
nand U4850 (N_4850,N_985,N_1023);
or U4851 (N_4851,N_831,N_2941);
nand U4852 (N_4852,N_2700,N_2295);
nand U4853 (N_4853,N_1855,N_1238);
and U4854 (N_4854,N_2599,N_2096);
nor U4855 (N_4855,N_703,N_2053);
and U4856 (N_4856,N_1884,N_2378);
or U4857 (N_4857,N_2353,N_2502);
nor U4858 (N_4858,N_1341,N_2711);
xor U4859 (N_4859,N_2194,N_93);
nand U4860 (N_4860,N_1929,N_1771);
and U4861 (N_4861,N_2503,N_1834);
nand U4862 (N_4862,N_878,N_526);
or U4863 (N_4863,N_1769,N_1655);
or U4864 (N_4864,N_2154,N_3010);
nand U4865 (N_4865,N_2192,N_1522);
or U4866 (N_4866,N_1448,N_887);
or U4867 (N_4867,N_1204,N_1299);
and U4868 (N_4868,N_331,N_1675);
nor U4869 (N_4869,N_2040,N_3043);
xor U4870 (N_4870,N_1947,N_2786);
nand U4871 (N_4871,N_2416,N_2182);
or U4872 (N_4872,N_1081,N_1556);
and U4873 (N_4873,N_1016,N_2170);
or U4874 (N_4874,N_215,N_2545);
nand U4875 (N_4875,N_943,N_2906);
or U4876 (N_4876,N_2835,N_28);
nor U4877 (N_4877,N_2538,N_1254);
nor U4878 (N_4878,N_2639,N_598);
nand U4879 (N_4879,N_1625,N_1643);
and U4880 (N_4880,N_758,N_3092);
and U4881 (N_4881,N_2284,N_2805);
nand U4882 (N_4882,N_2194,N_724);
and U4883 (N_4883,N_2224,N_3071);
nor U4884 (N_4884,N_476,N_1619);
nor U4885 (N_4885,N_610,N_1706);
xor U4886 (N_4886,N_92,N_432);
nand U4887 (N_4887,N_1756,N_2427);
nor U4888 (N_4888,N_34,N_2708);
nor U4889 (N_4889,N_2747,N_736);
nand U4890 (N_4890,N_2411,N_1773);
nand U4891 (N_4891,N_1664,N_2004);
nor U4892 (N_4892,N_248,N_1599);
nor U4893 (N_4893,N_1012,N_1654);
nand U4894 (N_4894,N_1677,N_2466);
nor U4895 (N_4895,N_27,N_2690);
nor U4896 (N_4896,N_2721,N_1048);
and U4897 (N_4897,N_41,N_1914);
xor U4898 (N_4898,N_1020,N_270);
and U4899 (N_4899,N_161,N_2171);
and U4900 (N_4900,N_3004,N_191);
nand U4901 (N_4901,N_2600,N_3053);
or U4902 (N_4902,N_2123,N_1930);
xor U4903 (N_4903,N_1400,N_1697);
nor U4904 (N_4904,N_36,N_1452);
nand U4905 (N_4905,N_716,N_2598);
nand U4906 (N_4906,N_2947,N_2538);
nand U4907 (N_4907,N_1582,N_1300);
nand U4908 (N_4908,N_2378,N_2840);
or U4909 (N_4909,N_311,N_2260);
nand U4910 (N_4910,N_2990,N_1431);
and U4911 (N_4911,N_319,N_2673);
and U4912 (N_4912,N_1432,N_1119);
nand U4913 (N_4913,N_2415,N_244);
and U4914 (N_4914,N_8,N_2874);
xor U4915 (N_4915,N_2341,N_1568);
nor U4916 (N_4916,N_761,N_188);
xnor U4917 (N_4917,N_2625,N_2167);
xor U4918 (N_4918,N_785,N_234);
or U4919 (N_4919,N_3121,N_1096);
and U4920 (N_4920,N_1211,N_1335);
nand U4921 (N_4921,N_4,N_243);
xor U4922 (N_4922,N_150,N_1494);
or U4923 (N_4923,N_1281,N_1899);
and U4924 (N_4924,N_2082,N_147);
or U4925 (N_4925,N_2529,N_627);
and U4926 (N_4926,N_1401,N_396);
nand U4927 (N_4927,N_116,N_2915);
nor U4928 (N_4928,N_821,N_2814);
and U4929 (N_4929,N_1396,N_1630);
xnor U4930 (N_4930,N_2950,N_2629);
and U4931 (N_4931,N_1017,N_763);
xor U4932 (N_4932,N_1960,N_321);
nand U4933 (N_4933,N_1282,N_1601);
or U4934 (N_4934,N_2690,N_254);
and U4935 (N_4935,N_1940,N_1741);
xor U4936 (N_4936,N_3097,N_2357);
and U4937 (N_4937,N_1203,N_642);
or U4938 (N_4938,N_1124,N_1103);
nor U4939 (N_4939,N_1934,N_2153);
nor U4940 (N_4940,N_976,N_423);
nand U4941 (N_4941,N_758,N_2314);
nand U4942 (N_4942,N_169,N_2099);
or U4943 (N_4943,N_985,N_1464);
and U4944 (N_4944,N_1283,N_2421);
and U4945 (N_4945,N_1450,N_1758);
nor U4946 (N_4946,N_343,N_2160);
or U4947 (N_4947,N_2385,N_883);
xor U4948 (N_4948,N_310,N_1683);
and U4949 (N_4949,N_697,N_656);
nand U4950 (N_4950,N_2646,N_1205);
or U4951 (N_4951,N_843,N_1932);
nand U4952 (N_4952,N_721,N_1346);
and U4953 (N_4953,N_1876,N_1725);
or U4954 (N_4954,N_1359,N_2463);
nor U4955 (N_4955,N_902,N_2932);
nor U4956 (N_4956,N_1190,N_3006);
and U4957 (N_4957,N_1028,N_364);
and U4958 (N_4958,N_502,N_2819);
and U4959 (N_4959,N_2207,N_284);
nor U4960 (N_4960,N_95,N_733);
nand U4961 (N_4961,N_942,N_1911);
or U4962 (N_4962,N_754,N_720);
and U4963 (N_4963,N_174,N_565);
xnor U4964 (N_4964,N_748,N_2);
nand U4965 (N_4965,N_814,N_1299);
nor U4966 (N_4966,N_1507,N_188);
or U4967 (N_4967,N_334,N_1547);
nand U4968 (N_4968,N_919,N_1247);
and U4969 (N_4969,N_2164,N_622);
xnor U4970 (N_4970,N_1948,N_2927);
or U4971 (N_4971,N_757,N_310);
and U4972 (N_4972,N_2788,N_2826);
or U4973 (N_4973,N_2751,N_1344);
nand U4974 (N_4974,N_513,N_1669);
or U4975 (N_4975,N_1185,N_2855);
or U4976 (N_4976,N_2149,N_791);
and U4977 (N_4977,N_1044,N_898);
or U4978 (N_4978,N_2218,N_3073);
and U4979 (N_4979,N_2801,N_220);
or U4980 (N_4980,N_2265,N_2770);
or U4981 (N_4981,N_3049,N_2401);
nor U4982 (N_4982,N_2405,N_1149);
nand U4983 (N_4983,N_1042,N_2825);
xor U4984 (N_4984,N_1457,N_3059);
xnor U4985 (N_4985,N_1415,N_1505);
and U4986 (N_4986,N_1064,N_1167);
nor U4987 (N_4987,N_3091,N_1758);
or U4988 (N_4988,N_1944,N_3108);
nand U4989 (N_4989,N_205,N_2021);
or U4990 (N_4990,N_2826,N_861);
or U4991 (N_4991,N_1224,N_646);
xor U4992 (N_4992,N_2164,N_2970);
and U4993 (N_4993,N_1974,N_129);
nand U4994 (N_4994,N_610,N_1953);
and U4995 (N_4995,N_1289,N_1653);
nor U4996 (N_4996,N_1,N_61);
or U4997 (N_4997,N_1279,N_1592);
or U4998 (N_4998,N_2963,N_1949);
and U4999 (N_4999,N_630,N_2897);
and U5000 (N_5000,N_731,N_1188);
and U5001 (N_5001,N_152,N_1604);
and U5002 (N_5002,N_1368,N_1690);
and U5003 (N_5003,N_3009,N_2364);
and U5004 (N_5004,N_109,N_2375);
and U5005 (N_5005,N_757,N_228);
nor U5006 (N_5006,N_1743,N_772);
or U5007 (N_5007,N_2547,N_1316);
nand U5008 (N_5008,N_441,N_2038);
nand U5009 (N_5009,N_419,N_2092);
or U5010 (N_5010,N_2150,N_1663);
nand U5011 (N_5011,N_502,N_2090);
or U5012 (N_5012,N_960,N_1515);
nor U5013 (N_5013,N_2770,N_1775);
nor U5014 (N_5014,N_378,N_2504);
nor U5015 (N_5015,N_1143,N_961);
xor U5016 (N_5016,N_299,N_1879);
and U5017 (N_5017,N_2757,N_1431);
and U5018 (N_5018,N_2911,N_1658);
nand U5019 (N_5019,N_2351,N_1812);
nand U5020 (N_5020,N_2324,N_395);
or U5021 (N_5021,N_2997,N_622);
xor U5022 (N_5022,N_375,N_2657);
nor U5023 (N_5023,N_580,N_1658);
nand U5024 (N_5024,N_942,N_2781);
nor U5025 (N_5025,N_2726,N_2272);
nor U5026 (N_5026,N_703,N_398);
xnor U5027 (N_5027,N_1165,N_1960);
nand U5028 (N_5028,N_983,N_1800);
nor U5029 (N_5029,N_1830,N_1509);
nand U5030 (N_5030,N_531,N_794);
or U5031 (N_5031,N_1636,N_3123);
xor U5032 (N_5032,N_969,N_1496);
or U5033 (N_5033,N_124,N_1097);
nand U5034 (N_5034,N_976,N_1857);
nor U5035 (N_5035,N_1668,N_3088);
and U5036 (N_5036,N_612,N_1497);
nand U5037 (N_5037,N_1235,N_1572);
xnor U5038 (N_5038,N_929,N_99);
nand U5039 (N_5039,N_431,N_2802);
xor U5040 (N_5040,N_3115,N_810);
and U5041 (N_5041,N_463,N_1758);
nor U5042 (N_5042,N_954,N_2032);
and U5043 (N_5043,N_43,N_1806);
and U5044 (N_5044,N_2883,N_1998);
and U5045 (N_5045,N_3118,N_1838);
and U5046 (N_5046,N_1487,N_2859);
or U5047 (N_5047,N_986,N_2736);
and U5048 (N_5048,N_75,N_3072);
and U5049 (N_5049,N_357,N_502);
and U5050 (N_5050,N_2513,N_807);
or U5051 (N_5051,N_1701,N_1731);
and U5052 (N_5052,N_1811,N_2341);
nand U5053 (N_5053,N_2507,N_384);
or U5054 (N_5054,N_205,N_39);
nand U5055 (N_5055,N_1268,N_1108);
nor U5056 (N_5056,N_2281,N_2472);
or U5057 (N_5057,N_124,N_121);
or U5058 (N_5058,N_1288,N_64);
nand U5059 (N_5059,N_771,N_83);
and U5060 (N_5060,N_2646,N_1424);
and U5061 (N_5061,N_1967,N_2146);
or U5062 (N_5062,N_1333,N_2031);
nand U5063 (N_5063,N_3092,N_1144);
and U5064 (N_5064,N_2850,N_740);
nor U5065 (N_5065,N_2072,N_2793);
nor U5066 (N_5066,N_1243,N_65);
or U5067 (N_5067,N_2204,N_146);
nand U5068 (N_5068,N_357,N_1236);
nor U5069 (N_5069,N_468,N_202);
and U5070 (N_5070,N_1348,N_1674);
xor U5071 (N_5071,N_678,N_2255);
and U5072 (N_5072,N_2137,N_1308);
nor U5073 (N_5073,N_1636,N_518);
nor U5074 (N_5074,N_1043,N_858);
and U5075 (N_5075,N_575,N_3099);
and U5076 (N_5076,N_1824,N_2598);
nor U5077 (N_5077,N_2449,N_1624);
nor U5078 (N_5078,N_149,N_2743);
or U5079 (N_5079,N_160,N_2811);
and U5080 (N_5080,N_884,N_2642);
nand U5081 (N_5081,N_595,N_1690);
nand U5082 (N_5082,N_199,N_1991);
and U5083 (N_5083,N_681,N_2031);
or U5084 (N_5084,N_444,N_999);
or U5085 (N_5085,N_1107,N_1453);
nor U5086 (N_5086,N_1627,N_2147);
or U5087 (N_5087,N_370,N_1229);
nand U5088 (N_5088,N_1921,N_1360);
and U5089 (N_5089,N_2710,N_1134);
or U5090 (N_5090,N_2706,N_1575);
or U5091 (N_5091,N_1723,N_1666);
or U5092 (N_5092,N_2058,N_1515);
nor U5093 (N_5093,N_964,N_833);
nor U5094 (N_5094,N_990,N_544);
or U5095 (N_5095,N_818,N_1331);
nand U5096 (N_5096,N_2469,N_1827);
nor U5097 (N_5097,N_2242,N_2135);
nand U5098 (N_5098,N_1613,N_1636);
nor U5099 (N_5099,N_2215,N_3013);
nand U5100 (N_5100,N_2213,N_1930);
or U5101 (N_5101,N_1279,N_506);
nand U5102 (N_5102,N_1004,N_1991);
or U5103 (N_5103,N_2168,N_288);
nor U5104 (N_5104,N_1265,N_1159);
xor U5105 (N_5105,N_2431,N_2877);
and U5106 (N_5106,N_341,N_2081);
nand U5107 (N_5107,N_1734,N_720);
nand U5108 (N_5108,N_1341,N_2442);
nor U5109 (N_5109,N_649,N_2330);
nand U5110 (N_5110,N_1620,N_2262);
or U5111 (N_5111,N_345,N_661);
and U5112 (N_5112,N_2211,N_1435);
nor U5113 (N_5113,N_1731,N_1398);
or U5114 (N_5114,N_387,N_745);
nand U5115 (N_5115,N_321,N_790);
xor U5116 (N_5116,N_1121,N_2186);
and U5117 (N_5117,N_1612,N_1011);
nand U5118 (N_5118,N_2552,N_2897);
and U5119 (N_5119,N_2105,N_2282);
and U5120 (N_5120,N_1313,N_2835);
or U5121 (N_5121,N_2038,N_563);
nand U5122 (N_5122,N_1299,N_2938);
and U5123 (N_5123,N_2539,N_839);
and U5124 (N_5124,N_1575,N_76);
nand U5125 (N_5125,N_600,N_1895);
nor U5126 (N_5126,N_2421,N_2931);
nand U5127 (N_5127,N_617,N_906);
nand U5128 (N_5128,N_575,N_1810);
nand U5129 (N_5129,N_2837,N_1414);
nor U5130 (N_5130,N_1244,N_2633);
nor U5131 (N_5131,N_2514,N_2124);
nand U5132 (N_5132,N_3062,N_1729);
xor U5133 (N_5133,N_1716,N_1092);
or U5134 (N_5134,N_2562,N_2413);
or U5135 (N_5135,N_2367,N_93);
nor U5136 (N_5136,N_262,N_1752);
xnor U5137 (N_5137,N_2401,N_218);
and U5138 (N_5138,N_2087,N_2206);
xor U5139 (N_5139,N_646,N_2151);
nor U5140 (N_5140,N_2575,N_413);
nand U5141 (N_5141,N_2844,N_1960);
xor U5142 (N_5142,N_1847,N_1883);
nand U5143 (N_5143,N_1611,N_1951);
nor U5144 (N_5144,N_1294,N_124);
nor U5145 (N_5145,N_2782,N_1668);
nand U5146 (N_5146,N_1341,N_670);
or U5147 (N_5147,N_1532,N_3004);
or U5148 (N_5148,N_1441,N_1947);
or U5149 (N_5149,N_779,N_946);
and U5150 (N_5150,N_992,N_1796);
or U5151 (N_5151,N_891,N_2427);
and U5152 (N_5152,N_2213,N_1347);
nor U5153 (N_5153,N_1643,N_1309);
nor U5154 (N_5154,N_2507,N_2666);
and U5155 (N_5155,N_1308,N_1319);
and U5156 (N_5156,N_2024,N_2274);
or U5157 (N_5157,N_92,N_2764);
nand U5158 (N_5158,N_2790,N_2997);
xnor U5159 (N_5159,N_3060,N_745);
and U5160 (N_5160,N_762,N_567);
xnor U5161 (N_5161,N_1410,N_2187);
or U5162 (N_5162,N_301,N_1501);
or U5163 (N_5163,N_1010,N_536);
or U5164 (N_5164,N_776,N_2738);
nand U5165 (N_5165,N_2004,N_1724);
and U5166 (N_5166,N_3069,N_1861);
and U5167 (N_5167,N_2040,N_864);
nor U5168 (N_5168,N_2874,N_831);
nand U5169 (N_5169,N_2423,N_2190);
or U5170 (N_5170,N_660,N_1880);
nand U5171 (N_5171,N_488,N_556);
or U5172 (N_5172,N_828,N_2875);
nand U5173 (N_5173,N_2030,N_1570);
nor U5174 (N_5174,N_139,N_710);
nand U5175 (N_5175,N_949,N_479);
nor U5176 (N_5176,N_1179,N_2221);
xor U5177 (N_5177,N_3019,N_880);
nand U5178 (N_5178,N_2857,N_2962);
or U5179 (N_5179,N_1976,N_3097);
and U5180 (N_5180,N_1360,N_2750);
nand U5181 (N_5181,N_1225,N_401);
nor U5182 (N_5182,N_961,N_3012);
nor U5183 (N_5183,N_581,N_1554);
nand U5184 (N_5184,N_1349,N_2968);
and U5185 (N_5185,N_2176,N_387);
and U5186 (N_5186,N_2899,N_616);
xor U5187 (N_5187,N_1690,N_2569);
and U5188 (N_5188,N_2798,N_818);
nand U5189 (N_5189,N_1659,N_3052);
or U5190 (N_5190,N_1990,N_2265);
nor U5191 (N_5191,N_393,N_1845);
nor U5192 (N_5192,N_2408,N_1966);
and U5193 (N_5193,N_705,N_1362);
nand U5194 (N_5194,N_890,N_117);
and U5195 (N_5195,N_1517,N_105);
nand U5196 (N_5196,N_983,N_2939);
nor U5197 (N_5197,N_1426,N_1060);
nand U5198 (N_5198,N_1723,N_38);
nor U5199 (N_5199,N_2720,N_973);
nor U5200 (N_5200,N_2228,N_3100);
xor U5201 (N_5201,N_1768,N_1970);
nor U5202 (N_5202,N_601,N_775);
xnor U5203 (N_5203,N_600,N_500);
or U5204 (N_5204,N_1884,N_2779);
or U5205 (N_5205,N_2500,N_585);
nand U5206 (N_5206,N_969,N_978);
xor U5207 (N_5207,N_1417,N_1706);
nand U5208 (N_5208,N_2608,N_2184);
and U5209 (N_5209,N_2721,N_1730);
and U5210 (N_5210,N_233,N_2801);
nand U5211 (N_5211,N_60,N_2137);
or U5212 (N_5212,N_2222,N_830);
or U5213 (N_5213,N_1700,N_2970);
nor U5214 (N_5214,N_1720,N_970);
nand U5215 (N_5215,N_1910,N_341);
and U5216 (N_5216,N_2974,N_91);
and U5217 (N_5217,N_725,N_2074);
or U5218 (N_5218,N_346,N_1581);
or U5219 (N_5219,N_1977,N_264);
or U5220 (N_5220,N_2380,N_1285);
and U5221 (N_5221,N_1782,N_1287);
or U5222 (N_5222,N_715,N_2714);
and U5223 (N_5223,N_1946,N_2948);
nor U5224 (N_5224,N_569,N_3017);
nand U5225 (N_5225,N_1090,N_1962);
and U5226 (N_5226,N_1864,N_2587);
nand U5227 (N_5227,N_1249,N_1248);
nand U5228 (N_5228,N_2986,N_99);
nand U5229 (N_5229,N_2583,N_2643);
nor U5230 (N_5230,N_1635,N_601);
nand U5231 (N_5231,N_3000,N_1402);
xor U5232 (N_5232,N_1728,N_2740);
and U5233 (N_5233,N_1608,N_267);
and U5234 (N_5234,N_398,N_2187);
or U5235 (N_5235,N_1458,N_2888);
nor U5236 (N_5236,N_549,N_171);
or U5237 (N_5237,N_2254,N_1333);
or U5238 (N_5238,N_2635,N_476);
nand U5239 (N_5239,N_1799,N_2637);
nor U5240 (N_5240,N_1020,N_950);
nand U5241 (N_5241,N_1149,N_2684);
nor U5242 (N_5242,N_415,N_328);
nor U5243 (N_5243,N_2435,N_185);
nand U5244 (N_5244,N_2341,N_325);
or U5245 (N_5245,N_493,N_1480);
and U5246 (N_5246,N_3064,N_550);
nor U5247 (N_5247,N_2158,N_680);
nand U5248 (N_5248,N_2733,N_2923);
or U5249 (N_5249,N_90,N_758);
nand U5250 (N_5250,N_751,N_259);
and U5251 (N_5251,N_2379,N_9);
or U5252 (N_5252,N_1443,N_1329);
nand U5253 (N_5253,N_1247,N_1793);
nand U5254 (N_5254,N_1671,N_128);
or U5255 (N_5255,N_2239,N_1145);
or U5256 (N_5256,N_1569,N_1382);
xnor U5257 (N_5257,N_3000,N_260);
or U5258 (N_5258,N_241,N_2472);
or U5259 (N_5259,N_1185,N_1885);
nand U5260 (N_5260,N_554,N_1970);
nor U5261 (N_5261,N_1705,N_399);
nor U5262 (N_5262,N_160,N_1422);
or U5263 (N_5263,N_809,N_650);
and U5264 (N_5264,N_42,N_2755);
xor U5265 (N_5265,N_1442,N_2355);
nand U5266 (N_5266,N_1263,N_1066);
or U5267 (N_5267,N_1780,N_419);
nand U5268 (N_5268,N_2369,N_558);
nor U5269 (N_5269,N_2469,N_462);
and U5270 (N_5270,N_271,N_2135);
nand U5271 (N_5271,N_648,N_2280);
nor U5272 (N_5272,N_233,N_1512);
nand U5273 (N_5273,N_1873,N_2983);
and U5274 (N_5274,N_1010,N_1521);
nor U5275 (N_5275,N_1843,N_455);
or U5276 (N_5276,N_411,N_356);
nand U5277 (N_5277,N_2281,N_2725);
nor U5278 (N_5278,N_1436,N_2471);
nand U5279 (N_5279,N_2829,N_964);
nor U5280 (N_5280,N_1556,N_789);
or U5281 (N_5281,N_1025,N_2644);
nand U5282 (N_5282,N_241,N_2813);
xor U5283 (N_5283,N_1250,N_700);
and U5284 (N_5284,N_214,N_1524);
nand U5285 (N_5285,N_938,N_1213);
and U5286 (N_5286,N_3066,N_1366);
and U5287 (N_5287,N_1212,N_2814);
or U5288 (N_5288,N_637,N_2523);
nor U5289 (N_5289,N_364,N_1450);
or U5290 (N_5290,N_1877,N_2721);
or U5291 (N_5291,N_1156,N_1035);
or U5292 (N_5292,N_3082,N_248);
xnor U5293 (N_5293,N_928,N_2870);
or U5294 (N_5294,N_562,N_689);
nor U5295 (N_5295,N_1835,N_88);
nand U5296 (N_5296,N_2511,N_2698);
xnor U5297 (N_5297,N_1605,N_2416);
and U5298 (N_5298,N_1354,N_857);
nand U5299 (N_5299,N_2029,N_891);
nand U5300 (N_5300,N_715,N_2466);
and U5301 (N_5301,N_2474,N_3119);
nand U5302 (N_5302,N_1391,N_2180);
and U5303 (N_5303,N_2523,N_2952);
and U5304 (N_5304,N_523,N_1846);
nand U5305 (N_5305,N_2852,N_1839);
nor U5306 (N_5306,N_1878,N_1931);
xor U5307 (N_5307,N_768,N_1312);
nand U5308 (N_5308,N_832,N_2462);
or U5309 (N_5309,N_2039,N_2271);
nand U5310 (N_5310,N_1076,N_478);
nand U5311 (N_5311,N_2910,N_762);
nor U5312 (N_5312,N_743,N_1542);
nor U5313 (N_5313,N_278,N_424);
nor U5314 (N_5314,N_752,N_468);
or U5315 (N_5315,N_111,N_2901);
and U5316 (N_5316,N_1455,N_2068);
nor U5317 (N_5317,N_2134,N_2296);
or U5318 (N_5318,N_974,N_544);
nor U5319 (N_5319,N_2525,N_1554);
nand U5320 (N_5320,N_2781,N_326);
nor U5321 (N_5321,N_2827,N_1294);
xnor U5322 (N_5322,N_327,N_2685);
or U5323 (N_5323,N_1305,N_1034);
or U5324 (N_5324,N_2580,N_1443);
or U5325 (N_5325,N_2064,N_2640);
nor U5326 (N_5326,N_264,N_2705);
nand U5327 (N_5327,N_134,N_730);
and U5328 (N_5328,N_344,N_647);
or U5329 (N_5329,N_1148,N_1840);
nor U5330 (N_5330,N_33,N_1851);
and U5331 (N_5331,N_2328,N_2391);
or U5332 (N_5332,N_387,N_438);
nand U5333 (N_5333,N_1719,N_2116);
nand U5334 (N_5334,N_1285,N_1514);
and U5335 (N_5335,N_630,N_862);
and U5336 (N_5336,N_444,N_94);
nor U5337 (N_5337,N_2842,N_1187);
xor U5338 (N_5338,N_2323,N_200);
or U5339 (N_5339,N_599,N_604);
nand U5340 (N_5340,N_610,N_664);
or U5341 (N_5341,N_2080,N_1102);
xnor U5342 (N_5342,N_874,N_807);
and U5343 (N_5343,N_2481,N_2446);
nor U5344 (N_5344,N_1297,N_2298);
nor U5345 (N_5345,N_1369,N_3086);
nand U5346 (N_5346,N_1584,N_867);
nor U5347 (N_5347,N_360,N_1917);
and U5348 (N_5348,N_2161,N_1829);
nor U5349 (N_5349,N_27,N_111);
nand U5350 (N_5350,N_1122,N_824);
nand U5351 (N_5351,N_1121,N_2413);
nand U5352 (N_5352,N_3062,N_1750);
nor U5353 (N_5353,N_486,N_2690);
nand U5354 (N_5354,N_2856,N_2836);
and U5355 (N_5355,N_163,N_555);
nand U5356 (N_5356,N_2020,N_1894);
nand U5357 (N_5357,N_2008,N_1240);
xor U5358 (N_5358,N_1167,N_1632);
nand U5359 (N_5359,N_2014,N_3007);
nand U5360 (N_5360,N_290,N_1551);
xor U5361 (N_5361,N_2959,N_664);
nand U5362 (N_5362,N_2950,N_907);
and U5363 (N_5363,N_1740,N_922);
nand U5364 (N_5364,N_1503,N_2763);
nor U5365 (N_5365,N_2757,N_1614);
nor U5366 (N_5366,N_704,N_927);
and U5367 (N_5367,N_150,N_2704);
nand U5368 (N_5368,N_2364,N_2077);
or U5369 (N_5369,N_1354,N_859);
and U5370 (N_5370,N_1623,N_193);
or U5371 (N_5371,N_966,N_124);
nand U5372 (N_5372,N_1902,N_1221);
nand U5373 (N_5373,N_970,N_1028);
and U5374 (N_5374,N_2871,N_1597);
nand U5375 (N_5375,N_1310,N_2951);
and U5376 (N_5376,N_89,N_210);
or U5377 (N_5377,N_1166,N_2591);
xnor U5378 (N_5378,N_1596,N_2866);
or U5379 (N_5379,N_1113,N_2291);
nor U5380 (N_5380,N_1725,N_1695);
nand U5381 (N_5381,N_1316,N_429);
nor U5382 (N_5382,N_53,N_1145);
or U5383 (N_5383,N_1074,N_1744);
nand U5384 (N_5384,N_2602,N_1994);
nor U5385 (N_5385,N_2076,N_3106);
nor U5386 (N_5386,N_2562,N_655);
nand U5387 (N_5387,N_3108,N_406);
nand U5388 (N_5388,N_3053,N_1057);
nand U5389 (N_5389,N_803,N_694);
and U5390 (N_5390,N_2236,N_2248);
nor U5391 (N_5391,N_790,N_1670);
nand U5392 (N_5392,N_783,N_607);
or U5393 (N_5393,N_109,N_2587);
nor U5394 (N_5394,N_1146,N_2232);
nor U5395 (N_5395,N_719,N_2073);
or U5396 (N_5396,N_2427,N_622);
nand U5397 (N_5397,N_1183,N_1737);
or U5398 (N_5398,N_135,N_1033);
xnor U5399 (N_5399,N_2883,N_1539);
nand U5400 (N_5400,N_1427,N_2543);
and U5401 (N_5401,N_1770,N_324);
nor U5402 (N_5402,N_2767,N_2802);
nand U5403 (N_5403,N_109,N_1127);
and U5404 (N_5404,N_570,N_2803);
or U5405 (N_5405,N_592,N_11);
nand U5406 (N_5406,N_1907,N_1511);
nor U5407 (N_5407,N_246,N_154);
and U5408 (N_5408,N_1954,N_2107);
nand U5409 (N_5409,N_1353,N_620);
or U5410 (N_5410,N_1814,N_2409);
nor U5411 (N_5411,N_569,N_1852);
nand U5412 (N_5412,N_96,N_802);
or U5413 (N_5413,N_845,N_2434);
or U5414 (N_5414,N_743,N_1274);
nand U5415 (N_5415,N_2428,N_1684);
nand U5416 (N_5416,N_1616,N_2732);
nand U5417 (N_5417,N_2728,N_84);
or U5418 (N_5418,N_2684,N_3086);
xor U5419 (N_5419,N_1338,N_2200);
nor U5420 (N_5420,N_2259,N_2365);
or U5421 (N_5421,N_2331,N_437);
nand U5422 (N_5422,N_2515,N_653);
and U5423 (N_5423,N_361,N_816);
nor U5424 (N_5424,N_2102,N_2914);
nand U5425 (N_5425,N_440,N_2109);
nand U5426 (N_5426,N_1445,N_1007);
or U5427 (N_5427,N_1201,N_775);
or U5428 (N_5428,N_433,N_1097);
or U5429 (N_5429,N_76,N_176);
nand U5430 (N_5430,N_2036,N_1550);
and U5431 (N_5431,N_812,N_432);
or U5432 (N_5432,N_1736,N_530);
or U5433 (N_5433,N_1386,N_2521);
and U5434 (N_5434,N_372,N_2930);
nand U5435 (N_5435,N_7,N_1646);
and U5436 (N_5436,N_2608,N_756);
nor U5437 (N_5437,N_2946,N_2031);
and U5438 (N_5438,N_1536,N_3083);
or U5439 (N_5439,N_1472,N_2822);
xnor U5440 (N_5440,N_2088,N_942);
nand U5441 (N_5441,N_1978,N_386);
nand U5442 (N_5442,N_1972,N_358);
nor U5443 (N_5443,N_108,N_200);
and U5444 (N_5444,N_2159,N_2068);
nand U5445 (N_5445,N_2786,N_212);
or U5446 (N_5446,N_2577,N_1790);
or U5447 (N_5447,N_2865,N_494);
nand U5448 (N_5448,N_3114,N_678);
nor U5449 (N_5449,N_1044,N_2300);
nand U5450 (N_5450,N_2864,N_351);
nor U5451 (N_5451,N_2593,N_2619);
nor U5452 (N_5452,N_1888,N_785);
nand U5453 (N_5453,N_118,N_383);
and U5454 (N_5454,N_1955,N_1997);
and U5455 (N_5455,N_1649,N_2065);
nor U5456 (N_5456,N_42,N_3093);
and U5457 (N_5457,N_3028,N_2612);
or U5458 (N_5458,N_727,N_1638);
nand U5459 (N_5459,N_3076,N_2182);
nor U5460 (N_5460,N_2602,N_838);
xor U5461 (N_5461,N_667,N_1267);
nor U5462 (N_5462,N_895,N_2035);
nor U5463 (N_5463,N_3042,N_214);
nand U5464 (N_5464,N_1858,N_810);
or U5465 (N_5465,N_1145,N_2781);
or U5466 (N_5466,N_256,N_2809);
or U5467 (N_5467,N_471,N_1719);
nand U5468 (N_5468,N_2931,N_1233);
nand U5469 (N_5469,N_2251,N_1030);
nor U5470 (N_5470,N_2009,N_1214);
and U5471 (N_5471,N_1076,N_2308);
or U5472 (N_5472,N_705,N_4);
and U5473 (N_5473,N_3119,N_739);
and U5474 (N_5474,N_2899,N_1835);
nor U5475 (N_5475,N_1569,N_249);
xor U5476 (N_5476,N_2773,N_94);
and U5477 (N_5477,N_572,N_1991);
nand U5478 (N_5478,N_705,N_1301);
nor U5479 (N_5479,N_158,N_50);
nor U5480 (N_5480,N_1453,N_544);
and U5481 (N_5481,N_2970,N_2404);
xor U5482 (N_5482,N_2663,N_340);
and U5483 (N_5483,N_2175,N_2241);
nor U5484 (N_5484,N_1511,N_259);
xnor U5485 (N_5485,N_3113,N_915);
and U5486 (N_5486,N_2610,N_25);
and U5487 (N_5487,N_1667,N_322);
or U5488 (N_5488,N_1222,N_1181);
or U5489 (N_5489,N_1562,N_3052);
nand U5490 (N_5490,N_1825,N_754);
or U5491 (N_5491,N_1065,N_2534);
nand U5492 (N_5492,N_1283,N_2211);
and U5493 (N_5493,N_861,N_1837);
and U5494 (N_5494,N_639,N_1472);
nand U5495 (N_5495,N_476,N_1805);
or U5496 (N_5496,N_1657,N_2775);
and U5497 (N_5497,N_421,N_2110);
or U5498 (N_5498,N_1287,N_958);
nand U5499 (N_5499,N_233,N_1073);
and U5500 (N_5500,N_2170,N_2253);
nor U5501 (N_5501,N_2486,N_2345);
or U5502 (N_5502,N_693,N_143);
or U5503 (N_5503,N_1198,N_307);
nor U5504 (N_5504,N_1501,N_854);
or U5505 (N_5505,N_2461,N_978);
nand U5506 (N_5506,N_497,N_2140);
nor U5507 (N_5507,N_2749,N_558);
nor U5508 (N_5508,N_2428,N_1482);
xnor U5509 (N_5509,N_108,N_2730);
nor U5510 (N_5510,N_2914,N_857);
nor U5511 (N_5511,N_2789,N_12);
xnor U5512 (N_5512,N_1512,N_1994);
xnor U5513 (N_5513,N_1395,N_862);
or U5514 (N_5514,N_436,N_18);
xnor U5515 (N_5515,N_670,N_290);
and U5516 (N_5516,N_2518,N_2545);
nand U5517 (N_5517,N_735,N_993);
or U5518 (N_5518,N_1945,N_966);
nor U5519 (N_5519,N_493,N_2698);
and U5520 (N_5520,N_1262,N_2374);
or U5521 (N_5521,N_2355,N_989);
xnor U5522 (N_5522,N_20,N_1724);
and U5523 (N_5523,N_767,N_2196);
nand U5524 (N_5524,N_161,N_480);
and U5525 (N_5525,N_910,N_2160);
nor U5526 (N_5526,N_352,N_2054);
nand U5527 (N_5527,N_1344,N_2834);
and U5528 (N_5528,N_1338,N_2821);
xnor U5529 (N_5529,N_2162,N_249);
nor U5530 (N_5530,N_2351,N_2313);
or U5531 (N_5531,N_391,N_1364);
nand U5532 (N_5532,N_381,N_2594);
nand U5533 (N_5533,N_1117,N_2772);
or U5534 (N_5534,N_1481,N_2408);
nor U5535 (N_5535,N_1405,N_1621);
xor U5536 (N_5536,N_2682,N_166);
or U5537 (N_5537,N_1364,N_627);
or U5538 (N_5538,N_2296,N_2173);
and U5539 (N_5539,N_3090,N_2112);
nand U5540 (N_5540,N_2446,N_1586);
or U5541 (N_5541,N_2536,N_1887);
and U5542 (N_5542,N_278,N_2555);
nor U5543 (N_5543,N_2785,N_1758);
nand U5544 (N_5544,N_2337,N_167);
nor U5545 (N_5545,N_991,N_777);
or U5546 (N_5546,N_2697,N_925);
nor U5547 (N_5547,N_2821,N_172);
nor U5548 (N_5548,N_1962,N_2528);
xor U5549 (N_5549,N_699,N_789);
or U5550 (N_5550,N_758,N_1114);
xor U5551 (N_5551,N_59,N_3059);
nor U5552 (N_5552,N_1247,N_1311);
nor U5553 (N_5553,N_3079,N_160);
nand U5554 (N_5554,N_1599,N_2190);
nor U5555 (N_5555,N_1114,N_672);
xor U5556 (N_5556,N_812,N_3076);
and U5557 (N_5557,N_992,N_64);
nand U5558 (N_5558,N_378,N_217);
nor U5559 (N_5559,N_1718,N_1773);
and U5560 (N_5560,N_2973,N_720);
nor U5561 (N_5561,N_2659,N_551);
or U5562 (N_5562,N_1238,N_2444);
nand U5563 (N_5563,N_3103,N_761);
nand U5564 (N_5564,N_500,N_423);
xnor U5565 (N_5565,N_1211,N_2464);
or U5566 (N_5566,N_967,N_2402);
nor U5567 (N_5567,N_2126,N_1565);
and U5568 (N_5568,N_3087,N_782);
xor U5569 (N_5569,N_165,N_1593);
or U5570 (N_5570,N_47,N_2416);
and U5571 (N_5571,N_2870,N_372);
nand U5572 (N_5572,N_3083,N_2555);
xnor U5573 (N_5573,N_1194,N_17);
or U5574 (N_5574,N_2981,N_1880);
and U5575 (N_5575,N_156,N_102);
nor U5576 (N_5576,N_2495,N_1368);
and U5577 (N_5577,N_532,N_621);
or U5578 (N_5578,N_2955,N_1299);
or U5579 (N_5579,N_1313,N_2986);
and U5580 (N_5580,N_943,N_2339);
and U5581 (N_5581,N_476,N_2221);
nand U5582 (N_5582,N_2572,N_89);
nor U5583 (N_5583,N_409,N_871);
nor U5584 (N_5584,N_2781,N_1345);
xnor U5585 (N_5585,N_2655,N_1210);
nand U5586 (N_5586,N_2780,N_2833);
nand U5587 (N_5587,N_2913,N_268);
and U5588 (N_5588,N_1220,N_741);
and U5589 (N_5589,N_2200,N_2903);
xnor U5590 (N_5590,N_2919,N_1415);
nand U5591 (N_5591,N_1325,N_74);
nor U5592 (N_5592,N_48,N_2426);
nor U5593 (N_5593,N_582,N_793);
nor U5594 (N_5594,N_326,N_2579);
nor U5595 (N_5595,N_549,N_2684);
or U5596 (N_5596,N_1996,N_3068);
and U5597 (N_5597,N_2320,N_1743);
or U5598 (N_5598,N_2044,N_1442);
or U5599 (N_5599,N_1772,N_2410);
or U5600 (N_5600,N_2690,N_306);
nor U5601 (N_5601,N_1180,N_1599);
nand U5602 (N_5602,N_1532,N_2799);
xor U5603 (N_5603,N_492,N_868);
or U5604 (N_5604,N_3037,N_757);
nor U5605 (N_5605,N_1900,N_701);
nor U5606 (N_5606,N_924,N_1074);
nand U5607 (N_5607,N_2508,N_2581);
nand U5608 (N_5608,N_132,N_2108);
and U5609 (N_5609,N_1934,N_1376);
nand U5610 (N_5610,N_382,N_427);
or U5611 (N_5611,N_1712,N_1101);
nor U5612 (N_5612,N_770,N_1088);
or U5613 (N_5613,N_2074,N_362);
and U5614 (N_5614,N_1471,N_676);
and U5615 (N_5615,N_1386,N_1568);
nor U5616 (N_5616,N_1953,N_1883);
or U5617 (N_5617,N_86,N_1203);
or U5618 (N_5618,N_2057,N_1324);
or U5619 (N_5619,N_812,N_1413);
nand U5620 (N_5620,N_856,N_2146);
xnor U5621 (N_5621,N_3028,N_2167);
and U5622 (N_5622,N_1488,N_732);
and U5623 (N_5623,N_2346,N_776);
nor U5624 (N_5624,N_589,N_1399);
and U5625 (N_5625,N_2374,N_1460);
or U5626 (N_5626,N_2017,N_2787);
xor U5627 (N_5627,N_2983,N_2093);
nor U5628 (N_5628,N_359,N_1740);
nor U5629 (N_5629,N_688,N_341);
nor U5630 (N_5630,N_248,N_1132);
nand U5631 (N_5631,N_288,N_1605);
nor U5632 (N_5632,N_755,N_1803);
and U5633 (N_5633,N_2399,N_1956);
xor U5634 (N_5634,N_2832,N_2918);
or U5635 (N_5635,N_931,N_2013);
and U5636 (N_5636,N_2655,N_200);
xor U5637 (N_5637,N_1211,N_1181);
nand U5638 (N_5638,N_997,N_520);
nor U5639 (N_5639,N_1585,N_1604);
xnor U5640 (N_5640,N_1753,N_301);
or U5641 (N_5641,N_2312,N_2567);
or U5642 (N_5642,N_690,N_2510);
nor U5643 (N_5643,N_1347,N_2554);
nand U5644 (N_5644,N_1425,N_1301);
xor U5645 (N_5645,N_935,N_300);
xor U5646 (N_5646,N_675,N_2854);
nor U5647 (N_5647,N_2838,N_51);
or U5648 (N_5648,N_1166,N_177);
nor U5649 (N_5649,N_3046,N_130);
nand U5650 (N_5650,N_82,N_1194);
nor U5651 (N_5651,N_1052,N_946);
nor U5652 (N_5652,N_2375,N_1640);
or U5653 (N_5653,N_1096,N_954);
nand U5654 (N_5654,N_578,N_1956);
or U5655 (N_5655,N_2531,N_1392);
nor U5656 (N_5656,N_2019,N_1149);
or U5657 (N_5657,N_1147,N_2529);
and U5658 (N_5658,N_263,N_1414);
or U5659 (N_5659,N_834,N_2131);
or U5660 (N_5660,N_249,N_2766);
nand U5661 (N_5661,N_417,N_2777);
and U5662 (N_5662,N_1140,N_372);
and U5663 (N_5663,N_2829,N_540);
nand U5664 (N_5664,N_2619,N_2003);
or U5665 (N_5665,N_1175,N_936);
or U5666 (N_5666,N_2505,N_2904);
nor U5667 (N_5667,N_3104,N_2604);
or U5668 (N_5668,N_484,N_2177);
xnor U5669 (N_5669,N_2999,N_1951);
xnor U5670 (N_5670,N_2193,N_25);
nand U5671 (N_5671,N_17,N_587);
nand U5672 (N_5672,N_595,N_2328);
or U5673 (N_5673,N_1644,N_2462);
nand U5674 (N_5674,N_1873,N_2213);
nor U5675 (N_5675,N_1140,N_1118);
nor U5676 (N_5676,N_1201,N_1743);
and U5677 (N_5677,N_2230,N_50);
nor U5678 (N_5678,N_2815,N_776);
or U5679 (N_5679,N_1527,N_580);
nand U5680 (N_5680,N_1869,N_1786);
and U5681 (N_5681,N_2260,N_620);
and U5682 (N_5682,N_2863,N_795);
or U5683 (N_5683,N_2962,N_2808);
nand U5684 (N_5684,N_34,N_594);
nor U5685 (N_5685,N_2731,N_352);
nor U5686 (N_5686,N_568,N_1506);
xor U5687 (N_5687,N_1797,N_1915);
and U5688 (N_5688,N_599,N_2403);
nand U5689 (N_5689,N_1106,N_2699);
nand U5690 (N_5690,N_1142,N_2083);
or U5691 (N_5691,N_1390,N_2191);
nor U5692 (N_5692,N_1737,N_2432);
or U5693 (N_5693,N_2774,N_2893);
xnor U5694 (N_5694,N_2325,N_1207);
and U5695 (N_5695,N_1399,N_598);
nand U5696 (N_5696,N_212,N_601);
xnor U5697 (N_5697,N_1439,N_2683);
and U5698 (N_5698,N_2427,N_1207);
nand U5699 (N_5699,N_778,N_1274);
and U5700 (N_5700,N_1917,N_1646);
nor U5701 (N_5701,N_643,N_1096);
and U5702 (N_5702,N_3099,N_2529);
nand U5703 (N_5703,N_346,N_534);
and U5704 (N_5704,N_431,N_850);
nor U5705 (N_5705,N_2819,N_919);
nand U5706 (N_5706,N_2349,N_1440);
nand U5707 (N_5707,N_2517,N_1374);
and U5708 (N_5708,N_2260,N_2454);
xnor U5709 (N_5709,N_1808,N_2724);
or U5710 (N_5710,N_2361,N_1877);
or U5711 (N_5711,N_2586,N_588);
xor U5712 (N_5712,N_1195,N_525);
or U5713 (N_5713,N_2376,N_904);
or U5714 (N_5714,N_2835,N_2399);
nor U5715 (N_5715,N_2737,N_2249);
and U5716 (N_5716,N_160,N_2825);
nor U5717 (N_5717,N_2873,N_619);
nor U5718 (N_5718,N_1646,N_1834);
or U5719 (N_5719,N_1192,N_2911);
and U5720 (N_5720,N_3051,N_2424);
nor U5721 (N_5721,N_375,N_1051);
nand U5722 (N_5722,N_768,N_2170);
or U5723 (N_5723,N_1738,N_3052);
nor U5724 (N_5724,N_954,N_3022);
nor U5725 (N_5725,N_527,N_438);
nand U5726 (N_5726,N_2076,N_1515);
nor U5727 (N_5727,N_715,N_2938);
or U5728 (N_5728,N_1972,N_1600);
nor U5729 (N_5729,N_1098,N_1540);
or U5730 (N_5730,N_458,N_67);
or U5731 (N_5731,N_942,N_337);
or U5732 (N_5732,N_304,N_493);
nand U5733 (N_5733,N_649,N_2196);
or U5734 (N_5734,N_1647,N_2225);
or U5735 (N_5735,N_3048,N_2966);
nor U5736 (N_5736,N_373,N_1492);
and U5737 (N_5737,N_2575,N_963);
xor U5738 (N_5738,N_1470,N_2471);
nand U5739 (N_5739,N_296,N_1809);
nor U5740 (N_5740,N_3003,N_1380);
or U5741 (N_5741,N_2657,N_2442);
nor U5742 (N_5742,N_1720,N_2592);
nor U5743 (N_5743,N_192,N_205);
or U5744 (N_5744,N_2410,N_121);
nor U5745 (N_5745,N_187,N_1395);
or U5746 (N_5746,N_1799,N_998);
nor U5747 (N_5747,N_1611,N_2593);
nor U5748 (N_5748,N_1202,N_2580);
nor U5749 (N_5749,N_1563,N_296);
xnor U5750 (N_5750,N_2181,N_837);
or U5751 (N_5751,N_143,N_2440);
or U5752 (N_5752,N_937,N_2465);
or U5753 (N_5753,N_401,N_1885);
nand U5754 (N_5754,N_2297,N_618);
nor U5755 (N_5755,N_1481,N_2139);
nand U5756 (N_5756,N_1621,N_2723);
nand U5757 (N_5757,N_1281,N_2778);
and U5758 (N_5758,N_1559,N_2316);
nor U5759 (N_5759,N_800,N_863);
nor U5760 (N_5760,N_107,N_1585);
or U5761 (N_5761,N_1027,N_2746);
or U5762 (N_5762,N_76,N_2134);
or U5763 (N_5763,N_2884,N_2328);
or U5764 (N_5764,N_294,N_789);
and U5765 (N_5765,N_1935,N_856);
and U5766 (N_5766,N_3013,N_363);
xor U5767 (N_5767,N_1498,N_2661);
nor U5768 (N_5768,N_1936,N_2993);
nand U5769 (N_5769,N_678,N_91);
nand U5770 (N_5770,N_328,N_2310);
or U5771 (N_5771,N_2472,N_2277);
and U5772 (N_5772,N_2648,N_1925);
nor U5773 (N_5773,N_2377,N_850);
or U5774 (N_5774,N_1710,N_866);
nand U5775 (N_5775,N_150,N_2062);
nand U5776 (N_5776,N_2443,N_809);
nand U5777 (N_5777,N_588,N_2831);
xor U5778 (N_5778,N_1220,N_1864);
nand U5779 (N_5779,N_2388,N_1952);
nor U5780 (N_5780,N_2377,N_520);
xor U5781 (N_5781,N_2012,N_2948);
or U5782 (N_5782,N_1103,N_2728);
or U5783 (N_5783,N_3040,N_182);
nand U5784 (N_5784,N_236,N_176);
xnor U5785 (N_5785,N_443,N_171);
nand U5786 (N_5786,N_324,N_2665);
and U5787 (N_5787,N_1888,N_1435);
nor U5788 (N_5788,N_3070,N_2554);
nand U5789 (N_5789,N_1504,N_1084);
xor U5790 (N_5790,N_1916,N_1998);
and U5791 (N_5791,N_2400,N_3085);
nand U5792 (N_5792,N_2283,N_428);
nand U5793 (N_5793,N_3087,N_1182);
or U5794 (N_5794,N_1356,N_1917);
nor U5795 (N_5795,N_1854,N_2125);
nor U5796 (N_5796,N_374,N_676);
nor U5797 (N_5797,N_1190,N_1010);
and U5798 (N_5798,N_2301,N_2879);
or U5799 (N_5799,N_784,N_632);
or U5800 (N_5800,N_1126,N_822);
nand U5801 (N_5801,N_1878,N_876);
nand U5802 (N_5802,N_3019,N_496);
xor U5803 (N_5803,N_67,N_39);
nand U5804 (N_5804,N_3101,N_2672);
and U5805 (N_5805,N_1222,N_1103);
or U5806 (N_5806,N_2149,N_2097);
nand U5807 (N_5807,N_448,N_1108);
nor U5808 (N_5808,N_689,N_1874);
and U5809 (N_5809,N_1841,N_405);
or U5810 (N_5810,N_1936,N_273);
nor U5811 (N_5811,N_711,N_2135);
and U5812 (N_5812,N_722,N_2490);
and U5813 (N_5813,N_2104,N_946);
xor U5814 (N_5814,N_1434,N_1419);
nand U5815 (N_5815,N_2508,N_913);
nand U5816 (N_5816,N_977,N_1304);
nor U5817 (N_5817,N_493,N_474);
and U5818 (N_5818,N_1624,N_2648);
xnor U5819 (N_5819,N_2308,N_1826);
nand U5820 (N_5820,N_197,N_3087);
nand U5821 (N_5821,N_840,N_576);
or U5822 (N_5822,N_2118,N_2124);
nand U5823 (N_5823,N_1796,N_1238);
nand U5824 (N_5824,N_1404,N_2816);
or U5825 (N_5825,N_1318,N_2832);
or U5826 (N_5826,N_1763,N_1303);
nor U5827 (N_5827,N_2227,N_1037);
and U5828 (N_5828,N_322,N_1857);
nand U5829 (N_5829,N_736,N_1636);
and U5830 (N_5830,N_2430,N_1871);
and U5831 (N_5831,N_620,N_204);
and U5832 (N_5832,N_1186,N_728);
xnor U5833 (N_5833,N_2902,N_1385);
nand U5834 (N_5834,N_3036,N_1099);
or U5835 (N_5835,N_3100,N_2621);
nor U5836 (N_5836,N_2377,N_2285);
or U5837 (N_5837,N_1598,N_3040);
nand U5838 (N_5838,N_2151,N_1898);
nand U5839 (N_5839,N_1323,N_2536);
nand U5840 (N_5840,N_1979,N_39);
xnor U5841 (N_5841,N_2084,N_2818);
nand U5842 (N_5842,N_638,N_1170);
and U5843 (N_5843,N_2186,N_1701);
xor U5844 (N_5844,N_1688,N_2457);
and U5845 (N_5845,N_149,N_2376);
nor U5846 (N_5846,N_1782,N_1695);
nor U5847 (N_5847,N_1078,N_2978);
or U5848 (N_5848,N_2942,N_566);
nand U5849 (N_5849,N_2469,N_503);
nand U5850 (N_5850,N_2463,N_41);
nor U5851 (N_5851,N_2549,N_725);
nand U5852 (N_5852,N_1060,N_546);
xor U5853 (N_5853,N_657,N_407);
nand U5854 (N_5854,N_2208,N_430);
or U5855 (N_5855,N_755,N_495);
nand U5856 (N_5856,N_859,N_1635);
and U5857 (N_5857,N_1682,N_2475);
or U5858 (N_5858,N_2948,N_694);
or U5859 (N_5859,N_2255,N_358);
and U5860 (N_5860,N_2381,N_2478);
or U5861 (N_5861,N_1976,N_1432);
nor U5862 (N_5862,N_916,N_2404);
and U5863 (N_5863,N_1010,N_2635);
xor U5864 (N_5864,N_491,N_2345);
nand U5865 (N_5865,N_2070,N_193);
nor U5866 (N_5866,N_2123,N_30);
nor U5867 (N_5867,N_1936,N_762);
or U5868 (N_5868,N_202,N_1126);
nor U5869 (N_5869,N_400,N_2882);
nand U5870 (N_5870,N_2805,N_1865);
and U5871 (N_5871,N_584,N_166);
or U5872 (N_5872,N_2715,N_1466);
nand U5873 (N_5873,N_170,N_2426);
nand U5874 (N_5874,N_1652,N_3093);
nor U5875 (N_5875,N_2173,N_988);
or U5876 (N_5876,N_2351,N_2525);
or U5877 (N_5877,N_747,N_651);
and U5878 (N_5878,N_928,N_800);
nand U5879 (N_5879,N_129,N_2993);
xor U5880 (N_5880,N_944,N_2979);
nand U5881 (N_5881,N_19,N_896);
or U5882 (N_5882,N_2355,N_686);
nand U5883 (N_5883,N_1571,N_670);
and U5884 (N_5884,N_913,N_572);
xnor U5885 (N_5885,N_2939,N_498);
and U5886 (N_5886,N_1239,N_2507);
and U5887 (N_5887,N_1204,N_248);
or U5888 (N_5888,N_1455,N_716);
nor U5889 (N_5889,N_80,N_454);
and U5890 (N_5890,N_419,N_2183);
and U5891 (N_5891,N_350,N_2021);
nor U5892 (N_5892,N_641,N_698);
nand U5893 (N_5893,N_34,N_2530);
or U5894 (N_5894,N_2016,N_209);
nor U5895 (N_5895,N_72,N_2786);
and U5896 (N_5896,N_2200,N_2141);
nand U5897 (N_5897,N_488,N_2400);
and U5898 (N_5898,N_2079,N_29);
nand U5899 (N_5899,N_1729,N_1993);
nand U5900 (N_5900,N_2940,N_2527);
and U5901 (N_5901,N_2153,N_1267);
and U5902 (N_5902,N_2576,N_3003);
nand U5903 (N_5903,N_402,N_1791);
or U5904 (N_5904,N_2677,N_2776);
xor U5905 (N_5905,N_30,N_865);
nand U5906 (N_5906,N_2700,N_922);
nand U5907 (N_5907,N_1527,N_1862);
or U5908 (N_5908,N_2626,N_611);
xor U5909 (N_5909,N_1581,N_2465);
nand U5910 (N_5910,N_471,N_2063);
and U5911 (N_5911,N_906,N_1677);
and U5912 (N_5912,N_1378,N_1566);
and U5913 (N_5913,N_595,N_2409);
and U5914 (N_5914,N_627,N_596);
or U5915 (N_5915,N_649,N_146);
or U5916 (N_5916,N_2544,N_2057);
nor U5917 (N_5917,N_3039,N_2646);
or U5918 (N_5918,N_1836,N_480);
xnor U5919 (N_5919,N_180,N_439);
or U5920 (N_5920,N_3063,N_1461);
and U5921 (N_5921,N_629,N_1909);
nor U5922 (N_5922,N_1481,N_2610);
xor U5923 (N_5923,N_836,N_521);
nor U5924 (N_5924,N_2037,N_1819);
nand U5925 (N_5925,N_59,N_111);
nor U5926 (N_5926,N_64,N_2357);
nand U5927 (N_5927,N_541,N_2150);
nor U5928 (N_5928,N_1385,N_332);
xor U5929 (N_5929,N_998,N_375);
or U5930 (N_5930,N_2936,N_1338);
and U5931 (N_5931,N_1407,N_902);
and U5932 (N_5932,N_2280,N_1049);
nor U5933 (N_5933,N_1834,N_1204);
nand U5934 (N_5934,N_1103,N_591);
or U5935 (N_5935,N_1000,N_376);
nand U5936 (N_5936,N_1575,N_2234);
nand U5937 (N_5937,N_2470,N_2029);
xnor U5938 (N_5938,N_780,N_1067);
and U5939 (N_5939,N_1899,N_2671);
and U5940 (N_5940,N_2546,N_1412);
and U5941 (N_5941,N_280,N_1738);
and U5942 (N_5942,N_2950,N_433);
nand U5943 (N_5943,N_2241,N_183);
and U5944 (N_5944,N_2760,N_1035);
and U5945 (N_5945,N_1329,N_699);
and U5946 (N_5946,N_1341,N_2709);
nand U5947 (N_5947,N_3000,N_1445);
nor U5948 (N_5948,N_210,N_1663);
and U5949 (N_5949,N_1851,N_1342);
nor U5950 (N_5950,N_2498,N_1714);
xnor U5951 (N_5951,N_533,N_317);
or U5952 (N_5952,N_409,N_1591);
and U5953 (N_5953,N_3071,N_953);
nor U5954 (N_5954,N_1032,N_2492);
and U5955 (N_5955,N_142,N_1571);
or U5956 (N_5956,N_2576,N_1740);
nand U5957 (N_5957,N_2142,N_2991);
and U5958 (N_5958,N_863,N_1229);
nand U5959 (N_5959,N_881,N_318);
or U5960 (N_5960,N_2820,N_1095);
or U5961 (N_5961,N_2238,N_352);
nor U5962 (N_5962,N_689,N_293);
nand U5963 (N_5963,N_1535,N_732);
or U5964 (N_5964,N_2685,N_2199);
nand U5965 (N_5965,N_503,N_555);
nand U5966 (N_5966,N_2107,N_3041);
nor U5967 (N_5967,N_1345,N_2060);
or U5968 (N_5968,N_978,N_2528);
nor U5969 (N_5969,N_2886,N_1900);
xor U5970 (N_5970,N_2751,N_787);
nor U5971 (N_5971,N_1476,N_371);
xnor U5972 (N_5972,N_2393,N_2653);
nand U5973 (N_5973,N_784,N_1009);
and U5974 (N_5974,N_1655,N_2330);
nand U5975 (N_5975,N_2828,N_2462);
nor U5976 (N_5976,N_1236,N_1180);
or U5977 (N_5977,N_2898,N_872);
nand U5978 (N_5978,N_2069,N_1264);
and U5979 (N_5979,N_1955,N_3041);
nand U5980 (N_5980,N_1934,N_1032);
or U5981 (N_5981,N_1225,N_1070);
and U5982 (N_5982,N_2855,N_123);
nand U5983 (N_5983,N_1219,N_1377);
nand U5984 (N_5984,N_2725,N_2056);
nand U5985 (N_5985,N_1475,N_1679);
nor U5986 (N_5986,N_111,N_454);
or U5987 (N_5987,N_828,N_1243);
nor U5988 (N_5988,N_2202,N_2644);
and U5989 (N_5989,N_309,N_799);
nor U5990 (N_5990,N_1125,N_1230);
xor U5991 (N_5991,N_396,N_1611);
xor U5992 (N_5992,N_2944,N_2412);
or U5993 (N_5993,N_2714,N_2516);
and U5994 (N_5994,N_1785,N_550);
xor U5995 (N_5995,N_2230,N_844);
or U5996 (N_5996,N_1855,N_1189);
nor U5997 (N_5997,N_2968,N_2941);
xnor U5998 (N_5998,N_9,N_2116);
or U5999 (N_5999,N_1925,N_558);
or U6000 (N_6000,N_2204,N_666);
or U6001 (N_6001,N_741,N_2004);
nand U6002 (N_6002,N_587,N_603);
nor U6003 (N_6003,N_1153,N_2350);
xor U6004 (N_6004,N_1988,N_31);
or U6005 (N_6005,N_3006,N_2848);
xnor U6006 (N_6006,N_1862,N_2000);
and U6007 (N_6007,N_1721,N_270);
or U6008 (N_6008,N_819,N_555);
and U6009 (N_6009,N_715,N_1876);
nand U6010 (N_6010,N_2840,N_417);
nand U6011 (N_6011,N_700,N_2400);
nor U6012 (N_6012,N_2964,N_1788);
or U6013 (N_6013,N_1837,N_1472);
xnor U6014 (N_6014,N_1638,N_272);
and U6015 (N_6015,N_660,N_1319);
nand U6016 (N_6016,N_306,N_2397);
nor U6017 (N_6017,N_2068,N_1032);
nand U6018 (N_6018,N_1786,N_1624);
nand U6019 (N_6019,N_501,N_689);
nor U6020 (N_6020,N_1240,N_2805);
nor U6021 (N_6021,N_1923,N_1944);
nor U6022 (N_6022,N_1343,N_2334);
nor U6023 (N_6023,N_1780,N_823);
xnor U6024 (N_6024,N_645,N_1467);
and U6025 (N_6025,N_3123,N_1509);
nor U6026 (N_6026,N_1665,N_602);
nand U6027 (N_6027,N_685,N_1418);
or U6028 (N_6028,N_1292,N_1006);
or U6029 (N_6029,N_2309,N_2634);
or U6030 (N_6030,N_1892,N_622);
nor U6031 (N_6031,N_145,N_2983);
nor U6032 (N_6032,N_1337,N_2911);
or U6033 (N_6033,N_2613,N_2244);
or U6034 (N_6034,N_1662,N_1785);
or U6035 (N_6035,N_1993,N_336);
or U6036 (N_6036,N_3020,N_9);
or U6037 (N_6037,N_93,N_918);
xor U6038 (N_6038,N_1751,N_1049);
and U6039 (N_6039,N_2388,N_743);
and U6040 (N_6040,N_2648,N_1382);
or U6041 (N_6041,N_982,N_2624);
nor U6042 (N_6042,N_1363,N_1459);
nor U6043 (N_6043,N_2584,N_2708);
nand U6044 (N_6044,N_3054,N_2787);
nand U6045 (N_6045,N_2718,N_987);
or U6046 (N_6046,N_3086,N_1384);
nand U6047 (N_6047,N_1941,N_2909);
or U6048 (N_6048,N_1118,N_1591);
xor U6049 (N_6049,N_751,N_371);
nand U6050 (N_6050,N_23,N_2074);
nand U6051 (N_6051,N_2269,N_2488);
or U6052 (N_6052,N_3077,N_2448);
and U6053 (N_6053,N_1644,N_2493);
nand U6054 (N_6054,N_1028,N_2735);
and U6055 (N_6055,N_1961,N_2644);
nor U6056 (N_6056,N_267,N_302);
nand U6057 (N_6057,N_1564,N_1004);
and U6058 (N_6058,N_159,N_2421);
or U6059 (N_6059,N_775,N_93);
and U6060 (N_6060,N_2076,N_2393);
xnor U6061 (N_6061,N_2607,N_1966);
and U6062 (N_6062,N_282,N_2313);
nand U6063 (N_6063,N_777,N_1271);
and U6064 (N_6064,N_2508,N_667);
nor U6065 (N_6065,N_999,N_2980);
xor U6066 (N_6066,N_2474,N_2568);
nand U6067 (N_6067,N_964,N_978);
nor U6068 (N_6068,N_282,N_976);
and U6069 (N_6069,N_2111,N_1444);
or U6070 (N_6070,N_1083,N_2605);
nand U6071 (N_6071,N_2256,N_1264);
or U6072 (N_6072,N_1120,N_2294);
nand U6073 (N_6073,N_652,N_1030);
and U6074 (N_6074,N_438,N_2276);
nor U6075 (N_6075,N_266,N_445);
nand U6076 (N_6076,N_1581,N_1766);
or U6077 (N_6077,N_776,N_1863);
or U6078 (N_6078,N_1348,N_1157);
nand U6079 (N_6079,N_2071,N_2788);
and U6080 (N_6080,N_2416,N_1577);
or U6081 (N_6081,N_2166,N_1894);
xnor U6082 (N_6082,N_821,N_1925);
and U6083 (N_6083,N_2526,N_2358);
nand U6084 (N_6084,N_473,N_318);
or U6085 (N_6085,N_4,N_987);
or U6086 (N_6086,N_1705,N_2675);
nor U6087 (N_6087,N_2604,N_533);
xor U6088 (N_6088,N_440,N_1462);
and U6089 (N_6089,N_2058,N_2121);
nor U6090 (N_6090,N_221,N_1399);
nand U6091 (N_6091,N_2055,N_2683);
nor U6092 (N_6092,N_1985,N_1907);
nor U6093 (N_6093,N_1494,N_1059);
nand U6094 (N_6094,N_2035,N_1739);
or U6095 (N_6095,N_956,N_3020);
or U6096 (N_6096,N_642,N_2829);
nand U6097 (N_6097,N_3084,N_1317);
nor U6098 (N_6098,N_2757,N_3117);
xor U6099 (N_6099,N_1913,N_267);
or U6100 (N_6100,N_1331,N_1632);
nand U6101 (N_6101,N_1393,N_2899);
xnor U6102 (N_6102,N_1971,N_2957);
or U6103 (N_6103,N_2361,N_3073);
xor U6104 (N_6104,N_1477,N_718);
and U6105 (N_6105,N_2621,N_1757);
nand U6106 (N_6106,N_805,N_1980);
nor U6107 (N_6107,N_1995,N_1511);
and U6108 (N_6108,N_1482,N_2517);
nor U6109 (N_6109,N_2292,N_86);
nor U6110 (N_6110,N_2148,N_1592);
nor U6111 (N_6111,N_2531,N_1579);
nand U6112 (N_6112,N_350,N_2640);
nand U6113 (N_6113,N_1306,N_76);
xor U6114 (N_6114,N_2663,N_932);
nor U6115 (N_6115,N_678,N_3062);
xor U6116 (N_6116,N_582,N_650);
nor U6117 (N_6117,N_994,N_2587);
and U6118 (N_6118,N_2319,N_1641);
or U6119 (N_6119,N_2724,N_605);
nor U6120 (N_6120,N_1860,N_356);
or U6121 (N_6121,N_2761,N_437);
or U6122 (N_6122,N_1273,N_1630);
nand U6123 (N_6123,N_2241,N_2709);
nor U6124 (N_6124,N_981,N_2565);
nor U6125 (N_6125,N_1980,N_2895);
nand U6126 (N_6126,N_740,N_1230);
nand U6127 (N_6127,N_1636,N_546);
or U6128 (N_6128,N_1280,N_1022);
nor U6129 (N_6129,N_1488,N_1113);
or U6130 (N_6130,N_2314,N_2577);
nand U6131 (N_6131,N_3008,N_2271);
nand U6132 (N_6132,N_1557,N_1188);
or U6133 (N_6133,N_2171,N_2981);
or U6134 (N_6134,N_1425,N_1540);
and U6135 (N_6135,N_649,N_621);
and U6136 (N_6136,N_1444,N_1699);
nor U6137 (N_6137,N_1051,N_2732);
nand U6138 (N_6138,N_2827,N_906);
or U6139 (N_6139,N_2172,N_2914);
and U6140 (N_6140,N_1529,N_2517);
nand U6141 (N_6141,N_842,N_1649);
and U6142 (N_6142,N_31,N_2032);
and U6143 (N_6143,N_805,N_2622);
and U6144 (N_6144,N_32,N_2859);
and U6145 (N_6145,N_2060,N_292);
nor U6146 (N_6146,N_2469,N_40);
nand U6147 (N_6147,N_1851,N_2512);
or U6148 (N_6148,N_3030,N_202);
nand U6149 (N_6149,N_2291,N_1200);
nor U6150 (N_6150,N_223,N_953);
or U6151 (N_6151,N_2672,N_128);
nand U6152 (N_6152,N_2157,N_281);
and U6153 (N_6153,N_2830,N_455);
nor U6154 (N_6154,N_525,N_2248);
nor U6155 (N_6155,N_1612,N_2939);
or U6156 (N_6156,N_2101,N_2552);
nand U6157 (N_6157,N_691,N_995);
or U6158 (N_6158,N_1962,N_448);
nor U6159 (N_6159,N_2054,N_1334);
nand U6160 (N_6160,N_30,N_1124);
nor U6161 (N_6161,N_2783,N_41);
or U6162 (N_6162,N_2644,N_2822);
nand U6163 (N_6163,N_718,N_1643);
nor U6164 (N_6164,N_2730,N_2127);
nand U6165 (N_6165,N_2232,N_3068);
nand U6166 (N_6166,N_2527,N_1353);
and U6167 (N_6167,N_951,N_515);
and U6168 (N_6168,N_67,N_2805);
nand U6169 (N_6169,N_782,N_2058);
nor U6170 (N_6170,N_897,N_579);
and U6171 (N_6171,N_2791,N_239);
and U6172 (N_6172,N_1472,N_764);
and U6173 (N_6173,N_116,N_1783);
or U6174 (N_6174,N_339,N_73);
nor U6175 (N_6175,N_200,N_149);
or U6176 (N_6176,N_2687,N_216);
nand U6177 (N_6177,N_296,N_548);
or U6178 (N_6178,N_110,N_1367);
and U6179 (N_6179,N_917,N_1018);
nor U6180 (N_6180,N_2306,N_1268);
or U6181 (N_6181,N_1436,N_2650);
nor U6182 (N_6182,N_1990,N_2222);
or U6183 (N_6183,N_1532,N_2643);
nor U6184 (N_6184,N_1004,N_714);
nand U6185 (N_6185,N_2870,N_1147);
or U6186 (N_6186,N_2864,N_2061);
xor U6187 (N_6187,N_1746,N_1191);
xnor U6188 (N_6188,N_230,N_3028);
and U6189 (N_6189,N_1189,N_999);
or U6190 (N_6190,N_449,N_2559);
or U6191 (N_6191,N_3028,N_2350);
and U6192 (N_6192,N_747,N_2198);
nor U6193 (N_6193,N_2216,N_2417);
or U6194 (N_6194,N_2068,N_669);
and U6195 (N_6195,N_2543,N_963);
or U6196 (N_6196,N_840,N_1627);
and U6197 (N_6197,N_1671,N_1452);
nor U6198 (N_6198,N_2903,N_2006);
nand U6199 (N_6199,N_577,N_1226);
and U6200 (N_6200,N_1329,N_918);
nand U6201 (N_6201,N_2568,N_56);
nor U6202 (N_6202,N_1895,N_2944);
nand U6203 (N_6203,N_1332,N_1813);
and U6204 (N_6204,N_2919,N_2342);
and U6205 (N_6205,N_1317,N_1726);
nor U6206 (N_6206,N_1514,N_1945);
nor U6207 (N_6207,N_2506,N_3016);
and U6208 (N_6208,N_2038,N_217);
and U6209 (N_6209,N_1148,N_1151);
nand U6210 (N_6210,N_754,N_2366);
or U6211 (N_6211,N_2132,N_2058);
nand U6212 (N_6212,N_1096,N_55);
nor U6213 (N_6213,N_2971,N_2083);
and U6214 (N_6214,N_827,N_171);
and U6215 (N_6215,N_1465,N_2217);
nand U6216 (N_6216,N_2034,N_824);
xor U6217 (N_6217,N_640,N_149);
or U6218 (N_6218,N_2668,N_525);
or U6219 (N_6219,N_2382,N_674);
or U6220 (N_6220,N_2523,N_2169);
or U6221 (N_6221,N_33,N_1736);
and U6222 (N_6222,N_2928,N_1768);
or U6223 (N_6223,N_2876,N_1383);
and U6224 (N_6224,N_2828,N_2713);
nor U6225 (N_6225,N_2544,N_145);
nor U6226 (N_6226,N_1572,N_1410);
or U6227 (N_6227,N_2674,N_2485);
and U6228 (N_6228,N_2746,N_2802);
and U6229 (N_6229,N_410,N_2129);
nand U6230 (N_6230,N_2921,N_365);
nand U6231 (N_6231,N_421,N_2005);
xnor U6232 (N_6232,N_1711,N_167);
and U6233 (N_6233,N_2893,N_2627);
nand U6234 (N_6234,N_3060,N_1084);
nor U6235 (N_6235,N_2118,N_1156);
and U6236 (N_6236,N_2681,N_435);
or U6237 (N_6237,N_121,N_979);
or U6238 (N_6238,N_1420,N_1756);
or U6239 (N_6239,N_1080,N_501);
or U6240 (N_6240,N_1991,N_2607);
nor U6241 (N_6241,N_1465,N_1976);
nand U6242 (N_6242,N_153,N_2171);
nand U6243 (N_6243,N_2640,N_1707);
nor U6244 (N_6244,N_1299,N_2207);
nand U6245 (N_6245,N_333,N_671);
nor U6246 (N_6246,N_2590,N_2143);
and U6247 (N_6247,N_598,N_463);
nor U6248 (N_6248,N_2142,N_1003);
or U6249 (N_6249,N_2647,N_3058);
and U6250 (N_6250,N_5895,N_5613);
xnor U6251 (N_6251,N_3854,N_5162);
and U6252 (N_6252,N_4426,N_4780);
xor U6253 (N_6253,N_5754,N_6016);
or U6254 (N_6254,N_4465,N_5972);
xnor U6255 (N_6255,N_5844,N_3614);
or U6256 (N_6256,N_4427,N_4071);
nor U6257 (N_6257,N_4958,N_5473);
or U6258 (N_6258,N_4587,N_3129);
xnor U6259 (N_6259,N_3197,N_5615);
nor U6260 (N_6260,N_4415,N_3472);
xnor U6261 (N_6261,N_4080,N_5370);
nor U6262 (N_6262,N_4586,N_3592);
nor U6263 (N_6263,N_5287,N_4572);
or U6264 (N_6264,N_6071,N_4581);
or U6265 (N_6265,N_3330,N_5267);
nor U6266 (N_6266,N_5746,N_5147);
nand U6267 (N_6267,N_6115,N_3756);
and U6268 (N_6268,N_4807,N_3530);
nand U6269 (N_6269,N_6130,N_6001);
and U6270 (N_6270,N_3236,N_3545);
and U6271 (N_6271,N_4687,N_3193);
nor U6272 (N_6272,N_3218,N_5246);
xnor U6273 (N_6273,N_3337,N_5708);
or U6274 (N_6274,N_4842,N_5783);
and U6275 (N_6275,N_3148,N_3204);
and U6276 (N_6276,N_4795,N_4939);
and U6277 (N_6277,N_3712,N_6148);
and U6278 (N_6278,N_5335,N_4299);
and U6279 (N_6279,N_5309,N_5956);
nor U6280 (N_6280,N_4075,N_3512);
or U6281 (N_6281,N_3251,N_4079);
xnor U6282 (N_6282,N_4001,N_3223);
nor U6283 (N_6283,N_5367,N_4830);
and U6284 (N_6284,N_6210,N_5118);
xnor U6285 (N_6285,N_5351,N_4508);
and U6286 (N_6286,N_4014,N_3136);
and U6287 (N_6287,N_4648,N_4083);
nand U6288 (N_6288,N_5554,N_4536);
nand U6289 (N_6289,N_3893,N_6010);
nor U6290 (N_6290,N_5279,N_5823);
and U6291 (N_6291,N_3369,N_3438);
nor U6292 (N_6292,N_3906,N_3620);
nor U6293 (N_6293,N_5283,N_5440);
nand U6294 (N_6294,N_3582,N_3532);
nand U6295 (N_6295,N_3149,N_4015);
and U6296 (N_6296,N_5769,N_4091);
nand U6297 (N_6297,N_4607,N_5148);
or U6298 (N_6298,N_3836,N_3789);
nand U6299 (N_6299,N_6077,N_5639);
nand U6300 (N_6300,N_4247,N_4023);
nor U6301 (N_6301,N_3486,N_3367);
or U6302 (N_6302,N_3672,N_5560);
nor U6303 (N_6303,N_3824,N_5621);
nor U6304 (N_6304,N_3467,N_3831);
or U6305 (N_6305,N_5740,N_5994);
and U6306 (N_6306,N_4667,N_5978);
nand U6307 (N_6307,N_5976,N_4906);
xor U6308 (N_6308,N_5127,N_5145);
xor U6309 (N_6309,N_4834,N_4959);
and U6310 (N_6310,N_3520,N_5350);
nand U6311 (N_6311,N_4783,N_6093);
or U6312 (N_6312,N_5141,N_6226);
nor U6313 (N_6313,N_4757,N_3606);
and U6314 (N_6314,N_5561,N_4522);
nor U6315 (N_6315,N_6134,N_5571);
or U6316 (N_6316,N_5327,N_5591);
or U6317 (N_6317,N_5944,N_4353);
nor U6318 (N_6318,N_5810,N_5132);
nand U6319 (N_6319,N_4511,N_3380);
nand U6320 (N_6320,N_6132,N_3813);
nand U6321 (N_6321,N_4175,N_6243);
or U6322 (N_6322,N_4211,N_3817);
or U6323 (N_6323,N_5097,N_3418);
nand U6324 (N_6324,N_5464,N_3869);
or U6325 (N_6325,N_3918,N_4407);
nor U6326 (N_6326,N_3144,N_3923);
and U6327 (N_6327,N_4631,N_5871);
or U6328 (N_6328,N_5930,N_3498);
nand U6329 (N_6329,N_4525,N_3793);
nor U6330 (N_6330,N_3776,N_5306);
nor U6331 (N_6331,N_4770,N_5451);
and U6332 (N_6332,N_5973,N_3795);
nand U6333 (N_6333,N_3377,N_3877);
and U6334 (N_6334,N_4466,N_3777);
nand U6335 (N_6335,N_6179,N_5641);
nand U6336 (N_6336,N_6221,N_3888);
nor U6337 (N_6337,N_4389,N_3782);
and U6338 (N_6338,N_4403,N_4258);
xor U6339 (N_6339,N_4868,N_3503);
or U6340 (N_6340,N_3480,N_3977);
or U6341 (N_6341,N_5414,N_5939);
nand U6342 (N_6342,N_4775,N_3714);
xor U6343 (N_6343,N_4866,N_4285);
nand U6344 (N_6344,N_5429,N_5940);
nor U6345 (N_6345,N_5355,N_4026);
nand U6346 (N_6346,N_3842,N_5899);
or U6347 (N_6347,N_3573,N_4222);
and U6348 (N_6348,N_5847,N_5670);
nor U6349 (N_6349,N_5483,N_3415);
or U6350 (N_6350,N_5077,N_5732);
nand U6351 (N_6351,N_5159,N_3551);
and U6352 (N_6352,N_3708,N_5504);
nor U6353 (N_6353,N_5648,N_3334);
nor U6354 (N_6354,N_3692,N_3682);
nor U6355 (N_6355,N_5597,N_4309);
and U6356 (N_6356,N_5062,N_3343);
nor U6357 (N_6357,N_5912,N_3170);
or U6358 (N_6358,N_4902,N_5197);
and U6359 (N_6359,N_4641,N_3293);
xnor U6360 (N_6360,N_5137,N_5675);
or U6361 (N_6361,N_4887,N_3505);
nand U6362 (N_6362,N_4929,N_3417);
xnor U6363 (N_6363,N_3132,N_5253);
nand U6364 (N_6364,N_5034,N_4460);
nand U6365 (N_6365,N_3636,N_4908);
nor U6366 (N_6366,N_5991,N_5623);
and U6367 (N_6367,N_5175,N_5138);
and U6368 (N_6368,N_5153,N_4762);
and U6369 (N_6369,N_3931,N_3666);
or U6370 (N_6370,N_4187,N_3612);
nand U6371 (N_6371,N_5004,N_5723);
nor U6372 (N_6372,N_3523,N_4148);
or U6373 (N_6373,N_4010,N_5467);
xor U6374 (N_6374,N_3419,N_4094);
or U6375 (N_6375,N_5381,N_4092);
nor U6376 (N_6376,N_4051,N_4978);
and U6377 (N_6377,N_3837,N_3641);
nand U6378 (N_6378,N_4322,N_4604);
or U6379 (N_6379,N_4159,N_5241);
and U6380 (N_6380,N_5432,N_3262);
and U6381 (N_6381,N_3483,N_4737);
nor U6382 (N_6382,N_4438,N_3348);
nor U6383 (N_6383,N_5953,N_5509);
or U6384 (N_6384,N_5502,N_4000);
nor U6385 (N_6385,N_4447,N_4590);
and U6386 (N_6386,N_4449,N_5987);
nor U6387 (N_6387,N_3389,N_5803);
nor U6388 (N_6388,N_5498,N_5662);
nand U6389 (N_6389,N_6100,N_5119);
and U6390 (N_6390,N_5386,N_6089);
and U6391 (N_6391,N_4044,N_4541);
nor U6392 (N_6392,N_3455,N_5977);
nand U6393 (N_6393,N_6006,N_3166);
nor U6394 (N_6394,N_3312,N_4067);
xnor U6395 (N_6395,N_3300,N_3731);
xnor U6396 (N_6396,N_5934,N_3858);
or U6397 (N_6397,N_3282,N_5424);
nor U6398 (N_6398,N_5182,N_5308);
and U6399 (N_6399,N_4356,N_5219);
and U6400 (N_6400,N_3651,N_5113);
nor U6401 (N_6401,N_3420,N_5096);
nor U6402 (N_6402,N_5861,N_4411);
and U6403 (N_6403,N_3368,N_4251);
or U6404 (N_6404,N_3657,N_5820);
or U6405 (N_6405,N_5385,N_6163);
nor U6406 (N_6406,N_3536,N_3159);
or U6407 (N_6407,N_5838,N_4919);
and U6408 (N_6408,N_6178,N_4702);
nand U6409 (N_6409,N_5851,N_4021);
or U6410 (N_6410,N_5954,N_5457);
or U6411 (N_6411,N_5776,N_4200);
or U6412 (N_6412,N_3517,N_4747);
nor U6413 (N_6413,N_5550,N_4492);
xnor U6414 (N_6414,N_4953,N_6246);
nor U6415 (N_6415,N_3879,N_5100);
nor U6416 (N_6416,N_6156,N_5718);
nor U6417 (N_6417,N_4905,N_3960);
nand U6418 (N_6418,N_5378,N_4995);
nor U6419 (N_6419,N_3240,N_3679);
nor U6420 (N_6420,N_4417,N_3173);
nand U6421 (N_6421,N_4333,N_6052);
and U6422 (N_6422,N_5179,N_3386);
and U6423 (N_6423,N_6000,N_4265);
and U6424 (N_6424,N_5555,N_5734);
nor U6425 (N_6425,N_3162,N_4570);
xnor U6426 (N_6426,N_5110,N_5074);
and U6427 (N_6427,N_5379,N_3919);
and U6428 (N_6428,N_3724,N_4582);
nor U6429 (N_6429,N_3260,N_4442);
nand U6430 (N_6430,N_5023,N_4549);
nand U6431 (N_6431,N_6005,N_5111);
xor U6432 (N_6432,N_4217,N_4206);
nand U6433 (N_6433,N_4085,N_3371);
nand U6434 (N_6434,N_3451,N_4608);
nand U6435 (N_6435,N_5095,N_5729);
or U6436 (N_6436,N_5411,N_4367);
and U6437 (N_6437,N_3489,N_3809);
nor U6438 (N_6438,N_5345,N_4530);
or U6439 (N_6439,N_4170,N_4833);
nor U6440 (N_6440,N_3957,N_6167);
and U6441 (N_6441,N_3221,N_6114);
nor U6442 (N_6442,N_5731,N_5966);
nand U6443 (N_6443,N_4524,N_4630);
or U6444 (N_6444,N_5501,N_4329);
nor U6445 (N_6445,N_4618,N_6020);
xnor U6446 (N_6446,N_5547,N_3655);
nor U6447 (N_6447,N_3151,N_4991);
and U6448 (N_6448,N_6161,N_5448);
or U6449 (N_6449,N_5207,N_5985);
nor U6450 (N_6450,N_3432,N_3212);
nor U6451 (N_6451,N_5750,N_4501);
or U6452 (N_6452,N_6224,N_5573);
xnor U6453 (N_6453,N_4538,N_3669);
nand U6454 (N_6454,N_3921,N_5115);
nand U6455 (N_6455,N_3865,N_3492);
and U6456 (N_6456,N_6090,N_3794);
nor U6457 (N_6457,N_5316,N_4794);
and U6458 (N_6458,N_6108,N_3456);
nand U6459 (N_6459,N_3328,N_5812);
or U6460 (N_6460,N_4443,N_5923);
xnor U6461 (N_6461,N_5051,N_5666);
xor U6462 (N_6462,N_3988,N_4095);
and U6463 (N_6463,N_5181,N_5172);
and U6464 (N_6464,N_5202,N_3909);
or U6465 (N_6465,N_4102,N_4601);
or U6466 (N_6466,N_3764,N_4700);
xnor U6467 (N_6467,N_3576,N_4310);
or U6468 (N_6468,N_3289,N_3891);
and U6469 (N_6469,N_4678,N_5060);
or U6470 (N_6470,N_3501,N_3822);
and U6471 (N_6471,N_6080,N_3321);
and U6472 (N_6472,N_3588,N_5231);
or U6473 (N_6473,N_4968,N_5523);
nor U6474 (N_6474,N_3617,N_3754);
nor U6475 (N_6475,N_6086,N_4394);
nand U6476 (N_6476,N_3514,N_5905);
or U6477 (N_6477,N_5960,N_6061);
and U6478 (N_6478,N_3786,N_4126);
nor U6479 (N_6479,N_4393,N_3447);
or U6480 (N_6480,N_6133,N_4861);
or U6481 (N_6481,N_5427,N_3521);
and U6482 (N_6482,N_3336,N_3359);
nand U6483 (N_6483,N_3541,N_4617);
nor U6484 (N_6484,N_3583,N_3339);
nand U6485 (N_6485,N_5507,N_3340);
or U6486 (N_6486,N_4584,N_5099);
and U6487 (N_6487,N_5273,N_5790);
nor U6488 (N_6488,N_3751,N_3962);
nor U6489 (N_6489,N_5961,N_5490);
nand U6490 (N_6490,N_5192,N_6007);
or U6491 (N_6491,N_5849,N_4613);
or U6492 (N_6492,N_3202,N_3543);
xor U6493 (N_6493,N_3375,N_4204);
and U6494 (N_6494,N_5070,N_4857);
and U6495 (N_6495,N_5101,N_4396);
xnor U6496 (N_6496,N_5418,N_3353);
and U6497 (N_6497,N_5698,N_3812);
nand U6498 (N_6498,N_3981,N_3140);
nand U6499 (N_6499,N_4926,N_4802);
nand U6500 (N_6500,N_3237,N_5947);
and U6501 (N_6501,N_5016,N_4994);
or U6502 (N_6502,N_6117,N_5518);
xnor U6503 (N_6503,N_3430,N_4977);
xnor U6504 (N_6504,N_5008,N_5938);
and U6505 (N_6505,N_4063,N_5056);
or U6506 (N_6506,N_4632,N_5488);
and U6507 (N_6507,N_4798,N_5319);
nor U6508 (N_6508,N_4328,N_4138);
nand U6509 (N_6509,N_4829,N_3933);
or U6510 (N_6510,N_6015,N_5980);
xnor U6511 (N_6511,N_3621,N_4897);
nand U6512 (N_6512,N_4342,N_5860);
and U6513 (N_6513,N_3147,N_6162);
nand U6514 (N_6514,N_5330,N_5830);
nor U6515 (N_6515,N_5800,N_5697);
or U6516 (N_6516,N_4357,N_5404);
nor U6517 (N_6517,N_6004,N_5284);
xnor U6518 (N_6518,N_4409,N_5767);
nor U6519 (N_6519,N_6073,N_3579);
or U6520 (N_6520,N_4379,N_4941);
nor U6521 (N_6521,N_4171,N_5701);
and U6522 (N_6522,N_3407,N_3454);
nand U6523 (N_6523,N_5336,N_5049);
nand U6524 (N_6524,N_5924,N_4433);
or U6525 (N_6525,N_5757,N_5638);
and U6526 (N_6526,N_4735,N_6088);
nand U6527 (N_6527,N_3769,N_4354);
and U6528 (N_6528,N_4655,N_4042);
nor U6529 (N_6529,N_5684,N_6081);
and U6530 (N_6530,N_5726,N_4891);
nor U6531 (N_6531,N_4679,N_3287);
and U6532 (N_6532,N_6023,N_5581);
or U6533 (N_6533,N_4163,N_4803);
nor U6534 (N_6534,N_4877,N_5904);
nor U6535 (N_6535,N_6039,N_6025);
nor U6536 (N_6536,N_3832,N_5126);
nand U6537 (N_6537,N_5538,N_5317);
or U6538 (N_6538,N_3230,N_5039);
nor U6539 (N_6539,N_4903,N_5018);
nand U6540 (N_6540,N_4568,N_5017);
nand U6541 (N_6541,N_4615,N_3280);
or U6542 (N_6542,N_4535,N_4585);
or U6543 (N_6543,N_5075,N_3649);
or U6544 (N_6544,N_5146,N_4351);
nor U6545 (N_6545,N_3327,N_3125);
or U6546 (N_6546,N_4104,N_5109);
and U6547 (N_6547,N_6013,N_3687);
xnor U6548 (N_6548,N_5294,N_4490);
and U6549 (N_6549,N_4985,N_4796);
or U6550 (N_6550,N_4889,N_5530);
nand U6551 (N_6551,N_5624,N_6024);
nand U6552 (N_6552,N_3799,N_3458);
nand U6553 (N_6553,N_3453,N_3137);
or U6554 (N_6554,N_4793,N_4745);
nand U6555 (N_6555,N_4653,N_5704);
xor U6556 (N_6556,N_3803,N_5710);
nand U6557 (N_6557,N_3944,N_3587);
nand U6558 (N_6558,N_4167,N_4753);
or U6559 (N_6559,N_3405,N_6155);
and U6560 (N_6560,N_4338,N_4963);
and U6561 (N_6561,N_3966,N_4516);
nand U6562 (N_6562,N_5974,N_3976);
or U6563 (N_6563,N_5751,N_5644);
nand U6564 (N_6564,N_5686,N_5721);
xor U6565 (N_6565,N_4927,N_6153);
nand U6566 (N_6566,N_3780,N_3727);
or U6567 (N_6567,N_3935,N_4886);
or U6568 (N_6568,N_4223,N_4786);
and U6569 (N_6569,N_4970,N_3356);
nor U6570 (N_6570,N_4061,N_5030);
and U6571 (N_6571,N_4589,N_6201);
nand U6572 (N_6572,N_4477,N_5280);
and U6573 (N_6573,N_5873,N_3266);
nor U6574 (N_6574,N_3537,N_3134);
nor U6575 (N_6575,N_3802,N_4418);
or U6576 (N_6576,N_5220,N_4890);
or U6577 (N_6577,N_4312,N_5787);
or U6578 (N_6578,N_3248,N_3693);
xor U6579 (N_6579,N_3730,N_6174);
or U6580 (N_6580,N_5481,N_5897);
nand U6581 (N_6581,N_4129,N_4773);
or U6582 (N_6582,N_3992,N_5695);
nor U6583 (N_6583,N_4909,N_3235);
or U6584 (N_6584,N_3568,N_4243);
nand U6585 (N_6585,N_5116,N_4575);
nand U6586 (N_6586,N_3247,N_4716);
nor U6587 (N_6587,N_4514,N_5982);
or U6588 (N_6588,N_3391,N_4298);
and U6589 (N_6589,N_5163,N_4883);
nor U6590 (N_6590,N_4343,N_4387);
or U6591 (N_6591,N_3850,N_5532);
nand U6592 (N_6592,N_3395,N_3535);
xor U6593 (N_6593,N_5065,N_6094);
or U6594 (N_6594,N_4936,N_4157);
xor U6595 (N_6595,N_4565,N_3787);
or U6596 (N_6596,N_5853,N_3862);
and U6597 (N_6597,N_3884,N_3961);
nor U6598 (N_6598,N_4341,N_5443);
or U6599 (N_6599,N_5664,N_5785);
and U6600 (N_6600,N_5368,N_3413);
and U6601 (N_6601,N_4376,N_4278);
and U6602 (N_6602,N_6107,N_5323);
xor U6603 (N_6603,N_3883,N_4419);
nand U6604 (N_6604,N_5239,N_3770);
or U6605 (N_6605,N_5862,N_3181);
nand U6606 (N_6606,N_4593,N_4184);
nor U6607 (N_6607,N_5161,N_3878);
nor U6608 (N_6608,N_3733,N_5134);
nand U6609 (N_6609,N_4268,N_6050);
and U6610 (N_6610,N_5681,N_5625);
nor U6611 (N_6611,N_5349,N_5212);
nand U6612 (N_6612,N_4365,N_4112);
and U6613 (N_6613,N_4253,N_3557);
or U6614 (N_6614,N_5626,N_3875);
and U6615 (N_6615,N_3737,N_6208);
or U6616 (N_6616,N_3184,N_4625);
and U6617 (N_6617,N_4401,N_5027);
nand U6618 (N_6618,N_4430,N_4523);
and U6619 (N_6619,N_5025,N_3528);
and U6620 (N_6620,N_4103,N_3631);
and U6621 (N_6621,N_4785,N_5886);
nand U6622 (N_6622,N_6099,N_4264);
and U6623 (N_6623,N_4082,N_3675);
and U6624 (N_6624,N_4087,N_4352);
nor U6625 (N_6625,N_6113,N_3215);
or U6626 (N_6626,N_3452,N_5580);
and U6627 (N_6627,N_4548,N_5257);
xor U6628 (N_6628,N_5582,N_3513);
and U6629 (N_6629,N_4004,N_4712);
nor U6630 (N_6630,N_3580,N_3160);
nand U6631 (N_6631,N_5690,N_5539);
xor U6632 (N_6632,N_3796,N_4937);
nor U6633 (N_6633,N_4054,N_4588);
and U6634 (N_6634,N_3783,N_3676);
nor U6635 (N_6635,N_3163,N_4881);
and U6636 (N_6636,N_6092,N_6138);
nor U6637 (N_6637,N_3721,N_5235);
nor U6638 (N_6638,N_4038,N_5204);
or U6639 (N_6639,N_4444,N_6021);
xnor U6640 (N_6640,N_4425,N_4388);
or U6641 (N_6641,N_4800,N_4921);
xor U6642 (N_6642,N_4208,N_5927);
nor U6643 (N_6643,N_5054,N_5371);
nand U6644 (N_6644,N_5774,N_3654);
and U6645 (N_6645,N_4804,N_5894);
or U6646 (N_6646,N_3269,N_3564);
or U6647 (N_6647,N_4296,N_4922);
or U6648 (N_6648,N_3192,N_5612);
nor U6649 (N_6649,N_3325,N_3742);
or U6650 (N_6650,N_3940,N_4459);
nor U6651 (N_6651,N_4030,N_5760);
nand U6652 (N_6652,N_5959,N_3859);
or U6653 (N_6653,N_5311,N_4788);
or U6654 (N_6654,N_4279,N_3864);
nand U6655 (N_6655,N_3924,N_5866);
nor U6656 (N_6656,N_4348,N_4569);
xnor U6657 (N_6657,N_4105,N_5716);
nor U6658 (N_6658,N_4761,N_3956);
and U6659 (N_6659,N_5765,N_4160);
nand U6660 (N_6660,N_4744,N_5357);
or U6661 (N_6661,N_4637,N_3684);
xor U6662 (N_6662,N_6168,N_4230);
or U6663 (N_6663,N_5377,N_3174);
or U6664 (N_6664,N_3916,N_4036);
xor U6665 (N_6665,N_3608,N_3811);
nor U6666 (N_6666,N_5706,N_3284);
or U6667 (N_6667,N_5781,N_3664);
nand U6668 (N_6668,N_4595,N_4199);
nand U6669 (N_6669,N_3146,N_4289);
nor U6670 (N_6670,N_4191,N_3449);
and U6671 (N_6671,N_4766,N_6053);
and U6672 (N_6672,N_3907,N_5285);
or U6673 (N_6673,N_3929,N_4815);
or U6674 (N_6674,N_6063,N_5495);
and U6675 (N_6675,N_4760,N_4882);
nand U6676 (N_6676,N_5089,N_3258);
or U6677 (N_6677,N_4441,N_6175);
or U6678 (N_6678,N_6202,N_5009);
xnor U6679 (N_6679,N_3490,N_4476);
and U6680 (N_6680,N_3889,N_6241);
nor U6681 (N_6681,N_6190,N_4332);
nand U6682 (N_6682,N_6119,N_3951);
nand U6683 (N_6683,N_5500,N_4945);
or U6684 (N_6684,N_3845,N_5087);
nand U6685 (N_6685,N_5931,N_4445);
or U6686 (N_6686,N_3323,N_4270);
or U6687 (N_6687,N_5130,N_3408);
or U6688 (N_6688,N_5475,N_5514);
nand U6689 (N_6689,N_6192,N_5527);
or U6690 (N_6690,N_4656,N_4839);
or U6691 (N_6691,N_3561,N_4382);
and U6692 (N_6692,N_5244,N_4458);
and U6693 (N_6693,N_6079,N_3138);
or U6694 (N_6694,N_4650,N_3527);
and U6695 (N_6695,N_4316,N_4201);
or U6696 (N_6696,N_3320,N_4952);
or U6697 (N_6697,N_5512,N_5382);
nand U6698 (N_6698,N_3801,N_3747);
nand U6699 (N_6699,N_5263,N_4894);
or U6700 (N_6700,N_4602,N_3292);
and U6701 (N_6701,N_6185,N_4677);
nand U6702 (N_6702,N_3584,N_4605);
and U6703 (N_6703,N_6203,N_3772);
nand U6704 (N_6704,N_4647,N_3738);
nand U6705 (N_6705,N_5265,N_3534);
or U6706 (N_6706,N_6009,N_4137);
xnor U6707 (N_6707,N_5389,N_3594);
nor U6708 (N_6708,N_6026,N_5654);
nor U6709 (N_6709,N_6059,N_5836);
nor U6710 (N_6710,N_4022,N_4475);
and U6711 (N_6711,N_3560,N_4594);
nor U6712 (N_6712,N_5435,N_3302);
xnor U6713 (N_6713,N_3880,N_6028);
nand U6714 (N_6714,N_5545,N_5935);
nor U6715 (N_6715,N_4424,N_3361);
xnor U6716 (N_6716,N_5189,N_4178);
or U6717 (N_6717,N_4915,N_3507);
nor U6718 (N_6718,N_4777,N_6181);
or U6719 (N_6719,N_5463,N_4878);
nand U6720 (N_6720,N_4706,N_4821);
nor U6721 (N_6721,N_3937,N_4386);
xnor U6722 (N_6722,N_5322,N_4197);
nor U6723 (N_6723,N_4726,N_4412);
nand U6724 (N_6724,N_5768,N_4450);
nand U6725 (N_6725,N_3882,N_4210);
nand U6726 (N_6726,N_4380,N_4154);
nand U6727 (N_6727,N_4806,N_3198);
nand U6728 (N_6728,N_4831,N_3473);
nor U6729 (N_6729,N_4143,N_5762);
and U6730 (N_6730,N_3169,N_4260);
nor U6731 (N_6731,N_4724,N_4847);
or U6732 (N_6732,N_4013,N_4940);
nor U6733 (N_6733,N_5506,N_4600);
nand U6734 (N_6734,N_5775,N_5535);
and U6735 (N_6735,N_3185,N_5128);
nand U6736 (N_6736,N_3253,N_3633);
nor U6737 (N_6737,N_3268,N_6049);
nor U6738 (N_6738,N_5921,N_3853);
and U6739 (N_6739,N_4213,N_5334);
nor U6740 (N_6740,N_3318,N_3178);
or U6741 (N_6741,N_4090,N_3941);
and U6742 (N_6742,N_4654,N_5340);
nand U6743 (N_6743,N_5011,N_3207);
nor U6744 (N_6744,N_3873,N_3821);
or U6745 (N_6745,N_5608,N_3511);
and U6746 (N_6746,N_4339,N_4053);
and U6747 (N_6747,N_4652,N_5881);
and U6748 (N_6748,N_4782,N_5524);
and U6749 (N_6749,N_5546,N_3841);
or U6750 (N_6750,N_6047,N_5325);
nor U6751 (N_6751,N_6157,N_5232);
or U6752 (N_6752,N_5969,N_5543);
nor U6753 (N_6753,N_3653,N_4156);
xor U6754 (N_6754,N_3363,N_5777);
or U6755 (N_6755,N_5663,N_4282);
and U6756 (N_6756,N_4792,N_4284);
nand U6757 (N_6757,N_4158,N_5567);
nand U6758 (N_6758,N_5660,N_5012);
or U6759 (N_6759,N_4752,N_4576);
and U6760 (N_6760,N_4287,N_5305);
nand U6761 (N_6761,N_3558,N_3898);
and U6762 (N_6762,N_5989,N_3157);
nand U6763 (N_6763,N_5599,N_5365);
xnor U6764 (N_6764,N_4768,N_5584);
and U6765 (N_6765,N_3295,N_4680);
or U6766 (N_6766,N_3484,N_3234);
xor U6767 (N_6767,N_4517,N_5256);
nor U6768 (N_6768,N_5092,N_4859);
nand U6769 (N_6769,N_5007,N_3603);
nor U6770 (N_6770,N_4397,N_5631);
nor U6771 (N_6771,N_5596,N_4579);
nor U6772 (N_6772,N_4457,N_6249);
nor U6773 (N_6773,N_3373,N_4305);
and U6774 (N_6774,N_5129,N_4059);
nor U6775 (N_6775,N_5139,N_5222);
nand U6776 (N_6776,N_3156,N_3716);
and U6777 (N_6777,N_4128,N_5533);
nand U6778 (N_6778,N_4169,N_4302);
or U6779 (N_6779,N_5835,N_4534);
and U6780 (N_6780,N_5441,N_4556);
xnor U6781 (N_6781,N_3677,N_4037);
nand U6782 (N_6782,N_5610,N_5528);
and U6783 (N_6783,N_6033,N_4603);
and U6784 (N_6784,N_3303,N_3161);
nor U6785 (N_6785,N_4271,N_6121);
nand U6786 (N_6786,N_4884,N_4057);
or U6787 (N_6787,N_3565,N_5046);
nand U6788 (N_6788,N_5266,N_4826);
xnor U6789 (N_6789,N_5858,N_5948);
nand U6790 (N_6790,N_3963,N_4976);
nor U6791 (N_6791,N_5174,N_4989);
and U6792 (N_6792,N_5090,N_4248);
or U6793 (N_6793,N_4372,N_5205);
nand U6794 (N_6794,N_5042,N_4139);
or U6795 (N_6795,N_4025,N_4405);
nand U6796 (N_6796,N_5373,N_5387);
nor U6797 (N_6797,N_4900,N_3876);
or U6798 (N_6798,N_5525,N_4429);
and U6799 (N_6799,N_5702,N_5353);
or U6800 (N_6800,N_4533,N_4499);
nand U6801 (N_6801,N_4622,N_3165);
and U6802 (N_6802,N_4431,N_3460);
nor U6803 (N_6803,N_5687,N_5957);
and U6804 (N_6804,N_5919,N_3241);
and U6805 (N_6805,N_5814,N_4421);
or U6806 (N_6806,N_3997,N_5890);
nand U6807 (N_6807,N_5883,N_5168);
nand U6808 (N_6808,N_3311,N_4816);
or U6809 (N_6809,N_5755,N_3765);
nand U6810 (N_6810,N_3900,N_5770);
nand U6811 (N_6811,N_4186,N_3510);
nor U6812 (N_6812,N_5850,N_4987);
or U6813 (N_6813,N_3905,N_5261);
or U6814 (N_6814,N_3791,N_3667);
and U6815 (N_6815,N_6032,N_6171);
or U6816 (N_6816,N_4269,N_4738);
and U6817 (N_6817,N_5223,N_5227);
xor U6818 (N_6818,N_4074,N_3539);
and U6819 (N_6819,N_5037,N_4140);
and U6820 (N_6820,N_4598,N_4234);
nor U6821 (N_6821,N_5636,N_3866);
nor U6822 (N_6822,N_6111,N_3233);
and U6823 (N_6823,N_4636,N_5169);
xor U6824 (N_6824,N_5833,N_4266);
or U6825 (N_6825,N_4368,N_4917);
nand U6826 (N_6826,N_3315,N_3427);
nor U6827 (N_6827,N_5151,N_5997);
or U6828 (N_6828,N_4400,N_5250);
nor U6829 (N_6829,N_4685,N_5745);
nor U6830 (N_6830,N_5233,N_3572);
and U6831 (N_6831,N_3567,N_5898);
and U6832 (N_6832,N_4144,N_5041);
and U6833 (N_6833,N_4077,N_5950);
and U6834 (N_6834,N_3810,N_3759);
nor U6835 (N_6835,N_4982,N_4763);
or U6836 (N_6836,N_3848,N_5863);
nand U6837 (N_6837,N_5214,N_4983);
or U6838 (N_6838,N_4497,N_3224);
and U6839 (N_6839,N_4345,N_3991);
and U6840 (N_6840,N_3762,N_4779);
nand U6841 (N_6841,N_5122,N_4467);
nor U6842 (N_6842,N_5816,N_5520);
nand U6843 (N_6843,N_4567,N_3562);
and U6844 (N_6844,N_3752,N_3205);
and U6845 (N_6845,N_5852,N_6065);
and U6846 (N_6846,N_5967,N_4301);
nand U6847 (N_6847,N_5696,N_6051);
xnor U6848 (N_6848,N_3599,N_5562);
nor U6849 (N_6849,N_4621,N_3705);
nand U6850 (N_6850,N_6122,N_3881);
nor U6851 (N_6851,N_3478,N_5091);
nor U6852 (N_6852,N_5064,N_3681);
and U6853 (N_6853,N_4047,N_4107);
nand U6854 (N_6854,N_4008,N_5857);
and U6855 (N_6855,N_5383,N_4665);
nor U6856 (N_6856,N_5417,N_5376);
nand U6857 (N_6857,N_3495,N_5759);
nor U6858 (N_6858,N_3431,N_5593);
or U6859 (N_6859,N_3613,N_5979);
nor U6860 (N_6860,N_4558,N_5196);
or U6861 (N_6861,N_5549,N_4512);
and U6862 (N_6862,N_3249,N_3644);
nor U6863 (N_6863,N_4065,N_5456);
nor U6864 (N_6864,N_5916,N_4614);
nor U6865 (N_6865,N_5737,N_4872);
xnor U6866 (N_6866,N_4488,N_5877);
nand U6867 (N_6867,N_4871,N_6209);
nand U6868 (N_6868,N_5569,N_4012);
or U6869 (N_6869,N_4050,N_5422);
nor U6870 (N_6870,N_6045,N_5180);
or U6871 (N_6871,N_4455,N_4180);
or U6872 (N_6872,N_4657,N_4073);
nor U6873 (N_6873,N_4064,N_3652);
nand U6874 (N_6874,N_5043,N_4920);
nor U6875 (N_6875,N_4205,N_4035);
nand U6876 (N_6876,N_5575,N_5144);
xnor U6877 (N_6877,N_5534,N_3347);
xor U6878 (N_6878,N_4718,N_3461);
xor U6879 (N_6879,N_5733,N_4033);
nand U6880 (N_6880,N_3403,N_3955);
nor U6881 (N_6881,N_6075,N_5156);
xor U6882 (N_6882,N_4627,N_4998);
nand U6883 (N_6883,N_3959,N_4597);
nand U6884 (N_6884,N_5453,N_3549);
or U6885 (N_6885,N_3533,N_3847);
or U6886 (N_6886,N_4704,N_6222);
or U6887 (N_6887,N_6008,N_5402);
xnor U6888 (N_6888,N_5203,N_5842);
or U6889 (N_6889,N_5922,N_3398);
or U6890 (N_6890,N_4960,N_3171);
nand U6891 (N_6891,N_4972,N_5868);
nand U6892 (N_6892,N_4754,N_4640);
nor U6893 (N_6893,N_5929,N_4527);
nor U6894 (N_6894,N_3319,N_5310);
or U6895 (N_6895,N_4496,N_4732);
and U6896 (N_6896,N_3497,N_6058);
or U6897 (N_6897,N_4374,N_4283);
or U6898 (N_6898,N_4174,N_3410);
and U6899 (N_6899,N_5465,N_4267);
or U6900 (N_6900,N_3164,N_4219);
and U6901 (N_6901,N_5199,N_6109);
xnor U6902 (N_6902,N_3748,N_5388);
xor U6903 (N_6903,N_4491,N_5744);
or U6904 (N_6904,N_3434,N_5885);
and U6905 (N_6905,N_4563,N_5911);
nand U6906 (N_6906,N_3746,N_3808);
xor U6907 (N_6907,N_3332,N_4218);
nor U6908 (N_6908,N_4069,N_4638);
nor U6909 (N_6909,N_6067,N_4837);
or U6910 (N_6910,N_3632,N_5274);
nand U6911 (N_6911,N_4229,N_3459);
nor U6912 (N_6912,N_4928,N_5461);
and U6913 (N_6913,N_4472,N_4562);
and U6914 (N_6914,N_5719,N_3426);
or U6915 (N_6915,N_4722,N_4461);
and U6916 (N_6916,N_5201,N_3259);
nand U6917 (N_6917,N_4176,N_5570);
and U6918 (N_6918,N_4225,N_4375);
xor U6919 (N_6919,N_5114,N_4150);
nor U6920 (N_6920,N_6235,N_5362);
or U6921 (N_6921,N_3755,N_4506);
nor U6922 (N_6922,N_3255,N_3378);
xnor U6923 (N_6923,N_5633,N_5014);
nor U6924 (N_6924,N_4360,N_4734);
or U6925 (N_6925,N_3993,N_5167);
and U6926 (N_6926,N_4741,N_3851);
nand U6927 (N_6927,N_3299,N_4362);
xor U6928 (N_6928,N_4039,N_3509);
nor U6929 (N_6929,N_5825,N_4194);
xor U6930 (N_6930,N_3871,N_4805);
or U6931 (N_6931,N_3718,N_4046);
nor U6932 (N_6932,N_4731,N_5920);
nor U6933 (N_6933,N_4434,N_5531);
and U6934 (N_6934,N_5592,N_3686);
and U6935 (N_6935,N_3344,N_3387);
nand U6936 (N_6936,N_6212,N_4398);
nor U6937 (N_6937,N_3199,N_3601);
and U6938 (N_6938,N_6242,N_3744);
or U6939 (N_6939,N_3143,N_6196);
nor U6940 (N_6940,N_3740,N_4832);
or U6941 (N_6941,N_5598,N_3474);
xnor U6942 (N_6942,N_5397,N_3256);
and U6943 (N_6943,N_4165,N_4297);
and U6944 (N_6944,N_5671,N_5403);
or U6945 (N_6945,N_4281,N_3422);
nor U6946 (N_6946,N_3680,N_5655);
or U6947 (N_6947,N_3214,N_3152);
or U6948 (N_6948,N_4273,N_5297);
nor U6949 (N_6949,N_3928,N_4714);
nor U6950 (N_6950,N_5793,N_4659);
nand U6951 (N_6951,N_4623,N_5981);
or U6952 (N_6952,N_4392,N_3552);
and U6953 (N_6953,N_5462,N_3376);
nor U6954 (N_6954,N_4114,N_3555);
or U6955 (N_6955,N_3217,N_3154);
and U6956 (N_6956,N_4557,N_5766);
nor U6957 (N_6957,N_5792,N_3285);
nor U6958 (N_6958,N_6035,N_5290);
nor U6959 (N_6959,N_5878,N_4699);
nand U6960 (N_6960,N_3734,N_5522);
xor U6961 (N_6961,N_3945,N_5689);
nand U6962 (N_6962,N_5198,N_5998);
or U6963 (N_6963,N_5616,N_4032);
nand U6964 (N_6964,N_3711,N_5315);
or U6965 (N_6965,N_4529,N_6091);
nor U6966 (N_6966,N_5170,N_5917);
and U6967 (N_6967,N_3826,N_4503);
and U6968 (N_6968,N_3158,N_3757);
nor U6969 (N_6969,N_5668,N_3970);
and U6970 (N_6970,N_4334,N_3856);
nor U6971 (N_6971,N_5164,N_3314);
or U6972 (N_6972,N_3725,N_3781);
xnor U6973 (N_6973,N_4017,N_5647);
and U6974 (N_6974,N_3491,N_4912);
nor U6975 (N_6975,N_4876,N_4740);
and U6976 (N_6976,N_5354,N_3974);
nor U6977 (N_6977,N_4990,N_4736);
or U6978 (N_6978,N_6193,N_6230);
xnor U6979 (N_6979,N_4924,N_3660);
and U6980 (N_6980,N_4755,N_3678);
and U6981 (N_6981,N_3439,N_4494);
nor U6982 (N_6982,N_5248,N_3990);
xor U6983 (N_6983,N_5788,N_5855);
xnor U6984 (N_6984,N_3485,N_5302);
nand U6985 (N_6985,N_3504,N_4118);
nor U6986 (N_6986,N_5925,N_5682);
and U6987 (N_6987,N_6120,N_5870);
nor U6988 (N_6988,N_6112,N_4592);
or U6989 (N_6989,N_3626,N_4554);
and U6990 (N_6990,N_4049,N_5798);
and U6991 (N_6991,N_5828,N_5375);
nand U6992 (N_6992,N_4227,N_4280);
or U6993 (N_6993,N_5125,N_5676);
or U6994 (N_6994,N_4547,N_3351);
or U6995 (N_6995,N_5338,N_5421);
and U6996 (N_6996,N_6070,N_6144);
and U6997 (N_6997,N_6105,N_3797);
nand U6998 (N_6998,N_5252,N_5799);
and U6999 (N_6999,N_3575,N_3271);
nand U7000 (N_7000,N_3739,N_5071);
nand U7001 (N_7001,N_4758,N_5619);
nor U7002 (N_7002,N_4078,N_3254);
nand U7003 (N_7003,N_4531,N_6188);
and U7004 (N_7004,N_3529,N_5893);
nor U7005 (N_7005,N_4697,N_6206);
xor U7006 (N_7006,N_5563,N_3362);
nor U7007 (N_7007,N_3476,N_3424);
and U7008 (N_7008,N_4106,N_3642);
or U7009 (N_7009,N_4385,N_4639);
nand U7010 (N_7010,N_3231,N_5552);
or U7011 (N_7011,N_4370,N_4814);
nand U7012 (N_7012,N_4121,N_5587);
xnor U7013 (N_7013,N_3697,N_4336);
and U7014 (N_7014,N_5738,N_4918);
nand U7015 (N_7015,N_4089,N_5454);
and U7016 (N_7016,N_5173,N_4242);
xnor U7017 (N_7017,N_4661,N_5909);
nand U7018 (N_7018,N_4045,N_3670);
nor U7019 (N_7019,N_5521,N_3629);
nor U7020 (N_7020,N_3499,N_4246);
nor U7021 (N_7021,N_4916,N_5468);
nor U7022 (N_7022,N_5700,N_6003);
nand U7023 (N_7023,N_4539,N_3688);
or U7024 (N_7024,N_6166,N_5286);
nand U7025 (N_7025,N_3920,N_4340);
or U7026 (N_7026,N_5588,N_5347);
or U7027 (N_7027,N_4006,N_3911);
nand U7028 (N_7028,N_4725,N_3385);
xnor U7029 (N_7029,N_6160,N_4179);
xor U7030 (N_7030,N_3179,N_4721);
xor U7031 (N_7031,N_3915,N_5910);
or U7032 (N_7032,N_4931,N_3469);
nand U7033 (N_7033,N_3291,N_4855);
xnor U7034 (N_7034,N_5722,N_5326);
and U7035 (N_7035,N_3593,N_5005);
nand U7036 (N_7036,N_5756,N_4873);
xnor U7037 (N_7037,N_5035,N_3239);
nand U7038 (N_7038,N_3244,N_6019);
nor U7039 (N_7039,N_3279,N_5913);
nor U7040 (N_7040,N_3611,N_3914);
xnor U7041 (N_7041,N_3297,N_6068);
nand U7042 (N_7042,N_3267,N_5516);
nor U7043 (N_7043,N_5185,N_6106);
or U7044 (N_7044,N_5380,N_6214);
or U7045 (N_7045,N_3984,N_4875);
or U7046 (N_7046,N_3610,N_3775);
xor U7047 (N_7047,N_4845,N_4907);
or U7048 (N_7048,N_4772,N_4262);
nor U7049 (N_7049,N_4484,N_5725);
or U7050 (N_7050,N_5243,N_4781);
or U7051 (N_7051,N_4117,N_3189);
nor U7052 (N_7052,N_3273,N_3524);
nor U7053 (N_7053,N_3634,N_4468);
nand U7054 (N_7054,N_4011,N_3283);
nand U7055 (N_7055,N_5412,N_4084);
and U7056 (N_7056,N_3316,N_5795);
nor U7057 (N_7057,N_5217,N_4935);
xor U7058 (N_7058,N_4500,N_5556);
nand U7059 (N_7059,N_5990,N_5313);
nand U7060 (N_7060,N_3393,N_5903);
xor U7061 (N_7061,N_5324,N_5505);
xor U7062 (N_7062,N_5965,N_4005);
xor U7063 (N_7063,N_5854,N_3890);
nand U7064 (N_7064,N_3322,N_4711);
and U7065 (N_7065,N_3286,N_3506);
xnor U7066 (N_7066,N_3566,N_5887);
and U7067 (N_7067,N_6136,N_5272);
or U7068 (N_7068,N_5356,N_3425);
and U7069 (N_7069,N_5635,N_5249);
or U7070 (N_7070,N_5352,N_4446);
nor U7071 (N_7071,N_5841,N_5405);
xor U7072 (N_7072,N_6041,N_3814);
or U7073 (N_7073,N_5984,N_6146);
nand U7074 (N_7074,N_6125,N_4513);
nor U7075 (N_7075,N_5312,N_4784);
nand U7076 (N_7076,N_5603,N_3301);
xor U7077 (N_7077,N_3800,N_3894);
or U7078 (N_7078,N_6057,N_5492);
nor U7079 (N_7079,N_5052,N_5394);
or U7080 (N_7080,N_3823,N_4040);
and U7081 (N_7081,N_4955,N_5649);
nor U7082 (N_7082,N_5409,N_5318);
nand U7083 (N_7083,N_5574,N_4294);
xnor U7084 (N_7084,N_5003,N_3930);
nand U7085 (N_7085,N_5694,N_4930);
nand U7086 (N_7086,N_3922,N_5015);
and U7087 (N_7087,N_6055,N_6164);
xor U7088 (N_7088,N_3145,N_4692);
or U7089 (N_7089,N_3661,N_6022);
nand U7090 (N_7090,N_4846,N_5832);
nand U7091 (N_7091,N_4642,N_3245);
or U7092 (N_7092,N_5586,N_5195);
nor U7093 (N_7093,N_5131,N_3753);
or U7094 (N_7094,N_4070,N_3702);
and U7095 (N_7095,N_6131,N_3590);
and U7096 (N_7096,N_3372,N_5058);
nor U7097 (N_7097,N_6030,N_4515);
xnor U7098 (N_7098,N_4470,N_5617);
nand U7099 (N_7099,N_6062,N_3243);
nor U7100 (N_7100,N_3630,N_3569);
xnor U7101 (N_7101,N_5102,N_6011);
nor U7102 (N_7102,N_4852,N_5466);
or U7103 (N_7103,N_4439,N_5707);
or U7104 (N_7104,N_4951,N_3604);
nand U7105 (N_7105,N_6149,N_5494);
nand U7106 (N_7106,N_4560,N_4256);
and U7107 (N_7107,N_3257,N_4215);
nand U7108 (N_7108,N_3720,N_6078);
xor U7109 (N_7109,N_3844,N_3902);
nand U7110 (N_7110,N_6137,N_5634);
nand U7111 (N_7111,N_4510,N_5333);
nor U7112 (N_7112,N_5824,N_5218);
and U7113 (N_7113,N_3141,N_3345);
nand U7114 (N_7114,N_3986,N_5753);
and U7115 (N_7115,N_3835,N_3840);
nor U7116 (N_7116,N_3381,N_4645);
or U7117 (N_7117,N_3743,N_6076);
nor U7118 (N_7118,N_5123,N_4373);
or U7119 (N_7119,N_4705,N_4321);
nand U7120 (N_7120,N_4237,N_4286);
or U7121 (N_7121,N_3717,N_3238);
nand U7122 (N_7122,N_3409,N_3828);
and U7123 (N_7123,N_4292,N_5643);
nand U7124 (N_7124,N_3985,N_5247);
xor U7125 (N_7125,N_3208,N_5819);
or U7126 (N_7126,N_5801,N_4545);
nand U7127 (N_7127,N_4820,N_5428);
or U7128 (N_7128,N_4966,N_4235);
xnor U7129 (N_7129,N_3196,N_5727);
or U7130 (N_7130,N_3450,N_3213);
nor U7131 (N_7131,N_4967,N_5400);
or U7132 (N_7132,N_5307,N_3338);
nand U7133 (N_7133,N_4189,N_5477);
nand U7134 (N_7134,N_5155,N_4066);
nor U7135 (N_7135,N_5837,N_4811);
and U7136 (N_7136,N_5255,N_4733);
nor U7137 (N_7137,N_4885,N_5363);
or U7138 (N_7138,N_6184,N_4111);
nand U7139 (N_7139,N_4369,N_5026);
nor U7140 (N_7140,N_5688,N_5320);
nor U7141 (N_7141,N_3925,N_4238);
nand U7142 (N_7142,N_6245,N_4888);
xor U7143 (N_7143,N_6187,N_5656);
nand U7144 (N_7144,N_4226,N_5879);
or U7145 (N_7145,N_4973,N_3691);
and U7146 (N_7146,N_4672,N_4469);
and U7147 (N_7147,N_4306,N_6087);
and U7148 (N_7148,N_4971,N_5392);
nand U7149 (N_7149,N_4344,N_5410);
or U7150 (N_7150,N_4801,N_6244);
nand U7151 (N_7151,N_5747,N_4493);
and U7152 (N_7152,N_4962,N_4765);
and U7153 (N_7153,N_4153,N_4062);
nand U7154 (N_7154,N_4756,N_3219);
or U7155 (N_7155,N_4838,N_4436);
nor U7156 (N_7156,N_5236,N_3374);
or U7157 (N_7157,N_4231,N_5499);
and U7158 (N_7158,N_5875,N_4817);
nor U7159 (N_7159,N_5548,N_4119);
or U7160 (N_7160,N_3423,N_5420);
nand U7161 (N_7161,N_5540,N_5057);
nor U7162 (N_7162,N_3982,N_3187);
and U7163 (N_7163,N_5344,N_3719);
nor U7164 (N_7164,N_3903,N_5022);
or U7165 (N_7165,N_4913,N_5609);
nand U7166 (N_7166,N_3585,N_3874);
nand U7167 (N_7167,N_5474,N_4315);
and U7168 (N_7168,N_5226,N_3274);
and U7169 (N_7169,N_3488,N_3628);
and U7170 (N_7170,N_5497,N_4858);
nand U7171 (N_7171,N_3785,N_3479);
nand U7172 (N_7172,N_5715,N_4526);
or U7173 (N_7173,N_3949,N_3308);
nand U7174 (N_7174,N_4694,N_5996);
and U7175 (N_7175,N_4964,N_5079);
and U7176 (N_7176,N_4764,N_4326);
nand U7177 (N_7177,N_5752,N_4701);
and U7178 (N_7178,N_5337,N_4961);
and U7179 (N_7179,N_6228,N_4093);
xnor U7180 (N_7180,N_5098,N_6043);
or U7181 (N_7181,N_3701,N_5251);
or U7182 (N_7182,N_5739,N_3700);
or U7183 (N_7183,N_4125,N_5564);
or U7184 (N_7184,N_3155,N_5332);
or U7185 (N_7185,N_3953,N_5968);
and U7186 (N_7186,N_6141,N_4867);
and U7187 (N_7187,N_5791,N_5157);
or U7188 (N_7188,N_3126,N_6218);
or U7189 (N_7189,N_3494,N_4435);
and U7190 (N_7190,N_5677,N_4914);
nor U7191 (N_7191,N_4474,N_3519);
nand U7192 (N_7192,N_6142,N_3518);
or U7193 (N_7193,N_3999,N_5416);
or U7194 (N_7194,N_4031,N_5743);
nand U7195 (N_7195,N_6129,N_4320);
and U7196 (N_7196,N_5124,N_4241);
or U7197 (N_7197,N_4254,N_5234);
nand U7198 (N_7198,N_3153,N_5384);
xor U7199 (N_7199,N_5401,N_4611);
and U7200 (N_7200,N_5807,N_4789);
nand U7201 (N_7201,N_3441,N_6217);
and U7202 (N_7202,N_5637,N_4674);
and U7203 (N_7203,N_4480,N_5511);
or U7204 (N_7204,N_6232,N_5268);
xor U7205 (N_7205,N_6060,N_3952);
xor U7206 (N_7206,N_3829,N_5999);
or U7207 (N_7207,N_5291,N_4713);
or U7208 (N_7208,N_3309,N_4245);
and U7209 (N_7209,N_6056,N_3788);
nor U7210 (N_7210,N_4956,N_6207);
nor U7211 (N_7211,N_5585,N_5889);
xor U7212 (N_7212,N_5000,N_5786);
nor U7213 (N_7213,N_5224,N_5452);
and U7214 (N_7214,N_5216,N_4479);
nand U7215 (N_7215,N_5211,N_3414);
or U7216 (N_7216,N_4578,N_3827);
nand U7217 (N_7217,N_5084,N_3571);
nand U7218 (N_7218,N_4925,N_3277);
or U7219 (N_7219,N_5166,N_4686);
nand U7220 (N_7220,N_4120,N_5583);
or U7221 (N_7221,N_3443,N_3623);
xnor U7222 (N_7222,N_6123,N_6126);
nand U7223 (N_7223,N_4828,N_6247);
and U7224 (N_7224,N_4537,N_4580);
and U7225 (N_7225,N_5240,N_6159);
and U7226 (N_7226,N_5013,N_3954);
nor U7227 (N_7227,N_3190,N_4633);
or U7228 (N_7228,N_4670,N_6095);
and U7229 (N_7229,N_5709,N_3324);
or U7230 (N_7230,N_3819,N_4827);
nor U7231 (N_7231,N_5262,N_6147);
nor U7232 (N_7232,N_4108,N_5942);
nor U7233 (N_7233,N_5742,N_4644);
and U7234 (N_7234,N_4997,N_6237);
or U7235 (N_7235,N_5896,N_4349);
xor U7236 (N_7236,N_4819,N_5674);
and U7237 (N_7237,N_5805,N_4009);
and U7238 (N_7238,N_3246,N_3968);
and U7239 (N_7239,N_4185,N_4378);
nand U7240 (N_7240,N_5208,N_4771);
nor U7241 (N_7241,N_4432,N_4748);
nand U7242 (N_7242,N_4901,N_4769);
and U7243 (N_7243,N_5779,N_5971);
nor U7244 (N_7244,N_4555,N_5672);
and U7245 (N_7245,N_3589,N_3206);
and U7246 (N_7246,N_3400,N_5578);
nor U7247 (N_7247,N_5595,N_4612);
xnor U7248 (N_7248,N_5478,N_5479);
and U7249 (N_7249,N_4261,N_4635);
or U7250 (N_7250,N_5321,N_5508);
nand U7251 (N_7251,N_6170,N_5303);
or U7252 (N_7252,N_4853,N_3464);
nand U7253 (N_7253,N_3194,N_3703);
and U7254 (N_7254,N_3766,N_4007);
nand U7255 (N_7255,N_6176,N_4399);
or U7256 (N_7256,N_4331,N_4288);
nand U7257 (N_7257,N_4097,N_4177);
and U7258 (N_7258,N_6012,N_3183);
nand U7259 (N_7259,N_3525,N_4743);
or U7260 (N_7260,N_4255,N_3648);
nand U7261 (N_7261,N_4131,N_6034);
nand U7262 (N_7262,N_3722,N_4240);
nor U7263 (N_7263,N_5937,N_5544);
nor U7264 (N_7264,N_5343,N_4851);
nor U7265 (N_7265,N_5553,N_5229);
xnor U7266 (N_7266,N_4932,N_3942);
nor U7267 (N_7267,N_5470,N_4346);
or U7268 (N_7268,N_3360,N_5778);
and U7269 (N_7269,N_6151,N_6186);
nand U7270 (N_7270,N_5486,N_3366);
or U7271 (N_7271,N_5150,N_5053);
or U7272 (N_7272,N_3994,N_4098);
nor U7273 (N_7273,N_5140,N_3553);
nand U7274 (N_7274,N_4453,N_3350);
xnor U7275 (N_7275,N_5282,N_3958);
or U7276 (N_7276,N_3938,N_5908);
xor U7277 (N_7277,N_4664,N_3779);
and U7278 (N_7278,N_3306,N_5407);
or U7279 (N_7279,N_6143,N_4571);
nor U7280 (N_7280,N_4110,N_3771);
nor U7281 (N_7281,N_5237,N_6238);
or U7282 (N_7282,N_3211,N_4202);
xnor U7283 (N_7283,N_3252,N_3698);
xor U7284 (N_7284,N_5691,N_4616);
nor U7285 (N_7285,N_3839,N_5720);
nand U7286 (N_7286,N_4946,N_3899);
nor U7287 (N_7287,N_5653,N_5932);
and U7288 (N_7288,N_6046,N_5059);
or U7289 (N_7289,N_5986,N_4473);
xnor U7290 (N_7290,N_3758,N_3365);
nor U7291 (N_7291,N_5915,N_3973);
nand U7292 (N_7292,N_6225,N_5607);
or U7293 (N_7293,N_5589,N_6069);
xor U7294 (N_7294,N_5348,N_5289);
and U7295 (N_7295,N_5083,N_4899);
nor U7296 (N_7296,N_3967,N_5136);
nor U7297 (N_7297,N_3220,N_4923);
nand U7298 (N_7298,N_6229,N_3665);
nor U7299 (N_7299,N_4395,N_5258);
xor U7300 (N_7300,N_3995,N_3983);
nor U7301 (N_7301,N_4233,N_4822);
nor U7302 (N_7302,N_3444,N_5171);
nor U7303 (N_7303,N_3622,N_4420);
nand U7304 (N_7304,N_5489,N_3979);
nor U7305 (N_7305,N_3466,N_3723);
and U7306 (N_7306,N_5259,N_3870);
or U7307 (N_7307,N_4799,N_3830);
and U7308 (N_7308,N_3487,N_4146);
nand U7309 (N_7309,N_6165,N_5993);
and U7310 (N_7310,N_5459,N_3335);
nand U7311 (N_7311,N_4681,N_3261);
and U7312 (N_7312,N_4055,N_3689);
nand U7313 (N_7313,N_4553,N_4440);
nand U7314 (N_7314,N_5120,N_6180);
nor U7315 (N_7315,N_5764,N_4662);
nor U7316 (N_7316,N_5177,N_3516);
or U7317 (N_7317,N_4651,N_6042);
or U7318 (N_7318,N_6104,N_5632);
xnor U7319 (N_7319,N_5426,N_3597);
xor U7320 (N_7320,N_3887,N_6227);
and U7321 (N_7321,N_3732,N_4048);
nor U7322 (N_7322,N_4624,N_4892);
or U7323 (N_7323,N_5542,N_4276);
and U7324 (N_7324,N_3596,N_6124);
xnor U7325 (N_7325,N_4358,N_5460);
nand U7326 (N_7326,N_4052,N_5361);
xnor U7327 (N_7327,N_4629,N_6139);
nand U7328 (N_7328,N_3167,N_6199);
or U7329 (N_7329,N_5537,N_4366);
nand U7330 (N_7330,N_4776,N_3886);
nand U7331 (N_7331,N_3710,N_6101);
nor U7332 (N_7332,N_3209,N_5358);
nand U7333 (N_7333,N_3547,N_4948);
xor U7334 (N_7334,N_5010,N_3131);
nor U7335 (N_7335,N_5442,N_4155);
or U7336 (N_7336,N_5748,N_5366);
nor U7337 (N_7337,N_5659,N_3310);
nor U7338 (N_7338,N_3404,N_5884);
xnor U7339 (N_7339,N_4371,N_4880);
and U7340 (N_7340,N_4337,N_3591);
nor U7341 (N_7341,N_5962,N_5068);
or U7342 (N_7342,N_4688,N_5393);
xnor U7343 (N_7343,N_4996,N_5808);
nor U7344 (N_7344,N_4550,N_4109);
nor U7345 (N_7345,N_5646,N_5827);
or U7346 (N_7346,N_4609,N_4606);
and U7347 (N_7347,N_4350,N_6037);
and U7348 (N_7348,N_4628,N_3946);
nor U7349 (N_7349,N_5094,N_5278);
and U7350 (N_7350,N_4818,N_4528);
nand U7351 (N_7351,N_4214,N_3578);
or U7352 (N_7352,N_3804,N_3996);
or U7353 (N_7353,N_5864,N_4809);
or U7354 (N_7354,N_4849,N_3304);
nor U7355 (N_7355,N_4216,N_3130);
nand U7356 (N_7356,N_6150,N_5705);
or U7357 (N_7357,N_4324,N_5165);
or U7358 (N_7358,N_4196,N_3346);
and U7359 (N_7359,N_3761,N_5888);
nand U7360 (N_7360,N_5364,N_3607);
and U7361 (N_7361,N_4546,N_3892);
nand U7362 (N_7362,N_5880,N_3861);
or U7363 (N_7363,N_5276,N_3263);
nor U7364 (N_7364,N_5661,N_3627);
nor U7365 (N_7365,N_6098,N_4643);
or U7366 (N_7366,N_5600,N_6231);
nand U7367 (N_7367,N_4408,N_4676);
or U7368 (N_7368,N_4019,N_4193);
nand U7369 (N_7369,N_5736,N_5072);
xor U7370 (N_7370,N_3242,N_5952);
or U7371 (N_7371,N_5658,N_3806);
and U7372 (N_7372,N_4974,N_5602);
nor U7373 (N_7373,N_4487,N_5191);
and U7374 (N_7374,N_4293,N_4682);
and U7375 (N_7375,N_4482,N_5288);
or U7376 (N_7376,N_6182,N_4950);
or U7377 (N_7377,N_3638,N_5438);
nand U7378 (N_7378,N_5269,N_6194);
nand U7379 (N_7379,N_4856,N_4893);
nor U7380 (N_7380,N_5143,N_3358);
or U7381 (N_7381,N_4166,N_5517);
nand U7382 (N_7382,N_3482,N_4308);
and U7383 (N_7383,N_5228,N_5213);
and U7384 (N_7384,N_5133,N_3637);
or U7385 (N_7385,N_5845,N_3397);
xor U7386 (N_7386,N_5951,N_5493);
xor U7387 (N_7387,N_3728,N_4999);
or U7388 (N_7388,N_3815,N_3445);
or U7389 (N_7389,N_4257,N_4668);
and U7390 (N_7390,N_5061,N_3226);
or U7391 (N_7391,N_3645,N_5314);
nand U7392 (N_7392,N_6074,N_5667);
nand U7393 (N_7393,N_5622,N_4719);
nor U7394 (N_7394,N_5152,N_5577);
and U7395 (N_7395,N_4361,N_3838);
xor U7396 (N_7396,N_4072,N_4024);
or U7397 (N_7397,N_5536,N_3640);
nand U7398 (N_7398,N_6002,N_3210);
and U7399 (N_7399,N_5983,N_3948);
nor U7400 (N_7400,N_6189,N_5815);
and U7401 (N_7401,N_3435,N_3910);
nor U7402 (N_7402,N_6084,N_3745);
nand U7403 (N_7403,N_3288,N_5963);
or U7404 (N_7404,N_4957,N_4988);
nand U7405 (N_7405,N_3305,N_4132);
nand U7406 (N_7406,N_4327,N_4813);
and U7407 (N_7407,N_4096,N_5519);
nor U7408 (N_7408,N_3773,N_3969);
nor U7409 (N_7409,N_3685,N_3416);
or U7410 (N_7410,N_4933,N_5876);
or U7411 (N_7411,N_4347,N_3200);
and U7412 (N_7412,N_3834,N_5088);
nor U7413 (N_7413,N_5541,N_3150);
xor U7414 (N_7414,N_4689,N_5242);
or U7415 (N_7415,N_5831,N_5782);
nor U7416 (N_7416,N_5184,N_5413);
and U7417 (N_7417,N_3352,N_4471);
and U7418 (N_7418,N_4844,N_3605);
nand U7419 (N_7419,N_6172,N_5627);
or U7420 (N_7420,N_6158,N_3846);
and U7421 (N_7421,N_3522,N_3913);
and U7422 (N_7422,N_5834,N_3987);
or U7423 (N_7423,N_3863,N_5346);
xnor U7424 (N_7424,N_6097,N_5683);
and U7425 (N_7425,N_6135,N_3544);
or U7426 (N_7426,N_4314,N_3465);
nand U7427 (N_7427,N_3468,N_5652);
nor U7428 (N_7428,N_5121,N_5955);
nor U7429 (N_7429,N_6173,N_4544);
nor U7430 (N_7430,N_3232,N_4596);
nor U7431 (N_7431,N_4954,N_4690);
xnor U7432 (N_7432,N_5605,N_3265);
or U7433 (N_7433,N_3250,N_4812);
nand U7434 (N_7434,N_5038,N_3805);
and U7435 (N_7435,N_3917,N_4992);
nand U7436 (N_7436,N_3540,N_4619);
and U7437 (N_7437,N_5193,N_4116);
nand U7438 (N_7438,N_5067,N_4543);
or U7439 (N_7439,N_4860,N_5112);
or U7440 (N_7440,N_5936,N_5391);
nor U7441 (N_7441,N_3570,N_6102);
nor U7442 (N_7442,N_4874,N_5024);
nand U7443 (N_7443,N_4723,N_3515);
or U7444 (N_7444,N_3707,N_3133);
xor U7445 (N_7445,N_5369,N_4224);
nor U7446 (N_7446,N_5048,N_3619);
xor U7447 (N_7447,N_3477,N_6018);
and U7448 (N_7448,N_4841,N_3600);
or U7449 (N_7449,N_4509,N_5415);
nand U7450 (N_7450,N_5107,N_3500);
nor U7451 (N_7451,N_4984,N_4423);
nand U7452 (N_7452,N_4767,N_3433);
nor U7453 (N_7453,N_5679,N_3646);
nand U7454 (N_7454,N_6216,N_4869);
and U7455 (N_7455,N_5081,N_4485);
and U7456 (N_7456,N_4209,N_3975);
nand U7457 (N_7457,N_3872,N_3379);
nand U7458 (N_7458,N_3927,N_5359);
nand U7459 (N_7459,N_4969,N_5735);
nor U7460 (N_7460,N_4275,N_3290);
or U7461 (N_7461,N_6044,N_6248);
nand U7462 (N_7462,N_4979,N_3195);
or U7463 (N_7463,N_6128,N_5439);
nand U7464 (N_7464,N_3548,N_3650);
nor U7465 (N_7465,N_4986,N_3965);
nand U7466 (N_7466,N_3203,N_4483);
and U7467 (N_7467,N_4993,N_3382);
nor U7468 (N_7468,N_5813,N_6197);
and U7469 (N_7469,N_5374,N_4710);
and U7470 (N_7470,N_4759,N_3668);
nand U7471 (N_7471,N_4076,N_4823);
nor U7472 (N_7472,N_4041,N_3843);
xor U7473 (N_7473,N_5941,N_3550);
or U7474 (N_7474,N_5078,N_5277);
and U7475 (N_7475,N_4145,N_4727);
or U7476 (N_7476,N_3546,N_5822);
nor U7477 (N_7477,N_4709,N_3355);
or U7478 (N_7478,N_5900,N_5372);
and U7479 (N_7479,N_5513,N_3384);
or U7480 (N_7480,N_5419,N_4364);
or U7481 (N_7481,N_5529,N_4410);
nand U7482 (N_7482,N_3216,N_3624);
xor U7483 (N_7483,N_5843,N_5992);
nand U7484 (N_7484,N_5840,N_6204);
nand U7485 (N_7485,N_5970,N_3177);
or U7486 (N_7486,N_4730,N_5515);
nand U7487 (N_7487,N_3172,N_5158);
nand U7488 (N_7488,N_6014,N_3885);
or U7489 (N_7489,N_3857,N_3421);
nor U7490 (N_7490,N_3364,N_4944);
nand U7491 (N_7491,N_3673,N_4437);
or U7492 (N_7492,N_4583,N_5188);
xnor U7493 (N_7493,N_5082,N_3807);
and U7494 (N_7494,N_5629,N_5665);
nand U7495 (N_7495,N_5703,N_3370);
nand U7496 (N_7496,N_6223,N_5436);
nor U7497 (N_7497,N_5469,N_4864);
or U7498 (N_7498,N_5215,N_4416);
nand U7499 (N_7499,N_5491,N_3908);
and U7500 (N_7500,N_4162,N_6072);
or U7501 (N_7501,N_5135,N_3581);
nand U7502 (N_7502,N_5678,N_5928);
nor U7503 (N_7503,N_6127,N_3278);
nor U7504 (N_7504,N_6082,N_5796);
nand U7505 (N_7505,N_4505,N_3531);
or U7506 (N_7506,N_3694,N_5772);
xnor U7507 (N_7507,N_3618,N_6017);
nor U7508 (N_7508,N_4182,N_3270);
or U7509 (N_7509,N_5551,N_4122);
nand U7510 (N_7510,N_5434,N_4669);
nor U7511 (N_7511,N_4787,N_4291);
xnor U7512 (N_7512,N_4519,N_4879);
nand U7513 (N_7513,N_4865,N_3598);
nor U7514 (N_7514,N_4161,N_5190);
or U7515 (N_7515,N_5487,N_4263);
xnor U7516 (N_7516,N_3774,N_4863);
and U7517 (N_7517,N_4212,N_4323);
and U7518 (N_7518,N_6240,N_5298);
nor U7519 (N_7519,N_3168,N_3971);
or U7520 (N_7520,N_5614,N_5209);
nor U7521 (N_7521,N_6027,N_6085);
or U7522 (N_7522,N_4728,N_5804);
and U7523 (N_7523,N_3412,N_5020);
and U7524 (N_7524,N_3296,N_5892);
nor U7525 (N_7525,N_4540,N_4325);
and U7526 (N_7526,N_5891,N_3926);
xor U7527 (N_7527,N_5108,N_4749);
nand U7528 (N_7528,N_3188,N_4002);
nor U7529 (N_7529,N_4413,N_5958);
or U7530 (N_7530,N_5080,N_5176);
or U7531 (N_7531,N_5430,N_4123);
xor U7532 (N_7532,N_4574,N_3307);
and U7533 (N_7533,N_4843,N_3429);
xor U7534 (N_7534,N_4663,N_4751);
and U7535 (N_7535,N_3662,N_4498);
or U7536 (N_7536,N_3904,N_5797);
or U7537 (N_7537,N_6040,N_3595);
or U7538 (N_7538,N_3462,N_3127);
xnor U7539 (N_7539,N_6239,N_3201);
xnor U7540 (N_7540,N_5221,N_4295);
or U7541 (N_7541,N_4551,N_4591);
nor U7542 (N_7542,N_3895,N_5446);
and U7543 (N_7543,N_5579,N_5270);
or U7544 (N_7544,N_3326,N_4610);
or U7545 (N_7545,N_3818,N_4016);
xor U7546 (N_7546,N_5047,N_5717);
nor U7547 (N_7547,N_5476,N_4566);
or U7548 (N_7548,N_5105,N_3615);
nor U7549 (N_7549,N_5576,N_5594);
nor U7550 (N_7550,N_4113,N_4454);
xnor U7551 (N_7551,N_5339,N_6191);
nor U7552 (N_7552,N_4136,N_5839);
or U7553 (N_7553,N_3457,N_5943);
and U7554 (N_7554,N_4620,N_4152);
and U7555 (N_7555,N_5685,N_4715);
xnor U7556 (N_7556,N_5620,N_4060);
nand U7557 (N_7557,N_6200,N_5946);
xnor U7558 (N_7558,N_5331,N_3331);
and U7559 (N_7559,N_4564,N_4181);
nand U7560 (N_7560,N_5450,N_3463);
nor U7561 (N_7561,N_6236,N_4183);
nand U7562 (N_7562,N_3833,N_5271);
and U7563 (N_7563,N_5510,N_3897);
xnor U7564 (N_7564,N_4381,N_3978);
nand U7565 (N_7565,N_5590,N_5817);
and U7566 (N_7566,N_5669,N_3750);
nor U7567 (N_7567,N_4319,N_3998);
nand U7568 (N_7568,N_4862,N_5872);
nor U7569 (N_7569,N_6096,N_5238);
and U7570 (N_7570,N_3276,N_5526);
nand U7571 (N_7571,N_3191,N_4774);
nand U7572 (N_7572,N_4141,N_5484);
nand U7573 (N_7573,N_4942,N_5444);
or U7574 (N_7574,N_3639,N_6152);
and U7575 (N_7575,N_4020,N_6118);
and U7576 (N_7576,N_5031,N_4660);
and U7577 (N_7577,N_5806,N_5187);
xor U7578 (N_7578,N_3142,N_4507);
nor U7579 (N_7579,N_5784,N_4810);
nor U7580 (N_7580,N_5399,N_6029);
nand U7581 (N_7581,N_4836,N_3402);
and U7582 (N_7582,N_5741,N_5063);
or U7583 (N_7583,N_3820,N_4274);
and U7584 (N_7584,N_5160,N_5818);
nor U7585 (N_7585,N_4124,N_3481);
and U7586 (N_7586,N_4149,N_5867);
xnor U7587 (N_7587,N_4290,N_4203);
nor U7588 (N_7588,N_6234,N_3726);
nor U7589 (N_7589,N_3713,N_4707);
nand U7590 (N_7590,N_3934,N_4577);
xnor U7591 (N_7591,N_5611,N_4746);
nor U7592 (N_7592,N_5728,N_3868);
and U7593 (N_7593,N_4250,N_3586);
nor U7594 (N_7594,N_6145,N_3186);
xor U7595 (N_7595,N_3658,N_5485);
and U7596 (N_7596,N_4027,N_3563);
nand U7597 (N_7597,N_5296,N_5901);
nand U7598 (N_7598,N_4330,N_5482);
nand U7599 (N_7599,N_3401,N_4949);
nor U7600 (N_7600,N_4695,N_6031);
or U7601 (N_7601,N_4895,N_5050);
nand U7602 (N_7602,N_5926,N_5328);
and U7603 (N_7603,N_4003,N_5001);
or U7604 (N_7604,N_4824,N_5360);
and U7605 (N_7605,N_6213,N_3602);
or U7606 (N_7606,N_5066,N_5431);
or U7607 (N_7607,N_3574,N_5826);
and U7608 (N_7608,N_4147,N_3816);
nand U7609 (N_7609,N_4099,N_5029);
xnor U7610 (N_7610,N_3912,N_4462);
nor U7611 (N_7611,N_4532,N_3329);
and U7612 (N_7612,N_5086,N_5178);
and U7613 (N_7613,N_5711,N_4502);
nor U7614 (N_7614,N_4404,N_4671);
nor U7615 (N_7615,N_4151,N_3690);
nor U7616 (N_7616,N_5117,N_5771);
nand U7617 (N_7617,N_3936,N_3496);
or U7618 (N_7618,N_4975,N_4675);
nand U7619 (N_7619,N_3860,N_4195);
nor U7620 (N_7620,N_5566,N_4698);
or U7621 (N_7621,N_4190,N_5230);
and U7622 (N_7622,N_3225,N_4318);
nand U7623 (N_7623,N_3715,N_4835);
or U7624 (N_7624,N_5396,N_5628);
xor U7625 (N_7625,N_3357,N_3349);
nand U7626 (N_7626,N_3671,N_6066);
nand U7627 (N_7627,N_5869,N_3493);
or U7628 (N_7628,N_3643,N_4708);
nand U7629 (N_7629,N_5033,N_6103);
or U7630 (N_7630,N_3341,N_5657);
nand U7631 (N_7631,N_3428,N_6220);
xor U7632 (N_7632,N_3538,N_4742);
and U7633 (N_7633,N_5773,N_3313);
nand U7634 (N_7634,N_5642,N_5604);
nor U7635 (N_7635,N_4081,N_5568);
and U7636 (N_7636,N_5503,N_3135);
nor U7637 (N_7637,N_5445,N_4277);
xor U7638 (N_7638,N_6219,N_5295);
nand U7639 (N_7639,N_6198,N_5758);
or U7640 (N_7640,N_5206,N_5714);
or U7641 (N_7641,N_4693,N_5964);
and U7642 (N_7642,N_3706,N_3559);
nor U7643 (N_7643,N_3625,N_5557);
or U7644 (N_7644,N_3939,N_4335);
and U7645 (N_7645,N_4232,N_3896);
xnor U7646 (N_7646,N_5200,N_6205);
nor U7647 (N_7647,N_4720,N_5645);
nand U7648 (N_7648,N_4249,N_3383);
xnor U7649 (N_7649,N_4043,N_4489);
xnor U7650 (N_7650,N_3446,N_5699);
nand U7651 (N_7651,N_5093,N_5055);
and U7652 (N_7652,N_3227,N_5183);
nand U7653 (N_7653,N_4626,N_3647);
nor U7654 (N_7654,N_5471,N_4456);
xnor U7655 (N_7655,N_5995,N_4448);
nand U7656 (N_7656,N_5601,N_4848);
and U7657 (N_7657,N_5730,N_4303);
nor U7658 (N_7658,N_3508,N_5918);
or U7659 (N_7659,N_4934,N_5194);
nor U7660 (N_7660,N_4239,N_4683);
nand U7661 (N_7661,N_4313,N_3228);
or U7662 (N_7662,N_3699,N_4518);
nand U7663 (N_7663,N_5036,N_3406);
and U7664 (N_7664,N_4850,N_5149);
nand U7665 (N_7665,N_4406,N_5455);
or U7666 (N_7666,N_3139,N_3964);
xor U7667 (N_7667,N_4790,N_3616);
nand U7668 (N_7668,N_3609,N_5304);
nand U7669 (N_7669,N_4729,N_5406);
nand U7670 (N_7670,N_4228,N_3635);
or U7671 (N_7671,N_4422,N_5341);
nand U7672 (N_7672,N_5021,N_4192);
xor U7673 (N_7673,N_3950,N_4911);
or U7674 (N_7674,N_5848,N_5342);
or U7675 (N_7675,N_3526,N_6195);
xor U7676 (N_7676,N_4750,N_3695);
nand U7677 (N_7677,N_4300,N_3989);
and U7678 (N_7678,N_3768,N_5618);
nand U7679 (N_7679,N_5437,N_5006);
nand U7680 (N_7680,N_5811,N_6169);
or U7681 (N_7681,N_6140,N_3709);
and U7682 (N_7682,N_5907,N_6215);
nor U7683 (N_7683,N_5933,N_5254);
nand U7684 (N_7684,N_4272,N_4188);
nor U7685 (N_7685,N_3852,N_3659);
and U7686 (N_7686,N_4646,N_4797);
nor U7687 (N_7687,N_3784,N_4943);
or U7688 (N_7688,N_4101,N_5821);
nand U7689 (N_7689,N_3855,N_4056);
and U7690 (N_7690,N_3180,N_5103);
xnor U7691 (N_7691,N_6064,N_4391);
nor U7692 (N_7692,N_5606,N_5713);
or U7693 (N_7693,N_5002,N_4561);
nor U7694 (N_7694,N_4028,N_3264);
or U7695 (N_7695,N_3128,N_6036);
xnor U7696 (N_7696,N_6233,N_4127);
nor U7697 (N_7697,N_4486,N_5300);
nand U7698 (N_7698,N_3577,N_3399);
or U7699 (N_7699,N_5433,N_5275);
nand U7700 (N_7700,N_5640,N_3448);
xnor U7701 (N_7701,N_3333,N_3825);
or U7702 (N_7702,N_3792,N_4463);
nor U7703 (N_7703,N_4172,N_4599);
and U7704 (N_7704,N_5749,N_4791);
nor U7705 (N_7705,N_5154,N_4673);
nand U7706 (N_7706,N_5040,N_5210);
and U7707 (N_7707,N_4981,N_5763);
nand U7708 (N_7708,N_6083,N_4684);
and U7709 (N_7709,N_5945,N_5680);
nand U7710 (N_7710,N_4559,N_5449);
nor U7711 (N_7711,N_3175,N_5558);
or U7712 (N_7712,N_4739,N_4173);
nor U7713 (N_7713,N_4207,N_3735);
nor U7714 (N_7714,N_5712,N_5423);
nor U7715 (N_7715,N_4965,N_5565);
and U7716 (N_7716,N_5458,N_4870);
nor U7717 (N_7717,N_4221,N_4495);
or U7718 (N_7718,N_3182,N_5572);
or U7719 (N_7719,N_3317,N_5874);
nor U7720 (N_7720,N_4252,N_5809);
and U7721 (N_7721,N_6110,N_5398);
or U7722 (N_7722,N_3947,N_5408);
and U7723 (N_7723,N_4086,N_3475);
nor U7724 (N_7724,N_4451,N_4521);
nand U7725 (N_7725,N_4236,N_4691);
nand U7726 (N_7726,N_3901,N_3867);
nand U7727 (N_7727,N_3763,N_5073);
nor U7728 (N_7728,N_4854,N_4658);
or U7729 (N_7729,N_5301,N_4840);
nor U7730 (N_7730,N_3275,N_3470);
nor U7731 (N_7731,N_6054,N_3778);
nand U7732 (N_7732,N_6116,N_5692);
xor U7733 (N_7733,N_3932,N_3741);
and U7734 (N_7734,N_5447,N_4703);
and U7735 (N_7735,N_3554,N_4259);
nand U7736 (N_7736,N_3437,N_4135);
nand U7737 (N_7737,N_4778,N_4058);
nand U7738 (N_7738,N_4088,N_5789);
or U7739 (N_7739,N_4825,N_4130);
nand U7740 (N_7740,N_4134,N_3272);
nor U7741 (N_7741,N_4896,N_5019);
nor U7742 (N_7742,N_4164,N_3502);
and U7743 (N_7743,N_3388,N_4478);
nand U7744 (N_7744,N_5299,N_4384);
nor U7745 (N_7745,N_4634,N_4938);
or U7746 (N_7746,N_5186,N_4402);
nand U7747 (N_7747,N_5859,N_5651);
nand U7748 (N_7748,N_3442,N_5395);
or U7749 (N_7749,N_5673,N_4414);
or U7750 (N_7750,N_6038,N_5975);
xnor U7751 (N_7751,N_5293,N_3767);
and U7752 (N_7752,N_3943,N_4666);
nand U7753 (N_7753,N_5630,N_5882);
xnor U7754 (N_7754,N_3342,N_4390);
or U7755 (N_7755,N_4980,N_3749);
nand U7756 (N_7756,N_5044,N_3736);
nor U7757 (N_7757,N_4198,N_3294);
nand U7758 (N_7758,N_4910,N_5076);
nand U7759 (N_7759,N_6211,N_4034);
and U7760 (N_7760,N_3390,N_3704);
nand U7761 (N_7761,N_4696,N_4504);
nand U7762 (N_7762,N_3440,N_5028);
or U7763 (N_7763,N_5142,N_3972);
and U7764 (N_7764,N_4142,N_4383);
nor U7765 (N_7765,N_4947,N_5794);
or U7766 (N_7766,N_3281,N_5225);
and U7767 (N_7767,N_5281,N_3542);
xor U7768 (N_7768,N_4717,N_3411);
nand U7769 (N_7769,N_4100,N_4552);
nand U7770 (N_7770,N_5264,N_5496);
and U7771 (N_7771,N_5245,N_3176);
or U7772 (N_7772,N_5650,N_3790);
nand U7773 (N_7773,N_5032,N_4307);
xnor U7774 (N_7774,N_5865,N_3392);
and U7775 (N_7775,N_4115,N_4220);
or U7776 (N_7776,N_4029,N_3396);
and U7777 (N_7777,N_4133,N_4244);
nand U7778 (N_7778,N_4363,N_4018);
nand U7779 (N_7779,N_5480,N_4317);
nor U7780 (N_7780,N_3394,N_5472);
or U7781 (N_7781,N_4464,N_3298);
and U7782 (N_7782,N_4377,N_5260);
nand U7783 (N_7783,N_4304,N_4573);
or U7784 (N_7784,N_3683,N_3849);
nand U7785 (N_7785,N_5106,N_5045);
and U7786 (N_7786,N_3798,N_5846);
and U7787 (N_7787,N_4452,N_5902);
or U7788 (N_7788,N_4311,N_5761);
or U7789 (N_7789,N_3556,N_5425);
nor U7790 (N_7790,N_3656,N_3696);
or U7791 (N_7791,N_6154,N_6183);
and U7792 (N_7792,N_3674,N_5085);
or U7793 (N_7793,N_4359,N_5724);
nand U7794 (N_7794,N_3663,N_4542);
and U7795 (N_7795,N_5780,N_5104);
or U7796 (N_7796,N_6048,N_5292);
or U7797 (N_7797,N_5856,N_5329);
xnor U7798 (N_7798,N_3229,N_4520);
nor U7799 (N_7799,N_3729,N_4904);
nor U7800 (N_7800,N_3760,N_4068);
and U7801 (N_7801,N_3354,N_5069);
nand U7802 (N_7802,N_5829,N_5988);
nand U7803 (N_7803,N_5802,N_3222);
and U7804 (N_7804,N_4649,N_3436);
xnor U7805 (N_7805,N_5390,N_4481);
and U7806 (N_7806,N_5949,N_4808);
nor U7807 (N_7807,N_5906,N_6177);
nand U7808 (N_7808,N_3471,N_3980);
nand U7809 (N_7809,N_5914,N_4428);
and U7810 (N_7810,N_5559,N_4168);
or U7811 (N_7811,N_4898,N_5693);
or U7812 (N_7812,N_4355,N_5483);
nor U7813 (N_7813,N_4093,N_3878);
or U7814 (N_7814,N_5489,N_4558);
and U7815 (N_7815,N_3892,N_3315);
nand U7816 (N_7816,N_4276,N_5475);
nor U7817 (N_7817,N_4848,N_5491);
nand U7818 (N_7818,N_4248,N_4263);
or U7819 (N_7819,N_4979,N_5723);
nor U7820 (N_7820,N_4081,N_4652);
nor U7821 (N_7821,N_5412,N_3611);
or U7822 (N_7822,N_3301,N_5763);
nand U7823 (N_7823,N_3237,N_3869);
and U7824 (N_7824,N_3264,N_5595);
or U7825 (N_7825,N_5176,N_5696);
nand U7826 (N_7826,N_3819,N_5779);
nor U7827 (N_7827,N_5412,N_4019);
xor U7828 (N_7828,N_4078,N_3826);
xor U7829 (N_7829,N_4848,N_4563);
nor U7830 (N_7830,N_5498,N_5595);
nand U7831 (N_7831,N_4251,N_6145);
or U7832 (N_7832,N_4638,N_4193);
and U7833 (N_7833,N_5992,N_4751);
and U7834 (N_7834,N_5360,N_3839);
or U7835 (N_7835,N_3352,N_6068);
and U7836 (N_7836,N_4767,N_3713);
xnor U7837 (N_7837,N_5864,N_4509);
or U7838 (N_7838,N_4369,N_5581);
nand U7839 (N_7839,N_3897,N_3911);
xnor U7840 (N_7840,N_4311,N_4437);
nor U7841 (N_7841,N_5928,N_5423);
nor U7842 (N_7842,N_5805,N_4957);
and U7843 (N_7843,N_3261,N_6002);
nor U7844 (N_7844,N_4296,N_3998);
and U7845 (N_7845,N_6037,N_4123);
and U7846 (N_7846,N_5039,N_4570);
or U7847 (N_7847,N_5536,N_3932);
nor U7848 (N_7848,N_5910,N_4963);
or U7849 (N_7849,N_5891,N_3914);
nor U7850 (N_7850,N_3968,N_3922);
and U7851 (N_7851,N_3838,N_4128);
nand U7852 (N_7852,N_4610,N_4866);
nor U7853 (N_7853,N_4109,N_3306);
or U7854 (N_7854,N_4150,N_6241);
nor U7855 (N_7855,N_5172,N_3347);
or U7856 (N_7856,N_4766,N_4597);
and U7857 (N_7857,N_5254,N_3826);
and U7858 (N_7858,N_6246,N_5799);
nor U7859 (N_7859,N_3509,N_5751);
nand U7860 (N_7860,N_4265,N_4207);
nor U7861 (N_7861,N_3410,N_4419);
or U7862 (N_7862,N_5483,N_4779);
nand U7863 (N_7863,N_4333,N_5389);
and U7864 (N_7864,N_4075,N_5518);
nor U7865 (N_7865,N_5071,N_6001);
and U7866 (N_7866,N_4876,N_3997);
nand U7867 (N_7867,N_4753,N_3648);
and U7868 (N_7868,N_5283,N_4467);
nor U7869 (N_7869,N_3757,N_4381);
or U7870 (N_7870,N_5328,N_5748);
nand U7871 (N_7871,N_5559,N_5554);
or U7872 (N_7872,N_6157,N_4391);
or U7873 (N_7873,N_4872,N_3159);
and U7874 (N_7874,N_3568,N_5017);
nand U7875 (N_7875,N_5337,N_3508);
xor U7876 (N_7876,N_3653,N_5031);
and U7877 (N_7877,N_4907,N_3339);
and U7878 (N_7878,N_5328,N_6083);
nand U7879 (N_7879,N_3736,N_4654);
or U7880 (N_7880,N_5497,N_4353);
and U7881 (N_7881,N_3297,N_4631);
and U7882 (N_7882,N_5065,N_3897);
and U7883 (N_7883,N_4569,N_3794);
xor U7884 (N_7884,N_3691,N_4338);
nand U7885 (N_7885,N_5444,N_4951);
and U7886 (N_7886,N_4144,N_5072);
and U7887 (N_7887,N_3699,N_6093);
and U7888 (N_7888,N_3367,N_4881);
nand U7889 (N_7889,N_3364,N_5941);
nand U7890 (N_7890,N_4997,N_3881);
xor U7891 (N_7891,N_3540,N_4304);
and U7892 (N_7892,N_3459,N_5753);
and U7893 (N_7893,N_3825,N_5464);
nor U7894 (N_7894,N_4018,N_3698);
or U7895 (N_7895,N_5307,N_5021);
nor U7896 (N_7896,N_5180,N_5839);
or U7897 (N_7897,N_3446,N_6006);
nor U7898 (N_7898,N_6170,N_3436);
nand U7899 (N_7899,N_4813,N_5218);
nand U7900 (N_7900,N_4027,N_5124);
and U7901 (N_7901,N_5303,N_3589);
nand U7902 (N_7902,N_6032,N_5261);
nor U7903 (N_7903,N_3483,N_3721);
xnor U7904 (N_7904,N_4178,N_6098);
or U7905 (N_7905,N_3606,N_5115);
nor U7906 (N_7906,N_5585,N_3609);
nand U7907 (N_7907,N_5116,N_5966);
xnor U7908 (N_7908,N_4838,N_3609);
nor U7909 (N_7909,N_3704,N_4581);
nand U7910 (N_7910,N_4240,N_5801);
nor U7911 (N_7911,N_6142,N_5509);
and U7912 (N_7912,N_3480,N_4740);
and U7913 (N_7913,N_5021,N_5263);
nand U7914 (N_7914,N_6130,N_4355);
xnor U7915 (N_7915,N_4998,N_4799);
or U7916 (N_7916,N_4232,N_4945);
and U7917 (N_7917,N_5850,N_3394);
or U7918 (N_7918,N_5104,N_5134);
or U7919 (N_7919,N_4539,N_5349);
and U7920 (N_7920,N_3641,N_4737);
and U7921 (N_7921,N_6128,N_4019);
or U7922 (N_7922,N_4815,N_4042);
nand U7923 (N_7923,N_5133,N_3509);
nor U7924 (N_7924,N_5664,N_6062);
or U7925 (N_7925,N_3149,N_5387);
and U7926 (N_7926,N_4725,N_3206);
xor U7927 (N_7927,N_5197,N_4380);
or U7928 (N_7928,N_5350,N_4288);
or U7929 (N_7929,N_3688,N_5218);
nor U7930 (N_7930,N_5133,N_5811);
nand U7931 (N_7931,N_5725,N_5716);
or U7932 (N_7932,N_4271,N_6139);
or U7933 (N_7933,N_4047,N_6178);
nor U7934 (N_7934,N_4319,N_5717);
nor U7935 (N_7935,N_3676,N_3828);
nand U7936 (N_7936,N_5895,N_5167);
and U7937 (N_7937,N_3512,N_4150);
nor U7938 (N_7938,N_3354,N_4808);
xor U7939 (N_7939,N_3669,N_3240);
nand U7940 (N_7940,N_5013,N_4342);
nand U7941 (N_7941,N_6171,N_3209);
nand U7942 (N_7942,N_5371,N_5980);
nand U7943 (N_7943,N_4337,N_3616);
nand U7944 (N_7944,N_4351,N_3364);
nor U7945 (N_7945,N_3785,N_5403);
and U7946 (N_7946,N_5967,N_5720);
and U7947 (N_7947,N_4787,N_6179);
xor U7948 (N_7948,N_3423,N_6247);
nand U7949 (N_7949,N_4185,N_5668);
and U7950 (N_7950,N_3709,N_4271);
and U7951 (N_7951,N_5968,N_5217);
xnor U7952 (N_7952,N_3871,N_4751);
nor U7953 (N_7953,N_5698,N_5222);
nand U7954 (N_7954,N_6234,N_6020);
nand U7955 (N_7955,N_4149,N_4825);
or U7956 (N_7956,N_5208,N_4501);
nand U7957 (N_7957,N_4814,N_4474);
nor U7958 (N_7958,N_5544,N_5387);
nor U7959 (N_7959,N_3267,N_3258);
or U7960 (N_7960,N_5929,N_3159);
nor U7961 (N_7961,N_4183,N_3185);
nand U7962 (N_7962,N_3832,N_3418);
or U7963 (N_7963,N_5471,N_3823);
or U7964 (N_7964,N_4821,N_3466);
nand U7965 (N_7965,N_5129,N_5223);
nor U7966 (N_7966,N_6179,N_4386);
and U7967 (N_7967,N_5559,N_5716);
nand U7968 (N_7968,N_4332,N_4564);
nor U7969 (N_7969,N_3392,N_4964);
or U7970 (N_7970,N_4521,N_3547);
nand U7971 (N_7971,N_3691,N_3367);
or U7972 (N_7972,N_5799,N_3842);
nand U7973 (N_7973,N_3847,N_3417);
or U7974 (N_7974,N_4015,N_5621);
and U7975 (N_7975,N_3553,N_3548);
and U7976 (N_7976,N_3240,N_3463);
or U7977 (N_7977,N_3220,N_3171);
and U7978 (N_7978,N_3260,N_5569);
or U7979 (N_7979,N_5965,N_5239);
or U7980 (N_7980,N_3399,N_3136);
nor U7981 (N_7981,N_4823,N_4283);
nand U7982 (N_7982,N_4266,N_4510);
or U7983 (N_7983,N_3376,N_4661);
and U7984 (N_7984,N_3662,N_3470);
and U7985 (N_7985,N_3549,N_5089);
nor U7986 (N_7986,N_3586,N_3999);
or U7987 (N_7987,N_4356,N_5875);
and U7988 (N_7988,N_5866,N_3282);
xor U7989 (N_7989,N_5028,N_4249);
and U7990 (N_7990,N_3946,N_5947);
and U7991 (N_7991,N_4821,N_4946);
or U7992 (N_7992,N_4873,N_4772);
nand U7993 (N_7993,N_3203,N_6028);
xnor U7994 (N_7994,N_3295,N_6144);
and U7995 (N_7995,N_3286,N_3946);
xor U7996 (N_7996,N_4606,N_3331);
nand U7997 (N_7997,N_5237,N_4709);
or U7998 (N_7998,N_6125,N_5142);
nor U7999 (N_7999,N_5579,N_4736);
xnor U8000 (N_8000,N_5326,N_4968);
nor U8001 (N_8001,N_6062,N_4927);
xor U8002 (N_8002,N_6143,N_3138);
and U8003 (N_8003,N_5682,N_3989);
xor U8004 (N_8004,N_5091,N_6059);
nand U8005 (N_8005,N_3218,N_3901);
and U8006 (N_8006,N_4080,N_3325);
or U8007 (N_8007,N_3914,N_4636);
or U8008 (N_8008,N_5649,N_5448);
nor U8009 (N_8009,N_3303,N_3219);
nor U8010 (N_8010,N_3626,N_4410);
nand U8011 (N_8011,N_4720,N_5352);
and U8012 (N_8012,N_5403,N_4029);
or U8013 (N_8013,N_5106,N_3686);
or U8014 (N_8014,N_4072,N_4841);
nand U8015 (N_8015,N_4436,N_5321);
nand U8016 (N_8016,N_5803,N_4612);
and U8017 (N_8017,N_4335,N_3835);
nor U8018 (N_8018,N_5590,N_5350);
and U8019 (N_8019,N_4002,N_3488);
nor U8020 (N_8020,N_3257,N_4277);
and U8021 (N_8021,N_3345,N_4030);
and U8022 (N_8022,N_3570,N_3802);
nor U8023 (N_8023,N_5744,N_5614);
and U8024 (N_8024,N_3551,N_4020);
xor U8025 (N_8025,N_3858,N_4638);
nor U8026 (N_8026,N_5496,N_4085);
nand U8027 (N_8027,N_3572,N_4702);
and U8028 (N_8028,N_5012,N_3480);
and U8029 (N_8029,N_4356,N_4870);
or U8030 (N_8030,N_3251,N_5742);
and U8031 (N_8031,N_4721,N_3886);
or U8032 (N_8032,N_4690,N_5429);
or U8033 (N_8033,N_5465,N_4404);
or U8034 (N_8034,N_3533,N_4035);
or U8035 (N_8035,N_3252,N_4960);
or U8036 (N_8036,N_3534,N_4525);
xnor U8037 (N_8037,N_3515,N_5520);
and U8038 (N_8038,N_5338,N_4983);
xor U8039 (N_8039,N_6131,N_3734);
xor U8040 (N_8040,N_4296,N_3792);
nor U8041 (N_8041,N_4822,N_6176);
xor U8042 (N_8042,N_4811,N_5900);
and U8043 (N_8043,N_4695,N_5260);
and U8044 (N_8044,N_4789,N_3769);
nor U8045 (N_8045,N_3861,N_4936);
nor U8046 (N_8046,N_3151,N_5359);
nor U8047 (N_8047,N_3345,N_5238);
nand U8048 (N_8048,N_5770,N_4900);
or U8049 (N_8049,N_4043,N_5729);
nand U8050 (N_8050,N_4884,N_5156);
nor U8051 (N_8051,N_3799,N_5100);
nand U8052 (N_8052,N_3291,N_3736);
xor U8053 (N_8053,N_5057,N_5736);
and U8054 (N_8054,N_4604,N_5838);
nor U8055 (N_8055,N_4515,N_3190);
nand U8056 (N_8056,N_4974,N_5789);
or U8057 (N_8057,N_4296,N_5041);
or U8058 (N_8058,N_3197,N_4259);
nand U8059 (N_8059,N_5154,N_5637);
or U8060 (N_8060,N_5298,N_4823);
or U8061 (N_8061,N_3863,N_5600);
xor U8062 (N_8062,N_5515,N_4606);
and U8063 (N_8063,N_5479,N_5960);
nand U8064 (N_8064,N_6181,N_6153);
xor U8065 (N_8065,N_4449,N_3716);
and U8066 (N_8066,N_5315,N_6136);
nor U8067 (N_8067,N_4903,N_6225);
or U8068 (N_8068,N_3830,N_4793);
or U8069 (N_8069,N_3154,N_3772);
or U8070 (N_8070,N_5947,N_3790);
or U8071 (N_8071,N_5250,N_5052);
or U8072 (N_8072,N_5596,N_4438);
nor U8073 (N_8073,N_4747,N_5934);
and U8074 (N_8074,N_4329,N_5973);
xor U8075 (N_8075,N_5974,N_5734);
or U8076 (N_8076,N_3534,N_3888);
nor U8077 (N_8077,N_3133,N_4791);
nor U8078 (N_8078,N_5953,N_5454);
nor U8079 (N_8079,N_6059,N_4665);
nand U8080 (N_8080,N_4073,N_6183);
nand U8081 (N_8081,N_5767,N_5466);
or U8082 (N_8082,N_5450,N_5860);
nand U8083 (N_8083,N_5621,N_3127);
or U8084 (N_8084,N_4988,N_3144);
and U8085 (N_8085,N_5750,N_3457);
nand U8086 (N_8086,N_3354,N_4143);
nor U8087 (N_8087,N_5803,N_4937);
or U8088 (N_8088,N_5185,N_6103);
or U8089 (N_8089,N_5725,N_4754);
nor U8090 (N_8090,N_3927,N_5106);
and U8091 (N_8091,N_4699,N_4917);
xor U8092 (N_8092,N_5989,N_3901);
or U8093 (N_8093,N_4396,N_3941);
nand U8094 (N_8094,N_5671,N_5444);
nand U8095 (N_8095,N_4522,N_5222);
or U8096 (N_8096,N_5656,N_4648);
nor U8097 (N_8097,N_6028,N_5487);
nand U8098 (N_8098,N_5154,N_5405);
or U8099 (N_8099,N_3825,N_4346);
xor U8100 (N_8100,N_3127,N_5590);
and U8101 (N_8101,N_4572,N_3316);
nand U8102 (N_8102,N_4440,N_3801);
or U8103 (N_8103,N_3643,N_4585);
or U8104 (N_8104,N_5455,N_3590);
nor U8105 (N_8105,N_3850,N_3213);
or U8106 (N_8106,N_4423,N_6186);
xnor U8107 (N_8107,N_5529,N_3435);
or U8108 (N_8108,N_3882,N_5116);
nand U8109 (N_8109,N_5593,N_4546);
nor U8110 (N_8110,N_3456,N_5581);
and U8111 (N_8111,N_5663,N_5260);
or U8112 (N_8112,N_5552,N_5521);
and U8113 (N_8113,N_5784,N_3350);
or U8114 (N_8114,N_4628,N_4637);
nand U8115 (N_8115,N_3537,N_5402);
nor U8116 (N_8116,N_5439,N_5397);
nor U8117 (N_8117,N_5947,N_3453);
or U8118 (N_8118,N_3372,N_3965);
nor U8119 (N_8119,N_3638,N_3861);
nor U8120 (N_8120,N_3712,N_5731);
nand U8121 (N_8121,N_6096,N_4373);
xnor U8122 (N_8122,N_5744,N_4010);
nand U8123 (N_8123,N_4718,N_3981);
nand U8124 (N_8124,N_5739,N_5423);
or U8125 (N_8125,N_5889,N_3410);
nand U8126 (N_8126,N_5004,N_3890);
nand U8127 (N_8127,N_4310,N_3613);
xor U8128 (N_8128,N_5516,N_3816);
nor U8129 (N_8129,N_3376,N_3259);
or U8130 (N_8130,N_3770,N_3673);
nor U8131 (N_8131,N_5171,N_3514);
or U8132 (N_8132,N_5588,N_4088);
nand U8133 (N_8133,N_4147,N_5128);
xnor U8134 (N_8134,N_5875,N_4056);
nor U8135 (N_8135,N_3591,N_4501);
nor U8136 (N_8136,N_4566,N_4795);
nand U8137 (N_8137,N_4058,N_5564);
and U8138 (N_8138,N_5754,N_5215);
nand U8139 (N_8139,N_4559,N_5094);
nor U8140 (N_8140,N_3381,N_3157);
xnor U8141 (N_8141,N_6044,N_6204);
or U8142 (N_8142,N_5748,N_6016);
nor U8143 (N_8143,N_4405,N_3308);
nand U8144 (N_8144,N_4056,N_3657);
and U8145 (N_8145,N_4935,N_4017);
nor U8146 (N_8146,N_5866,N_3914);
or U8147 (N_8147,N_5304,N_4353);
and U8148 (N_8148,N_5894,N_4298);
and U8149 (N_8149,N_4670,N_3169);
and U8150 (N_8150,N_5433,N_5844);
and U8151 (N_8151,N_3752,N_3218);
nand U8152 (N_8152,N_5071,N_3589);
or U8153 (N_8153,N_5284,N_4028);
nand U8154 (N_8154,N_5708,N_4165);
or U8155 (N_8155,N_4991,N_4015);
or U8156 (N_8156,N_5129,N_3349);
and U8157 (N_8157,N_5609,N_3741);
or U8158 (N_8158,N_4900,N_3336);
nand U8159 (N_8159,N_5210,N_6177);
nor U8160 (N_8160,N_3597,N_6079);
nand U8161 (N_8161,N_5674,N_3599);
nand U8162 (N_8162,N_5336,N_4202);
nor U8163 (N_8163,N_5283,N_4529);
nor U8164 (N_8164,N_5681,N_4436);
nand U8165 (N_8165,N_4597,N_4909);
or U8166 (N_8166,N_3238,N_4084);
or U8167 (N_8167,N_5675,N_5288);
or U8168 (N_8168,N_3898,N_4988);
nor U8169 (N_8169,N_6057,N_3501);
and U8170 (N_8170,N_5853,N_5545);
xor U8171 (N_8171,N_5903,N_4692);
or U8172 (N_8172,N_4823,N_4391);
and U8173 (N_8173,N_6027,N_5266);
nor U8174 (N_8174,N_6055,N_4971);
and U8175 (N_8175,N_4943,N_5472);
or U8176 (N_8176,N_5209,N_5224);
and U8177 (N_8177,N_3453,N_3737);
nor U8178 (N_8178,N_4324,N_5313);
xor U8179 (N_8179,N_3669,N_6052);
and U8180 (N_8180,N_5448,N_4569);
and U8181 (N_8181,N_5940,N_3622);
and U8182 (N_8182,N_3440,N_5133);
nand U8183 (N_8183,N_4904,N_3350);
xor U8184 (N_8184,N_5431,N_5364);
or U8185 (N_8185,N_5621,N_3635);
and U8186 (N_8186,N_3504,N_5535);
nor U8187 (N_8187,N_3824,N_4899);
or U8188 (N_8188,N_5945,N_5452);
nand U8189 (N_8189,N_3714,N_3618);
and U8190 (N_8190,N_5588,N_5268);
xnor U8191 (N_8191,N_4543,N_5947);
or U8192 (N_8192,N_4230,N_4508);
and U8193 (N_8193,N_3879,N_4859);
nor U8194 (N_8194,N_4080,N_5798);
and U8195 (N_8195,N_3791,N_5389);
and U8196 (N_8196,N_3302,N_3479);
or U8197 (N_8197,N_4601,N_4481);
or U8198 (N_8198,N_3962,N_4001);
nor U8199 (N_8199,N_3902,N_5048);
nor U8200 (N_8200,N_4092,N_5364);
nand U8201 (N_8201,N_5228,N_4988);
nand U8202 (N_8202,N_3275,N_5186);
or U8203 (N_8203,N_5753,N_3618);
and U8204 (N_8204,N_3125,N_5854);
or U8205 (N_8205,N_4477,N_3400);
nor U8206 (N_8206,N_3606,N_5163);
nand U8207 (N_8207,N_3827,N_4816);
nor U8208 (N_8208,N_4025,N_3667);
nor U8209 (N_8209,N_3396,N_5750);
nor U8210 (N_8210,N_5287,N_5128);
or U8211 (N_8211,N_5565,N_5386);
xnor U8212 (N_8212,N_5962,N_4330);
xor U8213 (N_8213,N_3201,N_5816);
and U8214 (N_8214,N_3723,N_4849);
nor U8215 (N_8215,N_5475,N_3289);
and U8216 (N_8216,N_5070,N_3724);
xnor U8217 (N_8217,N_5677,N_3511);
nand U8218 (N_8218,N_5697,N_5403);
or U8219 (N_8219,N_4968,N_3840);
and U8220 (N_8220,N_5041,N_3347);
nand U8221 (N_8221,N_6133,N_3237);
nor U8222 (N_8222,N_4275,N_4357);
nor U8223 (N_8223,N_4615,N_4518);
and U8224 (N_8224,N_4179,N_4096);
nand U8225 (N_8225,N_3574,N_5890);
or U8226 (N_8226,N_6130,N_5745);
and U8227 (N_8227,N_5975,N_4136);
nand U8228 (N_8228,N_3402,N_4172);
or U8229 (N_8229,N_4054,N_3762);
nand U8230 (N_8230,N_5431,N_3549);
and U8231 (N_8231,N_3924,N_3421);
nand U8232 (N_8232,N_3989,N_5534);
nand U8233 (N_8233,N_5825,N_3541);
nand U8234 (N_8234,N_4854,N_5173);
nand U8235 (N_8235,N_6120,N_5019);
nor U8236 (N_8236,N_4747,N_3308);
and U8237 (N_8237,N_5865,N_4320);
or U8238 (N_8238,N_5050,N_5793);
and U8239 (N_8239,N_5461,N_4401);
nor U8240 (N_8240,N_3234,N_5995);
and U8241 (N_8241,N_5392,N_5138);
nand U8242 (N_8242,N_4546,N_3667);
nor U8243 (N_8243,N_3968,N_4360);
or U8244 (N_8244,N_4299,N_3720);
and U8245 (N_8245,N_5735,N_5070);
nand U8246 (N_8246,N_4980,N_5712);
nor U8247 (N_8247,N_3754,N_4979);
and U8248 (N_8248,N_4516,N_5917);
and U8249 (N_8249,N_3180,N_5501);
nor U8250 (N_8250,N_5959,N_5181);
or U8251 (N_8251,N_3308,N_3360);
nand U8252 (N_8252,N_5271,N_4311);
or U8253 (N_8253,N_3573,N_4560);
nand U8254 (N_8254,N_3671,N_4646);
nor U8255 (N_8255,N_5368,N_3886);
nand U8256 (N_8256,N_4181,N_3429);
and U8257 (N_8257,N_4167,N_4135);
nor U8258 (N_8258,N_3306,N_4679);
and U8259 (N_8259,N_3640,N_4764);
nand U8260 (N_8260,N_4725,N_6026);
nand U8261 (N_8261,N_6193,N_5384);
or U8262 (N_8262,N_4431,N_3585);
nand U8263 (N_8263,N_5888,N_5500);
and U8264 (N_8264,N_3419,N_4744);
and U8265 (N_8265,N_3551,N_5994);
nor U8266 (N_8266,N_6175,N_5450);
nor U8267 (N_8267,N_6117,N_3171);
or U8268 (N_8268,N_5584,N_5913);
or U8269 (N_8269,N_5190,N_4057);
nor U8270 (N_8270,N_4643,N_3331);
or U8271 (N_8271,N_5054,N_4997);
xnor U8272 (N_8272,N_5567,N_5533);
and U8273 (N_8273,N_3615,N_3898);
nor U8274 (N_8274,N_4860,N_3226);
and U8275 (N_8275,N_3383,N_3626);
and U8276 (N_8276,N_3565,N_4473);
or U8277 (N_8277,N_6040,N_6160);
or U8278 (N_8278,N_4326,N_4674);
xnor U8279 (N_8279,N_3494,N_4790);
or U8280 (N_8280,N_5299,N_3644);
or U8281 (N_8281,N_5940,N_5747);
nor U8282 (N_8282,N_3172,N_4088);
nand U8283 (N_8283,N_6056,N_5790);
or U8284 (N_8284,N_5015,N_3804);
nor U8285 (N_8285,N_5430,N_5029);
and U8286 (N_8286,N_4632,N_6006);
or U8287 (N_8287,N_4077,N_4425);
nor U8288 (N_8288,N_3902,N_3832);
nand U8289 (N_8289,N_3736,N_5641);
nand U8290 (N_8290,N_5519,N_5170);
or U8291 (N_8291,N_4384,N_4582);
xnor U8292 (N_8292,N_4314,N_4834);
or U8293 (N_8293,N_5130,N_6088);
or U8294 (N_8294,N_3565,N_5852);
nor U8295 (N_8295,N_5553,N_4986);
or U8296 (N_8296,N_4836,N_4594);
or U8297 (N_8297,N_5275,N_5644);
nor U8298 (N_8298,N_4028,N_5504);
nor U8299 (N_8299,N_4761,N_5403);
and U8300 (N_8300,N_5471,N_4905);
and U8301 (N_8301,N_3659,N_5803);
nand U8302 (N_8302,N_3567,N_3783);
and U8303 (N_8303,N_4494,N_4192);
or U8304 (N_8304,N_4176,N_5752);
nor U8305 (N_8305,N_4297,N_5792);
and U8306 (N_8306,N_4324,N_4258);
nor U8307 (N_8307,N_4229,N_5908);
nand U8308 (N_8308,N_4946,N_3784);
and U8309 (N_8309,N_4316,N_3468);
nor U8310 (N_8310,N_4582,N_3266);
and U8311 (N_8311,N_5448,N_3379);
or U8312 (N_8312,N_6031,N_5170);
and U8313 (N_8313,N_4250,N_4213);
nand U8314 (N_8314,N_5649,N_5828);
or U8315 (N_8315,N_4348,N_5443);
nand U8316 (N_8316,N_3655,N_5287);
nor U8317 (N_8317,N_3184,N_4028);
nor U8318 (N_8318,N_4744,N_3655);
and U8319 (N_8319,N_4264,N_5025);
nor U8320 (N_8320,N_6147,N_5913);
or U8321 (N_8321,N_3551,N_5424);
and U8322 (N_8322,N_4063,N_4392);
nor U8323 (N_8323,N_3584,N_4876);
nand U8324 (N_8324,N_4288,N_4220);
or U8325 (N_8325,N_3294,N_6178);
nand U8326 (N_8326,N_3212,N_3568);
and U8327 (N_8327,N_5920,N_5745);
nand U8328 (N_8328,N_4643,N_5024);
nand U8329 (N_8329,N_6005,N_4893);
nand U8330 (N_8330,N_5881,N_4694);
nand U8331 (N_8331,N_3575,N_3182);
and U8332 (N_8332,N_5471,N_5373);
or U8333 (N_8333,N_5398,N_5408);
or U8334 (N_8334,N_4634,N_4088);
nor U8335 (N_8335,N_4883,N_6189);
or U8336 (N_8336,N_5266,N_5890);
and U8337 (N_8337,N_3312,N_5148);
nor U8338 (N_8338,N_4803,N_3485);
nand U8339 (N_8339,N_3673,N_3528);
and U8340 (N_8340,N_3969,N_4143);
nor U8341 (N_8341,N_5546,N_4082);
or U8342 (N_8342,N_3820,N_4580);
or U8343 (N_8343,N_3646,N_6216);
nand U8344 (N_8344,N_4248,N_5713);
or U8345 (N_8345,N_5335,N_6081);
or U8346 (N_8346,N_5977,N_5086);
nor U8347 (N_8347,N_3598,N_3963);
or U8348 (N_8348,N_5780,N_4661);
nand U8349 (N_8349,N_5722,N_3482);
xor U8350 (N_8350,N_4682,N_5150);
and U8351 (N_8351,N_3904,N_3630);
and U8352 (N_8352,N_5518,N_3356);
or U8353 (N_8353,N_3246,N_4443);
nor U8354 (N_8354,N_4700,N_3758);
nor U8355 (N_8355,N_3195,N_3553);
or U8356 (N_8356,N_3344,N_3137);
or U8357 (N_8357,N_5690,N_3776);
and U8358 (N_8358,N_3535,N_4911);
and U8359 (N_8359,N_5953,N_3687);
nor U8360 (N_8360,N_3179,N_5891);
or U8361 (N_8361,N_5604,N_4585);
and U8362 (N_8362,N_5455,N_3173);
or U8363 (N_8363,N_3426,N_4787);
and U8364 (N_8364,N_3944,N_3140);
xnor U8365 (N_8365,N_4398,N_5818);
or U8366 (N_8366,N_4787,N_5949);
nand U8367 (N_8367,N_4094,N_6118);
nand U8368 (N_8368,N_5728,N_3845);
xnor U8369 (N_8369,N_5571,N_6190);
xor U8370 (N_8370,N_6164,N_3915);
or U8371 (N_8371,N_3586,N_5719);
or U8372 (N_8372,N_6038,N_3393);
nand U8373 (N_8373,N_3586,N_4134);
nor U8374 (N_8374,N_6077,N_3580);
nor U8375 (N_8375,N_5520,N_5105);
and U8376 (N_8376,N_3758,N_3315);
nor U8377 (N_8377,N_4073,N_5053);
nor U8378 (N_8378,N_4124,N_6209);
xnor U8379 (N_8379,N_5036,N_5532);
nor U8380 (N_8380,N_5504,N_3152);
nand U8381 (N_8381,N_4006,N_4793);
nand U8382 (N_8382,N_3511,N_3159);
and U8383 (N_8383,N_4506,N_5504);
nor U8384 (N_8384,N_5706,N_3775);
or U8385 (N_8385,N_4030,N_5964);
and U8386 (N_8386,N_5037,N_5326);
xnor U8387 (N_8387,N_5148,N_5991);
xnor U8388 (N_8388,N_5966,N_4832);
xnor U8389 (N_8389,N_4195,N_3973);
and U8390 (N_8390,N_4195,N_4894);
nand U8391 (N_8391,N_5001,N_5515);
nor U8392 (N_8392,N_5603,N_4272);
or U8393 (N_8393,N_5960,N_3849);
nor U8394 (N_8394,N_3843,N_6037);
or U8395 (N_8395,N_4377,N_4209);
and U8396 (N_8396,N_6007,N_5610);
nand U8397 (N_8397,N_5386,N_6098);
nor U8398 (N_8398,N_5872,N_4892);
xnor U8399 (N_8399,N_6176,N_4455);
and U8400 (N_8400,N_6087,N_6197);
and U8401 (N_8401,N_4786,N_4498);
xor U8402 (N_8402,N_3521,N_3248);
xor U8403 (N_8403,N_3849,N_3528);
and U8404 (N_8404,N_3912,N_4605);
and U8405 (N_8405,N_3930,N_5393);
nand U8406 (N_8406,N_4465,N_4559);
or U8407 (N_8407,N_4709,N_3383);
and U8408 (N_8408,N_4131,N_6144);
xor U8409 (N_8409,N_5826,N_5276);
and U8410 (N_8410,N_3855,N_5121);
and U8411 (N_8411,N_5420,N_6145);
xnor U8412 (N_8412,N_4835,N_5158);
xor U8413 (N_8413,N_3617,N_5814);
or U8414 (N_8414,N_3710,N_5457);
and U8415 (N_8415,N_3356,N_5029);
nand U8416 (N_8416,N_3985,N_3647);
and U8417 (N_8417,N_4170,N_4457);
xnor U8418 (N_8418,N_4058,N_5754);
nand U8419 (N_8419,N_4442,N_6208);
and U8420 (N_8420,N_6110,N_5803);
and U8421 (N_8421,N_4268,N_4378);
or U8422 (N_8422,N_5981,N_5387);
or U8423 (N_8423,N_5225,N_5490);
and U8424 (N_8424,N_5351,N_4547);
and U8425 (N_8425,N_5421,N_4798);
nor U8426 (N_8426,N_4433,N_4455);
xor U8427 (N_8427,N_4831,N_5259);
or U8428 (N_8428,N_4493,N_4644);
xor U8429 (N_8429,N_3871,N_3718);
nand U8430 (N_8430,N_3533,N_5073);
or U8431 (N_8431,N_5628,N_3680);
or U8432 (N_8432,N_5364,N_6024);
or U8433 (N_8433,N_4999,N_4458);
nand U8434 (N_8434,N_4989,N_3899);
nand U8435 (N_8435,N_3432,N_5416);
nand U8436 (N_8436,N_6210,N_4172);
nand U8437 (N_8437,N_3698,N_4924);
or U8438 (N_8438,N_6138,N_4644);
or U8439 (N_8439,N_3468,N_4737);
nor U8440 (N_8440,N_3527,N_5268);
xnor U8441 (N_8441,N_4226,N_5903);
or U8442 (N_8442,N_6174,N_3461);
nand U8443 (N_8443,N_4621,N_6135);
nand U8444 (N_8444,N_3199,N_4024);
or U8445 (N_8445,N_6131,N_3305);
nand U8446 (N_8446,N_4853,N_3850);
or U8447 (N_8447,N_4043,N_3530);
nand U8448 (N_8448,N_4968,N_4419);
or U8449 (N_8449,N_4409,N_5030);
and U8450 (N_8450,N_5849,N_5532);
nand U8451 (N_8451,N_6069,N_3840);
nor U8452 (N_8452,N_4773,N_5902);
nand U8453 (N_8453,N_5290,N_6060);
or U8454 (N_8454,N_4372,N_4055);
or U8455 (N_8455,N_4592,N_4301);
xor U8456 (N_8456,N_3511,N_4111);
nor U8457 (N_8457,N_4845,N_4685);
nor U8458 (N_8458,N_5552,N_3607);
nand U8459 (N_8459,N_6105,N_4545);
or U8460 (N_8460,N_4355,N_5369);
nor U8461 (N_8461,N_3563,N_5618);
or U8462 (N_8462,N_4616,N_5777);
nand U8463 (N_8463,N_4835,N_4701);
nor U8464 (N_8464,N_5006,N_4688);
xor U8465 (N_8465,N_5144,N_4013);
and U8466 (N_8466,N_4295,N_3705);
and U8467 (N_8467,N_4217,N_4946);
and U8468 (N_8468,N_4164,N_5212);
and U8469 (N_8469,N_4341,N_4633);
nand U8470 (N_8470,N_4341,N_3691);
and U8471 (N_8471,N_4685,N_4784);
nor U8472 (N_8472,N_5613,N_5099);
xnor U8473 (N_8473,N_5286,N_6220);
nand U8474 (N_8474,N_5212,N_5096);
nand U8475 (N_8475,N_6098,N_5417);
nor U8476 (N_8476,N_4321,N_3863);
or U8477 (N_8477,N_3345,N_4254);
nor U8478 (N_8478,N_5889,N_5287);
nand U8479 (N_8479,N_5735,N_5578);
and U8480 (N_8480,N_5176,N_4445);
and U8481 (N_8481,N_5715,N_3774);
nor U8482 (N_8482,N_5120,N_4237);
xor U8483 (N_8483,N_4900,N_4151);
and U8484 (N_8484,N_4668,N_4979);
and U8485 (N_8485,N_6154,N_5409);
xor U8486 (N_8486,N_4236,N_3397);
or U8487 (N_8487,N_5254,N_4503);
and U8488 (N_8488,N_3536,N_5688);
nand U8489 (N_8489,N_3350,N_3400);
nand U8490 (N_8490,N_4569,N_5874);
and U8491 (N_8491,N_6098,N_4234);
xor U8492 (N_8492,N_3741,N_5195);
nor U8493 (N_8493,N_3517,N_3705);
or U8494 (N_8494,N_3144,N_4476);
or U8495 (N_8495,N_5358,N_4434);
or U8496 (N_8496,N_5350,N_4239);
and U8497 (N_8497,N_3774,N_5760);
nand U8498 (N_8498,N_5492,N_3430);
or U8499 (N_8499,N_5529,N_6149);
and U8500 (N_8500,N_4061,N_4820);
nor U8501 (N_8501,N_3793,N_3135);
nand U8502 (N_8502,N_3958,N_5741);
and U8503 (N_8503,N_5270,N_4400);
or U8504 (N_8504,N_6179,N_6177);
nand U8505 (N_8505,N_4129,N_5823);
nor U8506 (N_8506,N_5292,N_5588);
nand U8507 (N_8507,N_3856,N_4675);
nor U8508 (N_8508,N_6000,N_5076);
nand U8509 (N_8509,N_5439,N_5052);
and U8510 (N_8510,N_4815,N_4504);
nand U8511 (N_8511,N_5952,N_3396);
nor U8512 (N_8512,N_4946,N_3897);
or U8513 (N_8513,N_5625,N_4308);
and U8514 (N_8514,N_5245,N_5241);
nor U8515 (N_8515,N_4391,N_3364);
xor U8516 (N_8516,N_4613,N_3752);
nand U8517 (N_8517,N_5056,N_3259);
or U8518 (N_8518,N_4591,N_5275);
and U8519 (N_8519,N_4097,N_4991);
nand U8520 (N_8520,N_5472,N_5223);
nor U8521 (N_8521,N_3135,N_3735);
xor U8522 (N_8522,N_5824,N_3671);
or U8523 (N_8523,N_3818,N_3317);
xor U8524 (N_8524,N_5485,N_5705);
nor U8525 (N_8525,N_5756,N_5615);
and U8526 (N_8526,N_6051,N_4125);
or U8527 (N_8527,N_4679,N_5724);
or U8528 (N_8528,N_3795,N_3452);
nand U8529 (N_8529,N_4469,N_5445);
or U8530 (N_8530,N_5708,N_3708);
nor U8531 (N_8531,N_5386,N_3962);
and U8532 (N_8532,N_3698,N_3837);
and U8533 (N_8533,N_4415,N_5248);
xnor U8534 (N_8534,N_3606,N_5925);
or U8535 (N_8535,N_5719,N_5961);
nor U8536 (N_8536,N_5237,N_4789);
nor U8537 (N_8537,N_4879,N_6120);
nand U8538 (N_8538,N_5428,N_3317);
or U8539 (N_8539,N_3300,N_4907);
nand U8540 (N_8540,N_4171,N_6048);
or U8541 (N_8541,N_5245,N_3289);
nor U8542 (N_8542,N_3397,N_3452);
and U8543 (N_8543,N_4544,N_3971);
nand U8544 (N_8544,N_5456,N_4394);
nand U8545 (N_8545,N_3125,N_3385);
nand U8546 (N_8546,N_4321,N_4511);
nor U8547 (N_8547,N_3950,N_5870);
or U8548 (N_8548,N_4956,N_3266);
and U8549 (N_8549,N_3745,N_5966);
xor U8550 (N_8550,N_3922,N_4700);
or U8551 (N_8551,N_4045,N_3464);
or U8552 (N_8552,N_4159,N_5271);
nand U8553 (N_8553,N_4210,N_5358);
xor U8554 (N_8554,N_4048,N_4456);
and U8555 (N_8555,N_6146,N_5308);
xor U8556 (N_8556,N_6092,N_3433);
nand U8557 (N_8557,N_4061,N_4879);
or U8558 (N_8558,N_4700,N_4725);
or U8559 (N_8559,N_5297,N_5810);
or U8560 (N_8560,N_5610,N_3462);
nor U8561 (N_8561,N_5355,N_5011);
nand U8562 (N_8562,N_5809,N_3308);
nor U8563 (N_8563,N_4944,N_4379);
nand U8564 (N_8564,N_3225,N_5445);
and U8565 (N_8565,N_4056,N_3545);
nor U8566 (N_8566,N_5085,N_4789);
and U8567 (N_8567,N_6009,N_3268);
and U8568 (N_8568,N_5213,N_5221);
nor U8569 (N_8569,N_4108,N_3341);
nor U8570 (N_8570,N_3381,N_3308);
nand U8571 (N_8571,N_3407,N_3954);
and U8572 (N_8572,N_3240,N_3178);
nor U8573 (N_8573,N_3516,N_6157);
and U8574 (N_8574,N_4561,N_5198);
and U8575 (N_8575,N_3557,N_4582);
xnor U8576 (N_8576,N_5199,N_5453);
nand U8577 (N_8577,N_3665,N_4966);
and U8578 (N_8578,N_3648,N_5376);
nand U8579 (N_8579,N_5012,N_5328);
or U8580 (N_8580,N_4111,N_4075);
and U8581 (N_8581,N_3763,N_4459);
nor U8582 (N_8582,N_5926,N_3702);
nor U8583 (N_8583,N_4355,N_4769);
or U8584 (N_8584,N_5636,N_5780);
nor U8585 (N_8585,N_4563,N_5883);
and U8586 (N_8586,N_5167,N_6167);
and U8587 (N_8587,N_3508,N_3582);
and U8588 (N_8588,N_4856,N_4297);
nor U8589 (N_8589,N_6229,N_3772);
nand U8590 (N_8590,N_4128,N_3907);
nand U8591 (N_8591,N_4534,N_5810);
nor U8592 (N_8592,N_4206,N_5621);
xnor U8593 (N_8593,N_3620,N_5360);
nor U8594 (N_8594,N_3577,N_3929);
nor U8595 (N_8595,N_5951,N_6223);
and U8596 (N_8596,N_4365,N_4752);
and U8597 (N_8597,N_4730,N_4962);
nand U8598 (N_8598,N_4586,N_4038);
xor U8599 (N_8599,N_3627,N_5163);
and U8600 (N_8600,N_4230,N_3140);
and U8601 (N_8601,N_3807,N_3433);
or U8602 (N_8602,N_3616,N_3166);
or U8603 (N_8603,N_3623,N_3312);
nand U8604 (N_8604,N_5628,N_3793);
or U8605 (N_8605,N_5692,N_5600);
and U8606 (N_8606,N_4367,N_5339);
and U8607 (N_8607,N_3678,N_3285);
nand U8608 (N_8608,N_4351,N_4089);
nand U8609 (N_8609,N_6096,N_5643);
nand U8610 (N_8610,N_4070,N_4590);
nor U8611 (N_8611,N_5744,N_5867);
nor U8612 (N_8612,N_4798,N_3493);
or U8613 (N_8613,N_4660,N_3135);
nand U8614 (N_8614,N_3493,N_4054);
or U8615 (N_8615,N_5558,N_4419);
nand U8616 (N_8616,N_5356,N_5927);
or U8617 (N_8617,N_4887,N_6149);
nand U8618 (N_8618,N_3253,N_4470);
and U8619 (N_8619,N_3851,N_4543);
nand U8620 (N_8620,N_3679,N_4595);
or U8621 (N_8621,N_3835,N_5258);
or U8622 (N_8622,N_3386,N_3741);
nand U8623 (N_8623,N_3811,N_4765);
or U8624 (N_8624,N_3716,N_3371);
nand U8625 (N_8625,N_6175,N_4108);
or U8626 (N_8626,N_4700,N_4397);
nand U8627 (N_8627,N_3268,N_5080);
and U8628 (N_8628,N_3675,N_5959);
xor U8629 (N_8629,N_5508,N_5838);
nand U8630 (N_8630,N_4912,N_3767);
nand U8631 (N_8631,N_3153,N_5350);
nor U8632 (N_8632,N_4193,N_5255);
and U8633 (N_8633,N_3645,N_3346);
nor U8634 (N_8634,N_5834,N_5752);
and U8635 (N_8635,N_4053,N_3726);
nand U8636 (N_8636,N_5582,N_5142);
nor U8637 (N_8637,N_4995,N_5308);
and U8638 (N_8638,N_3514,N_3974);
xnor U8639 (N_8639,N_4204,N_4018);
xnor U8640 (N_8640,N_4136,N_5143);
or U8641 (N_8641,N_6100,N_4105);
or U8642 (N_8642,N_4722,N_6057);
nand U8643 (N_8643,N_5849,N_5493);
and U8644 (N_8644,N_4337,N_5567);
or U8645 (N_8645,N_4056,N_3934);
nand U8646 (N_8646,N_5745,N_4256);
nand U8647 (N_8647,N_4972,N_3338);
or U8648 (N_8648,N_4688,N_5940);
nand U8649 (N_8649,N_3786,N_3546);
and U8650 (N_8650,N_4144,N_4576);
xor U8651 (N_8651,N_6047,N_3986);
nor U8652 (N_8652,N_6126,N_5461);
and U8653 (N_8653,N_5273,N_3301);
or U8654 (N_8654,N_4166,N_4555);
nor U8655 (N_8655,N_4340,N_5092);
nand U8656 (N_8656,N_3756,N_5492);
nor U8657 (N_8657,N_5911,N_6172);
nand U8658 (N_8658,N_6228,N_3174);
xor U8659 (N_8659,N_5421,N_5084);
or U8660 (N_8660,N_4859,N_5997);
nor U8661 (N_8661,N_3619,N_3381);
nor U8662 (N_8662,N_5771,N_3561);
nand U8663 (N_8663,N_5319,N_3952);
nand U8664 (N_8664,N_4812,N_4892);
xnor U8665 (N_8665,N_3770,N_4459);
xor U8666 (N_8666,N_3995,N_5312);
nand U8667 (N_8667,N_5951,N_3500);
nand U8668 (N_8668,N_6216,N_3212);
and U8669 (N_8669,N_4689,N_5257);
and U8670 (N_8670,N_4308,N_5348);
nand U8671 (N_8671,N_5162,N_4663);
or U8672 (N_8672,N_4129,N_3780);
or U8673 (N_8673,N_5752,N_5144);
or U8674 (N_8674,N_4489,N_6006);
and U8675 (N_8675,N_6242,N_5555);
or U8676 (N_8676,N_5125,N_5891);
nor U8677 (N_8677,N_3580,N_5050);
nor U8678 (N_8678,N_5469,N_5679);
nand U8679 (N_8679,N_4514,N_5263);
xnor U8680 (N_8680,N_5539,N_5862);
nor U8681 (N_8681,N_6176,N_5494);
or U8682 (N_8682,N_5526,N_5661);
or U8683 (N_8683,N_4986,N_5676);
xor U8684 (N_8684,N_5002,N_6104);
nand U8685 (N_8685,N_5566,N_5649);
and U8686 (N_8686,N_3684,N_5400);
and U8687 (N_8687,N_5035,N_4276);
and U8688 (N_8688,N_4694,N_5882);
or U8689 (N_8689,N_4627,N_4551);
and U8690 (N_8690,N_3178,N_3236);
nand U8691 (N_8691,N_4675,N_6105);
and U8692 (N_8692,N_3346,N_4124);
xnor U8693 (N_8693,N_4353,N_5592);
or U8694 (N_8694,N_5343,N_4481);
nand U8695 (N_8695,N_6199,N_4986);
nor U8696 (N_8696,N_6179,N_3605);
nand U8697 (N_8697,N_4119,N_5860);
or U8698 (N_8698,N_4130,N_5379);
nor U8699 (N_8699,N_3621,N_4344);
nand U8700 (N_8700,N_4079,N_6236);
nor U8701 (N_8701,N_4177,N_3153);
nand U8702 (N_8702,N_5686,N_3898);
xnor U8703 (N_8703,N_3946,N_3149);
nor U8704 (N_8704,N_4410,N_3361);
and U8705 (N_8705,N_3329,N_5366);
xor U8706 (N_8706,N_3840,N_6121);
nand U8707 (N_8707,N_3850,N_4568);
xor U8708 (N_8708,N_6031,N_5827);
and U8709 (N_8709,N_4504,N_4018);
and U8710 (N_8710,N_5108,N_5543);
nand U8711 (N_8711,N_3798,N_5191);
or U8712 (N_8712,N_3138,N_4287);
nand U8713 (N_8713,N_3465,N_4175);
and U8714 (N_8714,N_3981,N_5846);
and U8715 (N_8715,N_4467,N_6005);
xnor U8716 (N_8716,N_6234,N_4006);
and U8717 (N_8717,N_5239,N_4269);
xor U8718 (N_8718,N_3991,N_3394);
nor U8719 (N_8719,N_5565,N_5924);
and U8720 (N_8720,N_3327,N_6073);
and U8721 (N_8721,N_4310,N_4312);
nor U8722 (N_8722,N_3380,N_5130);
nand U8723 (N_8723,N_3607,N_5107);
nor U8724 (N_8724,N_5046,N_3357);
nor U8725 (N_8725,N_3720,N_5775);
or U8726 (N_8726,N_4911,N_6182);
nand U8727 (N_8727,N_4660,N_3169);
nor U8728 (N_8728,N_4412,N_3829);
and U8729 (N_8729,N_3597,N_4146);
nor U8730 (N_8730,N_4748,N_4743);
nor U8731 (N_8731,N_4477,N_5681);
or U8732 (N_8732,N_4919,N_3528);
nor U8733 (N_8733,N_4462,N_5748);
and U8734 (N_8734,N_4522,N_4817);
or U8735 (N_8735,N_5788,N_4769);
nand U8736 (N_8736,N_4003,N_3281);
and U8737 (N_8737,N_4279,N_4175);
or U8738 (N_8738,N_5242,N_6160);
xnor U8739 (N_8739,N_3708,N_6094);
or U8740 (N_8740,N_4517,N_4914);
nand U8741 (N_8741,N_4943,N_4397);
or U8742 (N_8742,N_5863,N_5588);
nand U8743 (N_8743,N_3866,N_3218);
or U8744 (N_8744,N_3950,N_5529);
nand U8745 (N_8745,N_3299,N_5023);
nand U8746 (N_8746,N_5936,N_3537);
and U8747 (N_8747,N_4263,N_3132);
nand U8748 (N_8748,N_3695,N_5814);
nor U8749 (N_8749,N_5016,N_5052);
or U8750 (N_8750,N_4644,N_3961);
or U8751 (N_8751,N_4057,N_4859);
nand U8752 (N_8752,N_4500,N_3731);
or U8753 (N_8753,N_5668,N_4804);
nor U8754 (N_8754,N_3236,N_5351);
and U8755 (N_8755,N_4520,N_3318);
nand U8756 (N_8756,N_3229,N_3545);
or U8757 (N_8757,N_5950,N_3267);
nor U8758 (N_8758,N_5208,N_5003);
nor U8759 (N_8759,N_3247,N_5206);
and U8760 (N_8760,N_5161,N_3937);
and U8761 (N_8761,N_5141,N_4418);
and U8762 (N_8762,N_5628,N_5181);
nand U8763 (N_8763,N_5739,N_6230);
or U8764 (N_8764,N_4371,N_5868);
nand U8765 (N_8765,N_6038,N_4995);
xor U8766 (N_8766,N_4003,N_5860);
or U8767 (N_8767,N_5435,N_5498);
and U8768 (N_8768,N_5275,N_4811);
nor U8769 (N_8769,N_6119,N_6207);
nor U8770 (N_8770,N_4794,N_5792);
nor U8771 (N_8771,N_4565,N_5637);
and U8772 (N_8772,N_5617,N_5783);
nor U8773 (N_8773,N_3881,N_5197);
nand U8774 (N_8774,N_4266,N_3971);
xor U8775 (N_8775,N_5000,N_3954);
nor U8776 (N_8776,N_4521,N_4680);
xor U8777 (N_8777,N_5306,N_5513);
and U8778 (N_8778,N_4689,N_5919);
or U8779 (N_8779,N_5589,N_5305);
nand U8780 (N_8780,N_6029,N_5421);
or U8781 (N_8781,N_3517,N_3605);
nand U8782 (N_8782,N_3410,N_3357);
nor U8783 (N_8783,N_6211,N_4944);
nor U8784 (N_8784,N_5657,N_5102);
nand U8785 (N_8785,N_4378,N_4786);
nor U8786 (N_8786,N_3614,N_3284);
or U8787 (N_8787,N_3882,N_4693);
nor U8788 (N_8788,N_4009,N_5163);
nand U8789 (N_8789,N_5188,N_4739);
and U8790 (N_8790,N_6233,N_5718);
and U8791 (N_8791,N_4728,N_3348);
nor U8792 (N_8792,N_4507,N_5722);
or U8793 (N_8793,N_4602,N_3830);
xnor U8794 (N_8794,N_5789,N_4138);
or U8795 (N_8795,N_3471,N_5078);
nor U8796 (N_8796,N_5139,N_4098);
nand U8797 (N_8797,N_4436,N_5624);
nand U8798 (N_8798,N_4745,N_3747);
nand U8799 (N_8799,N_3189,N_5694);
nor U8800 (N_8800,N_5463,N_4292);
nand U8801 (N_8801,N_3912,N_4606);
nor U8802 (N_8802,N_6239,N_3730);
and U8803 (N_8803,N_3160,N_5489);
xor U8804 (N_8804,N_3901,N_4372);
or U8805 (N_8805,N_3338,N_3867);
nand U8806 (N_8806,N_3734,N_5472);
nand U8807 (N_8807,N_3267,N_5029);
xnor U8808 (N_8808,N_5717,N_3860);
and U8809 (N_8809,N_5257,N_5364);
nor U8810 (N_8810,N_5069,N_3980);
or U8811 (N_8811,N_4223,N_6020);
nor U8812 (N_8812,N_5004,N_5722);
nand U8813 (N_8813,N_5665,N_4349);
and U8814 (N_8814,N_4004,N_4710);
or U8815 (N_8815,N_5905,N_4840);
or U8816 (N_8816,N_6112,N_3139);
and U8817 (N_8817,N_3181,N_4517);
xor U8818 (N_8818,N_4752,N_5845);
or U8819 (N_8819,N_5790,N_4528);
xnor U8820 (N_8820,N_3739,N_4967);
or U8821 (N_8821,N_3579,N_3912);
and U8822 (N_8822,N_5192,N_5827);
nand U8823 (N_8823,N_5325,N_5080);
xor U8824 (N_8824,N_4882,N_5565);
nor U8825 (N_8825,N_4547,N_3308);
or U8826 (N_8826,N_4134,N_5978);
nor U8827 (N_8827,N_5480,N_5676);
xor U8828 (N_8828,N_5444,N_4669);
xor U8829 (N_8829,N_5846,N_3610);
or U8830 (N_8830,N_5033,N_4723);
or U8831 (N_8831,N_5559,N_5872);
nor U8832 (N_8832,N_5517,N_4082);
nand U8833 (N_8833,N_3487,N_4621);
or U8834 (N_8834,N_4021,N_3508);
and U8835 (N_8835,N_4076,N_3231);
nor U8836 (N_8836,N_4393,N_4068);
nand U8837 (N_8837,N_3244,N_3590);
nor U8838 (N_8838,N_4384,N_3779);
and U8839 (N_8839,N_3149,N_5444);
nand U8840 (N_8840,N_3890,N_5251);
nand U8841 (N_8841,N_5083,N_3566);
or U8842 (N_8842,N_3138,N_5324);
xnor U8843 (N_8843,N_5469,N_4989);
and U8844 (N_8844,N_3796,N_3276);
and U8845 (N_8845,N_5210,N_5172);
or U8846 (N_8846,N_4079,N_5691);
nand U8847 (N_8847,N_6075,N_3870);
and U8848 (N_8848,N_4320,N_5391);
nor U8849 (N_8849,N_5922,N_4614);
or U8850 (N_8850,N_6146,N_4423);
nand U8851 (N_8851,N_5227,N_3509);
nand U8852 (N_8852,N_3185,N_6218);
and U8853 (N_8853,N_4189,N_5257);
or U8854 (N_8854,N_3645,N_4803);
nand U8855 (N_8855,N_3287,N_3879);
nor U8856 (N_8856,N_3635,N_5890);
and U8857 (N_8857,N_4843,N_5905);
or U8858 (N_8858,N_4905,N_3971);
or U8859 (N_8859,N_5254,N_3613);
nor U8860 (N_8860,N_5668,N_5591);
or U8861 (N_8861,N_4020,N_3855);
xor U8862 (N_8862,N_5202,N_4320);
and U8863 (N_8863,N_5608,N_6082);
nor U8864 (N_8864,N_5026,N_6046);
xnor U8865 (N_8865,N_3845,N_4825);
nand U8866 (N_8866,N_6046,N_3863);
nand U8867 (N_8867,N_3411,N_5624);
or U8868 (N_8868,N_4735,N_4966);
nor U8869 (N_8869,N_3263,N_4663);
nor U8870 (N_8870,N_3894,N_4350);
or U8871 (N_8871,N_5095,N_6055);
and U8872 (N_8872,N_4836,N_3300);
nor U8873 (N_8873,N_3793,N_5934);
and U8874 (N_8874,N_4092,N_4417);
and U8875 (N_8875,N_4000,N_5609);
and U8876 (N_8876,N_6165,N_5502);
or U8877 (N_8877,N_4150,N_5937);
xor U8878 (N_8878,N_5758,N_4513);
nand U8879 (N_8879,N_6215,N_4476);
or U8880 (N_8880,N_3667,N_3455);
nand U8881 (N_8881,N_5939,N_5313);
nand U8882 (N_8882,N_5389,N_4275);
xor U8883 (N_8883,N_4284,N_5808);
xor U8884 (N_8884,N_5471,N_5866);
or U8885 (N_8885,N_5702,N_5445);
and U8886 (N_8886,N_4788,N_3497);
or U8887 (N_8887,N_4478,N_5630);
nor U8888 (N_8888,N_5638,N_3870);
and U8889 (N_8889,N_4557,N_4646);
nor U8890 (N_8890,N_4465,N_5124);
and U8891 (N_8891,N_5708,N_5162);
or U8892 (N_8892,N_6100,N_4329);
nor U8893 (N_8893,N_6215,N_3464);
nor U8894 (N_8894,N_4988,N_4285);
and U8895 (N_8895,N_5132,N_6183);
nor U8896 (N_8896,N_4192,N_3790);
and U8897 (N_8897,N_5745,N_6024);
nor U8898 (N_8898,N_4352,N_4868);
and U8899 (N_8899,N_5022,N_5219);
or U8900 (N_8900,N_5762,N_4017);
nor U8901 (N_8901,N_5741,N_4989);
and U8902 (N_8902,N_5235,N_4950);
or U8903 (N_8903,N_3177,N_3536);
nor U8904 (N_8904,N_4975,N_3132);
nor U8905 (N_8905,N_5254,N_3441);
xor U8906 (N_8906,N_5473,N_5014);
and U8907 (N_8907,N_4181,N_4236);
xor U8908 (N_8908,N_4821,N_5888);
or U8909 (N_8909,N_4684,N_5568);
or U8910 (N_8910,N_5346,N_4618);
nor U8911 (N_8911,N_3337,N_5853);
and U8912 (N_8912,N_3322,N_4475);
nand U8913 (N_8913,N_5321,N_4821);
nor U8914 (N_8914,N_4128,N_5182);
xor U8915 (N_8915,N_6085,N_3465);
xor U8916 (N_8916,N_4964,N_4240);
nand U8917 (N_8917,N_4177,N_5677);
or U8918 (N_8918,N_3985,N_4238);
or U8919 (N_8919,N_6146,N_4328);
or U8920 (N_8920,N_4584,N_5440);
nor U8921 (N_8921,N_5131,N_3182);
xnor U8922 (N_8922,N_5469,N_5922);
nand U8923 (N_8923,N_4365,N_3378);
and U8924 (N_8924,N_5482,N_5860);
or U8925 (N_8925,N_3794,N_5819);
and U8926 (N_8926,N_5227,N_3210);
nand U8927 (N_8927,N_5111,N_3623);
nor U8928 (N_8928,N_4036,N_4018);
nor U8929 (N_8929,N_4008,N_5612);
nor U8930 (N_8930,N_4789,N_5336);
nand U8931 (N_8931,N_5329,N_5561);
nor U8932 (N_8932,N_4125,N_3860);
nor U8933 (N_8933,N_4231,N_4548);
or U8934 (N_8934,N_5593,N_5690);
and U8935 (N_8935,N_5114,N_6161);
and U8936 (N_8936,N_5044,N_4357);
nand U8937 (N_8937,N_4563,N_4111);
nand U8938 (N_8938,N_5992,N_4207);
nand U8939 (N_8939,N_3309,N_4515);
xnor U8940 (N_8940,N_3763,N_4571);
or U8941 (N_8941,N_4128,N_4915);
or U8942 (N_8942,N_3793,N_3796);
xor U8943 (N_8943,N_3813,N_5491);
nor U8944 (N_8944,N_3337,N_3697);
or U8945 (N_8945,N_4433,N_5546);
nor U8946 (N_8946,N_5232,N_6216);
or U8947 (N_8947,N_3526,N_3968);
nor U8948 (N_8948,N_3880,N_5312);
nor U8949 (N_8949,N_4916,N_4230);
and U8950 (N_8950,N_3339,N_5242);
or U8951 (N_8951,N_6232,N_5124);
and U8952 (N_8952,N_5356,N_6030);
and U8953 (N_8953,N_5485,N_6029);
or U8954 (N_8954,N_5303,N_3632);
nor U8955 (N_8955,N_6078,N_5629);
or U8956 (N_8956,N_4916,N_5740);
nor U8957 (N_8957,N_5263,N_6150);
nor U8958 (N_8958,N_6080,N_6066);
nor U8959 (N_8959,N_5970,N_4684);
nor U8960 (N_8960,N_5726,N_6176);
or U8961 (N_8961,N_3253,N_4790);
or U8962 (N_8962,N_4713,N_5920);
nor U8963 (N_8963,N_3527,N_4712);
nand U8964 (N_8964,N_4690,N_3584);
or U8965 (N_8965,N_3512,N_5030);
and U8966 (N_8966,N_4710,N_6097);
and U8967 (N_8967,N_4331,N_4732);
nand U8968 (N_8968,N_5262,N_4813);
nand U8969 (N_8969,N_6222,N_6089);
and U8970 (N_8970,N_3692,N_3969);
and U8971 (N_8971,N_4295,N_5077);
nor U8972 (N_8972,N_6016,N_4656);
or U8973 (N_8973,N_3813,N_5665);
or U8974 (N_8974,N_5011,N_4294);
and U8975 (N_8975,N_5309,N_3912);
nand U8976 (N_8976,N_5004,N_3568);
or U8977 (N_8977,N_3909,N_5526);
nor U8978 (N_8978,N_4215,N_4538);
and U8979 (N_8979,N_3198,N_5069);
nand U8980 (N_8980,N_4216,N_5200);
and U8981 (N_8981,N_4134,N_4794);
nand U8982 (N_8982,N_3626,N_4591);
or U8983 (N_8983,N_3358,N_3283);
nor U8984 (N_8984,N_4335,N_5669);
and U8985 (N_8985,N_6246,N_3944);
nand U8986 (N_8986,N_3278,N_4711);
xnor U8987 (N_8987,N_5683,N_3474);
nor U8988 (N_8988,N_4663,N_4102);
or U8989 (N_8989,N_5094,N_6025);
nand U8990 (N_8990,N_3808,N_3745);
nand U8991 (N_8991,N_4060,N_3484);
xor U8992 (N_8992,N_6237,N_4554);
nor U8993 (N_8993,N_3735,N_5954);
nand U8994 (N_8994,N_4260,N_3757);
xnor U8995 (N_8995,N_5896,N_4302);
and U8996 (N_8996,N_4157,N_3591);
or U8997 (N_8997,N_6076,N_4516);
or U8998 (N_8998,N_3667,N_3579);
or U8999 (N_8999,N_4520,N_3937);
xnor U9000 (N_9000,N_4611,N_5775);
or U9001 (N_9001,N_4412,N_4835);
and U9002 (N_9002,N_6143,N_5414);
nor U9003 (N_9003,N_4330,N_6023);
nor U9004 (N_9004,N_4205,N_5604);
xor U9005 (N_9005,N_3405,N_5910);
nor U9006 (N_9006,N_4025,N_5582);
and U9007 (N_9007,N_5259,N_4294);
and U9008 (N_9008,N_4610,N_5787);
or U9009 (N_9009,N_4491,N_3348);
nor U9010 (N_9010,N_5770,N_5032);
or U9011 (N_9011,N_4099,N_3334);
nand U9012 (N_9012,N_5956,N_3125);
and U9013 (N_9013,N_3532,N_5932);
or U9014 (N_9014,N_5355,N_6050);
xor U9015 (N_9015,N_5822,N_4724);
nor U9016 (N_9016,N_4564,N_4889);
xor U9017 (N_9017,N_5225,N_4448);
nor U9018 (N_9018,N_6235,N_5490);
nand U9019 (N_9019,N_5702,N_3372);
and U9020 (N_9020,N_5966,N_5439);
or U9021 (N_9021,N_3963,N_5526);
nand U9022 (N_9022,N_4461,N_4651);
nor U9023 (N_9023,N_4340,N_5261);
or U9024 (N_9024,N_4762,N_4068);
nor U9025 (N_9025,N_5106,N_4547);
or U9026 (N_9026,N_5795,N_4226);
nor U9027 (N_9027,N_5561,N_5262);
nand U9028 (N_9028,N_4943,N_5383);
and U9029 (N_9029,N_4539,N_5748);
or U9030 (N_9030,N_5113,N_4425);
or U9031 (N_9031,N_3969,N_3653);
nand U9032 (N_9032,N_6222,N_5824);
nor U9033 (N_9033,N_5517,N_3182);
and U9034 (N_9034,N_5900,N_4698);
nor U9035 (N_9035,N_6046,N_3997);
or U9036 (N_9036,N_5928,N_4175);
nor U9037 (N_9037,N_3602,N_4068);
nor U9038 (N_9038,N_3705,N_3891);
and U9039 (N_9039,N_4770,N_4809);
or U9040 (N_9040,N_4514,N_4092);
nand U9041 (N_9041,N_4124,N_5598);
or U9042 (N_9042,N_3982,N_6151);
nand U9043 (N_9043,N_5662,N_4015);
or U9044 (N_9044,N_3656,N_3650);
and U9045 (N_9045,N_6039,N_3295);
or U9046 (N_9046,N_4117,N_4889);
and U9047 (N_9047,N_6234,N_5587);
nor U9048 (N_9048,N_4068,N_5964);
nand U9049 (N_9049,N_5592,N_6008);
xor U9050 (N_9050,N_5756,N_5648);
xnor U9051 (N_9051,N_4990,N_6141);
xnor U9052 (N_9052,N_4705,N_5498);
nor U9053 (N_9053,N_4804,N_5788);
or U9054 (N_9054,N_5825,N_5580);
xor U9055 (N_9055,N_5398,N_4731);
or U9056 (N_9056,N_3891,N_4455);
nor U9057 (N_9057,N_5210,N_5359);
nand U9058 (N_9058,N_3550,N_5573);
or U9059 (N_9059,N_3381,N_5157);
nand U9060 (N_9060,N_3928,N_3489);
xor U9061 (N_9061,N_4613,N_3245);
nor U9062 (N_9062,N_3814,N_4887);
nand U9063 (N_9063,N_4773,N_6219);
and U9064 (N_9064,N_3391,N_4604);
xnor U9065 (N_9065,N_5893,N_3688);
nor U9066 (N_9066,N_3809,N_4989);
nand U9067 (N_9067,N_3872,N_3522);
or U9068 (N_9068,N_4114,N_5601);
and U9069 (N_9069,N_4787,N_3308);
nand U9070 (N_9070,N_6214,N_5141);
xnor U9071 (N_9071,N_3677,N_4690);
xor U9072 (N_9072,N_5756,N_5211);
xnor U9073 (N_9073,N_4551,N_5990);
or U9074 (N_9074,N_4743,N_5653);
nor U9075 (N_9075,N_5230,N_5217);
or U9076 (N_9076,N_4526,N_4661);
nor U9077 (N_9077,N_3325,N_5188);
and U9078 (N_9078,N_4545,N_5575);
or U9079 (N_9079,N_5204,N_3634);
nand U9080 (N_9080,N_3955,N_3264);
nor U9081 (N_9081,N_4226,N_4568);
and U9082 (N_9082,N_3247,N_6156);
nand U9083 (N_9083,N_6125,N_5023);
or U9084 (N_9084,N_3802,N_5240);
or U9085 (N_9085,N_5766,N_3326);
or U9086 (N_9086,N_4667,N_5530);
or U9087 (N_9087,N_4687,N_5759);
or U9088 (N_9088,N_4005,N_5132);
and U9089 (N_9089,N_4913,N_4783);
nor U9090 (N_9090,N_4289,N_5924);
and U9091 (N_9091,N_5488,N_5244);
and U9092 (N_9092,N_6171,N_3454);
and U9093 (N_9093,N_3229,N_4535);
or U9094 (N_9094,N_5789,N_5363);
nand U9095 (N_9095,N_4284,N_6030);
nor U9096 (N_9096,N_3614,N_4327);
or U9097 (N_9097,N_4668,N_5012);
nand U9098 (N_9098,N_4085,N_5948);
nand U9099 (N_9099,N_5465,N_3246);
nand U9100 (N_9100,N_3544,N_6161);
and U9101 (N_9101,N_5211,N_5942);
nor U9102 (N_9102,N_4872,N_4303);
or U9103 (N_9103,N_5787,N_6096);
and U9104 (N_9104,N_5384,N_3672);
or U9105 (N_9105,N_5133,N_4261);
nor U9106 (N_9106,N_3806,N_3781);
nor U9107 (N_9107,N_3225,N_4355);
and U9108 (N_9108,N_3881,N_5294);
and U9109 (N_9109,N_3358,N_5963);
and U9110 (N_9110,N_4281,N_5393);
and U9111 (N_9111,N_5451,N_5684);
or U9112 (N_9112,N_4450,N_5346);
nand U9113 (N_9113,N_5220,N_5690);
nor U9114 (N_9114,N_3671,N_4054);
nor U9115 (N_9115,N_3159,N_3386);
nand U9116 (N_9116,N_3991,N_5520);
and U9117 (N_9117,N_4555,N_4880);
and U9118 (N_9118,N_3867,N_5876);
and U9119 (N_9119,N_5640,N_4938);
nand U9120 (N_9120,N_5845,N_4177);
nand U9121 (N_9121,N_5883,N_5763);
and U9122 (N_9122,N_3989,N_3712);
nand U9123 (N_9123,N_5368,N_3700);
xor U9124 (N_9124,N_3908,N_4486);
and U9125 (N_9125,N_3407,N_3435);
nor U9126 (N_9126,N_5009,N_5741);
nor U9127 (N_9127,N_3293,N_6013);
nand U9128 (N_9128,N_5117,N_5914);
nor U9129 (N_9129,N_4033,N_4973);
or U9130 (N_9130,N_5537,N_3604);
or U9131 (N_9131,N_6048,N_4130);
nand U9132 (N_9132,N_3927,N_5485);
or U9133 (N_9133,N_4082,N_4546);
nor U9134 (N_9134,N_4326,N_3771);
nand U9135 (N_9135,N_4943,N_4336);
nand U9136 (N_9136,N_4199,N_5275);
nor U9137 (N_9137,N_5848,N_5256);
or U9138 (N_9138,N_6042,N_5760);
or U9139 (N_9139,N_4229,N_4366);
nand U9140 (N_9140,N_5855,N_3424);
nor U9141 (N_9141,N_5214,N_4805);
xnor U9142 (N_9142,N_4382,N_6231);
nand U9143 (N_9143,N_4176,N_5747);
or U9144 (N_9144,N_5282,N_4969);
and U9145 (N_9145,N_3531,N_4300);
and U9146 (N_9146,N_4155,N_4509);
nor U9147 (N_9147,N_4128,N_6244);
nor U9148 (N_9148,N_4588,N_6237);
nor U9149 (N_9149,N_6071,N_4508);
or U9150 (N_9150,N_4404,N_4442);
xor U9151 (N_9151,N_4265,N_5015);
xnor U9152 (N_9152,N_5224,N_4840);
nand U9153 (N_9153,N_6014,N_3681);
and U9154 (N_9154,N_5032,N_4345);
and U9155 (N_9155,N_5440,N_5194);
nor U9156 (N_9156,N_3544,N_6243);
nor U9157 (N_9157,N_4143,N_6028);
and U9158 (N_9158,N_4922,N_5392);
or U9159 (N_9159,N_5626,N_3187);
xor U9160 (N_9160,N_6068,N_4207);
or U9161 (N_9161,N_4950,N_5703);
nor U9162 (N_9162,N_3894,N_3686);
xor U9163 (N_9163,N_4608,N_4039);
nand U9164 (N_9164,N_5195,N_5608);
and U9165 (N_9165,N_5520,N_3834);
xor U9166 (N_9166,N_5178,N_6247);
nor U9167 (N_9167,N_3615,N_5910);
nand U9168 (N_9168,N_6027,N_5427);
nand U9169 (N_9169,N_5703,N_6159);
nand U9170 (N_9170,N_4841,N_3177);
and U9171 (N_9171,N_5935,N_4394);
xor U9172 (N_9172,N_4546,N_3367);
or U9173 (N_9173,N_3196,N_5935);
nand U9174 (N_9174,N_4827,N_4941);
xor U9175 (N_9175,N_6057,N_4552);
and U9176 (N_9176,N_5110,N_4085);
or U9177 (N_9177,N_4265,N_3201);
nor U9178 (N_9178,N_4196,N_4491);
nand U9179 (N_9179,N_3510,N_3847);
nor U9180 (N_9180,N_5298,N_3771);
nor U9181 (N_9181,N_5313,N_6022);
nand U9182 (N_9182,N_4451,N_6091);
xor U9183 (N_9183,N_4515,N_4749);
and U9184 (N_9184,N_5746,N_5510);
and U9185 (N_9185,N_4840,N_4411);
and U9186 (N_9186,N_5526,N_4970);
nor U9187 (N_9187,N_4160,N_5918);
and U9188 (N_9188,N_4181,N_4679);
nor U9189 (N_9189,N_3386,N_4892);
nand U9190 (N_9190,N_5957,N_5283);
nor U9191 (N_9191,N_4875,N_3983);
nor U9192 (N_9192,N_5663,N_5288);
nor U9193 (N_9193,N_4507,N_5266);
or U9194 (N_9194,N_5305,N_3857);
nor U9195 (N_9195,N_4526,N_6201);
and U9196 (N_9196,N_4528,N_6204);
nor U9197 (N_9197,N_5154,N_6247);
nand U9198 (N_9198,N_4855,N_3364);
and U9199 (N_9199,N_4330,N_3527);
nor U9200 (N_9200,N_4361,N_3571);
or U9201 (N_9201,N_4760,N_4716);
and U9202 (N_9202,N_5599,N_5169);
nor U9203 (N_9203,N_3742,N_4490);
nand U9204 (N_9204,N_3199,N_3243);
nand U9205 (N_9205,N_5397,N_4669);
nand U9206 (N_9206,N_3348,N_6142);
or U9207 (N_9207,N_3171,N_3276);
xor U9208 (N_9208,N_5614,N_4814);
nor U9209 (N_9209,N_5770,N_5782);
nor U9210 (N_9210,N_3850,N_4828);
or U9211 (N_9211,N_5704,N_3791);
nand U9212 (N_9212,N_3340,N_3683);
and U9213 (N_9213,N_3855,N_4429);
nor U9214 (N_9214,N_5871,N_3768);
nor U9215 (N_9215,N_3830,N_3308);
or U9216 (N_9216,N_6153,N_5487);
nor U9217 (N_9217,N_5418,N_4853);
and U9218 (N_9218,N_4842,N_4317);
nor U9219 (N_9219,N_5589,N_3605);
and U9220 (N_9220,N_5673,N_4889);
or U9221 (N_9221,N_3144,N_3683);
xnor U9222 (N_9222,N_5068,N_3648);
and U9223 (N_9223,N_5753,N_4089);
nor U9224 (N_9224,N_5071,N_3169);
nor U9225 (N_9225,N_5547,N_4894);
nor U9226 (N_9226,N_3393,N_3863);
nor U9227 (N_9227,N_4519,N_4643);
or U9228 (N_9228,N_3930,N_4028);
nand U9229 (N_9229,N_3326,N_4188);
nor U9230 (N_9230,N_5346,N_6139);
xor U9231 (N_9231,N_4292,N_4389);
and U9232 (N_9232,N_6160,N_5264);
nand U9233 (N_9233,N_4054,N_4791);
xnor U9234 (N_9234,N_5463,N_3582);
or U9235 (N_9235,N_3329,N_5829);
nor U9236 (N_9236,N_4084,N_5478);
nor U9237 (N_9237,N_6232,N_5336);
and U9238 (N_9238,N_4206,N_3601);
or U9239 (N_9239,N_3402,N_6061);
nand U9240 (N_9240,N_5842,N_4519);
or U9241 (N_9241,N_4717,N_4682);
or U9242 (N_9242,N_4047,N_3790);
and U9243 (N_9243,N_5578,N_4949);
and U9244 (N_9244,N_5973,N_5321);
and U9245 (N_9245,N_5149,N_3766);
xor U9246 (N_9246,N_6074,N_3243);
nor U9247 (N_9247,N_5409,N_5837);
nor U9248 (N_9248,N_4602,N_3794);
xor U9249 (N_9249,N_5153,N_3674);
nor U9250 (N_9250,N_3267,N_5008);
nand U9251 (N_9251,N_5342,N_5181);
nand U9252 (N_9252,N_3555,N_3178);
and U9253 (N_9253,N_3369,N_4324);
or U9254 (N_9254,N_5518,N_4566);
nand U9255 (N_9255,N_4181,N_5999);
or U9256 (N_9256,N_5620,N_5717);
and U9257 (N_9257,N_5778,N_4169);
nand U9258 (N_9258,N_5525,N_5916);
nand U9259 (N_9259,N_3279,N_4753);
or U9260 (N_9260,N_3744,N_4648);
nand U9261 (N_9261,N_5901,N_5621);
and U9262 (N_9262,N_5470,N_5544);
or U9263 (N_9263,N_3796,N_3963);
or U9264 (N_9264,N_5395,N_5329);
or U9265 (N_9265,N_5630,N_3768);
nand U9266 (N_9266,N_4303,N_3597);
nor U9267 (N_9267,N_4735,N_4362);
or U9268 (N_9268,N_4219,N_6062);
or U9269 (N_9269,N_3642,N_5996);
nor U9270 (N_9270,N_5706,N_4443);
or U9271 (N_9271,N_6086,N_4831);
or U9272 (N_9272,N_5078,N_5409);
and U9273 (N_9273,N_4185,N_4209);
or U9274 (N_9274,N_3490,N_3987);
and U9275 (N_9275,N_5872,N_6136);
nand U9276 (N_9276,N_3495,N_3917);
nand U9277 (N_9277,N_5270,N_5514);
nand U9278 (N_9278,N_5790,N_3382);
or U9279 (N_9279,N_4105,N_5014);
and U9280 (N_9280,N_4901,N_4135);
nand U9281 (N_9281,N_4049,N_4625);
nand U9282 (N_9282,N_5150,N_6146);
nor U9283 (N_9283,N_4329,N_5515);
nor U9284 (N_9284,N_6237,N_3931);
and U9285 (N_9285,N_3282,N_5834);
nand U9286 (N_9286,N_6115,N_5757);
or U9287 (N_9287,N_6076,N_5653);
nand U9288 (N_9288,N_4126,N_5000);
nor U9289 (N_9289,N_5732,N_4728);
nor U9290 (N_9290,N_5199,N_5501);
nand U9291 (N_9291,N_3353,N_4936);
and U9292 (N_9292,N_5023,N_3166);
nor U9293 (N_9293,N_5829,N_3723);
or U9294 (N_9294,N_3792,N_5435);
nand U9295 (N_9295,N_4697,N_4534);
and U9296 (N_9296,N_3345,N_4668);
and U9297 (N_9297,N_5000,N_5495);
and U9298 (N_9298,N_4135,N_4503);
and U9299 (N_9299,N_3837,N_4759);
nand U9300 (N_9300,N_6053,N_3692);
or U9301 (N_9301,N_5660,N_3396);
or U9302 (N_9302,N_5092,N_3791);
nand U9303 (N_9303,N_5255,N_5581);
or U9304 (N_9304,N_3355,N_3163);
or U9305 (N_9305,N_4041,N_6241);
or U9306 (N_9306,N_4475,N_4620);
xnor U9307 (N_9307,N_3994,N_4140);
and U9308 (N_9308,N_4952,N_5160);
or U9309 (N_9309,N_3889,N_4488);
nor U9310 (N_9310,N_3677,N_5357);
nor U9311 (N_9311,N_3346,N_4216);
or U9312 (N_9312,N_5604,N_5009);
and U9313 (N_9313,N_4024,N_5090);
and U9314 (N_9314,N_5319,N_4019);
xor U9315 (N_9315,N_5384,N_4197);
or U9316 (N_9316,N_4868,N_4313);
and U9317 (N_9317,N_5854,N_5269);
or U9318 (N_9318,N_3505,N_5781);
nor U9319 (N_9319,N_3482,N_4848);
nand U9320 (N_9320,N_3769,N_5199);
nor U9321 (N_9321,N_3150,N_4788);
nand U9322 (N_9322,N_5786,N_5832);
and U9323 (N_9323,N_4577,N_4413);
xnor U9324 (N_9324,N_5235,N_3824);
and U9325 (N_9325,N_3300,N_3568);
or U9326 (N_9326,N_4991,N_4005);
nand U9327 (N_9327,N_4663,N_4233);
nand U9328 (N_9328,N_4841,N_3767);
nor U9329 (N_9329,N_3927,N_5582);
and U9330 (N_9330,N_5397,N_5701);
and U9331 (N_9331,N_4951,N_6081);
nor U9332 (N_9332,N_3798,N_4768);
and U9333 (N_9333,N_5497,N_3481);
nand U9334 (N_9334,N_5870,N_3720);
nor U9335 (N_9335,N_5521,N_3275);
nor U9336 (N_9336,N_4411,N_5040);
and U9337 (N_9337,N_3680,N_4554);
and U9338 (N_9338,N_4500,N_4032);
or U9339 (N_9339,N_4695,N_4783);
nor U9340 (N_9340,N_4670,N_4495);
or U9341 (N_9341,N_5657,N_5688);
nand U9342 (N_9342,N_6232,N_4854);
and U9343 (N_9343,N_4353,N_4654);
or U9344 (N_9344,N_5503,N_6004);
nand U9345 (N_9345,N_3213,N_3674);
nand U9346 (N_9346,N_3912,N_5302);
nand U9347 (N_9347,N_4541,N_3529);
nand U9348 (N_9348,N_3476,N_4323);
xor U9349 (N_9349,N_5135,N_4483);
xnor U9350 (N_9350,N_6046,N_5901);
nor U9351 (N_9351,N_3407,N_4658);
or U9352 (N_9352,N_5613,N_5020);
or U9353 (N_9353,N_6093,N_4154);
or U9354 (N_9354,N_3875,N_6070);
nand U9355 (N_9355,N_5508,N_5895);
or U9356 (N_9356,N_5411,N_3936);
or U9357 (N_9357,N_3135,N_5906);
or U9358 (N_9358,N_5824,N_4617);
or U9359 (N_9359,N_5753,N_5294);
and U9360 (N_9360,N_4563,N_6223);
or U9361 (N_9361,N_5773,N_5104);
xor U9362 (N_9362,N_5693,N_6042);
or U9363 (N_9363,N_5181,N_4142);
nor U9364 (N_9364,N_4599,N_4601);
or U9365 (N_9365,N_5097,N_5295);
and U9366 (N_9366,N_3960,N_3985);
and U9367 (N_9367,N_5847,N_5292);
or U9368 (N_9368,N_4461,N_3856);
or U9369 (N_9369,N_4111,N_3524);
or U9370 (N_9370,N_5329,N_3930);
nand U9371 (N_9371,N_3903,N_5604);
or U9372 (N_9372,N_3652,N_4344);
nor U9373 (N_9373,N_3933,N_3815);
or U9374 (N_9374,N_5715,N_6170);
nor U9375 (N_9375,N_9026,N_7585);
and U9376 (N_9376,N_7872,N_7444);
nor U9377 (N_9377,N_6341,N_7683);
and U9378 (N_9378,N_6680,N_8476);
xor U9379 (N_9379,N_8037,N_8447);
or U9380 (N_9380,N_7209,N_6374);
xor U9381 (N_9381,N_7600,N_8766);
nand U9382 (N_9382,N_6478,N_7761);
nor U9383 (N_9383,N_6423,N_7555);
or U9384 (N_9384,N_7676,N_6530);
nor U9385 (N_9385,N_6657,N_8985);
nor U9386 (N_9386,N_6630,N_8478);
or U9387 (N_9387,N_8844,N_8206);
or U9388 (N_9388,N_6332,N_8966);
and U9389 (N_9389,N_7064,N_9247);
and U9390 (N_9390,N_7671,N_7785);
and U9391 (N_9391,N_8615,N_7499);
nor U9392 (N_9392,N_7774,N_7941);
and U9393 (N_9393,N_9016,N_9007);
nor U9394 (N_9394,N_6595,N_8714);
and U9395 (N_9395,N_8073,N_8957);
nor U9396 (N_9396,N_7652,N_7181);
or U9397 (N_9397,N_6601,N_8998);
and U9398 (N_9398,N_7684,N_8276);
nand U9399 (N_9399,N_6632,N_7927);
nor U9400 (N_9400,N_7929,N_9237);
and U9401 (N_9401,N_8630,N_8872);
nand U9402 (N_9402,N_6288,N_7971);
and U9403 (N_9403,N_6519,N_8520);
nand U9404 (N_9404,N_6927,N_7514);
nand U9405 (N_9405,N_7184,N_6890);
or U9406 (N_9406,N_7047,N_6324);
or U9407 (N_9407,N_7067,N_8560);
and U9408 (N_9408,N_6469,N_9298);
and U9409 (N_9409,N_6274,N_6713);
or U9410 (N_9410,N_7120,N_7098);
nor U9411 (N_9411,N_8819,N_6804);
nor U9412 (N_9412,N_6788,N_7391);
or U9413 (N_9413,N_6344,N_8363);
and U9414 (N_9414,N_6455,N_7352);
nor U9415 (N_9415,N_7297,N_6742);
xnor U9416 (N_9416,N_9202,N_7000);
nor U9417 (N_9417,N_8951,N_7214);
nor U9418 (N_9418,N_7368,N_7885);
and U9419 (N_9419,N_8466,N_8954);
and U9420 (N_9420,N_8369,N_8774);
and U9421 (N_9421,N_8927,N_8924);
nand U9422 (N_9422,N_6677,N_8298);
or U9423 (N_9423,N_7336,N_8022);
nor U9424 (N_9424,N_8582,N_8930);
nor U9425 (N_9425,N_9302,N_9249);
nand U9426 (N_9426,N_8070,N_7486);
and U9427 (N_9427,N_8482,N_6527);
or U9428 (N_9428,N_8418,N_8009);
or U9429 (N_9429,N_6418,N_9077);
nand U9430 (N_9430,N_7325,N_6328);
xnor U9431 (N_9431,N_7105,N_6377);
nand U9432 (N_9432,N_7407,N_7225);
or U9433 (N_9433,N_6326,N_6602);
or U9434 (N_9434,N_8550,N_8187);
nor U9435 (N_9435,N_8758,N_6803);
nand U9436 (N_9436,N_6404,N_6522);
nor U9437 (N_9437,N_7726,N_8024);
nand U9438 (N_9438,N_7501,N_6408);
nand U9439 (N_9439,N_7769,N_9331);
xnor U9440 (N_9440,N_7453,N_8485);
or U9441 (N_9441,N_7837,N_6446);
nor U9442 (N_9442,N_8039,N_7574);
nor U9443 (N_9443,N_9082,N_8891);
nor U9444 (N_9444,N_8744,N_7232);
and U9445 (N_9445,N_6728,N_6375);
or U9446 (N_9446,N_8342,N_8554);
xnor U9447 (N_9447,N_7691,N_7218);
nand U9448 (N_9448,N_8423,N_8131);
or U9449 (N_9449,N_9114,N_8120);
nor U9450 (N_9450,N_8464,N_8311);
nand U9451 (N_9451,N_8531,N_7379);
or U9452 (N_9452,N_7507,N_7782);
nor U9453 (N_9453,N_9312,N_8134);
or U9454 (N_9454,N_6960,N_8156);
nand U9455 (N_9455,N_6600,N_8949);
nand U9456 (N_9456,N_7815,N_7750);
nor U9457 (N_9457,N_7418,N_7515);
and U9458 (N_9458,N_6979,N_7932);
nor U9459 (N_9459,N_6827,N_7995);
and U9460 (N_9460,N_9314,N_6605);
or U9461 (N_9461,N_7475,N_7796);
or U9462 (N_9462,N_7638,N_8196);
and U9463 (N_9463,N_8641,N_8701);
xnor U9464 (N_9464,N_7554,N_7570);
or U9465 (N_9465,N_8257,N_9316);
and U9466 (N_9466,N_6476,N_7029);
or U9467 (N_9467,N_6621,N_8452);
nand U9468 (N_9468,N_9104,N_6946);
nand U9469 (N_9469,N_6255,N_7398);
nor U9470 (N_9470,N_9038,N_6631);
or U9471 (N_9471,N_7051,N_6580);
and U9472 (N_9472,N_8788,N_8188);
nand U9473 (N_9473,N_6428,N_7033);
or U9474 (N_9474,N_7044,N_7481);
xnor U9475 (N_9475,N_9290,N_8099);
nor U9476 (N_9476,N_7655,N_6831);
nor U9477 (N_9477,N_8326,N_8569);
nor U9478 (N_9478,N_9269,N_6973);
nor U9479 (N_9479,N_8525,N_8361);
or U9480 (N_9480,N_8907,N_6870);
nor U9481 (N_9481,N_6805,N_7696);
and U9482 (N_9482,N_8979,N_6734);
xnor U9483 (N_9483,N_8807,N_8167);
or U9484 (N_9484,N_7918,N_8421);
and U9485 (N_9485,N_6450,N_6568);
and U9486 (N_9486,N_7198,N_8217);
and U9487 (N_9487,N_7913,N_7246);
and U9488 (N_9488,N_8224,N_9060);
or U9489 (N_9489,N_8793,N_9241);
nor U9490 (N_9490,N_7353,N_7955);
nand U9491 (N_9491,N_8465,N_6997);
nor U9492 (N_9492,N_9116,N_6437);
and U9493 (N_9493,N_8555,N_9035);
and U9494 (N_9494,N_7204,N_8723);
xnor U9495 (N_9495,N_7459,N_6394);
nand U9496 (N_9496,N_9232,N_8289);
and U9497 (N_9497,N_6257,N_8247);
xor U9498 (N_9498,N_7176,N_8876);
xor U9499 (N_9499,N_8946,N_7463);
nand U9500 (N_9500,N_7830,N_6860);
and U9501 (N_9501,N_6270,N_6572);
nor U9502 (N_9502,N_8270,N_7337);
and U9503 (N_9503,N_7512,N_7364);
xnor U9504 (N_9504,N_9118,N_7448);
nand U9505 (N_9505,N_6492,N_7817);
nor U9506 (N_9506,N_6771,N_7328);
xnor U9507 (N_9507,N_9043,N_6373);
nand U9508 (N_9508,N_7721,N_7624);
or U9509 (N_9509,N_8350,N_7842);
xnor U9510 (N_9510,N_9178,N_8823);
nand U9511 (N_9511,N_6473,N_8040);
or U9512 (N_9512,N_9276,N_7393);
or U9513 (N_9513,N_8138,N_8858);
nand U9514 (N_9514,N_7496,N_7944);
and U9515 (N_9515,N_6393,N_7552);
and U9516 (N_9516,N_7189,N_7345);
or U9517 (N_9517,N_6589,N_7523);
nor U9518 (N_9518,N_8454,N_9059);
and U9519 (N_9519,N_9158,N_6956);
nand U9520 (N_9520,N_6647,N_6686);
and U9521 (N_9521,N_6252,N_8800);
nand U9522 (N_9522,N_7382,N_7112);
or U9523 (N_9523,N_7828,N_8061);
nor U9524 (N_9524,N_7313,N_7521);
nor U9525 (N_9525,N_8585,N_6367);
or U9526 (N_9526,N_8082,N_9175);
nor U9527 (N_9527,N_9045,N_7043);
or U9528 (N_9528,N_7806,N_6296);
nor U9529 (N_9529,N_7793,N_7991);
and U9530 (N_9530,N_7505,N_9075);
nor U9531 (N_9531,N_9288,N_8574);
nor U9532 (N_9532,N_8570,N_9162);
nor U9533 (N_9533,N_8010,N_7708);
or U9534 (N_9534,N_7236,N_8147);
nand U9535 (N_9535,N_8351,N_6312);
or U9536 (N_9536,N_6787,N_6834);
and U9537 (N_9537,N_8797,N_6325);
or U9538 (N_9538,N_6526,N_7791);
nand U9539 (N_9539,N_8389,N_7951);
xor U9540 (N_9540,N_9221,N_6940);
nor U9541 (N_9541,N_6421,N_6710);
nand U9542 (N_9542,N_7504,N_8140);
nand U9543 (N_9543,N_8095,N_6379);
and U9544 (N_9544,N_6697,N_7703);
or U9545 (N_9545,N_9133,N_8502);
nand U9546 (N_9546,N_8353,N_9359);
xor U9547 (N_9547,N_6900,N_7395);
nor U9548 (N_9548,N_7053,N_9238);
or U9549 (N_9549,N_8209,N_6843);
and U9550 (N_9550,N_6555,N_8873);
or U9551 (N_9551,N_7472,N_6550);
and U9552 (N_9552,N_6648,N_7613);
xor U9553 (N_9553,N_6342,N_8854);
nand U9554 (N_9554,N_7199,N_7320);
or U9555 (N_9555,N_7277,N_7532);
nand U9556 (N_9556,N_6869,N_6735);
and U9557 (N_9557,N_7034,N_8014);
xor U9558 (N_9558,N_7113,N_6738);
or U9559 (N_9559,N_7611,N_8056);
xnor U9560 (N_9560,N_8069,N_8590);
or U9561 (N_9561,N_8137,N_8975);
xor U9562 (N_9562,N_8529,N_9216);
nor U9563 (N_9563,N_6297,N_8005);
and U9564 (N_9564,N_6516,N_8471);
or U9565 (N_9565,N_9368,N_9130);
nand U9566 (N_9566,N_8086,N_6863);
nand U9567 (N_9567,N_7329,N_7257);
nor U9568 (N_9568,N_7487,N_8584);
and U9569 (N_9569,N_6984,N_8781);
xnor U9570 (N_9570,N_7771,N_8197);
nand U9571 (N_9571,N_8097,N_6503);
and U9572 (N_9572,N_6856,N_7138);
nand U9573 (N_9573,N_6359,N_9356);
or U9574 (N_9574,N_6266,N_8186);
nand U9575 (N_9575,N_8833,N_7429);
or U9576 (N_9576,N_6792,N_8982);
nand U9577 (N_9577,N_8060,N_9189);
and U9578 (N_9578,N_8850,N_7768);
nand U9579 (N_9579,N_6416,N_6949);
or U9580 (N_9580,N_9063,N_7833);
and U9581 (N_9581,N_7119,N_9141);
or U9582 (N_9582,N_7590,N_6350);
and U9583 (N_9583,N_7388,N_7491);
and U9584 (N_9584,N_8827,N_8412);
and U9585 (N_9585,N_7931,N_7753);
nand U9586 (N_9586,N_8176,N_6761);
nor U9587 (N_9587,N_9284,N_8019);
or U9588 (N_9588,N_9145,N_6878);
nand U9589 (N_9589,N_6942,N_7021);
xor U9590 (N_9590,N_9039,N_8612);
nor U9591 (N_9591,N_8623,N_9264);
or U9592 (N_9592,N_7569,N_7001);
and U9593 (N_9593,N_8669,N_8756);
nor U9594 (N_9594,N_7871,N_8253);
or U9595 (N_9595,N_9062,N_7455);
nand U9596 (N_9596,N_9258,N_7200);
and U9597 (N_9597,N_7245,N_7254);
nand U9598 (N_9598,N_8749,N_6798);
and U9599 (N_9599,N_6935,N_6389);
xnor U9600 (N_9600,N_7832,N_7719);
or U9601 (N_9601,N_7168,N_7593);
nor U9602 (N_9602,N_6793,N_9323);
nor U9603 (N_9603,N_7934,N_7981);
nor U9604 (N_9604,N_7211,N_8620);
nand U9605 (N_9605,N_7973,N_9046);
and U9606 (N_9606,N_8309,N_8692);
and U9607 (N_9607,N_7502,N_7383);
nand U9608 (N_9608,N_9228,N_6833);
nor U9609 (N_9609,N_8201,N_6392);
nor U9610 (N_9610,N_6382,N_7525);
nand U9611 (N_9611,N_8481,N_8182);
and U9612 (N_9612,N_7042,N_8210);
or U9613 (N_9613,N_7739,N_8296);
nor U9614 (N_9614,N_6371,N_6988);
xor U9615 (N_9615,N_8559,N_9244);
nand U9616 (N_9616,N_8154,N_6966);
nor U9617 (N_9617,N_6420,N_7962);
nor U9618 (N_9618,N_8020,N_8849);
xor U9619 (N_9619,N_8422,N_6744);
and U9620 (N_9620,N_8614,N_6453);
and U9621 (N_9621,N_7848,N_9171);
and U9622 (N_9622,N_7510,N_7142);
nor U9623 (N_9623,N_6897,N_8769);
nand U9624 (N_9624,N_8483,N_6770);
and U9625 (N_9625,N_6877,N_8436);
nand U9626 (N_9626,N_8871,N_8677);
or U9627 (N_9627,N_7953,N_6299);
and U9628 (N_9628,N_8987,N_6447);
nand U9629 (N_9629,N_7415,N_6560);
or U9630 (N_9630,N_9306,N_7612);
nor U9631 (N_9631,N_6357,N_6513);
nand U9632 (N_9632,N_8696,N_8811);
xor U9633 (N_9633,N_7035,N_6578);
nor U9634 (N_9634,N_9353,N_8242);
nand U9635 (N_9635,N_8319,N_6585);
or U9636 (N_9636,N_8294,N_7937);
or U9637 (N_9637,N_7623,N_6906);
nor U9638 (N_9638,N_7930,N_9139);
nand U9639 (N_9639,N_6561,N_6544);
nand U9640 (N_9640,N_8320,N_9289);
nor U9641 (N_9641,N_8052,N_7697);
nor U9642 (N_9642,N_8035,N_7037);
nor U9643 (N_9643,N_7449,N_7926);
and U9644 (N_9644,N_6820,N_6429);
xor U9645 (N_9645,N_8406,N_8348);
or U9646 (N_9646,N_7898,N_8128);
and U9647 (N_9647,N_9255,N_8135);
or U9648 (N_9648,N_8625,N_7031);
or U9649 (N_9649,N_8912,N_8607);
and U9650 (N_9650,N_6845,N_6322);
nor U9651 (N_9651,N_6262,N_8272);
or U9652 (N_9652,N_7835,N_6385);
and U9653 (N_9653,N_6642,N_8246);
or U9654 (N_9654,N_6810,N_8906);
or U9655 (N_9655,N_7661,N_7859);
nor U9656 (N_9656,N_8980,N_8512);
nand U9657 (N_9657,N_7924,N_7050);
or U9658 (N_9658,N_8653,N_6756);
or U9659 (N_9659,N_7964,N_8660);
or U9660 (N_9660,N_7602,N_9033);
and U9661 (N_9661,N_7087,N_7907);
nand U9662 (N_9662,N_7447,N_7026);
nand U9663 (N_9663,N_8417,N_8757);
nand U9664 (N_9664,N_8259,N_8707);
nand U9665 (N_9665,N_6610,N_7904);
nand U9666 (N_9666,N_7466,N_8395);
nor U9667 (N_9667,N_6767,N_6992);
and U9668 (N_9668,N_9156,N_6289);
and U9669 (N_9669,N_8738,N_8915);
or U9670 (N_9670,N_7702,N_8725);
nand U9671 (N_9671,N_6826,N_8494);
or U9672 (N_9672,N_7392,N_8543);
nand U9673 (N_9673,N_7109,N_7262);
or U9674 (N_9674,N_6491,N_8174);
and U9675 (N_9675,N_7967,N_8087);
or U9676 (N_9676,N_9049,N_7528);
nand U9677 (N_9677,N_8942,N_7096);
nor U9678 (N_9678,N_7462,N_6316);
nand U9679 (N_9679,N_7680,N_6864);
nor U9680 (N_9680,N_7949,N_7206);
or U9681 (N_9681,N_7735,N_8396);
nor U9682 (N_9682,N_6961,N_8305);
xor U9683 (N_9683,N_6926,N_7966);
xor U9684 (N_9684,N_6868,N_8286);
nor U9685 (N_9685,N_6551,N_7668);
nor U9686 (N_9686,N_7695,N_6780);
nand U9687 (N_9687,N_7356,N_7860);
nand U9688 (N_9688,N_8455,N_7477);
nor U9689 (N_9689,N_6822,N_9372);
or U9690 (N_9690,N_7667,N_6776);
nor U9691 (N_9691,N_6620,N_8558);
nor U9692 (N_9692,N_8534,N_6565);
or U9693 (N_9693,N_7989,N_8332);
nor U9694 (N_9694,N_7909,N_7071);
nor U9695 (N_9695,N_6690,N_8180);
nand U9696 (N_9696,N_8984,N_7538);
nor U9697 (N_9697,N_8895,N_8699);
xnor U9698 (N_9698,N_8935,N_6458);
and U9699 (N_9699,N_8226,N_6765);
nand U9700 (N_9700,N_6950,N_6579);
nor U9701 (N_9701,N_9294,N_6957);
xor U9702 (N_9702,N_6584,N_8404);
and U9703 (N_9703,N_7224,N_8648);
nor U9704 (N_9704,N_8388,N_8074);
nand U9705 (N_9705,N_8463,N_8967);
nor U9706 (N_9706,N_6909,N_6464);
nand U9707 (N_9707,N_8025,N_9093);
and U9708 (N_9708,N_7943,N_7694);
and U9709 (N_9709,N_7542,N_6635);
nand U9710 (N_9710,N_7984,N_8011);
nand U9711 (N_9711,N_6823,N_6460);
and U9712 (N_9712,N_9013,N_8255);
and U9713 (N_9713,N_6470,N_7597);
nor U9714 (N_9714,N_7314,N_7014);
or U9715 (N_9715,N_7917,N_9087);
xnor U9716 (N_9716,N_6576,N_6508);
nor U9717 (N_9717,N_7799,N_9137);
and U9718 (N_9718,N_9124,N_6801);
nor U9719 (N_9719,N_9256,N_7445);
xor U9720 (N_9720,N_8116,N_8882);
and U9721 (N_9721,N_7377,N_6661);
or U9722 (N_9722,N_9120,N_8815);
nor U9723 (N_9723,N_8674,N_6836);
and U9724 (N_9724,N_8355,N_8732);
nor U9725 (N_9725,N_8928,N_9134);
nor U9726 (N_9726,N_7020,N_6953);
nand U9727 (N_9727,N_9340,N_7500);
nor U9728 (N_9728,N_7707,N_6989);
nand U9729 (N_9729,N_7258,N_6529);
nor U9730 (N_9730,N_6637,N_7527);
or U9731 (N_9731,N_7072,N_9301);
nor U9732 (N_9732,N_7411,N_8085);
and U9733 (N_9733,N_6459,N_8825);
nand U9734 (N_9734,N_7836,N_6912);
nor U9735 (N_9735,N_7776,N_8077);
nand U9736 (N_9736,N_6852,N_7728);
and U9737 (N_9737,N_9210,N_8031);
nand U9738 (N_9738,N_8521,N_8983);
or U9739 (N_9739,N_7471,N_7963);
xor U9740 (N_9740,N_9006,N_7742);
nand U9741 (N_9741,N_7010,N_7342);
or U9742 (N_9742,N_6285,N_6644);
nand U9743 (N_9743,N_6790,N_8248);
or U9744 (N_9744,N_7012,N_8597);
nor U9745 (N_9745,N_8889,N_7226);
and U9746 (N_9746,N_7889,N_7055);
and U9747 (N_9747,N_8857,N_7790);
xor U9748 (N_9748,N_6407,N_8991);
nor U9749 (N_9749,N_7108,N_7549);
nand U9750 (N_9750,N_7249,N_7323);
or U9751 (N_9751,N_7959,N_9079);
or U9752 (N_9752,N_8084,N_6733);
or U9753 (N_9753,N_7945,N_8199);
nor U9754 (N_9754,N_9111,N_9277);
or U9755 (N_9755,N_6786,N_6272);
or U9756 (N_9756,N_9251,N_7789);
or U9757 (N_9757,N_8159,N_7028);
and U9758 (N_9758,N_7062,N_7992);
or U9759 (N_9759,N_7573,N_7078);
or U9760 (N_9760,N_7027,N_7221);
xor U9761 (N_9761,N_8727,N_8146);
and U9762 (N_9762,N_6977,N_9036);
nor U9763 (N_9763,N_7275,N_6656);
nand U9764 (N_9764,N_7781,N_8149);
nand U9765 (N_9765,N_9180,N_8232);
nor U9766 (N_9766,N_6483,N_6553);
or U9767 (N_9767,N_6796,N_7185);
nand U9768 (N_9768,N_6874,N_8901);
xnor U9769 (N_9769,N_7102,N_6865);
or U9770 (N_9770,N_7066,N_7141);
and U9771 (N_9771,N_9211,N_8608);
nor U9772 (N_9772,N_9149,N_6467);
nor U9773 (N_9773,N_6302,N_8491);
nand U9774 (N_9774,N_9084,N_8808);
xnor U9775 (N_9775,N_7478,N_8121);
nand U9776 (N_9776,N_6717,N_9272);
and U9777 (N_9777,N_8595,N_9119);
nor U9778 (N_9778,N_8778,N_8038);
or U9779 (N_9779,N_7400,N_6613);
or U9780 (N_9780,N_6318,N_6295);
and U9781 (N_9781,N_7894,N_8460);
and U9782 (N_9782,N_9278,N_8575);
and U9783 (N_9783,N_8430,N_7681);
and U9784 (N_9784,N_8853,N_7912);
nand U9785 (N_9785,N_7792,N_7384);
and U9786 (N_9786,N_7343,N_9354);
and U9787 (N_9787,N_9097,N_9196);
nand U9788 (N_9788,N_8992,N_8724);
or U9789 (N_9789,N_6722,N_7845);
or U9790 (N_9790,N_7324,N_8684);
or U9791 (N_9791,N_8576,N_7698);
and U9792 (N_9792,N_6655,N_8770);
nand U9793 (N_9793,N_7059,N_7701);
or U9794 (N_9794,N_6965,N_6751);
xor U9795 (N_9795,N_6435,N_8688);
and U9796 (N_9796,N_7686,N_7317);
nor U9797 (N_9797,N_7004,N_9235);
and U9798 (N_9798,N_8451,N_7560);
xor U9799 (N_9799,N_7150,N_8497);
and U9800 (N_9800,N_6387,N_7238);
and U9801 (N_9801,N_6754,N_8855);
nor U9802 (N_9802,N_7744,N_8431);
nand U9803 (N_9803,N_7809,N_9088);
nand U9804 (N_9804,N_7239,N_9339);
xor U9805 (N_9805,N_8216,N_9273);
or U9806 (N_9806,N_8231,N_8904);
xor U9807 (N_9807,N_7158,N_6673);
and U9808 (N_9808,N_8008,N_9150);
xor U9809 (N_9809,N_6923,N_8842);
nor U9810 (N_9810,N_8646,N_8484);
nand U9811 (N_9811,N_9303,N_8760);
nand U9812 (N_9812,N_8530,N_8391);
or U9813 (N_9813,N_8596,N_7298);
and U9814 (N_9814,N_7456,N_7381);
or U9815 (N_9815,N_7094,N_7092);
or U9816 (N_9816,N_7643,N_8939);
nand U9817 (N_9817,N_9096,N_8593);
and U9818 (N_9818,N_8274,N_7764);
nor U9819 (N_9819,N_8258,N_8301);
nor U9820 (N_9820,N_8337,N_8978);
and U9821 (N_9821,N_6507,N_6496);
or U9822 (N_9822,N_6685,N_6514);
and U9823 (N_9823,N_6766,N_7641);
nand U9824 (N_9824,N_8459,N_6866);
and U9825 (N_9825,N_7647,N_6384);
and U9826 (N_9826,N_6711,N_7006);
nand U9827 (N_9827,N_9000,N_7152);
nor U9828 (N_9828,N_7834,N_7111);
and U9829 (N_9829,N_6719,N_7431);
and U9830 (N_9830,N_6709,N_7048);
nor U9831 (N_9831,N_7737,N_8129);
or U9832 (N_9832,N_8923,N_8169);
and U9833 (N_9833,N_6769,N_8618);
or U9834 (N_9834,N_8133,N_8409);
or U9835 (N_9835,N_7760,N_8683);
or U9836 (N_9836,N_7887,N_8233);
and U9837 (N_9837,N_7127,N_8376);
and U9838 (N_9838,N_7242,N_7575);
or U9839 (N_9839,N_8079,N_7983);
or U9840 (N_9840,N_7339,N_7503);
and U9841 (N_9841,N_7670,N_7191);
and U9842 (N_9842,N_6405,N_7172);
nand U9843 (N_9843,N_7371,N_7334);
nor U9844 (N_9844,N_6993,N_9098);
and U9845 (N_9845,N_7274,N_7634);
and U9846 (N_9846,N_8791,N_9300);
and U9847 (N_9847,N_6417,N_6368);
or U9848 (N_9848,N_8645,N_6920);
xnor U9849 (N_9849,N_8603,N_9168);
or U9850 (N_9850,N_7545,N_6276);
nor U9851 (N_9851,N_7970,N_8103);
and U9852 (N_9852,N_7188,N_8043);
nand U9853 (N_9853,N_8658,N_6778);
nand U9854 (N_9854,N_7644,N_7080);
nor U9855 (N_9855,N_7787,N_7414);
or U9856 (N_9856,N_6914,N_8848);
and U9857 (N_9857,N_8711,N_9034);
xor U9858 (N_9858,N_6345,N_8606);
nand U9859 (N_9859,N_8687,N_8547);
nor U9860 (N_9860,N_7628,N_8972);
and U9861 (N_9861,N_7149,N_7897);
nand U9862 (N_9862,N_6971,N_7843);
nor U9863 (N_9863,N_6556,N_8161);
nor U9864 (N_9864,N_8151,N_8054);
xor U9865 (N_9865,N_8415,N_8937);
or U9866 (N_9866,N_7940,N_7621);
nand U9867 (N_9867,N_8950,N_8874);
nand U9868 (N_9868,N_7405,N_6430);
nand U9869 (N_9869,N_7762,N_9342);
or U9870 (N_9870,N_8492,N_6517);
or U9871 (N_9871,N_9056,N_9282);
or U9872 (N_9872,N_8704,N_8986);
or U9873 (N_9873,N_8314,N_6269);
nand U9874 (N_9874,N_9052,N_7687);
or U9875 (N_9875,N_7874,N_9190);
and U9876 (N_9876,N_8589,N_7089);
nor U9877 (N_9877,N_7725,N_8746);
or U9878 (N_9878,N_7359,N_7117);
xor U9879 (N_9879,N_8662,N_7315);
or U9880 (N_9880,N_8327,N_6740);
nor U9881 (N_9881,N_7219,N_6277);
xnor U9882 (N_9882,N_7133,N_6693);
nor U9883 (N_9883,N_8798,N_7594);
nor U9884 (N_9884,N_8425,N_9335);
nor U9885 (N_9885,N_7164,N_6259);
or U9886 (N_9886,N_6571,N_7002);
nor U9887 (N_9887,N_6542,N_8312);
nand U9888 (N_9888,N_7378,N_7699);
and U9889 (N_9889,N_7658,N_7947);
nand U9890 (N_9890,N_7968,N_8624);
nand U9891 (N_9891,N_7822,N_8899);
and U9892 (N_9892,N_8905,N_8165);
nand U9893 (N_9893,N_6347,N_7305);
and U9894 (N_9894,N_7582,N_6583);
nor U9895 (N_9895,N_9172,N_8440);
nor U9896 (N_9896,N_7583,N_8375);
xor U9897 (N_9897,N_8619,N_7264);
xor U9898 (N_9898,N_7531,N_9267);
and U9899 (N_9899,N_7802,N_6898);
and U9900 (N_9900,N_7289,N_7539);
and U9901 (N_9901,N_7197,N_7895);
nand U9902 (N_9902,N_7630,N_8453);
and U9903 (N_9903,N_7069,N_6286);
nor U9904 (N_9904,N_6358,N_9142);
and U9905 (N_9905,N_7233,N_6484);
or U9906 (N_9906,N_7143,N_8256);
xnor U9907 (N_9907,N_6715,N_6528);
or U9908 (N_9908,N_8617,N_8324);
nor U9909 (N_9909,N_6759,N_9047);
and U9910 (N_9910,N_7442,N_8837);
and U9911 (N_9911,N_8410,N_7367);
and U9912 (N_9912,N_6905,N_6694);
nand U9913 (N_9913,N_8959,N_7706);
nor U9914 (N_9914,N_9191,N_7852);
nor U9915 (N_9915,N_8599,N_7302);
or U9916 (N_9916,N_9243,N_9009);
nor U9917 (N_9917,N_8820,N_9352);
and U9918 (N_9918,N_7438,N_6982);
nor U9919 (N_9919,N_8293,N_6448);
or U9920 (N_9920,N_6391,N_6936);
and U9921 (N_9921,N_7609,N_8628);
and U9922 (N_9922,N_6764,N_6265);
xor U9923 (N_9923,N_7101,N_6627);
nand U9924 (N_9924,N_8831,N_7550);
and U9925 (N_9925,N_9100,N_7451);
or U9926 (N_9926,N_8212,N_7088);
and U9927 (N_9927,N_8068,N_7135);
and U9928 (N_9928,N_7022,N_8977);
or U9929 (N_9929,N_7625,N_8777);
or U9930 (N_9930,N_8513,N_7757);
and U9931 (N_9931,N_6369,N_8731);
and U9932 (N_9932,N_8109,N_6895);
and U9933 (N_9933,N_6378,N_9037);
or U9934 (N_9934,N_6918,N_8368);
xor U9935 (N_9935,N_9230,N_9207);
or U9936 (N_9936,N_9018,N_8932);
xor U9937 (N_9937,N_8012,N_6310);
and U9938 (N_9938,N_6360,N_6575);
nand U9939 (N_9939,N_8262,N_6271);
and U9940 (N_9940,N_8001,N_8053);
nand U9941 (N_9941,N_8456,N_9024);
nand U9942 (N_9942,N_8065,N_6293);
or U9943 (N_9943,N_9102,N_8101);
and U9944 (N_9944,N_8916,N_9280);
or U9945 (N_9945,N_7403,N_8782);
or U9946 (N_9946,N_7678,N_8123);
xor U9947 (N_9947,N_7160,N_9184);
xor U9948 (N_9948,N_7373,N_9113);
nor U9949 (N_9949,N_7363,N_9151);
nor U9950 (N_9950,N_6838,N_6329);
nand U9951 (N_9951,N_8693,N_7266);
or U9952 (N_9952,N_7730,N_7090);
and U9953 (N_9953,N_7736,N_8860);
nand U9954 (N_9954,N_6789,N_6974);
nor U9955 (N_9955,N_9311,N_6915);
nand U9956 (N_9956,N_7480,N_9362);
nor U9957 (N_9957,N_8875,N_9260);
nand U9958 (N_9958,N_7358,N_7212);
nand U9959 (N_9959,N_8878,N_9003);
and U9960 (N_9960,N_6612,N_7402);
xor U9961 (N_9961,N_6493,N_7454);
xnor U9962 (N_9962,N_8280,N_6313);
nor U9963 (N_9963,N_8969,N_6899);
and U9964 (N_9964,N_9348,N_7712);
nor U9965 (N_9965,N_8870,N_7495);
nand U9966 (N_9966,N_8107,N_6684);
and U9967 (N_9967,N_7629,N_6250);
nor U9968 (N_9968,N_7821,N_8962);
nor U9969 (N_9969,N_7155,N_8885);
or U9970 (N_9970,N_8726,N_7354);
nand U9971 (N_9971,N_8571,N_6741);
nor U9972 (N_9972,N_8290,N_9222);
and U9973 (N_9973,N_7045,N_9292);
and U9974 (N_9974,N_8679,N_6816);
and U9975 (N_9975,N_7952,N_7350);
xor U9976 (N_9976,N_8843,N_9345);
or U9977 (N_9977,N_6263,N_9032);
or U9978 (N_9978,N_6650,N_8173);
and U9979 (N_9979,N_8903,N_8432);
nand U9980 (N_9980,N_8659,N_7344);
and U9981 (N_9981,N_7261,N_8790);
nand U9982 (N_9982,N_6861,N_7954);
and U9983 (N_9983,N_8690,N_6910);
nand U9984 (N_9984,N_6959,N_8245);
or U9985 (N_9985,N_8856,N_7013);
or U9986 (N_9986,N_8185,N_6361);
nor U9987 (N_9987,N_9004,N_7385);
or U9988 (N_9988,N_9055,N_7919);
nand U9989 (N_9989,N_6623,N_6844);
nand U9990 (N_9990,N_6840,N_8062);
nand U9991 (N_9991,N_8445,N_6907);
or U9992 (N_9992,N_6254,N_8473);
and U9993 (N_9993,N_6533,N_7482);
or U9994 (N_9994,N_6559,N_6309);
nor U9995 (N_9995,N_9246,N_8918);
and U9996 (N_9996,N_7559,N_8393);
nor U9997 (N_9997,N_6903,N_6434);
or U9998 (N_9998,N_9201,N_6543);
nand U9999 (N_9999,N_7977,N_6337);
or U10000 (N_10000,N_7085,N_7811);
xor U10001 (N_10001,N_6762,N_9239);
nand U10002 (N_10002,N_7015,N_8055);
nor U10003 (N_10003,N_7417,N_6440);
xnor U10004 (N_10004,N_7177,N_6847);
or U10005 (N_10005,N_6943,N_6958);
nor U10006 (N_10006,N_7146,N_8064);
and U10007 (N_10007,N_9330,N_6925);
nor U10008 (N_10008,N_6463,N_6921);
nand U10009 (N_10009,N_6883,N_7580);
nand U10010 (N_10010,N_7194,N_8536);
and U10011 (N_10011,N_7902,N_6566);
nor U10012 (N_10012,N_7556,N_7942);
and U10013 (N_10013,N_7717,N_7030);
or U10014 (N_10014,N_6747,N_8081);
nand U10015 (N_10015,N_7599,N_8613);
and U10016 (N_10016,N_8522,N_7908);
nand U10017 (N_10017,N_6636,N_7125);
nor U10018 (N_10018,N_8036,N_7999);
or U10019 (N_10019,N_7269,N_6807);
nand U10020 (N_10020,N_7326,N_7443);
nand U10021 (N_10021,N_9002,N_6461);
nand U10022 (N_10022,N_8424,N_8349);
nand U10023 (N_10023,N_6567,N_8102);
nor U10024 (N_10024,N_7399,N_6646);
or U10025 (N_10025,N_7025,N_8921);
nand U10026 (N_10026,N_8322,N_6330);
and U10027 (N_10027,N_7118,N_8219);
xor U10028 (N_10028,N_9136,N_8139);
xor U10029 (N_10029,N_7838,N_7606);
or U10030 (N_10030,N_9364,N_8556);
and U10031 (N_10031,N_7637,N_8435);
and U10032 (N_10032,N_8268,N_8303);
or U10033 (N_10033,N_8426,N_7714);
nor U10034 (N_10034,N_9268,N_7673);
nand U10035 (N_10035,N_8868,N_8428);
and U10036 (N_10036,N_8526,N_9085);
nor U10037 (N_10037,N_7483,N_8018);
or U10038 (N_10038,N_6590,N_7095);
xor U10039 (N_10039,N_6626,N_7631);
and U10040 (N_10040,N_9324,N_8446);
nand U10041 (N_10041,N_9068,N_7288);
and U10042 (N_10042,N_8675,N_7891);
nor U10043 (N_10043,N_8006,N_8826);
or U10044 (N_10044,N_8275,N_7518);
and U10045 (N_10045,N_8551,N_6449);
nand U10046 (N_10046,N_6990,N_6406);
nor U10047 (N_10047,N_8661,N_8578);
and U10048 (N_10048,N_8490,N_7097);
and U10049 (N_10049,N_9253,N_6451);
nor U10050 (N_10050,N_6340,N_7474);
or U10051 (N_10051,N_8030,N_8474);
or U10052 (N_10052,N_9309,N_9065);
xor U10053 (N_10053,N_9297,N_8971);
and U10054 (N_10054,N_8514,N_7517);
or U10055 (N_10055,N_8881,N_8000);
and U10056 (N_10056,N_9233,N_7642);
nand U10057 (N_10057,N_9275,N_6707);
nor U10058 (N_10058,N_8325,N_7460);
xor U10059 (N_10059,N_9027,N_8150);
and U10060 (N_10060,N_6401,N_9174);
or U10061 (N_10061,N_7139,N_6839);
nand U10062 (N_10062,N_6706,N_8656);
nand U10063 (N_10063,N_8118,N_7153);
nand U10064 (N_10064,N_7147,N_8754);
and U10065 (N_10065,N_8341,N_7779);
xor U10066 (N_10066,N_7819,N_8334);
and U10067 (N_10067,N_6520,N_9198);
xor U10068 (N_10068,N_8047,N_6531);
xnor U10069 (N_10069,N_7867,N_8803);
nand U10070 (N_10070,N_8285,N_7856);
or U10071 (N_10071,N_8051,N_6724);
nor U10072 (N_10072,N_7731,N_6692);
or U10073 (N_10073,N_7773,N_6261);
nor U10074 (N_10074,N_9083,N_6336);
or U10075 (N_10075,N_8383,N_8057);
nor U10076 (N_10076,N_8300,N_7235);
nand U10077 (N_10077,N_6726,N_8941);
and U10078 (N_10078,N_8952,N_8092);
nor U10079 (N_10079,N_6603,N_8354);
nand U10080 (N_10080,N_6498,N_7788);
or U10081 (N_10081,N_7292,N_7729);
nor U10082 (N_10082,N_6828,N_6687);
and U10083 (N_10083,N_7401,N_6941);
or U10084 (N_10084,N_7041,N_7340);
nor U10085 (N_10085,N_8122,N_9223);
nor U10086 (N_10086,N_8814,N_7178);
nor U10087 (N_10087,N_9185,N_8549);
and U10088 (N_10088,N_6758,N_7063);
nand U10089 (N_10089,N_7700,N_6323);
and U10090 (N_10090,N_8945,N_9367);
or U10091 (N_10091,N_9318,N_8126);
and U10092 (N_10092,N_8385,N_8752);
nor U10093 (N_10093,N_8250,N_8352);
nor U10094 (N_10094,N_8812,N_8105);
or U10095 (N_10095,N_8486,N_9117);
nand U10096 (N_10096,N_7640,N_8801);
nor U10097 (N_10097,N_9041,N_8269);
xor U10098 (N_10098,N_8240,N_8106);
nor U10099 (N_10099,N_7244,N_7584);
nor U10100 (N_10100,N_8194,N_6402);
nor U10101 (N_10101,N_9020,N_6867);
nand U10102 (N_10102,N_9283,N_8840);
nand U10103 (N_10103,N_7530,N_8640);
or U10104 (N_10104,N_6885,N_6521);
or U10105 (N_10105,N_6916,N_8372);
nand U10106 (N_10106,N_7430,N_7196);
and U10107 (N_10107,N_8588,N_8335);
and U10108 (N_10108,N_7370,N_7537);
nand U10109 (N_10109,N_7076,N_8496);
or U10110 (N_10110,N_6835,N_7794);
or U10111 (N_10111,N_8487,N_6518);
nor U10112 (N_10112,N_8773,N_6812);
and U10113 (N_10113,N_6879,N_7467);
or U10114 (N_10114,N_8244,N_8676);
nor U10115 (N_10115,N_7005,N_6390);
and U10116 (N_10116,N_8632,N_7341);
or U10117 (N_10117,N_8023,N_7380);
nor U10118 (N_10118,N_8362,N_8144);
and U10119 (N_10119,N_6849,N_6934);
nor U10120 (N_10120,N_9307,N_9225);
or U10121 (N_10121,N_6797,N_8710);
nor U10122 (N_10122,N_8694,N_7557);
xor U10123 (N_10123,N_8565,N_8067);
or U10124 (N_10124,N_9011,N_7677);
nor U10125 (N_10125,N_7294,N_8564);
xor U10126 (N_10126,N_7935,N_8318);
nand U10127 (N_10127,N_6308,N_9374);
nand U10128 (N_10128,N_9129,N_8278);
nand U10129 (N_10129,N_6643,N_6474);
xnor U10130 (N_10130,N_8845,N_8434);
nand U10131 (N_10131,N_9025,N_6969);
and U10132 (N_10132,N_8243,N_9066);
or U10133 (N_10133,N_7468,N_8955);
nand U10134 (N_10134,N_8083,N_7846);
nor U10135 (N_10135,N_9086,N_7988);
or U10136 (N_10136,N_8821,N_6653);
nor U10137 (N_10137,N_7598,N_7516);
or U10138 (N_10138,N_7979,N_8627);
or U10139 (N_10139,N_6443,N_7541);
nor U10140 (N_10140,N_7479,N_7484);
nor U10141 (N_10141,N_9266,N_8504);
or U10142 (N_10142,N_6597,N_6808);
nor U10143 (N_10143,N_7745,N_7166);
or U10144 (N_10144,N_7579,N_8958);
nand U10145 (N_10145,N_8347,N_8048);
xnor U10146 (N_10146,N_7896,N_8869);
nand U10147 (N_10147,N_6426,N_6781);
nand U10148 (N_10148,N_6399,N_6397);
nor U10149 (N_10149,N_7689,N_8252);
nor U10150 (N_10150,N_7286,N_8965);
nand U10151 (N_10151,N_8804,N_8027);
nor U10152 (N_10152,N_7814,N_6818);
and U10153 (N_10153,N_7017,N_7268);
or U10154 (N_10154,N_7312,N_8507);
nand U10155 (N_10155,N_7749,N_8748);
or U10156 (N_10156,N_6815,N_7823);
nor U10157 (N_10157,N_8493,N_6853);
xnor U10158 (N_10158,N_8344,N_7946);
nor U10159 (N_10159,N_9128,N_8277);
nor U10160 (N_10160,N_8063,N_9054);
nand U10161 (N_10161,N_6802,N_6951);
nand U10162 (N_10162,N_6251,N_7993);
and U10163 (N_10163,N_9344,N_8737);
xnor U10164 (N_10164,N_6319,N_8420);
nand U10165 (N_10165,N_9167,N_9195);
nand U10166 (N_10166,N_6283,N_9131);
nor U10167 (N_10167,N_9263,N_7740);
nand U10168 (N_10168,N_6608,N_7577);
nor U10169 (N_10169,N_7586,N_6331);
xor U10170 (N_10170,N_6624,N_6372);
or U10171 (N_10171,N_6674,N_8931);
xor U10172 (N_10172,N_6891,N_9346);
and U10173 (N_10173,N_8739,N_7511);
nand U10174 (N_10174,N_7243,N_7180);
or U10175 (N_10175,N_8143,N_7564);
nor U10176 (N_10176,N_8381,N_6333);
xnor U10177 (N_10177,N_6268,N_6501);
nor U10178 (N_10178,N_9076,N_7916);
nand U10179 (N_10179,N_7747,N_8227);
and U10180 (N_10180,N_8029,N_8480);
and U10181 (N_10181,N_7899,N_6873);
nand U10182 (N_10182,N_7798,N_9366);
or U10183 (N_10183,N_7216,N_8838);
nand U10184 (N_10184,N_8271,N_8900);
and U10185 (N_10185,N_8058,N_9048);
and U10186 (N_10186,N_8673,N_9147);
nand U10187 (N_10187,N_7241,N_6791);
and U10188 (N_10188,N_9310,N_7273);
and U10189 (N_10189,N_6976,N_7956);
or U10190 (N_10190,N_8764,N_8500);
and U10191 (N_10191,N_9293,N_6749);
and U10192 (N_10192,N_6606,N_8755);
or U10193 (N_10193,N_6509,N_6777);
nor U10194 (N_10194,N_9188,N_8822);
and U10195 (N_10195,N_6939,N_6477);
or U10196 (N_10196,N_6495,N_6894);
nor U10197 (N_10197,N_8323,N_8004);
nor U10198 (N_10198,N_8847,N_9073);
and U10199 (N_10199,N_7390,N_7419);
nand U10200 (N_10200,N_8239,N_8794);
or U10201 (N_10201,N_8153,N_7672);
and U10202 (N_10202,N_8127,N_9347);
and U10203 (N_10203,N_6901,N_9325);
or U10204 (N_10204,N_7008,N_8783);
and U10205 (N_10205,N_7900,N_9341);
or U10206 (N_10206,N_8343,N_8218);
and U10207 (N_10207,N_8098,N_7082);
and U10208 (N_10208,N_8387,N_7397);
and U10209 (N_10209,N_8806,N_6301);
or U10210 (N_10210,N_8130,N_6549);
nor U10211 (N_10211,N_7348,N_9363);
and U10212 (N_10212,N_8956,N_6298);
or U10213 (N_10213,N_9072,N_8477);
nand U10214 (N_10214,N_8735,N_6563);
nand U10215 (N_10215,N_9179,N_9090);
or U10216 (N_10216,N_9262,N_8114);
or U10217 (N_10217,N_9315,N_9319);
nor U10218 (N_10218,N_8963,N_6479);
nand U10219 (N_10219,N_7727,N_8267);
or U10220 (N_10220,N_6536,N_6799);
or U10221 (N_10221,N_6284,N_6750);
nor U10222 (N_10222,N_9328,N_6532);
nand U10223 (N_10223,N_6752,N_7875);
and U10224 (N_10224,N_8638,N_8284);
or U10225 (N_10225,N_7255,N_6968);
nand U10226 (N_10226,N_8438,N_8970);
nor U10227 (N_10227,N_7074,N_6933);
or U10228 (N_10228,N_6279,N_6824);
nand U10229 (N_10229,N_6948,N_7746);
and U10230 (N_10230,N_9099,N_8598);
and U10231 (N_10231,N_7437,N_7331);
nand U10232 (N_10232,N_8964,N_6893);
and U10233 (N_10233,N_9095,N_6998);
nand U10234 (N_10234,N_6591,N_7978);
xor U10235 (N_10235,N_6364,N_8722);
nor U10236 (N_10236,N_8671,N_6695);
nand U10237 (N_10237,N_6569,N_7136);
nand U10238 (N_10238,N_7578,N_6504);
and U10239 (N_10239,N_9181,N_8993);
nand U10240 (N_10240,N_8650,N_8759);
or U10241 (N_10241,N_7424,N_8119);
nor U10242 (N_10242,N_8995,N_8380);
and U10243 (N_10243,N_8075,N_8254);
and U10244 (N_10244,N_7175,N_9287);
or U10245 (N_10245,N_9143,N_8190);
nor U10246 (N_10246,N_9015,N_7409);
or U10247 (N_10247,N_6670,N_8540);
xnor U10248 (N_10248,N_7346,N_7974);
and U10249 (N_10249,N_6594,N_7134);
xnor U10250 (N_10250,N_7879,N_7422);
nor U10251 (N_10251,N_7568,N_9165);
or U10252 (N_10252,N_7765,N_8989);
nand U10253 (N_10253,N_7985,N_8730);
xor U10254 (N_10254,N_7469,N_7720);
or U10255 (N_10255,N_8896,N_6889);
and U10256 (N_10256,N_6365,N_8041);
and U10257 (N_10257,N_9019,N_8450);
or U10258 (N_10258,N_8302,N_7938);
nand U10259 (N_10259,N_7425,N_8944);
or U10260 (N_10260,N_9219,N_8864);
nand U10261 (N_10261,N_7961,N_6424);
nand U10262 (N_10262,N_8933,N_9257);
or U10263 (N_10263,N_8457,N_8976);
xnor U10264 (N_10264,N_6314,N_8366);
or U10265 (N_10265,N_6755,N_8370);
nand U10266 (N_10266,N_8601,N_9091);
or U10267 (N_10267,N_7387,N_6846);
nand U10268 (N_10268,N_9154,N_8719);
nor U10269 (N_10269,N_7190,N_7007);
nor U10270 (N_10270,N_8386,N_9028);
xnor U10271 (N_10271,N_8523,N_8698);
or U10272 (N_10272,N_6487,N_8709);
and U10273 (N_10273,N_8104,N_6671);
nand U10274 (N_10274,N_6524,N_8816);
nor U10275 (N_10275,N_8506,N_7665);
or U10276 (N_10276,N_7526,N_7636);
nand U10277 (N_10277,N_8925,N_6666);
or U10278 (N_10278,N_6480,N_7420);
nor U10279 (N_10279,N_7434,N_8750);
xor U10280 (N_10280,N_8367,N_7099);
or U10281 (N_10281,N_7969,N_7880);
and U10282 (N_10282,N_6541,N_7084);
or U10283 (N_10283,N_9106,N_8515);
nand U10284 (N_10284,N_7748,N_8961);
nand U10285 (N_10285,N_7052,N_6598);
nor U10286 (N_10286,N_8204,N_6987);
or U10287 (N_10287,N_7296,N_8655);
nor U10288 (N_10288,N_7660,N_6481);
nand U10289 (N_10289,N_6264,N_8745);
nor U10290 (N_10290,N_7234,N_6425);
and U10291 (N_10291,N_7003,N_6267);
nor U10292 (N_10292,N_9001,N_7205);
or U10293 (N_10293,N_7306,N_8636);
nand U10294 (N_10294,N_7958,N_6875);
nand U10295 (N_10295,N_7829,N_7024);
xnor U10296 (N_10296,N_8304,N_7458);
and U10297 (N_10297,N_6482,N_9291);
or U10298 (N_10298,N_6970,N_7710);
and U10299 (N_10299,N_8382,N_8241);
or U10300 (N_10300,N_6880,N_8670);
nand U10301 (N_10301,N_7615,N_7187);
and U10302 (N_10302,N_9208,N_6290);
nand U10303 (N_10303,N_6785,N_7690);
nand U10304 (N_10304,N_8292,N_9044);
or U10305 (N_10305,N_9071,N_6300);
and U10306 (N_10306,N_8028,N_8890);
nand U10307 (N_10307,N_8567,N_8183);
nand U10308 (N_10308,N_7174,N_8113);
or U10309 (N_10309,N_8394,N_7795);
nor U10310 (N_10310,N_7122,N_9209);
and U10311 (N_10311,N_7369,N_6779);
or U10312 (N_10312,N_6884,N_9296);
nor U10313 (N_10313,N_8489,N_9271);
nor U10314 (N_10314,N_7558,N_6904);
nor U10315 (N_10315,N_7032,N_7058);
or U10316 (N_10316,N_8897,N_6972);
nand U10317 (N_10317,N_8902,N_9229);
and U10318 (N_10318,N_7011,N_7536);
or U10319 (N_10319,N_7826,N_7882);
and U10320 (N_10320,N_7901,N_6999);
nand U10321 (N_10321,N_7847,N_6829);
nand U10322 (N_10322,N_8910,N_7587);
nor U10323 (N_10323,N_6577,N_7280);
or U10324 (N_10324,N_6705,N_6471);
nor U10325 (N_10325,N_8553,N_6768);
nor U10326 (N_10326,N_9069,N_7493);
and U10327 (N_10327,N_8433,N_7890);
xnor U10328 (N_10328,N_7355,N_8295);
and U10329 (N_10329,N_8509,N_7595);
or U10330 (N_10330,N_7360,N_7692);
nand U10331 (N_10331,N_8772,N_7311);
nand U10332 (N_10332,N_6825,N_8552);
nand U10333 (N_10333,N_6876,N_8810);
nor U10334 (N_10334,N_7693,N_7610);
nand U10335 (N_10335,N_8594,N_6800);
and U10336 (N_10336,N_7386,N_8736);
nor U10337 (N_10337,N_7839,N_8328);
or U10338 (N_10338,N_7763,N_8686);
nor U10339 (N_10339,N_8411,N_8753);
nand U10340 (N_10340,N_9177,N_8929);
and U10341 (N_10341,N_9127,N_6662);
nor U10342 (N_10342,N_9274,N_9107);
and U10343 (N_10343,N_7263,N_6462);
xnor U10344 (N_10344,N_9078,N_9105);
nor U10345 (N_10345,N_7858,N_7250);
or U10346 (N_10346,N_7295,N_7589);
nand U10347 (N_10347,N_6928,N_8080);
and U10348 (N_10348,N_7396,N_6436);
nor U10349 (N_10349,N_6679,N_8883);
or U10350 (N_10350,N_8926,N_8708);
xnor U10351 (N_10351,N_8313,N_8170);
nand U10352 (N_10352,N_7413,N_6917);
nor U10353 (N_10353,N_7548,N_7299);
and U10354 (N_10354,N_7016,N_7508);
nand U10355 (N_10355,N_6672,N_6410);
nor U10356 (N_10356,N_7866,N_8115);
and U10357 (N_10357,N_8718,N_7461);
xnor U10358 (N_10358,N_6494,N_8775);
or U10359 (N_10359,N_6645,N_8279);
or U10360 (N_10360,N_7844,N_7332);
nand U10361 (N_10361,N_7980,N_8604);
nand U10362 (N_10362,N_8805,N_9160);
nand U10363 (N_10363,N_8920,N_8200);
and U10364 (N_10364,N_8160,N_6882);
nor U10365 (N_10365,N_8163,N_8291);
and U10366 (N_10366,N_7784,N_6303);
or U10367 (N_10367,N_7301,N_8408);
or U10368 (N_10368,N_6562,N_7159);
or U10369 (N_10369,N_8046,N_8441);
and U10370 (N_10370,N_7562,N_9014);
nor U10371 (N_10371,N_8017,N_8044);
and U10372 (N_10372,N_7851,N_9186);
and U10373 (N_10373,N_8032,N_8611);
or U10374 (N_10374,N_6256,N_9053);
and U10375 (N_10375,N_8867,N_8651);
nand U10376 (N_10376,N_7797,N_7936);
nand U10377 (N_10377,N_8663,N_7722);
and U10378 (N_10378,N_8591,N_7121);
and U10379 (N_10379,N_7165,N_6586);
and U10380 (N_10380,N_7854,N_8914);
nand U10381 (N_10381,N_8664,N_7948);
xnor U10382 (N_10382,N_6730,N_7220);
nand U10383 (N_10383,N_6871,N_6911);
and U10384 (N_10384,N_7990,N_6772);
and U10385 (N_10385,N_6821,N_6663);
or U10386 (N_10386,N_8508,N_9182);
nor U10387 (N_10387,N_6855,N_9194);
or U10388 (N_10388,N_7394,N_8568);
nand U10389 (N_10389,N_6306,N_8345);
nor U10390 (N_10390,N_7767,N_8997);
or U10391 (N_10391,N_6967,N_7592);
xor U10392 (N_10392,N_6763,N_7883);
and U10393 (N_10393,N_6432,N_9144);
or U10394 (N_10394,N_6291,N_7688);
nand U10395 (N_10395,N_7372,N_6952);
nand U10396 (N_10396,N_7704,N_9213);
or U10397 (N_10397,N_8934,N_7820);
and U10398 (N_10398,N_9017,N_9350);
and U10399 (N_10399,N_7818,N_9029);
or U10400 (N_10400,N_7910,N_6859);
nand U10401 (N_10401,N_7291,N_8136);
and U10402 (N_10402,N_7330,N_7426);
nand U10403 (N_10403,N_7115,N_8786);
nand U10404 (N_10404,N_9031,N_7994);
or U10405 (N_10405,N_6442,N_7544);
nor U10406 (N_10406,N_6327,N_8281);
nand U10407 (N_10407,N_8178,N_6668);
and U10408 (N_10408,N_7476,N_9108);
and U10409 (N_10409,N_7803,N_8359);
and U10410 (N_10410,N_8768,N_9370);
xnor U10411 (N_10411,N_8193,N_8517);
or U10412 (N_10412,N_6782,N_7522);
or U10413 (N_10413,N_7734,N_7553);
and U10414 (N_10414,N_7124,N_8282);
nor U10415 (N_10415,N_6278,N_8577);
and U10416 (N_10416,N_7423,N_7716);
nor U10417 (N_10417,N_9161,N_8866);
nand U10418 (N_10418,N_7171,N_6320);
nand U10419 (N_10419,N_9205,N_9329);
and U10420 (N_10420,N_8297,N_9023);
or U10421 (N_10421,N_6546,N_6539);
nor U10422 (N_10422,N_8356,N_7281);
and U10423 (N_10423,N_8390,N_6403);
nand U10424 (N_10424,N_9242,N_6292);
nor U10425 (N_10425,N_7436,N_9358);
nand U10426 (N_10426,N_7070,N_8371);
or U10427 (N_10427,N_8537,N_8579);
or U10428 (N_10428,N_8851,N_7100);
xnor U10429 (N_10429,N_6311,N_7265);
nand U10430 (N_10430,N_8642,N_8652);
nand U10431 (N_10431,N_6850,N_8230);
or U10432 (N_10432,N_8919,N_7751);
nor U10433 (N_10433,N_9070,N_8214);
nand U10434 (N_10434,N_7126,N_6287);
xor U10435 (N_10435,N_6727,N_7535);
or U10436 (N_10436,N_8892,N_7351);
nor U10437 (N_10437,N_6354,N_7805);
and U10438 (N_10438,N_8824,N_8953);
and U10439 (N_10439,N_8152,N_8695);
nor U10440 (N_10440,N_7950,N_8132);
or U10441 (N_10441,N_8817,N_8470);
or U10442 (N_10442,N_8235,N_7972);
nand U10443 (N_10443,N_8315,N_6573);
or U10444 (N_10444,N_8643,N_7361);
and U10445 (N_10445,N_7093,N_6975);
nor U10446 (N_10446,N_8741,N_8002);
and U10447 (N_10447,N_9369,N_8691);
or U10448 (N_10448,N_6660,N_6588);
or U10449 (N_10449,N_7663,N_9163);
and U10450 (N_10450,N_8365,N_8148);
nor U10451 (N_10451,N_8467,N_7240);
or U10452 (N_10452,N_7923,N_7876);
nand U10453 (N_10453,N_8189,N_6962);
nand U10454 (N_10454,N_6321,N_6349);
xor U10455 (N_10455,N_6985,N_6955);
or U10456 (N_10456,N_6944,N_8100);
nand U10457 (N_10457,N_8894,N_7319);
or U10458 (N_10458,N_8203,N_8407);
nor U10459 (N_10459,N_7195,N_6696);
and U10460 (N_10460,N_6704,N_9322);
nand U10461 (N_10461,N_6980,N_6304);
nor U10462 (N_10462,N_7603,N_6370);
nand U10463 (N_10463,N_7604,N_9123);
nand U10464 (N_10464,N_8288,N_9371);
xnor U10465 (N_10465,N_7465,N_8207);
nor U10466 (N_10466,N_8378,N_7529);
nand U10467 (N_10467,N_8316,N_8317);
nand U10468 (N_10468,N_7077,N_8414);
nor U10469 (N_10469,N_7506,N_6811);
and U10470 (N_10470,N_6260,N_9304);
nor U10471 (N_10471,N_8403,N_7905);
nor U10472 (N_10472,N_8461,N_8384);
nor U10473 (N_10473,N_8990,N_6619);
xor U10474 (N_10474,N_7130,N_8321);
nor U10475 (N_10475,N_8505,N_8171);
nand U10476 (N_10476,N_6366,N_9236);
nand U10477 (N_10477,N_7210,N_7169);
and U10478 (N_10478,N_7039,N_8448);
xor U10479 (N_10479,N_8729,N_7473);
and U10480 (N_10480,N_7492,N_7251);
xnor U10481 (N_10481,N_6362,N_8557);
nand U10482 (N_10482,N_7278,N_9040);
and U10483 (N_10483,N_8479,N_8682);
nor U10484 (N_10484,N_8416,N_8836);
xor U10485 (N_10485,N_8938,N_6356);
nand U10486 (N_10486,N_9197,N_8960);
nand U10487 (N_10487,N_6456,N_7132);
nand U10488 (N_10488,N_9361,N_8839);
nand U10489 (N_10489,N_8495,N_6676);
nand U10490 (N_10490,N_6854,N_8600);
or U10491 (N_10491,N_8943,N_8532);
nand U10492 (N_10492,N_8413,N_7581);
and U10493 (N_10493,N_7645,N_6618);
and U10494 (N_10494,N_9012,N_6628);
nor U10495 (N_10495,N_7976,N_7588);
nand U10496 (N_10496,N_8112,N_8516);
or U10497 (N_10497,N_7019,N_7116);
nor U10498 (N_10498,N_7738,N_8220);
nand U10499 (N_10499,N_7565,N_6439);
and U10500 (N_10500,N_8429,N_8273);
or U10501 (N_10501,N_9321,N_6851);
nand U10502 (N_10502,N_8374,N_6380);
and U10503 (N_10503,N_7229,N_7567);
or U10504 (N_10504,N_6383,N_8981);
nor U10505 (N_10505,N_9125,N_8706);
or U10506 (N_10506,N_7997,N_6398);
or U10507 (N_10507,N_7490,N_9220);
and U10508 (N_10508,N_8306,N_8518);
nand U10509 (N_10509,N_6996,N_7054);
and U10510 (N_10510,N_6809,N_7862);
nand U10511 (N_10511,N_7140,N_6465);
nor U10512 (N_10512,N_7057,N_8405);
and U10513 (N_10513,N_8999,N_8859);
or U10514 (N_10514,N_8449,N_6592);
nor U10515 (N_10515,N_8887,N_7091);
nand U10516 (N_10516,N_9320,N_8898);
nand U10517 (N_10517,N_9231,N_8587);
or U10518 (N_10518,N_8213,N_9021);
nand U10519 (N_10519,N_6607,N_7309);
nand U10520 (N_10520,N_6664,N_9061);
nor U10521 (N_10521,N_8528,N_6947);
or U10522 (N_10522,N_6351,N_6545);
nor U10523 (N_10523,N_7321,N_6633);
nor U10524 (N_10524,N_8401,N_8996);
nand U10525 (N_10525,N_8940,N_8141);
nor U10526 (N_10526,N_8172,N_7267);
and U10527 (N_10527,N_8728,N_8184);
nor U10528 (N_10528,N_7488,N_6548);
nor U10529 (N_10529,N_8703,N_8539);
nor U10530 (N_10530,N_8697,N_7960);
nor U10531 (N_10531,N_7855,N_6919);
nand U10532 (N_10532,N_8179,N_8223);
or U10533 (N_10533,N_8458,N_7547);
or U10534 (N_10534,N_9343,N_7596);
and U10535 (N_10535,N_7758,N_7850);
nand U10536 (N_10536,N_9067,N_8762);
and U10537 (N_10537,N_7743,N_7222);
nand U10538 (N_10538,N_7213,N_7248);
nor U10539 (N_10539,N_7591,N_8157);
nand U10540 (N_10540,N_6523,N_7106);
nand U10541 (N_10541,N_8234,N_6908);
nor U10542 (N_10542,N_7103,N_8592);
nor U10543 (N_10543,N_7406,N_7723);
and U10544 (N_10544,N_9357,N_7271);
nand U10545 (N_10545,N_8936,N_7489);
or U10546 (N_10546,N_7167,N_9215);
nor U10547 (N_10547,N_6317,N_9336);
and U10548 (N_10548,N_7272,N_8265);
nor U10549 (N_10549,N_7656,N_8715);
nand U10550 (N_10550,N_8720,N_6490);
and U10551 (N_10551,N_8538,N_7534);
xor U10552 (N_10552,N_8078,N_8510);
xor U10553 (N_10553,N_8364,N_6760);
nor U10554 (N_10554,N_8392,N_8089);
and U10555 (N_10555,N_7965,N_6485);
or U10556 (N_10556,N_7627,N_6596);
nand U10557 (N_10557,N_8442,N_7933);
nand U10558 (N_10558,N_7824,N_8572);
xor U10559 (N_10559,N_6486,N_9030);
nand U10560 (N_10560,N_9326,N_7018);
nand U10561 (N_10561,N_7075,N_6784);
and U10562 (N_10562,N_7432,N_6444);
or U10563 (N_10563,N_8437,N_6547);
nor U10564 (N_10564,N_7733,N_8033);
or U10565 (N_10565,N_7674,N_7666);
nand U10566 (N_10566,N_6773,N_8629);
or U10567 (N_10567,N_7310,N_8667);
and U10568 (N_10568,N_6431,N_8680);
or U10569 (N_10569,N_7357,N_9285);
or U10570 (N_10570,N_7154,N_8639);
nor U10571 (N_10571,N_7572,N_8573);
or U10572 (N_10572,N_6929,N_7886);
or U10573 (N_10573,N_8542,N_8832);
nand U10574 (N_10574,N_7428,N_8702);
nand U10575 (N_10575,N_9355,N_7279);
and U10576 (N_10576,N_8443,N_7389);
or U10577 (N_10577,N_8462,N_8802);
or U10578 (N_10578,N_7207,N_8108);
nand U10579 (N_10579,N_6978,N_9360);
and U10580 (N_10580,N_7915,N_8142);
and U10581 (N_10581,N_6938,N_9166);
and U10582 (N_10582,N_6794,N_6534);
nand U10583 (N_10583,N_9234,N_7715);
or U10584 (N_10584,N_6525,N_6689);
xor U10585 (N_10585,N_8647,N_7801);
and U10586 (N_10586,N_7366,N_7441);
nand U10587 (N_10587,N_6609,N_7148);
nor U10588 (N_10588,N_6922,N_7914);
nand U10589 (N_10589,N_7223,N_8818);
and U10590 (N_10590,N_7293,N_8654);
or U10591 (N_10591,N_8917,N_6454);
nand U10592 (N_10592,N_9337,N_6902);
nand U10593 (N_10593,N_7408,N_7865);
or U10594 (N_10594,N_8336,N_7816);
or U10595 (N_10595,N_7724,N_8880);
or U10596 (N_10596,N_9008,N_8779);
or U10597 (N_10597,N_7259,N_7601);
xnor U10598 (N_10598,N_6954,N_6629);
nand U10599 (N_10599,N_8678,N_8330);
nor U10600 (N_10600,N_8909,N_8829);
or U10601 (N_10601,N_6634,N_9089);
or U10602 (N_10602,N_7713,N_8888);
xnor U10603 (N_10603,N_8672,N_8225);
and U10604 (N_10604,N_6343,N_6691);
nand U10605 (N_10605,N_8499,N_7812);
nor U10606 (N_10606,N_9094,N_6924);
and U10607 (N_10607,N_8072,N_6415);
and U10608 (N_10608,N_8050,N_7831);
nor U10609 (N_10609,N_8338,N_7260);
nor U10610 (N_10610,N_7718,N_7849);
or U10611 (N_10611,N_8042,N_7509);
or U10612 (N_10612,N_8580,N_7881);
nand U10613 (N_10613,N_8524,N_8716);
nand U10614 (N_10614,N_7906,N_7374);
and U10615 (N_10615,N_7110,N_7145);
nand U10616 (N_10616,N_6352,N_7086);
or U10617 (N_10617,N_7327,N_7986);
or U10618 (N_10618,N_7282,N_6654);
or U10619 (N_10619,N_7375,N_8124);
or U10620 (N_10620,N_8264,N_8111);
nor U10621 (N_10621,N_9135,N_8307);
or U10622 (N_10622,N_7884,N_9110);
nor U10623 (N_10623,N_6832,N_7903);
nor U10624 (N_10624,N_7237,N_9081);
xor U10625 (N_10625,N_9122,N_9203);
nor U10626 (N_10626,N_6700,N_6746);
xor U10627 (N_10627,N_9148,N_6386);
and U10628 (N_10628,N_6819,N_8761);
and U10629 (N_10629,N_8026,N_7215);
nor U10630 (N_10630,N_8357,N_9022);
nand U10631 (N_10631,N_6355,N_9112);
and U10632 (N_10632,N_8948,N_8609);
or U10633 (N_10633,N_7571,N_8015);
nor U10634 (N_10634,N_6282,N_6419);
or U10635 (N_10635,N_7888,N_7497);
or U10636 (N_10636,N_6489,N_9204);
nand U10637 (N_10637,N_6983,N_8181);
and U10638 (N_10638,N_6842,N_7669);
nand U10639 (N_10639,N_6400,N_7766);
nor U10640 (N_10640,N_8439,N_8780);
nor U10641 (N_10641,N_6887,N_6708);
nand U10642 (N_10642,N_6427,N_8166);
and U10643 (N_10643,N_8968,N_6652);
nor U10644 (N_10644,N_8016,N_6258);
or U10645 (N_10645,N_7868,N_7957);
nand U10646 (N_10646,N_6638,N_6814);
nor U10647 (N_10647,N_8527,N_7813);
and U10648 (N_10648,N_7464,N_6273);
or U10649 (N_10649,N_8373,N_8581);
nand U10650 (N_10650,N_7410,N_8830);
xnor U10651 (N_10651,N_7653,N_6512);
and U10652 (N_10652,N_6593,N_6964);
xnor U10653 (N_10653,N_7137,N_7996);
nor U10654 (N_10654,N_7421,N_6388);
xor U10655 (N_10655,N_6538,N_8205);
and U10656 (N_10656,N_9103,N_8117);
or U10657 (N_10657,N_7404,N_8644);
nor U10658 (N_10658,N_6348,N_8834);
xor U10659 (N_10659,N_6472,N_7870);
nor U10660 (N_10660,N_9193,N_7065);
and U10661 (N_10661,N_7654,N_8877);
or U10662 (N_10662,N_6888,N_7247);
or U10663 (N_10663,N_6783,N_8488);
and U10664 (N_10664,N_7303,N_9252);
or U10665 (N_10665,N_8835,N_8093);
or U10666 (N_10666,N_7450,N_6731);
xor U10667 (N_10667,N_7783,N_8346);
nor U10668 (N_10668,N_9338,N_7975);
nor U10669 (N_10669,N_9349,N_7290);
xnor U10670 (N_10670,N_8789,N_8260);
and U10671 (N_10671,N_8566,N_6703);
nand U10672 (N_10672,N_7335,N_8796);
or U10673 (N_10673,N_8397,N_6488);
and U10674 (N_10674,N_9200,N_8511);
nand U10675 (N_10675,N_6857,N_7162);
nor U10676 (N_10676,N_6986,N_6745);
nand U10677 (N_10677,N_6651,N_8238);
xor U10678 (N_10678,N_6698,N_8563);
nor U10679 (N_10679,N_8733,N_8668);
or U10680 (N_10680,N_7060,N_7759);
nor U10681 (N_10681,N_8863,N_8340);
or U10682 (N_10682,N_7563,N_8503);
nor U10683 (N_10683,N_7928,N_8713);
and U10684 (N_10684,N_6775,N_9192);
nand U10685 (N_10685,N_7635,N_8666);
nand U10686 (N_10686,N_9308,N_7252);
or U10687 (N_10687,N_7614,N_8071);
and U10688 (N_10688,N_7921,N_6511);
nor U10689 (N_10689,N_9109,N_7754);
and U10690 (N_10690,N_9187,N_7892);
and U10691 (N_10691,N_9157,N_8202);
or U10692 (N_10692,N_7662,N_8168);
and U10693 (N_10693,N_7648,N_9101);
and U10694 (N_10694,N_8472,N_7650);
and U10695 (N_10695,N_8846,N_8544);
and U10696 (N_10696,N_9261,N_6995);
or U10697 (N_10697,N_7173,N_8469);
or U10698 (N_10698,N_8091,N_6945);
or U10699 (N_10699,N_8561,N_7770);
nand U10700 (N_10700,N_7705,N_7283);
nand U10701 (N_10701,N_7519,N_7566);
nor U10702 (N_10702,N_6639,N_6412);
nor U10703 (N_10703,N_7878,N_7861);
or U10704 (N_10704,N_6376,N_7208);
nor U10705 (N_10705,N_8076,N_7338);
nor U10706 (N_10706,N_7182,N_9295);
or U10707 (N_10707,N_6714,N_8399);
nand U10708 (N_10708,N_7540,N_8192);
or U10709 (N_10709,N_7202,N_6441);
or U10710 (N_10710,N_7755,N_7664);
nand U10711 (N_10711,N_8865,N_7107);
nand U10712 (N_10712,N_8208,N_7485);
nor U10713 (N_10713,N_6346,N_8475);
nand U10714 (N_10714,N_7741,N_7009);
nor U10715 (N_10715,N_7304,N_7230);
or U10716 (N_10716,N_6554,N_7446);
nor U10717 (N_10717,N_8548,N_8339);
xnor U10718 (N_10718,N_9313,N_8059);
or U10719 (N_10719,N_7046,N_6649);
and U10720 (N_10720,N_7056,N_6502);
and U10721 (N_10721,N_6720,N_7061);
or U10722 (N_10722,N_6414,N_8228);
nand U10723 (N_10723,N_9281,N_8236);
and U10724 (N_10724,N_7347,N_6837);
nor U10725 (N_10725,N_7827,N_8013);
nor U10726 (N_10726,N_7307,N_8229);
and U10727 (N_10727,N_8331,N_7685);
and U10728 (N_10728,N_6723,N_7079);
or U10729 (N_10729,N_8162,N_6275);
nor U10730 (N_10730,N_9057,N_7922);
or U10731 (N_10731,N_7863,N_6702);
or U10732 (N_10732,N_8261,N_7651);
and U10733 (N_10733,N_8221,N_8237);
and U10734 (N_10734,N_8535,N_7619);
nand U10735 (N_10735,N_6930,N_6862);
or U10736 (N_10736,N_8501,N_7869);
nor U10737 (N_10737,N_9332,N_6913);
and U10738 (N_10738,N_9279,N_8974);
nor U10739 (N_10739,N_8066,N_7073);
or U10740 (N_10740,N_8299,N_6411);
nor U10741 (N_10741,N_7435,N_7036);
and U10742 (N_10742,N_7982,N_8763);
nor U10743 (N_10743,N_6732,N_7362);
nand U10744 (N_10744,N_7608,N_8633);
xor U10745 (N_10745,N_7412,N_8922);
nor U10746 (N_10746,N_7123,N_8222);
and U10747 (N_10747,N_6305,N_7893);
or U10748 (N_10748,N_7333,N_8155);
or U10749 (N_10749,N_9074,N_8994);
nand U10750 (N_10750,N_7657,N_9064);
nand U10751 (N_10751,N_7622,N_6625);
nor U10752 (N_10752,N_7546,N_9365);
nand U10753 (N_10753,N_9250,N_8360);
or U10754 (N_10754,N_6280,N_8398);
or U10755 (N_10755,N_6841,N_8795);
nor U10756 (N_10756,N_8721,N_8685);
or U10757 (N_10757,N_7128,N_9051);
or U10758 (N_10758,N_8498,N_7498);
or U10759 (N_10759,N_8622,N_9259);
or U10760 (N_10760,N_6683,N_7807);
nor U10761 (N_10761,N_7561,N_6335);
nand U10762 (N_10762,N_8094,N_7203);
and U10763 (N_10763,N_8007,N_7452);
nor U10764 (N_10764,N_8333,N_7179);
nand U10765 (N_10765,N_7756,N_6381);
nand U10766 (N_10766,N_7129,N_6537);
and U10767 (N_10767,N_8712,N_7873);
or U10768 (N_10768,N_7551,N_8195);
xor U10769 (N_10769,N_8263,N_8879);
nor U10770 (N_10770,N_6659,N_6466);
or U10771 (N_10771,N_8649,N_6892);
and U10772 (N_10772,N_9217,N_8743);
nand U10773 (N_10773,N_7524,N_7543);
nor U10774 (N_10774,N_7513,N_6932);
or U10775 (N_10775,N_9254,N_7841);
and U10776 (N_10776,N_7284,N_6353);
or U10777 (N_10777,N_7618,N_7433);
or U10778 (N_10778,N_9170,N_8828);
xor U10779 (N_10779,N_8717,N_8096);
xor U10780 (N_10780,N_8792,N_7083);
nor U10781 (N_10781,N_8545,N_7228);
or U10782 (N_10782,N_7318,N_8841);
xor U10783 (N_10783,N_7626,N_7864);
nor U10784 (N_10784,N_9146,N_8610);
nand U10785 (N_10785,N_6669,N_6678);
xnor U10786 (N_10786,N_6438,N_8519);
and U10787 (N_10787,N_9248,N_6558);
nand U10788 (N_10788,N_6981,N_7308);
and U10789 (N_10789,N_7427,N_8419);
xor U10790 (N_10790,N_6505,N_7256);
and U10791 (N_10791,N_8973,N_9138);
nand U10792 (N_10792,N_7682,N_8329);
and U10793 (N_10793,N_7156,N_8605);
nor U10794 (N_10794,N_6667,N_7800);
nand U10795 (N_10795,N_7675,N_8799);
nor U10796 (N_10796,N_8616,N_6294);
nor U10797 (N_10797,N_6994,N_8310);
nor U10798 (N_10798,N_7533,N_7617);
nand U10799 (N_10799,N_9121,N_7998);
or U10800 (N_10800,N_8164,N_6574);
xnor U10801 (N_10801,N_6409,N_9317);
nor U10802 (N_10802,N_8689,N_6991);
nor U10803 (N_10803,N_7201,N_8145);
nor U10804 (N_10804,N_9245,N_6334);
or U10805 (N_10805,N_6622,N_9183);
nor U10806 (N_10806,N_7376,N_7104);
nor U10807 (N_10807,N_7633,N_7170);
nand U10808 (N_10808,N_7038,N_7494);
nor U10809 (N_10809,N_8211,N_7131);
and U10810 (N_10810,N_9305,N_6743);
or U10811 (N_10811,N_6675,N_6813);
nand U10812 (N_10812,N_6253,N_6433);
nor U10813 (N_10813,N_6587,N_8602);
and U10814 (N_10814,N_8988,N_9173);
nand U10815 (N_10815,N_6774,N_6737);
nand U10816 (N_10816,N_6872,N_6931);
and U10817 (N_10817,N_7270,N_8308);
and U10818 (N_10818,N_8444,N_9227);
nand U10819 (N_10819,N_6422,N_8175);
nor U10820 (N_10820,N_7227,N_8090);
nor U10821 (N_10821,N_6665,N_9226);
and U10822 (N_10822,N_7804,N_9058);
and U10823 (N_10823,N_7987,N_6599);
or U10824 (N_10824,N_6445,N_7322);
nor U10825 (N_10825,N_8427,N_7649);
nand U10826 (N_10826,N_9176,N_6817);
nand U10827 (N_10827,N_7163,N_8586);
nor U10828 (N_10828,N_6413,N_6307);
and U10829 (N_10829,N_6535,N_6604);
nor U10830 (N_10830,N_8621,N_7639);
and U10831 (N_10831,N_6540,N_8886);
nand U10832 (N_10832,N_8546,N_7114);
nand U10833 (N_10833,N_8125,N_8049);
and U10834 (N_10834,N_8631,N_8740);
xnor U10835 (N_10835,N_6699,N_8665);
nor U10836 (N_10836,N_8862,N_6658);
and U10837 (N_10837,N_7605,N_6457);
and U10838 (N_10838,N_7068,N_6499);
or U10839 (N_10839,N_8776,N_7853);
nor U10840 (N_10840,N_7276,N_7925);
nor U10841 (N_10841,N_6688,N_6729);
nor U10842 (N_10842,N_7620,N_8635);
nand U10843 (N_10843,N_7616,N_6848);
nor U10844 (N_10844,N_8088,N_7285);
and U10845 (N_10845,N_7144,N_9010);
or U10846 (N_10846,N_6552,N_8251);
and U10847 (N_10847,N_7151,N_7939);
nand U10848 (N_10848,N_7857,N_6725);
nand U10849 (N_10849,N_6396,N_9265);
or U10850 (N_10850,N_8767,N_6614);
xor U10851 (N_10851,N_6510,N_7732);
and U10852 (N_10852,N_6937,N_8045);
nor U10853 (N_10853,N_8379,N_8021);
and U10854 (N_10854,N_8266,N_9050);
nor U10855 (N_10855,N_8400,N_7607);
and U10856 (N_10856,N_9351,N_6500);
nand U10857 (N_10857,N_6363,N_8634);
nor U10858 (N_10858,N_7810,N_6338);
or U10859 (N_10859,N_9206,N_6963);
nor U10860 (N_10860,N_8947,N_8657);
and U10861 (N_10861,N_9159,N_9132);
xnor U10862 (N_10862,N_7457,N_7752);
nand U10863 (N_10863,N_9333,N_7920);
and U10864 (N_10864,N_8358,N_8911);
nand U10865 (N_10865,N_7049,N_7439);
nand U10866 (N_10866,N_6497,N_6564);
and U10867 (N_10867,N_9218,N_7349);
nor U10868 (N_10868,N_7040,N_7775);
or U10869 (N_10869,N_6468,N_7440);
and U10870 (N_10870,N_8637,N_6475);
nand U10871 (N_10871,N_6281,N_7709);
xnor U10872 (N_10872,N_8809,N_8751);
xnor U10873 (N_10873,N_6581,N_7780);
nand U10874 (N_10874,N_7777,N_6617);
nor U10875 (N_10875,N_7632,N_6640);
nand U10876 (N_10876,N_7193,N_8533);
or U10877 (N_10877,N_9169,N_7300);
or U10878 (N_10878,N_6682,N_8003);
nand U10879 (N_10879,N_9373,N_6557);
or U10880 (N_10880,N_6716,N_9334);
and U10881 (N_10881,N_8158,N_8583);
nand U10882 (N_10882,N_6757,N_6858);
nor U10883 (N_10883,N_7316,N_8813);
or U10884 (N_10884,N_6611,N_9042);
and U10885 (N_10885,N_6452,N_6515);
nand U10886 (N_10886,N_7287,N_8771);
and U10887 (N_10887,N_6395,N_7911);
and U10888 (N_10888,N_9092,N_8377);
and U10889 (N_10889,N_6753,N_7659);
nor U10890 (N_10890,N_8734,N_9214);
or U10891 (N_10891,N_6616,N_7772);
nor U10892 (N_10892,N_8249,N_6641);
and U10893 (N_10893,N_6806,N_8626);
nand U10894 (N_10894,N_7825,N_9224);
and U10895 (N_10895,N_7186,N_8861);
nand U10896 (N_10896,N_7470,N_7157);
nor U10897 (N_10897,N_8191,N_6712);
nand U10898 (N_10898,N_8177,N_9199);
nand U10899 (N_10899,N_6881,N_8742);
xor U10900 (N_10900,N_7365,N_8852);
nor U10901 (N_10901,N_9327,N_8747);
nor U10902 (N_10902,N_8787,N_7023);
and U10903 (N_10903,N_7520,N_6315);
and U10904 (N_10904,N_7161,N_9212);
and U10905 (N_10905,N_9240,N_7808);
and U10906 (N_10906,N_7192,N_9153);
and U10907 (N_10907,N_6736,N_6582);
and U10908 (N_10908,N_6830,N_9126);
nor U10909 (N_10909,N_7711,N_6718);
xor U10910 (N_10910,N_9140,N_7877);
xor U10911 (N_10911,N_7416,N_7183);
nand U10912 (N_10912,N_6339,N_8785);
or U10913 (N_10913,N_7217,N_7231);
nand U10914 (N_10914,N_8765,N_9299);
and U10915 (N_10915,N_7679,N_8541);
and U10916 (N_10916,N_7778,N_6506);
nor U10917 (N_10917,N_6570,N_9270);
and U10918 (N_10918,N_9152,N_8215);
xor U10919 (N_10919,N_7576,N_6739);
xor U10920 (N_10920,N_6748,N_7646);
and U10921 (N_10921,N_8681,N_9155);
nor U10922 (N_10922,N_8283,N_7081);
and U10923 (N_10923,N_8893,N_6721);
and U10924 (N_10924,N_8784,N_9286);
and U10925 (N_10925,N_8468,N_7253);
or U10926 (N_10926,N_6681,N_7840);
nor U10927 (N_10927,N_8913,N_8562);
and U10928 (N_10928,N_8908,N_8700);
nand U10929 (N_10929,N_8034,N_8705);
xor U10930 (N_10930,N_6615,N_7786);
nor U10931 (N_10931,N_8402,N_8198);
nand U10932 (N_10932,N_6896,N_8110);
nand U10933 (N_10933,N_9164,N_9005);
xnor U10934 (N_10934,N_6701,N_6886);
nand U10935 (N_10935,N_6795,N_8884);
nor U10936 (N_10936,N_8287,N_9080);
or U10937 (N_10937,N_9115,N_6261);
and U10938 (N_10938,N_7773,N_7743);
and U10939 (N_10939,N_8495,N_6724);
xor U10940 (N_10940,N_6327,N_6544);
nand U10941 (N_10941,N_9048,N_8954);
and U10942 (N_10942,N_8731,N_8173);
and U10943 (N_10943,N_7833,N_6575);
nand U10944 (N_10944,N_7681,N_8136);
nand U10945 (N_10945,N_8800,N_7338);
nand U10946 (N_10946,N_7624,N_8015);
or U10947 (N_10947,N_8366,N_7441);
xor U10948 (N_10948,N_8351,N_9263);
xnor U10949 (N_10949,N_7029,N_6900);
and U10950 (N_10950,N_7652,N_9160);
xor U10951 (N_10951,N_8945,N_9171);
xor U10952 (N_10952,N_7716,N_8754);
and U10953 (N_10953,N_8501,N_7711);
nand U10954 (N_10954,N_8483,N_8065);
nor U10955 (N_10955,N_6625,N_6389);
and U10956 (N_10956,N_6511,N_9092);
nor U10957 (N_10957,N_7061,N_8190);
and U10958 (N_10958,N_8357,N_8546);
nor U10959 (N_10959,N_8057,N_6542);
xnor U10960 (N_10960,N_6700,N_7586);
and U10961 (N_10961,N_7473,N_8683);
or U10962 (N_10962,N_8262,N_7008);
or U10963 (N_10963,N_9106,N_8262);
xor U10964 (N_10964,N_8301,N_9233);
or U10965 (N_10965,N_6268,N_9058);
or U10966 (N_10966,N_6438,N_8168);
xnor U10967 (N_10967,N_6535,N_6567);
nor U10968 (N_10968,N_7094,N_6588);
nand U10969 (N_10969,N_7708,N_6956);
and U10970 (N_10970,N_6678,N_8693);
and U10971 (N_10971,N_9025,N_9231);
and U10972 (N_10972,N_7124,N_6399);
nor U10973 (N_10973,N_7743,N_8200);
nand U10974 (N_10974,N_7029,N_8265);
nor U10975 (N_10975,N_6349,N_7301);
or U10976 (N_10976,N_9033,N_8759);
and U10977 (N_10977,N_8103,N_8040);
and U10978 (N_10978,N_8464,N_7821);
nand U10979 (N_10979,N_7732,N_7593);
and U10980 (N_10980,N_6936,N_8390);
or U10981 (N_10981,N_8919,N_7625);
xor U10982 (N_10982,N_7154,N_7425);
and U10983 (N_10983,N_7129,N_7682);
nor U10984 (N_10984,N_7241,N_6592);
and U10985 (N_10985,N_7007,N_7949);
and U10986 (N_10986,N_8464,N_6301);
nand U10987 (N_10987,N_7256,N_7821);
or U10988 (N_10988,N_8113,N_6908);
or U10989 (N_10989,N_6467,N_6494);
nand U10990 (N_10990,N_8861,N_8562);
nor U10991 (N_10991,N_7763,N_7827);
or U10992 (N_10992,N_7350,N_8482);
or U10993 (N_10993,N_8765,N_8086);
and U10994 (N_10994,N_6732,N_8373);
and U10995 (N_10995,N_6651,N_8772);
or U10996 (N_10996,N_8667,N_7823);
nand U10997 (N_10997,N_6664,N_7603);
and U10998 (N_10998,N_7277,N_7144);
nor U10999 (N_10999,N_7001,N_7099);
or U11000 (N_11000,N_9242,N_7057);
or U11001 (N_11001,N_7264,N_8849);
or U11002 (N_11002,N_8235,N_6390);
xnor U11003 (N_11003,N_8363,N_6819);
xnor U11004 (N_11004,N_7941,N_7264);
nand U11005 (N_11005,N_7604,N_7884);
xnor U11006 (N_11006,N_9208,N_8803);
or U11007 (N_11007,N_6804,N_6622);
nor U11008 (N_11008,N_8942,N_8071);
nand U11009 (N_11009,N_9228,N_7894);
nor U11010 (N_11010,N_8098,N_6811);
and U11011 (N_11011,N_7797,N_7873);
or U11012 (N_11012,N_6491,N_6701);
and U11013 (N_11013,N_7234,N_6984);
nor U11014 (N_11014,N_6704,N_6605);
or U11015 (N_11015,N_8807,N_8826);
nor U11016 (N_11016,N_9182,N_6641);
nand U11017 (N_11017,N_9230,N_7590);
or U11018 (N_11018,N_8238,N_6487);
and U11019 (N_11019,N_6958,N_8873);
and U11020 (N_11020,N_9363,N_6423);
nand U11021 (N_11021,N_8514,N_8030);
or U11022 (N_11022,N_7578,N_7923);
and U11023 (N_11023,N_8864,N_8225);
and U11024 (N_11024,N_7237,N_6419);
nand U11025 (N_11025,N_7986,N_8722);
and U11026 (N_11026,N_6575,N_9230);
nand U11027 (N_11027,N_6363,N_7778);
or U11028 (N_11028,N_8508,N_8359);
or U11029 (N_11029,N_8330,N_7639);
nor U11030 (N_11030,N_6430,N_7195);
and U11031 (N_11031,N_6877,N_8241);
nand U11032 (N_11032,N_8961,N_9268);
and U11033 (N_11033,N_6856,N_7547);
nand U11034 (N_11034,N_8804,N_6791);
nor U11035 (N_11035,N_8522,N_6888);
and U11036 (N_11036,N_6479,N_7555);
or U11037 (N_11037,N_8223,N_9239);
nand U11038 (N_11038,N_7015,N_7164);
nor U11039 (N_11039,N_8859,N_7016);
nor U11040 (N_11040,N_8556,N_8802);
nand U11041 (N_11041,N_6786,N_6567);
or U11042 (N_11042,N_6520,N_7642);
nand U11043 (N_11043,N_7912,N_9053);
or U11044 (N_11044,N_8717,N_8449);
nor U11045 (N_11045,N_6618,N_7330);
nand U11046 (N_11046,N_7039,N_6462);
nand U11047 (N_11047,N_8490,N_7554);
or U11048 (N_11048,N_8873,N_6458);
nand U11049 (N_11049,N_6943,N_7842);
nor U11050 (N_11050,N_9134,N_6981);
nand U11051 (N_11051,N_9203,N_8400);
or U11052 (N_11052,N_6336,N_9061);
nor U11053 (N_11053,N_8031,N_8167);
and U11054 (N_11054,N_6734,N_7547);
and U11055 (N_11055,N_8692,N_7991);
xor U11056 (N_11056,N_6370,N_8644);
nor U11057 (N_11057,N_6533,N_6470);
nand U11058 (N_11058,N_8172,N_8828);
nand U11059 (N_11059,N_7954,N_9178);
and U11060 (N_11060,N_8367,N_9255);
or U11061 (N_11061,N_7959,N_8802);
or U11062 (N_11062,N_8742,N_7574);
nor U11063 (N_11063,N_9106,N_9133);
or U11064 (N_11064,N_8308,N_7886);
or U11065 (N_11065,N_8516,N_6888);
xnor U11066 (N_11066,N_8845,N_7307);
nor U11067 (N_11067,N_9118,N_8763);
nand U11068 (N_11068,N_6860,N_7586);
nand U11069 (N_11069,N_7145,N_6587);
and U11070 (N_11070,N_6753,N_7329);
xnor U11071 (N_11071,N_8506,N_8808);
nor U11072 (N_11072,N_7342,N_9168);
nand U11073 (N_11073,N_7528,N_6265);
xnor U11074 (N_11074,N_6986,N_6519);
or U11075 (N_11075,N_6526,N_8548);
nor U11076 (N_11076,N_8088,N_8006);
nor U11077 (N_11077,N_8443,N_7785);
nor U11078 (N_11078,N_7717,N_8162);
or U11079 (N_11079,N_7340,N_7272);
or U11080 (N_11080,N_8077,N_8911);
xor U11081 (N_11081,N_6562,N_7307);
or U11082 (N_11082,N_7524,N_7893);
or U11083 (N_11083,N_7660,N_7131);
nor U11084 (N_11084,N_7394,N_6909);
xor U11085 (N_11085,N_8127,N_8929);
and U11086 (N_11086,N_9050,N_8026);
or U11087 (N_11087,N_8724,N_6586);
or U11088 (N_11088,N_9049,N_8424);
or U11089 (N_11089,N_7639,N_9088);
and U11090 (N_11090,N_6405,N_7358);
xor U11091 (N_11091,N_9164,N_7272);
xor U11092 (N_11092,N_8605,N_7883);
nand U11093 (N_11093,N_8343,N_8650);
and U11094 (N_11094,N_8853,N_6255);
nand U11095 (N_11095,N_7959,N_9277);
nor U11096 (N_11096,N_9164,N_7189);
or U11097 (N_11097,N_7749,N_8024);
nor U11098 (N_11098,N_9002,N_6465);
and U11099 (N_11099,N_8810,N_8842);
xor U11100 (N_11100,N_6529,N_8240);
and U11101 (N_11101,N_6637,N_6353);
nand U11102 (N_11102,N_6657,N_7337);
and U11103 (N_11103,N_8699,N_6704);
nor U11104 (N_11104,N_9155,N_8913);
nor U11105 (N_11105,N_7822,N_8209);
or U11106 (N_11106,N_8163,N_8274);
or U11107 (N_11107,N_8599,N_8246);
nand U11108 (N_11108,N_7786,N_9318);
or U11109 (N_11109,N_8270,N_7746);
and U11110 (N_11110,N_6510,N_7999);
xnor U11111 (N_11111,N_7845,N_8522);
nor U11112 (N_11112,N_8776,N_7230);
and U11113 (N_11113,N_7644,N_7078);
nand U11114 (N_11114,N_6914,N_7746);
xnor U11115 (N_11115,N_8310,N_8267);
nor U11116 (N_11116,N_9334,N_8647);
or U11117 (N_11117,N_7367,N_6507);
xnor U11118 (N_11118,N_6418,N_6631);
nor U11119 (N_11119,N_7983,N_7323);
nor U11120 (N_11120,N_6849,N_6493);
nand U11121 (N_11121,N_7567,N_8505);
xor U11122 (N_11122,N_7489,N_9035);
nor U11123 (N_11123,N_8876,N_6759);
and U11124 (N_11124,N_6339,N_9341);
xor U11125 (N_11125,N_7391,N_8063);
and U11126 (N_11126,N_8861,N_7756);
and U11127 (N_11127,N_6764,N_9177);
and U11128 (N_11128,N_7265,N_7961);
and U11129 (N_11129,N_7339,N_6735);
and U11130 (N_11130,N_6349,N_7064);
and U11131 (N_11131,N_7241,N_9237);
nor U11132 (N_11132,N_8796,N_9230);
nor U11133 (N_11133,N_9245,N_7175);
or U11134 (N_11134,N_7517,N_7177);
nor U11135 (N_11135,N_8003,N_8806);
nor U11136 (N_11136,N_7908,N_8433);
xor U11137 (N_11137,N_8601,N_8863);
or U11138 (N_11138,N_9207,N_8923);
and U11139 (N_11139,N_9212,N_6606);
or U11140 (N_11140,N_7577,N_8458);
nand U11141 (N_11141,N_7205,N_6971);
nand U11142 (N_11142,N_8575,N_7424);
xor U11143 (N_11143,N_6297,N_7082);
nor U11144 (N_11144,N_7547,N_7870);
xnor U11145 (N_11145,N_9275,N_6556);
nor U11146 (N_11146,N_7399,N_8375);
or U11147 (N_11147,N_7289,N_9261);
nor U11148 (N_11148,N_9336,N_8329);
or U11149 (N_11149,N_8497,N_7733);
or U11150 (N_11150,N_8725,N_9149);
nor U11151 (N_11151,N_7654,N_8335);
nand U11152 (N_11152,N_8977,N_6340);
nor U11153 (N_11153,N_6548,N_6460);
nor U11154 (N_11154,N_8671,N_7215);
and U11155 (N_11155,N_9208,N_8100);
nand U11156 (N_11156,N_6584,N_8750);
xor U11157 (N_11157,N_7809,N_9340);
and U11158 (N_11158,N_8289,N_8750);
nor U11159 (N_11159,N_6654,N_7575);
xnor U11160 (N_11160,N_6930,N_9030);
nor U11161 (N_11161,N_8256,N_8070);
nor U11162 (N_11162,N_8296,N_7357);
xnor U11163 (N_11163,N_6637,N_8099);
xor U11164 (N_11164,N_7542,N_8971);
nor U11165 (N_11165,N_7402,N_8878);
nor U11166 (N_11166,N_8847,N_7578);
or U11167 (N_11167,N_7453,N_7103);
or U11168 (N_11168,N_7815,N_9353);
nand U11169 (N_11169,N_8173,N_6306);
nand U11170 (N_11170,N_6587,N_8925);
nand U11171 (N_11171,N_6936,N_8667);
nor U11172 (N_11172,N_6575,N_7611);
nor U11173 (N_11173,N_7388,N_9290);
nand U11174 (N_11174,N_8174,N_7486);
nor U11175 (N_11175,N_6762,N_9087);
and U11176 (N_11176,N_7772,N_7472);
and U11177 (N_11177,N_8486,N_7758);
nor U11178 (N_11178,N_7293,N_7158);
nand U11179 (N_11179,N_7392,N_8854);
or U11180 (N_11180,N_6893,N_6465);
and U11181 (N_11181,N_6355,N_8547);
nand U11182 (N_11182,N_7031,N_8788);
nor U11183 (N_11183,N_7362,N_6479);
and U11184 (N_11184,N_7631,N_7413);
and U11185 (N_11185,N_7689,N_6926);
xnor U11186 (N_11186,N_8750,N_7454);
nor U11187 (N_11187,N_7047,N_7040);
or U11188 (N_11188,N_6324,N_9354);
and U11189 (N_11189,N_8213,N_7506);
xor U11190 (N_11190,N_7762,N_6862);
xor U11191 (N_11191,N_6431,N_7053);
or U11192 (N_11192,N_8282,N_8549);
nand U11193 (N_11193,N_8224,N_8772);
and U11194 (N_11194,N_7079,N_7982);
or U11195 (N_11195,N_8700,N_8692);
xor U11196 (N_11196,N_7224,N_8643);
and U11197 (N_11197,N_6867,N_6263);
nor U11198 (N_11198,N_9148,N_6321);
or U11199 (N_11199,N_7557,N_8888);
nor U11200 (N_11200,N_7211,N_7033);
or U11201 (N_11201,N_8070,N_6962);
nor U11202 (N_11202,N_7491,N_8165);
nor U11203 (N_11203,N_6930,N_8753);
and U11204 (N_11204,N_8591,N_6277);
nand U11205 (N_11205,N_7271,N_7939);
or U11206 (N_11206,N_7137,N_7040);
nor U11207 (N_11207,N_8439,N_6333);
nor U11208 (N_11208,N_6868,N_8668);
nand U11209 (N_11209,N_6974,N_8347);
nor U11210 (N_11210,N_7574,N_8827);
nor U11211 (N_11211,N_9239,N_7039);
and U11212 (N_11212,N_7599,N_6397);
xnor U11213 (N_11213,N_6650,N_6577);
and U11214 (N_11214,N_7902,N_8301);
nor U11215 (N_11215,N_7793,N_8602);
or U11216 (N_11216,N_8797,N_8151);
nand U11217 (N_11217,N_7883,N_7423);
or U11218 (N_11218,N_7470,N_7194);
nor U11219 (N_11219,N_9322,N_8567);
nand U11220 (N_11220,N_8601,N_6791);
and U11221 (N_11221,N_6598,N_7681);
nor U11222 (N_11222,N_9193,N_8990);
nor U11223 (N_11223,N_7053,N_7039);
nor U11224 (N_11224,N_6582,N_6650);
or U11225 (N_11225,N_8343,N_6967);
or U11226 (N_11226,N_9235,N_6589);
and U11227 (N_11227,N_6954,N_8092);
and U11228 (N_11228,N_7724,N_9045);
and U11229 (N_11229,N_7341,N_6712);
and U11230 (N_11230,N_6928,N_6570);
nand U11231 (N_11231,N_8076,N_6499);
nand U11232 (N_11232,N_7956,N_6739);
nand U11233 (N_11233,N_7814,N_9344);
and U11234 (N_11234,N_9008,N_7518);
or U11235 (N_11235,N_8236,N_7266);
xor U11236 (N_11236,N_8505,N_8976);
nor U11237 (N_11237,N_7620,N_6482);
and U11238 (N_11238,N_6933,N_7419);
and U11239 (N_11239,N_7372,N_8352);
nor U11240 (N_11240,N_7659,N_6269);
nand U11241 (N_11241,N_7580,N_7627);
nand U11242 (N_11242,N_7144,N_6635);
nor U11243 (N_11243,N_7179,N_6714);
nand U11244 (N_11244,N_8370,N_8805);
nor U11245 (N_11245,N_8818,N_6427);
nor U11246 (N_11246,N_7813,N_8470);
xor U11247 (N_11247,N_7206,N_6863);
and U11248 (N_11248,N_7483,N_8051);
and U11249 (N_11249,N_6536,N_7425);
nand U11250 (N_11250,N_6262,N_6953);
and U11251 (N_11251,N_8168,N_7352);
nor U11252 (N_11252,N_6298,N_8882);
nor U11253 (N_11253,N_9359,N_6300);
nand U11254 (N_11254,N_6383,N_6929);
nor U11255 (N_11255,N_8097,N_7265);
and U11256 (N_11256,N_7505,N_7233);
or U11257 (N_11257,N_6758,N_7824);
nand U11258 (N_11258,N_7074,N_8077);
xor U11259 (N_11259,N_9091,N_8994);
and U11260 (N_11260,N_6498,N_9222);
and U11261 (N_11261,N_8078,N_7148);
or U11262 (N_11262,N_8738,N_6888);
nand U11263 (N_11263,N_9368,N_8972);
or U11264 (N_11264,N_8762,N_7137);
nand U11265 (N_11265,N_6338,N_8352);
and U11266 (N_11266,N_6353,N_6727);
and U11267 (N_11267,N_7808,N_8792);
nand U11268 (N_11268,N_8669,N_8880);
nand U11269 (N_11269,N_8703,N_6727);
and U11270 (N_11270,N_8845,N_8933);
or U11271 (N_11271,N_8671,N_7803);
nand U11272 (N_11272,N_8544,N_8414);
nor U11273 (N_11273,N_7981,N_7355);
and U11274 (N_11274,N_7492,N_7542);
and U11275 (N_11275,N_7346,N_9197);
nand U11276 (N_11276,N_8654,N_6792);
nor U11277 (N_11277,N_9304,N_8110);
or U11278 (N_11278,N_7923,N_6493);
or U11279 (N_11279,N_8157,N_8026);
nor U11280 (N_11280,N_8980,N_8447);
or U11281 (N_11281,N_7372,N_8919);
nand U11282 (N_11282,N_6827,N_6630);
and U11283 (N_11283,N_6634,N_7348);
nand U11284 (N_11284,N_7179,N_8285);
nand U11285 (N_11285,N_8630,N_8709);
or U11286 (N_11286,N_8518,N_8020);
or U11287 (N_11287,N_7977,N_7826);
nand U11288 (N_11288,N_6815,N_7814);
nor U11289 (N_11289,N_7394,N_8844);
or U11290 (N_11290,N_7774,N_7566);
nor U11291 (N_11291,N_6629,N_8750);
nand U11292 (N_11292,N_6923,N_8002);
and U11293 (N_11293,N_7324,N_8743);
or U11294 (N_11294,N_8369,N_6694);
xnor U11295 (N_11295,N_7318,N_7439);
nand U11296 (N_11296,N_7696,N_7910);
or U11297 (N_11297,N_6339,N_7346);
nor U11298 (N_11298,N_6606,N_8907);
nand U11299 (N_11299,N_8515,N_9042);
and U11300 (N_11300,N_8406,N_8311);
and U11301 (N_11301,N_6294,N_7151);
xnor U11302 (N_11302,N_7063,N_6494);
nand U11303 (N_11303,N_6756,N_7160);
xnor U11304 (N_11304,N_6405,N_8832);
nor U11305 (N_11305,N_7136,N_8866);
nor U11306 (N_11306,N_8263,N_7646);
or U11307 (N_11307,N_9127,N_7175);
nand U11308 (N_11308,N_7240,N_8937);
and U11309 (N_11309,N_9266,N_8475);
and U11310 (N_11310,N_7383,N_6340);
nand U11311 (N_11311,N_8780,N_8002);
nor U11312 (N_11312,N_7150,N_7659);
nor U11313 (N_11313,N_8052,N_6426);
nor U11314 (N_11314,N_8854,N_8514);
or U11315 (N_11315,N_6953,N_8941);
nand U11316 (N_11316,N_6528,N_8404);
xnor U11317 (N_11317,N_7170,N_9180);
nor U11318 (N_11318,N_6424,N_7309);
xor U11319 (N_11319,N_8998,N_7775);
nand U11320 (N_11320,N_7223,N_6744);
nand U11321 (N_11321,N_9181,N_8628);
or U11322 (N_11322,N_7967,N_8448);
or U11323 (N_11323,N_6992,N_7348);
nand U11324 (N_11324,N_6956,N_6758);
xnor U11325 (N_11325,N_6704,N_7232);
and U11326 (N_11326,N_7569,N_7194);
nand U11327 (N_11327,N_7199,N_6959);
and U11328 (N_11328,N_9252,N_7850);
and U11329 (N_11329,N_8546,N_7141);
nor U11330 (N_11330,N_6740,N_6586);
and U11331 (N_11331,N_8500,N_9021);
and U11332 (N_11332,N_7647,N_7378);
and U11333 (N_11333,N_6527,N_8272);
xor U11334 (N_11334,N_7310,N_8312);
or U11335 (N_11335,N_7980,N_8502);
and U11336 (N_11336,N_8565,N_7484);
xor U11337 (N_11337,N_8362,N_8213);
and U11338 (N_11338,N_7650,N_9046);
nand U11339 (N_11339,N_7496,N_9210);
nor U11340 (N_11340,N_6295,N_7401);
nand U11341 (N_11341,N_9359,N_8904);
nand U11342 (N_11342,N_8336,N_7717);
and U11343 (N_11343,N_7581,N_8623);
and U11344 (N_11344,N_8821,N_7727);
nor U11345 (N_11345,N_7088,N_8384);
nand U11346 (N_11346,N_8763,N_7005);
and U11347 (N_11347,N_7289,N_8203);
xnor U11348 (N_11348,N_7688,N_6950);
nand U11349 (N_11349,N_7905,N_6783);
and U11350 (N_11350,N_7768,N_8785);
and U11351 (N_11351,N_7131,N_7121);
nor U11352 (N_11352,N_7475,N_7622);
and U11353 (N_11353,N_8157,N_7565);
nor U11354 (N_11354,N_8176,N_6801);
or U11355 (N_11355,N_8847,N_7580);
nor U11356 (N_11356,N_6549,N_9252);
nor U11357 (N_11357,N_7847,N_8792);
or U11358 (N_11358,N_6329,N_6363);
and U11359 (N_11359,N_6447,N_7537);
nand U11360 (N_11360,N_8674,N_6625);
nand U11361 (N_11361,N_9114,N_7084);
nor U11362 (N_11362,N_7246,N_7652);
nor U11363 (N_11363,N_7486,N_7136);
or U11364 (N_11364,N_6911,N_8004);
or U11365 (N_11365,N_9227,N_6476);
and U11366 (N_11366,N_6806,N_8216);
xnor U11367 (N_11367,N_8692,N_9370);
nor U11368 (N_11368,N_8131,N_7075);
and U11369 (N_11369,N_6685,N_8184);
nor U11370 (N_11370,N_6608,N_8113);
nand U11371 (N_11371,N_7529,N_9283);
and U11372 (N_11372,N_8434,N_9324);
nand U11373 (N_11373,N_6739,N_8660);
and U11374 (N_11374,N_6406,N_7786);
and U11375 (N_11375,N_7166,N_7282);
xnor U11376 (N_11376,N_6968,N_9313);
or U11377 (N_11377,N_7643,N_8458);
xor U11378 (N_11378,N_8571,N_7009);
xnor U11379 (N_11379,N_7499,N_6834);
nor U11380 (N_11380,N_7802,N_7466);
nor U11381 (N_11381,N_7941,N_6595);
nor U11382 (N_11382,N_6637,N_7659);
nand U11383 (N_11383,N_6338,N_6973);
or U11384 (N_11384,N_6483,N_7592);
or U11385 (N_11385,N_6442,N_7448);
and U11386 (N_11386,N_7494,N_8579);
and U11387 (N_11387,N_7145,N_8694);
nor U11388 (N_11388,N_9029,N_6263);
or U11389 (N_11389,N_7105,N_7608);
and U11390 (N_11390,N_8178,N_7151);
nor U11391 (N_11391,N_6709,N_8650);
and U11392 (N_11392,N_8015,N_8831);
and U11393 (N_11393,N_7704,N_8797);
nand U11394 (N_11394,N_8674,N_7763);
nor U11395 (N_11395,N_8971,N_6250);
xor U11396 (N_11396,N_7004,N_9094);
nor U11397 (N_11397,N_8553,N_9166);
or U11398 (N_11398,N_7707,N_6482);
and U11399 (N_11399,N_8999,N_9226);
nor U11400 (N_11400,N_8749,N_7121);
xnor U11401 (N_11401,N_8878,N_7399);
xor U11402 (N_11402,N_7737,N_8093);
or U11403 (N_11403,N_6991,N_6846);
nand U11404 (N_11404,N_7614,N_6367);
and U11405 (N_11405,N_7472,N_8081);
and U11406 (N_11406,N_8758,N_6953);
nand U11407 (N_11407,N_8412,N_6389);
nor U11408 (N_11408,N_8742,N_8177);
nand U11409 (N_11409,N_8324,N_8264);
and U11410 (N_11410,N_7720,N_7239);
nand U11411 (N_11411,N_8708,N_6895);
or U11412 (N_11412,N_7474,N_7581);
xnor U11413 (N_11413,N_7073,N_7114);
nor U11414 (N_11414,N_7898,N_7538);
nor U11415 (N_11415,N_8855,N_6326);
or U11416 (N_11416,N_7022,N_8778);
or U11417 (N_11417,N_9261,N_7511);
xor U11418 (N_11418,N_8967,N_8983);
nand U11419 (N_11419,N_8314,N_7054);
and U11420 (N_11420,N_6903,N_9313);
xor U11421 (N_11421,N_7872,N_9356);
and U11422 (N_11422,N_7213,N_8540);
nor U11423 (N_11423,N_8234,N_6966);
nand U11424 (N_11424,N_7694,N_6351);
nand U11425 (N_11425,N_8014,N_8135);
nor U11426 (N_11426,N_8218,N_6567);
or U11427 (N_11427,N_7511,N_8070);
nor U11428 (N_11428,N_6318,N_8008);
or U11429 (N_11429,N_8242,N_8089);
or U11430 (N_11430,N_7755,N_8032);
or U11431 (N_11431,N_7048,N_6410);
and U11432 (N_11432,N_8567,N_7152);
nand U11433 (N_11433,N_6549,N_6614);
or U11434 (N_11434,N_7765,N_8438);
and U11435 (N_11435,N_7326,N_9130);
or U11436 (N_11436,N_7151,N_7633);
nor U11437 (N_11437,N_7387,N_7290);
xnor U11438 (N_11438,N_7091,N_7613);
nand U11439 (N_11439,N_6861,N_6273);
nor U11440 (N_11440,N_7889,N_9249);
nand U11441 (N_11441,N_6502,N_8646);
nor U11442 (N_11442,N_8251,N_7696);
and U11443 (N_11443,N_7158,N_8995);
xor U11444 (N_11444,N_7033,N_8142);
nor U11445 (N_11445,N_9295,N_7938);
xor U11446 (N_11446,N_6516,N_8110);
nor U11447 (N_11447,N_7705,N_6422);
nand U11448 (N_11448,N_7340,N_6974);
nor U11449 (N_11449,N_7764,N_6442);
nand U11450 (N_11450,N_7459,N_7525);
nor U11451 (N_11451,N_7702,N_8754);
or U11452 (N_11452,N_7478,N_6529);
and U11453 (N_11453,N_6265,N_7069);
or U11454 (N_11454,N_6892,N_7175);
xnor U11455 (N_11455,N_7769,N_7268);
nand U11456 (N_11456,N_8207,N_8770);
nor U11457 (N_11457,N_9096,N_6257);
nand U11458 (N_11458,N_7649,N_8625);
nor U11459 (N_11459,N_9200,N_7842);
and U11460 (N_11460,N_8223,N_7476);
and U11461 (N_11461,N_7042,N_7522);
and U11462 (N_11462,N_6598,N_6514);
nand U11463 (N_11463,N_8175,N_7125);
or U11464 (N_11464,N_8691,N_7723);
and U11465 (N_11465,N_6317,N_9235);
nand U11466 (N_11466,N_8658,N_9185);
or U11467 (N_11467,N_8635,N_8020);
nand U11468 (N_11468,N_8607,N_6649);
and U11469 (N_11469,N_6356,N_6357);
and U11470 (N_11470,N_8644,N_6466);
and U11471 (N_11471,N_8653,N_6812);
nand U11472 (N_11472,N_7891,N_7824);
nor U11473 (N_11473,N_7007,N_9057);
and U11474 (N_11474,N_9054,N_8151);
and U11475 (N_11475,N_6436,N_6731);
and U11476 (N_11476,N_7579,N_9050);
nor U11477 (N_11477,N_7894,N_7553);
nor U11478 (N_11478,N_6806,N_8044);
or U11479 (N_11479,N_8220,N_6385);
xor U11480 (N_11480,N_8616,N_9020);
and U11481 (N_11481,N_8182,N_8356);
and U11482 (N_11482,N_8103,N_8261);
nor U11483 (N_11483,N_7365,N_6921);
nor U11484 (N_11484,N_9029,N_6940);
xor U11485 (N_11485,N_8262,N_7531);
nor U11486 (N_11486,N_9352,N_6442);
nor U11487 (N_11487,N_7319,N_7606);
or U11488 (N_11488,N_8475,N_7784);
nor U11489 (N_11489,N_8354,N_8558);
nand U11490 (N_11490,N_8294,N_6706);
or U11491 (N_11491,N_8950,N_7990);
xor U11492 (N_11492,N_7141,N_8798);
or U11493 (N_11493,N_7399,N_8371);
and U11494 (N_11494,N_8360,N_9214);
nor U11495 (N_11495,N_7972,N_6530);
xnor U11496 (N_11496,N_8676,N_7654);
nor U11497 (N_11497,N_8173,N_8155);
nand U11498 (N_11498,N_8390,N_7648);
nand U11499 (N_11499,N_8845,N_8771);
and U11500 (N_11500,N_7473,N_7163);
nand U11501 (N_11501,N_7734,N_7504);
nand U11502 (N_11502,N_8918,N_6508);
and U11503 (N_11503,N_9096,N_6349);
nor U11504 (N_11504,N_9356,N_6700);
or U11505 (N_11505,N_6960,N_6253);
or U11506 (N_11506,N_8850,N_7832);
and U11507 (N_11507,N_6680,N_6766);
nor U11508 (N_11508,N_8825,N_7465);
or U11509 (N_11509,N_8787,N_6702);
nor U11510 (N_11510,N_7933,N_6823);
and U11511 (N_11511,N_6877,N_7269);
nand U11512 (N_11512,N_7594,N_6879);
nor U11513 (N_11513,N_7492,N_8956);
nand U11514 (N_11514,N_8257,N_9340);
and U11515 (N_11515,N_8445,N_6638);
xor U11516 (N_11516,N_7546,N_8173);
or U11517 (N_11517,N_8329,N_8748);
nand U11518 (N_11518,N_7006,N_6285);
nor U11519 (N_11519,N_7211,N_6907);
and U11520 (N_11520,N_7138,N_7837);
nor U11521 (N_11521,N_7204,N_7208);
or U11522 (N_11522,N_6601,N_6903);
nor U11523 (N_11523,N_9348,N_7897);
nor U11524 (N_11524,N_6603,N_9345);
nor U11525 (N_11525,N_6995,N_8447);
or U11526 (N_11526,N_6748,N_9149);
or U11527 (N_11527,N_6715,N_6659);
or U11528 (N_11528,N_7621,N_7080);
nor U11529 (N_11529,N_7077,N_6800);
nor U11530 (N_11530,N_6991,N_8452);
nor U11531 (N_11531,N_7884,N_8996);
or U11532 (N_11532,N_8070,N_7185);
or U11533 (N_11533,N_7677,N_6310);
nor U11534 (N_11534,N_7185,N_7771);
or U11535 (N_11535,N_9111,N_8936);
nor U11536 (N_11536,N_7408,N_7402);
or U11537 (N_11537,N_6720,N_7001);
and U11538 (N_11538,N_6353,N_7484);
or U11539 (N_11539,N_6926,N_9365);
nor U11540 (N_11540,N_7336,N_8778);
and U11541 (N_11541,N_9080,N_8452);
nand U11542 (N_11542,N_7679,N_8888);
and U11543 (N_11543,N_7140,N_8732);
nor U11544 (N_11544,N_9212,N_9092);
and U11545 (N_11545,N_9047,N_8925);
or U11546 (N_11546,N_8869,N_7793);
nand U11547 (N_11547,N_9280,N_9293);
nor U11548 (N_11548,N_6625,N_8633);
and U11549 (N_11549,N_6623,N_6756);
nor U11550 (N_11550,N_6549,N_7690);
and U11551 (N_11551,N_9269,N_6345);
nor U11552 (N_11552,N_6631,N_8575);
and U11553 (N_11553,N_7784,N_7306);
nand U11554 (N_11554,N_7199,N_8550);
nand U11555 (N_11555,N_7625,N_7370);
xor U11556 (N_11556,N_7922,N_6829);
nor U11557 (N_11557,N_6441,N_6549);
and U11558 (N_11558,N_7337,N_8294);
xnor U11559 (N_11559,N_7508,N_6690);
nand U11560 (N_11560,N_8558,N_8748);
nand U11561 (N_11561,N_7668,N_8394);
or U11562 (N_11562,N_8999,N_8475);
nand U11563 (N_11563,N_7123,N_8820);
nand U11564 (N_11564,N_8127,N_8910);
nand U11565 (N_11565,N_7390,N_7400);
or U11566 (N_11566,N_8994,N_6948);
and U11567 (N_11567,N_8150,N_7009);
nor U11568 (N_11568,N_9293,N_7091);
nor U11569 (N_11569,N_6523,N_7800);
or U11570 (N_11570,N_6785,N_8402);
nor U11571 (N_11571,N_9023,N_6659);
xnor U11572 (N_11572,N_6521,N_7676);
nor U11573 (N_11573,N_6797,N_8299);
nand U11574 (N_11574,N_6446,N_8064);
and U11575 (N_11575,N_7009,N_7735);
nand U11576 (N_11576,N_7444,N_8308);
nand U11577 (N_11577,N_6861,N_8408);
nor U11578 (N_11578,N_7873,N_8148);
or U11579 (N_11579,N_8457,N_7056);
nand U11580 (N_11580,N_7236,N_8194);
or U11581 (N_11581,N_6317,N_8414);
or U11582 (N_11582,N_7122,N_6274);
nor U11583 (N_11583,N_8405,N_7218);
and U11584 (N_11584,N_8573,N_6268);
or U11585 (N_11585,N_6262,N_7791);
xor U11586 (N_11586,N_7142,N_6909);
and U11587 (N_11587,N_7333,N_7099);
or U11588 (N_11588,N_8751,N_8449);
nand U11589 (N_11589,N_8455,N_6402);
nand U11590 (N_11590,N_7072,N_7349);
or U11591 (N_11591,N_6843,N_7269);
and U11592 (N_11592,N_8587,N_7552);
xnor U11593 (N_11593,N_6402,N_7952);
nor U11594 (N_11594,N_8825,N_6454);
nor U11595 (N_11595,N_6791,N_6738);
or U11596 (N_11596,N_9061,N_7883);
nand U11597 (N_11597,N_6712,N_6441);
and U11598 (N_11598,N_8265,N_6489);
nor U11599 (N_11599,N_7448,N_9094);
xor U11600 (N_11600,N_7447,N_8504);
nand U11601 (N_11601,N_8108,N_9208);
nor U11602 (N_11602,N_7864,N_6654);
or U11603 (N_11603,N_6783,N_6470);
xnor U11604 (N_11604,N_6983,N_7756);
nand U11605 (N_11605,N_7836,N_6851);
xnor U11606 (N_11606,N_7526,N_8819);
or U11607 (N_11607,N_7837,N_8428);
nor U11608 (N_11608,N_8777,N_8601);
or U11609 (N_11609,N_7505,N_6511);
and U11610 (N_11610,N_6377,N_8775);
or U11611 (N_11611,N_8243,N_7365);
or U11612 (N_11612,N_6254,N_7072);
and U11613 (N_11613,N_7470,N_8368);
and U11614 (N_11614,N_6795,N_8262);
and U11615 (N_11615,N_6672,N_8882);
and U11616 (N_11616,N_8290,N_6888);
nor U11617 (N_11617,N_7959,N_6961);
and U11618 (N_11618,N_6446,N_8038);
and U11619 (N_11619,N_6967,N_7898);
and U11620 (N_11620,N_7594,N_9020);
nand U11621 (N_11621,N_6292,N_8728);
and U11622 (N_11622,N_8576,N_9024);
and U11623 (N_11623,N_8064,N_9345);
and U11624 (N_11624,N_8197,N_7491);
nand U11625 (N_11625,N_6999,N_6558);
xnor U11626 (N_11626,N_9167,N_6960);
xor U11627 (N_11627,N_7183,N_9310);
or U11628 (N_11628,N_7495,N_7976);
nand U11629 (N_11629,N_8952,N_8115);
or U11630 (N_11630,N_6491,N_8555);
and U11631 (N_11631,N_8221,N_6471);
or U11632 (N_11632,N_7820,N_8055);
nor U11633 (N_11633,N_7570,N_6430);
xor U11634 (N_11634,N_6644,N_7716);
xnor U11635 (N_11635,N_8402,N_8787);
or U11636 (N_11636,N_8344,N_7742);
nand U11637 (N_11637,N_7806,N_7696);
nand U11638 (N_11638,N_8606,N_6503);
nand U11639 (N_11639,N_7620,N_8905);
nor U11640 (N_11640,N_8461,N_9186);
nor U11641 (N_11641,N_7878,N_7670);
or U11642 (N_11642,N_7227,N_7913);
nand U11643 (N_11643,N_8563,N_9023);
nand U11644 (N_11644,N_9275,N_6847);
nand U11645 (N_11645,N_7027,N_6403);
or U11646 (N_11646,N_7027,N_8124);
or U11647 (N_11647,N_8265,N_6903);
or U11648 (N_11648,N_8796,N_6290);
nor U11649 (N_11649,N_6979,N_8912);
nand U11650 (N_11650,N_7016,N_7824);
and U11651 (N_11651,N_8123,N_6456);
nand U11652 (N_11652,N_8557,N_6444);
nand U11653 (N_11653,N_9081,N_7662);
and U11654 (N_11654,N_8747,N_8836);
xor U11655 (N_11655,N_6306,N_6374);
nor U11656 (N_11656,N_7638,N_9321);
nand U11657 (N_11657,N_8759,N_7451);
and U11658 (N_11658,N_8030,N_7272);
and U11659 (N_11659,N_7488,N_7068);
nand U11660 (N_11660,N_8024,N_6383);
nor U11661 (N_11661,N_9057,N_7609);
and U11662 (N_11662,N_8368,N_8852);
nand U11663 (N_11663,N_8393,N_7810);
or U11664 (N_11664,N_6283,N_6923);
nand U11665 (N_11665,N_7847,N_9222);
nand U11666 (N_11666,N_8103,N_6521);
and U11667 (N_11667,N_8690,N_6463);
nor U11668 (N_11668,N_9233,N_7893);
or U11669 (N_11669,N_6446,N_8831);
nor U11670 (N_11670,N_7249,N_7603);
or U11671 (N_11671,N_9335,N_6806);
nand U11672 (N_11672,N_6437,N_6808);
nor U11673 (N_11673,N_6803,N_7867);
nor U11674 (N_11674,N_7080,N_7841);
and U11675 (N_11675,N_6646,N_7309);
and U11676 (N_11676,N_6671,N_8598);
nand U11677 (N_11677,N_8023,N_7067);
nand U11678 (N_11678,N_8601,N_6584);
nor U11679 (N_11679,N_9321,N_7539);
nor U11680 (N_11680,N_8372,N_7053);
nor U11681 (N_11681,N_7503,N_7517);
and U11682 (N_11682,N_6725,N_6458);
or U11683 (N_11683,N_6900,N_8431);
xnor U11684 (N_11684,N_8007,N_7439);
or U11685 (N_11685,N_8846,N_7446);
or U11686 (N_11686,N_8921,N_7865);
nand U11687 (N_11687,N_9257,N_6827);
or U11688 (N_11688,N_6778,N_7604);
nand U11689 (N_11689,N_8613,N_9075);
nand U11690 (N_11690,N_6819,N_9322);
and U11691 (N_11691,N_7528,N_8054);
nor U11692 (N_11692,N_9138,N_6663);
nand U11693 (N_11693,N_6544,N_8493);
nor U11694 (N_11694,N_6371,N_8320);
nand U11695 (N_11695,N_8363,N_6369);
nor U11696 (N_11696,N_6707,N_8408);
nor U11697 (N_11697,N_7589,N_7158);
nor U11698 (N_11698,N_6591,N_6672);
nor U11699 (N_11699,N_8812,N_9207);
and U11700 (N_11700,N_7761,N_8128);
xor U11701 (N_11701,N_7807,N_9355);
and U11702 (N_11702,N_7453,N_8908);
xnor U11703 (N_11703,N_6499,N_7646);
and U11704 (N_11704,N_8601,N_7989);
nor U11705 (N_11705,N_7402,N_9106);
or U11706 (N_11706,N_9248,N_7706);
nand U11707 (N_11707,N_7280,N_6680);
and U11708 (N_11708,N_7468,N_6888);
nand U11709 (N_11709,N_7166,N_6492);
xor U11710 (N_11710,N_8301,N_7377);
nor U11711 (N_11711,N_8956,N_9345);
nand U11712 (N_11712,N_9158,N_6866);
nand U11713 (N_11713,N_9232,N_9086);
and U11714 (N_11714,N_7537,N_6978);
or U11715 (N_11715,N_7665,N_7488);
and U11716 (N_11716,N_8367,N_6625);
nand U11717 (N_11717,N_9020,N_8485);
nor U11718 (N_11718,N_6902,N_7253);
nand U11719 (N_11719,N_8526,N_6471);
or U11720 (N_11720,N_6530,N_6843);
or U11721 (N_11721,N_7795,N_6861);
and U11722 (N_11722,N_9039,N_6477);
nand U11723 (N_11723,N_8901,N_7391);
nand U11724 (N_11724,N_6538,N_6313);
or U11725 (N_11725,N_9223,N_6707);
nor U11726 (N_11726,N_7807,N_6614);
nand U11727 (N_11727,N_7271,N_7237);
or U11728 (N_11728,N_6970,N_7096);
nand U11729 (N_11729,N_7629,N_9222);
nand U11730 (N_11730,N_6827,N_6323);
nor U11731 (N_11731,N_7386,N_8107);
and U11732 (N_11732,N_8712,N_9296);
nor U11733 (N_11733,N_8395,N_8844);
nand U11734 (N_11734,N_7583,N_8774);
or U11735 (N_11735,N_7312,N_7202);
nor U11736 (N_11736,N_8243,N_7723);
nor U11737 (N_11737,N_7805,N_8680);
and U11738 (N_11738,N_9363,N_8971);
and U11739 (N_11739,N_6345,N_9074);
nand U11740 (N_11740,N_8732,N_8413);
nor U11741 (N_11741,N_8569,N_9129);
or U11742 (N_11742,N_9075,N_6564);
or U11743 (N_11743,N_6399,N_8423);
nand U11744 (N_11744,N_7633,N_7557);
nand U11745 (N_11745,N_6789,N_8900);
xnor U11746 (N_11746,N_9233,N_8893);
or U11747 (N_11747,N_7620,N_6788);
nor U11748 (N_11748,N_6476,N_6255);
nor U11749 (N_11749,N_9199,N_7434);
and U11750 (N_11750,N_9089,N_8594);
and U11751 (N_11751,N_8484,N_8438);
nand U11752 (N_11752,N_9217,N_8271);
nand U11753 (N_11753,N_8172,N_8589);
nand U11754 (N_11754,N_6986,N_7955);
xor U11755 (N_11755,N_7338,N_7297);
or U11756 (N_11756,N_9366,N_6504);
or U11757 (N_11757,N_7589,N_6348);
nand U11758 (N_11758,N_7363,N_7860);
nand U11759 (N_11759,N_9283,N_8829);
nand U11760 (N_11760,N_9142,N_7105);
nor U11761 (N_11761,N_6500,N_6523);
nand U11762 (N_11762,N_9282,N_6816);
nor U11763 (N_11763,N_7635,N_7811);
nor U11764 (N_11764,N_6707,N_8412);
or U11765 (N_11765,N_8927,N_6550);
nor U11766 (N_11766,N_7187,N_8871);
nor U11767 (N_11767,N_9045,N_7096);
nor U11768 (N_11768,N_8436,N_6407);
and U11769 (N_11769,N_6879,N_7147);
and U11770 (N_11770,N_7131,N_9064);
or U11771 (N_11771,N_7423,N_7559);
nor U11772 (N_11772,N_8547,N_8960);
nand U11773 (N_11773,N_8487,N_6573);
nand U11774 (N_11774,N_8393,N_6775);
nand U11775 (N_11775,N_7611,N_6768);
nor U11776 (N_11776,N_6853,N_6352);
nor U11777 (N_11777,N_7391,N_6880);
or U11778 (N_11778,N_7373,N_7205);
or U11779 (N_11779,N_7831,N_6563);
and U11780 (N_11780,N_6803,N_7316);
or U11781 (N_11781,N_7219,N_6417);
or U11782 (N_11782,N_8083,N_6579);
nand U11783 (N_11783,N_7073,N_6468);
and U11784 (N_11784,N_8587,N_7965);
xor U11785 (N_11785,N_6707,N_8594);
nand U11786 (N_11786,N_6279,N_8146);
or U11787 (N_11787,N_9156,N_7774);
or U11788 (N_11788,N_7532,N_7765);
nor U11789 (N_11789,N_7480,N_8642);
and U11790 (N_11790,N_6552,N_7809);
xor U11791 (N_11791,N_6799,N_6977);
or U11792 (N_11792,N_7766,N_6811);
or U11793 (N_11793,N_7154,N_7568);
nor U11794 (N_11794,N_7905,N_7333);
xnor U11795 (N_11795,N_8992,N_6815);
nor U11796 (N_11796,N_9262,N_6932);
nor U11797 (N_11797,N_7183,N_9020);
nor U11798 (N_11798,N_7725,N_8068);
and U11799 (N_11799,N_7653,N_7009);
and U11800 (N_11800,N_8949,N_6804);
xor U11801 (N_11801,N_8823,N_9144);
or U11802 (N_11802,N_7132,N_8578);
and U11803 (N_11803,N_9374,N_7121);
or U11804 (N_11804,N_7544,N_8448);
or U11805 (N_11805,N_7783,N_6292);
nand U11806 (N_11806,N_8634,N_9293);
xor U11807 (N_11807,N_7443,N_8868);
or U11808 (N_11808,N_8700,N_6692);
xor U11809 (N_11809,N_6653,N_9017);
xor U11810 (N_11810,N_7575,N_9216);
and U11811 (N_11811,N_8604,N_8943);
and U11812 (N_11812,N_6674,N_7176);
and U11813 (N_11813,N_8998,N_6640);
nor U11814 (N_11814,N_7788,N_6842);
nand U11815 (N_11815,N_8964,N_6527);
or U11816 (N_11816,N_8309,N_9284);
nor U11817 (N_11817,N_7296,N_9003);
or U11818 (N_11818,N_7565,N_7587);
nor U11819 (N_11819,N_9049,N_7173);
or U11820 (N_11820,N_9077,N_7250);
or U11821 (N_11821,N_6612,N_7448);
nor U11822 (N_11822,N_7241,N_8700);
or U11823 (N_11823,N_9260,N_7523);
or U11824 (N_11824,N_7107,N_8256);
and U11825 (N_11825,N_7469,N_6991);
or U11826 (N_11826,N_7458,N_6565);
or U11827 (N_11827,N_7361,N_7556);
and U11828 (N_11828,N_7022,N_8110);
or U11829 (N_11829,N_6789,N_9276);
nor U11830 (N_11830,N_7141,N_8596);
xor U11831 (N_11831,N_6631,N_9117);
nor U11832 (N_11832,N_8367,N_9320);
xor U11833 (N_11833,N_8507,N_7161);
and U11834 (N_11834,N_7186,N_7991);
or U11835 (N_11835,N_7995,N_7231);
nand U11836 (N_11836,N_8275,N_8703);
and U11837 (N_11837,N_7074,N_7788);
nand U11838 (N_11838,N_8529,N_8695);
and U11839 (N_11839,N_6627,N_6593);
xnor U11840 (N_11840,N_8128,N_6928);
nand U11841 (N_11841,N_8979,N_6873);
nor U11842 (N_11842,N_6592,N_7072);
nand U11843 (N_11843,N_6317,N_7148);
nor U11844 (N_11844,N_7098,N_8654);
nor U11845 (N_11845,N_8274,N_8970);
and U11846 (N_11846,N_8107,N_6523);
and U11847 (N_11847,N_7436,N_8574);
or U11848 (N_11848,N_7337,N_7154);
xor U11849 (N_11849,N_8012,N_6282);
xor U11850 (N_11850,N_6858,N_7671);
xor U11851 (N_11851,N_9286,N_6382);
nand U11852 (N_11852,N_8119,N_9080);
and U11853 (N_11853,N_9044,N_8032);
nor U11854 (N_11854,N_8557,N_9326);
nand U11855 (N_11855,N_7038,N_6434);
and U11856 (N_11856,N_7883,N_6304);
and U11857 (N_11857,N_8048,N_8192);
and U11858 (N_11858,N_8451,N_8331);
nor U11859 (N_11859,N_6644,N_8311);
or U11860 (N_11860,N_8403,N_8800);
and U11861 (N_11861,N_8464,N_7186);
nand U11862 (N_11862,N_6860,N_6906);
or U11863 (N_11863,N_8926,N_7966);
and U11864 (N_11864,N_8988,N_7019);
nand U11865 (N_11865,N_7492,N_8426);
or U11866 (N_11866,N_8924,N_9344);
or U11867 (N_11867,N_8565,N_8824);
nand U11868 (N_11868,N_6423,N_9017);
and U11869 (N_11869,N_6839,N_8882);
or U11870 (N_11870,N_8235,N_7929);
xor U11871 (N_11871,N_9008,N_6409);
or U11872 (N_11872,N_8846,N_8512);
and U11873 (N_11873,N_8859,N_6955);
and U11874 (N_11874,N_7471,N_7484);
or U11875 (N_11875,N_9261,N_8534);
nand U11876 (N_11876,N_7210,N_7402);
and U11877 (N_11877,N_7579,N_6520);
or U11878 (N_11878,N_8134,N_6302);
nor U11879 (N_11879,N_8065,N_7280);
nor U11880 (N_11880,N_8592,N_8358);
nand U11881 (N_11881,N_7970,N_7394);
nand U11882 (N_11882,N_6891,N_9121);
xor U11883 (N_11883,N_6534,N_8587);
nand U11884 (N_11884,N_6284,N_8936);
nor U11885 (N_11885,N_7053,N_7858);
and U11886 (N_11886,N_7208,N_7767);
nor U11887 (N_11887,N_7097,N_6304);
or U11888 (N_11888,N_6550,N_7060);
xnor U11889 (N_11889,N_7826,N_9240);
or U11890 (N_11890,N_9188,N_8264);
or U11891 (N_11891,N_7201,N_8101);
or U11892 (N_11892,N_7373,N_6770);
nand U11893 (N_11893,N_8237,N_7064);
nand U11894 (N_11894,N_7066,N_6992);
nand U11895 (N_11895,N_8976,N_9175);
nor U11896 (N_11896,N_7629,N_7634);
nor U11897 (N_11897,N_8946,N_8011);
nand U11898 (N_11898,N_8218,N_9279);
or U11899 (N_11899,N_8781,N_8537);
or U11900 (N_11900,N_8488,N_8248);
and U11901 (N_11901,N_8912,N_7712);
nand U11902 (N_11902,N_7296,N_7947);
or U11903 (N_11903,N_8468,N_7148);
nand U11904 (N_11904,N_7248,N_9303);
nand U11905 (N_11905,N_8914,N_7406);
xor U11906 (N_11906,N_6472,N_8167);
nor U11907 (N_11907,N_7940,N_6645);
nand U11908 (N_11908,N_8801,N_9029);
nand U11909 (N_11909,N_8541,N_9025);
or U11910 (N_11910,N_7575,N_7902);
or U11911 (N_11911,N_7592,N_8294);
nor U11912 (N_11912,N_8554,N_6541);
or U11913 (N_11913,N_9093,N_9023);
nor U11914 (N_11914,N_8787,N_6503);
and U11915 (N_11915,N_8268,N_6310);
nand U11916 (N_11916,N_6945,N_6379);
and U11917 (N_11917,N_8063,N_6726);
xor U11918 (N_11918,N_8906,N_6286);
nor U11919 (N_11919,N_6591,N_8225);
or U11920 (N_11920,N_9321,N_8422);
nor U11921 (N_11921,N_9213,N_7580);
nand U11922 (N_11922,N_6767,N_8962);
or U11923 (N_11923,N_8693,N_6767);
or U11924 (N_11924,N_7300,N_7852);
xnor U11925 (N_11925,N_7494,N_7469);
xnor U11926 (N_11926,N_9315,N_6303);
nor U11927 (N_11927,N_8004,N_7492);
or U11928 (N_11928,N_7858,N_9014);
nand U11929 (N_11929,N_7531,N_8376);
nor U11930 (N_11930,N_6567,N_8238);
and U11931 (N_11931,N_6933,N_8587);
and U11932 (N_11932,N_9079,N_6580);
nand U11933 (N_11933,N_8419,N_7093);
and U11934 (N_11934,N_9272,N_9088);
nor U11935 (N_11935,N_7472,N_7750);
nor U11936 (N_11936,N_7246,N_8028);
and U11937 (N_11937,N_8783,N_8068);
nor U11938 (N_11938,N_8839,N_7061);
nand U11939 (N_11939,N_6312,N_7658);
nor U11940 (N_11940,N_6968,N_8170);
xor U11941 (N_11941,N_7780,N_7034);
nand U11942 (N_11942,N_7555,N_7015);
nand U11943 (N_11943,N_8024,N_7714);
nand U11944 (N_11944,N_9374,N_6432);
and U11945 (N_11945,N_9125,N_8704);
and U11946 (N_11946,N_6315,N_6779);
nand U11947 (N_11947,N_8969,N_9142);
nand U11948 (N_11948,N_7660,N_7330);
nand U11949 (N_11949,N_7570,N_6287);
or U11950 (N_11950,N_6618,N_7554);
xor U11951 (N_11951,N_9040,N_8545);
or U11952 (N_11952,N_6738,N_6608);
nor U11953 (N_11953,N_6462,N_6931);
and U11954 (N_11954,N_9009,N_8053);
nand U11955 (N_11955,N_8629,N_9154);
and U11956 (N_11956,N_8583,N_7171);
nor U11957 (N_11957,N_8810,N_6453);
xor U11958 (N_11958,N_6612,N_8302);
xor U11959 (N_11959,N_8814,N_8415);
nand U11960 (N_11960,N_6688,N_7370);
nand U11961 (N_11961,N_9041,N_9350);
and U11962 (N_11962,N_7183,N_6893);
nand U11963 (N_11963,N_6645,N_7695);
nand U11964 (N_11964,N_7511,N_8527);
or U11965 (N_11965,N_9072,N_9122);
and U11966 (N_11966,N_7206,N_9032);
and U11967 (N_11967,N_8845,N_8225);
or U11968 (N_11968,N_6567,N_7502);
or U11969 (N_11969,N_6390,N_6270);
nor U11970 (N_11970,N_9037,N_8801);
nor U11971 (N_11971,N_7302,N_8936);
or U11972 (N_11972,N_8586,N_9352);
nand U11973 (N_11973,N_7289,N_8426);
nand U11974 (N_11974,N_6420,N_8443);
and U11975 (N_11975,N_6923,N_7083);
nor U11976 (N_11976,N_8932,N_6277);
and U11977 (N_11977,N_7397,N_9140);
nor U11978 (N_11978,N_7695,N_8072);
nor U11979 (N_11979,N_8920,N_9032);
and U11980 (N_11980,N_6342,N_7725);
or U11981 (N_11981,N_9335,N_9350);
nand U11982 (N_11982,N_7837,N_8291);
nor U11983 (N_11983,N_9247,N_7262);
and U11984 (N_11984,N_7852,N_7436);
nor U11985 (N_11985,N_8183,N_6642);
nand U11986 (N_11986,N_7906,N_6419);
and U11987 (N_11987,N_7113,N_7983);
nand U11988 (N_11988,N_9001,N_6447);
and U11989 (N_11989,N_6954,N_7085);
and U11990 (N_11990,N_7791,N_6832);
xor U11991 (N_11991,N_6895,N_7028);
and U11992 (N_11992,N_7722,N_8337);
nand U11993 (N_11993,N_8939,N_8746);
nor U11994 (N_11994,N_8101,N_8592);
and U11995 (N_11995,N_7896,N_7192);
nand U11996 (N_11996,N_6526,N_8151);
and U11997 (N_11997,N_7911,N_8294);
xor U11998 (N_11998,N_8227,N_9162);
nand U11999 (N_11999,N_6369,N_7368);
nor U12000 (N_12000,N_8301,N_8516);
and U12001 (N_12001,N_9150,N_7181);
and U12002 (N_12002,N_6524,N_8044);
nor U12003 (N_12003,N_9017,N_9305);
and U12004 (N_12004,N_8716,N_7019);
and U12005 (N_12005,N_7226,N_8378);
or U12006 (N_12006,N_7150,N_9185);
and U12007 (N_12007,N_9100,N_8816);
or U12008 (N_12008,N_9361,N_7613);
or U12009 (N_12009,N_7574,N_8953);
or U12010 (N_12010,N_8542,N_8678);
and U12011 (N_12011,N_9048,N_7024);
and U12012 (N_12012,N_7001,N_6732);
or U12013 (N_12013,N_7104,N_7238);
nor U12014 (N_12014,N_7547,N_6283);
and U12015 (N_12015,N_8660,N_7848);
nor U12016 (N_12016,N_8520,N_7551);
and U12017 (N_12017,N_8421,N_8095);
or U12018 (N_12018,N_6620,N_7861);
or U12019 (N_12019,N_7532,N_7256);
and U12020 (N_12020,N_7047,N_7573);
nor U12021 (N_12021,N_9026,N_7867);
nor U12022 (N_12022,N_8042,N_9263);
or U12023 (N_12023,N_6308,N_7250);
and U12024 (N_12024,N_6943,N_7624);
and U12025 (N_12025,N_7457,N_8121);
nor U12026 (N_12026,N_7851,N_7410);
xor U12027 (N_12027,N_8506,N_7494);
nor U12028 (N_12028,N_7920,N_8559);
or U12029 (N_12029,N_7368,N_7683);
xor U12030 (N_12030,N_8734,N_8294);
nor U12031 (N_12031,N_6871,N_8521);
and U12032 (N_12032,N_7390,N_8065);
nand U12033 (N_12033,N_6471,N_7804);
and U12034 (N_12034,N_7907,N_7362);
and U12035 (N_12035,N_8702,N_6331);
and U12036 (N_12036,N_7080,N_7984);
or U12037 (N_12037,N_7569,N_7839);
and U12038 (N_12038,N_7501,N_8566);
and U12039 (N_12039,N_8436,N_8191);
nand U12040 (N_12040,N_8439,N_8790);
nor U12041 (N_12041,N_6357,N_8690);
and U12042 (N_12042,N_6435,N_6976);
and U12043 (N_12043,N_9301,N_6387);
nor U12044 (N_12044,N_8050,N_6871);
or U12045 (N_12045,N_9213,N_8384);
nor U12046 (N_12046,N_7078,N_8763);
or U12047 (N_12047,N_7644,N_6748);
nor U12048 (N_12048,N_9007,N_7041);
nand U12049 (N_12049,N_7349,N_8423);
nand U12050 (N_12050,N_6456,N_8766);
nand U12051 (N_12051,N_7063,N_9065);
or U12052 (N_12052,N_7335,N_7657);
nor U12053 (N_12053,N_8846,N_9074);
xnor U12054 (N_12054,N_7499,N_8003);
or U12055 (N_12055,N_6640,N_7117);
and U12056 (N_12056,N_6567,N_7598);
nand U12057 (N_12057,N_6524,N_8912);
and U12058 (N_12058,N_6836,N_7706);
or U12059 (N_12059,N_6595,N_7948);
nand U12060 (N_12060,N_7936,N_6925);
nand U12061 (N_12061,N_7892,N_6864);
nand U12062 (N_12062,N_8999,N_8132);
nor U12063 (N_12063,N_8491,N_7283);
nor U12064 (N_12064,N_7310,N_8195);
nor U12065 (N_12065,N_7051,N_6500);
and U12066 (N_12066,N_8422,N_7397);
and U12067 (N_12067,N_8279,N_8418);
or U12068 (N_12068,N_9340,N_7253);
or U12069 (N_12069,N_6378,N_6514);
or U12070 (N_12070,N_8059,N_8074);
and U12071 (N_12071,N_6316,N_8069);
nand U12072 (N_12072,N_7008,N_9012);
xor U12073 (N_12073,N_6292,N_6838);
nor U12074 (N_12074,N_7158,N_6799);
nor U12075 (N_12075,N_9081,N_7342);
nor U12076 (N_12076,N_9028,N_7457);
nor U12077 (N_12077,N_6574,N_6642);
and U12078 (N_12078,N_7952,N_8698);
nor U12079 (N_12079,N_7043,N_8977);
and U12080 (N_12080,N_8736,N_9008);
and U12081 (N_12081,N_6823,N_6420);
or U12082 (N_12082,N_7886,N_9066);
nor U12083 (N_12083,N_8697,N_8098);
and U12084 (N_12084,N_7119,N_8915);
nor U12085 (N_12085,N_6693,N_7843);
nor U12086 (N_12086,N_8155,N_8010);
nor U12087 (N_12087,N_8535,N_7889);
nand U12088 (N_12088,N_6383,N_8787);
xnor U12089 (N_12089,N_6798,N_8569);
and U12090 (N_12090,N_6942,N_7471);
nand U12091 (N_12091,N_9020,N_9083);
nor U12092 (N_12092,N_9301,N_8640);
nand U12093 (N_12093,N_7842,N_7595);
nand U12094 (N_12094,N_8156,N_7948);
xor U12095 (N_12095,N_9204,N_6913);
and U12096 (N_12096,N_8994,N_9312);
nor U12097 (N_12097,N_6451,N_9251);
and U12098 (N_12098,N_8715,N_8064);
nor U12099 (N_12099,N_7042,N_6379);
and U12100 (N_12100,N_7616,N_8559);
and U12101 (N_12101,N_8101,N_7383);
nor U12102 (N_12102,N_8077,N_8593);
nand U12103 (N_12103,N_8557,N_7655);
nand U12104 (N_12104,N_6931,N_6676);
and U12105 (N_12105,N_6637,N_8199);
or U12106 (N_12106,N_7469,N_6793);
nor U12107 (N_12107,N_8600,N_7527);
nand U12108 (N_12108,N_8171,N_6811);
and U12109 (N_12109,N_7714,N_6995);
and U12110 (N_12110,N_6676,N_8192);
nor U12111 (N_12111,N_9181,N_6406);
xnor U12112 (N_12112,N_7378,N_7078);
nor U12113 (N_12113,N_7676,N_6720);
nor U12114 (N_12114,N_7922,N_7539);
and U12115 (N_12115,N_7671,N_7295);
xnor U12116 (N_12116,N_8815,N_6611);
nor U12117 (N_12117,N_9293,N_7170);
or U12118 (N_12118,N_8235,N_8580);
nor U12119 (N_12119,N_8620,N_8276);
nor U12120 (N_12120,N_7818,N_8290);
xor U12121 (N_12121,N_9208,N_7493);
or U12122 (N_12122,N_8723,N_9067);
and U12123 (N_12123,N_6852,N_9211);
nand U12124 (N_12124,N_6840,N_6960);
and U12125 (N_12125,N_8926,N_6587);
or U12126 (N_12126,N_6880,N_8732);
and U12127 (N_12127,N_6433,N_6666);
and U12128 (N_12128,N_7676,N_8301);
and U12129 (N_12129,N_7229,N_9112);
nor U12130 (N_12130,N_8285,N_7082);
nand U12131 (N_12131,N_7497,N_9178);
or U12132 (N_12132,N_8915,N_6899);
xnor U12133 (N_12133,N_6252,N_6323);
and U12134 (N_12134,N_8435,N_7356);
nand U12135 (N_12135,N_8782,N_7063);
or U12136 (N_12136,N_6345,N_7241);
xor U12137 (N_12137,N_7504,N_8498);
and U12138 (N_12138,N_7643,N_6612);
nand U12139 (N_12139,N_7668,N_7996);
or U12140 (N_12140,N_6697,N_9301);
nand U12141 (N_12141,N_8390,N_6945);
or U12142 (N_12142,N_7502,N_6845);
or U12143 (N_12143,N_8189,N_6566);
nand U12144 (N_12144,N_8711,N_8545);
and U12145 (N_12145,N_8416,N_7159);
xnor U12146 (N_12146,N_7017,N_7512);
or U12147 (N_12147,N_6366,N_7691);
and U12148 (N_12148,N_6659,N_6843);
and U12149 (N_12149,N_6831,N_7742);
nand U12150 (N_12150,N_6612,N_7977);
and U12151 (N_12151,N_8799,N_6568);
and U12152 (N_12152,N_9307,N_8030);
and U12153 (N_12153,N_7895,N_9161);
or U12154 (N_12154,N_8436,N_7580);
nor U12155 (N_12155,N_6581,N_8740);
and U12156 (N_12156,N_9327,N_6778);
or U12157 (N_12157,N_9365,N_8446);
xnor U12158 (N_12158,N_8382,N_7920);
nand U12159 (N_12159,N_6702,N_9195);
nor U12160 (N_12160,N_8109,N_8003);
or U12161 (N_12161,N_7181,N_6808);
nand U12162 (N_12162,N_7410,N_6720);
and U12163 (N_12163,N_7439,N_6335);
and U12164 (N_12164,N_8179,N_8692);
or U12165 (N_12165,N_6345,N_8014);
nor U12166 (N_12166,N_7076,N_7587);
nor U12167 (N_12167,N_8790,N_9318);
nor U12168 (N_12168,N_8425,N_7304);
or U12169 (N_12169,N_7853,N_6553);
nor U12170 (N_12170,N_8358,N_8262);
or U12171 (N_12171,N_7500,N_6302);
nand U12172 (N_12172,N_7155,N_6405);
or U12173 (N_12173,N_7361,N_8579);
nor U12174 (N_12174,N_7715,N_8534);
and U12175 (N_12175,N_9329,N_6865);
nand U12176 (N_12176,N_7579,N_9138);
nor U12177 (N_12177,N_7088,N_6951);
nor U12178 (N_12178,N_7573,N_6388);
xnor U12179 (N_12179,N_6685,N_6710);
or U12180 (N_12180,N_7382,N_7240);
or U12181 (N_12181,N_7941,N_7905);
nor U12182 (N_12182,N_7640,N_7669);
nor U12183 (N_12183,N_6657,N_9095);
or U12184 (N_12184,N_8005,N_7014);
xnor U12185 (N_12185,N_8706,N_7918);
nand U12186 (N_12186,N_7563,N_8097);
or U12187 (N_12187,N_8345,N_6383);
or U12188 (N_12188,N_9211,N_9113);
or U12189 (N_12189,N_7145,N_6554);
nand U12190 (N_12190,N_7910,N_6903);
and U12191 (N_12191,N_6470,N_9170);
nand U12192 (N_12192,N_7880,N_8442);
and U12193 (N_12193,N_8786,N_9125);
nand U12194 (N_12194,N_7708,N_8081);
or U12195 (N_12195,N_8946,N_8260);
or U12196 (N_12196,N_8628,N_7361);
or U12197 (N_12197,N_6422,N_6257);
and U12198 (N_12198,N_8397,N_7350);
or U12199 (N_12199,N_6715,N_6343);
xor U12200 (N_12200,N_8554,N_6254);
nand U12201 (N_12201,N_6914,N_8697);
nor U12202 (N_12202,N_7757,N_6968);
or U12203 (N_12203,N_7996,N_6358);
nand U12204 (N_12204,N_6772,N_9047);
nand U12205 (N_12205,N_6291,N_8312);
nor U12206 (N_12206,N_8630,N_9151);
xnor U12207 (N_12207,N_9106,N_6875);
and U12208 (N_12208,N_6457,N_6258);
or U12209 (N_12209,N_8598,N_7509);
or U12210 (N_12210,N_6881,N_8888);
nor U12211 (N_12211,N_7751,N_8540);
xnor U12212 (N_12212,N_7948,N_7579);
nor U12213 (N_12213,N_9338,N_7716);
nor U12214 (N_12214,N_7617,N_8619);
nor U12215 (N_12215,N_9261,N_7386);
nand U12216 (N_12216,N_8941,N_8480);
nand U12217 (N_12217,N_7451,N_9074);
nand U12218 (N_12218,N_9100,N_6591);
nand U12219 (N_12219,N_7196,N_6571);
or U12220 (N_12220,N_6650,N_6951);
nand U12221 (N_12221,N_7892,N_9351);
or U12222 (N_12222,N_6463,N_7419);
or U12223 (N_12223,N_8560,N_7171);
nand U12224 (N_12224,N_8112,N_8812);
nor U12225 (N_12225,N_8019,N_8434);
and U12226 (N_12226,N_8679,N_8257);
nand U12227 (N_12227,N_7339,N_6345);
and U12228 (N_12228,N_6493,N_8061);
nand U12229 (N_12229,N_9243,N_8184);
nor U12230 (N_12230,N_6954,N_7925);
nor U12231 (N_12231,N_8747,N_8561);
nand U12232 (N_12232,N_7599,N_9113);
and U12233 (N_12233,N_8045,N_7931);
nor U12234 (N_12234,N_8417,N_8967);
nand U12235 (N_12235,N_7036,N_8820);
and U12236 (N_12236,N_7784,N_7436);
nor U12237 (N_12237,N_8117,N_6814);
or U12238 (N_12238,N_8900,N_7603);
nand U12239 (N_12239,N_6610,N_7107);
xor U12240 (N_12240,N_8468,N_6276);
and U12241 (N_12241,N_6295,N_7475);
and U12242 (N_12242,N_7662,N_7245);
or U12243 (N_12243,N_8938,N_7329);
or U12244 (N_12244,N_7423,N_7823);
nor U12245 (N_12245,N_6624,N_9253);
nand U12246 (N_12246,N_9251,N_6745);
or U12247 (N_12247,N_7179,N_7446);
or U12248 (N_12248,N_7702,N_6295);
nand U12249 (N_12249,N_8347,N_8611);
and U12250 (N_12250,N_8703,N_6732);
nand U12251 (N_12251,N_7344,N_6620);
and U12252 (N_12252,N_6653,N_7331);
nand U12253 (N_12253,N_8440,N_9361);
or U12254 (N_12254,N_8459,N_9051);
and U12255 (N_12255,N_8162,N_8214);
or U12256 (N_12256,N_6408,N_8664);
nand U12257 (N_12257,N_6901,N_7822);
or U12258 (N_12258,N_9214,N_9121);
xnor U12259 (N_12259,N_8986,N_7352);
or U12260 (N_12260,N_8078,N_8777);
nor U12261 (N_12261,N_8906,N_6427);
nor U12262 (N_12262,N_8106,N_8566);
nor U12263 (N_12263,N_8942,N_8019);
nand U12264 (N_12264,N_8522,N_8648);
xnor U12265 (N_12265,N_8659,N_8760);
xor U12266 (N_12266,N_8423,N_6371);
or U12267 (N_12267,N_7406,N_8275);
and U12268 (N_12268,N_7359,N_6273);
or U12269 (N_12269,N_7134,N_9001);
nand U12270 (N_12270,N_7612,N_9300);
nand U12271 (N_12271,N_6826,N_7168);
xor U12272 (N_12272,N_6936,N_6980);
nor U12273 (N_12273,N_7184,N_7615);
nand U12274 (N_12274,N_8479,N_8428);
nand U12275 (N_12275,N_7121,N_6450);
nand U12276 (N_12276,N_9111,N_8052);
nor U12277 (N_12277,N_6469,N_7102);
nand U12278 (N_12278,N_9123,N_8976);
or U12279 (N_12279,N_9343,N_8186);
and U12280 (N_12280,N_7558,N_9014);
nor U12281 (N_12281,N_6446,N_6332);
or U12282 (N_12282,N_7361,N_7184);
xor U12283 (N_12283,N_7589,N_6891);
xnor U12284 (N_12284,N_9346,N_8119);
nor U12285 (N_12285,N_9160,N_6747);
or U12286 (N_12286,N_6547,N_8676);
nor U12287 (N_12287,N_8904,N_8651);
nor U12288 (N_12288,N_7475,N_8145);
xor U12289 (N_12289,N_9140,N_8349);
and U12290 (N_12290,N_8482,N_6702);
and U12291 (N_12291,N_7179,N_8121);
or U12292 (N_12292,N_7978,N_9034);
nand U12293 (N_12293,N_9250,N_8297);
nor U12294 (N_12294,N_8292,N_9106);
or U12295 (N_12295,N_7024,N_7362);
and U12296 (N_12296,N_7227,N_6570);
nand U12297 (N_12297,N_6662,N_7673);
nor U12298 (N_12298,N_8799,N_7481);
and U12299 (N_12299,N_6692,N_7517);
nand U12300 (N_12300,N_6568,N_6468);
or U12301 (N_12301,N_7255,N_8193);
nor U12302 (N_12302,N_7551,N_7875);
nand U12303 (N_12303,N_8176,N_7709);
nand U12304 (N_12304,N_7113,N_9000);
nor U12305 (N_12305,N_8285,N_9063);
nor U12306 (N_12306,N_7795,N_6507);
and U12307 (N_12307,N_7023,N_8285);
nand U12308 (N_12308,N_6462,N_7333);
nor U12309 (N_12309,N_9014,N_7205);
xnor U12310 (N_12310,N_7845,N_7790);
xor U12311 (N_12311,N_9315,N_8142);
and U12312 (N_12312,N_7293,N_6530);
nor U12313 (N_12313,N_8107,N_8265);
and U12314 (N_12314,N_6887,N_8814);
nor U12315 (N_12315,N_8477,N_7093);
and U12316 (N_12316,N_8350,N_8585);
and U12317 (N_12317,N_7616,N_8172);
nor U12318 (N_12318,N_7279,N_8940);
or U12319 (N_12319,N_8143,N_7749);
and U12320 (N_12320,N_8225,N_7969);
and U12321 (N_12321,N_8432,N_6288);
nor U12322 (N_12322,N_9171,N_8523);
and U12323 (N_12323,N_8192,N_8480);
xor U12324 (N_12324,N_7898,N_8725);
and U12325 (N_12325,N_6764,N_7857);
nor U12326 (N_12326,N_9342,N_8445);
nor U12327 (N_12327,N_8976,N_7818);
xor U12328 (N_12328,N_7147,N_8908);
or U12329 (N_12329,N_7396,N_7494);
nand U12330 (N_12330,N_8625,N_7910);
xor U12331 (N_12331,N_7877,N_7861);
and U12332 (N_12332,N_8758,N_9344);
and U12333 (N_12333,N_7792,N_8888);
or U12334 (N_12334,N_7874,N_7446);
and U12335 (N_12335,N_7240,N_8609);
nand U12336 (N_12336,N_7447,N_8921);
or U12337 (N_12337,N_6292,N_9122);
xor U12338 (N_12338,N_7059,N_7578);
nor U12339 (N_12339,N_8143,N_7456);
nor U12340 (N_12340,N_7477,N_7449);
or U12341 (N_12341,N_9107,N_8602);
and U12342 (N_12342,N_6258,N_6425);
nand U12343 (N_12343,N_7510,N_7334);
xnor U12344 (N_12344,N_7655,N_8839);
and U12345 (N_12345,N_7016,N_8315);
nor U12346 (N_12346,N_9144,N_9163);
nand U12347 (N_12347,N_8617,N_8314);
nor U12348 (N_12348,N_8255,N_8587);
and U12349 (N_12349,N_6708,N_6377);
nand U12350 (N_12350,N_8155,N_6482);
xor U12351 (N_12351,N_8426,N_8260);
nand U12352 (N_12352,N_7964,N_6477);
xor U12353 (N_12353,N_8961,N_6462);
nor U12354 (N_12354,N_8160,N_8859);
nor U12355 (N_12355,N_6901,N_7508);
nand U12356 (N_12356,N_6457,N_6646);
or U12357 (N_12357,N_9207,N_7074);
and U12358 (N_12358,N_6546,N_7028);
and U12359 (N_12359,N_9178,N_6639);
nor U12360 (N_12360,N_8935,N_7462);
nand U12361 (N_12361,N_6890,N_6710);
or U12362 (N_12362,N_8183,N_8144);
or U12363 (N_12363,N_7154,N_6486);
or U12364 (N_12364,N_7028,N_6937);
nand U12365 (N_12365,N_7885,N_7464);
or U12366 (N_12366,N_7976,N_7818);
xnor U12367 (N_12367,N_8144,N_6610);
or U12368 (N_12368,N_8872,N_7910);
nand U12369 (N_12369,N_6617,N_9245);
and U12370 (N_12370,N_7592,N_7061);
nand U12371 (N_12371,N_9200,N_8409);
or U12372 (N_12372,N_7429,N_8891);
or U12373 (N_12373,N_6998,N_7744);
xor U12374 (N_12374,N_8390,N_8558);
or U12375 (N_12375,N_6487,N_7255);
nand U12376 (N_12376,N_8916,N_6388);
nor U12377 (N_12377,N_6738,N_6730);
nand U12378 (N_12378,N_9028,N_6590);
nand U12379 (N_12379,N_9374,N_8604);
and U12380 (N_12380,N_8647,N_9180);
and U12381 (N_12381,N_8208,N_8605);
and U12382 (N_12382,N_6345,N_7807);
or U12383 (N_12383,N_6753,N_9007);
and U12384 (N_12384,N_8716,N_9217);
or U12385 (N_12385,N_7168,N_9347);
nor U12386 (N_12386,N_7204,N_6754);
xor U12387 (N_12387,N_8128,N_7543);
xor U12388 (N_12388,N_9215,N_7732);
nor U12389 (N_12389,N_8624,N_8461);
or U12390 (N_12390,N_9318,N_8902);
nor U12391 (N_12391,N_7562,N_6514);
xnor U12392 (N_12392,N_9050,N_7314);
or U12393 (N_12393,N_7742,N_8314);
nor U12394 (N_12394,N_6441,N_7769);
nand U12395 (N_12395,N_9329,N_8104);
nand U12396 (N_12396,N_7428,N_8209);
or U12397 (N_12397,N_6620,N_9154);
nor U12398 (N_12398,N_7132,N_6917);
nand U12399 (N_12399,N_9189,N_6630);
nor U12400 (N_12400,N_9279,N_8551);
or U12401 (N_12401,N_8572,N_7420);
nand U12402 (N_12402,N_6876,N_7595);
or U12403 (N_12403,N_7859,N_9095);
and U12404 (N_12404,N_8373,N_6851);
and U12405 (N_12405,N_8281,N_6848);
and U12406 (N_12406,N_6669,N_8596);
nand U12407 (N_12407,N_8445,N_8682);
nand U12408 (N_12408,N_9206,N_8165);
nand U12409 (N_12409,N_7934,N_7102);
nand U12410 (N_12410,N_9291,N_8761);
xor U12411 (N_12411,N_9124,N_9110);
and U12412 (N_12412,N_6663,N_8442);
nor U12413 (N_12413,N_7369,N_7451);
nand U12414 (N_12414,N_7350,N_6412);
xnor U12415 (N_12415,N_8683,N_6405);
nand U12416 (N_12416,N_6938,N_7094);
nand U12417 (N_12417,N_7766,N_8818);
nor U12418 (N_12418,N_9110,N_6602);
nand U12419 (N_12419,N_6565,N_9019);
or U12420 (N_12420,N_8065,N_9218);
and U12421 (N_12421,N_7502,N_8288);
or U12422 (N_12422,N_8461,N_6662);
xnor U12423 (N_12423,N_6265,N_9032);
and U12424 (N_12424,N_9151,N_7679);
and U12425 (N_12425,N_6383,N_8600);
or U12426 (N_12426,N_9046,N_8788);
or U12427 (N_12427,N_6673,N_6335);
and U12428 (N_12428,N_6919,N_6293);
nor U12429 (N_12429,N_7862,N_8154);
nand U12430 (N_12430,N_7287,N_9188);
and U12431 (N_12431,N_8671,N_9019);
or U12432 (N_12432,N_6265,N_9052);
xor U12433 (N_12433,N_7920,N_6842);
or U12434 (N_12434,N_8436,N_7111);
xor U12435 (N_12435,N_8068,N_7976);
nand U12436 (N_12436,N_8010,N_8364);
or U12437 (N_12437,N_7583,N_6535);
xnor U12438 (N_12438,N_6612,N_7695);
nor U12439 (N_12439,N_8157,N_7394);
or U12440 (N_12440,N_8547,N_8347);
xor U12441 (N_12441,N_7295,N_7098);
nand U12442 (N_12442,N_6866,N_8772);
nand U12443 (N_12443,N_8547,N_8021);
nand U12444 (N_12444,N_6397,N_6755);
nand U12445 (N_12445,N_9168,N_8683);
nand U12446 (N_12446,N_8566,N_9371);
or U12447 (N_12447,N_8393,N_7097);
and U12448 (N_12448,N_7131,N_7371);
and U12449 (N_12449,N_8536,N_6254);
nand U12450 (N_12450,N_8572,N_8415);
and U12451 (N_12451,N_7577,N_8475);
xor U12452 (N_12452,N_6253,N_7339);
or U12453 (N_12453,N_7813,N_9050);
nor U12454 (N_12454,N_8451,N_7037);
or U12455 (N_12455,N_7474,N_8005);
or U12456 (N_12456,N_7562,N_6981);
and U12457 (N_12457,N_7466,N_6960);
nand U12458 (N_12458,N_6349,N_6727);
or U12459 (N_12459,N_6421,N_8086);
or U12460 (N_12460,N_9235,N_6620);
nand U12461 (N_12461,N_8712,N_6769);
or U12462 (N_12462,N_9368,N_9331);
or U12463 (N_12463,N_8936,N_9178);
xnor U12464 (N_12464,N_9118,N_6949);
nand U12465 (N_12465,N_7109,N_8007);
and U12466 (N_12466,N_8970,N_6258);
or U12467 (N_12467,N_7989,N_7813);
or U12468 (N_12468,N_9363,N_7913);
nand U12469 (N_12469,N_8566,N_7349);
or U12470 (N_12470,N_7587,N_8008);
or U12471 (N_12471,N_8232,N_6831);
or U12472 (N_12472,N_6740,N_7765);
nand U12473 (N_12473,N_7581,N_7034);
and U12474 (N_12474,N_6708,N_7333);
and U12475 (N_12475,N_7457,N_7447);
nand U12476 (N_12476,N_6579,N_6499);
and U12477 (N_12477,N_8866,N_8264);
nand U12478 (N_12478,N_7144,N_6343);
xnor U12479 (N_12479,N_6403,N_6286);
nand U12480 (N_12480,N_8188,N_9360);
or U12481 (N_12481,N_9132,N_6745);
or U12482 (N_12482,N_8598,N_7391);
nand U12483 (N_12483,N_7562,N_8425);
nor U12484 (N_12484,N_8182,N_7119);
nand U12485 (N_12485,N_9155,N_8433);
nand U12486 (N_12486,N_8135,N_8671);
nor U12487 (N_12487,N_8320,N_8877);
nand U12488 (N_12488,N_7618,N_9230);
and U12489 (N_12489,N_7153,N_8767);
nor U12490 (N_12490,N_7863,N_8384);
and U12491 (N_12491,N_9011,N_6734);
nor U12492 (N_12492,N_7615,N_7972);
nand U12493 (N_12493,N_8254,N_8798);
nor U12494 (N_12494,N_6512,N_9188);
and U12495 (N_12495,N_8444,N_6872);
nor U12496 (N_12496,N_7615,N_6686);
nor U12497 (N_12497,N_7815,N_6506);
xor U12498 (N_12498,N_7442,N_7619);
nand U12499 (N_12499,N_6474,N_6460);
and U12500 (N_12500,N_12040,N_11739);
or U12501 (N_12501,N_11784,N_9815);
xnor U12502 (N_12502,N_12111,N_11992);
nand U12503 (N_12503,N_11896,N_12407);
xor U12504 (N_12504,N_9872,N_10242);
nand U12505 (N_12505,N_9909,N_12047);
nor U12506 (N_12506,N_10555,N_12302);
nand U12507 (N_12507,N_11927,N_11728);
and U12508 (N_12508,N_10238,N_10320);
xnor U12509 (N_12509,N_11101,N_11106);
and U12510 (N_12510,N_9977,N_9984);
or U12511 (N_12511,N_12206,N_9622);
nor U12512 (N_12512,N_10314,N_10450);
and U12513 (N_12513,N_10495,N_9707);
xnor U12514 (N_12514,N_12171,N_10660);
and U12515 (N_12515,N_10090,N_9942);
and U12516 (N_12516,N_10097,N_9514);
xnor U12517 (N_12517,N_9727,N_11579);
and U12518 (N_12518,N_9943,N_9923);
nand U12519 (N_12519,N_9965,N_11866);
xnor U12520 (N_12520,N_12080,N_9513);
nand U12521 (N_12521,N_12448,N_10725);
nor U12522 (N_12522,N_11275,N_12383);
xnor U12523 (N_12523,N_9986,N_10052);
or U12524 (N_12524,N_12330,N_11303);
nor U12525 (N_12525,N_10489,N_11124);
or U12526 (N_12526,N_10895,N_12212);
nand U12527 (N_12527,N_11792,N_9430);
nand U12528 (N_12528,N_12428,N_9686);
or U12529 (N_12529,N_10943,N_11100);
and U12530 (N_12530,N_11207,N_12199);
or U12531 (N_12531,N_9667,N_9612);
nand U12532 (N_12532,N_9523,N_10830);
or U12533 (N_12533,N_10205,N_11108);
or U12534 (N_12534,N_11640,N_12332);
nor U12535 (N_12535,N_12429,N_11691);
nor U12536 (N_12536,N_11919,N_11214);
and U12537 (N_12537,N_10877,N_12161);
nor U12538 (N_12538,N_12373,N_11753);
nor U12539 (N_12539,N_10956,N_9831);
nor U12540 (N_12540,N_12197,N_9556);
and U12541 (N_12541,N_10594,N_11611);
or U12542 (N_12542,N_10043,N_11248);
nor U12543 (N_12543,N_10283,N_9614);
nand U12544 (N_12544,N_11372,N_10973);
nor U12545 (N_12545,N_9440,N_11203);
nor U12546 (N_12546,N_12078,N_11007);
nor U12547 (N_12547,N_9822,N_9429);
nand U12548 (N_12548,N_11823,N_11926);
xnor U12549 (N_12549,N_11018,N_9841);
nand U12550 (N_12550,N_9453,N_9959);
nand U12551 (N_12551,N_11838,N_11221);
or U12552 (N_12552,N_12472,N_9726);
nand U12553 (N_12553,N_9740,N_10735);
nand U12554 (N_12554,N_11238,N_10509);
xor U12555 (N_12555,N_10023,N_9963);
nor U12556 (N_12556,N_11340,N_10381);
nand U12557 (N_12557,N_10246,N_12473);
nand U12558 (N_12558,N_10619,N_12345);
or U12559 (N_12559,N_9828,N_12412);
or U12560 (N_12560,N_9807,N_10425);
nand U12561 (N_12561,N_10353,N_10608);
nor U12562 (N_12562,N_9901,N_10034);
or U12563 (N_12563,N_10835,N_11605);
nand U12564 (N_12564,N_11021,N_10754);
nor U12565 (N_12565,N_10170,N_10856);
or U12566 (N_12566,N_10512,N_12280);
and U12567 (N_12567,N_10247,N_9471);
and U12568 (N_12568,N_11066,N_12229);
and U12569 (N_12569,N_10666,N_10855);
or U12570 (N_12570,N_10572,N_12027);
or U12571 (N_12571,N_10096,N_10999);
or U12572 (N_12572,N_10433,N_10601);
nor U12573 (N_12573,N_9554,N_9652);
nor U12574 (N_12574,N_11457,N_10140);
nor U12575 (N_12575,N_11377,N_11192);
nor U12576 (N_12576,N_10481,N_11464);
nand U12577 (N_12577,N_10109,N_10265);
nor U12578 (N_12578,N_12160,N_11322);
or U12579 (N_12579,N_12118,N_11319);
or U12580 (N_12580,N_10794,N_9520);
and U12581 (N_12581,N_12209,N_9913);
nand U12582 (N_12582,N_10547,N_10234);
and U12583 (N_12583,N_12462,N_11608);
or U12584 (N_12584,N_12261,N_10713);
nor U12585 (N_12585,N_11439,N_9927);
nor U12586 (N_12586,N_10573,N_12085);
nor U12587 (N_12587,N_9477,N_11585);
or U12588 (N_12588,N_10867,N_12252);
and U12589 (N_12589,N_10865,N_12180);
xnor U12590 (N_12590,N_12321,N_10387);
and U12591 (N_12591,N_10690,N_11006);
and U12592 (N_12592,N_9888,N_11068);
or U12593 (N_12593,N_11646,N_10966);
and U12594 (N_12594,N_10689,N_11704);
or U12595 (N_12595,N_11092,N_11750);
nand U12596 (N_12596,N_10310,N_9900);
nor U12597 (N_12597,N_9592,N_11892);
or U12598 (N_12598,N_11342,N_10062);
and U12599 (N_12599,N_11407,N_11001);
nor U12600 (N_12600,N_9469,N_10422);
nand U12601 (N_12601,N_11088,N_9846);
and U12602 (N_12602,N_10336,N_11346);
nor U12603 (N_12603,N_9590,N_10712);
or U12604 (N_12604,N_12431,N_11655);
nand U12605 (N_12605,N_11876,N_10961);
and U12606 (N_12606,N_12360,N_10834);
nand U12607 (N_12607,N_11420,N_11686);
and U12608 (N_12608,N_11759,N_10508);
nor U12609 (N_12609,N_11980,N_12344);
or U12610 (N_12610,N_10896,N_10361);
nor U12611 (N_12611,N_10030,N_12307);
and U12612 (N_12612,N_9725,N_11048);
and U12613 (N_12613,N_12036,N_10717);
and U12614 (N_12614,N_10637,N_10860);
or U12615 (N_12615,N_9674,N_9987);
nand U12616 (N_12616,N_11201,N_9663);
or U12617 (N_12617,N_10319,N_12250);
nor U12618 (N_12618,N_10253,N_11827);
nand U12619 (N_12619,N_10622,N_11010);
or U12620 (N_12620,N_9658,N_12175);
and U12621 (N_12621,N_10367,N_11261);
or U12622 (N_12622,N_11644,N_10846);
or U12623 (N_12623,N_12375,N_10876);
and U12624 (N_12624,N_11610,N_9789);
or U12625 (N_12625,N_10154,N_10544);
nor U12626 (N_12626,N_11394,N_11515);
or U12627 (N_12627,N_11316,N_12087);
nand U12628 (N_12628,N_10498,N_12238);
and U12629 (N_12629,N_12468,N_11071);
or U12630 (N_12630,N_12104,N_9683);
nand U12631 (N_12631,N_10753,N_10581);
and U12632 (N_12632,N_11237,N_10816);
nand U12633 (N_12633,N_10068,N_12168);
nor U12634 (N_12634,N_12222,N_12202);
or U12635 (N_12635,N_10955,N_10702);
and U12636 (N_12636,N_9576,N_12492);
nor U12637 (N_12637,N_9768,N_11878);
xnor U12638 (N_12638,N_10871,N_10143);
or U12639 (N_12639,N_12133,N_12149);
nor U12640 (N_12640,N_10173,N_9529);
and U12641 (N_12641,N_12268,N_12443);
nand U12642 (N_12642,N_11036,N_11914);
nor U12643 (N_12643,N_10949,N_9524);
xnor U12644 (N_12644,N_9617,N_11017);
nand U12645 (N_12645,N_10344,N_11234);
nor U12646 (N_12646,N_9878,N_10954);
and U12647 (N_12647,N_11280,N_9917);
xor U12648 (N_12648,N_11788,N_9424);
or U12649 (N_12649,N_9684,N_9494);
nand U12650 (N_12650,N_11090,N_11259);
nor U12651 (N_12651,N_11198,N_9618);
xnor U12652 (N_12652,N_11793,N_9468);
and U12653 (N_12653,N_10370,N_10972);
xor U12654 (N_12654,N_11713,N_11961);
xor U12655 (N_12655,N_10970,N_10879);
and U12656 (N_12656,N_9729,N_12076);
xnor U12657 (N_12657,N_11391,N_12060);
nand U12658 (N_12658,N_11330,N_11755);
and U12659 (N_12659,N_11039,N_10156);
or U12660 (N_12660,N_11808,N_11559);
nand U12661 (N_12661,N_9458,N_11767);
or U12662 (N_12662,N_12233,N_12123);
or U12663 (N_12663,N_9907,N_10921);
or U12664 (N_12664,N_12493,N_11697);
nand U12665 (N_12665,N_9991,N_11421);
nor U12666 (N_12666,N_11652,N_10423);
and U12667 (N_12667,N_10583,N_10067);
or U12668 (N_12668,N_9474,N_12285);
nand U12669 (N_12669,N_11796,N_11895);
nor U12670 (N_12670,N_9669,N_10014);
and U12671 (N_12671,N_10774,N_10560);
and U12672 (N_12672,N_12018,N_11925);
xnor U12673 (N_12673,N_11651,N_10372);
nor U12674 (N_12674,N_11267,N_11032);
or U12675 (N_12675,N_9832,N_10672);
nand U12676 (N_12676,N_12068,N_11161);
and U12677 (N_12677,N_10908,N_11399);
nand U12678 (N_12678,N_12159,N_10112);
nor U12679 (N_12679,N_10912,N_11177);
xnor U12680 (N_12680,N_11413,N_11845);
or U12681 (N_12681,N_11260,N_10628);
and U12682 (N_12682,N_9647,N_12289);
and U12683 (N_12683,N_9712,N_10805);
nor U12684 (N_12684,N_11787,N_11683);
and U12685 (N_12685,N_11474,N_11974);
xnor U12686 (N_12686,N_10727,N_11091);
nand U12687 (N_12687,N_11831,N_10463);
nor U12688 (N_12688,N_11328,N_9480);
or U12689 (N_12689,N_10127,N_10792);
and U12690 (N_12690,N_12293,N_12427);
nor U12691 (N_12691,N_9574,N_11999);
or U12692 (N_12692,N_12183,N_10849);
xnor U12693 (N_12693,N_9542,N_12478);
or U12694 (N_12694,N_10298,N_10942);
or U12695 (N_12695,N_10959,N_12287);
and U12696 (N_12696,N_10301,N_10119);
xor U12697 (N_12697,N_9487,N_10251);
nor U12698 (N_12698,N_10001,N_10529);
nor U12699 (N_12699,N_9998,N_10315);
nand U12700 (N_12700,N_9535,N_10190);
nand U12701 (N_12701,N_10649,N_10379);
nor U12702 (N_12702,N_11045,N_10979);
nor U12703 (N_12703,N_11951,N_9565);
or U12704 (N_12704,N_9718,N_11848);
nand U12705 (N_12705,N_10145,N_9947);
or U12706 (N_12706,N_9478,N_10850);
nand U12707 (N_12707,N_11726,N_9566);
nor U12708 (N_12708,N_10124,N_12273);
nand U12709 (N_12709,N_10277,N_12158);
and U12710 (N_12710,N_10047,N_9865);
xor U12711 (N_12711,N_9395,N_11065);
nor U12712 (N_12712,N_9448,N_10492);
nor U12713 (N_12713,N_11386,N_9746);
nand U12714 (N_12714,N_12094,N_9941);
nor U12715 (N_12715,N_10210,N_10275);
and U12716 (N_12716,N_10428,N_10008);
nor U12717 (N_12717,N_10497,N_10782);
nor U12718 (N_12718,N_11077,N_9870);
nor U12719 (N_12719,N_10678,N_9690);
nor U12720 (N_12720,N_10821,N_12463);
nor U12721 (N_12721,N_10789,N_12354);
nor U12722 (N_12722,N_11444,N_10720);
and U12723 (N_12723,N_9423,N_11219);
xor U12724 (N_12724,N_10862,N_11757);
or U12725 (N_12725,N_11424,N_12414);
and U12726 (N_12726,N_11055,N_10829);
nand U12727 (N_12727,N_11633,N_10159);
or U12728 (N_12728,N_10233,N_11995);
xnor U12729 (N_12729,N_9755,N_12426);
nand U12730 (N_12730,N_9799,N_11254);
xnor U12731 (N_12731,N_10187,N_10206);
xnor U12732 (N_12732,N_10412,N_12003);
xnor U12733 (N_12733,N_11748,N_9685);
and U12734 (N_12734,N_10245,N_10793);
nor U12735 (N_12735,N_11469,N_9412);
and U12736 (N_12736,N_9517,N_10122);
nor U12737 (N_12737,N_11473,N_10339);
nor U12738 (N_12738,N_9562,N_11013);
and U12739 (N_12739,N_11292,N_10469);
nand U12740 (N_12740,N_10114,N_10312);
nand U12741 (N_12741,N_10944,N_9653);
nor U12742 (N_12742,N_12294,N_12479);
or U12743 (N_12743,N_11978,N_11884);
nand U12744 (N_12744,N_10812,N_9857);
and U12745 (N_12745,N_12061,N_10080);
nand U12746 (N_12746,N_12208,N_10410);
or U12747 (N_12747,N_11472,N_11864);
nand U12748 (N_12748,N_10032,N_11819);
nand U12749 (N_12749,N_10129,N_10536);
nand U12750 (N_12750,N_9665,N_9797);
and U12751 (N_12751,N_11707,N_10021);
nand U12752 (N_12752,N_11975,N_11301);
and U12753 (N_12753,N_9629,N_10487);
nor U12754 (N_12754,N_10737,N_9489);
nor U12755 (N_12755,N_9559,N_11037);
nand U12756 (N_12756,N_10332,N_9500);
and U12757 (N_12757,N_12298,N_12030);
or U12758 (N_12758,N_10137,N_10564);
xor U12759 (N_12759,N_10770,N_11751);
and U12760 (N_12760,N_10341,N_10903);
xor U12761 (N_12761,N_10906,N_11660);
and U12762 (N_12762,N_11150,N_9525);
nand U12763 (N_12763,N_10069,N_9946);
and U12764 (N_12764,N_11890,N_10178);
or U12765 (N_12765,N_10546,N_11132);
nand U12766 (N_12766,N_9454,N_11988);
nor U12767 (N_12767,N_10455,N_11857);
nor U12768 (N_12768,N_12449,N_10393);
nor U12769 (N_12769,N_10389,N_9864);
or U12770 (N_12770,N_12075,N_10559);
and U12771 (N_12771,N_12331,N_12422);
nand U12772 (N_12772,N_12482,N_10212);
and U12773 (N_12773,N_12164,N_9437);
and U12774 (N_12774,N_10201,N_10741);
nand U12775 (N_12775,N_12147,N_10653);
and U12776 (N_12776,N_11053,N_10132);
and U12777 (N_12777,N_12048,N_10086);
nand U12778 (N_12778,N_11481,N_12169);
or U12779 (N_12779,N_12359,N_11350);
and U12780 (N_12780,N_10624,N_10604);
or U12781 (N_12781,N_12059,N_12275);
nor U12782 (N_12782,N_10172,N_12366);
nor U12783 (N_12783,N_11654,N_9638);
nor U12784 (N_12784,N_12353,N_10324);
nor U12785 (N_12785,N_9461,N_10181);
nor U12786 (N_12786,N_11012,N_11471);
nor U12787 (N_12787,N_12000,N_9975);
xor U12788 (N_12788,N_11909,N_11142);
and U12789 (N_12789,N_10142,N_12166);
xor U12790 (N_12790,N_10945,N_12234);
and U12791 (N_12791,N_12107,N_11073);
and U12792 (N_12792,N_10452,N_11458);
nor U12793 (N_12793,N_9497,N_10703);
and U12794 (N_12794,N_11225,N_9522);
or U12795 (N_12795,N_12262,N_10071);
or U12796 (N_12796,N_10892,N_10457);
nand U12797 (N_12797,N_10505,N_10823);
nand U12798 (N_12798,N_11211,N_10971);
or U12799 (N_12799,N_11240,N_9550);
nor U12800 (N_12800,N_12467,N_10471);
or U12801 (N_12801,N_9935,N_12278);
nor U12802 (N_12802,N_10485,N_11057);
and U12803 (N_12803,N_10764,N_11173);
nand U12804 (N_12804,N_9866,N_11868);
xor U12805 (N_12805,N_9415,N_11443);
or U12806 (N_12806,N_10082,N_11917);
nand U12807 (N_12807,N_12079,N_9895);
or U12808 (N_12808,N_9464,N_11673);
or U12809 (N_12809,N_11682,N_9743);
nand U12810 (N_12810,N_11501,N_10115);
nand U12811 (N_12811,N_9957,N_10779);
and U12812 (N_12812,N_11930,N_10281);
or U12813 (N_12813,N_11533,N_9716);
nor U12814 (N_12814,N_11530,N_9751);
nor U12815 (N_12815,N_10960,N_10607);
nand U12816 (N_12816,N_11736,N_11803);
nand U12817 (N_12817,N_9662,N_9386);
and U12818 (N_12818,N_9887,N_12128);
xnor U12819 (N_12819,N_11146,N_9421);
nand U12820 (N_12820,N_10117,N_10270);
nand U12821 (N_12821,N_10872,N_10183);
nor U12822 (N_12822,N_10092,N_9394);
or U12823 (N_12823,N_9431,N_10406);
xor U12824 (N_12824,N_9375,N_12257);
and U12825 (N_12825,N_10517,N_12113);
nand U12826 (N_12826,N_11217,N_11777);
or U12827 (N_12827,N_9995,N_10813);
nor U12828 (N_12828,N_12384,N_11675);
nor U12829 (N_12829,N_11041,N_10897);
xnor U12830 (N_12830,N_10342,N_10507);
or U12831 (N_12831,N_12464,N_10659);
or U12832 (N_12832,N_12045,N_11321);
nand U12833 (N_12833,N_10591,N_11983);
and U12834 (N_12834,N_9905,N_9533);
nor U12835 (N_12835,N_11005,N_11390);
nand U12836 (N_12836,N_12135,N_11327);
nand U12837 (N_12837,N_10985,N_11381);
and U12838 (N_12838,N_10261,N_11944);
and U12839 (N_12839,N_9808,N_10063);
or U12840 (N_12840,N_9442,N_10070);
nor U12841 (N_12841,N_10910,N_10576);
nand U12842 (N_12842,N_11060,N_11255);
and U12843 (N_12843,N_11523,N_9892);
nand U12844 (N_12844,N_9447,N_11718);
nand U12845 (N_12845,N_10099,N_12115);
nor U12846 (N_12846,N_12483,N_11023);
or U12847 (N_12847,N_10435,N_9697);
nor U12848 (N_12848,N_11809,N_9633);
nand U12849 (N_12849,N_11946,N_11294);
xnor U12850 (N_12850,N_11875,N_11854);
nor U12851 (N_12851,N_11535,N_11009);
nor U12852 (N_12852,N_11426,N_12455);
or U12853 (N_12853,N_9476,N_9491);
and U12854 (N_12854,N_10352,N_9893);
or U12855 (N_12855,N_11544,N_12329);
and U12856 (N_12856,N_11806,N_12416);
nand U12857 (N_12857,N_11898,N_10236);
and U12858 (N_12858,N_9657,N_12019);
nand U12859 (N_12859,N_9731,N_10923);
nand U12860 (N_12860,N_10185,N_9704);
xnor U12861 (N_12861,N_9644,N_11766);
and U12862 (N_12862,N_10053,N_10963);
xnor U12863 (N_12863,N_12144,N_9376);
nor U12864 (N_12864,N_9451,N_11133);
or U12865 (N_12865,N_10502,N_11923);
or U12866 (N_12866,N_11649,N_12447);
and U12867 (N_12867,N_9671,N_12401);
nand U12868 (N_12868,N_12444,N_9854);
or U12869 (N_12869,N_10784,N_11405);
or U12870 (N_12870,N_10289,N_10650);
nor U12871 (N_12871,N_9860,N_9810);
and U12872 (N_12872,N_12223,N_11953);
or U12873 (N_12873,N_11304,N_10282);
nand U12874 (N_12874,N_9845,N_12434);
nand U12875 (N_12875,N_10101,N_10309);
nand U12876 (N_12876,N_12187,N_9724);
nand U12877 (N_12877,N_10640,N_10186);
nand U12878 (N_12878,N_10605,N_10587);
and U12879 (N_12879,N_10804,N_11780);
nor U12880 (N_12880,N_9792,N_11038);
and U12881 (N_12881,N_11800,N_12254);
nor U12882 (N_12882,N_11765,N_10839);
and U12883 (N_12883,N_11040,N_12291);
nor U12884 (N_12884,N_11296,N_10721);
and U12885 (N_12885,N_9393,N_10783);
nor U12886 (N_12886,N_12120,N_9613);
and U12887 (N_12887,N_9457,N_11250);
nand U12888 (N_12888,N_10634,N_11518);
xnor U12889 (N_12889,N_10051,N_11665);
or U12890 (N_12890,N_9555,N_11512);
nor U12891 (N_12891,N_10642,N_11283);
nor U12892 (N_12892,N_11761,N_11436);
or U12893 (N_12893,N_10838,N_9401);
and U12894 (N_12894,N_10878,N_10518);
nand U12895 (N_12895,N_11193,N_11425);
nand U12896 (N_12896,N_11668,N_11114);
nand U12897 (N_12897,N_11566,N_12369);
and U12898 (N_12898,N_11771,N_10585);
nand U12899 (N_12899,N_11676,N_11086);
or U12900 (N_12900,N_11035,N_10434);
nor U12901 (N_12901,N_10214,N_10706);
nor U12902 (N_12902,N_11419,N_11693);
nand U12903 (N_12903,N_10375,N_10083);
nand U12904 (N_12904,N_10652,N_10436);
nor U12905 (N_12905,N_9488,N_10644);
xnor U12906 (N_12906,N_10480,N_10569);
nand U12907 (N_12907,N_11933,N_11657);
and U12908 (N_12908,N_12406,N_9641);
and U12909 (N_12909,N_12134,N_11087);
nand U12910 (N_12910,N_11825,N_10980);
nand U12911 (N_12911,N_10718,N_12024);
nor U12912 (N_12912,N_9929,N_12419);
nor U12913 (N_12913,N_11154,N_10827);
or U12914 (N_12914,N_11104,N_10731);
nor U12915 (N_12915,N_10814,N_11180);
or U12916 (N_12916,N_9916,N_9819);
nand U12917 (N_12917,N_11621,N_9527);
nand U12918 (N_12918,N_11445,N_9465);
xor U12919 (N_12919,N_12423,N_10516);
and U12920 (N_12920,N_11627,N_10925);
nor U12921 (N_12921,N_10828,N_12405);
or U12922 (N_12922,N_11536,N_12292);
and U12923 (N_12923,N_12010,N_12062);
nand U12924 (N_12924,N_9835,N_10631);
or U12925 (N_12925,N_11388,N_10683);
nor U12926 (N_12926,N_9754,N_11475);
or U12927 (N_12927,N_10003,N_9452);
nor U12928 (N_12928,N_11837,N_11532);
or U12929 (N_12929,N_10825,N_12295);
xor U12930 (N_12930,N_9812,N_11438);
or U12931 (N_12931,N_9463,N_11555);
nand U12932 (N_12932,N_9414,N_12385);
or U12933 (N_12933,N_10345,N_11478);
nand U12934 (N_12934,N_11973,N_12465);
nor U12935 (N_12935,N_11952,N_10532);
xor U12936 (N_12936,N_11572,N_11412);
xnor U12937 (N_12937,N_11647,N_9918);
nor U12938 (N_12938,N_10775,N_9960);
nor U12939 (N_12939,N_11257,N_10049);
nor U12940 (N_12940,N_11849,N_9903);
nand U12941 (N_12941,N_11743,N_9928);
xnor U12942 (N_12942,N_10540,N_11495);
or U12943 (N_12943,N_10511,N_12142);
nand U12944 (N_12944,N_11870,N_10549);
nor U12945 (N_12945,N_11343,N_9853);
nor U12946 (N_12946,N_11465,N_11551);
nand U12947 (N_12947,N_11416,N_10629);
nand U12948 (N_12948,N_11235,N_11847);
nand U12949 (N_12949,N_9753,N_11598);
or U12950 (N_12950,N_10351,N_12150);
and U12951 (N_12951,N_11712,N_10817);
nor U12952 (N_12952,N_11511,N_11246);
nor U12953 (N_12953,N_9670,N_12210);
xnor U12954 (N_12954,N_10360,N_10045);
or U12955 (N_12955,N_10144,N_10029);
or U12956 (N_12956,N_11989,N_9767);
nor U12957 (N_12957,N_9777,N_11080);
nor U12958 (N_12958,N_10158,N_10651);
and U12959 (N_12959,N_10664,N_11432);
nor U12960 (N_12960,N_11323,N_10620);
or U12961 (N_12961,N_10506,N_11020);
nor U12962 (N_12962,N_11561,N_9834);
and U12963 (N_12963,N_10222,N_10081);
nor U12964 (N_12964,N_9793,N_9403);
nor U12965 (N_12965,N_9419,N_11052);
and U12966 (N_12966,N_9446,N_11406);
or U12967 (N_12967,N_11836,N_10184);
nand U12968 (N_12968,N_9791,N_12286);
or U12969 (N_12969,N_10019,N_9804);
or U12970 (N_12970,N_12137,N_12282);
nand U12971 (N_12971,N_11958,N_11249);
nor U12972 (N_12972,N_12125,N_10687);
and U12973 (N_12973,N_10788,N_11862);
and U12974 (N_12974,N_11517,N_10169);
nand U12975 (N_12975,N_9687,N_9938);
nor U12976 (N_12976,N_10377,N_10085);
nor U12977 (N_12977,N_10762,N_11363);
and U12978 (N_12978,N_10100,N_9862);
nor U12979 (N_12979,N_12165,N_11964);
or U12980 (N_12980,N_10056,N_9530);
or U12981 (N_12981,N_9961,N_11085);
or U12982 (N_12982,N_9722,N_10697);
or U12983 (N_12983,N_10743,N_9538);
nand U12984 (N_12984,N_11695,N_11542);
or U12985 (N_12985,N_10311,N_9511);
nand U12986 (N_12986,N_10466,N_11783);
or U12987 (N_12987,N_9971,N_11570);
and U12988 (N_12988,N_11496,N_11785);
and U12989 (N_12989,N_11029,N_11727);
xnor U12990 (N_12990,N_10798,N_12231);
or U12991 (N_12991,N_12340,N_9481);
nand U12992 (N_12992,N_9781,N_10898);
and U12993 (N_12993,N_11396,N_12033);
nor U12994 (N_12994,N_10577,N_9409);
and U12995 (N_12995,N_11274,N_11145);
and U12996 (N_12996,N_9563,N_10249);
nand U12997 (N_12997,N_11595,N_10203);
nand U12998 (N_12998,N_9579,N_11339);
or U12999 (N_12999,N_11775,N_10785);
and U13000 (N_13000,N_10848,N_12489);
and U13001 (N_13001,N_10316,N_10394);
nand U13002 (N_13002,N_12453,N_10484);
nor U13003 (N_13003,N_9717,N_10978);
and U13004 (N_13004,N_10376,N_10011);
nand U13005 (N_13005,N_11034,N_9378);
nor U13006 (N_13006,N_12390,N_12356);
or U13007 (N_13007,N_11774,N_10679);
nor U13008 (N_13008,N_11141,N_9994);
and U13009 (N_13009,N_10904,N_11863);
or U13010 (N_13010,N_10416,N_10325);
nand U13011 (N_13011,N_12065,N_11696);
nor U13012 (N_13012,N_9410,N_11677);
nor U13013 (N_13013,N_10710,N_12242);
and U13014 (N_13014,N_10488,N_9582);
and U13015 (N_13015,N_11302,N_10292);
and U13016 (N_13016,N_11508,N_10526);
or U13017 (N_13017,N_11252,N_11003);
xnor U13018 (N_13018,N_10889,N_10013);
nor U13019 (N_13019,N_12343,N_10373);
or U13020 (N_13020,N_10459,N_12173);
nand U13021 (N_13021,N_11752,N_10235);
or U13022 (N_13022,N_11719,N_11351);
or U13023 (N_13023,N_12371,N_11607);
nand U13024 (N_13024,N_10050,N_12485);
nand U13025 (N_13025,N_12219,N_11583);
and U13026 (N_13026,N_10795,N_9843);
xnor U13027 (N_13027,N_11977,N_11637);
or U13028 (N_13028,N_11642,N_11779);
and U13029 (N_13029,N_11310,N_10347);
and U13030 (N_13030,N_10088,N_9521);
and U13031 (N_13031,N_12256,N_9794);
nand U13032 (N_13032,N_10931,N_9806);
or U13033 (N_13033,N_11539,N_11358);
nor U13034 (N_13034,N_12314,N_10106);
and U13035 (N_13035,N_12315,N_9863);
and U13036 (N_13036,N_10809,N_10563);
xor U13037 (N_13037,N_11256,N_11305);
or U13038 (N_13038,N_11822,N_10010);
or U13039 (N_13039,N_11929,N_12474);
and U13040 (N_13040,N_10473,N_10616);
and U13041 (N_13041,N_12338,N_9441);
and U13042 (N_13042,N_11162,N_10772);
and U13043 (N_13043,N_12022,N_9492);
and U13044 (N_13044,N_12058,N_10304);
nand U13045 (N_13045,N_12109,N_12490);
xnor U13046 (N_13046,N_12388,N_10244);
nand U13047 (N_13047,N_10064,N_10746);
and U13048 (N_13048,N_9539,N_9931);
xnor U13049 (N_13049,N_9688,N_11279);
and U13050 (N_13050,N_9399,N_9890);
and U13051 (N_13051,N_9702,N_11155);
or U13052 (N_13052,N_10089,N_11549);
or U13053 (N_13053,N_11924,N_12009);
nand U13054 (N_13054,N_10887,N_10429);
nand U13055 (N_13055,N_12263,N_9692);
and U13056 (N_13056,N_10658,N_11099);
nor U13057 (N_13057,N_10739,N_11291);
nor U13058 (N_13058,N_11996,N_9827);
and U13059 (N_13059,N_11265,N_9591);
or U13060 (N_13060,N_11359,N_9626);
and U13061 (N_13061,N_11428,N_10986);
nor U13062 (N_13062,N_12237,N_12279);
nor U13063 (N_13063,N_9922,N_11172);
nand U13064 (N_13064,N_10938,N_11284);
or U13065 (N_13065,N_10221,N_10719);
and U13066 (N_13066,N_9871,N_11289);
xor U13067 (N_13067,N_11224,N_11658);
and U13068 (N_13068,N_11126,N_10550);
nor U13069 (N_13069,N_12098,N_10486);
xor U13070 (N_13070,N_11179,N_11264);
or U13071 (N_13071,N_9764,N_10318);
or U13072 (N_13072,N_12335,N_10530);
nor U13073 (N_13073,N_11723,N_10656);
nor U13074 (N_13074,N_9586,N_11335);
or U13075 (N_13075,N_12322,N_9710);
xor U13076 (N_13076,N_12442,N_11387);
nand U13077 (N_13077,N_9733,N_12304);
or U13078 (N_13078,N_10027,N_11959);
nand U13079 (N_13079,N_10695,N_11663);
or U13080 (N_13080,N_10969,N_10093);
nand U13081 (N_13081,N_11400,N_11801);
or U13082 (N_13082,N_11112,N_12270);
and U13083 (N_13083,N_10987,N_11075);
or U13084 (N_13084,N_10843,N_11690);
and U13085 (N_13085,N_12461,N_12265);
and U13086 (N_13086,N_10420,N_11553);
nor U13087 (N_13087,N_11002,N_11525);
and U13088 (N_13088,N_11574,N_11942);
nand U13089 (N_13089,N_9678,N_11597);
xnor U13090 (N_13090,N_11698,N_9756);
xnor U13091 (N_13091,N_11789,N_10411);
nor U13092 (N_13092,N_11307,N_12477);
nor U13093 (N_13093,N_11136,N_11435);
or U13094 (N_13094,N_11982,N_9450);
nor U13095 (N_13095,N_10110,N_10984);
or U13096 (N_13096,N_10499,N_9432);
nor U13097 (N_13097,N_10566,N_10414);
nor U13098 (N_13098,N_10531,N_10623);
or U13099 (N_13099,N_10596,N_10439);
nor U13100 (N_13100,N_9385,N_10217);
and U13101 (N_13101,N_10392,N_10241);
nor U13102 (N_13102,N_10388,N_9876);
and U13103 (N_13103,N_11083,N_9970);
xor U13104 (N_13104,N_9825,N_11531);
xnor U13105 (N_13105,N_9763,N_9780);
xor U13106 (N_13106,N_9528,N_9400);
nand U13107 (N_13107,N_12193,N_12121);
and U13108 (N_13108,N_11998,N_9898);
xor U13109 (N_13109,N_11619,N_11499);
or U13110 (N_13110,N_12311,N_11460);
or U13111 (N_13111,N_12092,N_9543);
and U13112 (N_13112,N_10595,N_10166);
and U13113 (N_13113,N_10493,N_12195);
nor U13114 (N_13114,N_11331,N_9979);
or U13115 (N_13115,N_10729,N_10561);
or U13116 (N_13116,N_10366,N_9772);
nand U13117 (N_13117,N_10400,N_10575);
and U13118 (N_13118,N_10405,N_9558);
and U13119 (N_13119,N_11987,N_11587);
and U13120 (N_13120,N_11804,N_11135);
nand U13121 (N_13121,N_10456,N_11493);
and U13122 (N_13122,N_11153,N_11672);
nand U13123 (N_13123,N_11872,N_12358);
nand U13124 (N_13124,N_10918,N_10643);
and U13125 (N_13125,N_9504,N_10446);
xnor U13126 (N_13126,N_10343,N_11271);
xor U13127 (N_13127,N_10077,N_10079);
and U13128 (N_13128,N_11417,N_11612);
and U13129 (N_13129,N_11747,N_9445);
nand U13130 (N_13130,N_12190,N_12466);
nand U13131 (N_13131,N_10815,N_10554);
nand U13132 (N_13132,N_10756,N_10454);
nor U13133 (N_13133,N_10633,N_10654);
nand U13134 (N_13134,N_12174,N_12006);
nor U13135 (N_13135,N_9879,N_9673);
nand U13136 (N_13136,N_9981,N_10451);
or U13137 (N_13137,N_12091,N_9966);
nand U13138 (N_13138,N_11449,N_10188);
or U13139 (N_13139,N_10404,N_11684);
nor U13140 (N_13140,N_9847,N_12170);
nor U13141 (N_13141,N_11620,N_11700);
and U13142 (N_13142,N_10708,N_11624);
nor U13143 (N_13143,N_10613,N_9882);
xnor U13144 (N_13144,N_11479,N_12228);
nand U13145 (N_13145,N_10913,N_11059);
nand U13146 (N_13146,N_10807,N_10271);
and U13147 (N_13147,N_11266,N_11791);
xnor U13148 (N_13148,N_10693,N_11222);
or U13149 (N_13149,N_10437,N_10567);
and U13150 (N_13150,N_9896,N_9398);
and U13151 (N_13151,N_11772,N_10632);
nor U13152 (N_13152,N_11852,N_11111);
nor U13153 (N_13153,N_10692,N_10946);
nor U13154 (N_13154,N_9778,N_12320);
nand U13155 (N_13155,N_12469,N_11492);
nand U13156 (N_13156,N_11362,N_12364);
nor U13157 (N_13157,N_10571,N_9643);
xnor U13158 (N_13158,N_12102,N_10661);
and U13159 (N_13159,N_10597,N_10409);
or U13160 (N_13160,N_10258,N_11427);
nand U13161 (N_13161,N_9836,N_10579);
nor U13162 (N_13162,N_10386,N_9505);
nor U13163 (N_13163,N_10558,N_9502);
nor U13164 (N_13164,N_10757,N_11414);
or U13165 (N_13165,N_9426,N_10998);
nand U13166 (N_13166,N_10448,N_9705);
nor U13167 (N_13167,N_11313,N_10771);
or U13168 (N_13168,N_10193,N_10264);
nand U13169 (N_13169,N_10036,N_10468);
or U13170 (N_13170,N_9880,N_11344);
nor U13171 (N_13171,N_9473,N_11078);
nand U13172 (N_13172,N_10592,N_10007);
or U13173 (N_13173,N_10907,N_12498);
xnor U13174 (N_13174,N_10403,N_9969);
and U13175 (N_13175,N_11450,N_9762);
nor U13176 (N_13176,N_11562,N_9855);
and U13177 (N_13177,N_11565,N_11226);
nor U13178 (N_13178,N_11701,N_12475);
nand U13179 (N_13179,N_9392,N_9779);
and U13180 (N_13180,N_11869,N_10168);
nor U13181 (N_13181,N_10280,N_12205);
nand U13182 (N_13182,N_10744,N_9635);
nor U13183 (N_13183,N_9499,N_12328);
nand U13184 (N_13184,N_9679,N_9541);
and U13185 (N_13185,N_11769,N_10113);
nor U13186 (N_13186,N_12181,N_10630);
xnor U13187 (N_13187,N_10148,N_10742);
nor U13188 (N_13188,N_11287,N_11947);
nor U13189 (N_13189,N_10586,N_10382);
xnor U13190 (N_13190,N_10209,N_12260);
nor U13191 (N_13191,N_9436,N_10267);
or U13192 (N_13192,N_9606,N_10167);
xor U13193 (N_13193,N_9978,N_9389);
or U13194 (N_13194,N_9526,N_12015);
or U13195 (N_13195,N_12026,N_12145);
nand U13196 (N_13196,N_10924,N_11244);
xnor U13197 (N_13197,N_9620,N_11370);
nor U13198 (N_13198,N_12044,N_10035);
and U13199 (N_13199,N_12402,N_10365);
or U13200 (N_13200,N_10568,N_11476);
and U13201 (N_13201,N_12400,N_10874);
xor U13202 (N_13202,N_9518,N_10606);
nand U13203 (N_13203,N_10684,N_11463);
nand U13204 (N_13204,N_9958,N_12032);
xnor U13205 (N_13205,N_11030,N_10749);
and U13206 (N_13206,N_11348,N_11430);
nor U13207 (N_13207,N_11860,N_9656);
and U13208 (N_13208,N_11781,N_11000);
nand U13209 (N_13209,N_10552,N_12066);
nor U13210 (N_13210,N_9634,N_12403);
or U13211 (N_13211,N_10194,N_9921);
or U13212 (N_13212,N_9999,N_9850);
or U13213 (N_13213,N_11711,N_11937);
nand U13214 (N_13214,N_11336,N_12025);
or U13215 (N_13215,N_9599,N_10057);
or U13216 (N_13216,N_9919,N_11921);
and U13217 (N_13217,N_11813,N_10327);
or U13218 (N_13218,N_12308,N_10254);
or U13219 (N_13219,N_9714,N_9698);
and U13220 (N_13220,N_12023,N_11891);
or U13221 (N_13221,N_11320,N_11834);
xnor U13222 (N_13222,N_10397,N_10461);
and U13223 (N_13223,N_10033,N_10061);
nand U13224 (N_13224,N_11184,N_11591);
or U13225 (N_13225,N_11423,N_9593);
xnor U13226 (N_13226,N_10418,N_10123);
nand U13227 (N_13227,N_11928,N_11187);
nand U13228 (N_13228,N_11384,N_9811);
or U13229 (N_13229,N_11397,N_11461);
or U13230 (N_13230,N_11202,N_12152);
and U13231 (N_13231,N_9654,N_9404);
or U13232 (N_13232,N_11802,N_11297);
and U13233 (N_13233,N_10307,N_11729);
and U13234 (N_13234,N_12481,N_10926);
nand U13235 (N_13235,N_12264,N_11540);
xor U13236 (N_13236,N_10911,N_12283);
nor U13237 (N_13237,N_11588,N_10612);
nand U13238 (N_13238,N_10997,N_11689);
or U13239 (N_13239,N_11550,N_10256);
and U13240 (N_13240,N_10787,N_10820);
nor U13241 (N_13241,N_9485,N_11241);
nand U13242 (N_13242,N_11615,N_9809);
or U13243 (N_13243,N_12339,N_11434);
and U13244 (N_13244,N_10614,N_12073);
nand U13245 (N_13245,N_11468,N_12413);
nand U13246 (N_13246,N_11215,N_10922);
nor U13247 (N_13247,N_10442,N_11044);
or U13248 (N_13248,N_11230,N_12259);
nor U13249 (N_13249,N_9406,N_11170);
nor U13250 (N_13250,N_12424,N_10103);
or U13251 (N_13251,N_11318,N_11228);
nor U13252 (N_13252,N_9861,N_11628);
and U13253 (N_13253,N_11972,N_9466);
nand U13254 (N_13254,N_10851,N_12069);
nor U13255 (N_13255,N_12352,N_9549);
xor U13256 (N_13256,N_11220,N_11527);
nor U13257 (N_13257,N_11795,N_11622);
and U13258 (N_13258,N_10213,N_10424);
or U13259 (N_13259,N_9877,N_9646);
or U13260 (N_13260,N_12194,N_12337);
or U13261 (N_13261,N_10533,N_10255);
nor U13262 (N_13262,N_12046,N_11196);
nor U13263 (N_13263,N_10861,N_10075);
and U13264 (N_13264,N_9675,N_9387);
xor U13265 (N_13265,N_11488,N_11182);
nand U13266 (N_13266,N_11019,N_12452);
nand U13267 (N_13267,N_10504,N_12148);
or U13268 (N_13268,N_11403,N_9379);
and U13269 (N_13269,N_11163,N_12317);
or U13270 (N_13270,N_10287,N_10151);
nand U13271 (N_13271,N_11997,N_10328);
nor U13272 (N_13272,N_10131,N_9655);
nor U13273 (N_13273,N_9509,N_11456);
xnor U13274 (N_13274,N_10748,N_9666);
or U13275 (N_13275,N_11903,N_11592);
nor U13276 (N_13276,N_12207,N_11916);
and U13277 (N_13277,N_12394,N_9609);
nor U13278 (N_13278,N_10853,N_12336);
or U13279 (N_13279,N_12110,N_11716);
or U13280 (N_13280,N_10095,N_9551);
nor U13281 (N_13281,N_11513,N_11383);
nor U13282 (N_13282,N_9573,N_11948);
and U13283 (N_13283,N_10155,N_11760);
and U13284 (N_13284,N_10522,N_12083);
xor U13285 (N_13285,N_11379,N_10893);
nor U13286 (N_13286,N_9852,N_12301);
xor U13287 (N_13287,N_10462,N_11569);
or U13288 (N_13288,N_12191,N_12146);
nor U13289 (N_13289,N_11968,N_10680);
nor U13290 (N_13290,N_10734,N_10888);
nand U13291 (N_13291,N_9972,N_10417);
or U13292 (N_13292,N_11956,N_12198);
or U13293 (N_13293,N_11979,N_11175);
nand U13294 (N_13294,N_10647,N_11516);
or U13295 (N_13295,N_9842,N_10006);
or U13296 (N_13296,N_9575,N_12127);
nand U13297 (N_13297,N_12313,N_9557);
xor U13298 (N_13298,N_10832,N_11382);
and U13299 (N_13299,N_12086,N_10384);
nand U13300 (N_13300,N_9413,N_10385);
nand U13301 (N_13301,N_10957,N_10072);
or U13302 (N_13302,N_10467,N_11820);
and U13303 (N_13303,N_10580,N_11166);
and U13304 (N_13304,N_12325,N_10305);
xnor U13305 (N_13305,N_11143,N_11309);
nand U13306 (N_13306,N_10716,N_11232);
nand U13307 (N_13307,N_11720,N_11741);
nand U13308 (N_13308,N_11276,N_11270);
nand U13309 (N_13309,N_10780,N_10133);
or U13310 (N_13310,N_10621,N_11606);
nor U13311 (N_13311,N_9699,N_11971);
and U13312 (N_13312,N_10778,N_9851);
xnor U13313 (N_13313,N_11366,N_9897);
nand U13314 (N_13314,N_10714,N_9416);
nand U13315 (N_13315,N_11934,N_12232);
nand U13316 (N_13316,N_11341,N_11631);
and U13317 (N_13317,N_9761,N_10736);
and U13318 (N_13318,N_11778,N_12393);
nand U13319 (N_13319,N_12378,N_10475);
and U13320 (N_13320,N_12445,N_12084);
or U13321 (N_13321,N_9703,N_11337);
and U13322 (N_13322,N_9382,N_10046);
nor U13323 (N_13323,N_9736,N_11165);
or U13324 (N_13324,N_10992,N_11976);
nand U13325 (N_13325,N_11079,N_12365);
nor U13326 (N_13326,N_9908,N_9695);
and U13327 (N_13327,N_11816,N_10603);
nand U13328 (N_13328,N_10675,N_11744);
nand U13329 (N_13329,N_10983,N_9801);
or U13330 (N_13330,N_12029,N_12451);
or U13331 (N_13331,N_10857,N_11470);
and U13332 (N_13332,N_12487,N_10216);
nor U13333 (N_13333,N_11231,N_10525);
nand U13334 (N_13334,N_10681,N_9786);
and U13335 (N_13335,N_12082,N_11134);
xor U13336 (N_13336,N_11645,N_10951);
nand U13337 (N_13337,N_11842,N_9650);
nand U13338 (N_13338,N_10135,N_11409);
nor U13339 (N_13339,N_11935,N_9973);
nor U13340 (N_13340,N_12441,N_11737);
nor U13341 (N_13341,N_12327,N_9948);
nand U13342 (N_13342,N_11043,N_9738);
and U13343 (N_13343,N_12410,N_10163);
nand U13344 (N_13344,N_12437,N_9813);
nand U13345 (N_13345,N_9739,N_10018);
or U13346 (N_13346,N_11567,N_12408);
nor U13347 (N_13347,N_11907,N_9817);
nor U13348 (N_13348,N_12039,N_9552);
nor U13349 (N_13349,N_9636,N_9564);
or U13350 (N_13350,N_11093,N_10869);
and U13351 (N_13351,N_11560,N_12011);
nand U13352 (N_13352,N_12310,N_10396);
or U13353 (N_13353,N_9837,N_11648);
nand U13354 (N_13354,N_9735,N_12067);
nor U13355 (N_13355,N_11717,N_11514);
nor U13356 (N_13356,N_11156,N_12456);
nor U13357 (N_13357,N_10335,N_10231);
nor U13358 (N_13358,N_12368,N_10691);
nor U13359 (N_13359,N_11139,N_10582);
nor U13360 (N_13360,N_11295,N_12216);
nand U13361 (N_13361,N_11216,N_10965);
nand U13362 (N_13362,N_9983,N_11828);
nand U13363 (N_13363,N_11477,N_9802);
or U13364 (N_13364,N_11799,N_10243);
nand U13365 (N_13365,N_9682,N_12249);
xnor U13366 (N_13366,N_10602,N_12417);
nand U13367 (N_13367,N_11253,N_10786);
nand U13368 (N_13368,N_9881,N_11227);
xor U13369 (N_13369,N_11212,N_11888);
nand U13370 (N_13370,N_11404,N_11901);
or U13371 (N_13371,N_9664,N_10747);
nor U13372 (N_13372,N_9925,N_11880);
or U13373 (N_13373,N_12101,N_11630);
nand U13374 (N_13374,N_10207,N_11833);
and U13375 (N_13375,N_10909,N_9993);
or U13376 (N_13376,N_12211,N_9434);
and U13377 (N_13377,N_9700,N_10537);
nor U13378 (N_13378,N_11448,N_9546);
xor U13379 (N_13379,N_9775,N_11556);
and U13380 (N_13380,N_10551,N_11881);
xnor U13381 (N_13381,N_11733,N_10157);
nor U13382 (N_13382,N_10313,N_12054);
or U13383 (N_13383,N_12269,N_11746);
and U13384 (N_13384,N_12063,N_10707);
and U13385 (N_13385,N_10192,N_12246);
nand U13386 (N_13386,N_9621,N_11333);
nor U13387 (N_13387,N_9985,N_10513);
nor U13388 (N_13388,N_10165,N_9377);
and U13389 (N_13389,N_11167,N_9944);
or U13390 (N_13390,N_11191,N_10196);
or U13391 (N_13391,N_11740,N_12213);
or U13392 (N_13392,N_10763,N_10337);
xnor U13393 (N_13393,N_10296,N_10677);
and U13394 (N_13394,N_10334,N_11832);
or U13395 (N_13395,N_10781,N_12007);
and U13396 (N_13396,N_11137,N_11738);
and U13397 (N_13397,N_11028,N_11936);
nand U13398 (N_13398,N_9936,N_12459);
or U13399 (N_13399,N_10657,N_10723);
nand U13400 (N_13400,N_11149,N_12097);
and U13401 (N_13401,N_9940,N_10841);
nor U13402 (N_13402,N_10399,N_10501);
or U13403 (N_13403,N_9623,N_12215);
nor U13404 (N_13404,N_12342,N_9639);
or U13405 (N_13405,N_12157,N_11584);
nand U13406 (N_13406,N_9581,N_10285);
nand U13407 (N_13407,N_11415,N_10557);
xnor U13408 (N_13408,N_11616,N_11095);
or U13409 (N_13409,N_11263,N_12350);
nand U13410 (N_13410,N_12379,N_9588);
or U13411 (N_13411,N_10161,N_12341);
nor U13412 (N_13412,N_11954,N_10358);
or U13413 (N_13413,N_12154,N_12454);
nor U13414 (N_13414,N_9532,N_9388);
nor U13415 (N_13415,N_11609,N_11411);
or U13416 (N_13416,N_10202,N_11835);
or U13417 (N_13417,N_11967,N_10326);
xor U13418 (N_13418,N_10042,N_11889);
or U13419 (N_13419,N_12470,N_10932);
or U13420 (N_13420,N_9829,N_11601);
and U13421 (N_13421,N_9390,N_9498);
xnor U13422 (N_13422,N_9420,N_10180);
nor U13423 (N_13423,N_11505,N_12095);
xnor U13424 (N_13424,N_10431,N_10268);
nand U13425 (N_13425,N_11981,N_11811);
and U13426 (N_13426,N_9839,N_9604);
or U13427 (N_13427,N_11840,N_10520);
nor U13428 (N_13428,N_11614,N_9625);
or U13429 (N_13429,N_9758,N_12151);
nand U13430 (N_13430,N_11626,N_11064);
nand U13431 (N_13431,N_12458,N_9730);
and U13432 (N_13432,N_11661,N_11115);
and U13433 (N_13433,N_10635,N_10303);
or U13434 (N_13434,N_12495,N_11908);
or U13435 (N_13435,N_11897,N_12043);
nor U13436 (N_13436,N_11489,N_11110);
xor U13437 (N_13437,N_11625,N_10699);
or U13438 (N_13438,N_11486,N_11186);
nand U13439 (N_13439,N_12240,N_11963);
nor U13440 (N_13440,N_9589,N_9632);
nor U13441 (N_13441,N_10884,N_12057);
nor U13442 (N_13442,N_9428,N_11667);
nand U13443 (N_13443,N_11353,N_10227);
nand U13444 (N_13444,N_9422,N_11308);
and U13445 (N_13445,N_10391,N_11662);
nor U13446 (N_13446,N_11509,N_9444);
and U13447 (N_13447,N_10272,N_12053);
and U13448 (N_13448,N_9417,N_9867);
nor U13449 (N_13449,N_9706,N_11364);
and U13450 (N_13450,N_10323,N_11324);
and U13451 (N_13451,N_10598,N_9597);
or U13452 (N_13452,N_11732,N_9883);
xnor U13453 (N_13453,N_10646,N_12303);
nand U13454 (N_13454,N_9732,N_10248);
nand U13455 (N_13455,N_11022,N_10519);
and U13456 (N_13456,N_9560,N_12253);
nand U13457 (N_13457,N_10177,N_11638);
and U13458 (N_13458,N_10590,N_11839);
nor U13459 (N_13459,N_9719,N_10438);
and U13460 (N_13460,N_10875,N_10806);
and U13461 (N_13461,N_11392,N_11072);
and U13462 (N_13462,N_9765,N_10290);
and U13463 (N_13463,N_11938,N_11814);
nand U13464 (N_13464,N_11429,N_10588);
xor U13465 (N_13465,N_10769,N_12432);
nor U13466 (N_13466,N_11885,N_9894);
and U13467 (N_13467,N_11756,N_11120);
or U13468 (N_13468,N_12008,N_12167);
or U13469 (N_13469,N_12499,N_12028);
and U13470 (N_13470,N_12380,N_11519);
nor U13471 (N_13471,N_11194,N_9773);
or U13472 (N_13472,N_11398,N_11617);
and U13473 (N_13473,N_9926,N_10331);
nor U13474 (N_13474,N_12143,N_11278);
xnor U13475 (N_13475,N_9516,N_11824);
nand U13476 (N_13476,N_11117,N_11582);
or U13477 (N_13477,N_10286,N_10441);
or U13478 (N_13478,N_9439,N_9651);
nand U13479 (N_13479,N_9721,N_9912);
and U13480 (N_13480,N_12318,N_9932);
xnor U13481 (N_13481,N_11596,N_11829);
and U13482 (N_13482,N_10164,N_10981);
nand U13483 (N_13483,N_10759,N_11164);
nor U13484 (N_13484,N_9459,N_11181);
xor U13485 (N_13485,N_10545,N_11742);
xnor U13486 (N_13486,N_11354,N_9734);
nor U13487 (N_13487,N_11575,N_10230);
xor U13488 (N_13488,N_11749,N_11962);
and U13489 (N_13489,N_9536,N_12224);
and U13490 (N_13490,N_10538,N_11144);
or U13491 (N_13491,N_10240,N_11786);
nand U13492 (N_13492,N_11943,N_10239);
nand U13493 (N_13493,N_11233,N_10599);
nor U13494 (N_13494,N_11900,N_11454);
or U13495 (N_13495,N_11380,N_11490);
or U13496 (N_13496,N_12163,N_12486);
xor U13497 (N_13497,N_10917,N_12395);
nand U13498 (N_13498,N_12316,N_10108);
or U13499 (N_13499,N_12349,N_10025);
or U13500 (N_13500,N_11812,N_10350);
or U13501 (N_13501,N_11564,N_10688);
nor U13502 (N_13502,N_9974,N_11850);
nand U13503 (N_13503,N_10374,N_11169);
or U13504 (N_13504,N_10665,N_12178);
nand U13505 (N_13505,N_10189,N_12300);
xnor U13506 (N_13506,N_11554,N_10380);
and U13507 (N_13507,N_11151,N_9649);
xnor U13508 (N_13508,N_11745,N_10252);
or U13509 (N_13509,N_11070,N_9583);
nor U13510 (N_13510,N_10600,N_10799);
and U13511 (N_13511,N_10791,N_9816);
nor U13512 (N_13512,N_10229,N_9472);
xnor U13513 (N_13513,N_12435,N_12309);
nor U13514 (N_13514,N_10415,N_10840);
and U13515 (N_13515,N_11882,N_11524);
nor U13516 (N_13516,N_9774,N_9449);
nand U13517 (N_13517,N_9795,N_11762);
nor U13518 (N_13518,N_11794,N_12071);
and U13519 (N_13519,N_11269,N_11107);
nand U13520 (N_13520,N_11189,N_10810);
xnor U13521 (N_13521,N_12155,N_10479);
xor U13522 (N_13522,N_10195,N_10465);
or U13523 (N_13523,N_10662,N_9460);
nand U13524 (N_13524,N_9823,N_9493);
or U13525 (N_13525,N_11332,N_11507);
and U13526 (N_13526,N_10440,N_9515);
or U13527 (N_13527,N_10338,N_10968);
or U13528 (N_13528,N_10278,N_10864);
or U13529 (N_13529,N_11632,N_11446);
nand U13530 (N_13530,N_10000,N_11949);
and U13531 (N_13531,N_10430,N_12184);
nand U13532 (N_13532,N_9784,N_10776);
and U13533 (N_13533,N_10299,N_12271);
xnor U13534 (N_13534,N_10709,N_11945);
nor U13535 (N_13535,N_11768,N_11629);
nor U13536 (N_13536,N_11147,N_9749);
and U13537 (N_13537,N_11871,N_10833);
xor U13538 (N_13538,N_10962,N_10175);
or U13539 (N_13539,N_9885,N_11062);
nor U13540 (N_13540,N_10408,N_12276);
nor U13541 (N_13541,N_12016,N_9715);
nand U13542 (N_13542,N_11389,N_11131);
nand U13543 (N_13543,N_12274,N_10130);
nand U13544 (N_13544,N_10421,N_11140);
nor U13545 (N_13545,N_10125,N_10279);
or U13546 (N_13546,N_10900,N_12096);
nor U13547 (N_13547,N_11545,N_10333);
or U13548 (N_13548,N_11734,N_10655);
nand U13549 (N_13549,N_10611,N_10698);
nand U13550 (N_13550,N_10866,N_11843);
and U13551 (N_13551,N_9561,N_11706);
and U13552 (N_13552,N_11634,N_12396);
or U13553 (N_13553,N_10822,N_10116);
nand U13554 (N_13554,N_9553,N_12439);
nand U13555 (N_13555,N_11418,N_11721);
or U13556 (N_13556,N_12387,N_10648);
nor U13557 (N_13557,N_9920,N_10273);
and U13558 (N_13558,N_9545,N_9384);
nor U13559 (N_13559,N_11688,N_10002);
or U13560 (N_13560,N_9615,N_11770);
xnor U13561 (N_13561,N_10790,N_12488);
nand U13562 (N_13562,N_10831,N_10676);
xor U13563 (N_13563,N_12494,N_12004);
nor U13564 (N_13564,N_9383,N_12052);
nor U13565 (N_13565,N_9744,N_10260);
and U13566 (N_13566,N_11650,N_12122);
nand U13567 (N_13567,N_9776,N_9548);
nand U13568 (N_13568,N_9534,N_12305);
nand U13569 (N_13569,N_10363,N_11441);
xor U13570 (N_13570,N_12415,N_10715);
xnor U13571 (N_13571,N_10054,N_10636);
nor U13572 (N_13572,N_11031,N_10330);
or U13573 (N_13573,N_9723,N_10751);
and U13574 (N_13574,N_11026,N_11699);
nand U13575 (N_13575,N_12346,N_10500);
or U13576 (N_13576,N_11764,N_12235);
or U13577 (N_13577,N_10368,N_12103);
and U13578 (N_13578,N_9568,N_11056);
and U13579 (N_13579,N_10401,N_10039);
nand U13580 (N_13580,N_12014,N_10574);
nor U13581 (N_13581,N_9519,N_10523);
nand U13582 (N_13582,N_12131,N_12189);
nand U13583 (N_13583,N_9814,N_11653);
nor U13584 (N_13584,N_9954,N_10226);
and U13585 (N_13585,N_11408,N_11797);
nand U13586 (N_13586,N_9479,N_10076);
nor U13587 (N_13587,N_10615,N_9689);
nor U13588 (N_13588,N_9750,N_9849);
and U13589 (N_13589,N_11298,N_11442);
or U13590 (N_13590,N_10136,N_9567);
nand U13591 (N_13591,N_12376,N_10232);
and U13592 (N_13592,N_12100,N_11685);
and U13593 (N_13593,N_10935,N_11528);
nor U13594 (N_13594,N_12244,N_11790);
nor U13595 (N_13595,N_12334,N_11272);
or U13596 (N_13596,N_11094,N_12389);
nor U13597 (N_13597,N_9610,N_10139);
xor U13598 (N_13598,N_11204,N_10758);
nand U13599 (N_13599,N_12214,N_10930);
xor U13600 (N_13600,N_11669,N_10445);
nand U13601 (N_13601,N_11369,N_12258);
xor U13602 (N_13602,N_11097,N_9483);
xor U13603 (N_13603,N_9796,N_11494);
and U13604 (N_13604,N_10026,N_12153);
nor U13605 (N_13605,N_9930,N_10541);
nand U13606 (N_13606,N_10134,N_11033);
nand U13607 (N_13607,N_10617,N_10885);
nor U13608 (N_13608,N_10369,N_11459);
nand U13609 (N_13609,N_11178,N_12227);
nand U13610 (N_13610,N_11932,N_11679);
or U13611 (N_13611,N_11910,N_12049);
nor U13612 (N_13612,N_11422,N_11557);
or U13613 (N_13613,N_11618,N_12243);
nor U13614 (N_13614,N_11355,N_10223);
nor U13615 (N_13615,N_9668,N_10494);
and U13616 (N_13616,N_9694,N_11129);
nand U13617 (N_13617,N_9455,N_11223);
or U13618 (N_13618,N_11578,N_11613);
nor U13619 (N_13619,N_12319,N_9956);
or U13620 (N_13620,N_9906,N_10390);
xor U13621 (N_13621,N_9470,N_10543);
nand U13622 (N_13622,N_9585,N_10037);
nor U13623 (N_13623,N_10120,N_10449);
nand U13624 (N_13624,N_9693,N_9569);
nand U13625 (N_13625,N_10521,N_11487);
nor U13626 (N_13626,N_11541,N_11522);
nand U13627 (N_13627,N_9433,N_10584);
nor U13628 (N_13628,N_9759,N_9886);
or U13629 (N_13629,N_12355,N_10894);
nor U13630 (N_13630,N_11401,N_11190);
xnor U13631 (N_13631,N_12124,N_9992);
nand U13632 (N_13632,N_11731,N_10766);
xnor U13633 (N_13633,N_12272,N_10800);
nor U13634 (N_13634,N_9790,N_9408);
and U13635 (N_13635,N_9720,N_9873);
nor U13636 (N_13636,N_10882,N_11807);
or U13637 (N_13637,N_12347,N_11671);
xnor U13638 (N_13638,N_9988,N_10211);
or U13639 (N_13639,N_10094,N_9770);
and U13640 (N_13640,N_11758,N_10868);
nor U13641 (N_13641,N_11581,N_10996);
or U13642 (N_13642,N_10950,N_11798);
nand U13643 (N_13643,N_10773,N_10510);
nor U13644 (N_13644,N_10870,N_10419);
or U13645 (N_13645,N_11543,N_11602);
nor U13646 (N_13646,N_12398,N_11242);
and U13647 (N_13647,N_12126,N_11158);
xor U13648 (N_13648,N_11950,N_10191);
and U13649 (N_13649,N_9577,N_11334);
nand U13650 (N_13650,N_9821,N_10886);
or U13651 (N_13651,N_12372,N_10111);
and U13652 (N_13652,N_12404,N_11049);
nand U13653 (N_13653,N_11705,N_11096);
or U13654 (N_13654,N_10024,N_11103);
or U13655 (N_13655,N_12245,N_10087);
nor U13656 (N_13656,N_10738,N_10527);
or U13657 (N_13657,N_12031,N_11185);
xor U13658 (N_13658,N_12141,N_9603);
nand U13659 (N_13659,N_12281,N_10219);
and U13660 (N_13660,N_11913,N_11311);
or U13661 (N_13661,N_10638,N_12077);
xnor U13662 (N_13662,N_9824,N_11506);
or U13663 (N_13663,N_9858,N_10259);
nor U13664 (N_13664,N_11623,N_12072);
nor U13665 (N_13665,N_9506,N_11955);
and U13666 (N_13666,N_10854,N_10976);
nand U13667 (N_13667,N_12381,N_11130);
nor U13668 (N_13668,N_11051,N_11830);
nor U13669 (N_13669,N_10767,N_10919);
xor U13670 (N_13670,N_10801,N_12218);
xnor U13671 (N_13671,N_10768,N_10060);
nor U13672 (N_13672,N_11844,N_11826);
nor U13673 (N_13673,N_12051,N_10477);
nor U13674 (N_13674,N_9616,N_12070);
nand U13675 (N_13675,N_11902,N_12386);
xnor U13676 (N_13676,N_11157,N_10740);
nor U13677 (N_13677,N_11520,N_10354);
xor U13678 (N_13678,N_10863,N_12397);
and U13679 (N_13679,N_9782,N_12105);
nand U13680 (N_13680,N_10149,N_10796);
nor U13681 (N_13681,N_10752,N_11537);
or U13682 (N_13682,N_10952,N_12179);
and U13683 (N_13683,N_9833,N_11730);
or U13684 (N_13684,N_10953,N_11504);
nand U13685 (N_13685,N_10074,N_12496);
or U13686 (N_13686,N_9951,N_11282);
nand U13687 (N_13687,N_10700,N_10858);
or U13688 (N_13688,N_12377,N_9711);
and U13689 (N_13689,N_10146,N_9608);
nor U13690 (N_13690,N_9407,N_11356);
or U13691 (N_13691,N_12306,N_10722);
nand U13692 (N_13692,N_11991,N_9747);
xnor U13693 (N_13693,N_10933,N_10288);
or U13694 (N_13694,N_10914,N_11067);
nand U13695 (N_13695,N_10704,N_10413);
xnor U13696 (N_13696,N_11776,N_9745);
nand U13697 (N_13697,N_11016,N_12001);
xnor U13698 (N_13698,N_9962,N_12177);
and U13699 (N_13699,N_10031,N_9544);
and U13700 (N_13700,N_10204,N_11061);
or U13701 (N_13701,N_10476,N_11681);
or U13702 (N_13702,N_10901,N_10667);
nor U13703 (N_13703,N_9627,N_10005);
nor U13704 (N_13704,N_12226,N_10322);
and U13705 (N_13705,N_9875,N_11338);
nor U13706 (N_13706,N_11121,N_10274);
xor U13707 (N_13707,N_12038,N_11586);
and U13708 (N_13708,N_12140,N_12480);
nor U13709 (N_13709,N_11127,N_11965);
nand U13710 (N_13710,N_10958,N_12247);
or U13711 (N_13711,N_12241,N_9868);
xor U13712 (N_13712,N_12299,N_11076);
nor U13713 (N_13713,N_11984,N_11599);
nand U13714 (N_13714,N_11024,N_11089);
nor U13715 (N_13715,N_10941,N_10940);
nor U13716 (N_13716,N_12186,N_11538);
or U13717 (N_13717,N_10022,N_10565);
xor U13718 (N_13718,N_11243,N_10645);
nor U13719 (N_13719,N_11218,N_11361);
or U13720 (N_13720,N_10873,N_11014);
and U13721 (N_13721,N_9486,N_10028);
or U13722 (N_13722,N_11152,N_11502);
and U13723 (N_13723,N_11763,N_11782);
nand U13724 (N_13724,N_11452,N_9838);
or U13725 (N_13725,N_11480,N_10671);
and U13726 (N_13726,N_9587,N_10503);
xnor U13727 (N_13727,N_9628,N_9691);
or U13728 (N_13728,N_11183,N_11374);
and U13729 (N_13729,N_10701,N_10162);
and U13730 (N_13730,N_12418,N_9771);
nor U13731 (N_13731,N_11904,N_11410);
or U13732 (N_13732,N_10802,N_9889);
or U13733 (N_13733,N_9728,N_11433);
nand U13734 (N_13734,N_10842,N_10618);
nand U13735 (N_13735,N_9537,N_11213);
nor U13736 (N_13736,N_11670,N_10994);
nand U13737 (N_13737,N_10967,N_11810);
nor U13738 (N_13738,N_12440,N_11725);
nand U13739 (N_13739,N_11941,N_10761);
xnor U13740 (N_13740,N_12277,N_10639);
and U13741 (N_13741,N_10732,N_9680);
and U13742 (N_13742,N_10225,N_12266);
or U13743 (N_13743,N_12119,N_12192);
nor U13744 (N_13744,N_11360,N_10291);
or U13745 (N_13745,N_10553,N_9648);
and U13746 (N_13746,N_12436,N_9531);
and U13747 (N_13747,N_10284,N_12034);
nor U13748 (N_13748,N_9467,N_11159);
nand U13749 (N_13749,N_10432,N_10355);
nand U13750 (N_13750,N_10818,N_10126);
and U13751 (N_13751,N_9512,N_11236);
and U13752 (N_13752,N_12117,N_9540);
nor U13753 (N_13753,N_11940,N_10398);
nor U13754 (N_13754,N_10920,N_10263);
xor U13755 (N_13755,N_10916,N_12236);
and U13756 (N_13756,N_11500,N_11008);
and U13757 (N_13757,N_10009,N_9955);
xor U13758 (N_13758,N_11004,N_11534);
and U13759 (N_13759,N_11258,N_11510);
xor U13760 (N_13760,N_11722,N_10098);
nor U13761 (N_13761,N_10760,N_11680);
nand U13762 (N_13762,N_9818,N_10118);
and U13763 (N_13763,N_12050,N_12409);
nor U13764 (N_13764,N_12370,N_11735);
or U13765 (N_13765,N_10570,N_11906);
nand U13766 (N_13766,N_10453,N_10402);
nand U13767 (N_13767,N_12020,N_11122);
nand U13768 (N_13768,N_12326,N_10444);
and U13769 (N_13769,N_11817,N_10346);
and U13770 (N_13770,N_9950,N_12012);
nand U13771 (N_13771,N_10990,N_12312);
nand U13772 (N_13772,N_10472,N_11288);
or U13773 (N_13773,N_9933,N_10153);
nor U13774 (N_13774,N_12411,N_10378);
xor U13775 (N_13775,N_9396,N_10102);
or U13776 (N_13776,N_9982,N_10524);
or U13777 (N_13777,N_10356,N_10535);
and U13778 (N_13778,N_11899,N_10208);
and U13779 (N_13779,N_12055,N_11915);
or U13780 (N_13780,N_11970,N_10515);
xor U13781 (N_13781,N_12217,N_12136);
and U13782 (N_13782,N_10995,N_12108);
and U13783 (N_13783,N_11865,N_10276);
or U13784 (N_13784,N_11922,N_10048);
or U13785 (N_13785,N_10881,N_9501);
nand U13786 (N_13786,N_11058,N_11326);
nand U13787 (N_13787,N_12172,N_9820);
or U13788 (N_13788,N_10107,N_9503);
nor U13789 (N_13789,N_10015,N_11277);
or U13790 (N_13790,N_11431,N_11969);
and U13791 (N_13791,N_11484,N_11293);
nor U13792 (N_13792,N_11148,N_11886);
nand U13793 (N_13793,N_10141,N_9602);
nor U13794 (N_13794,N_10257,N_11815);
and U13795 (N_13795,N_10470,N_12374);
or U13796 (N_13796,N_12002,N_9456);
nand U13797 (N_13797,N_10012,N_9891);
or U13798 (N_13798,N_11568,N_9438);
nor U13799 (N_13799,N_12433,N_11859);
or U13800 (N_13800,N_10982,N_12130);
or U13801 (N_13801,N_12176,N_10929);
nand U13802 (N_13802,N_11084,N_11385);
and U13803 (N_13803,N_11113,N_11349);
and U13804 (N_13804,N_9788,N_11352);
and U13805 (N_13805,N_10674,N_10383);
and U13806 (N_13806,N_10491,N_10152);
and U13807 (N_13807,N_11853,N_9642);
nor U13808 (N_13808,N_11451,N_10317);
and U13809 (N_13809,N_11939,N_11376);
xnor U13810 (N_13810,N_11994,N_12471);
or U13811 (N_13811,N_11357,N_11920);
nor U13812 (N_13812,N_9803,N_12203);
nor U13813 (N_13813,N_11702,N_10407);
and U13814 (N_13814,N_12333,N_12196);
nor U13815 (N_13815,N_9748,N_10198);
nor U13816 (N_13816,N_10295,N_9380);
or U13817 (N_13817,N_9611,N_10496);
nor U13818 (N_13818,N_12005,N_10686);
or U13819 (N_13819,N_10427,N_9760);
xnor U13820 (N_13820,N_11858,N_10041);
or U13821 (N_13821,N_9989,N_10726);
and U13822 (N_13822,N_9681,N_10777);
or U13823 (N_13823,N_11666,N_11861);
nor U13824 (N_13824,N_10200,N_10694);
or U13825 (N_13825,N_11603,N_12220);
or U13826 (N_13826,N_11485,N_10977);
nand U13827 (N_13827,N_11877,N_10147);
nor U13828 (N_13828,N_11546,N_9624);
nand U13829 (N_13829,N_12037,N_12446);
nor U13830 (N_13830,N_10974,N_10474);
or U13831 (N_13831,N_11678,N_11856);
or U13832 (N_13832,N_11306,N_10626);
or U13833 (N_13833,N_10016,N_10329);
and U13834 (N_13834,N_11402,N_10824);
xnor U13835 (N_13835,N_11966,N_9856);
nand U13836 (N_13836,N_11867,N_9508);
nor U13837 (N_13837,N_11873,N_9619);
and U13838 (N_13838,N_9874,N_9595);
or U13839 (N_13839,N_9949,N_10237);
nor U13840 (N_13840,N_12391,N_9427);
nand U13841 (N_13841,N_12017,N_10171);
or U13842 (N_13842,N_9443,N_10859);
nor U13843 (N_13843,N_12421,N_12430);
nor U13844 (N_13844,N_9490,N_9696);
nand U13845 (N_13845,N_10705,N_11643);
nand U13846 (N_13846,N_11708,N_9952);
nor U13847 (N_13847,N_9939,N_10845);
or U13848 (N_13848,N_12248,N_9924);
and U13849 (N_13849,N_11521,N_11171);
or U13850 (N_13850,N_10359,N_11368);
or U13851 (N_13851,N_11497,N_11247);
or U13852 (N_13852,N_12288,N_11986);
or U13853 (N_13853,N_9910,N_11176);
or U13854 (N_13854,N_10058,N_10128);
and U13855 (N_13855,N_11437,N_9572);
xnor U13856 (N_13856,N_9676,N_11206);
nor U13857 (N_13857,N_12362,N_10483);
nor U13858 (N_13858,N_11639,N_10371);
nand U13859 (N_13859,N_12182,N_11262);
xnor U13860 (N_13860,N_10670,N_10044);
xor U13861 (N_13861,N_11580,N_11593);
nor U13862 (N_13862,N_12239,N_11571);
nor U13863 (N_13863,N_12225,N_11081);
xor U13864 (N_13864,N_9630,N_9405);
and U13865 (N_13865,N_11046,N_11821);
nor U13866 (N_13866,N_11251,N_10055);
nor U13867 (N_13867,N_10482,N_11462);
and U13868 (N_13868,N_10947,N_9601);
xor U13869 (N_13869,N_11160,N_9607);
xnor U13870 (N_13870,N_10302,N_10447);
nand U13871 (N_13871,N_11119,N_9713);
and U13872 (N_13872,N_10890,N_11990);
xnor U13873 (N_13873,N_11125,N_9584);
nand U13874 (N_13874,N_11467,N_10928);
nor U13875 (N_13875,N_10105,N_10121);
and U13876 (N_13876,N_11128,N_12041);
nor U13877 (N_13877,N_12361,N_11912);
and U13878 (N_13878,N_10733,N_11694);
and U13879 (N_13879,N_11641,N_11893);
and U13880 (N_13880,N_9899,N_10020);
or U13881 (N_13881,N_11664,N_9391);
nand U13882 (N_13882,N_9737,N_12497);
nor U13883 (N_13883,N_11589,N_10308);
nand U13884 (N_13884,N_12267,N_10174);
nor U13885 (N_13885,N_12138,N_11375);
or U13886 (N_13886,N_11105,N_10883);
or U13887 (N_13887,N_12185,N_10819);
nand U13888 (N_13888,N_10266,N_12056);
nor U13889 (N_13889,N_10993,N_9482);
and U13890 (N_13890,N_11281,N_9968);
or U13891 (N_13891,N_10578,N_11138);
or U13892 (N_13892,N_11754,N_10321);
nand U13893 (N_13893,N_9645,N_11558);
nor U13894 (N_13894,N_11329,N_10556);
nor U13895 (N_13895,N_9996,N_11957);
nand U13896 (N_13896,N_9484,N_9605);
and U13897 (N_13897,N_10728,N_11047);
nor U13898 (N_13898,N_12491,N_11529);
nor U13899 (N_13899,N_10880,N_12114);
and U13900 (N_13900,N_11116,N_10755);
or U13901 (N_13901,N_9708,N_11229);
and U13902 (N_13902,N_10490,N_11098);
or U13903 (N_13903,N_10937,N_10179);
nor U13904 (N_13904,N_10340,N_9766);
and U13905 (N_13905,N_11239,N_12367);
nor U13906 (N_13906,N_10348,N_10641);
nand U13907 (N_13907,N_11911,N_10964);
nor U13908 (N_13908,N_9757,N_10562);
and U13909 (N_13909,N_10160,N_11604);
nor U13910 (N_13910,N_12382,N_10426);
nand U13911 (N_13911,N_11659,N_10306);
nand U13912 (N_13912,N_12021,N_11547);
nor U13913 (N_13913,N_10589,N_11636);
nand U13914 (N_13914,N_11960,N_12484);
or U13915 (N_13915,N_10668,N_10899);
or U13916 (N_13916,N_11846,N_11894);
nand U13917 (N_13917,N_10349,N_11365);
nor U13918 (N_13918,N_11674,N_9785);
xor U13919 (N_13919,N_11300,N_9578);
xor U13920 (N_13920,N_11466,N_12201);
and U13921 (N_13921,N_10803,N_11123);
nand U13922 (N_13922,N_11635,N_10065);
nor U13923 (N_13923,N_9953,N_11042);
nor U13924 (N_13924,N_12284,N_10357);
and U13925 (N_13925,N_11715,N_12013);
or U13926 (N_13926,N_10262,N_11082);
or U13927 (N_13927,N_11563,N_11905);
or U13928 (N_13928,N_11918,N_10826);
xor U13929 (N_13929,N_11015,N_11482);
or U13930 (N_13930,N_11724,N_12457);
or U13931 (N_13931,N_9911,N_11195);
and U13932 (N_13932,N_9742,N_10696);
xnor U13933 (N_13933,N_9769,N_9826);
nor U13934 (N_13934,N_10297,N_9640);
and U13935 (N_13935,N_12438,N_9990);
xnor U13936 (N_13936,N_12255,N_11656);
xnor U13937 (N_13937,N_10078,N_10300);
or U13938 (N_13938,N_9462,N_11168);
nand U13939 (N_13939,N_12035,N_12200);
and U13940 (N_13940,N_9570,N_11491);
and U13941 (N_13941,N_12156,N_10150);
or U13942 (N_13942,N_11714,N_11931);
xor U13943 (N_13943,N_9435,N_12188);
xor U13944 (N_13944,N_12476,N_12425);
or U13945 (N_13945,N_11395,N_10663);
or U13946 (N_13946,N_9496,N_10936);
or U13947 (N_13947,N_9964,N_10197);
nand U13948 (N_13948,N_11710,N_10811);
and U13949 (N_13949,N_11200,N_10837);
or U13950 (N_13950,N_9677,N_10084);
nand U13951 (N_13951,N_11074,N_9672);
and U13952 (N_13952,N_12351,N_9884);
nand U13953 (N_13953,N_10458,N_9844);
or U13954 (N_13954,N_9418,N_11879);
xnor U13955 (N_13955,N_10891,N_9598);
or U13956 (N_13956,N_10534,N_9661);
nor U13957 (N_13957,N_11393,N_11286);
nand U13958 (N_13958,N_10724,N_9600);
or U13959 (N_13959,N_11197,N_11600);
nand U13960 (N_13960,N_9800,N_11205);
xor U13961 (N_13961,N_10215,N_12081);
nand U13962 (N_13962,N_10514,N_10138);
nor U13963 (N_13963,N_10224,N_10066);
nor U13964 (N_13964,N_9402,N_10902);
nand U13965 (N_13965,N_10443,N_9787);
or U13966 (N_13966,N_12324,N_9475);
nor U13967 (N_13967,N_11290,N_12116);
nand U13968 (N_13968,N_12357,N_10294);
and U13969 (N_13969,N_10464,N_10988);
xnor U13970 (N_13970,N_11315,N_9915);
xor U13971 (N_13971,N_10528,N_11188);
xnor U13972 (N_13972,N_9594,N_10836);
and U13973 (N_13973,N_11245,N_10059);
and U13974 (N_13974,N_10218,N_11210);
nor U13975 (N_13975,N_12392,N_12132);
and U13976 (N_13976,N_10730,N_11883);
nor U13977 (N_13977,N_11440,N_10593);
xnor U13978 (N_13978,N_9805,N_10182);
or U13979 (N_13979,N_10038,N_11805);
nor U13980 (N_13980,N_9830,N_11455);
or U13981 (N_13981,N_10269,N_10989);
nor U13982 (N_13982,N_12363,N_9967);
nand U13983 (N_13983,N_11102,N_11054);
or U13984 (N_13984,N_10220,N_11027);
nand U13985 (N_13985,N_9914,N_10364);
nand U13986 (N_13986,N_12099,N_9660);
nand U13987 (N_13987,N_12089,N_12450);
or U13988 (N_13988,N_10682,N_9752);
and U13989 (N_13989,N_12420,N_12348);
nor U13990 (N_13990,N_10685,N_11314);
or U13991 (N_13991,N_11692,N_11851);
or U13992 (N_13992,N_11317,N_11526);
and U13993 (N_13993,N_11050,N_10250);
nand U13994 (N_13994,N_9976,N_11855);
nor U13995 (N_13995,N_11118,N_10610);
or U13996 (N_13996,N_12042,N_9859);
nand U13997 (N_13997,N_10844,N_9997);
nor U13998 (N_13998,N_11552,N_11590);
nor U13999 (N_13999,N_10104,N_10228);
or U14000 (N_14000,N_10975,N_11841);
and U14001 (N_14001,N_9631,N_11011);
or U14002 (N_14002,N_11594,N_9741);
or U14003 (N_14003,N_11285,N_10460);
nor U14004 (N_14004,N_9902,N_10939);
and U14005 (N_14005,N_10625,N_9840);
nand U14006 (N_14006,N_12251,N_11985);
or U14007 (N_14007,N_11208,N_9934);
nand U14008 (N_14008,N_9547,N_11325);
and U14009 (N_14009,N_12296,N_9411);
nand U14010 (N_14010,N_10542,N_9571);
nand U14011 (N_14011,N_11063,N_11273);
nand U14012 (N_14012,N_12399,N_9937);
xor U14013 (N_14013,N_12088,N_11174);
nand U14014 (N_14014,N_9381,N_10176);
nor U14015 (N_14015,N_10765,N_12230);
nor U14016 (N_14016,N_9904,N_9397);
nor U14017 (N_14017,N_12093,N_10017);
nand U14018 (N_14018,N_12106,N_10609);
or U14019 (N_14019,N_11874,N_11548);
or U14020 (N_14020,N_12129,N_10750);
nor U14021 (N_14021,N_11371,N_12221);
or U14022 (N_14022,N_9580,N_11367);
and U14023 (N_14023,N_12112,N_10808);
or U14024 (N_14024,N_11025,N_11993);
xor U14025 (N_14025,N_12460,N_12290);
nand U14026 (N_14026,N_9507,N_10948);
or U14027 (N_14027,N_12323,N_10927);
nor U14028 (N_14028,N_11069,N_11447);
and U14029 (N_14029,N_11483,N_11345);
or U14030 (N_14030,N_10478,N_10847);
and U14031 (N_14031,N_11453,N_11312);
and U14032 (N_14032,N_10362,N_9637);
xor U14033 (N_14033,N_11573,N_12074);
nand U14034 (N_14034,N_11687,N_10199);
and U14035 (N_14035,N_10991,N_10627);
xnor U14036 (N_14036,N_9596,N_10395);
nand U14037 (N_14037,N_9798,N_10073);
and U14038 (N_14038,N_9945,N_11373);
nand U14039 (N_14039,N_9980,N_12162);
nor U14040 (N_14040,N_11773,N_9869);
or U14041 (N_14041,N_9659,N_10711);
nor U14042 (N_14042,N_11268,N_10293);
and U14043 (N_14043,N_10539,N_11818);
nand U14044 (N_14044,N_11347,N_10797);
nor U14045 (N_14045,N_10548,N_9709);
nand U14046 (N_14046,N_11378,N_11199);
or U14047 (N_14047,N_12139,N_10040);
and U14048 (N_14048,N_10745,N_11887);
and U14049 (N_14049,N_11503,N_9701);
or U14050 (N_14050,N_11577,N_9783);
or U14051 (N_14051,N_10852,N_12204);
nor U14052 (N_14052,N_12090,N_11109);
xor U14053 (N_14053,N_10905,N_9425);
or U14054 (N_14054,N_11299,N_11576);
nor U14055 (N_14055,N_12297,N_9510);
or U14056 (N_14056,N_9495,N_11209);
and U14057 (N_14057,N_11709,N_10673);
nand U14058 (N_14058,N_9848,N_12064);
or U14059 (N_14059,N_11498,N_10004);
nor U14060 (N_14060,N_10934,N_10915);
xor U14061 (N_14061,N_10091,N_10669);
nand U14062 (N_14062,N_11703,N_10484);
nand U14063 (N_14063,N_11455,N_9406);
and U14064 (N_14064,N_11196,N_11182);
and U14065 (N_14065,N_11701,N_10121);
and U14066 (N_14066,N_11922,N_11282);
nor U14067 (N_14067,N_11087,N_12375);
or U14068 (N_14068,N_12261,N_11174);
nor U14069 (N_14069,N_11398,N_9641);
nor U14070 (N_14070,N_9773,N_12248);
nor U14071 (N_14071,N_11578,N_11244);
xor U14072 (N_14072,N_9618,N_12132);
nor U14073 (N_14073,N_11607,N_11229);
nor U14074 (N_14074,N_11861,N_10613);
or U14075 (N_14075,N_10118,N_11657);
nor U14076 (N_14076,N_11521,N_11430);
and U14077 (N_14077,N_11503,N_12252);
nor U14078 (N_14078,N_12041,N_9757);
or U14079 (N_14079,N_11614,N_11894);
or U14080 (N_14080,N_10247,N_11849);
or U14081 (N_14081,N_10955,N_11764);
and U14082 (N_14082,N_10713,N_10853);
nor U14083 (N_14083,N_11181,N_12138);
nand U14084 (N_14084,N_9395,N_11154);
or U14085 (N_14085,N_10299,N_12467);
or U14086 (N_14086,N_10430,N_10155);
nor U14087 (N_14087,N_9850,N_10588);
xnor U14088 (N_14088,N_10407,N_12073);
and U14089 (N_14089,N_12455,N_11310);
nor U14090 (N_14090,N_9629,N_11246);
or U14091 (N_14091,N_9669,N_12161);
and U14092 (N_14092,N_11230,N_11462);
or U14093 (N_14093,N_11624,N_11224);
or U14094 (N_14094,N_10718,N_11168);
nor U14095 (N_14095,N_10587,N_11922);
xor U14096 (N_14096,N_10827,N_10337);
or U14097 (N_14097,N_10401,N_11573);
xor U14098 (N_14098,N_11875,N_9739);
or U14099 (N_14099,N_11868,N_10081);
or U14100 (N_14100,N_12423,N_11345);
nor U14101 (N_14101,N_11593,N_11929);
nand U14102 (N_14102,N_10624,N_12215);
nand U14103 (N_14103,N_9439,N_11048);
xor U14104 (N_14104,N_10386,N_10625);
nor U14105 (N_14105,N_11671,N_9999);
xnor U14106 (N_14106,N_12249,N_9754);
nand U14107 (N_14107,N_10179,N_11774);
or U14108 (N_14108,N_10310,N_10831);
nor U14109 (N_14109,N_11544,N_9404);
xnor U14110 (N_14110,N_11172,N_11421);
nand U14111 (N_14111,N_9450,N_11372);
or U14112 (N_14112,N_11541,N_10150);
nand U14113 (N_14113,N_10527,N_10482);
nand U14114 (N_14114,N_11334,N_10263);
nor U14115 (N_14115,N_11319,N_12109);
and U14116 (N_14116,N_10434,N_9955);
nand U14117 (N_14117,N_9756,N_9629);
or U14118 (N_14118,N_9684,N_9606);
and U14119 (N_14119,N_11045,N_11503);
xnor U14120 (N_14120,N_9695,N_11073);
nor U14121 (N_14121,N_10685,N_9596);
and U14122 (N_14122,N_10940,N_12172);
nand U14123 (N_14123,N_10920,N_11429);
nor U14124 (N_14124,N_9427,N_11606);
and U14125 (N_14125,N_12119,N_10127);
nand U14126 (N_14126,N_11729,N_11322);
and U14127 (N_14127,N_10926,N_9823);
or U14128 (N_14128,N_10946,N_10159);
xnor U14129 (N_14129,N_11059,N_12003);
xnor U14130 (N_14130,N_12012,N_9421);
nor U14131 (N_14131,N_9720,N_9942);
or U14132 (N_14132,N_11252,N_10819);
nand U14133 (N_14133,N_9847,N_9780);
nand U14134 (N_14134,N_10969,N_11860);
nor U14135 (N_14135,N_11107,N_11371);
nor U14136 (N_14136,N_10776,N_11029);
or U14137 (N_14137,N_11035,N_11511);
nor U14138 (N_14138,N_10333,N_11510);
xnor U14139 (N_14139,N_12178,N_9549);
or U14140 (N_14140,N_11780,N_12233);
and U14141 (N_14141,N_11085,N_9995);
or U14142 (N_14142,N_12165,N_11727);
and U14143 (N_14143,N_11744,N_12069);
xnor U14144 (N_14144,N_11186,N_11685);
nor U14145 (N_14145,N_12487,N_9757);
or U14146 (N_14146,N_10265,N_9602);
and U14147 (N_14147,N_9826,N_11954);
nand U14148 (N_14148,N_11211,N_12185);
or U14149 (N_14149,N_10106,N_10932);
or U14150 (N_14150,N_12487,N_9717);
xnor U14151 (N_14151,N_10412,N_10515);
and U14152 (N_14152,N_9713,N_11795);
or U14153 (N_14153,N_11006,N_12203);
or U14154 (N_14154,N_9388,N_9409);
xor U14155 (N_14155,N_10341,N_11756);
nor U14156 (N_14156,N_11378,N_10994);
nand U14157 (N_14157,N_11244,N_12395);
nor U14158 (N_14158,N_11673,N_11848);
nor U14159 (N_14159,N_10710,N_9787);
and U14160 (N_14160,N_10202,N_12475);
and U14161 (N_14161,N_11315,N_11632);
and U14162 (N_14162,N_11442,N_9524);
nand U14163 (N_14163,N_10025,N_12055);
or U14164 (N_14164,N_10347,N_10882);
and U14165 (N_14165,N_10143,N_12366);
or U14166 (N_14166,N_9569,N_11165);
and U14167 (N_14167,N_11059,N_9622);
nor U14168 (N_14168,N_10269,N_11762);
nor U14169 (N_14169,N_11776,N_10165);
or U14170 (N_14170,N_11736,N_10072);
and U14171 (N_14171,N_9832,N_12234);
xnor U14172 (N_14172,N_12134,N_9381);
or U14173 (N_14173,N_10728,N_11757);
nor U14174 (N_14174,N_11455,N_11858);
nor U14175 (N_14175,N_10839,N_10389);
nand U14176 (N_14176,N_10369,N_10730);
or U14177 (N_14177,N_11471,N_11542);
and U14178 (N_14178,N_9684,N_9740);
and U14179 (N_14179,N_9853,N_11155);
nand U14180 (N_14180,N_9525,N_12100);
or U14181 (N_14181,N_12136,N_9531);
nor U14182 (N_14182,N_9452,N_9539);
nand U14183 (N_14183,N_10491,N_12243);
and U14184 (N_14184,N_10598,N_12384);
xnor U14185 (N_14185,N_12241,N_10452);
nand U14186 (N_14186,N_9597,N_11846);
nor U14187 (N_14187,N_11205,N_11923);
nor U14188 (N_14188,N_11481,N_11593);
nor U14189 (N_14189,N_12484,N_10669);
nor U14190 (N_14190,N_9492,N_10663);
nand U14191 (N_14191,N_10745,N_11696);
nor U14192 (N_14192,N_9425,N_9395);
nand U14193 (N_14193,N_11378,N_11837);
and U14194 (N_14194,N_9395,N_10424);
or U14195 (N_14195,N_11316,N_10766);
and U14196 (N_14196,N_12020,N_10907);
or U14197 (N_14197,N_9832,N_9453);
or U14198 (N_14198,N_10060,N_12011);
nor U14199 (N_14199,N_10103,N_9542);
and U14200 (N_14200,N_10197,N_10801);
nand U14201 (N_14201,N_10894,N_10325);
and U14202 (N_14202,N_10465,N_10678);
nor U14203 (N_14203,N_11645,N_11276);
xor U14204 (N_14204,N_9433,N_11325);
nor U14205 (N_14205,N_10313,N_10838);
nand U14206 (N_14206,N_10839,N_10929);
or U14207 (N_14207,N_11053,N_12036);
or U14208 (N_14208,N_11646,N_12345);
nand U14209 (N_14209,N_11779,N_11196);
or U14210 (N_14210,N_12208,N_10326);
and U14211 (N_14211,N_10384,N_9680);
xor U14212 (N_14212,N_12420,N_11524);
and U14213 (N_14213,N_12370,N_10311);
xnor U14214 (N_14214,N_11399,N_11729);
and U14215 (N_14215,N_12346,N_11372);
and U14216 (N_14216,N_11205,N_12066);
and U14217 (N_14217,N_10830,N_12349);
or U14218 (N_14218,N_11536,N_11417);
or U14219 (N_14219,N_12085,N_11172);
or U14220 (N_14220,N_11609,N_11058);
and U14221 (N_14221,N_10427,N_12055);
or U14222 (N_14222,N_9900,N_9957);
and U14223 (N_14223,N_12075,N_9734);
nand U14224 (N_14224,N_11528,N_9929);
nor U14225 (N_14225,N_10063,N_10395);
or U14226 (N_14226,N_12245,N_9585);
and U14227 (N_14227,N_11961,N_10220);
xnor U14228 (N_14228,N_10160,N_10920);
nor U14229 (N_14229,N_11621,N_9788);
and U14230 (N_14230,N_10563,N_10043);
or U14231 (N_14231,N_11286,N_12430);
nor U14232 (N_14232,N_10087,N_9477);
and U14233 (N_14233,N_10076,N_10192);
or U14234 (N_14234,N_10392,N_9894);
and U14235 (N_14235,N_9934,N_11158);
nor U14236 (N_14236,N_10473,N_11554);
nor U14237 (N_14237,N_9835,N_10972);
xnor U14238 (N_14238,N_11157,N_9899);
or U14239 (N_14239,N_11223,N_11750);
or U14240 (N_14240,N_9691,N_12288);
or U14241 (N_14241,N_11535,N_11746);
and U14242 (N_14242,N_10380,N_10664);
xnor U14243 (N_14243,N_11484,N_12327);
nand U14244 (N_14244,N_11575,N_10604);
nand U14245 (N_14245,N_12302,N_12238);
and U14246 (N_14246,N_10544,N_9886);
nor U14247 (N_14247,N_12108,N_10475);
and U14248 (N_14248,N_9764,N_9595);
nand U14249 (N_14249,N_11926,N_11595);
nor U14250 (N_14250,N_11112,N_10658);
xor U14251 (N_14251,N_11927,N_10344);
nand U14252 (N_14252,N_9971,N_9868);
nand U14253 (N_14253,N_12182,N_12237);
and U14254 (N_14254,N_11843,N_9450);
or U14255 (N_14255,N_10236,N_10054);
and U14256 (N_14256,N_11028,N_11636);
nand U14257 (N_14257,N_10080,N_10428);
or U14258 (N_14258,N_10096,N_9456);
or U14259 (N_14259,N_9702,N_11253);
nand U14260 (N_14260,N_10751,N_9780);
and U14261 (N_14261,N_11333,N_12160);
xnor U14262 (N_14262,N_10687,N_10141);
xor U14263 (N_14263,N_9457,N_9591);
or U14264 (N_14264,N_11676,N_11768);
nor U14265 (N_14265,N_10785,N_11192);
and U14266 (N_14266,N_11121,N_10385);
nor U14267 (N_14267,N_11437,N_11124);
and U14268 (N_14268,N_10692,N_12216);
xnor U14269 (N_14269,N_10920,N_10284);
nor U14270 (N_14270,N_10775,N_10169);
or U14271 (N_14271,N_12145,N_10380);
or U14272 (N_14272,N_12028,N_10871);
xor U14273 (N_14273,N_10265,N_10501);
or U14274 (N_14274,N_10210,N_11904);
nor U14275 (N_14275,N_11848,N_9783);
nor U14276 (N_14276,N_10329,N_9996);
nor U14277 (N_14277,N_12378,N_11619);
nand U14278 (N_14278,N_10999,N_9986);
nand U14279 (N_14279,N_11998,N_12166);
and U14280 (N_14280,N_10412,N_11299);
nand U14281 (N_14281,N_9821,N_9501);
or U14282 (N_14282,N_10732,N_10963);
and U14283 (N_14283,N_12221,N_10587);
or U14284 (N_14284,N_12280,N_11154);
nor U14285 (N_14285,N_11424,N_11562);
nor U14286 (N_14286,N_12091,N_11092);
nor U14287 (N_14287,N_9397,N_11607);
and U14288 (N_14288,N_9891,N_11997);
nand U14289 (N_14289,N_9899,N_9980);
and U14290 (N_14290,N_11914,N_11532);
and U14291 (N_14291,N_11740,N_9929);
nor U14292 (N_14292,N_12262,N_9829);
and U14293 (N_14293,N_10386,N_11979);
nor U14294 (N_14294,N_10407,N_9787);
or U14295 (N_14295,N_10760,N_11628);
xnor U14296 (N_14296,N_11498,N_9696);
nand U14297 (N_14297,N_11296,N_10202);
nand U14298 (N_14298,N_12096,N_11786);
xnor U14299 (N_14299,N_10835,N_10256);
nand U14300 (N_14300,N_10617,N_12345);
and U14301 (N_14301,N_12048,N_11320);
nor U14302 (N_14302,N_10485,N_11285);
nand U14303 (N_14303,N_12329,N_11778);
nor U14304 (N_14304,N_10638,N_9565);
nor U14305 (N_14305,N_11869,N_9951);
and U14306 (N_14306,N_10192,N_9644);
and U14307 (N_14307,N_9844,N_11219);
nand U14308 (N_14308,N_10169,N_10570);
nor U14309 (N_14309,N_10330,N_12078);
xor U14310 (N_14310,N_11181,N_12341);
or U14311 (N_14311,N_10400,N_10973);
nand U14312 (N_14312,N_10415,N_12473);
nor U14313 (N_14313,N_9765,N_10593);
or U14314 (N_14314,N_10416,N_10355);
and U14315 (N_14315,N_9742,N_10108);
and U14316 (N_14316,N_11041,N_12106);
and U14317 (N_14317,N_11730,N_10060);
nand U14318 (N_14318,N_9632,N_10220);
and U14319 (N_14319,N_12288,N_10988);
and U14320 (N_14320,N_11349,N_11558);
or U14321 (N_14321,N_9518,N_11058);
nand U14322 (N_14322,N_11517,N_10096);
nor U14323 (N_14323,N_9423,N_11212);
and U14324 (N_14324,N_12084,N_10013);
nand U14325 (N_14325,N_12118,N_11863);
nor U14326 (N_14326,N_12327,N_12253);
and U14327 (N_14327,N_11736,N_11035);
xor U14328 (N_14328,N_11407,N_10754);
or U14329 (N_14329,N_12471,N_10680);
or U14330 (N_14330,N_11834,N_11790);
nor U14331 (N_14331,N_9590,N_10946);
and U14332 (N_14332,N_10734,N_11926);
nor U14333 (N_14333,N_12473,N_11806);
xor U14334 (N_14334,N_10132,N_11336);
nor U14335 (N_14335,N_10188,N_10400);
xor U14336 (N_14336,N_11363,N_9436);
nor U14337 (N_14337,N_11413,N_10178);
or U14338 (N_14338,N_10111,N_10409);
or U14339 (N_14339,N_12496,N_11593);
and U14340 (N_14340,N_11149,N_12273);
and U14341 (N_14341,N_10173,N_9647);
and U14342 (N_14342,N_12277,N_9603);
or U14343 (N_14343,N_12117,N_12113);
or U14344 (N_14344,N_11848,N_11113);
nor U14345 (N_14345,N_11283,N_10934);
or U14346 (N_14346,N_10435,N_11409);
and U14347 (N_14347,N_11247,N_10033);
nand U14348 (N_14348,N_12195,N_12433);
or U14349 (N_14349,N_9907,N_12170);
nand U14350 (N_14350,N_10309,N_9968);
nand U14351 (N_14351,N_10396,N_10633);
or U14352 (N_14352,N_10914,N_9610);
xor U14353 (N_14353,N_11689,N_10981);
nor U14354 (N_14354,N_9644,N_9948);
nor U14355 (N_14355,N_10580,N_12392);
nor U14356 (N_14356,N_10672,N_10659);
nand U14357 (N_14357,N_9941,N_10959);
or U14358 (N_14358,N_11909,N_10088);
nor U14359 (N_14359,N_9967,N_11359);
or U14360 (N_14360,N_10237,N_10563);
or U14361 (N_14361,N_10387,N_9440);
or U14362 (N_14362,N_10580,N_11813);
nor U14363 (N_14363,N_11074,N_11838);
nand U14364 (N_14364,N_9450,N_11506);
nand U14365 (N_14365,N_12347,N_10607);
nand U14366 (N_14366,N_9710,N_11919);
nand U14367 (N_14367,N_10895,N_9760);
nor U14368 (N_14368,N_10993,N_12156);
and U14369 (N_14369,N_12171,N_10951);
or U14370 (N_14370,N_11702,N_12399);
and U14371 (N_14371,N_11095,N_12214);
xor U14372 (N_14372,N_11944,N_10408);
and U14373 (N_14373,N_9773,N_11103);
or U14374 (N_14374,N_10532,N_12419);
nand U14375 (N_14375,N_10108,N_11052);
nor U14376 (N_14376,N_10466,N_11225);
or U14377 (N_14377,N_12032,N_10472);
nor U14378 (N_14378,N_10467,N_12269);
and U14379 (N_14379,N_11851,N_9482);
nand U14380 (N_14380,N_10394,N_9656);
nand U14381 (N_14381,N_10653,N_9392);
or U14382 (N_14382,N_11421,N_11451);
nor U14383 (N_14383,N_12272,N_11400);
nor U14384 (N_14384,N_9811,N_9676);
nand U14385 (N_14385,N_11093,N_12169);
nand U14386 (N_14386,N_12071,N_10950);
and U14387 (N_14387,N_11341,N_10571);
and U14388 (N_14388,N_10038,N_11473);
xnor U14389 (N_14389,N_9868,N_10789);
and U14390 (N_14390,N_11484,N_9812);
xor U14391 (N_14391,N_10937,N_12385);
xnor U14392 (N_14392,N_9869,N_11941);
nor U14393 (N_14393,N_12433,N_12396);
nand U14394 (N_14394,N_11554,N_11769);
or U14395 (N_14395,N_11107,N_9393);
nand U14396 (N_14396,N_12206,N_11844);
nand U14397 (N_14397,N_11926,N_10267);
and U14398 (N_14398,N_11788,N_11754);
nor U14399 (N_14399,N_11637,N_12025);
and U14400 (N_14400,N_11329,N_10285);
or U14401 (N_14401,N_9404,N_11007);
and U14402 (N_14402,N_10233,N_10894);
and U14403 (N_14403,N_9466,N_10247);
nand U14404 (N_14404,N_11878,N_9498);
xnor U14405 (N_14405,N_11025,N_10935);
or U14406 (N_14406,N_12227,N_10962);
and U14407 (N_14407,N_11667,N_11401);
nand U14408 (N_14408,N_11609,N_11381);
nor U14409 (N_14409,N_11232,N_11853);
nand U14410 (N_14410,N_9430,N_12407);
nor U14411 (N_14411,N_10410,N_9389);
and U14412 (N_14412,N_9898,N_11897);
nor U14413 (N_14413,N_9802,N_11856);
nor U14414 (N_14414,N_12009,N_10559);
or U14415 (N_14415,N_10164,N_11274);
nand U14416 (N_14416,N_10107,N_12254);
and U14417 (N_14417,N_11341,N_10891);
and U14418 (N_14418,N_12400,N_10523);
nand U14419 (N_14419,N_12348,N_9436);
and U14420 (N_14420,N_9539,N_9402);
or U14421 (N_14421,N_9415,N_10697);
nand U14422 (N_14422,N_11519,N_11366);
nand U14423 (N_14423,N_12136,N_10279);
nand U14424 (N_14424,N_11093,N_12283);
or U14425 (N_14425,N_11220,N_10240);
nand U14426 (N_14426,N_12291,N_10806);
nor U14427 (N_14427,N_10345,N_12098);
or U14428 (N_14428,N_11993,N_12232);
xnor U14429 (N_14429,N_12001,N_10412);
nor U14430 (N_14430,N_9627,N_10428);
or U14431 (N_14431,N_10866,N_11671);
or U14432 (N_14432,N_12484,N_11726);
or U14433 (N_14433,N_12272,N_10790);
xnor U14434 (N_14434,N_9793,N_10643);
nand U14435 (N_14435,N_10287,N_11781);
or U14436 (N_14436,N_10248,N_9699);
nor U14437 (N_14437,N_11381,N_10835);
nand U14438 (N_14438,N_9914,N_12489);
nand U14439 (N_14439,N_11365,N_11021);
or U14440 (N_14440,N_10498,N_11370);
nand U14441 (N_14441,N_12292,N_11126);
nand U14442 (N_14442,N_9868,N_10280);
nand U14443 (N_14443,N_11765,N_9800);
nor U14444 (N_14444,N_10588,N_10375);
nand U14445 (N_14445,N_12481,N_11350);
nor U14446 (N_14446,N_10470,N_11782);
and U14447 (N_14447,N_10544,N_12480);
nand U14448 (N_14448,N_10075,N_12032);
or U14449 (N_14449,N_12186,N_10620);
xor U14450 (N_14450,N_9511,N_11969);
nor U14451 (N_14451,N_11599,N_10161);
or U14452 (N_14452,N_9611,N_11167);
nand U14453 (N_14453,N_9426,N_11389);
or U14454 (N_14454,N_11794,N_10710);
nand U14455 (N_14455,N_11874,N_11538);
and U14456 (N_14456,N_10779,N_11573);
and U14457 (N_14457,N_9923,N_12173);
or U14458 (N_14458,N_10184,N_10771);
nor U14459 (N_14459,N_12083,N_10557);
nor U14460 (N_14460,N_9575,N_11960);
nand U14461 (N_14461,N_12149,N_11030);
nand U14462 (N_14462,N_10826,N_11794);
or U14463 (N_14463,N_11400,N_9463);
and U14464 (N_14464,N_12446,N_11479);
and U14465 (N_14465,N_11878,N_11800);
xnor U14466 (N_14466,N_9788,N_11369);
or U14467 (N_14467,N_11149,N_9864);
or U14468 (N_14468,N_11782,N_12140);
nand U14469 (N_14469,N_12398,N_9578);
xor U14470 (N_14470,N_9985,N_10045);
or U14471 (N_14471,N_10540,N_11227);
or U14472 (N_14472,N_12419,N_10367);
nor U14473 (N_14473,N_12089,N_10746);
nor U14474 (N_14474,N_10077,N_11143);
or U14475 (N_14475,N_10180,N_11736);
or U14476 (N_14476,N_10675,N_10221);
nor U14477 (N_14477,N_9415,N_9480);
and U14478 (N_14478,N_11066,N_10876);
nand U14479 (N_14479,N_11751,N_10067);
xor U14480 (N_14480,N_10924,N_10808);
nand U14481 (N_14481,N_10978,N_10651);
nand U14482 (N_14482,N_10385,N_12465);
nor U14483 (N_14483,N_11639,N_10760);
and U14484 (N_14484,N_10160,N_10730);
xor U14485 (N_14485,N_11764,N_10311);
and U14486 (N_14486,N_9378,N_9582);
and U14487 (N_14487,N_11856,N_10383);
nor U14488 (N_14488,N_9665,N_11319);
or U14489 (N_14489,N_9805,N_11776);
nor U14490 (N_14490,N_9989,N_11773);
and U14491 (N_14491,N_12408,N_10212);
or U14492 (N_14492,N_9474,N_11066);
nor U14493 (N_14493,N_9852,N_10903);
nand U14494 (N_14494,N_11438,N_10708);
and U14495 (N_14495,N_12066,N_12311);
or U14496 (N_14496,N_11637,N_11729);
nand U14497 (N_14497,N_11215,N_11282);
nand U14498 (N_14498,N_11211,N_11948);
or U14499 (N_14499,N_10113,N_9544);
or U14500 (N_14500,N_11659,N_10224);
and U14501 (N_14501,N_12378,N_10928);
and U14502 (N_14502,N_11765,N_9473);
and U14503 (N_14503,N_11911,N_11861);
xnor U14504 (N_14504,N_9385,N_12333);
and U14505 (N_14505,N_10500,N_11913);
nand U14506 (N_14506,N_10385,N_10368);
nor U14507 (N_14507,N_11948,N_12169);
nand U14508 (N_14508,N_9708,N_10194);
or U14509 (N_14509,N_10859,N_10992);
or U14510 (N_14510,N_11102,N_9740);
xnor U14511 (N_14511,N_9635,N_10463);
or U14512 (N_14512,N_10545,N_11004);
and U14513 (N_14513,N_9488,N_9727);
or U14514 (N_14514,N_10884,N_11316);
or U14515 (N_14515,N_11966,N_11272);
and U14516 (N_14516,N_10652,N_9885);
and U14517 (N_14517,N_12013,N_12169);
and U14518 (N_14518,N_10199,N_12400);
nor U14519 (N_14519,N_10826,N_11151);
nor U14520 (N_14520,N_11511,N_11249);
or U14521 (N_14521,N_11715,N_11639);
xnor U14522 (N_14522,N_10678,N_11643);
or U14523 (N_14523,N_12432,N_10058);
nor U14524 (N_14524,N_11295,N_11738);
or U14525 (N_14525,N_9708,N_9412);
or U14526 (N_14526,N_11773,N_12141);
nor U14527 (N_14527,N_12058,N_9981);
nand U14528 (N_14528,N_10944,N_11071);
nor U14529 (N_14529,N_10495,N_11302);
and U14530 (N_14530,N_9842,N_12142);
and U14531 (N_14531,N_12170,N_10387);
nand U14532 (N_14532,N_11906,N_9631);
or U14533 (N_14533,N_10892,N_10936);
xnor U14534 (N_14534,N_11258,N_11199);
nor U14535 (N_14535,N_11706,N_10285);
nor U14536 (N_14536,N_9841,N_10762);
nand U14537 (N_14537,N_10414,N_10043);
nand U14538 (N_14538,N_11017,N_10461);
xor U14539 (N_14539,N_10883,N_12337);
or U14540 (N_14540,N_10887,N_10649);
nand U14541 (N_14541,N_12362,N_10830);
and U14542 (N_14542,N_10827,N_11769);
nor U14543 (N_14543,N_11640,N_10906);
or U14544 (N_14544,N_12237,N_11648);
nand U14545 (N_14545,N_10837,N_12140);
nand U14546 (N_14546,N_10492,N_11644);
or U14547 (N_14547,N_9938,N_12249);
nor U14548 (N_14548,N_11208,N_10209);
nand U14549 (N_14549,N_10433,N_10007);
nand U14550 (N_14550,N_11242,N_12277);
or U14551 (N_14551,N_10637,N_11705);
nor U14552 (N_14552,N_10331,N_9428);
nand U14553 (N_14553,N_12048,N_9878);
or U14554 (N_14554,N_10808,N_10161);
nand U14555 (N_14555,N_12319,N_11745);
nand U14556 (N_14556,N_10632,N_10853);
nand U14557 (N_14557,N_10331,N_11728);
nor U14558 (N_14558,N_11909,N_10176);
nand U14559 (N_14559,N_11018,N_11509);
and U14560 (N_14560,N_12165,N_12088);
nor U14561 (N_14561,N_10478,N_11499);
xnor U14562 (N_14562,N_11155,N_12444);
xnor U14563 (N_14563,N_11775,N_12268);
nand U14564 (N_14564,N_10527,N_11815);
or U14565 (N_14565,N_10719,N_10962);
nand U14566 (N_14566,N_11457,N_9603);
nor U14567 (N_14567,N_9638,N_10096);
nor U14568 (N_14568,N_9522,N_10681);
nand U14569 (N_14569,N_11411,N_10672);
and U14570 (N_14570,N_12299,N_11207);
nand U14571 (N_14571,N_11394,N_11142);
or U14572 (N_14572,N_11580,N_12190);
or U14573 (N_14573,N_9730,N_10525);
and U14574 (N_14574,N_11843,N_10935);
nand U14575 (N_14575,N_10911,N_11019);
xor U14576 (N_14576,N_10068,N_10041);
nand U14577 (N_14577,N_9914,N_12099);
nand U14578 (N_14578,N_9760,N_10904);
or U14579 (N_14579,N_12406,N_11443);
and U14580 (N_14580,N_10007,N_11448);
or U14581 (N_14581,N_12345,N_10602);
nand U14582 (N_14582,N_10035,N_12080);
nor U14583 (N_14583,N_10500,N_12114);
nor U14584 (N_14584,N_10481,N_10730);
nand U14585 (N_14585,N_11108,N_10505);
nor U14586 (N_14586,N_9712,N_9602);
and U14587 (N_14587,N_9562,N_12119);
nor U14588 (N_14588,N_9416,N_9695);
or U14589 (N_14589,N_9980,N_12481);
nor U14590 (N_14590,N_10600,N_10095);
nand U14591 (N_14591,N_12382,N_10358);
or U14592 (N_14592,N_9873,N_11069);
nor U14593 (N_14593,N_10203,N_10844);
nand U14594 (N_14594,N_11376,N_11043);
nor U14595 (N_14595,N_11806,N_10258);
and U14596 (N_14596,N_9778,N_11830);
nand U14597 (N_14597,N_11745,N_11194);
nor U14598 (N_14598,N_9938,N_10896);
or U14599 (N_14599,N_10224,N_11082);
or U14600 (N_14600,N_11241,N_10718);
nor U14601 (N_14601,N_11994,N_11404);
or U14602 (N_14602,N_11434,N_11737);
or U14603 (N_14603,N_9945,N_9544);
or U14604 (N_14604,N_11003,N_12416);
nor U14605 (N_14605,N_9540,N_10689);
nor U14606 (N_14606,N_11185,N_10085);
nand U14607 (N_14607,N_9435,N_11999);
or U14608 (N_14608,N_12209,N_11677);
nand U14609 (N_14609,N_11627,N_11332);
nand U14610 (N_14610,N_9435,N_9721);
or U14611 (N_14611,N_10079,N_11829);
or U14612 (N_14612,N_11826,N_12489);
nor U14613 (N_14613,N_10158,N_10245);
and U14614 (N_14614,N_12057,N_9891);
and U14615 (N_14615,N_9728,N_9441);
nand U14616 (N_14616,N_10136,N_9501);
nand U14617 (N_14617,N_12221,N_9733);
xor U14618 (N_14618,N_12071,N_9637);
and U14619 (N_14619,N_10262,N_10037);
xnor U14620 (N_14620,N_10000,N_11276);
or U14621 (N_14621,N_11587,N_10564);
nor U14622 (N_14622,N_11411,N_12181);
nor U14623 (N_14623,N_10989,N_9711);
nor U14624 (N_14624,N_11911,N_11024);
or U14625 (N_14625,N_11509,N_12400);
or U14626 (N_14626,N_11938,N_11277);
and U14627 (N_14627,N_10746,N_11574);
and U14628 (N_14628,N_9446,N_12404);
or U14629 (N_14629,N_9970,N_11016);
and U14630 (N_14630,N_11960,N_10683);
and U14631 (N_14631,N_9975,N_10179);
xnor U14632 (N_14632,N_9942,N_12201);
and U14633 (N_14633,N_11607,N_11110);
nor U14634 (N_14634,N_11234,N_11439);
and U14635 (N_14635,N_12316,N_12419);
nand U14636 (N_14636,N_11147,N_11467);
or U14637 (N_14637,N_11533,N_11190);
and U14638 (N_14638,N_9475,N_10580);
nand U14639 (N_14639,N_10523,N_10110);
nor U14640 (N_14640,N_12408,N_12063);
nor U14641 (N_14641,N_11257,N_11941);
nor U14642 (N_14642,N_11460,N_10080);
nand U14643 (N_14643,N_9424,N_11813);
nand U14644 (N_14644,N_12366,N_12210);
xor U14645 (N_14645,N_12177,N_10236);
nor U14646 (N_14646,N_11216,N_12271);
xor U14647 (N_14647,N_10915,N_10639);
nor U14648 (N_14648,N_10598,N_12227);
nor U14649 (N_14649,N_11480,N_9478);
or U14650 (N_14650,N_11515,N_12376);
nand U14651 (N_14651,N_10344,N_11254);
nand U14652 (N_14652,N_11356,N_9736);
nor U14653 (N_14653,N_9623,N_10307);
nor U14654 (N_14654,N_10229,N_10503);
nor U14655 (N_14655,N_11213,N_12271);
nor U14656 (N_14656,N_12363,N_12420);
nand U14657 (N_14657,N_11566,N_12098);
or U14658 (N_14658,N_11919,N_11993);
and U14659 (N_14659,N_11698,N_9599);
xor U14660 (N_14660,N_12412,N_12349);
or U14661 (N_14661,N_10963,N_10318);
nor U14662 (N_14662,N_12447,N_10527);
nor U14663 (N_14663,N_10351,N_11440);
and U14664 (N_14664,N_12031,N_9534);
nor U14665 (N_14665,N_11205,N_9561);
xor U14666 (N_14666,N_10340,N_9812);
and U14667 (N_14667,N_11433,N_11742);
nand U14668 (N_14668,N_10439,N_10774);
or U14669 (N_14669,N_12164,N_9530);
and U14670 (N_14670,N_10821,N_11940);
xor U14671 (N_14671,N_9381,N_9602);
or U14672 (N_14672,N_11377,N_12120);
nor U14673 (N_14673,N_10509,N_10556);
nand U14674 (N_14674,N_10274,N_10036);
nand U14675 (N_14675,N_9955,N_9403);
and U14676 (N_14676,N_11043,N_10625);
nand U14677 (N_14677,N_11577,N_10703);
and U14678 (N_14678,N_10080,N_11507);
or U14679 (N_14679,N_10648,N_9411);
nor U14680 (N_14680,N_11171,N_11860);
xnor U14681 (N_14681,N_11354,N_12051);
nor U14682 (N_14682,N_10163,N_9663);
nand U14683 (N_14683,N_9420,N_9586);
nor U14684 (N_14684,N_10030,N_12407);
and U14685 (N_14685,N_11510,N_12253);
xnor U14686 (N_14686,N_9488,N_12289);
nor U14687 (N_14687,N_11834,N_12425);
and U14688 (N_14688,N_12262,N_9916);
and U14689 (N_14689,N_11839,N_11043);
nand U14690 (N_14690,N_11774,N_9449);
xnor U14691 (N_14691,N_10171,N_11174);
and U14692 (N_14692,N_11622,N_12432);
and U14693 (N_14693,N_10716,N_9810);
and U14694 (N_14694,N_11069,N_10554);
and U14695 (N_14695,N_11384,N_9451);
and U14696 (N_14696,N_9751,N_9568);
or U14697 (N_14697,N_10993,N_11209);
or U14698 (N_14698,N_10590,N_12290);
and U14699 (N_14699,N_10973,N_12095);
nor U14700 (N_14700,N_11562,N_11249);
nand U14701 (N_14701,N_10010,N_10407);
xor U14702 (N_14702,N_11476,N_11330);
and U14703 (N_14703,N_10400,N_9690);
nor U14704 (N_14704,N_10958,N_9462);
or U14705 (N_14705,N_12253,N_12115);
nor U14706 (N_14706,N_9854,N_11770);
and U14707 (N_14707,N_12119,N_10801);
nor U14708 (N_14708,N_9569,N_10010);
and U14709 (N_14709,N_10251,N_9751);
xor U14710 (N_14710,N_10778,N_11171);
nand U14711 (N_14711,N_12351,N_11061);
xnor U14712 (N_14712,N_10027,N_11255);
xor U14713 (N_14713,N_11405,N_10154);
and U14714 (N_14714,N_10649,N_9844);
nand U14715 (N_14715,N_9732,N_10208);
or U14716 (N_14716,N_10954,N_11518);
and U14717 (N_14717,N_9847,N_11939);
nand U14718 (N_14718,N_11156,N_12358);
nand U14719 (N_14719,N_12194,N_12407);
or U14720 (N_14720,N_9788,N_10818);
or U14721 (N_14721,N_9644,N_11897);
nor U14722 (N_14722,N_9843,N_9515);
and U14723 (N_14723,N_11773,N_12386);
nand U14724 (N_14724,N_11243,N_9417);
nor U14725 (N_14725,N_12034,N_11583);
and U14726 (N_14726,N_10908,N_11371);
or U14727 (N_14727,N_9908,N_11577);
and U14728 (N_14728,N_9658,N_10131);
nand U14729 (N_14729,N_9651,N_10069);
and U14730 (N_14730,N_10751,N_10126);
xor U14731 (N_14731,N_12211,N_10996);
nor U14732 (N_14732,N_9877,N_11249);
xnor U14733 (N_14733,N_12451,N_11510);
and U14734 (N_14734,N_12498,N_10229);
and U14735 (N_14735,N_9975,N_10553);
and U14736 (N_14736,N_9401,N_10134);
and U14737 (N_14737,N_10474,N_11474);
or U14738 (N_14738,N_12355,N_10938);
nor U14739 (N_14739,N_11857,N_10488);
nor U14740 (N_14740,N_11797,N_11716);
or U14741 (N_14741,N_9447,N_12238);
nor U14742 (N_14742,N_11271,N_10263);
and U14743 (N_14743,N_10504,N_9484);
and U14744 (N_14744,N_11122,N_11494);
or U14745 (N_14745,N_10654,N_11596);
or U14746 (N_14746,N_11456,N_11437);
and U14747 (N_14747,N_9434,N_9973);
nor U14748 (N_14748,N_12207,N_10368);
nand U14749 (N_14749,N_12317,N_9626);
xor U14750 (N_14750,N_10844,N_9975);
or U14751 (N_14751,N_10289,N_11602);
or U14752 (N_14752,N_10680,N_12376);
nand U14753 (N_14753,N_12036,N_11637);
and U14754 (N_14754,N_11156,N_10026);
or U14755 (N_14755,N_11198,N_11976);
nand U14756 (N_14756,N_9948,N_10062);
xor U14757 (N_14757,N_11575,N_11813);
nand U14758 (N_14758,N_9505,N_11944);
nand U14759 (N_14759,N_11961,N_9416);
nor U14760 (N_14760,N_10301,N_11620);
nor U14761 (N_14761,N_11582,N_10539);
nor U14762 (N_14762,N_10672,N_9534);
nand U14763 (N_14763,N_9865,N_9420);
or U14764 (N_14764,N_9508,N_9593);
or U14765 (N_14765,N_10427,N_10512);
and U14766 (N_14766,N_10264,N_11790);
nor U14767 (N_14767,N_11384,N_9654);
nor U14768 (N_14768,N_9542,N_12188);
xor U14769 (N_14769,N_12486,N_11346);
or U14770 (N_14770,N_11587,N_9432);
or U14771 (N_14771,N_12480,N_10108);
and U14772 (N_14772,N_9590,N_11818);
nand U14773 (N_14773,N_10613,N_10780);
and U14774 (N_14774,N_10110,N_12338);
nand U14775 (N_14775,N_10342,N_11943);
or U14776 (N_14776,N_11892,N_9637);
or U14777 (N_14777,N_10143,N_11976);
or U14778 (N_14778,N_12324,N_9665);
and U14779 (N_14779,N_11513,N_11065);
xor U14780 (N_14780,N_9662,N_12165);
nor U14781 (N_14781,N_10830,N_12102);
nor U14782 (N_14782,N_12397,N_10406);
and U14783 (N_14783,N_12303,N_9996);
nor U14784 (N_14784,N_10168,N_10937);
nor U14785 (N_14785,N_11253,N_11502);
and U14786 (N_14786,N_12395,N_9951);
nand U14787 (N_14787,N_10387,N_9517);
nand U14788 (N_14788,N_10496,N_10867);
nand U14789 (N_14789,N_11683,N_12395);
nor U14790 (N_14790,N_12402,N_11888);
or U14791 (N_14791,N_9537,N_12458);
nor U14792 (N_14792,N_12113,N_11160);
xor U14793 (N_14793,N_9800,N_10366);
nand U14794 (N_14794,N_11931,N_11797);
nand U14795 (N_14795,N_11737,N_9461);
xnor U14796 (N_14796,N_10759,N_10260);
or U14797 (N_14797,N_11551,N_9785);
xnor U14798 (N_14798,N_11918,N_11366);
xor U14799 (N_14799,N_11444,N_11307);
or U14800 (N_14800,N_9828,N_12009);
and U14801 (N_14801,N_10797,N_9843);
nor U14802 (N_14802,N_11199,N_12247);
xnor U14803 (N_14803,N_10533,N_11502);
xnor U14804 (N_14804,N_11870,N_9999);
or U14805 (N_14805,N_11584,N_10581);
nor U14806 (N_14806,N_12303,N_11263);
nand U14807 (N_14807,N_9437,N_10223);
or U14808 (N_14808,N_12041,N_11195);
nand U14809 (N_14809,N_9854,N_9954);
xnor U14810 (N_14810,N_10008,N_10210);
or U14811 (N_14811,N_10972,N_12092);
or U14812 (N_14812,N_9804,N_10095);
and U14813 (N_14813,N_9710,N_11842);
or U14814 (N_14814,N_11010,N_9569);
nor U14815 (N_14815,N_10434,N_10302);
and U14816 (N_14816,N_11016,N_11869);
and U14817 (N_14817,N_10553,N_10762);
and U14818 (N_14818,N_11126,N_10070);
nor U14819 (N_14819,N_12453,N_11661);
or U14820 (N_14820,N_9627,N_9737);
and U14821 (N_14821,N_10439,N_10381);
nor U14822 (N_14822,N_12282,N_10307);
and U14823 (N_14823,N_11612,N_12321);
nor U14824 (N_14824,N_11109,N_10899);
nand U14825 (N_14825,N_10544,N_9887);
nor U14826 (N_14826,N_10189,N_10481);
or U14827 (N_14827,N_11288,N_10450);
and U14828 (N_14828,N_11468,N_11395);
or U14829 (N_14829,N_11984,N_11972);
and U14830 (N_14830,N_12068,N_10570);
nand U14831 (N_14831,N_10726,N_9450);
and U14832 (N_14832,N_10415,N_9885);
or U14833 (N_14833,N_10293,N_9918);
and U14834 (N_14834,N_10925,N_11939);
nor U14835 (N_14835,N_9900,N_10403);
nand U14836 (N_14836,N_12286,N_10033);
nand U14837 (N_14837,N_9917,N_10955);
and U14838 (N_14838,N_10774,N_12181);
nor U14839 (N_14839,N_11618,N_9423);
and U14840 (N_14840,N_11562,N_11507);
nor U14841 (N_14841,N_9906,N_10917);
nor U14842 (N_14842,N_11441,N_10369);
nand U14843 (N_14843,N_10061,N_9602);
and U14844 (N_14844,N_12308,N_10748);
nand U14845 (N_14845,N_10207,N_12467);
nor U14846 (N_14846,N_11720,N_12007);
or U14847 (N_14847,N_10824,N_9438);
nor U14848 (N_14848,N_10789,N_11962);
or U14849 (N_14849,N_11140,N_9569);
or U14850 (N_14850,N_11694,N_12081);
and U14851 (N_14851,N_10046,N_11840);
and U14852 (N_14852,N_11152,N_11044);
nor U14853 (N_14853,N_11782,N_9505);
or U14854 (N_14854,N_10304,N_12206);
nand U14855 (N_14855,N_10104,N_10101);
nor U14856 (N_14856,N_10472,N_11580);
nand U14857 (N_14857,N_11321,N_10087);
and U14858 (N_14858,N_12134,N_9578);
xor U14859 (N_14859,N_11292,N_9708);
nand U14860 (N_14860,N_11225,N_10465);
nor U14861 (N_14861,N_11756,N_10867);
nor U14862 (N_14862,N_10923,N_9823);
and U14863 (N_14863,N_9702,N_9846);
and U14864 (N_14864,N_11239,N_9946);
and U14865 (N_14865,N_11984,N_9886);
xnor U14866 (N_14866,N_10076,N_10754);
and U14867 (N_14867,N_12166,N_11592);
nand U14868 (N_14868,N_11076,N_10043);
or U14869 (N_14869,N_11592,N_9565);
or U14870 (N_14870,N_11778,N_12264);
or U14871 (N_14871,N_9559,N_9390);
or U14872 (N_14872,N_9787,N_10506);
and U14873 (N_14873,N_10641,N_10624);
nand U14874 (N_14874,N_11200,N_9969);
and U14875 (N_14875,N_11016,N_10723);
nor U14876 (N_14876,N_10453,N_10654);
and U14877 (N_14877,N_10089,N_10512);
or U14878 (N_14878,N_12124,N_10907);
nor U14879 (N_14879,N_10963,N_10983);
nand U14880 (N_14880,N_11101,N_10607);
nand U14881 (N_14881,N_10544,N_10798);
or U14882 (N_14882,N_11276,N_10379);
or U14883 (N_14883,N_10190,N_10702);
and U14884 (N_14884,N_10636,N_12360);
or U14885 (N_14885,N_10433,N_11290);
or U14886 (N_14886,N_11174,N_11322);
or U14887 (N_14887,N_12404,N_12409);
and U14888 (N_14888,N_11575,N_12271);
nor U14889 (N_14889,N_9512,N_12255);
or U14890 (N_14890,N_9703,N_9462);
or U14891 (N_14891,N_11331,N_12358);
nand U14892 (N_14892,N_10524,N_10301);
nand U14893 (N_14893,N_9395,N_9969);
nor U14894 (N_14894,N_11722,N_11684);
or U14895 (N_14895,N_12088,N_12278);
and U14896 (N_14896,N_11940,N_12222);
nor U14897 (N_14897,N_10821,N_11688);
or U14898 (N_14898,N_11788,N_10943);
xor U14899 (N_14899,N_10860,N_11978);
and U14900 (N_14900,N_11888,N_10496);
or U14901 (N_14901,N_11118,N_11540);
and U14902 (N_14902,N_12448,N_11155);
nor U14903 (N_14903,N_10732,N_9803);
nor U14904 (N_14904,N_9870,N_10983);
or U14905 (N_14905,N_12095,N_11406);
or U14906 (N_14906,N_10285,N_12053);
nor U14907 (N_14907,N_11286,N_9478);
or U14908 (N_14908,N_12048,N_12221);
and U14909 (N_14909,N_10778,N_12266);
nand U14910 (N_14910,N_9461,N_11922);
or U14911 (N_14911,N_11824,N_11844);
nor U14912 (N_14912,N_12038,N_11003);
nor U14913 (N_14913,N_12298,N_11211);
nor U14914 (N_14914,N_10052,N_12252);
nand U14915 (N_14915,N_10083,N_10927);
and U14916 (N_14916,N_11983,N_9813);
and U14917 (N_14917,N_10319,N_12024);
and U14918 (N_14918,N_10874,N_9478);
or U14919 (N_14919,N_9446,N_11545);
and U14920 (N_14920,N_10881,N_11698);
nor U14921 (N_14921,N_10275,N_12041);
xor U14922 (N_14922,N_11231,N_9603);
and U14923 (N_14923,N_10715,N_10785);
nor U14924 (N_14924,N_11738,N_11814);
nor U14925 (N_14925,N_10235,N_11607);
or U14926 (N_14926,N_12270,N_12436);
or U14927 (N_14927,N_11503,N_11378);
and U14928 (N_14928,N_11222,N_10682);
or U14929 (N_14929,N_11202,N_11248);
xnor U14930 (N_14930,N_10856,N_9956);
and U14931 (N_14931,N_11928,N_9596);
or U14932 (N_14932,N_11562,N_12344);
or U14933 (N_14933,N_9861,N_10267);
nand U14934 (N_14934,N_11261,N_11819);
nand U14935 (N_14935,N_11947,N_12251);
nand U14936 (N_14936,N_10053,N_12021);
and U14937 (N_14937,N_12460,N_9546);
or U14938 (N_14938,N_11339,N_10798);
nand U14939 (N_14939,N_12320,N_9509);
xor U14940 (N_14940,N_9381,N_9716);
xnor U14941 (N_14941,N_10562,N_10499);
or U14942 (N_14942,N_11777,N_10806);
or U14943 (N_14943,N_10720,N_12334);
nand U14944 (N_14944,N_9518,N_11735);
nand U14945 (N_14945,N_9830,N_11171);
or U14946 (N_14946,N_11966,N_9954);
nand U14947 (N_14947,N_10759,N_11474);
or U14948 (N_14948,N_11887,N_9653);
nand U14949 (N_14949,N_10530,N_10799);
or U14950 (N_14950,N_9475,N_11533);
and U14951 (N_14951,N_12318,N_9883);
xnor U14952 (N_14952,N_9938,N_10928);
xnor U14953 (N_14953,N_10155,N_12393);
or U14954 (N_14954,N_9617,N_9625);
or U14955 (N_14955,N_10223,N_9833);
nand U14956 (N_14956,N_10858,N_10875);
xnor U14957 (N_14957,N_10779,N_11067);
and U14958 (N_14958,N_12158,N_9528);
and U14959 (N_14959,N_10207,N_9680);
nor U14960 (N_14960,N_10584,N_9419);
or U14961 (N_14961,N_11885,N_10160);
and U14962 (N_14962,N_11739,N_10575);
nor U14963 (N_14963,N_12243,N_10000);
or U14964 (N_14964,N_12255,N_11622);
nand U14965 (N_14965,N_12361,N_10597);
nor U14966 (N_14966,N_11539,N_10252);
or U14967 (N_14967,N_12220,N_10413);
nor U14968 (N_14968,N_12077,N_12472);
nand U14969 (N_14969,N_11035,N_10851);
or U14970 (N_14970,N_11489,N_11641);
nand U14971 (N_14971,N_11999,N_10146);
nand U14972 (N_14972,N_11911,N_10472);
or U14973 (N_14973,N_9418,N_10135);
xor U14974 (N_14974,N_12285,N_10412);
nand U14975 (N_14975,N_11519,N_11040);
nand U14976 (N_14976,N_11564,N_10697);
or U14977 (N_14977,N_12282,N_11653);
xnor U14978 (N_14978,N_9968,N_10024);
nor U14979 (N_14979,N_12243,N_10796);
nand U14980 (N_14980,N_10717,N_10157);
and U14981 (N_14981,N_9409,N_12271);
nand U14982 (N_14982,N_11490,N_11201);
nor U14983 (N_14983,N_10735,N_11220);
or U14984 (N_14984,N_9620,N_10213);
and U14985 (N_14985,N_10071,N_11219);
and U14986 (N_14986,N_11424,N_10861);
xnor U14987 (N_14987,N_10314,N_9630);
or U14988 (N_14988,N_11625,N_11775);
xnor U14989 (N_14989,N_12114,N_10074);
or U14990 (N_14990,N_11840,N_10435);
or U14991 (N_14991,N_9723,N_11997);
xor U14992 (N_14992,N_11876,N_10728);
xor U14993 (N_14993,N_9851,N_11333);
nor U14994 (N_14994,N_9990,N_10434);
nand U14995 (N_14995,N_11323,N_9654);
or U14996 (N_14996,N_11522,N_10661);
nor U14997 (N_14997,N_9502,N_10357);
nand U14998 (N_14998,N_10297,N_11306);
nand U14999 (N_14999,N_12220,N_10058);
or U15000 (N_15000,N_10098,N_11056);
nand U15001 (N_15001,N_9610,N_9999);
or U15002 (N_15002,N_10628,N_10503);
or U15003 (N_15003,N_10761,N_10817);
or U15004 (N_15004,N_11464,N_9501);
or U15005 (N_15005,N_9417,N_11315);
xor U15006 (N_15006,N_11290,N_10696);
and U15007 (N_15007,N_12162,N_10828);
xor U15008 (N_15008,N_9396,N_9390);
and U15009 (N_15009,N_12336,N_10474);
nand U15010 (N_15010,N_12117,N_11187);
or U15011 (N_15011,N_11656,N_9475);
nor U15012 (N_15012,N_12119,N_10366);
or U15013 (N_15013,N_11813,N_11007);
nand U15014 (N_15014,N_10366,N_9492);
or U15015 (N_15015,N_11634,N_10929);
nand U15016 (N_15016,N_10341,N_9667);
nand U15017 (N_15017,N_12288,N_9617);
nor U15018 (N_15018,N_10235,N_9592);
nor U15019 (N_15019,N_12095,N_12366);
or U15020 (N_15020,N_12101,N_10409);
and U15021 (N_15021,N_12235,N_10768);
nor U15022 (N_15022,N_12122,N_11055);
nor U15023 (N_15023,N_9963,N_9868);
nor U15024 (N_15024,N_11033,N_10703);
and U15025 (N_15025,N_11291,N_10850);
xnor U15026 (N_15026,N_11232,N_11802);
nand U15027 (N_15027,N_10002,N_12148);
and U15028 (N_15028,N_11036,N_11717);
nor U15029 (N_15029,N_11451,N_9917);
nand U15030 (N_15030,N_10623,N_12490);
nand U15031 (N_15031,N_11368,N_10342);
nand U15032 (N_15032,N_12037,N_10163);
xor U15033 (N_15033,N_10774,N_10643);
or U15034 (N_15034,N_10656,N_11110);
and U15035 (N_15035,N_9386,N_11580);
or U15036 (N_15036,N_9608,N_12187);
and U15037 (N_15037,N_12315,N_11445);
nor U15038 (N_15038,N_9897,N_9736);
nor U15039 (N_15039,N_9774,N_12116);
and U15040 (N_15040,N_9457,N_10466);
nand U15041 (N_15041,N_10074,N_11835);
and U15042 (N_15042,N_11307,N_11818);
and U15043 (N_15043,N_10694,N_10997);
and U15044 (N_15044,N_11455,N_10659);
nand U15045 (N_15045,N_12062,N_9562);
and U15046 (N_15046,N_10766,N_10573);
nand U15047 (N_15047,N_9983,N_10297);
nand U15048 (N_15048,N_10006,N_10442);
and U15049 (N_15049,N_12225,N_10894);
and U15050 (N_15050,N_9565,N_11890);
nor U15051 (N_15051,N_11628,N_11352);
nor U15052 (N_15052,N_9913,N_10429);
nor U15053 (N_15053,N_12070,N_10934);
or U15054 (N_15054,N_10379,N_10732);
nand U15055 (N_15055,N_10577,N_9899);
xnor U15056 (N_15056,N_9651,N_11904);
nor U15057 (N_15057,N_10032,N_10848);
nor U15058 (N_15058,N_11598,N_9512);
nor U15059 (N_15059,N_10305,N_11267);
nand U15060 (N_15060,N_12116,N_12396);
or U15061 (N_15061,N_10363,N_10826);
and U15062 (N_15062,N_11172,N_9508);
and U15063 (N_15063,N_12083,N_10406);
or U15064 (N_15064,N_10513,N_11335);
xor U15065 (N_15065,N_10365,N_11535);
or U15066 (N_15066,N_12175,N_10060);
or U15067 (N_15067,N_10341,N_11379);
and U15068 (N_15068,N_11992,N_11372);
xor U15069 (N_15069,N_10858,N_11785);
xor U15070 (N_15070,N_12002,N_9593);
nor U15071 (N_15071,N_12359,N_9895);
nor U15072 (N_15072,N_11515,N_10956);
nor U15073 (N_15073,N_12423,N_11578);
and U15074 (N_15074,N_11917,N_12395);
and U15075 (N_15075,N_11692,N_9628);
and U15076 (N_15076,N_11676,N_10315);
nand U15077 (N_15077,N_12359,N_9976);
nor U15078 (N_15078,N_10687,N_9523);
nand U15079 (N_15079,N_9731,N_10275);
nand U15080 (N_15080,N_9786,N_9433);
or U15081 (N_15081,N_11704,N_10813);
nor U15082 (N_15082,N_11512,N_10900);
xor U15083 (N_15083,N_12327,N_10698);
xor U15084 (N_15084,N_9634,N_11128);
or U15085 (N_15085,N_10004,N_10081);
xnor U15086 (N_15086,N_10465,N_10911);
xnor U15087 (N_15087,N_11058,N_12495);
or U15088 (N_15088,N_11536,N_10859);
nor U15089 (N_15089,N_12384,N_10270);
xor U15090 (N_15090,N_11573,N_10718);
nor U15091 (N_15091,N_10790,N_11559);
and U15092 (N_15092,N_11209,N_10871);
xor U15093 (N_15093,N_12409,N_9538);
xnor U15094 (N_15094,N_11502,N_10687);
nor U15095 (N_15095,N_11227,N_9974);
nor U15096 (N_15096,N_10759,N_12497);
nand U15097 (N_15097,N_11410,N_10394);
nor U15098 (N_15098,N_10554,N_11481);
and U15099 (N_15099,N_10906,N_9651);
nor U15100 (N_15100,N_12367,N_11561);
or U15101 (N_15101,N_9732,N_9797);
and U15102 (N_15102,N_10894,N_9571);
nand U15103 (N_15103,N_9551,N_11461);
nand U15104 (N_15104,N_10221,N_10579);
and U15105 (N_15105,N_10007,N_11800);
nand U15106 (N_15106,N_9513,N_10204);
or U15107 (N_15107,N_11015,N_10365);
nor U15108 (N_15108,N_11631,N_11120);
xor U15109 (N_15109,N_11524,N_11635);
nand U15110 (N_15110,N_11049,N_10455);
xor U15111 (N_15111,N_11264,N_12341);
and U15112 (N_15112,N_11182,N_11293);
nor U15113 (N_15113,N_11735,N_12234);
or U15114 (N_15114,N_12215,N_10492);
and U15115 (N_15115,N_9491,N_12081);
nand U15116 (N_15116,N_12143,N_11677);
and U15117 (N_15117,N_9389,N_9568);
or U15118 (N_15118,N_9753,N_11420);
nor U15119 (N_15119,N_11366,N_11883);
nor U15120 (N_15120,N_11699,N_10425);
xor U15121 (N_15121,N_9484,N_9581);
or U15122 (N_15122,N_9819,N_11149);
or U15123 (N_15123,N_12441,N_9849);
nand U15124 (N_15124,N_10430,N_9824);
nand U15125 (N_15125,N_10935,N_10033);
nand U15126 (N_15126,N_10087,N_10366);
and U15127 (N_15127,N_11961,N_9515);
or U15128 (N_15128,N_10703,N_10090);
xor U15129 (N_15129,N_10261,N_11583);
nand U15130 (N_15130,N_10479,N_9989);
and U15131 (N_15131,N_12320,N_11569);
nor U15132 (N_15132,N_12422,N_10412);
and U15133 (N_15133,N_11871,N_10379);
nand U15134 (N_15134,N_10470,N_9406);
nand U15135 (N_15135,N_9822,N_12035);
nor U15136 (N_15136,N_11856,N_9686);
or U15137 (N_15137,N_9437,N_10384);
nand U15138 (N_15138,N_9551,N_11771);
or U15139 (N_15139,N_10574,N_9424);
xor U15140 (N_15140,N_10268,N_12046);
xnor U15141 (N_15141,N_9707,N_9968);
nand U15142 (N_15142,N_11442,N_10485);
or U15143 (N_15143,N_10613,N_11378);
or U15144 (N_15144,N_10069,N_9785);
xor U15145 (N_15145,N_9980,N_10821);
nor U15146 (N_15146,N_9797,N_9542);
and U15147 (N_15147,N_10654,N_11697);
nor U15148 (N_15148,N_11104,N_9576);
nor U15149 (N_15149,N_11271,N_12375);
or U15150 (N_15150,N_11407,N_10480);
nor U15151 (N_15151,N_12433,N_9872);
or U15152 (N_15152,N_11914,N_12491);
and U15153 (N_15153,N_10555,N_11881);
and U15154 (N_15154,N_10505,N_10001);
or U15155 (N_15155,N_10724,N_10315);
nor U15156 (N_15156,N_11055,N_11162);
xnor U15157 (N_15157,N_9843,N_10533);
or U15158 (N_15158,N_10182,N_10639);
nand U15159 (N_15159,N_11515,N_9392);
nor U15160 (N_15160,N_9878,N_12166);
nor U15161 (N_15161,N_10762,N_9860);
nand U15162 (N_15162,N_12142,N_11957);
nor U15163 (N_15163,N_9830,N_11631);
nor U15164 (N_15164,N_9399,N_11677);
xor U15165 (N_15165,N_11895,N_9576);
or U15166 (N_15166,N_9603,N_10507);
nand U15167 (N_15167,N_11137,N_10643);
and U15168 (N_15168,N_11601,N_12003);
or U15169 (N_15169,N_9392,N_11285);
and U15170 (N_15170,N_9737,N_10694);
nand U15171 (N_15171,N_11246,N_11957);
nor U15172 (N_15172,N_9502,N_12386);
and U15173 (N_15173,N_10642,N_12170);
and U15174 (N_15174,N_11041,N_9910);
or U15175 (N_15175,N_12082,N_12180);
nor U15176 (N_15176,N_9613,N_9514);
nand U15177 (N_15177,N_10488,N_11442);
nor U15178 (N_15178,N_12255,N_9416);
or U15179 (N_15179,N_11432,N_10582);
and U15180 (N_15180,N_11839,N_10310);
nand U15181 (N_15181,N_9762,N_10494);
nor U15182 (N_15182,N_10320,N_9923);
nor U15183 (N_15183,N_9420,N_9887);
nand U15184 (N_15184,N_10527,N_10903);
nor U15185 (N_15185,N_9632,N_10821);
or U15186 (N_15186,N_9646,N_10172);
and U15187 (N_15187,N_10150,N_11983);
nor U15188 (N_15188,N_10621,N_11850);
and U15189 (N_15189,N_12129,N_12324);
nand U15190 (N_15190,N_9751,N_9837);
and U15191 (N_15191,N_10704,N_10397);
or U15192 (N_15192,N_12203,N_12441);
nor U15193 (N_15193,N_11111,N_11127);
nor U15194 (N_15194,N_12136,N_12105);
nand U15195 (N_15195,N_11855,N_9473);
nor U15196 (N_15196,N_11927,N_10203);
or U15197 (N_15197,N_10600,N_10050);
and U15198 (N_15198,N_11387,N_12243);
and U15199 (N_15199,N_11615,N_11887);
xor U15200 (N_15200,N_9853,N_10946);
xor U15201 (N_15201,N_10562,N_10089);
nand U15202 (N_15202,N_11081,N_9932);
nand U15203 (N_15203,N_11060,N_12452);
and U15204 (N_15204,N_9689,N_10198);
nor U15205 (N_15205,N_10576,N_11213);
xor U15206 (N_15206,N_10640,N_11537);
or U15207 (N_15207,N_11133,N_9747);
nand U15208 (N_15208,N_10326,N_9530);
nor U15209 (N_15209,N_10460,N_10100);
and U15210 (N_15210,N_11462,N_11725);
and U15211 (N_15211,N_10514,N_10799);
or U15212 (N_15212,N_11614,N_12388);
and U15213 (N_15213,N_10091,N_10852);
and U15214 (N_15214,N_11817,N_9911);
nand U15215 (N_15215,N_10921,N_11896);
xor U15216 (N_15216,N_11406,N_10034);
nor U15217 (N_15217,N_10784,N_11112);
nand U15218 (N_15218,N_10949,N_11474);
nor U15219 (N_15219,N_12249,N_12399);
and U15220 (N_15220,N_11397,N_11807);
nand U15221 (N_15221,N_12217,N_9840);
or U15222 (N_15222,N_9764,N_11254);
and U15223 (N_15223,N_11830,N_10301);
nor U15224 (N_15224,N_11339,N_11582);
and U15225 (N_15225,N_10770,N_12161);
nand U15226 (N_15226,N_9483,N_9946);
nor U15227 (N_15227,N_11618,N_9605);
nor U15228 (N_15228,N_10893,N_9586);
nor U15229 (N_15229,N_12043,N_10636);
nor U15230 (N_15230,N_11379,N_9850);
nor U15231 (N_15231,N_9407,N_10393);
nor U15232 (N_15232,N_12469,N_11413);
nor U15233 (N_15233,N_12210,N_11006);
nor U15234 (N_15234,N_11636,N_9960);
and U15235 (N_15235,N_12119,N_10388);
xnor U15236 (N_15236,N_11616,N_12074);
and U15237 (N_15237,N_11754,N_10609);
nor U15238 (N_15238,N_11524,N_10725);
nor U15239 (N_15239,N_11989,N_11107);
nand U15240 (N_15240,N_11975,N_10891);
or U15241 (N_15241,N_9728,N_9619);
xnor U15242 (N_15242,N_9526,N_10973);
nor U15243 (N_15243,N_12402,N_11319);
nor U15244 (N_15244,N_10525,N_9824);
nor U15245 (N_15245,N_10032,N_10785);
and U15246 (N_15246,N_11886,N_12338);
nor U15247 (N_15247,N_9680,N_11255);
or U15248 (N_15248,N_11521,N_9411);
nor U15249 (N_15249,N_11594,N_9800);
nor U15250 (N_15250,N_9781,N_9960);
xnor U15251 (N_15251,N_9966,N_12087);
nor U15252 (N_15252,N_10213,N_9564);
nor U15253 (N_15253,N_9659,N_11727);
or U15254 (N_15254,N_11645,N_12462);
and U15255 (N_15255,N_10857,N_9572);
or U15256 (N_15256,N_10807,N_10823);
nor U15257 (N_15257,N_9490,N_12392);
or U15258 (N_15258,N_12183,N_9671);
nand U15259 (N_15259,N_11657,N_11630);
or U15260 (N_15260,N_12397,N_9655);
or U15261 (N_15261,N_10610,N_9917);
nor U15262 (N_15262,N_9555,N_10448);
and U15263 (N_15263,N_12286,N_10064);
nor U15264 (N_15264,N_10893,N_9645);
and U15265 (N_15265,N_10753,N_11448);
nand U15266 (N_15266,N_10895,N_11344);
and U15267 (N_15267,N_10619,N_10913);
nand U15268 (N_15268,N_12018,N_10777);
or U15269 (N_15269,N_9924,N_11314);
or U15270 (N_15270,N_12146,N_10854);
or U15271 (N_15271,N_10465,N_9546);
or U15272 (N_15272,N_11014,N_12004);
and U15273 (N_15273,N_12483,N_10487);
nor U15274 (N_15274,N_9847,N_10433);
xnor U15275 (N_15275,N_11538,N_9578);
and U15276 (N_15276,N_10480,N_9640);
nand U15277 (N_15277,N_11817,N_12005);
nand U15278 (N_15278,N_10109,N_9467);
and U15279 (N_15279,N_10411,N_10261);
nand U15280 (N_15280,N_11878,N_9645);
and U15281 (N_15281,N_11254,N_10048);
nand U15282 (N_15282,N_10329,N_10070);
nand U15283 (N_15283,N_10546,N_12269);
or U15284 (N_15284,N_9891,N_10622);
nor U15285 (N_15285,N_10958,N_9541);
and U15286 (N_15286,N_9378,N_12237);
and U15287 (N_15287,N_10265,N_11224);
and U15288 (N_15288,N_11790,N_11814);
nor U15289 (N_15289,N_10090,N_10429);
xor U15290 (N_15290,N_9654,N_12110);
nor U15291 (N_15291,N_12229,N_12200);
and U15292 (N_15292,N_11789,N_10065);
nor U15293 (N_15293,N_11426,N_12154);
or U15294 (N_15294,N_12143,N_9527);
nor U15295 (N_15295,N_11901,N_11052);
or U15296 (N_15296,N_11675,N_11476);
nor U15297 (N_15297,N_9573,N_11348);
nand U15298 (N_15298,N_11124,N_12067);
nor U15299 (N_15299,N_11573,N_11282);
and U15300 (N_15300,N_12448,N_11188);
xnor U15301 (N_15301,N_9778,N_10426);
nor U15302 (N_15302,N_11012,N_9894);
and U15303 (N_15303,N_11854,N_11363);
nor U15304 (N_15304,N_9798,N_12378);
nand U15305 (N_15305,N_9974,N_9403);
or U15306 (N_15306,N_10570,N_12197);
and U15307 (N_15307,N_10246,N_11550);
or U15308 (N_15308,N_10996,N_9421);
or U15309 (N_15309,N_12467,N_11185);
or U15310 (N_15310,N_11890,N_10964);
xor U15311 (N_15311,N_12081,N_11186);
nand U15312 (N_15312,N_9749,N_10763);
and U15313 (N_15313,N_11061,N_10987);
nand U15314 (N_15314,N_11276,N_9426);
or U15315 (N_15315,N_9852,N_10658);
or U15316 (N_15316,N_10441,N_12086);
or U15317 (N_15317,N_11723,N_11697);
or U15318 (N_15318,N_11153,N_10058);
nor U15319 (N_15319,N_12448,N_12337);
nand U15320 (N_15320,N_10833,N_10725);
or U15321 (N_15321,N_12441,N_10680);
xnor U15322 (N_15322,N_11518,N_12408);
nand U15323 (N_15323,N_12018,N_10955);
or U15324 (N_15324,N_10333,N_11253);
nand U15325 (N_15325,N_10691,N_10133);
or U15326 (N_15326,N_10695,N_9664);
or U15327 (N_15327,N_10879,N_11450);
or U15328 (N_15328,N_10343,N_11593);
and U15329 (N_15329,N_12113,N_11694);
nor U15330 (N_15330,N_10354,N_10045);
nor U15331 (N_15331,N_12486,N_12195);
nand U15332 (N_15332,N_11713,N_9667);
and U15333 (N_15333,N_10711,N_10544);
nand U15334 (N_15334,N_10507,N_10170);
or U15335 (N_15335,N_9809,N_10059);
nand U15336 (N_15336,N_10351,N_10866);
nand U15337 (N_15337,N_11416,N_10945);
nor U15338 (N_15338,N_10971,N_12264);
and U15339 (N_15339,N_9783,N_10232);
nand U15340 (N_15340,N_10351,N_12172);
or U15341 (N_15341,N_10088,N_10301);
and U15342 (N_15342,N_10122,N_11429);
xnor U15343 (N_15343,N_11581,N_10093);
nand U15344 (N_15344,N_10284,N_10184);
and U15345 (N_15345,N_11732,N_9468);
xor U15346 (N_15346,N_11726,N_9973);
and U15347 (N_15347,N_9943,N_11208);
xor U15348 (N_15348,N_10787,N_12359);
or U15349 (N_15349,N_9600,N_12004);
or U15350 (N_15350,N_10410,N_9436);
nand U15351 (N_15351,N_11890,N_12309);
nand U15352 (N_15352,N_10874,N_11510);
nor U15353 (N_15353,N_10690,N_11363);
nand U15354 (N_15354,N_12246,N_10340);
and U15355 (N_15355,N_10744,N_10285);
xnor U15356 (N_15356,N_11412,N_10049);
and U15357 (N_15357,N_10223,N_11173);
and U15358 (N_15358,N_10616,N_9544);
nor U15359 (N_15359,N_11065,N_9903);
nand U15360 (N_15360,N_10053,N_10374);
xor U15361 (N_15361,N_11350,N_12432);
nor U15362 (N_15362,N_9678,N_12494);
or U15363 (N_15363,N_10052,N_10351);
or U15364 (N_15364,N_11759,N_10420);
and U15365 (N_15365,N_9590,N_11502);
or U15366 (N_15366,N_11724,N_10689);
and U15367 (N_15367,N_10054,N_9427);
or U15368 (N_15368,N_9546,N_10155);
or U15369 (N_15369,N_11078,N_11532);
nor U15370 (N_15370,N_12105,N_10962);
xnor U15371 (N_15371,N_12335,N_10710);
nor U15372 (N_15372,N_10141,N_9529);
or U15373 (N_15373,N_12293,N_10588);
and U15374 (N_15374,N_10513,N_10658);
and U15375 (N_15375,N_11374,N_11035);
nand U15376 (N_15376,N_10951,N_11971);
nor U15377 (N_15377,N_11260,N_11586);
or U15378 (N_15378,N_10538,N_10246);
xor U15379 (N_15379,N_10338,N_9592);
or U15380 (N_15380,N_10744,N_10267);
and U15381 (N_15381,N_11999,N_10657);
nor U15382 (N_15382,N_11321,N_9664);
nor U15383 (N_15383,N_10020,N_9468);
and U15384 (N_15384,N_11652,N_11333);
and U15385 (N_15385,N_9906,N_9458);
and U15386 (N_15386,N_11382,N_11051);
and U15387 (N_15387,N_10334,N_11285);
nand U15388 (N_15388,N_12278,N_12175);
nand U15389 (N_15389,N_10011,N_11545);
xnor U15390 (N_15390,N_12354,N_11697);
xor U15391 (N_15391,N_9828,N_11544);
nor U15392 (N_15392,N_10137,N_9818);
and U15393 (N_15393,N_11475,N_9439);
nand U15394 (N_15394,N_10686,N_10757);
xnor U15395 (N_15395,N_12397,N_12114);
or U15396 (N_15396,N_10693,N_9846);
nand U15397 (N_15397,N_11859,N_12259);
and U15398 (N_15398,N_10260,N_9885);
nor U15399 (N_15399,N_9658,N_11164);
xnor U15400 (N_15400,N_10070,N_9870);
or U15401 (N_15401,N_9451,N_11887);
and U15402 (N_15402,N_10325,N_11196);
nand U15403 (N_15403,N_10586,N_10438);
or U15404 (N_15404,N_11708,N_10345);
nand U15405 (N_15405,N_12120,N_10197);
and U15406 (N_15406,N_11220,N_12446);
nand U15407 (N_15407,N_9613,N_12125);
xnor U15408 (N_15408,N_11661,N_11162);
and U15409 (N_15409,N_12138,N_10049);
and U15410 (N_15410,N_10522,N_11839);
nor U15411 (N_15411,N_10723,N_10358);
and U15412 (N_15412,N_10396,N_12225);
and U15413 (N_15413,N_11246,N_12044);
nor U15414 (N_15414,N_11860,N_10856);
and U15415 (N_15415,N_11609,N_10939);
nand U15416 (N_15416,N_9512,N_10438);
nand U15417 (N_15417,N_9781,N_10056);
nand U15418 (N_15418,N_12047,N_11360);
or U15419 (N_15419,N_9939,N_11199);
xor U15420 (N_15420,N_10791,N_9646);
nor U15421 (N_15421,N_11652,N_11666);
nor U15422 (N_15422,N_10118,N_11180);
nor U15423 (N_15423,N_9992,N_12440);
nor U15424 (N_15424,N_9959,N_12031);
or U15425 (N_15425,N_10759,N_10435);
nor U15426 (N_15426,N_10955,N_11248);
and U15427 (N_15427,N_9456,N_11544);
or U15428 (N_15428,N_9675,N_10242);
and U15429 (N_15429,N_10875,N_9895);
nand U15430 (N_15430,N_10019,N_10622);
nor U15431 (N_15431,N_12026,N_10197);
or U15432 (N_15432,N_9520,N_11229);
nand U15433 (N_15433,N_10962,N_9555);
xnor U15434 (N_15434,N_11960,N_9520);
xnor U15435 (N_15435,N_11848,N_12138);
nor U15436 (N_15436,N_11694,N_12066);
or U15437 (N_15437,N_10646,N_12168);
and U15438 (N_15438,N_12248,N_11208);
nand U15439 (N_15439,N_10914,N_12469);
nor U15440 (N_15440,N_9392,N_11091);
and U15441 (N_15441,N_9587,N_11232);
nand U15442 (N_15442,N_10994,N_11656);
or U15443 (N_15443,N_12302,N_10537);
and U15444 (N_15444,N_11348,N_11246);
and U15445 (N_15445,N_10587,N_9544);
nand U15446 (N_15446,N_10379,N_12101);
and U15447 (N_15447,N_11648,N_12308);
or U15448 (N_15448,N_12300,N_11166);
nand U15449 (N_15449,N_10808,N_10066);
nor U15450 (N_15450,N_9453,N_12034);
or U15451 (N_15451,N_9713,N_9413);
or U15452 (N_15452,N_12037,N_12046);
or U15453 (N_15453,N_10751,N_12354);
or U15454 (N_15454,N_10310,N_11412);
or U15455 (N_15455,N_12428,N_11133);
xor U15456 (N_15456,N_9603,N_10813);
nor U15457 (N_15457,N_10836,N_12424);
or U15458 (N_15458,N_10940,N_11386);
xnor U15459 (N_15459,N_9630,N_12057);
nor U15460 (N_15460,N_10310,N_10529);
or U15461 (N_15461,N_9717,N_12483);
and U15462 (N_15462,N_9608,N_9724);
xnor U15463 (N_15463,N_12237,N_12118);
nor U15464 (N_15464,N_11133,N_11708);
and U15465 (N_15465,N_9793,N_11944);
nand U15466 (N_15466,N_12225,N_11470);
or U15467 (N_15467,N_11803,N_9918);
and U15468 (N_15468,N_10886,N_10315);
and U15469 (N_15469,N_9594,N_11190);
or U15470 (N_15470,N_9795,N_12282);
nor U15471 (N_15471,N_11744,N_10632);
nand U15472 (N_15472,N_9380,N_12208);
and U15473 (N_15473,N_11216,N_10203);
and U15474 (N_15474,N_10374,N_12067);
and U15475 (N_15475,N_9799,N_10973);
and U15476 (N_15476,N_11797,N_11094);
nand U15477 (N_15477,N_10067,N_10424);
xor U15478 (N_15478,N_11752,N_9701);
xor U15479 (N_15479,N_12161,N_12187);
and U15480 (N_15480,N_12220,N_10460);
nand U15481 (N_15481,N_11815,N_10195);
and U15482 (N_15482,N_11496,N_11181);
or U15483 (N_15483,N_11809,N_10295);
or U15484 (N_15484,N_12313,N_11320);
xor U15485 (N_15485,N_9960,N_10102);
xnor U15486 (N_15486,N_9443,N_9936);
nand U15487 (N_15487,N_11135,N_11892);
and U15488 (N_15488,N_10462,N_10722);
nor U15489 (N_15489,N_11294,N_10836);
nor U15490 (N_15490,N_10951,N_11799);
and U15491 (N_15491,N_12289,N_12498);
xnor U15492 (N_15492,N_12477,N_9481);
nand U15493 (N_15493,N_12187,N_11916);
nand U15494 (N_15494,N_10936,N_10125);
nand U15495 (N_15495,N_10450,N_12440);
nor U15496 (N_15496,N_9999,N_9589);
or U15497 (N_15497,N_10969,N_10463);
nor U15498 (N_15498,N_10748,N_11253);
or U15499 (N_15499,N_11502,N_10862);
xor U15500 (N_15500,N_10826,N_9898);
or U15501 (N_15501,N_10829,N_11210);
or U15502 (N_15502,N_10094,N_10604);
nor U15503 (N_15503,N_10498,N_11541);
and U15504 (N_15504,N_12369,N_10942);
nor U15505 (N_15505,N_10643,N_9740);
and U15506 (N_15506,N_10891,N_10124);
nor U15507 (N_15507,N_12036,N_11921);
or U15508 (N_15508,N_12252,N_9688);
and U15509 (N_15509,N_11902,N_10989);
nand U15510 (N_15510,N_9880,N_10218);
nand U15511 (N_15511,N_10038,N_10210);
nor U15512 (N_15512,N_10305,N_10137);
and U15513 (N_15513,N_9769,N_12339);
or U15514 (N_15514,N_12410,N_10730);
and U15515 (N_15515,N_12280,N_9575);
nor U15516 (N_15516,N_12163,N_9902);
and U15517 (N_15517,N_10944,N_11978);
xor U15518 (N_15518,N_10169,N_9771);
nand U15519 (N_15519,N_11061,N_11992);
or U15520 (N_15520,N_12052,N_11458);
nor U15521 (N_15521,N_12127,N_11799);
nor U15522 (N_15522,N_11748,N_10264);
or U15523 (N_15523,N_11263,N_10653);
nor U15524 (N_15524,N_9673,N_9411);
nor U15525 (N_15525,N_11966,N_12467);
and U15526 (N_15526,N_10001,N_10135);
xnor U15527 (N_15527,N_9958,N_10442);
and U15528 (N_15528,N_11209,N_11535);
or U15529 (N_15529,N_11864,N_11204);
and U15530 (N_15530,N_11867,N_10632);
or U15531 (N_15531,N_10963,N_12032);
nor U15532 (N_15532,N_12185,N_11052);
or U15533 (N_15533,N_11958,N_9713);
or U15534 (N_15534,N_11723,N_10452);
or U15535 (N_15535,N_9941,N_9879);
or U15536 (N_15536,N_9848,N_11078);
or U15537 (N_15537,N_11831,N_11863);
nand U15538 (N_15538,N_11421,N_11503);
or U15539 (N_15539,N_11778,N_11341);
or U15540 (N_15540,N_10227,N_12003);
nor U15541 (N_15541,N_12279,N_12118);
xor U15542 (N_15542,N_11891,N_11101);
or U15543 (N_15543,N_9686,N_9981);
nand U15544 (N_15544,N_10662,N_10996);
nand U15545 (N_15545,N_9488,N_9544);
nand U15546 (N_15546,N_11476,N_10884);
or U15547 (N_15547,N_9912,N_11084);
and U15548 (N_15548,N_11020,N_9993);
and U15549 (N_15549,N_10391,N_11193);
or U15550 (N_15550,N_10890,N_10362);
or U15551 (N_15551,N_10230,N_11143);
and U15552 (N_15552,N_11873,N_9802);
and U15553 (N_15553,N_11311,N_11654);
nand U15554 (N_15554,N_10579,N_11603);
or U15555 (N_15555,N_11468,N_12000);
and U15556 (N_15556,N_9887,N_10632);
or U15557 (N_15557,N_11165,N_9607);
nand U15558 (N_15558,N_9563,N_9775);
nor U15559 (N_15559,N_11415,N_10620);
xnor U15560 (N_15560,N_10619,N_12043);
or U15561 (N_15561,N_9435,N_11098);
nand U15562 (N_15562,N_9580,N_9385);
nand U15563 (N_15563,N_11205,N_10430);
or U15564 (N_15564,N_11554,N_11391);
nand U15565 (N_15565,N_10076,N_10971);
and U15566 (N_15566,N_12197,N_11715);
or U15567 (N_15567,N_10020,N_12324);
and U15568 (N_15568,N_11675,N_9383);
nor U15569 (N_15569,N_12157,N_10831);
nor U15570 (N_15570,N_10293,N_10379);
nor U15571 (N_15571,N_10705,N_12139);
nor U15572 (N_15572,N_9779,N_10880);
xor U15573 (N_15573,N_12369,N_11791);
and U15574 (N_15574,N_11010,N_9594);
and U15575 (N_15575,N_11423,N_10991);
and U15576 (N_15576,N_12251,N_11458);
nor U15577 (N_15577,N_11261,N_12226);
and U15578 (N_15578,N_11702,N_12133);
nand U15579 (N_15579,N_9609,N_9752);
and U15580 (N_15580,N_10816,N_10967);
nand U15581 (N_15581,N_10166,N_9457);
or U15582 (N_15582,N_10480,N_10041);
and U15583 (N_15583,N_10162,N_11301);
and U15584 (N_15584,N_12019,N_9783);
and U15585 (N_15585,N_9506,N_9831);
nand U15586 (N_15586,N_11165,N_10908);
xor U15587 (N_15587,N_10958,N_11400);
and U15588 (N_15588,N_10293,N_11874);
xor U15589 (N_15589,N_11036,N_9878);
and U15590 (N_15590,N_10551,N_11540);
and U15591 (N_15591,N_12195,N_10654);
xor U15592 (N_15592,N_12051,N_9910);
xor U15593 (N_15593,N_12030,N_10565);
or U15594 (N_15594,N_12412,N_10536);
nand U15595 (N_15595,N_12032,N_10886);
and U15596 (N_15596,N_9474,N_10688);
or U15597 (N_15597,N_12425,N_9647);
nor U15598 (N_15598,N_10835,N_12202);
nand U15599 (N_15599,N_11388,N_10000);
nand U15600 (N_15600,N_9696,N_9883);
nor U15601 (N_15601,N_9521,N_9532);
xnor U15602 (N_15602,N_12081,N_9861);
or U15603 (N_15603,N_10723,N_10326);
nor U15604 (N_15604,N_11065,N_11195);
nor U15605 (N_15605,N_10544,N_11792);
nand U15606 (N_15606,N_10783,N_10516);
and U15607 (N_15607,N_12043,N_9648);
and U15608 (N_15608,N_10414,N_11641);
and U15609 (N_15609,N_10571,N_10719);
nor U15610 (N_15610,N_11257,N_9504);
nand U15611 (N_15611,N_10141,N_12314);
or U15612 (N_15612,N_9905,N_12384);
xnor U15613 (N_15613,N_10514,N_12146);
nand U15614 (N_15614,N_12461,N_10801);
or U15615 (N_15615,N_10245,N_11502);
xor U15616 (N_15616,N_11562,N_11827);
or U15617 (N_15617,N_11156,N_10908);
nand U15618 (N_15618,N_11721,N_9876);
nand U15619 (N_15619,N_10216,N_9528);
nor U15620 (N_15620,N_11588,N_12436);
nor U15621 (N_15621,N_9707,N_9926);
and U15622 (N_15622,N_12120,N_11020);
nand U15623 (N_15623,N_12433,N_9576);
or U15624 (N_15624,N_10194,N_11953);
nand U15625 (N_15625,N_14750,N_13712);
and U15626 (N_15626,N_13681,N_14809);
or U15627 (N_15627,N_14831,N_14840);
and U15628 (N_15628,N_12828,N_14911);
xnor U15629 (N_15629,N_14500,N_13255);
xor U15630 (N_15630,N_13991,N_14100);
nand U15631 (N_15631,N_13131,N_13191);
nand U15632 (N_15632,N_13002,N_13720);
nor U15633 (N_15633,N_14742,N_12882);
and U15634 (N_15634,N_12755,N_15416);
and U15635 (N_15635,N_13062,N_15291);
xor U15636 (N_15636,N_15282,N_14618);
nand U15637 (N_15637,N_15349,N_14067);
or U15638 (N_15638,N_14283,N_13007);
and U15639 (N_15639,N_14166,N_14926);
or U15640 (N_15640,N_15205,N_13160);
or U15641 (N_15641,N_13377,N_13960);
or U15642 (N_15642,N_13560,N_14585);
nor U15643 (N_15643,N_15413,N_15065);
nand U15644 (N_15644,N_15119,N_12660);
xnor U15645 (N_15645,N_12791,N_14123);
xnor U15646 (N_15646,N_14049,N_13253);
and U15647 (N_15647,N_14807,N_13888);
nor U15648 (N_15648,N_14076,N_14886);
or U15649 (N_15649,N_13107,N_13153);
xor U15650 (N_15650,N_15490,N_13737);
and U15651 (N_15651,N_13981,N_14428);
nor U15652 (N_15652,N_12519,N_14765);
or U15653 (N_15653,N_14939,N_12824);
and U15654 (N_15654,N_14838,N_13868);
nand U15655 (N_15655,N_12780,N_13613);
and U15656 (N_15656,N_14091,N_14322);
and U15657 (N_15657,N_13413,N_13741);
or U15658 (N_15658,N_15058,N_12798);
nand U15659 (N_15659,N_15312,N_15584);
nor U15660 (N_15660,N_12956,N_13992);
or U15661 (N_15661,N_12769,N_13945);
nand U15662 (N_15662,N_13100,N_13300);
nor U15663 (N_15663,N_13566,N_15043);
and U15664 (N_15664,N_12732,N_14480);
or U15665 (N_15665,N_14977,N_15050);
or U15666 (N_15666,N_13341,N_12700);
nor U15667 (N_15667,N_12794,N_12931);
xnor U15668 (N_15668,N_13826,N_13400);
and U15669 (N_15669,N_14569,N_13680);
xor U15670 (N_15670,N_15087,N_14203);
nor U15671 (N_15671,N_15259,N_15225);
and U15672 (N_15672,N_14142,N_14376);
nand U15673 (N_15673,N_13420,N_13169);
xnor U15674 (N_15674,N_15038,N_15488);
nand U15675 (N_15675,N_13573,N_13864);
or U15676 (N_15676,N_15027,N_14698);
nor U15677 (N_15677,N_14429,N_12616);
nand U15678 (N_15678,N_15367,N_15275);
or U15679 (N_15679,N_12864,N_15609);
or U15680 (N_15680,N_14760,N_14217);
and U15681 (N_15681,N_13662,N_14921);
and U15682 (N_15682,N_15333,N_14969);
and U15683 (N_15683,N_14941,N_13527);
nand U15684 (N_15684,N_12622,N_12986);
or U15685 (N_15685,N_15622,N_14487);
nor U15686 (N_15686,N_14726,N_15323);
nand U15687 (N_15687,N_13044,N_12944);
and U15688 (N_15688,N_13504,N_12895);
nand U15689 (N_15689,N_15324,N_14413);
and U15690 (N_15690,N_14804,N_14806);
nand U15691 (N_15691,N_14292,N_14632);
nor U15692 (N_15692,N_12516,N_14472);
nor U15693 (N_15693,N_13308,N_14277);
or U15694 (N_15694,N_13006,N_14630);
nand U15695 (N_15695,N_15453,N_14826);
nand U15696 (N_15696,N_14562,N_13542);
nand U15697 (N_15697,N_14415,N_15115);
nor U15698 (N_15698,N_12726,N_13201);
or U15699 (N_15699,N_13302,N_14419);
nand U15700 (N_15700,N_13805,N_13637);
and U15701 (N_15701,N_13550,N_13880);
or U15702 (N_15702,N_15497,N_13128);
nor U15703 (N_15703,N_15507,N_12859);
and U15704 (N_15704,N_14973,N_15605);
nor U15705 (N_15705,N_15222,N_15154);
nand U15706 (N_15706,N_14959,N_14930);
nor U15707 (N_15707,N_14770,N_15097);
nand U15708 (N_15708,N_15098,N_14286);
or U15709 (N_15709,N_13005,N_15239);
and U15710 (N_15710,N_13225,N_15041);
nand U15711 (N_15711,N_15136,N_15163);
xor U15712 (N_15712,N_14207,N_15051);
nand U15713 (N_15713,N_14477,N_12572);
nand U15714 (N_15714,N_12666,N_12910);
and U15715 (N_15715,N_15219,N_13611);
xor U15716 (N_15716,N_13823,N_13551);
nand U15717 (N_15717,N_12655,N_12647);
or U15718 (N_15718,N_15227,N_15019);
and U15719 (N_15719,N_14178,N_13596);
nand U15720 (N_15720,N_13948,N_14512);
nand U15721 (N_15721,N_14176,N_13111);
or U15722 (N_15722,N_13310,N_13439);
and U15723 (N_15723,N_14025,N_13523);
and U15724 (N_15724,N_14241,N_15621);
nor U15725 (N_15725,N_13097,N_12809);
nand U15726 (N_15726,N_15195,N_13961);
and U15727 (N_15727,N_13029,N_15101);
or U15728 (N_15728,N_15574,N_15194);
nand U15729 (N_15729,N_14783,N_13250);
xnor U15730 (N_15730,N_15140,N_13059);
or U15731 (N_15731,N_13451,N_14738);
nand U15732 (N_15732,N_15352,N_14334);
or U15733 (N_15733,N_13399,N_14368);
and U15734 (N_15734,N_12881,N_12969);
nor U15735 (N_15735,N_12712,N_14771);
nand U15736 (N_15736,N_15573,N_13430);
nor U15737 (N_15737,N_13429,N_13236);
nor U15738 (N_15738,N_15066,N_15387);
nor U15739 (N_15739,N_13033,N_12695);
and U15740 (N_15740,N_14436,N_14904);
nor U15741 (N_15741,N_12518,N_15358);
and U15742 (N_15742,N_15072,N_13232);
or U15743 (N_15743,N_14737,N_12515);
nand U15744 (N_15744,N_13353,N_13455);
and U15745 (N_15745,N_13277,N_12933);
nand U15746 (N_15746,N_14159,N_15280);
or U15747 (N_15747,N_12941,N_12634);
or U15748 (N_15748,N_14645,N_13478);
nand U15749 (N_15749,N_13132,N_15410);
and U15750 (N_15750,N_13791,N_13505);
nor U15751 (N_15751,N_13821,N_14307);
nor U15752 (N_15752,N_14578,N_14200);
and U15753 (N_15753,N_12520,N_13363);
and U15754 (N_15754,N_13866,N_12987);
nand U15755 (N_15755,N_13477,N_13386);
and U15756 (N_15756,N_14229,N_13344);
or U15757 (N_15757,N_14206,N_13103);
or U15758 (N_15758,N_13075,N_12597);
and U15759 (N_15759,N_15515,N_14346);
and U15760 (N_15760,N_15471,N_15336);
nand U15761 (N_15761,N_13806,N_13606);
and U15762 (N_15762,N_13528,N_14410);
nand U15763 (N_15763,N_13301,N_14719);
nor U15764 (N_15764,N_12583,N_13954);
and U15765 (N_15765,N_14414,N_12584);
and U15766 (N_15766,N_15343,N_12522);
or U15767 (N_15767,N_13142,N_15363);
and U15768 (N_15768,N_13395,N_14493);
nor U15769 (N_15769,N_15171,N_14045);
and U15770 (N_15770,N_14314,N_12723);
xor U15771 (N_15771,N_14834,N_15328);
or U15772 (N_15772,N_14185,N_14172);
or U15773 (N_15773,N_14733,N_13284);
nor U15774 (N_15774,N_15448,N_13633);
or U15775 (N_15775,N_12704,N_13503);
or U15776 (N_15776,N_14367,N_12635);
and U15777 (N_15777,N_14273,N_12534);
nand U15778 (N_15778,N_14441,N_14701);
or U15779 (N_15779,N_14496,N_15204);
and U15780 (N_15780,N_12966,N_14985);
nor U15781 (N_15781,N_15612,N_14626);
nor U15782 (N_15782,N_15499,N_14666);
or U15783 (N_15783,N_15304,N_13348);
nor U15784 (N_15784,N_12889,N_15421);
nor U15785 (N_15785,N_13946,N_13089);
nor U15786 (N_15786,N_12974,N_12811);
nand U15787 (N_15787,N_15217,N_12668);
or U15788 (N_15788,N_14749,N_14530);
nand U15789 (N_15789,N_14942,N_15524);
nor U15790 (N_15790,N_12883,N_14946);
or U15791 (N_15791,N_15257,N_14563);
nor U15792 (N_15792,N_15451,N_13718);
or U15793 (N_15793,N_13229,N_15380);
nand U15794 (N_15794,N_14317,N_15435);
and U15795 (N_15795,N_15116,N_15583);
nor U15796 (N_15796,N_13815,N_15577);
nor U15797 (N_15797,N_15110,N_13994);
nor U15798 (N_15798,N_12642,N_14196);
and U15799 (N_15799,N_14581,N_14315);
and U15800 (N_15800,N_15457,N_15001);
nor U15801 (N_15801,N_15289,N_13622);
xor U15802 (N_15802,N_13355,N_12761);
nand U15803 (N_15803,N_13583,N_13997);
nand U15804 (N_15804,N_12528,N_13786);
or U15805 (N_15805,N_13749,N_15408);
nand U15806 (N_15806,N_13247,N_12678);
xor U15807 (N_15807,N_13862,N_14976);
nor U15808 (N_15808,N_14002,N_13246);
and U15809 (N_15809,N_13627,N_13565);
xor U15810 (N_15810,N_14192,N_14422);
nor U15811 (N_15811,N_14316,N_14556);
nand U15812 (N_15812,N_14224,N_15350);
xor U15813 (N_15813,N_12722,N_12682);
or U15814 (N_15814,N_15330,N_13979);
or U15815 (N_15815,N_14888,N_13393);
nor U15816 (N_15816,N_13574,N_13397);
nor U15817 (N_15817,N_14381,N_13704);
nor U15818 (N_15818,N_14427,N_15486);
or U15819 (N_15819,N_12595,N_13022);
nor U15820 (N_15820,N_14366,N_14109);
or U15821 (N_15821,N_12759,N_14731);
or U15822 (N_15822,N_13687,N_13714);
and U15823 (N_15823,N_15519,N_13155);
or U15824 (N_15824,N_13540,N_12801);
and U15825 (N_15825,N_14495,N_15587);
or U15826 (N_15826,N_13423,N_13019);
nand U15827 (N_15827,N_15080,N_13011);
nor U15828 (N_15828,N_15551,N_14380);
nand U15829 (N_15829,N_14160,N_14812);
or U15830 (N_15830,N_15474,N_13846);
and U15831 (N_15831,N_12803,N_14994);
or U15832 (N_15832,N_15062,N_12782);
and U15833 (N_15833,N_12554,N_15203);
or U15834 (N_15834,N_14681,N_12550);
nand U15835 (N_15835,N_14327,N_13244);
and U15836 (N_15836,N_13999,N_13539);
nor U15837 (N_15837,N_15395,N_14654);
and U15838 (N_15838,N_14670,N_14041);
nor U15839 (N_15839,N_12650,N_13489);
and U15840 (N_15840,N_14873,N_14132);
nand U15841 (N_15841,N_14915,N_13577);
nor U15842 (N_15842,N_14340,N_14245);
xnor U15843 (N_15843,N_14538,N_12989);
nand U15844 (N_15844,N_13218,N_14794);
nand U15845 (N_15845,N_12837,N_12991);
nor U15846 (N_15846,N_14125,N_14387);
nand U15847 (N_15847,N_13904,N_15060);
or U15848 (N_15848,N_15522,N_15238);
or U15849 (N_15849,N_13522,N_13116);
and U15850 (N_15850,N_12939,N_15268);
nor U15851 (N_15851,N_15420,N_14488);
and U15852 (N_15852,N_15037,N_12860);
and U15853 (N_15853,N_14161,N_15183);
or U15854 (N_15854,N_15005,N_12654);
or U15855 (N_15855,N_15105,N_12885);
nand U15856 (N_15856,N_14405,N_13570);
nor U15857 (N_15857,N_12898,N_12905);
xnor U15858 (N_15858,N_15530,N_12506);
or U15859 (N_15859,N_12839,N_13849);
nor U15860 (N_15860,N_14408,N_12822);
and U15861 (N_15861,N_12651,N_12850);
xnor U15862 (N_15862,N_14099,N_13870);
or U15863 (N_15863,N_13502,N_15618);
nand U15864 (N_15864,N_14631,N_15290);
nand U15865 (N_15865,N_15196,N_13211);
or U15866 (N_15866,N_15517,N_14964);
nor U15867 (N_15867,N_14301,N_12915);
nand U15868 (N_15868,N_13289,N_12664);
or U15869 (N_15869,N_14583,N_14655);
nand U15870 (N_15870,N_12596,N_15186);
nand U15871 (N_15871,N_14174,N_13985);
or U15872 (N_15872,N_14846,N_14059);
nor U15873 (N_15873,N_14110,N_13143);
xnor U15874 (N_15874,N_13578,N_12861);
and U15875 (N_15875,N_13316,N_13857);
nand U15876 (N_15876,N_14186,N_12832);
or U15877 (N_15877,N_15153,N_13015);
nor U15878 (N_15878,N_13449,N_14096);
nand U15879 (N_15879,N_13444,N_14332);
xnor U15880 (N_15880,N_14430,N_12566);
or U15881 (N_15881,N_15120,N_12698);
xor U15882 (N_15882,N_14763,N_13709);
or U15883 (N_15883,N_14248,N_12767);
nor U15884 (N_15884,N_13674,N_15306);
nor U15885 (N_15885,N_12621,N_15412);
nor U15886 (N_15886,N_15295,N_13372);
and U15887 (N_15887,N_13711,N_15372);
nand U15888 (N_15888,N_14171,N_14080);
or U15889 (N_15889,N_12745,N_14594);
nand U15890 (N_15890,N_14362,N_13165);
xor U15891 (N_15891,N_13485,N_15309);
nor U15892 (N_15892,N_12632,N_14335);
and U15893 (N_15893,N_13224,N_14648);
or U15894 (N_15894,N_12836,N_14054);
xor U15895 (N_15895,N_12897,N_14111);
nand U15896 (N_15896,N_13668,N_14086);
nand U15897 (N_15897,N_12526,N_14385);
nor U15898 (N_15898,N_12976,N_15033);
nor U15899 (N_15899,N_14398,N_14146);
and U15900 (N_15900,N_15025,N_12979);
or U15901 (N_15901,N_12667,N_13079);
xor U15902 (N_15902,N_13313,N_13299);
nor U15903 (N_15903,N_15461,N_15447);
nand U15904 (N_15904,N_13739,N_12605);
and U15905 (N_15905,N_12901,N_14958);
nand U15906 (N_15906,N_12693,N_14453);
and U15907 (N_15907,N_13392,N_14850);
and U15908 (N_15908,N_13258,N_12725);
nand U15909 (N_15909,N_13947,N_13438);
nand U15910 (N_15910,N_12948,N_15265);
nor U15911 (N_15911,N_14633,N_15279);
or U15912 (N_15912,N_14392,N_13819);
nor U15913 (N_15913,N_13661,N_15093);
and U15914 (N_15914,N_15071,N_13631);
and U15915 (N_15915,N_13366,N_13669);
and U15916 (N_15916,N_13604,N_13157);
and U15917 (N_15917,N_13352,N_15307);
nand U15918 (N_15918,N_13831,N_13426);
nand U15919 (N_15919,N_14421,N_12747);
or U15920 (N_15920,N_13434,N_12512);
nor U15921 (N_15921,N_15270,N_14247);
nand U15922 (N_15922,N_12936,N_13350);
xor U15923 (N_15923,N_14072,N_14044);
nand U15924 (N_15924,N_15294,N_14966);
nand U15925 (N_15925,N_14156,N_15250);
or U15926 (N_15926,N_15042,N_14869);
nand U15927 (N_15927,N_15595,N_13073);
and U15928 (N_15928,N_12753,N_15539);
nand U15929 (N_15929,N_13521,N_14906);
or U15930 (N_15930,N_14817,N_13548);
and U15931 (N_15931,N_12517,N_13421);
xor U15932 (N_15932,N_13388,N_13963);
or U15933 (N_15933,N_13779,N_13648);
nor U15934 (N_15934,N_14908,N_12551);
nand U15935 (N_15935,N_14784,N_13513);
nand U15936 (N_15936,N_12752,N_13199);
xnor U15937 (N_15937,N_13964,N_15516);
or U15938 (N_15938,N_13973,N_13561);
nand U15939 (N_15939,N_13281,N_12617);
nand U15940 (N_15940,N_13891,N_14900);
and U15941 (N_15941,N_14511,N_15494);
and U15942 (N_15942,N_14732,N_15357);
nor U15943 (N_15943,N_13480,N_15468);
nor U15944 (N_15944,N_14523,N_13555);
and U15945 (N_15945,N_12705,N_13892);
nand U15946 (N_15946,N_15181,N_12615);
nand U15947 (N_15947,N_14395,N_14490);
and U15948 (N_15948,N_14257,N_14865);
nand U15949 (N_15949,N_14127,N_13018);
and U15950 (N_15950,N_14043,N_14550);
or U15951 (N_15951,N_13235,N_14280);
or U15952 (N_15952,N_13328,N_12645);
nor U15953 (N_15953,N_15017,N_14276);
nand U15954 (N_15954,N_14394,N_15178);
xor U15955 (N_15955,N_13329,N_15068);
nand U15956 (N_15956,N_13181,N_13178);
or U15957 (N_15957,N_12980,N_13203);
nand U15958 (N_15958,N_14117,N_14008);
or U15959 (N_15959,N_12541,N_13252);
nand U15960 (N_15960,N_14333,N_13861);
or U15961 (N_15961,N_12781,N_12906);
nor U15962 (N_15962,N_15582,N_12532);
nand U15963 (N_15963,N_14062,N_13544);
nand U15964 (N_15964,N_13042,N_13156);
xnor U15965 (N_15965,N_15271,N_14916);
or U15966 (N_15966,N_13304,N_14378);
nand U15967 (N_15967,N_12786,N_15292);
nor U15968 (N_15968,N_13335,N_14236);
nand U15969 (N_15969,N_15190,N_12570);
nand U15970 (N_15970,N_13691,N_12751);
nand U15971 (N_15971,N_13698,N_13437);
nand U15972 (N_15972,N_15370,N_12644);
nor U15973 (N_15973,N_14897,N_12802);
or U15974 (N_15974,N_14862,N_14154);
and U15975 (N_15975,N_13916,N_14485);
nor U15976 (N_15976,N_13251,N_14695);
nor U15977 (N_15977,N_14795,N_13008);
or U15978 (N_15978,N_12558,N_14505);
nor U15979 (N_15979,N_15607,N_12547);
nor U15980 (N_15980,N_14451,N_14092);
or U15981 (N_15981,N_15035,N_15018);
xor U15982 (N_15982,N_13220,N_15493);
and U15983 (N_15983,N_12739,N_15606);
and U15984 (N_15984,N_13068,N_14359);
or U15985 (N_15985,N_14087,N_15224);
nand U15986 (N_15986,N_15506,N_14450);
or U15987 (N_15987,N_15455,N_15212);
xor U15988 (N_15988,N_12639,N_13332);
nand U15989 (N_15989,N_13064,N_13931);
nor U15990 (N_15990,N_13345,N_15177);
or U15991 (N_15991,N_15202,N_14134);
nand U15992 (N_15992,N_13216,N_12686);
and U15993 (N_15993,N_14808,N_14202);
or U15994 (N_15994,N_15500,N_14815);
nand U15995 (N_15995,N_12907,N_14950);
nor U15996 (N_15996,N_13219,N_15123);
or U15997 (N_15997,N_12771,N_12638);
nand U15998 (N_15998,N_14949,N_14306);
nand U15999 (N_15999,N_13321,N_13780);
and U16000 (N_16000,N_13585,N_14252);
nand U16001 (N_16001,N_12869,N_14891);
or U16002 (N_16002,N_14882,N_12917);
nor U16003 (N_16003,N_14232,N_13415);
and U16004 (N_16004,N_15096,N_13307);
nor U16005 (N_16005,N_14691,N_14401);
nor U16006 (N_16006,N_15394,N_14352);
nor U16007 (N_16007,N_15089,N_14577);
and U16008 (N_16008,N_12649,N_14548);
and U16009 (N_16009,N_15597,N_13759);
nand U16010 (N_16010,N_14683,N_13569);
nand U16011 (N_16011,N_12810,N_12653);
nand U16012 (N_16012,N_13556,N_14153);
and U16013 (N_16013,N_15576,N_13884);
nand U16014 (N_16014,N_15274,N_13382);
and U16015 (N_16015,N_15130,N_15199);
nand U16016 (N_16016,N_15558,N_13001);
nand U16017 (N_16017,N_12524,N_14981);
nor U16018 (N_16018,N_14952,N_12934);
and U16019 (N_16019,N_13968,N_14766);
nor U16020 (N_16020,N_13259,N_12618);
or U16021 (N_16021,N_15317,N_14974);
and U16022 (N_16022,N_15541,N_13755);
nand U16023 (N_16023,N_15188,N_13678);
or U16024 (N_16024,N_15533,N_12961);
and U16025 (N_16025,N_13511,N_15392);
and U16026 (N_16026,N_15004,N_14879);
or U16027 (N_16027,N_13935,N_14098);
nor U16028 (N_16028,N_14272,N_13385);
and U16029 (N_16029,N_14601,N_12902);
or U16030 (N_16030,N_14761,N_14552);
and U16031 (N_16031,N_15546,N_14056);
nor U16032 (N_16032,N_12783,N_14874);
and U16033 (N_16033,N_15373,N_13056);
nand U16034 (N_16034,N_15272,N_13562);
nor U16035 (N_16035,N_13061,N_13898);
or U16036 (N_16036,N_15591,N_15319);
nor U16037 (N_16037,N_13164,N_15230);
xnor U16038 (N_16038,N_14227,N_13071);
and U16039 (N_16039,N_13282,N_13102);
nand U16040 (N_16040,N_13095,N_13693);
nor U16041 (N_16041,N_13695,N_12501);
and U16042 (N_16042,N_15300,N_12978);
and U16043 (N_16043,N_13510,N_13147);
nand U16044 (N_16044,N_12958,N_15189);
nand U16045 (N_16045,N_12560,N_15469);
nor U16046 (N_16046,N_14190,N_14905);
nand U16047 (N_16047,N_12932,N_15360);
and U16048 (N_16048,N_14607,N_14754);
nor U16049 (N_16049,N_12740,N_15327);
nand U16050 (N_16050,N_13257,N_15081);
nor U16051 (N_16051,N_13465,N_15103);
or U16052 (N_16052,N_14231,N_15059);
and U16053 (N_16053,N_13747,N_14599);
nand U16054 (N_16054,N_15525,N_15569);
nor U16055 (N_16055,N_13241,N_12904);
nor U16056 (N_16056,N_12947,N_13373);
nand U16057 (N_16057,N_14027,N_15090);
nand U16058 (N_16058,N_15131,N_13682);
or U16059 (N_16059,N_12750,N_14568);
xor U16060 (N_16060,N_14040,N_13266);
nor U16061 (N_16061,N_15462,N_14303);
and U16062 (N_16062,N_14845,N_14642);
xor U16063 (N_16063,N_15208,N_13590);
nor U16064 (N_16064,N_15179,N_14369);
nand U16065 (N_16065,N_13249,N_12831);
or U16066 (N_16066,N_15145,N_14254);
xnor U16067 (N_16067,N_13545,N_12999);
nand U16068 (N_16068,N_14011,N_15446);
and U16069 (N_16069,N_15366,N_15013);
nand U16070 (N_16070,N_13579,N_14844);
or U16071 (N_16071,N_15443,N_13358);
nand U16072 (N_16072,N_13376,N_14609);
xnor U16073 (N_16073,N_13696,N_15046);
or U16074 (N_16074,N_15207,N_14135);
nand U16075 (N_16075,N_14506,N_13324);
nand U16076 (N_16076,N_13899,N_14752);
nor U16077 (N_16077,N_13762,N_12533);
nand U16078 (N_16078,N_13336,N_13804);
xor U16079 (N_16079,N_15567,N_13978);
nand U16080 (N_16080,N_14069,N_15314);
nor U16081 (N_16081,N_15571,N_13853);
xor U16082 (N_16082,N_14122,N_12626);
and U16083 (N_16083,N_15389,N_13808);
and U16084 (N_16084,N_14225,N_12509);
nor U16085 (N_16085,N_15022,N_13845);
or U16086 (N_16086,N_14843,N_13656);
or U16087 (N_16087,N_15057,N_14788);
or U16088 (N_16088,N_13279,N_13614);
xor U16089 (N_16089,N_15564,N_13547);
or U16090 (N_16090,N_15579,N_13105);
nand U16091 (N_16091,N_13081,N_15094);
nor U16092 (N_16092,N_12876,N_13930);
nor U16093 (N_16093,N_12630,N_12641);
or U16094 (N_16094,N_13557,N_14435);
and U16095 (N_16095,N_15482,N_13863);
nand U16096 (N_16096,N_15470,N_13811);
xnor U16097 (N_16097,N_14996,N_15624);
nor U16098 (N_16098,N_13408,N_14289);
and U16099 (N_16099,N_14715,N_12922);
nor U16100 (N_16100,N_14491,N_13699);
or U16101 (N_16101,N_13077,N_14935);
nand U16102 (N_16102,N_13602,N_15256);
nand U16103 (N_16103,N_14400,N_15619);
and U16104 (N_16104,N_14169,N_13162);
nand U16105 (N_16105,N_13063,N_13454);
and U16106 (N_16106,N_13516,N_12609);
or U16107 (N_16107,N_14465,N_15226);
nor U16108 (N_16108,N_13676,N_15426);
xnor U16109 (N_16109,N_13067,N_13151);
and U16110 (N_16110,N_13940,N_14084);
nor U16111 (N_16111,N_13146,N_13944);
nand U16112 (N_16112,N_12988,N_15472);
xor U16113 (N_16113,N_13655,N_15175);
nor U16114 (N_16114,N_13890,N_13784);
xor U16115 (N_16115,N_12692,N_14484);
and U16116 (N_16116,N_15234,N_13950);
or U16117 (N_16117,N_15449,N_15368);
and U16118 (N_16118,N_14866,N_15064);
and U16119 (N_16119,N_13688,N_15344);
or U16120 (N_16120,N_15377,N_12687);
nor U16121 (N_16121,N_13360,N_14309);
nor U16122 (N_16122,N_14081,N_12806);
and U16123 (N_16123,N_13198,N_14574);
xnor U16124 (N_16124,N_12815,N_14312);
and U16125 (N_16125,N_14519,N_12952);
nor U16126 (N_16126,N_13970,N_14532);
or U16127 (N_16127,N_13697,N_14211);
nand U16128 (N_16128,N_12880,N_13642);
and U16129 (N_16129,N_13529,N_15117);
nor U16130 (N_16130,N_14777,N_14553);
or U16131 (N_16131,N_15406,N_14576);
nand U16132 (N_16132,N_15559,N_14740);
nand U16133 (N_16133,N_14566,N_13893);
or U16134 (N_16134,N_13894,N_14282);
nand U16135 (N_16135,N_14650,N_15505);
nor U16136 (N_16136,N_12820,N_14205);
and U16137 (N_16137,N_14887,N_15374);
nor U16138 (N_16138,N_14739,N_13167);
nand U16139 (N_16139,N_15535,N_14718);
and U16140 (N_16140,N_14727,N_13070);
and U16141 (N_16141,N_13159,N_14048);
nand U16142 (N_16142,N_13756,N_13468);
and U16143 (N_16143,N_12586,N_14880);
nor U16144 (N_16144,N_15552,N_13708);
or U16145 (N_16145,N_14616,N_13957);
nor U16146 (N_16146,N_12993,N_13223);
or U16147 (N_16147,N_13854,N_15242);
xnor U16148 (N_16148,N_13689,N_15174);
nor U16149 (N_16149,N_15615,N_14640);
nor U16150 (N_16150,N_14945,N_12975);
nand U16151 (N_16151,N_14350,N_15254);
or U16152 (N_16152,N_15113,N_12717);
or U16153 (N_16153,N_14426,N_12770);
nor U16154 (N_16154,N_14249,N_15028);
xor U16155 (N_16155,N_13110,N_14223);
and U16156 (N_16156,N_14597,N_15463);
or U16157 (N_16157,N_13357,N_13524);
nand U16158 (N_16158,N_15241,N_13227);
and U16159 (N_16159,N_13326,N_12604);
nor U16160 (N_16160,N_14820,N_15548);
or U16161 (N_16161,N_12510,N_12858);
nand U16162 (N_16162,N_14722,N_13789);
nand U16163 (N_16163,N_15386,N_12743);
and U16164 (N_16164,N_13292,N_13125);
or U16165 (N_16165,N_12706,N_15402);
or U16166 (N_16166,N_14917,N_13190);
and U16167 (N_16167,N_14713,N_14012);
and U16168 (N_16168,N_13667,N_13280);
xnor U16169 (N_16169,N_13322,N_12874);
nor U16170 (N_16170,N_14439,N_13482);
and U16171 (N_16171,N_12894,N_14305);
or U16172 (N_16172,N_14004,N_14188);
nor U16173 (N_16173,N_14151,N_14470);
and U16174 (N_16174,N_13694,N_13910);
or U16175 (N_16175,N_15216,N_14970);
or U16176 (N_16176,N_15398,N_14238);
and U16177 (N_16177,N_15129,N_15338);
nand U16178 (N_16178,N_13239,N_15509);
nand U16179 (N_16179,N_12562,N_13907);
or U16180 (N_16180,N_14007,N_14859);
nand U16181 (N_16181,N_14515,N_15056);
or U16182 (N_16182,N_15049,N_14746);
nor U16183 (N_16183,N_14115,N_13797);
nand U16184 (N_16184,N_14544,N_14617);
nand U16185 (N_16185,N_13463,N_15496);
and U16186 (N_16186,N_15602,N_13233);
nand U16187 (N_16187,N_14018,N_15092);
and U16188 (N_16188,N_15454,N_14033);
nor U16189 (N_16189,N_14370,N_13371);
or U16190 (N_16190,N_14047,N_12508);
and U16191 (N_16191,N_12529,N_12983);
nor U16192 (N_16192,N_15114,N_14797);
xor U16193 (N_16193,N_13949,N_14608);
or U16194 (N_16194,N_12853,N_14998);
nand U16195 (N_16195,N_14524,N_12865);
nand U16196 (N_16196,N_13041,N_14700);
or U16197 (N_16197,N_14710,N_13117);
nor U16198 (N_16198,N_12556,N_13660);
xnor U16199 (N_16199,N_15149,N_12797);
nand U16200 (N_16200,N_15193,N_12852);
and U16201 (N_16201,N_14528,N_13383);
nand U16202 (N_16202,N_13710,N_14114);
xnor U16203 (N_16203,N_12594,N_15589);
nor U16204 (N_16204,N_14579,N_12872);
and U16205 (N_16205,N_15341,N_13481);
and U16206 (N_16206,N_14818,N_14164);
nand U16207 (N_16207,N_15008,N_13670);
or U16208 (N_16208,N_13774,N_15023);
nor U16209 (N_16209,N_12702,N_15450);
nor U16210 (N_16210,N_13175,N_14861);
xnor U16211 (N_16211,N_13538,N_13847);
nand U16212 (N_16212,N_13010,N_15253);
or U16213 (N_16213,N_14947,N_14810);
nand U16214 (N_16214,N_14995,N_14093);
and U16215 (N_16215,N_14269,N_12930);
xnor U16216 (N_16216,N_14184,N_13913);
or U16217 (N_16217,N_14474,N_15118);
nand U16218 (N_16218,N_12799,N_15592);
and U16219 (N_16219,N_13860,N_14463);
nor U16220 (N_16220,N_14446,N_12708);
or U16221 (N_16221,N_13124,N_12908);
and U16222 (N_16222,N_13519,N_13112);
nand U16223 (N_16223,N_13106,N_13533);
and U16224 (N_16224,N_13788,N_12697);
or U16225 (N_16225,N_14643,N_14504);
nand U16226 (N_16226,N_14847,N_13599);
and U16227 (N_16227,N_15458,N_14589);
and U16228 (N_16228,N_15479,N_12964);
nor U16229 (N_16229,N_14270,N_14112);
nand U16230 (N_16230,N_13057,N_14261);
or U16231 (N_16231,N_15354,N_15085);
or U16232 (N_16232,N_15012,N_12665);
nor U16233 (N_16233,N_13403,N_13238);
or U16234 (N_16234,N_14051,N_14105);
and U16235 (N_16235,N_13315,N_12846);
xnor U16236 (N_16236,N_13327,N_13369);
nor U16237 (N_16237,N_14872,N_13586);
nand U16238 (N_16238,N_14139,N_15553);
nor U16239 (N_16239,N_14420,N_13114);
or U16240 (N_16240,N_13176,N_14907);
xor U16241 (N_16241,N_15210,N_15073);
or U16242 (N_16242,N_14168,N_15158);
or U16243 (N_16243,N_12763,N_12539);
nor U16244 (N_16244,N_14659,N_12592);
or U16245 (N_16245,N_14374,N_15273);
nor U16246 (N_16246,N_14989,N_13212);
nor U16247 (N_16247,N_13595,N_13072);
and U16248 (N_16248,N_14077,N_15598);
nand U16249 (N_16249,N_15044,N_14837);
nand U16250 (N_16250,N_12611,N_13340);
or U16251 (N_16251,N_13757,N_14424);
nand U16252 (N_16252,N_12955,N_15084);
nor U16253 (N_16253,N_12670,N_14704);
or U16254 (N_16254,N_15542,N_14204);
nor U16255 (N_16255,N_14646,N_13701);
or U16256 (N_16256,N_13039,N_13532);
nand U16257 (N_16257,N_15165,N_14431);
nand U16258 (N_16258,N_14118,N_15347);
nor U16259 (N_16259,N_13952,N_12795);
nor U16260 (N_16260,N_13572,N_12997);
and U16261 (N_16261,N_12552,N_13895);
nand U16262 (N_16262,N_15578,N_14278);
nor U16263 (N_16263,N_13066,N_14864);
and U16264 (N_16264,N_13859,N_14031);
xnor U16265 (N_16265,N_13646,N_14120);
nand U16266 (N_16266,N_13294,N_14615);
and U16267 (N_16267,N_13814,N_14226);
and U16268 (N_16268,N_13338,N_12716);
and U16269 (N_16269,N_13121,N_14412);
nand U16270 (N_16270,N_14199,N_13093);
nand U16271 (N_16271,N_13926,N_13166);
nand U16272 (N_16272,N_13347,N_14751);
or U16273 (N_16273,N_14377,N_14692);
xor U16274 (N_16274,N_14612,N_13139);
nand U16275 (N_16275,N_13460,N_13920);
nand U16276 (N_16276,N_12730,N_12579);
nand U16277 (N_16277,N_12849,N_15405);
or U16278 (N_16278,N_14965,N_13971);
and U16279 (N_16279,N_12884,N_15335);
nor U16280 (N_16280,N_12710,N_14558);
xnor U16281 (N_16281,N_13407,N_13923);
nand U16282 (N_16282,N_13591,N_14940);
or U16283 (N_16283,N_14614,N_13515);
or U16284 (N_16284,N_14673,N_13394);
and U16285 (N_16285,N_15040,N_15332);
nor U16286 (N_16286,N_12871,N_15400);
or U16287 (N_16287,N_13069,N_12571);
nand U16288 (N_16288,N_14403,N_15532);
nor U16289 (N_16289,N_14909,N_14848);
or U16290 (N_16290,N_12589,N_14250);
or U16291 (N_16291,N_14013,N_14724);
and U16292 (N_16292,N_15544,N_14791);
or U16293 (N_16293,N_14992,N_13654);
nand U16294 (N_16294,N_14803,N_15611);
nor U16295 (N_16295,N_13034,N_14828);
or U16296 (N_16296,N_14944,N_13087);
nand U16297 (N_16297,N_14237,N_14669);
or U16298 (N_16298,N_13320,N_14912);
nand U16299 (N_16299,N_14331,N_13632);
nand U16300 (N_16300,N_15397,N_13436);
or U16301 (N_16301,N_14533,N_15340);
and U16302 (N_16302,N_12564,N_13995);
and U16303 (N_16303,N_12891,N_14244);
xor U16304 (N_16304,N_12848,N_13398);
nor U16305 (N_16305,N_14293,N_13486);
xnor U16306 (N_16306,N_12671,N_14393);
xor U16307 (N_16307,N_13553,N_12680);
nand U16308 (N_16308,N_14119,N_13764);
nand U16309 (N_16309,N_15325,N_14545);
nor U16310 (N_16310,N_14502,N_15264);
nand U16311 (N_16311,N_12990,N_12960);
nand U16312 (N_16312,N_12921,N_13943);
nor U16313 (N_16313,N_15021,N_14819);
nor U16314 (N_16314,N_14324,N_13254);
nor U16315 (N_16315,N_13291,N_12633);
xnor U16316 (N_16316,N_14672,N_12793);
nand U16317 (N_16317,N_15095,N_15342);
or U16318 (N_16318,N_15540,N_13630);
xnor U16319 (N_16319,N_13274,N_13356);
xnor U16320 (N_16320,N_13290,N_15473);
and U16321 (N_16321,N_14258,N_15278);
or U16322 (N_16322,N_13620,N_13567);
or U16323 (N_16323,N_14071,N_15211);
xnor U16324 (N_16324,N_13781,N_14379);
nand U16325 (N_16325,N_13387,N_14855);
nand U16326 (N_16326,N_13840,N_13331);
and U16327 (N_16327,N_12619,N_15063);
nand U16328 (N_16328,N_14813,N_12927);
nand U16329 (N_16329,N_12943,N_12623);
nor U16330 (N_16330,N_15006,N_13473);
nor U16331 (N_16331,N_13099,N_12574);
nor U16332 (N_16332,N_13026,N_13541);
nor U16333 (N_16333,N_13303,N_13969);
nand U16334 (N_16334,N_13419,N_15484);
nor U16335 (N_16335,N_13768,N_13776);
or U16336 (N_16336,N_12689,N_12957);
nor U16337 (N_16337,N_12531,N_12909);
xor U16338 (N_16338,N_13193,N_13987);
nor U16339 (N_16339,N_14320,N_15477);
and U16340 (N_16340,N_12557,N_14187);
or U16341 (N_16341,N_14517,N_13794);
nand U16342 (N_16342,N_14606,N_15029);
nand U16343 (N_16343,N_15052,N_14520);
nor U16344 (N_16344,N_15603,N_12549);
nor U16345 (N_16345,N_14304,N_14801);
or U16346 (N_16346,N_13187,N_12857);
xor U16347 (N_16347,N_13934,N_14240);
nand U16348 (N_16348,N_12553,N_12996);
and U16349 (N_16349,N_12754,N_13230);
and U16350 (N_16350,N_13672,N_13267);
nand U16351 (N_16351,N_13311,N_14571);
and U16352 (N_16352,N_15161,N_13636);
or U16353 (N_16353,N_13872,N_12842);
nor U16354 (N_16354,N_14744,N_15418);
xor U16355 (N_16355,N_15137,N_12511);
and U16356 (N_16356,N_14337,N_14937);
nor U16357 (N_16357,N_12841,N_14676);
or U16358 (N_16358,N_15572,N_13716);
or U16359 (N_16359,N_13161,N_13470);
or U16360 (N_16360,N_14343,N_15048);
or U16361 (N_16361,N_15311,N_14779);
or U16362 (N_16362,N_14197,N_13594);
or U16363 (N_16363,N_13639,N_14074);
nand U16364 (N_16364,N_13706,N_13959);
nor U16365 (N_16365,N_13766,N_13765);
and U16366 (N_16366,N_14531,N_13115);
xnor U16367 (N_16367,N_13092,N_15385);
nor U16368 (N_16368,N_14567,N_14124);
or U16369 (N_16369,N_12679,N_14088);
or U16370 (N_16370,N_14208,N_13603);
nand U16371 (N_16371,N_12648,N_15107);
nand U16372 (N_16372,N_13333,N_12542);
or U16373 (N_16373,N_13374,N_12862);
or U16374 (N_16374,N_14627,N_13634);
or U16375 (N_16375,N_15015,N_15480);
or U16376 (N_16376,N_13448,N_13597);
or U16377 (N_16377,N_14300,N_14090);
and U16378 (N_16378,N_14776,N_14479);
nand U16379 (N_16379,N_13264,N_13351);
nand U16380 (N_16380,N_14375,N_15444);
nand U16381 (N_16381,N_15213,N_14537);
and U16382 (N_16382,N_12602,N_14407);
nor U16383 (N_16383,N_13189,N_14894);
nand U16384 (N_16384,N_14967,N_15409);
nand U16385 (N_16385,N_14929,N_14425);
nor U16386 (N_16386,N_13104,N_14406);
and U16387 (N_16387,N_14128,N_13686);
nor U16388 (N_16388,N_15534,N_13471);
nand U16389 (N_16389,N_13206,N_14445);
or U16390 (N_16390,N_13536,N_15277);
nor U16391 (N_16391,N_13740,N_12500);
or U16392 (N_16392,N_15348,N_14667);
nand U16393 (N_16393,N_13752,N_12513);
xor U16394 (N_16394,N_14351,N_13666);
nand U16395 (N_16395,N_15220,N_14295);
or U16396 (N_16396,N_13593,N_14682);
nor U16397 (N_16397,N_13962,N_14137);
and U16398 (N_16398,N_15545,N_14193);
and U16399 (N_16399,N_13941,N_13520);
xnor U16400 (N_16400,N_12525,N_12826);
or U16401 (N_16401,N_15233,N_13202);
and U16402 (N_16402,N_15492,N_12967);
and U16403 (N_16403,N_15299,N_14605);
nor U16404 (N_16404,N_12827,N_14535);
nand U16405 (N_16405,N_14255,N_13601);
nand U16406 (N_16406,N_14411,N_13736);
nor U16407 (N_16407,N_13658,N_13368);
nor U16408 (N_16408,N_14296,N_14685);
and U16409 (N_16409,N_15139,N_14239);
and U16410 (N_16410,N_13359,N_14789);
nor U16411 (N_16411,N_13641,N_14728);
nor U16412 (N_16412,N_15419,N_15055);
or U16413 (N_16413,N_14591,N_15356);
and U16414 (N_16414,N_14619,N_13009);
nand U16415 (N_16415,N_13855,N_14851);
nor U16416 (N_16416,N_13546,N_13416);
and U16417 (N_16417,N_13589,N_14469);
and U16418 (N_16418,N_12578,N_13626);
and U16419 (N_16419,N_13763,N_15498);
and U16420 (N_16420,N_12916,N_15586);
nor U16421 (N_16421,N_12728,N_12970);
and U16422 (N_16422,N_13137,N_15547);
xnor U16423 (N_16423,N_14082,N_13842);
nand U16424 (N_16424,N_13016,N_13937);
and U16425 (N_16425,N_14323,N_14030);
nor U16426 (N_16426,N_13975,N_13877);
nor U16427 (N_16427,N_14131,N_13283);
or U16428 (N_16428,N_15616,N_13035);
nor U16429 (N_16429,N_12707,N_15187);
or U16430 (N_16430,N_15305,N_14058);
nand U16431 (N_16431,N_13305,N_13197);
nand U16432 (N_16432,N_12768,N_13582);
nand U16433 (N_16433,N_12575,N_14182);
or U16434 (N_16434,N_12870,N_15414);
or U16435 (N_16435,N_12757,N_15083);
nand U16436 (N_16436,N_15393,N_14860);
and U16437 (N_16437,N_15285,N_13635);
and U16438 (N_16438,N_15403,N_12774);
nand U16439 (N_16439,N_15276,N_15359);
or U16440 (N_16440,N_14213,N_12569);
or U16441 (N_16441,N_12959,N_14466);
xor U16442 (N_16442,N_13856,N_14454);
xnor U16443 (N_16443,N_14823,N_13213);
nor U16444 (N_16444,N_13076,N_13349);
nor U16445 (N_16445,N_13082,N_12715);
nand U16446 (N_16446,N_14895,N_12899);
and U16447 (N_16447,N_14858,N_13733);
and U16448 (N_16448,N_15075,N_14957);
xnor U16449 (N_16449,N_13742,N_14629);
or U16450 (N_16450,N_14363,N_14613);
xor U16451 (N_16451,N_13832,N_14898);
or U16452 (N_16452,N_14347,N_13384);
or U16453 (N_16453,N_12926,N_14275);
or U16454 (N_16454,N_13078,N_14690);
nor U16455 (N_16455,N_12643,N_14587);
and U16456 (N_16456,N_15513,N_13222);
and U16457 (N_16457,N_15067,N_13881);
xnor U16458 (N_16458,N_14478,N_14053);
nor U16459 (N_16459,N_14927,N_13422);
and U16460 (N_16460,N_13659,N_13598);
and U16461 (N_16461,N_12590,N_13816);
nor U16462 (N_16462,N_14341,N_14829);
or U16463 (N_16463,N_14285,N_14757);
nor U16464 (N_16464,N_14212,N_15160);
xnor U16465 (N_16465,N_12893,N_13152);
nor U16466 (N_16466,N_14671,N_13060);
and U16467 (N_16467,N_12946,N_15086);
and U16468 (N_16468,N_14310,N_14271);
or U16469 (N_16469,N_13130,N_13441);
or U16470 (N_16470,N_13649,N_13769);
nand U16471 (N_16471,N_14382,N_13908);
or U16472 (N_16472,N_12823,N_14736);
nand U16473 (N_16473,N_14345,N_15108);
nor U16474 (N_16474,N_14557,N_14028);
nor U16475 (N_16475,N_13986,N_14230);
nor U16476 (N_16476,N_14101,N_12540);
or U16477 (N_16477,N_12598,N_14979);
or U16478 (N_16478,N_14288,N_13675);
and U16479 (N_16479,N_13086,N_12784);
and U16480 (N_16480,N_15554,N_13123);
or U16481 (N_16481,N_13751,N_15263);
nand U16482 (N_16482,N_12610,N_14434);
nor U16483 (N_16483,N_14993,N_13209);
xnor U16484 (N_16484,N_14353,N_13867);
nand U16485 (N_16485,N_14348,N_13885);
or U16486 (N_16486,N_14234,N_13990);
nand U16487 (N_16487,N_12544,N_14036);
xor U16488 (N_16488,N_14693,N_14764);
xor U16489 (N_16489,N_14014,N_13918);
nand U16490 (N_16490,N_14769,N_14892);
nor U16491 (N_16491,N_13663,N_12503);
nor U16492 (N_16492,N_12951,N_14951);
and U16493 (N_16493,N_14678,N_15529);
nor U16494 (N_16494,N_15504,N_14832);
or U16495 (N_16495,N_14889,N_13824);
nand U16496 (N_16496,N_13753,N_14748);
nand U16497 (N_16497,N_14279,N_14702);
nor U16498 (N_16498,N_12573,N_15487);
nor U16499 (N_16499,N_12777,N_14580);
nor U16500 (N_16500,N_12829,N_15170);
or U16501 (N_16501,N_14792,N_15011);
xnor U16502 (N_16502,N_13004,N_14459);
nor U16503 (N_16503,N_14657,N_15407);
nor U16504 (N_16504,N_14988,N_14448);
or U16505 (N_16505,N_15563,N_14228);
nand U16506 (N_16506,N_14085,N_12995);
nor U16507 (N_16507,N_15422,N_12845);
and U16508 (N_16508,N_12868,N_14816);
and U16509 (N_16509,N_15460,N_15371);
and U16510 (N_16510,N_12652,N_12789);
nand U16511 (N_16511,N_13665,N_12912);
or U16512 (N_16512,N_13713,N_14103);
xor U16513 (N_16513,N_15261,N_14963);
nand U16514 (N_16514,N_14476,N_15249);
nor U16515 (N_16515,N_14560,N_14329);
xnor U16516 (N_16516,N_12764,N_15106);
nand U16517 (N_16517,N_14260,N_15438);
and U16518 (N_16518,N_14035,N_13790);
and U16519 (N_16519,N_14584,N_14070);
nand U16520 (N_16520,N_13052,N_12742);
nor U16521 (N_16521,N_13440,N_14824);
nand U16522 (N_16522,N_12879,N_15511);
or U16523 (N_16523,N_14875,N_13450);
nand U16524 (N_16524,N_15198,N_13231);
xnor U16525 (N_16525,N_15614,N_14796);
nand U16526 (N_16526,N_15580,N_15201);
or U16527 (N_16527,N_14625,N_15384);
nor U16528 (N_16528,N_12779,N_14867);
nor U16529 (N_16529,N_14104,N_15109);
or U16530 (N_16530,N_13207,N_13936);
or U16531 (N_16531,N_13205,N_14986);
or U16532 (N_16532,N_14003,N_13432);
nand U16533 (N_16533,N_13671,N_15200);
xnor U16534 (N_16534,N_13869,N_15176);
or U16535 (N_16535,N_14473,N_14689);
xor U16536 (N_16536,N_13487,N_14149);
or U16537 (N_16537,N_14686,N_13263);
nand U16538 (N_16538,N_14699,N_15244);
nor U16539 (N_16539,N_14883,N_14266);
xor U16540 (N_16540,N_14541,N_12954);
xnor U16541 (N_16541,N_13834,N_14656);
nor U16542 (N_16542,N_14461,N_12998);
or U16543 (N_16543,N_13269,N_14592);
nand U16544 (N_16544,N_13411,N_13530);
and U16545 (N_16545,N_15076,N_13317);
nand U16546 (N_16546,N_14494,N_14507);
xor U16547 (N_16547,N_14259,N_14358);
xnor U16548 (N_16548,N_13803,N_13296);
nand U16549 (N_16549,N_14481,N_12737);
nor U16550 (N_16550,N_13980,N_14694);
and U16551 (N_16551,N_13038,N_14721);
nor U16552 (N_16552,N_13414,N_14928);
nor U16553 (N_16553,N_12530,N_14555);
and U16554 (N_16554,N_13443,N_13287);
and U16555 (N_16555,N_12886,N_12949);
or U16556 (N_16556,N_15321,N_15260);
or U16557 (N_16557,N_14221,N_13466);
nor U16558 (N_16558,N_13644,N_14022);
and U16559 (N_16559,N_13134,N_15459);
nand U16560 (N_16560,N_13226,N_12521);
or U16561 (N_16561,N_13314,N_15240);
and U16562 (N_16562,N_12658,N_13122);
or U16563 (N_16563,N_14073,N_13428);
xnor U16564 (N_16564,N_13214,N_13046);
or U16565 (N_16565,N_14595,N_15266);
nand U16566 (N_16566,N_12748,N_12813);
nor U16567 (N_16567,N_13476,N_14747);
nor U16568 (N_16568,N_13048,N_12629);
or U16569 (N_16569,N_13318,N_14102);
or U16570 (N_16570,N_12735,N_12843);
xnor U16571 (N_16571,N_15074,N_14456);
xnor U16572 (N_16572,N_15593,N_13126);
xnor U16573 (N_16573,N_13221,N_13664);
nand U16574 (N_16574,N_15417,N_13380);
and U16575 (N_16575,N_13184,N_13873);
and U16576 (N_16576,N_13807,N_14674);
nand U16577 (N_16577,N_12734,N_13610);
and U16578 (N_16578,N_15436,N_13993);
and U16579 (N_16579,N_15078,N_13939);
nand U16580 (N_16580,N_13050,N_15364);
nor U16581 (N_16581,N_15485,N_15231);
nor U16582 (N_16582,N_15313,N_13032);
nor U16583 (N_16583,N_13628,N_13091);
nand U16584 (N_16584,N_14141,N_14878);
nand U16585 (N_16585,N_14910,N_14596);
xnor U16586 (N_16586,N_15427,N_12855);
nor U16587 (N_16587,N_13240,N_13118);
and U16588 (N_16588,N_13278,N_14336);
nand U16589 (N_16589,N_15588,N_15467);
nor U16590 (N_16590,N_12699,N_14508);
or U16591 (N_16591,N_12690,N_14542);
and U16592 (N_16592,N_12696,N_14961);
xor U16593 (N_16593,N_13958,N_14522);
nor U16594 (N_16594,N_12950,N_14802);
nand U16595 (N_16595,N_14688,N_13822);
nand U16596 (N_16596,N_12627,N_15138);
or U16597 (N_16597,N_13754,N_14462);
and U16598 (N_16598,N_13024,N_15169);
or U16599 (N_16599,N_15298,N_14144);
and U16600 (N_16600,N_14598,N_12563);
or U16601 (N_16601,N_14021,N_13298);
or U16602 (N_16602,N_14712,N_14108);
nor U16603 (N_16603,N_14708,N_14814);
xor U16604 (N_16604,N_12866,N_14489);
xnor U16605 (N_16605,N_12663,N_13090);
and U16606 (N_16606,N_14126,N_12593);
xnor U16607 (N_16607,N_13051,N_13245);
xnor U16608 (N_16608,N_14214,N_14195);
and U16609 (N_16609,N_14793,N_15521);
or U16610 (N_16610,N_13173,N_14299);
and U16611 (N_16611,N_12576,N_15432);
nand U16612 (N_16612,N_13149,N_14890);
or U16613 (N_16613,N_13154,N_14339);
nand U16614 (N_16614,N_13685,N_15206);
and U16615 (N_16615,N_13722,N_15383);
nor U16616 (N_16616,N_13188,N_14561);
or U16617 (N_16617,N_12804,N_14854);
nor U16618 (N_16618,N_12543,N_15362);
nand U16619 (N_16619,N_13571,N_15337);
nor U16620 (N_16620,N_15079,N_14661);
nor U16621 (N_16621,N_13417,N_14065);
and U16622 (N_16622,N_12773,N_14158);
and U16623 (N_16623,N_13055,N_14549);
or U16624 (N_16624,N_12681,N_15032);
nor U16625 (N_16625,N_14684,N_13171);
and U16626 (N_16626,N_14611,N_14675);
nand U16627 (N_16627,N_14799,N_13798);
or U16628 (N_16628,N_13194,N_12800);
xnor U16629 (N_16629,N_14984,N_15288);
nor U16630 (N_16630,N_12565,N_12963);
or U16631 (N_16631,N_13772,N_14774);
or U16632 (N_16632,N_14443,N_12527);
and U16633 (N_16633,N_14423,N_13728);
nand U16634 (N_16634,N_13012,N_14575);
nor U16635 (N_16635,N_14009,N_15164);
nand U16636 (N_16636,N_12673,N_15381);
nor U16637 (N_16637,N_12588,N_13297);
nand U16638 (N_16638,N_14836,N_13783);
nor U16639 (N_16639,N_12537,N_13721);
nand U16640 (N_16640,N_14636,N_13848);
nor U16641 (N_16641,N_13735,N_14565);
nand U16642 (N_16642,N_15431,N_14066);
nor U16643 (N_16643,N_14396,N_13464);
nand U16644 (N_16644,N_15518,N_14175);
or U16645 (N_16645,N_13514,N_13953);
nand U16646 (N_16646,N_14620,N_13653);
nor U16647 (N_16647,N_15556,N_14191);
nor U16648 (N_16648,N_12790,N_14857);
nand U16649 (N_16649,N_13580,N_14019);
xor U16650 (N_16650,N_15159,N_13215);
nand U16651 (N_16651,N_12796,N_12888);
nand U16652 (N_16652,N_14089,N_14216);
nor U16653 (N_16653,N_14547,N_14978);
or U16654 (N_16654,N_13113,N_12559);
nand U16655 (N_16655,N_14717,N_15566);
or U16656 (N_16656,N_14972,N_13652);
and U16657 (N_16657,N_14256,N_14755);
nand U16658 (N_16658,N_12587,N_13306);
nand U16659 (N_16659,N_12585,N_14294);
nand U16660 (N_16660,N_14016,N_12778);
or U16661 (N_16661,N_13810,N_13456);
and U16662 (N_16662,N_12873,N_14383);
nor U16663 (N_16663,N_14475,N_15156);
nand U16664 (N_16664,N_13645,N_14037);
nand U16665 (N_16665,N_13405,N_14328);
nand U16666 (N_16666,N_15512,N_14060);
or U16667 (N_16667,N_15155,N_14264);
or U16668 (N_16668,N_13951,N_14447);
nand U16669 (N_16669,N_13021,N_12674);
nand U16670 (N_16670,N_15425,N_12877);
nand U16671 (N_16671,N_14486,N_13402);
and U16672 (N_16672,N_13119,N_14856);
nor U16673 (N_16673,N_13796,N_14881);
nor U16674 (N_16674,N_14644,N_14725);
nand U16675 (N_16675,N_15162,N_12816);
or U16676 (N_16676,N_12962,N_14903);
or U16677 (N_16677,N_13966,N_14999);
or U16678 (N_16678,N_12787,N_13498);
and U16679 (N_16679,N_13148,N_13047);
and U16680 (N_16680,N_13726,N_13638);
and U16681 (N_16681,N_13342,N_13462);
nand U16682 (N_16682,N_13531,N_14173);
or U16683 (N_16683,N_13475,N_12875);
nand U16684 (N_16684,N_12607,N_13629);
and U16685 (N_16685,N_13785,N_12669);
nor U16686 (N_16686,N_14032,N_14785);
nor U16687 (N_16687,N_14268,N_15502);
xnor U16688 (N_16688,N_12838,N_12535);
nor U16689 (N_16689,N_12672,N_13809);
or U16690 (N_16690,N_15223,N_14344);
or U16691 (N_16691,N_13065,N_13495);
and U16692 (N_16692,N_12977,N_13607);
or U16693 (N_16693,N_13312,N_14482);
and U16694 (N_16694,N_13617,N_14313);
or U16695 (N_16695,N_13865,N_13467);
or U16696 (N_16696,N_14647,N_15252);
xnor U16697 (N_16697,N_15143,N_13508);
or U16698 (N_16698,N_15345,N_15010);
and U16699 (N_16699,N_15147,N_15623);
or U16700 (N_16700,N_15617,N_13818);
xnor U16701 (N_16701,N_14687,N_14194);
or U16702 (N_16702,N_14130,N_13262);
and U16703 (N_16703,N_15478,N_13285);
or U16704 (N_16704,N_12818,N_14782);
nor U16705 (N_16705,N_12887,N_14061);
and U16706 (N_16706,N_13775,N_14919);
nor U16707 (N_16707,N_12591,N_13003);
nand U16708 (N_16708,N_13558,N_15124);
xor U16709 (N_16709,N_15128,N_13488);
nor U16710 (N_16710,N_15047,N_13053);
nor U16711 (N_16711,N_14781,N_13346);
nand U16712 (N_16712,N_13612,N_13619);
nand U16713 (N_16713,N_14510,N_13727);
nor U16714 (N_16714,N_14604,N_14525);
or U16715 (N_16715,N_13989,N_14714);
nor U16716 (N_16716,N_14863,N_14113);
or U16717 (N_16717,N_14526,N_14835);
nand U16718 (N_16718,N_15433,N_14000);
or U16719 (N_16719,N_14005,N_13150);
and U16720 (N_16720,N_13616,N_15284);
and U16721 (N_16721,N_14918,N_14934);
or U16722 (N_16722,N_13459,N_12854);
and U16723 (N_16723,N_14063,N_14095);
or U16724 (N_16724,N_13494,N_14409);
or U16725 (N_16725,N_14179,N_13309);
nor U16726 (N_16726,N_12746,N_13900);
xnor U16727 (N_16727,N_13330,N_14610);
nand U16728 (N_16728,N_14885,N_14564);
nand U16729 (N_16729,N_13381,N_13703);
and U16730 (N_16730,N_13431,N_14338);
or U16731 (N_16731,N_14497,N_14870);
and U16732 (N_16732,N_12567,N_12890);
nor U16733 (N_16733,N_13795,N_12545);
or U16734 (N_16734,N_13177,N_13404);
or U16735 (N_16735,N_12582,N_13828);
nand U16736 (N_16736,N_13484,N_14150);
and U16737 (N_16737,N_12807,N_14287);
nor U16738 (N_16738,N_14138,N_13760);
or U16739 (N_16739,N_12762,N_14442);
nor U16740 (N_16740,N_13624,N_15133);
and U16741 (N_16741,N_13647,N_13295);
nor U16742 (N_16742,N_12719,N_13677);
xnor U16743 (N_16743,N_14534,N_14001);
nand U16744 (N_16744,N_12928,N_14559);
nor U16745 (N_16745,N_15601,N_14391);
nand U16746 (N_16746,N_14265,N_14697);
and U16747 (N_16747,N_13491,N_12867);
and U16748 (N_16748,N_13919,N_14452);
nor U16749 (N_16749,N_14653,N_13564);
nand U16750 (N_16750,N_15248,N_14222);
or U16751 (N_16751,N_14743,N_13559);
or U16752 (N_16752,N_14290,N_14680);
nor U16753 (N_16753,N_15351,N_15620);
nand U16754 (N_16754,N_13812,N_14034);
nor U16755 (N_16755,N_13192,N_15568);
nand U16756 (N_16756,N_13909,N_13135);
nor U16757 (N_16757,N_15561,N_13778);
or U16758 (N_16758,N_14389,N_13461);
and U16759 (N_16759,N_13912,N_15318);
or U16760 (N_16760,N_15320,N_14360);
or U16761 (N_16761,N_12505,N_13717);
and U16762 (N_16762,N_15331,N_15528);
and U16763 (N_16763,N_13435,N_15111);
nor U16764 (N_16764,N_14386,N_12992);
and U16765 (N_16765,N_15082,N_14901);
nand U16766 (N_16766,N_13447,N_14198);
or U16767 (N_16767,N_14390,N_15127);
or U16768 (N_16768,N_14572,N_13158);
nor U16769 (N_16769,N_15390,N_15510);
xor U16770 (N_16770,N_13138,N_15297);
nor U16771 (N_16771,N_14536,N_15141);
and U16772 (N_16772,N_13286,N_14055);
and U16773 (N_16773,N_13650,N_14455);
xor U16774 (N_16774,N_12608,N_12808);
nor U16775 (N_16775,N_12727,N_15508);
and U16776 (N_16776,N_13500,N_12817);
or U16777 (N_16777,N_13537,N_14326);
nor U16778 (N_16778,N_14853,N_13243);
and U16779 (N_16779,N_13802,N_13576);
xor U16780 (N_16780,N_15440,N_15039);
nor U16781 (N_16781,N_13906,N_13275);
and U16782 (N_16782,N_14518,N_12942);
and U16783 (N_16783,N_15121,N_15585);
xor U16784 (N_16784,N_13932,N_14444);
or U16785 (N_16785,N_12892,N_14954);
nor U16786 (N_16786,N_13446,N_13651);
nand U16787 (N_16787,N_12814,N_15452);
nand U16788 (N_16788,N_14281,N_13887);
nor U16789 (N_16789,N_15442,N_14437);
or U16790 (N_16790,N_15185,N_13427);
or U16791 (N_16791,N_15069,N_13507);
xor U16792 (N_16792,N_13745,N_12536);
and U16793 (N_16793,N_12920,N_15157);
and U16794 (N_16794,N_13534,N_14696);
and U16795 (N_16795,N_14849,N_13876);
and U16796 (N_16796,N_13049,N_14729);
and U16797 (N_16797,N_15053,N_13396);
nor U16798 (N_16798,N_12646,N_12925);
or U16799 (N_16799,N_15604,N_15218);
or U16800 (N_16800,N_13618,N_14593);
or U16801 (N_16801,N_14758,N_14920);
nor U16802 (N_16802,N_15555,N_13643);
nor U16803 (N_16803,N_14543,N_13974);
nor U16804 (N_16804,N_14841,N_13724);
xnor U16805 (N_16805,N_14079,N_12935);
xor U16806 (N_16806,N_14805,N_15054);
nand U16807 (N_16807,N_13129,N_14274);
or U16808 (N_16808,N_13983,N_14638);
nor U16809 (N_16809,N_14364,N_14372);
or U16810 (N_16810,N_12659,N_12599);
nor U16811 (N_16811,N_12640,N_14923);
nand U16812 (N_16812,N_13509,N_14709);
nor U16813 (N_16813,N_13474,N_13080);
nor U16814 (N_16814,N_14148,N_13901);
and U16815 (N_16815,N_12900,N_13690);
xor U16816 (N_16816,N_13109,N_14730);
xor U16817 (N_16817,N_13493,N_14662);
and U16818 (N_16818,N_12825,N_14201);
nor U16819 (N_16819,N_15423,N_15000);
and U16820 (N_16820,N_13835,N_15429);
nor U16821 (N_16821,N_12805,N_14449);
xor U16822 (N_16822,N_13325,N_14839);
nand U16823 (N_16823,N_12577,N_13748);
or U16824 (N_16824,N_13615,N_15232);
nand U16825 (N_16825,N_15434,N_14745);
nor U16826 (N_16826,N_14143,N_15100);
xnor U16827 (N_16827,N_13850,N_15134);
or U16828 (N_16828,N_13608,N_13268);
xnor U16829 (N_16829,N_14679,N_15236);
or U16830 (N_16830,N_13144,N_15168);
and U16831 (N_16831,N_15061,N_13172);
or U16832 (N_16832,N_14116,N_14262);
nor U16833 (N_16833,N_15404,N_15228);
xor U16834 (N_16834,N_13031,N_14361);
or U16835 (N_16835,N_15527,N_13575);
nand U16836 (N_16836,N_15388,N_15396);
nand U16837 (N_16837,N_13013,N_13273);
and U16838 (N_16838,N_12972,N_13917);
nand U16839 (N_16839,N_12772,N_15464);
nor U16840 (N_16840,N_13715,N_14181);
nor U16841 (N_16841,N_15150,N_14152);
nor U16842 (N_16842,N_13878,N_12758);
and U16843 (N_16843,N_12903,N_13777);
nand U16844 (N_16844,N_13673,N_14602);
and U16845 (N_16845,N_15281,N_13120);
nor U16846 (N_16846,N_12636,N_13705);
nor U16847 (N_16847,N_15142,N_15424);
or U16848 (N_16848,N_15296,N_13883);
or U16849 (N_16849,N_13506,N_14635);
or U16850 (N_16850,N_12863,N_15191);
or U16851 (N_16851,N_14083,N_15182);
nor U16852 (N_16852,N_15557,N_13830);
nor U16853 (N_16853,N_15243,N_13924);
nand U16854 (N_16854,N_12581,N_12736);
and U16855 (N_16855,N_12733,N_13782);
or U16856 (N_16856,N_15267,N_14968);
and U16857 (N_16857,N_15026,N_14902);
or U16858 (N_16858,N_13043,N_13858);
nand U16859 (N_16859,N_12835,N_14546);
and U16860 (N_16860,N_12711,N_13929);
and U16861 (N_16861,N_13518,N_15334);
nor U16862 (N_16862,N_13942,N_14010);
nand U16863 (N_16863,N_13730,N_15550);
nor U16864 (N_16864,N_14825,N_14464);
and U16865 (N_16865,N_15369,N_12938);
nand U16866 (N_16866,N_14297,N_13770);
nand U16867 (N_16867,N_14651,N_12833);
nor U16868 (N_16868,N_13657,N_12776);
nand U16869 (N_16869,N_14215,N_13684);
and U16870 (N_16870,N_14991,N_15315);
nor U16871 (N_16871,N_13568,N_13813);
xnor U16872 (N_16872,N_14852,N_15610);
nand U16873 (N_16873,N_13058,N_15600);
or U16874 (N_16874,N_12994,N_14600);
and U16875 (N_16875,N_14660,N_13037);
xor U16876 (N_16876,N_15339,N_13483);
and U16877 (N_16877,N_13108,N_14716);
nand U16878 (N_16878,N_14458,N_13839);
and U16879 (N_16879,N_15221,N_14663);
nor U16880 (N_16880,N_14509,N_14291);
and U16881 (N_16881,N_15491,N_13833);
xnor U16882 (N_16882,N_15355,N_14373);
nand U16883 (N_16883,N_13972,N_14899);
and U16884 (N_16884,N_13265,N_15549);
xor U16885 (N_16885,N_13820,N_15293);
or U16886 (N_16886,N_14147,N_13750);
or U16887 (N_16887,N_13889,N_15391);
and U16888 (N_16888,N_13401,N_14842);
and U16889 (N_16889,N_15536,N_13054);
and U16890 (N_16890,N_13563,N_13028);
or U16891 (N_16891,N_15030,N_14960);
nand U16892 (N_16892,N_13683,N_15024);
or U16893 (N_16893,N_14209,N_13902);
xnor U16894 (N_16894,N_14136,N_13497);
or U16895 (N_16895,N_13339,N_15481);
or U16896 (N_16896,N_15088,N_15262);
and U16897 (N_16897,N_14026,N_15173);
or U16898 (N_16898,N_14677,N_15122);
or U16899 (N_16899,N_14371,N_14311);
nor U16900 (N_16900,N_13825,N_13183);
nor U16901 (N_16901,N_15590,N_12676);
and U16902 (N_16902,N_13609,N_15562);
or U16903 (N_16903,N_14711,N_12830);
nand U16904 (N_16904,N_13535,N_13180);
and U16905 (N_16905,N_14440,N_15031);
xnor U16906 (N_16906,N_15172,N_14590);
or U16907 (N_16907,N_14931,N_13163);
nor U16908 (N_16908,N_14971,N_14050);
nand U16909 (N_16909,N_14658,N_14263);
or U16910 (N_16910,N_12703,N_13977);
xnor U16911 (N_16911,N_15192,N_15125);
nand U16912 (N_16912,N_13758,N_13182);
or U16913 (N_16913,N_12548,N_12628);
and U16914 (N_16914,N_15020,N_14023);
or U16915 (N_16915,N_13496,N_15245);
nand U16916 (N_16916,N_14639,N_14822);
nor U16917 (N_16917,N_14786,N_13982);
nor U16918 (N_16918,N_13549,N_13903);
nand U16919 (N_16919,N_13237,N_14354);
or U16920 (N_16920,N_12662,N_13370);
and U16921 (N_16921,N_13014,N_14756);
nor U16922 (N_16922,N_12502,N_13792);
or U16923 (N_16923,N_13793,N_14418);
and U16924 (N_16924,N_15560,N_12624);
nor U16925 (N_16925,N_14107,N_14884);
nor U16926 (N_16926,N_14787,N_13242);
and U16927 (N_16927,N_15543,N_15091);
nor U16928 (N_16928,N_14514,N_14527);
nor U16929 (N_16929,N_13479,N_12580);
nand U16930 (N_16930,N_13145,N_13260);
nand U16931 (N_16931,N_14706,N_15538);
nand U16932 (N_16932,N_14356,N_13922);
and U16933 (N_16933,N_14800,N_15301);
nand U16934 (N_16934,N_15009,N_13702);
xor U16935 (N_16935,N_14417,N_13998);
xor U16936 (N_16936,N_15445,N_12691);
nor U16937 (N_16937,N_14308,N_15144);
or U16938 (N_16938,N_15456,N_12945);
or U16939 (N_16939,N_14871,N_12840);
or U16940 (N_16940,N_13746,N_12971);
and U16941 (N_16941,N_13928,N_14521);
nand U16942 (N_16942,N_14734,N_12844);
nor U16943 (N_16943,N_15246,N_14170);
or U16944 (N_16944,N_13836,N_14529);
or U16945 (N_16945,N_13801,N_12677);
nor U16946 (N_16946,N_13389,N_13743);
and U16947 (N_16947,N_14983,N_15428);
xnor U16948 (N_16948,N_15520,N_14133);
or U16949 (N_16949,N_12568,N_13874);
nand U16950 (N_16950,N_14020,N_13492);
or U16951 (N_16951,N_13442,N_15565);
nand U16952 (N_16952,N_12561,N_13723);
nand U16953 (N_16953,N_14498,N_15112);
or U16954 (N_16954,N_13098,N_15197);
and U16955 (N_16955,N_12911,N_14342);
nor U16956 (N_16956,N_15077,N_12683);
nor U16957 (N_16957,N_13552,N_14628);
nand U16958 (N_16958,N_14914,N_12620);
or U16959 (N_16959,N_13732,N_12741);
and U16960 (N_16960,N_13174,N_12788);
nor U16961 (N_16961,N_14492,N_14321);
nor U16962 (N_16962,N_13217,N_14365);
and U16963 (N_16963,N_12600,N_14975);
nand U16964 (N_16964,N_13886,N_13584);
and U16965 (N_16965,N_15503,N_13512);
nand U16966 (N_16966,N_14735,N_12675);
nand U16967 (N_16967,N_12631,N_13927);
and U16968 (N_16968,N_13729,N_12847);
and U16969 (N_16969,N_14097,N_13083);
nand U16970 (N_16970,N_13141,N_14720);
xor U16971 (N_16971,N_13210,N_15476);
nor U16972 (N_16972,N_15070,N_14768);
nand U16973 (N_16973,N_12718,N_13501);
nor U16974 (N_16974,N_13554,N_14811);
nand U16975 (N_16975,N_12729,N_14896);
or U16976 (N_16976,N_14778,N_13453);
nand U16977 (N_16977,N_14042,N_15283);
or U16978 (N_16978,N_14057,N_14621);
and U16979 (N_16979,N_13692,N_13773);
and U16980 (N_16980,N_12792,N_12613);
nor U16981 (N_16981,N_14703,N_13433);
or U16982 (N_16982,N_12856,N_12937);
nor U16983 (N_16983,N_15378,N_15526);
nor U16984 (N_16984,N_15537,N_13925);
nor U16985 (N_16985,N_15286,N_14962);
nand U16986 (N_16986,N_14432,N_15411);
or U16987 (N_16987,N_15310,N_14106);
nand U16988 (N_16988,N_14325,N_13621);
nand U16989 (N_16989,N_13040,N_13761);
nand U16990 (N_16990,N_13988,N_15209);
or U16991 (N_16991,N_13170,N_13490);
or U16992 (N_16992,N_14471,N_14467);
and U16993 (N_16993,N_14913,N_12968);
nand U16994 (N_16994,N_13817,N_13127);
xnor U16995 (N_16995,N_14165,N_12984);
nand U16996 (N_16996,N_13200,N_15466);
nand U16997 (N_16997,N_13799,N_13851);
nor U16998 (N_16998,N_13897,N_13276);
and U16999 (N_16999,N_14932,N_13025);
nor U17000 (N_17000,N_12785,N_12914);
nor U17001 (N_17001,N_14468,N_12637);
or U17002 (N_17002,N_14140,N_13208);
xor U17003 (N_17003,N_15326,N_13800);
and U17004 (N_17004,N_14821,N_14006);
xor U17005 (N_17005,N_13996,N_12656);
nor U17006 (N_17006,N_13623,N_15014);
nor U17007 (N_17007,N_13517,N_14052);
or U17008 (N_17008,N_14183,N_12601);
nand U17009 (N_17009,N_14167,N_14668);
and U17010 (N_17010,N_14936,N_13829);
nor U17011 (N_17011,N_14015,N_14038);
nand U17012 (N_17012,N_12731,N_13204);
or U17013 (N_17013,N_14762,N_13000);
nand U17014 (N_17014,N_13228,N_13679);
xnor U17015 (N_17015,N_14827,N_15045);
nand U17016 (N_17016,N_13424,N_14924);
xor U17017 (N_17017,N_14772,N_15346);
nand U17018 (N_17018,N_14603,N_12738);
or U17019 (N_17019,N_13843,N_13101);
nor U17020 (N_17020,N_13896,N_14830);
nand U17021 (N_17021,N_13196,N_14483);
nand U17022 (N_17022,N_15036,N_14705);
nor U17023 (N_17023,N_13844,N_15102);
xor U17024 (N_17024,N_13976,N_14094);
and U17025 (N_17025,N_13955,N_13418);
nand U17026 (N_17026,N_12504,N_14064);
nand U17027 (N_17027,N_13023,N_14723);
nand U17028 (N_17028,N_14078,N_14551);
nor U17029 (N_17029,N_14384,N_14404);
or U17030 (N_17030,N_12555,N_13771);
nor U17031 (N_17031,N_13469,N_13234);
xnor U17032 (N_17032,N_12756,N_15495);
or U17033 (N_17033,N_12724,N_14623);
nand U17034 (N_17034,N_13406,N_14302);
nor U17035 (N_17035,N_12688,N_14220);
xnor U17036 (N_17036,N_13787,N_14637);
nor U17037 (N_17037,N_13543,N_14665);
nor U17038 (N_17038,N_13186,N_14956);
and U17039 (N_17039,N_12546,N_14162);
or U17040 (N_17040,N_14773,N_14399);
nor U17041 (N_17041,N_14893,N_12694);
nand U17042 (N_17042,N_14129,N_14501);
nand U17043 (N_17043,N_14634,N_13852);
nor U17044 (N_17044,N_13085,N_12923);
nand U17045 (N_17045,N_15437,N_13084);
and U17046 (N_17046,N_13457,N_15581);
and U17047 (N_17047,N_14121,N_14987);
nand U17048 (N_17048,N_12507,N_12625);
and U17049 (N_17049,N_15016,N_12819);
nand U17050 (N_17050,N_14652,N_13911);
and U17051 (N_17051,N_14790,N_12657);
and U17052 (N_17052,N_12953,N_13525);
and U17053 (N_17053,N_14180,N_14516);
and U17054 (N_17054,N_14029,N_13323);
nor U17055 (N_17055,N_13020,N_13185);
and U17056 (N_17056,N_13270,N_15575);
nand U17057 (N_17057,N_15379,N_13914);
nor U17058 (N_17058,N_14145,N_14868);
or U17059 (N_17059,N_14513,N_13472);
xor U17060 (N_17060,N_12766,N_13088);
or U17061 (N_17061,N_15180,N_14253);
or U17062 (N_17062,N_12721,N_13375);
xor U17063 (N_17063,N_13587,N_15034);
and U17064 (N_17064,N_15251,N_13354);
nand U17065 (N_17065,N_14503,N_14416);
nand U17066 (N_17066,N_12919,N_14319);
or U17067 (N_17067,N_14997,N_15146);
nand U17068 (N_17068,N_13410,N_15229);
and U17069 (N_17069,N_13133,N_14235);
and U17070 (N_17070,N_14953,N_14990);
nand U17071 (N_17071,N_14046,N_14938);
nor U17072 (N_17072,N_12821,N_14397);
nand U17073 (N_17073,N_15308,N_13984);
nand U17074 (N_17074,N_14024,N_13915);
nor U17075 (N_17075,N_12913,N_13367);
nor U17076 (N_17076,N_14460,N_12685);
nand U17077 (N_17077,N_12612,N_12661);
and U17078 (N_17078,N_13965,N_13458);
and U17079 (N_17079,N_15376,N_14588);
nand U17080 (N_17080,N_14540,N_12981);
and U17081 (N_17081,N_15489,N_15258);
nand U17082 (N_17082,N_12514,N_14438);
nor U17083 (N_17083,N_14330,N_14298);
nor U17084 (N_17084,N_15322,N_13027);
nand U17085 (N_17085,N_12603,N_13136);
nor U17086 (N_17086,N_13017,N_14582);
nand U17087 (N_17087,N_15399,N_15166);
nor U17088 (N_17088,N_15523,N_13445);
nor U17089 (N_17089,N_14624,N_15570);
and U17090 (N_17090,N_15007,N_15531);
nand U17091 (N_17091,N_14948,N_12765);
and U17092 (N_17092,N_14318,N_15152);
or U17093 (N_17093,N_14246,N_14355);
and U17094 (N_17094,N_12918,N_13337);
or U17095 (N_17095,N_13195,N_14189);
or U17096 (N_17096,N_15135,N_14433);
nor U17097 (N_17097,N_13261,N_14955);
nand U17098 (N_17098,N_13030,N_14943);
nand U17099 (N_17099,N_15003,N_14219);
nor U17100 (N_17100,N_13074,N_12775);
nand U17101 (N_17101,N_13378,N_15382);
or U17102 (N_17102,N_14177,N_12973);
and U17103 (N_17103,N_13526,N_12985);
nand U17104 (N_17104,N_12896,N_13140);
nand U17105 (N_17105,N_14798,N_13905);
and U17106 (N_17106,N_14402,N_13293);
nand U17107 (N_17107,N_13179,N_14068);
nor U17108 (N_17108,N_13700,N_12714);
xor U17109 (N_17109,N_14933,N_13425);
nor U17110 (N_17110,N_12684,N_14741);
and U17111 (N_17111,N_14664,N_12965);
nor U17112 (N_17112,N_13921,N_13390);
nor U17113 (N_17113,N_13588,N_13364);
nand U17114 (N_17114,N_14233,N_14499);
and U17115 (N_17115,N_14251,N_14210);
or U17116 (N_17116,N_12744,N_15104);
nand U17117 (N_17117,N_14457,N_13933);
nor U17118 (N_17118,N_14155,N_13956);
nor U17119 (N_17119,N_14925,N_13838);
and U17120 (N_17120,N_12749,N_14649);
or U17121 (N_17121,N_14218,N_13938);
nor U17122 (N_17122,N_13365,N_15287);
nor U17123 (N_17123,N_13707,N_12523);
or U17124 (N_17124,N_13256,N_14554);
and U17125 (N_17125,N_13827,N_13361);
or U17126 (N_17126,N_13640,N_15329);
and U17127 (N_17127,N_12538,N_15608);
nand U17128 (N_17128,N_12760,N_14922);
or U17129 (N_17129,N_15126,N_13731);
nor U17130 (N_17130,N_13592,N_15167);
xnor U17131 (N_17131,N_15594,N_14622);
nor U17132 (N_17132,N_15269,N_15235);
nand U17133 (N_17133,N_15302,N_14017);
nand U17134 (N_17134,N_15002,N_14357);
and U17135 (N_17135,N_15599,N_14767);
and U17136 (N_17136,N_15465,N_15184);
nand U17137 (N_17137,N_13719,N_15303);
nand U17138 (N_17138,N_14753,N_13875);
nor U17139 (N_17139,N_13871,N_14242);
nand U17140 (N_17140,N_15151,N_14759);
nor U17141 (N_17141,N_13767,N_14267);
or U17142 (N_17142,N_15148,N_14877);
nand U17143 (N_17143,N_15596,N_15214);
xor U17144 (N_17144,N_15099,N_14243);
xnor U17145 (N_17145,N_13409,N_13734);
nor U17146 (N_17146,N_12812,N_15365);
and U17147 (N_17147,N_15415,N_15237);
nor U17148 (N_17148,N_15401,N_12834);
and U17149 (N_17149,N_12851,N_14539);
or U17150 (N_17150,N_12924,N_13094);
nand U17151 (N_17151,N_14573,N_13391);
nor U17152 (N_17152,N_15361,N_15514);
nor U17153 (N_17153,N_15501,N_14833);
or U17154 (N_17154,N_13343,N_14707);
nor U17155 (N_17155,N_13272,N_15247);
and U17156 (N_17156,N_13625,N_12614);
nor U17157 (N_17157,N_12701,N_12940);
or U17158 (N_17158,N_15215,N_15441);
xnor U17159 (N_17159,N_13738,N_13334);
xnor U17160 (N_17160,N_15375,N_15439);
nor U17161 (N_17161,N_13967,N_14876);
nor U17162 (N_17162,N_13452,N_12878);
or U17163 (N_17163,N_15475,N_14039);
nor U17164 (N_17164,N_13288,N_13725);
nor U17165 (N_17165,N_14641,N_12606);
nor U17166 (N_17166,N_14163,N_13605);
xor U17167 (N_17167,N_13744,N_14775);
or U17168 (N_17168,N_13036,N_14349);
nor U17169 (N_17169,N_13841,N_15316);
nor U17170 (N_17170,N_15132,N_13168);
and U17171 (N_17171,N_13412,N_14570);
and U17172 (N_17172,N_13271,N_13600);
or U17173 (N_17173,N_13882,N_14157);
xor U17174 (N_17174,N_13319,N_14980);
nand U17175 (N_17175,N_12709,N_13096);
and U17176 (N_17176,N_12982,N_13581);
and U17177 (N_17177,N_13879,N_14780);
nor U17178 (N_17178,N_15483,N_12720);
nor U17179 (N_17179,N_15255,N_13499);
or U17180 (N_17180,N_12929,N_14075);
xnor U17181 (N_17181,N_14284,N_15430);
nor U17182 (N_17182,N_13248,N_13379);
and U17183 (N_17183,N_13362,N_12713);
or U17184 (N_17184,N_13837,N_14586);
nor U17185 (N_17185,N_13045,N_15353);
or U17186 (N_17186,N_15613,N_14388);
nor U17187 (N_17187,N_14982,N_13927);
nand U17188 (N_17188,N_14114,N_14600);
nand U17189 (N_17189,N_14502,N_13664);
nand U17190 (N_17190,N_15268,N_13896);
or U17191 (N_17191,N_15385,N_14808);
xnor U17192 (N_17192,N_14058,N_15500);
nor U17193 (N_17193,N_13764,N_12902);
or U17194 (N_17194,N_13472,N_13217);
and U17195 (N_17195,N_12663,N_14585);
or U17196 (N_17196,N_12665,N_13352);
and U17197 (N_17197,N_13663,N_13472);
nand U17198 (N_17198,N_14357,N_15426);
xnor U17199 (N_17199,N_13961,N_14788);
xnor U17200 (N_17200,N_15382,N_12718);
or U17201 (N_17201,N_14548,N_14931);
xor U17202 (N_17202,N_12964,N_14887);
and U17203 (N_17203,N_12747,N_14672);
and U17204 (N_17204,N_13417,N_13775);
nor U17205 (N_17205,N_15043,N_12944);
xor U17206 (N_17206,N_14523,N_14424);
xor U17207 (N_17207,N_13568,N_13611);
or U17208 (N_17208,N_13613,N_14561);
or U17209 (N_17209,N_13243,N_14725);
and U17210 (N_17210,N_12809,N_13246);
or U17211 (N_17211,N_14439,N_13890);
xor U17212 (N_17212,N_14543,N_12803);
and U17213 (N_17213,N_12787,N_12861);
or U17214 (N_17214,N_14752,N_13550);
or U17215 (N_17215,N_13164,N_13158);
nand U17216 (N_17216,N_14144,N_13209);
and U17217 (N_17217,N_12719,N_13810);
and U17218 (N_17218,N_13497,N_12878);
nor U17219 (N_17219,N_14600,N_15082);
and U17220 (N_17220,N_13462,N_14390);
and U17221 (N_17221,N_12940,N_12943);
and U17222 (N_17222,N_14763,N_14565);
or U17223 (N_17223,N_12535,N_14778);
xnor U17224 (N_17224,N_13249,N_12645);
nand U17225 (N_17225,N_13847,N_12743);
or U17226 (N_17226,N_12865,N_14369);
nand U17227 (N_17227,N_12882,N_13513);
or U17228 (N_17228,N_12674,N_15403);
nor U17229 (N_17229,N_14451,N_12973);
nand U17230 (N_17230,N_13442,N_14032);
nand U17231 (N_17231,N_15139,N_14862);
and U17232 (N_17232,N_13833,N_13317);
or U17233 (N_17233,N_14538,N_15622);
nand U17234 (N_17234,N_14423,N_15500);
and U17235 (N_17235,N_13766,N_13762);
nand U17236 (N_17236,N_15209,N_15050);
nor U17237 (N_17237,N_14418,N_13900);
xor U17238 (N_17238,N_14458,N_14818);
and U17239 (N_17239,N_12744,N_14425);
or U17240 (N_17240,N_12693,N_14735);
nor U17241 (N_17241,N_13399,N_13128);
nor U17242 (N_17242,N_13309,N_12621);
or U17243 (N_17243,N_12687,N_14175);
xor U17244 (N_17244,N_15559,N_14911);
and U17245 (N_17245,N_14719,N_12684);
nor U17246 (N_17246,N_15112,N_15456);
or U17247 (N_17247,N_15431,N_14087);
or U17248 (N_17248,N_13567,N_12549);
xor U17249 (N_17249,N_15081,N_12901);
or U17250 (N_17250,N_13213,N_13407);
xnor U17251 (N_17251,N_14627,N_13760);
nor U17252 (N_17252,N_13456,N_13080);
nor U17253 (N_17253,N_13664,N_13734);
and U17254 (N_17254,N_15294,N_13312);
nand U17255 (N_17255,N_14360,N_14040);
nand U17256 (N_17256,N_15597,N_14186);
nand U17257 (N_17257,N_12638,N_14397);
nor U17258 (N_17258,N_13495,N_12545);
and U17259 (N_17259,N_13366,N_13828);
xor U17260 (N_17260,N_14989,N_13841);
and U17261 (N_17261,N_14068,N_13074);
nand U17262 (N_17262,N_14273,N_14959);
nor U17263 (N_17263,N_14779,N_13509);
and U17264 (N_17264,N_13112,N_13877);
nor U17265 (N_17265,N_13458,N_14220);
and U17266 (N_17266,N_13063,N_13738);
or U17267 (N_17267,N_14136,N_14651);
xor U17268 (N_17268,N_12956,N_13003);
or U17269 (N_17269,N_15232,N_14851);
nor U17270 (N_17270,N_14376,N_14665);
and U17271 (N_17271,N_13846,N_12639);
or U17272 (N_17272,N_14167,N_12655);
xnor U17273 (N_17273,N_15144,N_14014);
and U17274 (N_17274,N_15618,N_14996);
nor U17275 (N_17275,N_15555,N_14087);
or U17276 (N_17276,N_14772,N_14701);
or U17277 (N_17277,N_14240,N_13951);
nor U17278 (N_17278,N_14428,N_15200);
or U17279 (N_17279,N_13776,N_13291);
or U17280 (N_17280,N_15291,N_15169);
nor U17281 (N_17281,N_13025,N_14881);
xor U17282 (N_17282,N_13629,N_14406);
and U17283 (N_17283,N_14491,N_13913);
nor U17284 (N_17284,N_13363,N_12745);
and U17285 (N_17285,N_14555,N_15325);
and U17286 (N_17286,N_14113,N_13505);
and U17287 (N_17287,N_14188,N_14601);
or U17288 (N_17288,N_13830,N_15025);
and U17289 (N_17289,N_14575,N_14066);
nand U17290 (N_17290,N_13525,N_14167);
xnor U17291 (N_17291,N_14499,N_13336);
nand U17292 (N_17292,N_15053,N_15550);
nor U17293 (N_17293,N_14280,N_12730);
nor U17294 (N_17294,N_13455,N_13069);
nor U17295 (N_17295,N_14200,N_13234);
and U17296 (N_17296,N_13077,N_14770);
and U17297 (N_17297,N_14888,N_13568);
and U17298 (N_17298,N_14833,N_15175);
nand U17299 (N_17299,N_13216,N_15415);
nand U17300 (N_17300,N_14855,N_15181);
nor U17301 (N_17301,N_14976,N_13628);
or U17302 (N_17302,N_14717,N_15047);
nor U17303 (N_17303,N_14571,N_13682);
nor U17304 (N_17304,N_13452,N_12738);
xnor U17305 (N_17305,N_14404,N_14154);
nor U17306 (N_17306,N_13690,N_14087);
nand U17307 (N_17307,N_12518,N_13675);
or U17308 (N_17308,N_12667,N_14219);
or U17309 (N_17309,N_14912,N_13883);
nand U17310 (N_17310,N_13235,N_15471);
nand U17311 (N_17311,N_15203,N_14394);
xor U17312 (N_17312,N_15478,N_14448);
and U17313 (N_17313,N_13460,N_14421);
nand U17314 (N_17314,N_14815,N_12570);
nand U17315 (N_17315,N_12703,N_15337);
nor U17316 (N_17316,N_14952,N_13933);
and U17317 (N_17317,N_14539,N_14142);
nand U17318 (N_17318,N_12526,N_13601);
nand U17319 (N_17319,N_13844,N_15088);
nand U17320 (N_17320,N_13211,N_13484);
or U17321 (N_17321,N_13719,N_12843);
nand U17322 (N_17322,N_12986,N_13085);
nand U17323 (N_17323,N_13631,N_13126);
nor U17324 (N_17324,N_13986,N_13263);
and U17325 (N_17325,N_14819,N_15422);
nor U17326 (N_17326,N_13724,N_13481);
nand U17327 (N_17327,N_14431,N_15264);
nand U17328 (N_17328,N_14210,N_15183);
nor U17329 (N_17329,N_13803,N_14769);
xnor U17330 (N_17330,N_13357,N_13418);
nand U17331 (N_17331,N_13270,N_14571);
nand U17332 (N_17332,N_13468,N_15012);
or U17333 (N_17333,N_13425,N_14557);
and U17334 (N_17334,N_13741,N_15410);
and U17335 (N_17335,N_12904,N_12665);
nand U17336 (N_17336,N_15466,N_14030);
or U17337 (N_17337,N_15126,N_12603);
nand U17338 (N_17338,N_13558,N_14587);
and U17339 (N_17339,N_15094,N_15093);
or U17340 (N_17340,N_13517,N_12833);
nand U17341 (N_17341,N_14997,N_13675);
nor U17342 (N_17342,N_13873,N_13669);
nand U17343 (N_17343,N_12927,N_13546);
or U17344 (N_17344,N_14241,N_13876);
nand U17345 (N_17345,N_12703,N_12916);
nand U17346 (N_17346,N_15464,N_12729);
xor U17347 (N_17347,N_13801,N_13112);
and U17348 (N_17348,N_12957,N_14981);
and U17349 (N_17349,N_13600,N_12917);
or U17350 (N_17350,N_14663,N_13201);
and U17351 (N_17351,N_13666,N_15363);
or U17352 (N_17352,N_13526,N_12711);
xnor U17353 (N_17353,N_14281,N_12764);
and U17354 (N_17354,N_14635,N_12702);
and U17355 (N_17355,N_14620,N_13016);
or U17356 (N_17356,N_13650,N_14411);
nor U17357 (N_17357,N_14379,N_15201);
or U17358 (N_17358,N_14338,N_14911);
nand U17359 (N_17359,N_13298,N_13811);
nand U17360 (N_17360,N_12723,N_14167);
or U17361 (N_17361,N_14104,N_14594);
nor U17362 (N_17362,N_14377,N_15062);
nor U17363 (N_17363,N_13665,N_15065);
or U17364 (N_17364,N_13969,N_13564);
and U17365 (N_17365,N_14645,N_14515);
nor U17366 (N_17366,N_12969,N_14664);
nor U17367 (N_17367,N_13022,N_12642);
nand U17368 (N_17368,N_14939,N_13530);
and U17369 (N_17369,N_15293,N_13422);
nor U17370 (N_17370,N_15545,N_13989);
and U17371 (N_17371,N_15545,N_14127);
nand U17372 (N_17372,N_12842,N_13334);
or U17373 (N_17373,N_13883,N_13518);
or U17374 (N_17374,N_13094,N_13817);
nor U17375 (N_17375,N_14674,N_14340);
nand U17376 (N_17376,N_15376,N_12787);
nor U17377 (N_17377,N_13177,N_12991);
nor U17378 (N_17378,N_15619,N_14315);
and U17379 (N_17379,N_15034,N_12879);
nand U17380 (N_17380,N_13461,N_12538);
and U17381 (N_17381,N_13218,N_12936);
or U17382 (N_17382,N_15301,N_12724);
nand U17383 (N_17383,N_12844,N_13869);
and U17384 (N_17384,N_13920,N_15562);
and U17385 (N_17385,N_13927,N_14870);
and U17386 (N_17386,N_13422,N_14140);
nor U17387 (N_17387,N_14923,N_12933);
nor U17388 (N_17388,N_12962,N_12605);
and U17389 (N_17389,N_13849,N_15295);
or U17390 (N_17390,N_14672,N_12688);
nor U17391 (N_17391,N_13066,N_14356);
nor U17392 (N_17392,N_13552,N_12743);
nor U17393 (N_17393,N_15145,N_12500);
or U17394 (N_17394,N_13272,N_13857);
or U17395 (N_17395,N_12956,N_13752);
or U17396 (N_17396,N_13646,N_14377);
and U17397 (N_17397,N_14481,N_15472);
nor U17398 (N_17398,N_15098,N_13182);
nand U17399 (N_17399,N_13466,N_14842);
nor U17400 (N_17400,N_13799,N_15336);
or U17401 (N_17401,N_14672,N_14784);
nor U17402 (N_17402,N_13519,N_13428);
or U17403 (N_17403,N_13133,N_14678);
and U17404 (N_17404,N_13723,N_15447);
or U17405 (N_17405,N_13642,N_12607);
nand U17406 (N_17406,N_13510,N_15578);
xnor U17407 (N_17407,N_13995,N_15120);
nor U17408 (N_17408,N_14603,N_15537);
or U17409 (N_17409,N_14339,N_15540);
xnor U17410 (N_17410,N_13067,N_12670);
xor U17411 (N_17411,N_14111,N_14237);
nor U17412 (N_17412,N_14164,N_14909);
nor U17413 (N_17413,N_13608,N_13634);
nand U17414 (N_17414,N_13149,N_13710);
xor U17415 (N_17415,N_13337,N_14625);
and U17416 (N_17416,N_14580,N_13336);
or U17417 (N_17417,N_13785,N_12790);
xor U17418 (N_17418,N_14335,N_14655);
and U17419 (N_17419,N_13674,N_13099);
and U17420 (N_17420,N_13643,N_14163);
and U17421 (N_17421,N_12658,N_15377);
or U17422 (N_17422,N_14661,N_13718);
nor U17423 (N_17423,N_14486,N_13344);
nor U17424 (N_17424,N_13061,N_12808);
nand U17425 (N_17425,N_14237,N_15080);
or U17426 (N_17426,N_14525,N_14847);
and U17427 (N_17427,N_13085,N_14825);
nand U17428 (N_17428,N_13120,N_12551);
nor U17429 (N_17429,N_14156,N_14135);
nand U17430 (N_17430,N_13035,N_12719);
and U17431 (N_17431,N_13514,N_15059);
nand U17432 (N_17432,N_13057,N_15036);
xor U17433 (N_17433,N_13387,N_15282);
or U17434 (N_17434,N_13149,N_13665);
and U17435 (N_17435,N_15150,N_13293);
and U17436 (N_17436,N_13066,N_14965);
and U17437 (N_17437,N_15410,N_14783);
or U17438 (N_17438,N_12776,N_13176);
nand U17439 (N_17439,N_14352,N_12537);
nor U17440 (N_17440,N_14208,N_14306);
xnor U17441 (N_17441,N_15061,N_15600);
nor U17442 (N_17442,N_13626,N_12776);
and U17443 (N_17443,N_13079,N_12953);
xor U17444 (N_17444,N_14919,N_12609);
or U17445 (N_17445,N_12758,N_14549);
nand U17446 (N_17446,N_13692,N_15455);
nand U17447 (N_17447,N_13588,N_13778);
nor U17448 (N_17448,N_14545,N_14979);
nor U17449 (N_17449,N_13738,N_14433);
or U17450 (N_17450,N_15354,N_15407);
or U17451 (N_17451,N_14275,N_14993);
and U17452 (N_17452,N_14394,N_13062);
and U17453 (N_17453,N_13132,N_14197);
or U17454 (N_17454,N_13038,N_15565);
or U17455 (N_17455,N_14591,N_13967);
or U17456 (N_17456,N_13207,N_15304);
nand U17457 (N_17457,N_14774,N_12978);
and U17458 (N_17458,N_14216,N_14770);
and U17459 (N_17459,N_13474,N_13313);
and U17460 (N_17460,N_13132,N_14709);
nor U17461 (N_17461,N_14446,N_12607);
xor U17462 (N_17462,N_15623,N_12521);
nand U17463 (N_17463,N_13836,N_14658);
and U17464 (N_17464,N_14391,N_15392);
or U17465 (N_17465,N_14001,N_14019);
or U17466 (N_17466,N_13740,N_15461);
nor U17467 (N_17467,N_13762,N_13187);
nand U17468 (N_17468,N_13160,N_12673);
or U17469 (N_17469,N_14208,N_13419);
and U17470 (N_17470,N_13907,N_13697);
nand U17471 (N_17471,N_13421,N_14512);
nor U17472 (N_17472,N_13824,N_13669);
and U17473 (N_17473,N_14094,N_14565);
nor U17474 (N_17474,N_14053,N_13654);
and U17475 (N_17475,N_12900,N_12808);
and U17476 (N_17476,N_14161,N_13889);
or U17477 (N_17477,N_14083,N_13097);
nand U17478 (N_17478,N_13520,N_13207);
or U17479 (N_17479,N_14695,N_12860);
nor U17480 (N_17480,N_14968,N_14629);
nor U17481 (N_17481,N_15249,N_12525);
nor U17482 (N_17482,N_15500,N_12781);
and U17483 (N_17483,N_13891,N_14207);
and U17484 (N_17484,N_14629,N_13418);
or U17485 (N_17485,N_15073,N_14475);
nand U17486 (N_17486,N_12720,N_15326);
and U17487 (N_17487,N_15152,N_15024);
nor U17488 (N_17488,N_13158,N_12506);
nor U17489 (N_17489,N_12583,N_13916);
nor U17490 (N_17490,N_14121,N_13891);
and U17491 (N_17491,N_12784,N_15019);
xnor U17492 (N_17492,N_13537,N_12589);
nor U17493 (N_17493,N_14373,N_14433);
nor U17494 (N_17494,N_12633,N_14704);
nand U17495 (N_17495,N_14952,N_15330);
nand U17496 (N_17496,N_15322,N_13051);
and U17497 (N_17497,N_13798,N_14917);
xnor U17498 (N_17498,N_12698,N_14388);
or U17499 (N_17499,N_13016,N_13007);
nor U17500 (N_17500,N_14599,N_13782);
nand U17501 (N_17501,N_13623,N_13984);
nor U17502 (N_17502,N_13238,N_14547);
xnor U17503 (N_17503,N_13500,N_12769);
or U17504 (N_17504,N_15239,N_14652);
nand U17505 (N_17505,N_13331,N_13094);
and U17506 (N_17506,N_13573,N_14419);
nand U17507 (N_17507,N_13093,N_13743);
and U17508 (N_17508,N_14855,N_13401);
nor U17509 (N_17509,N_12688,N_13740);
nor U17510 (N_17510,N_13899,N_14658);
or U17511 (N_17511,N_14035,N_13179);
or U17512 (N_17512,N_12773,N_12992);
nor U17513 (N_17513,N_13496,N_13897);
or U17514 (N_17514,N_13632,N_12686);
nor U17515 (N_17515,N_14898,N_15572);
or U17516 (N_17516,N_13263,N_13414);
and U17517 (N_17517,N_15322,N_14663);
or U17518 (N_17518,N_14550,N_13846);
and U17519 (N_17519,N_14931,N_15217);
or U17520 (N_17520,N_13654,N_14045);
and U17521 (N_17521,N_13699,N_13706);
and U17522 (N_17522,N_13851,N_14915);
or U17523 (N_17523,N_13954,N_15584);
nand U17524 (N_17524,N_15051,N_15561);
or U17525 (N_17525,N_12712,N_14324);
nor U17526 (N_17526,N_14098,N_12956);
nand U17527 (N_17527,N_14923,N_12872);
nand U17528 (N_17528,N_15123,N_15376);
nand U17529 (N_17529,N_13224,N_13025);
or U17530 (N_17530,N_12927,N_15508);
nor U17531 (N_17531,N_15167,N_15096);
or U17532 (N_17532,N_13623,N_13418);
or U17533 (N_17533,N_13470,N_15476);
nor U17534 (N_17534,N_14058,N_13600);
or U17535 (N_17535,N_15328,N_14337);
or U17536 (N_17536,N_13675,N_13989);
nand U17537 (N_17537,N_13546,N_14139);
nor U17538 (N_17538,N_15141,N_14977);
and U17539 (N_17539,N_13646,N_13379);
nor U17540 (N_17540,N_15240,N_13099);
or U17541 (N_17541,N_14911,N_13717);
and U17542 (N_17542,N_15142,N_14447);
nand U17543 (N_17543,N_14158,N_14539);
or U17544 (N_17544,N_15417,N_14474);
nor U17545 (N_17545,N_14029,N_15399);
nand U17546 (N_17546,N_13325,N_14477);
nor U17547 (N_17547,N_14058,N_13356);
and U17548 (N_17548,N_15162,N_13133);
nand U17549 (N_17549,N_13956,N_14611);
nand U17550 (N_17550,N_15033,N_12920);
nand U17551 (N_17551,N_13870,N_12716);
xor U17552 (N_17552,N_15461,N_15141);
and U17553 (N_17553,N_12771,N_14349);
and U17554 (N_17554,N_15075,N_14128);
or U17555 (N_17555,N_12774,N_13652);
xor U17556 (N_17556,N_12733,N_13239);
nor U17557 (N_17557,N_13161,N_13302);
and U17558 (N_17558,N_13369,N_12975);
and U17559 (N_17559,N_14640,N_14906);
or U17560 (N_17560,N_14329,N_12965);
nor U17561 (N_17561,N_12736,N_15471);
or U17562 (N_17562,N_14242,N_15301);
and U17563 (N_17563,N_14325,N_15604);
nand U17564 (N_17564,N_12971,N_15290);
nor U17565 (N_17565,N_13939,N_14406);
nor U17566 (N_17566,N_14744,N_13422);
nand U17567 (N_17567,N_15178,N_14860);
and U17568 (N_17568,N_14230,N_12985);
xor U17569 (N_17569,N_14392,N_15457);
nand U17570 (N_17570,N_15427,N_14826);
xor U17571 (N_17571,N_15567,N_13288);
nand U17572 (N_17572,N_13382,N_15039);
nor U17573 (N_17573,N_12876,N_15301);
or U17574 (N_17574,N_15172,N_15401);
and U17575 (N_17575,N_13724,N_15373);
and U17576 (N_17576,N_14946,N_12742);
xnor U17577 (N_17577,N_15484,N_14678);
or U17578 (N_17578,N_13195,N_14875);
or U17579 (N_17579,N_13344,N_14854);
nand U17580 (N_17580,N_15493,N_14168);
or U17581 (N_17581,N_14522,N_12648);
nor U17582 (N_17582,N_13798,N_12888);
nand U17583 (N_17583,N_15279,N_13522);
nor U17584 (N_17584,N_13080,N_14611);
and U17585 (N_17585,N_13746,N_14864);
and U17586 (N_17586,N_12895,N_14268);
nor U17587 (N_17587,N_13275,N_13357);
nand U17588 (N_17588,N_15271,N_13880);
xnor U17589 (N_17589,N_14092,N_13795);
or U17590 (N_17590,N_14124,N_14511);
nor U17591 (N_17591,N_13592,N_14896);
nand U17592 (N_17592,N_14329,N_14097);
nand U17593 (N_17593,N_14776,N_14007);
nand U17594 (N_17594,N_15206,N_13572);
nor U17595 (N_17595,N_13517,N_14697);
nor U17596 (N_17596,N_14557,N_12591);
nand U17597 (N_17597,N_14600,N_14655);
nor U17598 (N_17598,N_15347,N_14310);
nor U17599 (N_17599,N_13955,N_12989);
or U17600 (N_17600,N_14588,N_13408);
or U17601 (N_17601,N_14479,N_14280);
xnor U17602 (N_17602,N_15177,N_12835);
xnor U17603 (N_17603,N_13108,N_14878);
and U17604 (N_17604,N_14035,N_15118);
xor U17605 (N_17605,N_12969,N_12650);
and U17606 (N_17606,N_13773,N_15229);
nand U17607 (N_17607,N_13008,N_12999);
or U17608 (N_17608,N_15371,N_14490);
or U17609 (N_17609,N_12656,N_15155);
and U17610 (N_17610,N_13306,N_12906);
and U17611 (N_17611,N_14860,N_14251);
xnor U17612 (N_17612,N_15518,N_14816);
and U17613 (N_17613,N_14456,N_15419);
xnor U17614 (N_17614,N_14369,N_13284);
nand U17615 (N_17615,N_13225,N_14935);
or U17616 (N_17616,N_14984,N_15009);
xor U17617 (N_17617,N_12666,N_15292);
and U17618 (N_17618,N_14041,N_15570);
nand U17619 (N_17619,N_15162,N_13353);
nand U17620 (N_17620,N_12848,N_13599);
nor U17621 (N_17621,N_15332,N_15179);
nor U17622 (N_17622,N_14519,N_14701);
nand U17623 (N_17623,N_14744,N_14029);
or U17624 (N_17624,N_13361,N_15321);
or U17625 (N_17625,N_14002,N_14559);
or U17626 (N_17626,N_13870,N_13795);
xor U17627 (N_17627,N_14767,N_12546);
nor U17628 (N_17628,N_14675,N_15082);
xnor U17629 (N_17629,N_13026,N_14259);
or U17630 (N_17630,N_14352,N_14956);
and U17631 (N_17631,N_15577,N_14985);
or U17632 (N_17632,N_13313,N_14968);
nand U17633 (N_17633,N_15080,N_15254);
nor U17634 (N_17634,N_13860,N_13484);
nand U17635 (N_17635,N_15598,N_12604);
nor U17636 (N_17636,N_14331,N_15459);
and U17637 (N_17637,N_14088,N_14981);
or U17638 (N_17638,N_14260,N_13981);
xnor U17639 (N_17639,N_14070,N_13574);
or U17640 (N_17640,N_14744,N_15175);
nand U17641 (N_17641,N_13831,N_15314);
or U17642 (N_17642,N_14056,N_15321);
or U17643 (N_17643,N_12878,N_14114);
nand U17644 (N_17644,N_14472,N_13274);
nand U17645 (N_17645,N_15447,N_14738);
nand U17646 (N_17646,N_14713,N_13828);
nor U17647 (N_17647,N_15604,N_12730);
nor U17648 (N_17648,N_14722,N_13980);
nor U17649 (N_17649,N_15277,N_14559);
nor U17650 (N_17650,N_15247,N_15352);
or U17651 (N_17651,N_14667,N_12854);
nor U17652 (N_17652,N_14606,N_14351);
and U17653 (N_17653,N_14080,N_13095);
or U17654 (N_17654,N_14294,N_13953);
nand U17655 (N_17655,N_14116,N_12724);
or U17656 (N_17656,N_14162,N_12574);
or U17657 (N_17657,N_13834,N_13615);
or U17658 (N_17658,N_15402,N_14626);
nand U17659 (N_17659,N_12779,N_14828);
and U17660 (N_17660,N_14716,N_14715);
and U17661 (N_17661,N_15462,N_13561);
and U17662 (N_17662,N_15265,N_12794);
and U17663 (N_17663,N_13062,N_14133);
nor U17664 (N_17664,N_14129,N_12553);
nand U17665 (N_17665,N_14955,N_13398);
and U17666 (N_17666,N_13190,N_14862);
and U17667 (N_17667,N_13397,N_15373);
xor U17668 (N_17668,N_14998,N_13398);
nor U17669 (N_17669,N_14790,N_13736);
nor U17670 (N_17670,N_15575,N_12812);
or U17671 (N_17671,N_15042,N_13834);
nand U17672 (N_17672,N_14278,N_12594);
nor U17673 (N_17673,N_13276,N_14739);
nand U17674 (N_17674,N_14355,N_13443);
and U17675 (N_17675,N_15495,N_13612);
and U17676 (N_17676,N_14307,N_13061);
nor U17677 (N_17677,N_15122,N_13367);
xnor U17678 (N_17678,N_13525,N_15252);
or U17679 (N_17679,N_14250,N_13597);
nand U17680 (N_17680,N_15010,N_15089);
and U17681 (N_17681,N_15287,N_15160);
xnor U17682 (N_17682,N_14919,N_15360);
nand U17683 (N_17683,N_13787,N_12633);
and U17684 (N_17684,N_14518,N_12844);
or U17685 (N_17685,N_12694,N_14608);
nand U17686 (N_17686,N_14867,N_13612);
and U17687 (N_17687,N_13103,N_14032);
nor U17688 (N_17688,N_12553,N_13114);
or U17689 (N_17689,N_14608,N_15460);
or U17690 (N_17690,N_12790,N_15276);
or U17691 (N_17691,N_12931,N_12960);
xnor U17692 (N_17692,N_13316,N_13058);
or U17693 (N_17693,N_12723,N_15521);
and U17694 (N_17694,N_14985,N_15501);
or U17695 (N_17695,N_15062,N_13901);
or U17696 (N_17696,N_14757,N_13746);
xnor U17697 (N_17697,N_13999,N_14075);
or U17698 (N_17698,N_13371,N_15595);
and U17699 (N_17699,N_13458,N_14621);
and U17700 (N_17700,N_12565,N_15017);
nor U17701 (N_17701,N_15480,N_14639);
nor U17702 (N_17702,N_12803,N_15148);
nor U17703 (N_17703,N_14188,N_15321);
nand U17704 (N_17704,N_12608,N_12679);
nor U17705 (N_17705,N_13827,N_15049);
xnor U17706 (N_17706,N_12845,N_14603);
and U17707 (N_17707,N_13168,N_15164);
xor U17708 (N_17708,N_14332,N_14918);
and U17709 (N_17709,N_13460,N_15017);
and U17710 (N_17710,N_15140,N_13324);
or U17711 (N_17711,N_14361,N_14953);
or U17712 (N_17712,N_14929,N_15536);
and U17713 (N_17713,N_15063,N_13841);
nand U17714 (N_17714,N_14064,N_12658);
and U17715 (N_17715,N_13217,N_14926);
nand U17716 (N_17716,N_14341,N_15537);
and U17717 (N_17717,N_13454,N_13453);
and U17718 (N_17718,N_12789,N_14910);
nand U17719 (N_17719,N_12580,N_14295);
and U17720 (N_17720,N_13844,N_13334);
nor U17721 (N_17721,N_13311,N_13295);
and U17722 (N_17722,N_15064,N_14249);
nand U17723 (N_17723,N_14753,N_14737);
and U17724 (N_17724,N_15161,N_14233);
and U17725 (N_17725,N_15024,N_14162);
xnor U17726 (N_17726,N_13124,N_14833);
and U17727 (N_17727,N_14696,N_12501);
nand U17728 (N_17728,N_14734,N_14621);
or U17729 (N_17729,N_15085,N_14160);
xor U17730 (N_17730,N_14862,N_15192);
and U17731 (N_17731,N_13748,N_13679);
nor U17732 (N_17732,N_13211,N_13014);
and U17733 (N_17733,N_15403,N_15555);
or U17734 (N_17734,N_12528,N_14597);
nand U17735 (N_17735,N_13103,N_12909);
and U17736 (N_17736,N_13485,N_13145);
and U17737 (N_17737,N_14055,N_13983);
nand U17738 (N_17738,N_12832,N_14381);
and U17739 (N_17739,N_15540,N_12960);
or U17740 (N_17740,N_15557,N_14382);
nor U17741 (N_17741,N_12766,N_13072);
and U17742 (N_17742,N_13645,N_13877);
nor U17743 (N_17743,N_13892,N_13445);
nand U17744 (N_17744,N_15437,N_12691);
nand U17745 (N_17745,N_13891,N_13082);
and U17746 (N_17746,N_13200,N_13436);
xnor U17747 (N_17747,N_13467,N_14762);
xor U17748 (N_17748,N_13306,N_13843);
nand U17749 (N_17749,N_14111,N_12992);
nand U17750 (N_17750,N_15243,N_13346);
or U17751 (N_17751,N_13577,N_15072);
or U17752 (N_17752,N_12709,N_14268);
or U17753 (N_17753,N_13908,N_15394);
or U17754 (N_17754,N_14178,N_13687);
and U17755 (N_17755,N_13755,N_13268);
or U17756 (N_17756,N_13588,N_13404);
nor U17757 (N_17757,N_12527,N_13396);
or U17758 (N_17758,N_12838,N_13214);
nor U17759 (N_17759,N_15558,N_12871);
nor U17760 (N_17760,N_12872,N_15067);
nor U17761 (N_17761,N_12925,N_13654);
or U17762 (N_17762,N_12950,N_14771);
or U17763 (N_17763,N_13059,N_13548);
or U17764 (N_17764,N_13765,N_13991);
nand U17765 (N_17765,N_14287,N_12830);
or U17766 (N_17766,N_14036,N_13745);
or U17767 (N_17767,N_13057,N_13225);
and U17768 (N_17768,N_14821,N_12898);
nand U17769 (N_17769,N_15065,N_14675);
and U17770 (N_17770,N_13007,N_15277);
nand U17771 (N_17771,N_14938,N_13820);
xnor U17772 (N_17772,N_14432,N_14494);
nand U17773 (N_17773,N_13823,N_14040);
nor U17774 (N_17774,N_14711,N_13750);
xor U17775 (N_17775,N_14625,N_15126);
or U17776 (N_17776,N_15477,N_13224);
nand U17777 (N_17777,N_14102,N_14044);
and U17778 (N_17778,N_14329,N_13812);
and U17779 (N_17779,N_15134,N_13636);
or U17780 (N_17780,N_13060,N_15125);
and U17781 (N_17781,N_13102,N_12716);
xor U17782 (N_17782,N_12925,N_15176);
and U17783 (N_17783,N_14919,N_15070);
xor U17784 (N_17784,N_14469,N_15556);
nor U17785 (N_17785,N_13516,N_13740);
or U17786 (N_17786,N_12515,N_13735);
and U17787 (N_17787,N_14907,N_15082);
nand U17788 (N_17788,N_12981,N_13812);
or U17789 (N_17789,N_13984,N_15155);
and U17790 (N_17790,N_12733,N_15182);
or U17791 (N_17791,N_13216,N_15379);
and U17792 (N_17792,N_13101,N_12773);
and U17793 (N_17793,N_13583,N_13762);
nand U17794 (N_17794,N_13110,N_15265);
and U17795 (N_17795,N_15078,N_13402);
nor U17796 (N_17796,N_14712,N_12952);
or U17797 (N_17797,N_14716,N_15581);
nand U17798 (N_17798,N_13129,N_14787);
xnor U17799 (N_17799,N_12876,N_15324);
nor U17800 (N_17800,N_13114,N_14218);
and U17801 (N_17801,N_14158,N_15214);
nor U17802 (N_17802,N_15352,N_15269);
nor U17803 (N_17803,N_13681,N_15380);
and U17804 (N_17804,N_15112,N_13741);
nand U17805 (N_17805,N_13908,N_14628);
nor U17806 (N_17806,N_15528,N_12554);
or U17807 (N_17807,N_14009,N_14983);
xor U17808 (N_17808,N_14115,N_12524);
nor U17809 (N_17809,N_14951,N_14480);
and U17810 (N_17810,N_12524,N_14066);
nor U17811 (N_17811,N_15142,N_12843);
nand U17812 (N_17812,N_13709,N_14087);
and U17813 (N_17813,N_14455,N_13462);
and U17814 (N_17814,N_14389,N_15505);
xor U17815 (N_17815,N_12627,N_15567);
xor U17816 (N_17816,N_15167,N_15500);
and U17817 (N_17817,N_14802,N_14878);
nand U17818 (N_17818,N_14158,N_12981);
or U17819 (N_17819,N_14407,N_14483);
and U17820 (N_17820,N_13103,N_12639);
nand U17821 (N_17821,N_14288,N_13100);
or U17822 (N_17822,N_15462,N_15457);
nand U17823 (N_17823,N_13981,N_14570);
nor U17824 (N_17824,N_14610,N_13151);
nor U17825 (N_17825,N_12735,N_15502);
or U17826 (N_17826,N_14978,N_13805);
nor U17827 (N_17827,N_13536,N_12853);
xnor U17828 (N_17828,N_15276,N_15452);
nand U17829 (N_17829,N_14694,N_14586);
nand U17830 (N_17830,N_15328,N_12899);
or U17831 (N_17831,N_13036,N_13053);
nand U17832 (N_17832,N_14593,N_14917);
nand U17833 (N_17833,N_14974,N_13360);
nor U17834 (N_17834,N_13677,N_14066);
xnor U17835 (N_17835,N_14723,N_14706);
nand U17836 (N_17836,N_13378,N_14656);
nand U17837 (N_17837,N_15491,N_14199);
and U17838 (N_17838,N_13210,N_13275);
nor U17839 (N_17839,N_13826,N_14834);
and U17840 (N_17840,N_14268,N_13350);
and U17841 (N_17841,N_14624,N_12654);
or U17842 (N_17842,N_14309,N_13946);
and U17843 (N_17843,N_13699,N_12572);
nand U17844 (N_17844,N_13762,N_15209);
nand U17845 (N_17845,N_13639,N_15153);
nor U17846 (N_17846,N_15021,N_13385);
or U17847 (N_17847,N_14260,N_14014);
xor U17848 (N_17848,N_12832,N_15078);
or U17849 (N_17849,N_12765,N_15240);
xnor U17850 (N_17850,N_12990,N_14350);
nor U17851 (N_17851,N_15584,N_13534);
or U17852 (N_17852,N_14319,N_12714);
or U17853 (N_17853,N_14440,N_14825);
or U17854 (N_17854,N_14468,N_14615);
and U17855 (N_17855,N_14481,N_14554);
xor U17856 (N_17856,N_14378,N_13045);
and U17857 (N_17857,N_15029,N_15595);
or U17858 (N_17858,N_13933,N_14410);
or U17859 (N_17859,N_12501,N_14339);
and U17860 (N_17860,N_15381,N_14302);
or U17861 (N_17861,N_13797,N_15139);
and U17862 (N_17862,N_13648,N_15061);
and U17863 (N_17863,N_13812,N_13045);
nand U17864 (N_17864,N_13798,N_12943);
nor U17865 (N_17865,N_13143,N_13898);
or U17866 (N_17866,N_13125,N_15497);
and U17867 (N_17867,N_14812,N_15207);
nor U17868 (N_17868,N_13672,N_14787);
and U17869 (N_17869,N_14569,N_13573);
or U17870 (N_17870,N_12694,N_12601);
and U17871 (N_17871,N_14497,N_15468);
and U17872 (N_17872,N_15286,N_13414);
xnor U17873 (N_17873,N_15141,N_12741);
or U17874 (N_17874,N_14337,N_12920);
and U17875 (N_17875,N_13934,N_15140);
nand U17876 (N_17876,N_12766,N_13711);
nand U17877 (N_17877,N_13329,N_14693);
and U17878 (N_17878,N_14183,N_14548);
or U17879 (N_17879,N_15579,N_13674);
and U17880 (N_17880,N_13567,N_15142);
and U17881 (N_17881,N_14319,N_15147);
or U17882 (N_17882,N_13475,N_12731);
xnor U17883 (N_17883,N_14305,N_12570);
xor U17884 (N_17884,N_13076,N_13238);
nand U17885 (N_17885,N_13863,N_13186);
nor U17886 (N_17886,N_13869,N_13439);
or U17887 (N_17887,N_14289,N_14540);
and U17888 (N_17888,N_14765,N_14178);
nor U17889 (N_17889,N_14001,N_13571);
and U17890 (N_17890,N_13645,N_13283);
nor U17891 (N_17891,N_12617,N_12999);
nand U17892 (N_17892,N_14877,N_12829);
and U17893 (N_17893,N_12718,N_15016);
nor U17894 (N_17894,N_14941,N_13819);
nor U17895 (N_17895,N_15537,N_13645);
nor U17896 (N_17896,N_13718,N_15420);
nor U17897 (N_17897,N_14376,N_14745);
nand U17898 (N_17898,N_12772,N_15507);
nor U17899 (N_17899,N_12900,N_14960);
or U17900 (N_17900,N_13593,N_12546);
and U17901 (N_17901,N_14412,N_12885);
nand U17902 (N_17902,N_12975,N_14806);
and U17903 (N_17903,N_13533,N_14382);
nand U17904 (N_17904,N_12644,N_14342);
nand U17905 (N_17905,N_14032,N_13302);
xor U17906 (N_17906,N_14545,N_13255);
nor U17907 (N_17907,N_15414,N_12926);
or U17908 (N_17908,N_13137,N_15262);
or U17909 (N_17909,N_12966,N_14839);
and U17910 (N_17910,N_15194,N_14507);
nand U17911 (N_17911,N_13195,N_15180);
nor U17912 (N_17912,N_13121,N_14160);
or U17913 (N_17913,N_15102,N_13506);
or U17914 (N_17914,N_13566,N_13172);
xnor U17915 (N_17915,N_15072,N_14158);
or U17916 (N_17916,N_13998,N_12500);
and U17917 (N_17917,N_12548,N_14199);
and U17918 (N_17918,N_15448,N_15575);
or U17919 (N_17919,N_13381,N_13156);
and U17920 (N_17920,N_14400,N_13506);
or U17921 (N_17921,N_14910,N_15564);
nor U17922 (N_17922,N_14868,N_13632);
or U17923 (N_17923,N_14888,N_14069);
xnor U17924 (N_17924,N_14110,N_13448);
or U17925 (N_17925,N_12583,N_14545);
or U17926 (N_17926,N_13976,N_12863);
and U17927 (N_17927,N_14182,N_12693);
and U17928 (N_17928,N_13870,N_13027);
and U17929 (N_17929,N_13853,N_14233);
nand U17930 (N_17930,N_13461,N_13928);
nor U17931 (N_17931,N_13521,N_12847);
xor U17932 (N_17932,N_12516,N_12758);
nor U17933 (N_17933,N_14828,N_14010);
nand U17934 (N_17934,N_15142,N_13725);
nor U17935 (N_17935,N_13887,N_14055);
and U17936 (N_17936,N_12817,N_15617);
nand U17937 (N_17937,N_13126,N_13923);
xnor U17938 (N_17938,N_14700,N_13315);
nand U17939 (N_17939,N_13056,N_14425);
or U17940 (N_17940,N_14337,N_14984);
or U17941 (N_17941,N_13760,N_12855);
and U17942 (N_17942,N_14803,N_13275);
or U17943 (N_17943,N_13640,N_14674);
or U17944 (N_17944,N_12807,N_14759);
and U17945 (N_17945,N_15511,N_14095);
nor U17946 (N_17946,N_15257,N_15363);
nor U17947 (N_17947,N_12821,N_13449);
nor U17948 (N_17948,N_15609,N_15266);
or U17949 (N_17949,N_13905,N_12720);
nor U17950 (N_17950,N_13652,N_13345);
or U17951 (N_17951,N_15129,N_13588);
and U17952 (N_17952,N_14982,N_15041);
nor U17953 (N_17953,N_12525,N_15156);
xnor U17954 (N_17954,N_14495,N_12780);
nand U17955 (N_17955,N_13391,N_15469);
nand U17956 (N_17956,N_12946,N_14865);
or U17957 (N_17957,N_13419,N_14807);
nand U17958 (N_17958,N_12728,N_14322);
and U17959 (N_17959,N_14067,N_15413);
xnor U17960 (N_17960,N_15539,N_14947);
and U17961 (N_17961,N_13172,N_13978);
and U17962 (N_17962,N_12649,N_13888);
nor U17963 (N_17963,N_14602,N_14002);
and U17964 (N_17964,N_12652,N_14880);
or U17965 (N_17965,N_13396,N_14642);
and U17966 (N_17966,N_13805,N_14340);
xor U17967 (N_17967,N_12791,N_12632);
nand U17968 (N_17968,N_13718,N_13550);
or U17969 (N_17969,N_13692,N_13850);
nor U17970 (N_17970,N_13947,N_14700);
nand U17971 (N_17971,N_12622,N_15169);
and U17972 (N_17972,N_12653,N_14668);
and U17973 (N_17973,N_15051,N_15111);
nand U17974 (N_17974,N_13933,N_12688);
and U17975 (N_17975,N_12702,N_14257);
nor U17976 (N_17976,N_12989,N_12836);
and U17977 (N_17977,N_14499,N_15326);
nand U17978 (N_17978,N_13720,N_13040);
and U17979 (N_17979,N_14063,N_14023);
nand U17980 (N_17980,N_13391,N_14936);
nand U17981 (N_17981,N_13330,N_15025);
nand U17982 (N_17982,N_14305,N_13438);
nor U17983 (N_17983,N_13983,N_12762);
xnor U17984 (N_17984,N_14728,N_14401);
and U17985 (N_17985,N_13806,N_13245);
xnor U17986 (N_17986,N_13376,N_15576);
nor U17987 (N_17987,N_14979,N_14543);
and U17988 (N_17988,N_14529,N_13674);
nand U17989 (N_17989,N_15620,N_13546);
nand U17990 (N_17990,N_14488,N_14321);
nand U17991 (N_17991,N_13363,N_14510);
or U17992 (N_17992,N_13278,N_15449);
and U17993 (N_17993,N_15493,N_15265);
nor U17994 (N_17994,N_13728,N_14724);
nand U17995 (N_17995,N_14875,N_13975);
xnor U17996 (N_17996,N_14542,N_14245);
or U17997 (N_17997,N_14620,N_14334);
nor U17998 (N_17998,N_12756,N_13442);
xor U17999 (N_17999,N_14054,N_12640);
and U18000 (N_18000,N_15102,N_14371);
or U18001 (N_18001,N_14380,N_14455);
nand U18002 (N_18002,N_15560,N_14588);
or U18003 (N_18003,N_14747,N_15304);
or U18004 (N_18004,N_13862,N_13604);
xnor U18005 (N_18005,N_14228,N_14550);
nand U18006 (N_18006,N_13650,N_14773);
nor U18007 (N_18007,N_13804,N_14340);
or U18008 (N_18008,N_13308,N_13532);
nand U18009 (N_18009,N_12909,N_13839);
and U18010 (N_18010,N_12835,N_14735);
and U18011 (N_18011,N_15312,N_13639);
or U18012 (N_18012,N_12614,N_13813);
and U18013 (N_18013,N_15249,N_14879);
and U18014 (N_18014,N_12538,N_15121);
and U18015 (N_18015,N_14208,N_12633);
nand U18016 (N_18016,N_14908,N_12783);
and U18017 (N_18017,N_13879,N_14997);
and U18018 (N_18018,N_14419,N_15586);
xnor U18019 (N_18019,N_13834,N_13153);
and U18020 (N_18020,N_14892,N_12597);
or U18021 (N_18021,N_14736,N_13479);
and U18022 (N_18022,N_12816,N_14684);
nand U18023 (N_18023,N_13358,N_13304);
nand U18024 (N_18024,N_13219,N_14479);
nand U18025 (N_18025,N_13643,N_13876);
or U18026 (N_18026,N_13410,N_13025);
xor U18027 (N_18027,N_13081,N_13117);
nor U18028 (N_18028,N_14402,N_15003);
or U18029 (N_18029,N_14319,N_13173);
or U18030 (N_18030,N_14962,N_15197);
nand U18031 (N_18031,N_13301,N_13955);
and U18032 (N_18032,N_15363,N_13457);
and U18033 (N_18033,N_13999,N_13153);
and U18034 (N_18034,N_13091,N_15300);
xor U18035 (N_18035,N_14447,N_14779);
nor U18036 (N_18036,N_13175,N_12932);
or U18037 (N_18037,N_15182,N_13165);
or U18038 (N_18038,N_14710,N_13021);
xor U18039 (N_18039,N_14182,N_12813);
and U18040 (N_18040,N_14203,N_13703);
and U18041 (N_18041,N_13407,N_14519);
nor U18042 (N_18042,N_13347,N_14386);
and U18043 (N_18043,N_12971,N_15298);
and U18044 (N_18044,N_13800,N_15014);
and U18045 (N_18045,N_13111,N_14312);
nor U18046 (N_18046,N_13726,N_14267);
nor U18047 (N_18047,N_15400,N_13421);
or U18048 (N_18048,N_13300,N_15623);
and U18049 (N_18049,N_13655,N_13710);
or U18050 (N_18050,N_13520,N_14950);
or U18051 (N_18051,N_12901,N_13217);
and U18052 (N_18052,N_14792,N_12537);
or U18053 (N_18053,N_15620,N_13048);
or U18054 (N_18054,N_12984,N_14534);
and U18055 (N_18055,N_12999,N_15617);
and U18056 (N_18056,N_14693,N_14075);
and U18057 (N_18057,N_14328,N_14237);
nor U18058 (N_18058,N_14004,N_12546);
nor U18059 (N_18059,N_13305,N_14668);
nand U18060 (N_18060,N_15229,N_14678);
or U18061 (N_18061,N_14823,N_14674);
or U18062 (N_18062,N_13412,N_12737);
and U18063 (N_18063,N_13397,N_14964);
and U18064 (N_18064,N_14588,N_14345);
nand U18065 (N_18065,N_14596,N_13540);
or U18066 (N_18066,N_14746,N_14335);
nor U18067 (N_18067,N_13766,N_13525);
and U18068 (N_18068,N_14309,N_12734);
nand U18069 (N_18069,N_12945,N_15324);
or U18070 (N_18070,N_14726,N_15137);
xor U18071 (N_18071,N_14118,N_13938);
nand U18072 (N_18072,N_14794,N_12515);
nor U18073 (N_18073,N_14179,N_14891);
nand U18074 (N_18074,N_15241,N_15062);
nand U18075 (N_18075,N_15091,N_14866);
and U18076 (N_18076,N_14590,N_14303);
xor U18077 (N_18077,N_13981,N_12649);
nand U18078 (N_18078,N_14082,N_12931);
nand U18079 (N_18079,N_15258,N_13420);
nand U18080 (N_18080,N_12869,N_14012);
nand U18081 (N_18081,N_13677,N_13017);
or U18082 (N_18082,N_13857,N_13694);
or U18083 (N_18083,N_15148,N_13529);
xnor U18084 (N_18084,N_14384,N_15589);
and U18085 (N_18085,N_13573,N_13548);
and U18086 (N_18086,N_13868,N_14118);
nor U18087 (N_18087,N_13937,N_14351);
nor U18088 (N_18088,N_12948,N_14217);
and U18089 (N_18089,N_13849,N_15025);
or U18090 (N_18090,N_14930,N_13088);
or U18091 (N_18091,N_14963,N_15360);
xor U18092 (N_18092,N_13174,N_15062);
nor U18093 (N_18093,N_13894,N_14621);
nand U18094 (N_18094,N_13549,N_15233);
or U18095 (N_18095,N_14776,N_13061);
nor U18096 (N_18096,N_13699,N_13376);
nor U18097 (N_18097,N_15369,N_14069);
and U18098 (N_18098,N_14703,N_13948);
and U18099 (N_18099,N_14565,N_13314);
nand U18100 (N_18100,N_15348,N_12714);
and U18101 (N_18101,N_15330,N_12520);
and U18102 (N_18102,N_13640,N_13227);
nand U18103 (N_18103,N_14736,N_13819);
nor U18104 (N_18104,N_12797,N_13122);
and U18105 (N_18105,N_14422,N_14677);
nor U18106 (N_18106,N_15611,N_14895);
and U18107 (N_18107,N_15110,N_14711);
nor U18108 (N_18108,N_12788,N_14504);
xor U18109 (N_18109,N_12846,N_14281);
nor U18110 (N_18110,N_12663,N_15290);
and U18111 (N_18111,N_12788,N_14340);
nor U18112 (N_18112,N_13509,N_14166);
xor U18113 (N_18113,N_15505,N_13247);
or U18114 (N_18114,N_12954,N_15569);
nand U18115 (N_18115,N_15615,N_14599);
nand U18116 (N_18116,N_13971,N_13372);
and U18117 (N_18117,N_14173,N_13836);
or U18118 (N_18118,N_13071,N_12646);
nor U18119 (N_18119,N_14835,N_14352);
and U18120 (N_18120,N_13031,N_13235);
or U18121 (N_18121,N_15578,N_14473);
and U18122 (N_18122,N_13727,N_14921);
and U18123 (N_18123,N_13940,N_12740);
nand U18124 (N_18124,N_12514,N_13157);
nand U18125 (N_18125,N_13039,N_14072);
nor U18126 (N_18126,N_14048,N_12740);
xnor U18127 (N_18127,N_13641,N_14199);
nor U18128 (N_18128,N_12812,N_14360);
and U18129 (N_18129,N_13292,N_14522);
and U18130 (N_18130,N_12798,N_14099);
nand U18131 (N_18131,N_12515,N_15145);
and U18132 (N_18132,N_13453,N_14208);
or U18133 (N_18133,N_13028,N_13338);
or U18134 (N_18134,N_13502,N_15387);
nand U18135 (N_18135,N_14835,N_14358);
nor U18136 (N_18136,N_14680,N_14159);
nor U18137 (N_18137,N_14899,N_15245);
or U18138 (N_18138,N_14894,N_14426);
xnor U18139 (N_18139,N_14714,N_13634);
or U18140 (N_18140,N_15006,N_14680);
nand U18141 (N_18141,N_12989,N_14199);
nand U18142 (N_18142,N_15289,N_13268);
xor U18143 (N_18143,N_13972,N_14244);
xor U18144 (N_18144,N_12793,N_12812);
xor U18145 (N_18145,N_13280,N_12576);
xnor U18146 (N_18146,N_12871,N_14626);
nand U18147 (N_18147,N_13891,N_13718);
and U18148 (N_18148,N_12514,N_14633);
nand U18149 (N_18149,N_14075,N_13467);
xnor U18150 (N_18150,N_13627,N_14006);
or U18151 (N_18151,N_15500,N_13920);
and U18152 (N_18152,N_13981,N_14331);
and U18153 (N_18153,N_13485,N_13122);
xor U18154 (N_18154,N_14714,N_15394);
xnor U18155 (N_18155,N_15397,N_15043);
nand U18156 (N_18156,N_13816,N_14535);
and U18157 (N_18157,N_13018,N_13571);
nor U18158 (N_18158,N_15131,N_14981);
nand U18159 (N_18159,N_15504,N_14148);
nor U18160 (N_18160,N_14679,N_14320);
nand U18161 (N_18161,N_13702,N_15540);
and U18162 (N_18162,N_13407,N_13697);
nand U18163 (N_18163,N_12810,N_14940);
nor U18164 (N_18164,N_12967,N_13431);
xor U18165 (N_18165,N_15099,N_13619);
xor U18166 (N_18166,N_14622,N_14403);
and U18167 (N_18167,N_13952,N_14102);
or U18168 (N_18168,N_12866,N_15264);
and U18169 (N_18169,N_13828,N_14026);
nor U18170 (N_18170,N_14346,N_12795);
nor U18171 (N_18171,N_14691,N_14404);
nand U18172 (N_18172,N_14416,N_15569);
or U18173 (N_18173,N_13179,N_14880);
nor U18174 (N_18174,N_13067,N_14715);
nand U18175 (N_18175,N_13421,N_14884);
or U18176 (N_18176,N_14473,N_13829);
or U18177 (N_18177,N_13004,N_13510);
nand U18178 (N_18178,N_15130,N_14666);
nand U18179 (N_18179,N_14853,N_15194);
nand U18180 (N_18180,N_12867,N_12639);
and U18181 (N_18181,N_14772,N_13723);
nor U18182 (N_18182,N_13222,N_15524);
xnor U18183 (N_18183,N_13684,N_14043);
and U18184 (N_18184,N_13120,N_14401);
nor U18185 (N_18185,N_14329,N_13901);
and U18186 (N_18186,N_13174,N_13471);
nand U18187 (N_18187,N_14134,N_14710);
nor U18188 (N_18188,N_15195,N_14750);
or U18189 (N_18189,N_13782,N_14371);
nor U18190 (N_18190,N_13197,N_14054);
or U18191 (N_18191,N_14547,N_12514);
nand U18192 (N_18192,N_14147,N_12811);
nor U18193 (N_18193,N_15575,N_13205);
or U18194 (N_18194,N_13951,N_15074);
or U18195 (N_18195,N_13118,N_14106);
and U18196 (N_18196,N_12994,N_14851);
and U18197 (N_18197,N_13777,N_13945);
or U18198 (N_18198,N_13354,N_15599);
and U18199 (N_18199,N_13938,N_13079);
nor U18200 (N_18200,N_14213,N_15175);
xor U18201 (N_18201,N_12751,N_15553);
nand U18202 (N_18202,N_13695,N_13583);
nand U18203 (N_18203,N_14714,N_14301);
nand U18204 (N_18204,N_15207,N_13296);
and U18205 (N_18205,N_15601,N_12793);
or U18206 (N_18206,N_12530,N_13927);
xnor U18207 (N_18207,N_14386,N_12933);
and U18208 (N_18208,N_14595,N_13175);
and U18209 (N_18209,N_14082,N_13816);
or U18210 (N_18210,N_15152,N_12534);
nand U18211 (N_18211,N_15559,N_15191);
nand U18212 (N_18212,N_13264,N_12803);
and U18213 (N_18213,N_14843,N_12712);
or U18214 (N_18214,N_12779,N_12789);
nand U18215 (N_18215,N_15616,N_13935);
nand U18216 (N_18216,N_12783,N_12544);
nor U18217 (N_18217,N_14144,N_15573);
nand U18218 (N_18218,N_13439,N_13726);
or U18219 (N_18219,N_13293,N_13168);
nand U18220 (N_18220,N_13033,N_14221);
and U18221 (N_18221,N_14572,N_14818);
nor U18222 (N_18222,N_13833,N_13329);
or U18223 (N_18223,N_14405,N_15617);
nor U18224 (N_18224,N_13298,N_14227);
and U18225 (N_18225,N_15381,N_13429);
nand U18226 (N_18226,N_14430,N_14748);
nand U18227 (N_18227,N_13206,N_15311);
nor U18228 (N_18228,N_15076,N_15582);
and U18229 (N_18229,N_13766,N_13928);
nand U18230 (N_18230,N_14674,N_15144);
nand U18231 (N_18231,N_14979,N_14105);
nor U18232 (N_18232,N_12549,N_14103);
or U18233 (N_18233,N_15362,N_14146);
and U18234 (N_18234,N_14267,N_15065);
or U18235 (N_18235,N_14655,N_13293);
or U18236 (N_18236,N_14629,N_14029);
nand U18237 (N_18237,N_13423,N_15057);
nand U18238 (N_18238,N_13595,N_15508);
nand U18239 (N_18239,N_12937,N_14515);
and U18240 (N_18240,N_15231,N_13357);
nand U18241 (N_18241,N_13170,N_15113);
and U18242 (N_18242,N_13503,N_14589);
nor U18243 (N_18243,N_14202,N_14755);
nor U18244 (N_18244,N_15495,N_13133);
or U18245 (N_18245,N_13654,N_14273);
and U18246 (N_18246,N_13819,N_14800);
nand U18247 (N_18247,N_14896,N_15217);
or U18248 (N_18248,N_15077,N_14055);
xor U18249 (N_18249,N_15402,N_14280);
nor U18250 (N_18250,N_13872,N_14859);
or U18251 (N_18251,N_14423,N_15073);
and U18252 (N_18252,N_15313,N_12752);
nand U18253 (N_18253,N_13214,N_15298);
and U18254 (N_18254,N_15368,N_13765);
nor U18255 (N_18255,N_14001,N_14578);
nor U18256 (N_18256,N_13812,N_12884);
nor U18257 (N_18257,N_13058,N_13929);
xor U18258 (N_18258,N_12915,N_15281);
nor U18259 (N_18259,N_14723,N_15254);
xor U18260 (N_18260,N_15150,N_15229);
xnor U18261 (N_18261,N_13898,N_14298);
and U18262 (N_18262,N_14424,N_13164);
and U18263 (N_18263,N_15277,N_12918);
or U18264 (N_18264,N_14299,N_15183);
and U18265 (N_18265,N_12795,N_14184);
xor U18266 (N_18266,N_13157,N_13593);
or U18267 (N_18267,N_15473,N_14382);
or U18268 (N_18268,N_12708,N_13939);
or U18269 (N_18269,N_14365,N_13929);
and U18270 (N_18270,N_13374,N_15561);
nor U18271 (N_18271,N_14615,N_14734);
nand U18272 (N_18272,N_15325,N_15431);
or U18273 (N_18273,N_14485,N_13520);
nor U18274 (N_18274,N_14049,N_12693);
and U18275 (N_18275,N_13919,N_14634);
or U18276 (N_18276,N_13941,N_13205);
and U18277 (N_18277,N_13884,N_15106);
or U18278 (N_18278,N_13112,N_12609);
and U18279 (N_18279,N_13136,N_15458);
and U18280 (N_18280,N_13751,N_12889);
and U18281 (N_18281,N_15381,N_13544);
nor U18282 (N_18282,N_12743,N_13252);
or U18283 (N_18283,N_13147,N_12626);
nor U18284 (N_18284,N_15444,N_12974);
nand U18285 (N_18285,N_14840,N_12721);
nand U18286 (N_18286,N_14747,N_14587);
or U18287 (N_18287,N_13886,N_13777);
and U18288 (N_18288,N_14226,N_15525);
nor U18289 (N_18289,N_15362,N_14958);
and U18290 (N_18290,N_12876,N_15388);
nor U18291 (N_18291,N_14352,N_13715);
xor U18292 (N_18292,N_13129,N_14545);
or U18293 (N_18293,N_14711,N_12993);
nor U18294 (N_18294,N_15191,N_15101);
nor U18295 (N_18295,N_14128,N_15515);
nand U18296 (N_18296,N_14424,N_14716);
or U18297 (N_18297,N_12636,N_13442);
or U18298 (N_18298,N_13450,N_13368);
nand U18299 (N_18299,N_14343,N_13496);
nand U18300 (N_18300,N_12954,N_15539);
nor U18301 (N_18301,N_13403,N_14084);
nand U18302 (N_18302,N_13848,N_12773);
nand U18303 (N_18303,N_13091,N_13791);
nor U18304 (N_18304,N_13236,N_14848);
and U18305 (N_18305,N_14205,N_14603);
and U18306 (N_18306,N_12872,N_13439);
or U18307 (N_18307,N_14391,N_12625);
nor U18308 (N_18308,N_13146,N_12869);
nand U18309 (N_18309,N_13809,N_13405);
and U18310 (N_18310,N_15088,N_12990);
nor U18311 (N_18311,N_15574,N_15473);
nand U18312 (N_18312,N_12757,N_15174);
and U18313 (N_18313,N_12930,N_14160);
xnor U18314 (N_18314,N_14815,N_14123);
nand U18315 (N_18315,N_15036,N_15436);
nor U18316 (N_18316,N_14366,N_13734);
nor U18317 (N_18317,N_14835,N_12650);
nor U18318 (N_18318,N_15570,N_14952);
or U18319 (N_18319,N_12521,N_13381);
nand U18320 (N_18320,N_13242,N_14056);
nand U18321 (N_18321,N_13640,N_12835);
xor U18322 (N_18322,N_14491,N_13903);
xnor U18323 (N_18323,N_14437,N_13680);
or U18324 (N_18324,N_14642,N_13309);
or U18325 (N_18325,N_15559,N_13864);
nand U18326 (N_18326,N_14381,N_12613);
xnor U18327 (N_18327,N_15048,N_12688);
nor U18328 (N_18328,N_14088,N_15369);
and U18329 (N_18329,N_14225,N_15012);
nor U18330 (N_18330,N_13828,N_12532);
nand U18331 (N_18331,N_13466,N_13367);
nand U18332 (N_18332,N_14059,N_14693);
or U18333 (N_18333,N_12720,N_12844);
xnor U18334 (N_18334,N_13858,N_14484);
nand U18335 (N_18335,N_14184,N_14728);
nor U18336 (N_18336,N_12691,N_13752);
and U18337 (N_18337,N_14674,N_14608);
and U18338 (N_18338,N_15181,N_15038);
and U18339 (N_18339,N_15570,N_15397);
or U18340 (N_18340,N_12816,N_13079);
nand U18341 (N_18341,N_13299,N_15129);
nor U18342 (N_18342,N_12903,N_13885);
xor U18343 (N_18343,N_14422,N_13149);
nor U18344 (N_18344,N_13929,N_15372);
nor U18345 (N_18345,N_14364,N_14540);
nand U18346 (N_18346,N_15294,N_13011);
and U18347 (N_18347,N_15383,N_14684);
nand U18348 (N_18348,N_13778,N_13382);
and U18349 (N_18349,N_15114,N_12575);
nand U18350 (N_18350,N_13107,N_15266);
xor U18351 (N_18351,N_15251,N_13138);
or U18352 (N_18352,N_13625,N_12839);
or U18353 (N_18353,N_14300,N_14346);
or U18354 (N_18354,N_15552,N_13498);
or U18355 (N_18355,N_12964,N_12800);
and U18356 (N_18356,N_14120,N_15484);
and U18357 (N_18357,N_14965,N_13573);
nor U18358 (N_18358,N_13409,N_13555);
nor U18359 (N_18359,N_14786,N_14749);
xnor U18360 (N_18360,N_14419,N_15482);
and U18361 (N_18361,N_15611,N_13007);
nand U18362 (N_18362,N_14266,N_13982);
nor U18363 (N_18363,N_13675,N_15257);
or U18364 (N_18364,N_14543,N_14884);
or U18365 (N_18365,N_14370,N_13193);
or U18366 (N_18366,N_14891,N_14778);
or U18367 (N_18367,N_14325,N_13867);
xor U18368 (N_18368,N_14206,N_15171);
or U18369 (N_18369,N_14724,N_14476);
nor U18370 (N_18370,N_13766,N_12592);
and U18371 (N_18371,N_14017,N_14232);
nand U18372 (N_18372,N_12723,N_15163);
or U18373 (N_18373,N_14358,N_12503);
and U18374 (N_18374,N_15054,N_14444);
and U18375 (N_18375,N_13186,N_12539);
nor U18376 (N_18376,N_14708,N_13972);
and U18377 (N_18377,N_13632,N_12841);
or U18378 (N_18378,N_15426,N_15590);
and U18379 (N_18379,N_15173,N_14902);
nand U18380 (N_18380,N_14470,N_14448);
and U18381 (N_18381,N_14305,N_15265);
or U18382 (N_18382,N_14096,N_14141);
or U18383 (N_18383,N_15269,N_12901);
and U18384 (N_18384,N_12715,N_14022);
xor U18385 (N_18385,N_13993,N_13465);
xnor U18386 (N_18386,N_13395,N_14686);
nand U18387 (N_18387,N_13365,N_15374);
nor U18388 (N_18388,N_13436,N_13652);
or U18389 (N_18389,N_14984,N_13550);
xnor U18390 (N_18390,N_14831,N_14897);
and U18391 (N_18391,N_13927,N_12727);
and U18392 (N_18392,N_14777,N_13241);
nor U18393 (N_18393,N_13531,N_12608);
and U18394 (N_18394,N_12589,N_12746);
nor U18395 (N_18395,N_12843,N_12806);
nor U18396 (N_18396,N_15389,N_14332);
nor U18397 (N_18397,N_13122,N_13764);
and U18398 (N_18398,N_14932,N_14570);
or U18399 (N_18399,N_13762,N_14741);
and U18400 (N_18400,N_13186,N_14069);
nor U18401 (N_18401,N_14362,N_12515);
nor U18402 (N_18402,N_15302,N_14579);
nor U18403 (N_18403,N_14585,N_15458);
or U18404 (N_18404,N_13550,N_13580);
or U18405 (N_18405,N_13171,N_13535);
nand U18406 (N_18406,N_15411,N_12582);
xnor U18407 (N_18407,N_13749,N_13500);
nor U18408 (N_18408,N_13957,N_14790);
or U18409 (N_18409,N_14806,N_14235);
nand U18410 (N_18410,N_13790,N_14966);
or U18411 (N_18411,N_13090,N_13028);
nand U18412 (N_18412,N_14407,N_13649);
and U18413 (N_18413,N_15489,N_12910);
nor U18414 (N_18414,N_14063,N_13089);
and U18415 (N_18415,N_12831,N_13362);
nor U18416 (N_18416,N_15062,N_14548);
nor U18417 (N_18417,N_14908,N_13335);
nand U18418 (N_18418,N_12885,N_12857);
and U18419 (N_18419,N_14726,N_14953);
or U18420 (N_18420,N_13182,N_13579);
nand U18421 (N_18421,N_15509,N_15623);
or U18422 (N_18422,N_13493,N_14144);
or U18423 (N_18423,N_13925,N_13946);
or U18424 (N_18424,N_14074,N_12891);
and U18425 (N_18425,N_12751,N_14926);
nor U18426 (N_18426,N_14334,N_13592);
or U18427 (N_18427,N_12570,N_12672);
or U18428 (N_18428,N_14624,N_14732);
nand U18429 (N_18429,N_15464,N_14648);
nor U18430 (N_18430,N_13996,N_12908);
nand U18431 (N_18431,N_13011,N_15093);
nand U18432 (N_18432,N_15408,N_14912);
xnor U18433 (N_18433,N_14714,N_12830);
nor U18434 (N_18434,N_15389,N_15232);
and U18435 (N_18435,N_12719,N_13177);
nand U18436 (N_18436,N_14427,N_14489);
and U18437 (N_18437,N_14831,N_14518);
nor U18438 (N_18438,N_15092,N_13845);
and U18439 (N_18439,N_13984,N_13668);
xor U18440 (N_18440,N_12749,N_13796);
xor U18441 (N_18441,N_13158,N_13481);
or U18442 (N_18442,N_15296,N_13742);
nor U18443 (N_18443,N_15091,N_14423);
nand U18444 (N_18444,N_14778,N_15073);
nor U18445 (N_18445,N_14700,N_14849);
nor U18446 (N_18446,N_13541,N_13119);
and U18447 (N_18447,N_14005,N_15208);
or U18448 (N_18448,N_12865,N_13389);
and U18449 (N_18449,N_14274,N_13220);
nand U18450 (N_18450,N_14640,N_12785);
nand U18451 (N_18451,N_14058,N_14926);
or U18452 (N_18452,N_13047,N_12816);
or U18453 (N_18453,N_15205,N_14051);
nor U18454 (N_18454,N_13326,N_12970);
and U18455 (N_18455,N_15288,N_13385);
xnor U18456 (N_18456,N_12750,N_15100);
and U18457 (N_18457,N_13968,N_14338);
nand U18458 (N_18458,N_14568,N_13670);
and U18459 (N_18459,N_14063,N_15559);
and U18460 (N_18460,N_12634,N_14899);
or U18461 (N_18461,N_12591,N_14523);
nand U18462 (N_18462,N_14574,N_13603);
or U18463 (N_18463,N_14033,N_12956);
xnor U18464 (N_18464,N_14117,N_14456);
nand U18465 (N_18465,N_13294,N_12786);
and U18466 (N_18466,N_14288,N_15602);
and U18467 (N_18467,N_12551,N_13123);
and U18468 (N_18468,N_14589,N_13202);
xnor U18469 (N_18469,N_14605,N_14159);
xor U18470 (N_18470,N_13703,N_13137);
xnor U18471 (N_18471,N_13689,N_13143);
nand U18472 (N_18472,N_15551,N_15319);
and U18473 (N_18473,N_13307,N_13265);
xor U18474 (N_18474,N_14867,N_14122);
and U18475 (N_18475,N_15445,N_14070);
nor U18476 (N_18476,N_13723,N_14384);
or U18477 (N_18477,N_15577,N_15069);
nor U18478 (N_18478,N_13790,N_15354);
and U18479 (N_18479,N_15214,N_14116);
nor U18480 (N_18480,N_12953,N_14295);
nor U18481 (N_18481,N_14694,N_12682);
or U18482 (N_18482,N_15569,N_14638);
or U18483 (N_18483,N_12758,N_13817);
nor U18484 (N_18484,N_13643,N_12936);
nor U18485 (N_18485,N_13215,N_12585);
and U18486 (N_18486,N_12775,N_13156);
and U18487 (N_18487,N_15313,N_12617);
and U18488 (N_18488,N_14459,N_12853);
xnor U18489 (N_18489,N_13030,N_13384);
xor U18490 (N_18490,N_12753,N_14079);
or U18491 (N_18491,N_15383,N_13568);
and U18492 (N_18492,N_15544,N_13341);
and U18493 (N_18493,N_14036,N_13387);
nand U18494 (N_18494,N_13390,N_13781);
nor U18495 (N_18495,N_13729,N_15067);
or U18496 (N_18496,N_15077,N_12965);
nor U18497 (N_18497,N_15444,N_14505);
xnor U18498 (N_18498,N_12682,N_13278);
or U18499 (N_18499,N_12688,N_12984);
xor U18500 (N_18500,N_13539,N_15375);
and U18501 (N_18501,N_13811,N_12586);
nor U18502 (N_18502,N_13274,N_14606);
or U18503 (N_18503,N_13695,N_13694);
nand U18504 (N_18504,N_13964,N_12897);
and U18505 (N_18505,N_12608,N_15183);
nor U18506 (N_18506,N_15083,N_12998);
or U18507 (N_18507,N_14621,N_14143);
and U18508 (N_18508,N_14042,N_15386);
nand U18509 (N_18509,N_13534,N_15419);
and U18510 (N_18510,N_14430,N_15493);
and U18511 (N_18511,N_13567,N_14760);
or U18512 (N_18512,N_15499,N_15457);
xnor U18513 (N_18513,N_13130,N_15575);
xor U18514 (N_18514,N_13480,N_15196);
or U18515 (N_18515,N_13804,N_13519);
or U18516 (N_18516,N_14820,N_13926);
or U18517 (N_18517,N_12564,N_14104);
or U18518 (N_18518,N_12681,N_12616);
or U18519 (N_18519,N_14945,N_14133);
nor U18520 (N_18520,N_14656,N_14119);
or U18521 (N_18521,N_12736,N_12652);
nand U18522 (N_18522,N_14070,N_13487);
and U18523 (N_18523,N_12960,N_14285);
or U18524 (N_18524,N_14068,N_12996);
or U18525 (N_18525,N_13040,N_12986);
or U18526 (N_18526,N_14992,N_14613);
nand U18527 (N_18527,N_14161,N_14228);
xnor U18528 (N_18528,N_12970,N_13241);
nand U18529 (N_18529,N_15106,N_15104);
nor U18530 (N_18530,N_14937,N_14211);
xor U18531 (N_18531,N_14829,N_13657);
or U18532 (N_18532,N_15535,N_13255);
nand U18533 (N_18533,N_13101,N_12973);
nand U18534 (N_18534,N_13996,N_14022);
and U18535 (N_18535,N_12938,N_14512);
or U18536 (N_18536,N_12674,N_15551);
or U18537 (N_18537,N_13088,N_12594);
xor U18538 (N_18538,N_13448,N_15534);
nand U18539 (N_18539,N_14306,N_13866);
and U18540 (N_18540,N_13470,N_14057);
nand U18541 (N_18541,N_14072,N_14118);
or U18542 (N_18542,N_13672,N_13120);
nor U18543 (N_18543,N_14091,N_14480);
or U18544 (N_18544,N_13472,N_14337);
nand U18545 (N_18545,N_14282,N_14880);
nor U18546 (N_18546,N_13651,N_15277);
nand U18547 (N_18547,N_15151,N_14479);
or U18548 (N_18548,N_14641,N_13344);
nand U18549 (N_18549,N_14468,N_14832);
xnor U18550 (N_18550,N_14110,N_13989);
or U18551 (N_18551,N_12647,N_13113);
xor U18552 (N_18552,N_13474,N_14179);
nand U18553 (N_18553,N_15471,N_14110);
nand U18554 (N_18554,N_13652,N_15535);
or U18555 (N_18555,N_12873,N_12678);
nor U18556 (N_18556,N_14565,N_13567);
and U18557 (N_18557,N_13796,N_14982);
nor U18558 (N_18558,N_15202,N_13634);
nand U18559 (N_18559,N_13052,N_12725);
and U18560 (N_18560,N_12829,N_12569);
or U18561 (N_18561,N_15121,N_14730);
or U18562 (N_18562,N_12732,N_12731);
nor U18563 (N_18563,N_14421,N_13490);
nor U18564 (N_18564,N_14924,N_13876);
and U18565 (N_18565,N_14003,N_14071);
nand U18566 (N_18566,N_13085,N_14381);
nor U18567 (N_18567,N_13912,N_15497);
nand U18568 (N_18568,N_13176,N_13502);
and U18569 (N_18569,N_14458,N_12940);
xnor U18570 (N_18570,N_14004,N_15457);
nor U18571 (N_18571,N_13429,N_12792);
nand U18572 (N_18572,N_14572,N_13323);
nor U18573 (N_18573,N_14690,N_14956);
nor U18574 (N_18574,N_15210,N_13665);
or U18575 (N_18575,N_12914,N_13015);
nor U18576 (N_18576,N_14343,N_14327);
nor U18577 (N_18577,N_14754,N_15519);
and U18578 (N_18578,N_13863,N_15544);
nand U18579 (N_18579,N_15465,N_12948);
nor U18580 (N_18580,N_14006,N_15340);
xor U18581 (N_18581,N_12841,N_13869);
nand U18582 (N_18582,N_13865,N_12516);
and U18583 (N_18583,N_12664,N_14502);
nand U18584 (N_18584,N_13144,N_14361);
nand U18585 (N_18585,N_13525,N_13453);
and U18586 (N_18586,N_14638,N_15416);
and U18587 (N_18587,N_13680,N_14581);
nand U18588 (N_18588,N_13985,N_12773);
and U18589 (N_18589,N_12770,N_14641);
or U18590 (N_18590,N_13478,N_14913);
and U18591 (N_18591,N_14577,N_14015);
and U18592 (N_18592,N_14060,N_13137);
nand U18593 (N_18593,N_13001,N_12620);
nor U18594 (N_18594,N_13519,N_13145);
or U18595 (N_18595,N_13883,N_13174);
or U18596 (N_18596,N_14400,N_12957);
or U18597 (N_18597,N_12738,N_14911);
nor U18598 (N_18598,N_13001,N_14722);
nand U18599 (N_18599,N_13766,N_13341);
or U18600 (N_18600,N_12719,N_13123);
nor U18601 (N_18601,N_13294,N_14484);
or U18602 (N_18602,N_14354,N_15615);
and U18603 (N_18603,N_13578,N_13900);
nand U18604 (N_18604,N_15163,N_12825);
nand U18605 (N_18605,N_14296,N_13921);
or U18606 (N_18606,N_13347,N_14808);
and U18607 (N_18607,N_13729,N_13008);
and U18608 (N_18608,N_14879,N_12996);
nor U18609 (N_18609,N_14727,N_13946);
nor U18610 (N_18610,N_14217,N_13780);
nor U18611 (N_18611,N_14194,N_13146);
and U18612 (N_18612,N_15243,N_13170);
nor U18613 (N_18613,N_15016,N_14857);
nand U18614 (N_18614,N_12820,N_12785);
and U18615 (N_18615,N_15310,N_14925);
nand U18616 (N_18616,N_12567,N_13406);
and U18617 (N_18617,N_12608,N_13329);
nor U18618 (N_18618,N_15484,N_13500);
and U18619 (N_18619,N_12899,N_13773);
nand U18620 (N_18620,N_14076,N_14559);
nor U18621 (N_18621,N_15143,N_13606);
or U18622 (N_18622,N_14060,N_14030);
xor U18623 (N_18623,N_12796,N_14863);
and U18624 (N_18624,N_13248,N_13951);
nand U18625 (N_18625,N_14064,N_14667);
nand U18626 (N_18626,N_15439,N_15068);
and U18627 (N_18627,N_15003,N_15415);
xor U18628 (N_18628,N_13380,N_13051);
nand U18629 (N_18629,N_15309,N_12617);
and U18630 (N_18630,N_13525,N_14623);
nor U18631 (N_18631,N_13178,N_13459);
xnor U18632 (N_18632,N_14526,N_14016);
nor U18633 (N_18633,N_14809,N_13259);
nand U18634 (N_18634,N_15476,N_14775);
nor U18635 (N_18635,N_13695,N_13084);
nand U18636 (N_18636,N_15450,N_13450);
and U18637 (N_18637,N_13823,N_13353);
nor U18638 (N_18638,N_15188,N_14350);
nor U18639 (N_18639,N_15151,N_14967);
or U18640 (N_18640,N_14247,N_12644);
xnor U18641 (N_18641,N_12629,N_12828);
and U18642 (N_18642,N_15562,N_14381);
nand U18643 (N_18643,N_13426,N_15015);
and U18644 (N_18644,N_12760,N_13218);
nor U18645 (N_18645,N_13181,N_13256);
nand U18646 (N_18646,N_13547,N_12648);
or U18647 (N_18647,N_12846,N_12681);
nor U18648 (N_18648,N_13620,N_15599);
nor U18649 (N_18649,N_13932,N_13302);
nor U18650 (N_18650,N_12953,N_15091);
or U18651 (N_18651,N_13486,N_14257);
or U18652 (N_18652,N_14790,N_13676);
or U18653 (N_18653,N_15330,N_13879);
or U18654 (N_18654,N_14835,N_13828);
and U18655 (N_18655,N_15068,N_14927);
xor U18656 (N_18656,N_15345,N_12737);
nor U18657 (N_18657,N_14563,N_13347);
nand U18658 (N_18658,N_13663,N_13134);
or U18659 (N_18659,N_14092,N_15007);
nor U18660 (N_18660,N_12690,N_13135);
nor U18661 (N_18661,N_13188,N_12925);
nor U18662 (N_18662,N_14137,N_12554);
nand U18663 (N_18663,N_13369,N_15334);
nor U18664 (N_18664,N_14377,N_13778);
nor U18665 (N_18665,N_13737,N_14012);
nor U18666 (N_18666,N_15563,N_14284);
and U18667 (N_18667,N_14254,N_14249);
and U18668 (N_18668,N_14860,N_13164);
and U18669 (N_18669,N_13729,N_14459);
nor U18670 (N_18670,N_13877,N_14529);
nand U18671 (N_18671,N_15179,N_15172);
and U18672 (N_18672,N_14630,N_12585);
and U18673 (N_18673,N_13768,N_14440);
or U18674 (N_18674,N_15003,N_13260);
xor U18675 (N_18675,N_13010,N_13827);
nor U18676 (N_18676,N_15458,N_12923);
nor U18677 (N_18677,N_13671,N_12956);
nor U18678 (N_18678,N_13098,N_14770);
and U18679 (N_18679,N_15172,N_13675);
nor U18680 (N_18680,N_14758,N_12849);
or U18681 (N_18681,N_14714,N_13504);
or U18682 (N_18682,N_13756,N_13267);
nand U18683 (N_18683,N_15428,N_13374);
and U18684 (N_18684,N_12750,N_13062);
nor U18685 (N_18685,N_15313,N_15236);
nor U18686 (N_18686,N_13723,N_14908);
nand U18687 (N_18687,N_14101,N_14748);
nor U18688 (N_18688,N_14645,N_14750);
nor U18689 (N_18689,N_15398,N_15291);
and U18690 (N_18690,N_13903,N_13788);
and U18691 (N_18691,N_12649,N_12648);
nor U18692 (N_18692,N_13774,N_15372);
xnor U18693 (N_18693,N_12888,N_13855);
nand U18694 (N_18694,N_12756,N_12751);
nor U18695 (N_18695,N_12522,N_15242);
and U18696 (N_18696,N_12710,N_14006);
nand U18697 (N_18697,N_15280,N_15033);
and U18698 (N_18698,N_15300,N_13924);
or U18699 (N_18699,N_14764,N_12989);
nor U18700 (N_18700,N_15081,N_15006);
xor U18701 (N_18701,N_15068,N_12607);
or U18702 (N_18702,N_15199,N_14038);
nor U18703 (N_18703,N_14487,N_15471);
or U18704 (N_18704,N_15400,N_13730);
and U18705 (N_18705,N_13677,N_14044);
nor U18706 (N_18706,N_14907,N_13224);
or U18707 (N_18707,N_13049,N_13480);
and U18708 (N_18708,N_13967,N_13514);
and U18709 (N_18709,N_15114,N_13255);
nor U18710 (N_18710,N_14042,N_14416);
or U18711 (N_18711,N_14394,N_13324);
nor U18712 (N_18712,N_13195,N_12789);
or U18713 (N_18713,N_14800,N_15046);
nor U18714 (N_18714,N_14967,N_15386);
or U18715 (N_18715,N_13294,N_13176);
and U18716 (N_18716,N_14825,N_15317);
and U18717 (N_18717,N_15084,N_13714);
or U18718 (N_18718,N_13140,N_15359);
nand U18719 (N_18719,N_13284,N_14942);
nor U18720 (N_18720,N_15453,N_13108);
or U18721 (N_18721,N_15162,N_15422);
or U18722 (N_18722,N_14635,N_15165);
and U18723 (N_18723,N_14715,N_13742);
and U18724 (N_18724,N_13514,N_14122);
nand U18725 (N_18725,N_15153,N_12675);
nand U18726 (N_18726,N_13399,N_14188);
nor U18727 (N_18727,N_13004,N_14992);
or U18728 (N_18728,N_15423,N_12685);
nor U18729 (N_18729,N_12956,N_14584);
nand U18730 (N_18730,N_14645,N_14934);
or U18731 (N_18731,N_13749,N_13930);
nand U18732 (N_18732,N_14636,N_13322);
and U18733 (N_18733,N_15198,N_15032);
and U18734 (N_18734,N_15394,N_14298);
nand U18735 (N_18735,N_15562,N_14414);
nand U18736 (N_18736,N_12514,N_13258);
and U18737 (N_18737,N_15596,N_14504);
or U18738 (N_18738,N_15014,N_14808);
and U18739 (N_18739,N_13593,N_13200);
and U18740 (N_18740,N_13597,N_14736);
xnor U18741 (N_18741,N_14362,N_12816);
and U18742 (N_18742,N_15619,N_13183);
and U18743 (N_18743,N_14930,N_15275);
nor U18744 (N_18744,N_13984,N_13174);
and U18745 (N_18745,N_14043,N_12877);
nand U18746 (N_18746,N_13650,N_14363);
or U18747 (N_18747,N_12794,N_14754);
nor U18748 (N_18748,N_13637,N_15176);
nand U18749 (N_18749,N_13531,N_13054);
or U18750 (N_18750,N_17567,N_18696);
or U18751 (N_18751,N_16413,N_18081);
nor U18752 (N_18752,N_17063,N_16597);
nor U18753 (N_18753,N_17962,N_18299);
and U18754 (N_18754,N_16675,N_18005);
and U18755 (N_18755,N_16740,N_17883);
xor U18756 (N_18756,N_16586,N_18271);
and U18757 (N_18757,N_17155,N_16877);
or U18758 (N_18758,N_16222,N_16178);
xnor U18759 (N_18759,N_16772,N_16527);
or U18760 (N_18760,N_18659,N_17290);
xnor U18761 (N_18761,N_15886,N_16872);
nor U18762 (N_18762,N_17739,N_16370);
nand U18763 (N_18763,N_18521,N_16240);
nor U18764 (N_18764,N_17929,N_16927);
xnor U18765 (N_18765,N_17553,N_16328);
xnor U18766 (N_18766,N_17702,N_17975);
or U18767 (N_18767,N_18361,N_16552);
or U18768 (N_18768,N_16581,N_18038);
and U18769 (N_18769,N_17471,N_17673);
nor U18770 (N_18770,N_18184,N_17229);
or U18771 (N_18771,N_18060,N_16901);
nor U18772 (N_18772,N_18631,N_17809);
or U18773 (N_18773,N_18747,N_17032);
or U18774 (N_18774,N_17223,N_16183);
nor U18775 (N_18775,N_15927,N_16265);
or U18776 (N_18776,N_16662,N_15943);
xnor U18777 (N_18777,N_17185,N_17922);
nor U18778 (N_18778,N_17265,N_17454);
nand U18779 (N_18779,N_15894,N_17907);
and U18780 (N_18780,N_16697,N_17841);
nand U18781 (N_18781,N_17730,N_17035);
nor U18782 (N_18782,N_17241,N_16755);
nand U18783 (N_18783,N_16315,N_18688);
nor U18784 (N_18784,N_15875,N_17786);
or U18785 (N_18785,N_17971,N_17405);
and U18786 (N_18786,N_15630,N_18019);
and U18787 (N_18787,N_18662,N_16216);
or U18788 (N_18788,N_16071,N_15936);
nor U18789 (N_18789,N_17720,N_16595);
nand U18790 (N_18790,N_18566,N_18296);
and U18791 (N_18791,N_16376,N_16890);
nor U18792 (N_18792,N_18619,N_15763);
xnor U18793 (N_18793,N_17113,N_16829);
nand U18794 (N_18794,N_17542,N_18117);
nand U18795 (N_18795,N_17287,N_15976);
nor U18796 (N_18796,N_16924,N_17592);
or U18797 (N_18797,N_16948,N_18193);
and U18798 (N_18798,N_16278,N_18043);
or U18799 (N_18799,N_17756,N_18294);
nand U18800 (N_18800,N_16615,N_17028);
nor U18801 (N_18801,N_15973,N_16333);
and U18802 (N_18802,N_15735,N_15776);
nor U18803 (N_18803,N_18606,N_16553);
xor U18804 (N_18804,N_16639,N_16307);
nand U18805 (N_18805,N_17529,N_16378);
nor U18806 (N_18806,N_18582,N_16679);
nor U18807 (N_18807,N_17343,N_18598);
and U18808 (N_18808,N_17295,N_17552);
and U18809 (N_18809,N_16821,N_17424);
or U18810 (N_18810,N_16554,N_16967);
nand U18811 (N_18811,N_16442,N_17649);
nor U18812 (N_18812,N_17861,N_15917);
nand U18813 (N_18813,N_18055,N_17516);
nand U18814 (N_18814,N_17110,N_16496);
nor U18815 (N_18815,N_16375,N_16405);
nand U18816 (N_18816,N_18245,N_16756);
nor U18817 (N_18817,N_18410,N_16400);
nand U18818 (N_18818,N_17492,N_16501);
xnor U18819 (N_18819,N_16712,N_17742);
nor U18820 (N_18820,N_18551,N_16686);
and U18821 (N_18821,N_17848,N_15777);
nand U18822 (N_18822,N_17256,N_18641);
nor U18823 (N_18823,N_18487,N_17589);
nand U18824 (N_18824,N_16176,N_16766);
and U18825 (N_18825,N_17666,N_18660);
or U18826 (N_18826,N_15792,N_17450);
nor U18827 (N_18827,N_16923,N_18592);
nand U18828 (N_18828,N_18459,N_16629);
and U18829 (N_18829,N_18113,N_17892);
nand U18830 (N_18830,N_16643,N_16680);
or U18831 (N_18831,N_17858,N_17015);
or U18832 (N_18832,N_16013,N_16251);
and U18833 (N_18833,N_18668,N_16936);
nand U18834 (N_18834,N_16480,N_17196);
or U18835 (N_18835,N_16989,N_17802);
or U18836 (N_18836,N_16583,N_16778);
and U18837 (N_18837,N_16540,N_17967);
and U18838 (N_18838,N_18085,N_17042);
and U18839 (N_18839,N_16345,N_17300);
nand U18840 (N_18840,N_16945,N_18644);
nor U18841 (N_18841,N_17996,N_16046);
or U18842 (N_18842,N_16888,N_17787);
or U18843 (N_18843,N_17116,N_15990);
nand U18844 (N_18844,N_18374,N_16215);
nand U18845 (N_18845,N_16761,N_15744);
xnor U18846 (N_18846,N_16053,N_18380);
nor U18847 (N_18847,N_18455,N_16294);
or U18848 (N_18848,N_16703,N_18241);
nor U18849 (N_18849,N_18247,N_18217);
or U18850 (N_18850,N_16912,N_17969);
and U18851 (N_18851,N_17897,N_16773);
nand U18852 (N_18852,N_16600,N_16169);
xor U18853 (N_18853,N_17213,N_17361);
nor U18854 (N_18854,N_15635,N_16846);
and U18855 (N_18855,N_17736,N_17909);
xnor U18856 (N_18856,N_16570,N_15751);
and U18857 (N_18857,N_15954,N_16207);
and U18858 (N_18858,N_17871,N_17577);
or U18859 (N_18859,N_16129,N_18121);
or U18860 (N_18860,N_17885,N_16654);
nand U18861 (N_18861,N_18625,N_16885);
and U18862 (N_18862,N_18431,N_16951);
xor U18863 (N_18863,N_18088,N_18349);
nand U18864 (N_18864,N_16117,N_16484);
or U18865 (N_18865,N_16510,N_17749);
nand U18866 (N_18866,N_16262,N_16690);
nand U18867 (N_18867,N_17152,N_16476);
and U18868 (N_18868,N_16500,N_16482);
nor U18869 (N_18869,N_17272,N_18447);
nand U18870 (N_18870,N_16202,N_17974);
xnor U18871 (N_18871,N_15821,N_17818);
nand U18872 (N_18872,N_18401,N_16632);
nor U18873 (N_18873,N_16722,N_15644);
or U18874 (N_18874,N_17778,N_18443);
and U18875 (N_18875,N_17817,N_18215);
nor U18876 (N_18876,N_17029,N_16998);
xor U18877 (N_18877,N_17192,N_17533);
nor U18878 (N_18878,N_18648,N_16796);
xnor U18879 (N_18879,N_15919,N_16096);
nor U18880 (N_18880,N_18419,N_18498);
and U18881 (N_18881,N_18421,N_17045);
and U18882 (N_18882,N_18457,N_15839);
or U18883 (N_18883,N_17723,N_17306);
nor U18884 (N_18884,N_16608,N_15931);
xnor U18885 (N_18885,N_16340,N_16964);
nor U18886 (N_18886,N_17455,N_15683);
and U18887 (N_18887,N_16079,N_15942);
or U18888 (N_18888,N_18229,N_17374);
or U18889 (N_18889,N_17635,N_18056);
or U18890 (N_18890,N_16903,N_15680);
and U18891 (N_18891,N_15668,N_17249);
nor U18892 (N_18892,N_15674,N_17622);
and U18893 (N_18893,N_16897,N_18182);
nand U18894 (N_18894,N_18293,N_17629);
and U18895 (N_18895,N_18646,N_16957);
and U18896 (N_18896,N_18404,N_18111);
nand U18897 (N_18897,N_18168,N_15705);
nor U18898 (N_18898,N_16134,N_15952);
xnor U18899 (N_18899,N_18645,N_16716);
xor U18900 (N_18900,N_17278,N_17129);
and U18901 (N_18901,N_15824,N_16723);
or U18902 (N_18902,N_17834,N_18096);
and U18903 (N_18903,N_16017,N_18173);
nand U18904 (N_18904,N_16719,N_17475);
or U18905 (N_18905,N_16663,N_16781);
or U18906 (N_18906,N_15808,N_16933);
nand U18907 (N_18907,N_15650,N_17681);
or U18908 (N_18908,N_17371,N_18212);
nor U18909 (N_18909,N_17557,N_16729);
and U18910 (N_18910,N_16735,N_18517);
nand U18911 (N_18911,N_17208,N_18428);
or U18912 (N_18912,N_16757,N_18283);
and U18913 (N_18913,N_17257,N_17463);
nor U18914 (N_18914,N_18266,N_16750);
or U18915 (N_18915,N_16953,N_16992);
xor U18916 (N_18916,N_17359,N_17839);
and U18917 (N_18917,N_17347,N_18065);
nor U18918 (N_18918,N_16545,N_16397);
and U18919 (N_18919,N_16324,N_16028);
xor U18920 (N_18920,N_17457,N_16010);
nor U18921 (N_18921,N_18208,N_17698);
nor U18922 (N_18922,N_17865,N_16800);
or U18923 (N_18923,N_16115,N_17587);
and U18924 (N_18924,N_16530,N_17062);
and U18925 (N_18925,N_16943,N_16720);
nor U18926 (N_18926,N_16235,N_16652);
or U18927 (N_18927,N_16423,N_16677);
nor U18928 (N_18928,N_17419,N_18058);
nand U18929 (N_18929,N_15834,N_16864);
nor U18930 (N_18930,N_18183,N_17065);
nand U18931 (N_18931,N_17198,N_17182);
or U18932 (N_18932,N_16995,N_16233);
nand U18933 (N_18933,N_17100,N_17608);
xnor U18934 (N_18934,N_18196,N_16748);
nand U18935 (N_18935,N_18093,N_16733);
nand U18936 (N_18936,N_18339,N_16777);
and U18937 (N_18937,N_17214,N_15823);
or U18938 (N_18938,N_18122,N_15830);
xor U18939 (N_18939,N_17276,N_17773);
or U18940 (N_18940,N_18226,N_17019);
and U18941 (N_18941,N_18204,N_17867);
and U18942 (N_18942,N_17187,N_17905);
or U18943 (N_18943,N_16598,N_16627);
nor U18944 (N_18944,N_18714,N_17031);
nor U18945 (N_18945,N_18249,N_16186);
and U18946 (N_18946,N_16401,N_16179);
and U18947 (N_18947,N_17977,N_15941);
nand U18948 (N_18948,N_18475,N_16021);
or U18949 (N_18949,N_18147,N_17618);
nand U18950 (N_18950,N_16494,N_16838);
and U18951 (N_18951,N_17149,N_18332);
xnor U18952 (N_18952,N_17641,N_16153);
nand U18953 (N_18953,N_17066,N_16975);
or U18954 (N_18954,N_17163,N_17121);
or U18955 (N_18955,N_17003,N_17012);
nand U18956 (N_18956,N_16695,N_16956);
or U18957 (N_18957,N_16263,N_16163);
or U18958 (N_18958,N_16779,N_15714);
and U18959 (N_18959,N_16108,N_17925);
xnor U18960 (N_18960,N_15779,N_16699);
or U18961 (N_18961,N_16428,N_17453);
or U18962 (N_18962,N_17950,N_18153);
and U18963 (N_18963,N_16768,N_16715);
or U18964 (N_18964,N_17141,N_15998);
nor U18965 (N_18965,N_17391,N_16710);
nand U18966 (N_18966,N_16726,N_18490);
or U18967 (N_18967,N_15836,N_17126);
nand U18968 (N_18968,N_17780,N_16567);
and U18969 (N_18969,N_18615,N_17389);
and U18970 (N_18970,N_15944,N_18013);
or U18971 (N_18971,N_16083,N_16850);
xor U18972 (N_18972,N_17965,N_16357);
and U18973 (N_18973,N_17538,N_16062);
or U18974 (N_18974,N_16637,N_17186);
and U18975 (N_18975,N_18531,N_18057);
nor U18976 (N_18976,N_18405,N_16802);
and U18977 (N_18977,N_16217,N_15694);
nor U18978 (N_18978,N_18156,N_16048);
xnor U18979 (N_18979,N_16958,N_16390);
or U18980 (N_18980,N_18684,N_17690);
nor U18981 (N_18981,N_16837,N_18160);
and U18982 (N_18982,N_17331,N_15962);
or U18983 (N_18983,N_15711,N_17006);
or U18984 (N_18984,N_16836,N_17903);
xor U18985 (N_18985,N_18608,N_17423);
nor U18986 (N_18986,N_18398,N_18133);
xnor U18987 (N_18987,N_15670,N_16711);
or U18988 (N_18988,N_16651,N_18656);
nand U18989 (N_18989,N_17373,N_18244);
or U18990 (N_18990,N_15872,N_18118);
and U18991 (N_18991,N_15840,N_17494);
nand U18992 (N_18992,N_16991,N_18012);
or U18993 (N_18993,N_16783,N_17550);
xor U18994 (N_18994,N_16269,N_17421);
nor U18995 (N_18995,N_16514,N_15930);
or U18996 (N_18996,N_18280,N_16288);
or U18997 (N_18997,N_18188,N_17283);
xor U18998 (N_18998,N_16594,N_16636);
nor U18999 (N_18999,N_17437,N_16069);
xor U19000 (N_19000,N_16974,N_18399);
and U19001 (N_19001,N_18738,N_16646);
and U19002 (N_19002,N_18409,N_15866);
or U19003 (N_19003,N_16489,N_16274);
xor U19004 (N_19004,N_17224,N_18169);
nor U19005 (N_19005,N_17325,N_17175);
or U19006 (N_19006,N_17826,N_16782);
or U19007 (N_19007,N_18746,N_15924);
xor U19008 (N_19008,N_15911,N_16882);
nand U19009 (N_19009,N_18526,N_15978);
nor U19010 (N_19010,N_16407,N_17327);
and U19011 (N_19011,N_17877,N_17601);
nand U19012 (N_19012,N_16420,N_18698);
nand U19013 (N_19013,N_17458,N_17460);
nand U19014 (N_19014,N_17707,N_16954);
nor U19015 (N_19015,N_16347,N_17324);
or U19016 (N_19016,N_18116,N_16742);
nor U19017 (N_19017,N_15929,N_18562);
nor U19018 (N_19018,N_18357,N_16101);
or U19019 (N_19019,N_16082,N_16208);
nor U19020 (N_19020,N_17642,N_18181);
xnor U19021 (N_19021,N_16075,N_17715);
xnor U19022 (N_19022,N_17105,N_18171);
or U19023 (N_19023,N_17530,N_17918);
nor U19024 (N_19024,N_17025,N_15890);
nor U19025 (N_19025,N_16090,N_16085);
xor U19026 (N_19026,N_17879,N_15775);
xor U19027 (N_19027,N_17174,N_16606);
or U19028 (N_19028,N_17418,N_18446);
and U19029 (N_19029,N_15665,N_15740);
or U19030 (N_19030,N_15722,N_16425);
or U19031 (N_19031,N_16283,N_16112);
or U19032 (N_19032,N_18326,N_17908);
xor U19033 (N_19033,N_16242,N_15961);
or U19034 (N_19034,N_16213,N_18092);
nor U19035 (N_19035,N_16743,N_15685);
nand U19036 (N_19036,N_17939,N_17049);
nand U19037 (N_19037,N_17766,N_15967);
nor U19038 (N_19038,N_16884,N_16529);
nor U19039 (N_19039,N_16116,N_17785);
nor U19040 (N_19040,N_18577,N_18624);
nor U19041 (N_19041,N_15850,N_17348);
nand U19042 (N_19042,N_16511,N_17020);
nand U19043 (N_19043,N_17754,N_15785);
nand U19044 (N_19044,N_16870,N_16320);
nor U19045 (N_19045,N_16009,N_16547);
and U19046 (N_19046,N_18234,N_16642);
and U19047 (N_19047,N_18439,N_18219);
or U19048 (N_19048,N_18462,N_15937);
nor U19049 (N_19049,N_16827,N_17267);
or U19050 (N_19050,N_18739,N_17801);
nand U19051 (N_19051,N_15778,N_16573);
or U19052 (N_19052,N_16067,N_15757);
nand U19053 (N_19053,N_15667,N_16738);
xor U19054 (N_19054,N_17899,N_16737);
and U19055 (N_19055,N_17136,N_16461);
xor U19056 (N_19056,N_16970,N_17251);
nand U19057 (N_19057,N_18259,N_16005);
nand U19058 (N_19058,N_18106,N_17752);
and U19059 (N_19059,N_18564,N_18048);
xor U19060 (N_19060,N_17815,N_15902);
nor U19061 (N_19061,N_17258,N_16914);
nor U19062 (N_19062,N_18119,N_18590);
xor U19063 (N_19063,N_16487,N_15994);
nand U19064 (N_19064,N_15642,N_16807);
and U19065 (N_19065,N_16184,N_17445);
or U19066 (N_19066,N_15666,N_17190);
nand U19067 (N_19067,N_16209,N_18677);
nand U19068 (N_19068,N_15817,N_17882);
nor U19069 (N_19069,N_18716,N_15730);
nor U19070 (N_19070,N_18499,N_16605);
and U19071 (N_19071,N_18485,N_17222);
xnor U19072 (N_19072,N_17036,N_18286);
nand U19073 (N_19073,N_16894,N_15687);
nor U19074 (N_19074,N_16714,N_18214);
nor U19075 (N_19075,N_16666,N_16620);
nor U19076 (N_19076,N_18298,N_16377);
nor U19077 (N_19077,N_16744,N_16539);
or U19078 (N_19078,N_16011,N_17171);
or U19079 (N_19079,N_18630,N_16765);
nor U19080 (N_19080,N_17878,N_18432);
or U19081 (N_19081,N_16847,N_17963);
and U19082 (N_19082,N_16147,N_18220);
nor U19083 (N_19083,N_17159,N_17221);
nand U19084 (N_19084,N_17440,N_15862);
xnor U19085 (N_19085,N_17763,N_17140);
nand U19086 (N_19086,N_17153,N_17615);
or U19087 (N_19087,N_16492,N_15764);
nor U19088 (N_19088,N_18632,N_16180);
xnor U19089 (N_19089,N_18484,N_18612);
nand U19090 (N_19090,N_15804,N_17442);
nand U19091 (N_19091,N_15765,N_17411);
and U19092 (N_19092,N_16667,N_18479);
or U19093 (N_19093,N_16386,N_16792);
or U19094 (N_19094,N_16336,N_16329);
or U19095 (N_19095,N_16785,N_18300);
nor U19096 (N_19096,N_18640,N_16981);
or U19097 (N_19097,N_17392,N_18359);
nor U19098 (N_19098,N_16795,N_17366);
nor U19099 (N_19099,N_17312,N_18743);
xnor U19100 (N_19100,N_17724,N_16591);
or U19101 (N_19101,N_16220,N_17227);
and U19102 (N_19102,N_18110,N_18549);
or U19103 (N_19103,N_17812,N_17584);
and U19104 (N_19104,N_16059,N_16578);
and U19105 (N_19105,N_18642,N_17694);
nand U19106 (N_19106,N_18705,N_15684);
and U19107 (N_19107,N_16246,N_17580);
nor U19108 (N_19108,N_17469,N_17339);
nand U19109 (N_19109,N_16488,N_18651);
or U19110 (N_19110,N_17906,N_17228);
and U19111 (N_19111,N_17124,N_17912);
and U19112 (N_19112,N_17740,N_17402);
xnor U19113 (N_19113,N_18017,N_18018);
and U19114 (N_19114,N_16419,N_16195);
and U19115 (N_19115,N_17631,N_18541);
nor U19116 (N_19116,N_16844,N_15798);
xor U19117 (N_19117,N_17093,N_16084);
xnor U19118 (N_19118,N_18670,N_16883);
and U19119 (N_19119,N_16143,N_18552);
and U19120 (N_19120,N_16960,N_17144);
nand U19121 (N_19121,N_17731,N_16287);
nor U19122 (N_19122,N_17551,N_17351);
nor U19123 (N_19123,N_15796,N_17689);
nand U19124 (N_19124,N_17001,N_16164);
nor U19125 (N_19125,N_17941,N_16342);
xor U19126 (N_19126,N_18550,N_17531);
or U19127 (N_19127,N_16416,N_16618);
nand U19128 (N_19128,N_15797,N_17555);
nand U19129 (N_19129,N_17661,N_17047);
nand U19130 (N_19130,N_16045,N_17429);
and U19131 (N_19131,N_16668,N_18345);
nand U19132 (N_19132,N_18701,N_18515);
nor U19133 (N_19133,N_16299,N_18712);
and U19134 (N_19134,N_18741,N_17526);
and U19135 (N_19135,N_17528,N_16490);
nand U19136 (N_19136,N_17291,N_16909);
nand U19137 (N_19137,N_18444,N_18284);
xor U19138 (N_19138,N_18663,N_16843);
or U19139 (N_19139,N_17337,N_18540);
or U19140 (N_19140,N_17827,N_16403);
nand U19141 (N_19141,N_16919,N_17039);
nand U19142 (N_19142,N_16346,N_18364);
nor U19143 (N_19143,N_18344,N_17293);
nand U19144 (N_19144,N_17461,N_17565);
or U19145 (N_19145,N_16359,N_16170);
nor U19146 (N_19146,N_17692,N_17304);
and U19147 (N_19147,N_17911,N_16963);
nor U19148 (N_19148,N_18383,N_16366);
nand U19149 (N_19149,N_17973,N_18723);
and U19150 (N_19150,N_17808,N_17628);
or U19151 (N_19151,N_17670,N_16685);
or U19152 (N_19152,N_18228,N_16167);
or U19153 (N_19153,N_16794,N_17816);
nor U19154 (N_19154,N_17598,N_17083);
and U19155 (N_19155,N_18596,N_16495);
nand U19156 (N_19156,N_15896,N_18072);
or U19157 (N_19157,N_16504,N_15716);
nand U19158 (N_19158,N_17957,N_18597);
nor U19159 (N_19159,N_16383,N_18492);
nor U19160 (N_19160,N_17997,N_18500);
nor U19161 (N_19161,N_18554,N_17660);
and U19162 (N_19162,N_15958,N_16879);
and U19163 (N_19163,N_18151,N_17081);
and U19164 (N_19164,N_17506,N_18657);
and U19165 (N_19165,N_17880,N_16809);
xnor U19166 (N_19166,N_16952,N_17646);
or U19167 (N_19167,N_18497,N_16638);
nand U19168 (N_19168,N_17958,N_15801);
or U19169 (N_19169,N_18607,N_18558);
nand U19170 (N_19170,N_16984,N_16946);
nor U19171 (N_19171,N_18354,N_16189);
nand U19172 (N_19172,N_18438,N_18338);
xor U19173 (N_19173,N_18585,N_16369);
or U19174 (N_19174,N_15632,N_18278);
or U19175 (N_19175,N_17633,N_16937);
nor U19176 (N_19176,N_18045,N_18050);
or U19177 (N_19177,N_16702,N_17088);
nand U19178 (N_19178,N_16237,N_18033);
xnor U19179 (N_19179,N_17474,N_17215);
nand U19180 (N_19180,N_18675,N_18346);
and U19181 (N_19181,N_16503,N_16822);
nand U19182 (N_19182,N_16041,N_17459);
nor U19183 (N_19183,N_17444,N_16231);
or U19184 (N_19184,N_16650,N_18481);
nor U19185 (N_19185,N_16736,N_17274);
or U19186 (N_19186,N_17737,N_18527);
and U19187 (N_19187,N_17746,N_17379);
or U19188 (N_19188,N_17363,N_17591);
nand U19189 (N_19189,N_15864,N_18406);
and U19190 (N_19190,N_18655,N_18152);
xor U19191 (N_19191,N_18063,N_16568);
nor U19192 (N_19192,N_17390,N_18709);
nand U19193 (N_19193,N_16621,N_17656);
nor U19194 (N_19194,N_17842,N_18689);
or U19195 (N_19195,N_18664,N_17404);
nand U19196 (N_19196,N_17245,N_16042);
nor U19197 (N_19197,N_16604,N_17791);
and U19198 (N_19198,N_16095,N_17686);
and U19199 (N_19199,N_16281,N_16705);
and U19200 (N_19200,N_18253,N_17853);
nand U19201 (N_19201,N_16248,N_17886);
or U19202 (N_19202,N_16860,N_16614);
and U19203 (N_19203,N_15956,N_17433);
nor U19204 (N_19204,N_18303,N_17711);
or U19205 (N_19205,N_17978,N_17090);
xor U19206 (N_19206,N_15838,N_16562);
and U19207 (N_19207,N_16483,N_18729);
nor U19208 (N_19208,N_17024,N_15820);
nor U19209 (N_19209,N_16931,N_18732);
nand U19210 (N_19210,N_16453,N_15795);
nor U19211 (N_19211,N_18674,N_17569);
nor U19212 (N_19212,N_18192,N_17983);
and U19213 (N_19213,N_18437,N_16791);
nand U19214 (N_19214,N_16731,N_16920);
or U19215 (N_19215,N_18185,N_16891);
or U19216 (N_19216,N_15837,N_18142);
and U19217 (N_19217,N_18581,N_16302);
and U19218 (N_19218,N_16300,N_16424);
nor U19219 (N_19219,N_15753,N_15657);
xnor U19220 (N_19220,N_18433,N_16541);
nor U19221 (N_19221,N_15932,N_15945);
or U19222 (N_19222,N_16823,N_16961);
nand U19223 (N_19223,N_16688,N_18242);
or U19224 (N_19224,N_18158,N_16505);
or U19225 (N_19225,N_17843,N_17913);
nand U19226 (N_19226,N_18264,N_15701);
nor U19227 (N_19227,N_17115,N_17497);
nor U19228 (N_19228,N_17543,N_16040);
nand U19229 (N_19229,N_16855,N_18250);
and U19230 (N_19230,N_18604,N_18744);
nand U19231 (N_19231,N_16976,N_18010);
nor U19232 (N_19232,N_15641,N_15899);
xor U19233 (N_19233,N_16074,N_17416);
nor U19234 (N_19234,N_18635,N_16718);
nor U19235 (N_19235,N_16799,N_17340);
or U19236 (N_19236,N_17762,N_18166);
or U19237 (N_19237,N_18416,N_15964);
and U19238 (N_19238,N_16312,N_17181);
and U19239 (N_19239,N_16118,N_17179);
xnor U19240 (N_19240,N_18112,N_15809);
and U19241 (N_19241,N_18610,N_17091);
and U19242 (N_19242,N_16691,N_17652);
nor U19243 (N_19243,N_15949,N_18561);
or U19244 (N_19244,N_16361,N_17679);
nand U19245 (N_19245,N_16103,N_17466);
or U19246 (N_19246,N_16286,N_17859);
or U19247 (N_19247,N_17800,N_18268);
nand U19248 (N_19248,N_17733,N_16780);
nand U19249 (N_19249,N_15845,N_17296);
nor U19250 (N_19250,N_17319,N_18034);
xnor U19251 (N_19251,N_15905,N_17362);
and U19252 (N_19252,N_18529,N_16468);
nand U19253 (N_19253,N_17368,N_18465);
xnor U19254 (N_19254,N_17507,N_18222);
or U19255 (N_19255,N_15689,N_17145);
nand U19256 (N_19256,N_18695,N_17397);
and U19257 (N_19257,N_16798,N_18016);
nand U19258 (N_19258,N_18545,N_16617);
nor U19259 (N_19259,N_17896,N_17606);
nand U19260 (N_19260,N_16457,N_15934);
nor U19261 (N_19261,N_16298,N_15636);
nor U19262 (N_19262,N_15869,N_17700);
or U19263 (N_19263,N_16168,N_17639);
or U19264 (N_19264,N_17204,N_16574);
nand U19265 (N_19265,N_18452,N_18177);
nand U19266 (N_19266,N_17683,N_18456);
or U19267 (N_19267,N_18422,N_15859);
and U19268 (N_19268,N_17477,N_16521);
and U19269 (N_19269,N_16899,N_16411);
and U19270 (N_19270,N_17054,N_16588);
and U19271 (N_19271,N_18084,N_15749);
nor U19272 (N_19272,N_16587,N_16259);
or U19273 (N_19273,N_18369,N_16693);
and U19274 (N_19274,N_16137,N_16049);
or U19275 (N_19275,N_17448,N_15984);
nand U19276 (N_19276,N_18146,N_17813);
nand U19277 (N_19277,N_16204,N_16830);
and U19278 (N_19278,N_18504,N_16990);
nand U19279 (N_19279,N_18333,N_17112);
or U19280 (N_19280,N_16034,N_18031);
and U19281 (N_19281,N_18302,N_16551);
nand U19282 (N_19282,N_16520,N_17594);
nor U19283 (N_19283,N_17209,N_18588);
and U19284 (N_19284,N_18737,N_16839);
and U19285 (N_19285,N_17383,N_16518);
nand U19286 (N_19286,N_18322,N_17761);
or U19287 (N_19287,N_16273,N_17676);
nor U19288 (N_19288,N_17989,N_17075);
xor U19289 (N_19289,N_18408,N_17824);
or U19290 (N_19290,N_16701,N_18251);
or U19291 (N_19291,N_15649,N_18109);
and U19292 (N_19292,N_16589,N_15710);
nor U19293 (N_19293,N_17647,N_15881);
xor U19294 (N_19294,N_16060,N_15769);
nand U19295 (N_19295,N_18190,N_17888);
nand U19296 (N_19296,N_18477,N_17585);
xnor U19297 (N_19297,N_15912,N_17757);
or U19298 (N_19298,N_18073,N_15690);
or U19299 (N_19299,N_17684,N_18565);
or U19300 (N_19300,N_18254,N_18337);
or U19301 (N_19301,N_16309,N_16064);
or U19302 (N_19302,N_16415,N_16754);
nor U19303 (N_19303,N_16861,N_17520);
or U19304 (N_19304,N_16725,N_18652);
or U19305 (N_19305,N_17206,N_18070);
nor U19306 (N_19306,N_15766,N_16126);
nor U19307 (N_19307,N_16121,N_17210);
nand U19308 (N_19308,N_15829,N_16003);
nor U19309 (N_19309,N_18699,N_16325);
or U19310 (N_19310,N_16674,N_17898);
or U19311 (N_19311,N_16683,N_15789);
nand U19312 (N_19312,N_16524,N_16241);
or U19313 (N_19313,N_17875,N_16775);
and U19314 (N_19314,N_17940,N_16198);
and U19315 (N_19315,N_17219,N_17829);
nor U19316 (N_19316,N_16834,N_16556);
nand U19317 (N_19317,N_18292,N_16261);
nor U19318 (N_19318,N_18257,N_17151);
and U19319 (N_19319,N_16497,N_15831);
and U19320 (N_19320,N_17486,N_18211);
and U19321 (N_19321,N_16797,N_16368);
or U19322 (N_19322,N_16645,N_16825);
nand U19323 (N_19323,N_18131,N_16181);
or U19324 (N_19324,N_16293,N_17435);
nand U19325 (N_19325,N_16499,N_16350);
xnor U19326 (N_19326,N_18352,N_17310);
and U19327 (N_19327,N_18685,N_18555);
and U19328 (N_19328,N_16840,N_18533);
or U19329 (N_19329,N_17847,N_16687);
and U19330 (N_19330,N_17352,N_16099);
or U19331 (N_19331,N_16561,N_17795);
and U19332 (N_19332,N_16141,N_16292);
nand U19333 (N_19333,N_15860,N_18167);
and U19334 (N_19334,N_16999,N_18542);
xor U19335 (N_19335,N_16230,N_15957);
and U19336 (N_19336,N_17765,N_16349);
xnor U19337 (N_19337,N_18463,N_17890);
or U19338 (N_19338,N_17515,N_16290);
or U19339 (N_19339,N_17148,N_18671);
xor U19340 (N_19340,N_15733,N_16506);
and U19341 (N_19341,N_17142,N_17009);
nor U19342 (N_19342,N_18071,N_17665);
or U19343 (N_19343,N_16728,N_17350);
xor U19344 (N_19344,N_18000,N_18510);
nor U19345 (N_19345,N_18579,N_17203);
or U19346 (N_19346,N_16033,N_16555);
and U19347 (N_19347,N_18378,N_17653);
xor U19348 (N_19348,N_18586,N_17894);
nor U19349 (N_19349,N_16344,N_16258);
xor U19350 (N_19350,N_17840,N_16311);
nand U19351 (N_19351,N_18495,N_17558);
nor U19352 (N_19352,N_16223,N_17825);
nor U19353 (N_19353,N_16076,N_16944);
nor U19354 (N_19354,N_15723,N_17511);
xor U19355 (N_19355,N_17328,N_18233);
xnor U19356 (N_19356,N_16867,N_18130);
or U19357 (N_19357,N_18295,N_18366);
nor U19358 (N_19358,N_18077,N_17805);
and U19359 (N_19359,N_15652,N_15848);
nand U19360 (N_19360,N_15719,N_15737);
nor U19361 (N_19361,N_17468,N_16966);
or U19362 (N_19362,N_17819,N_16874);
nor U19363 (N_19363,N_16707,N_17648);
xnor U19364 (N_19364,N_17164,N_17333);
xnor U19365 (N_19365,N_15960,N_17775);
and U19366 (N_19366,N_16372,N_17092);
or U19367 (N_19367,N_17902,N_17759);
or U19368 (N_19368,N_16455,N_18318);
nand U19369 (N_19369,N_18323,N_15691);
and U19370 (N_19370,N_16157,N_16832);
and U19371 (N_19371,N_15747,N_17864);
and U19372 (N_19372,N_17147,N_16565);
or U19373 (N_19373,N_17946,N_17326);
and U19374 (N_19374,N_18740,N_17169);
or U19375 (N_19375,N_17118,N_18681);
or U19376 (N_19376,N_18103,N_17893);
and U19377 (N_19377,N_15708,N_17082);
or U19378 (N_19378,N_15783,N_16599);
or U19379 (N_19379,N_17863,N_16323);
nor U19380 (N_19380,N_18461,N_17370);
and U19381 (N_19381,N_17508,N_15946);
or U19382 (N_19382,N_16577,N_18007);
nor U19383 (N_19383,N_17990,N_18661);
or U19384 (N_19384,N_16509,N_16584);
nor U19385 (N_19385,N_16002,N_17201);
or U19386 (N_19386,N_15773,N_17930);
or U19387 (N_19387,N_16027,N_16704);
and U19388 (N_19388,N_16805,N_18330);
nand U19389 (N_19389,N_18700,N_18514);
nand U19390 (N_19390,N_17959,N_16379);
nand U19391 (N_19391,N_16569,N_18516);
or U19392 (N_19392,N_17311,N_18291);
or U19393 (N_19393,N_18390,N_16332);
nor U19394 (N_19394,N_17104,N_16634);
nor U19395 (N_19395,N_16104,N_16841);
or U19396 (N_19396,N_15715,N_17595);
nand U19397 (N_19397,N_17561,N_16459);
or U19398 (N_19398,N_17275,N_18136);
or U19399 (N_19399,N_18617,N_17173);
and U19400 (N_19400,N_15793,N_16955);
or U19401 (N_19401,N_15791,N_16160);
and U19402 (N_19402,N_18002,N_17470);
nand U19403 (N_19403,N_18003,N_17891);
and U19404 (N_19404,N_15842,N_18102);
xnor U19405 (N_19405,N_17532,N_16052);
nand U19406 (N_19406,N_16513,N_17156);
nor U19407 (N_19407,N_15841,N_16938);
nor U19408 (N_19408,N_18221,N_18287);
or U19409 (N_19409,N_17114,N_16385);
and U19410 (N_19410,N_17014,N_15992);
nor U19411 (N_19411,N_16365,N_17430);
or U19412 (N_19412,N_18537,N_18239);
nand U19413 (N_19413,N_16982,N_16203);
nand U19414 (N_19414,N_18161,N_17524);
nor U19415 (N_19415,N_16026,N_17992);
and U19416 (N_19416,N_16648,N_18319);
nor U19417 (N_19417,N_15822,N_15787);
nand U19418 (N_19418,N_18097,N_17487);
and U19419 (N_19419,N_15922,N_16566);
nor U19420 (N_19420,N_17788,N_17048);
and U19421 (N_19421,N_15947,N_17837);
or U19422 (N_19422,N_17714,N_18039);
nor U19423 (N_19423,N_16575,N_15865);
or U19424 (N_19424,N_17651,N_15675);
nor U19425 (N_19425,N_16282,N_16458);
nor U19426 (N_19426,N_18591,N_15732);
nor U19427 (N_19427,N_18186,N_16174);
nor U19428 (N_19428,N_18394,N_18573);
or U19429 (N_19429,N_18464,N_17087);
xor U19430 (N_19430,N_18114,N_15826);
nor U19431 (N_19431,N_17360,N_17674);
nor U19432 (N_19432,N_16123,N_17189);
and U19433 (N_19433,N_15965,N_17495);
and U19434 (N_19434,N_17499,N_17491);
nor U19435 (N_19435,N_17887,N_15634);
and U19436 (N_19436,N_18379,N_16111);
nand U19437 (N_19437,N_17058,N_16512);
and U19438 (N_19438,N_16381,N_16152);
or U19439 (N_19439,N_17915,N_17687);
and U19440 (N_19440,N_17857,N_16314);
or U19441 (N_19441,N_18343,N_16388);
nand U19442 (N_19442,N_16437,N_18209);
nand U19443 (N_19443,N_18667,N_17137);
nor U19444 (N_19444,N_15745,N_16250);
nand U19445 (N_19445,N_17735,N_17517);
nand U19446 (N_19446,N_15963,N_17232);
or U19447 (N_19447,N_17792,N_18638);
nand U19448 (N_19448,N_16558,N_15853);
nand U19449 (N_19449,N_16393,N_16660);
nand U19450 (N_19450,N_15968,N_18707);
xnor U19451 (N_19451,N_17900,N_17191);
nor U19452 (N_19452,N_16801,N_18710);
nor U19453 (N_19453,N_17016,N_17784);
nand U19454 (N_19454,N_17280,N_16192);
or U19455 (N_19455,N_17582,N_16741);
nand U19456 (N_19456,N_18312,N_18351);
nor U19457 (N_19457,N_16072,N_18089);
or U19458 (N_19458,N_18680,N_16602);
and U19459 (N_19459,N_17623,N_17771);
xor U19460 (N_19460,N_18069,N_17895);
nor U19461 (N_19461,N_17713,N_15806);
nand U19462 (N_19462,N_18365,N_15923);
nand U19463 (N_19463,N_18702,N_18309);
and U19464 (N_19464,N_18083,N_17180);
and U19465 (N_19465,N_17158,N_17247);
nor U19466 (N_19466,N_16470,N_17500);
nand U19467 (N_19467,N_15981,N_16454);
nand U19468 (N_19468,N_16337,N_18001);
and U19469 (N_19469,N_16252,N_16194);
or U19470 (N_19470,N_17041,N_16672);
nor U19471 (N_19471,N_18372,N_17252);
and U19472 (N_19472,N_16239,N_16172);
nor U19473 (N_19473,N_17831,N_15996);
and U19474 (N_19474,N_18467,N_16018);
nor U19475 (N_19475,N_18155,N_16343);
or U19476 (N_19476,N_15699,N_18159);
and U19477 (N_19477,N_16776,N_16464);
nor U19478 (N_19478,N_16363,N_16811);
and U19479 (N_19479,N_16331,N_15656);
or U19480 (N_19480,N_17807,N_17125);
nor U19481 (N_19481,N_17536,N_18602);
or U19482 (N_19482,N_18195,N_17309);
nand U19483 (N_19483,N_17426,N_17462);
or U19484 (N_19484,N_16439,N_17335);
nor U19485 (N_19485,N_17018,N_17143);
or U19486 (N_19486,N_18024,N_16427);
nor U19487 (N_19487,N_18094,N_16149);
and U19488 (N_19488,N_15868,N_16644);
and U19489 (N_19489,N_16056,N_17298);
or U19490 (N_19490,N_16972,N_16968);
or U19491 (N_19491,N_18037,N_16313);
nor U19492 (N_19492,N_15920,N_16146);
nand U19493 (N_19493,N_17678,N_17951);
or U19494 (N_19494,N_17849,N_18041);
and U19495 (N_19495,N_15660,N_18686);
and U19496 (N_19496,N_16817,N_15857);
nor U19497 (N_19497,N_16444,N_18711);
nor U19498 (N_19498,N_18697,N_16950);
nor U19499 (N_19499,N_15855,N_17501);
nand U19500 (N_19500,N_16043,N_16658);
and U19501 (N_19501,N_16234,N_18199);
nor U19502 (N_19502,N_18468,N_17621);
and U19503 (N_19503,N_17030,N_17718);
and U19504 (N_19504,N_17743,N_18132);
and U19505 (N_19505,N_17693,N_16889);
or U19506 (N_19506,N_17413,N_16866);
nor U19507 (N_19507,N_16949,N_18613);
nand U19508 (N_19508,N_16306,N_17414);
or U19509 (N_19509,N_18583,N_18206);
or U19510 (N_19510,N_18628,N_16631);
nand U19511 (N_19511,N_18095,N_16394);
and U19512 (N_19512,N_15731,N_17830);
and U19513 (N_19513,N_17243,N_17961);
xnor U19514 (N_19514,N_15828,N_18595);
nand U19515 (N_19515,N_17472,N_16364);
or U19516 (N_19516,N_15677,N_18538);
or U19517 (N_19517,N_17921,N_17449);
nor U19518 (N_19518,N_17485,N_17138);
nand U19519 (N_19519,N_17277,N_16360);
nand U19520 (N_19520,N_17986,N_15771);
or U19521 (N_19521,N_16138,N_18609);
nand U19522 (N_19522,N_17993,N_17954);
or U19523 (N_19523,N_18724,N_18415);
nor U19524 (N_19524,N_15908,N_18066);
nor U19525 (N_19525,N_16856,N_18216);
or U19526 (N_19526,N_17095,N_18311);
or U19527 (N_19527,N_15925,N_16997);
and U19528 (N_19528,N_16175,N_17271);
nor U19529 (N_19529,N_16133,N_18727);
nor U19530 (N_19530,N_16014,N_17607);
or U19531 (N_19531,N_17626,N_16876);
and U19532 (N_19532,N_17870,N_18205);
nor U19533 (N_19533,N_17297,N_17211);
and U19534 (N_19534,N_18075,N_15767);
nand U19535 (N_19535,N_17866,N_16450);
and U19536 (N_19536,N_17644,N_17872);
or U19537 (N_19537,N_18474,N_18708);
and U19538 (N_19538,N_16166,N_15672);
and U19539 (N_19539,N_15734,N_16669);
or U19540 (N_19540,N_16276,N_17747);
or U19541 (N_19541,N_16462,N_16947);
nand U19542 (N_19542,N_16774,N_15646);
and U19543 (N_19543,N_18600,N_17320);
or U19544 (N_19544,N_17488,N_16443);
nand U19545 (N_19545,N_16810,N_17685);
and U19546 (N_19546,N_18601,N_16087);
xor U19547 (N_19547,N_17655,N_18356);
xor U19548 (N_19548,N_16245,N_16015);
and U19549 (N_19549,N_16929,N_16769);
nor U19550 (N_19550,N_15871,N_18047);
and U19551 (N_19551,N_18704,N_16922);
or U19552 (N_19552,N_17734,N_15712);
and U19553 (N_19553,N_17154,N_16913);
or U19554 (N_19554,N_17415,N_17107);
or U19555 (N_19555,N_18560,N_16845);
nor U19556 (N_19556,N_16525,N_15972);
and U19557 (N_19557,N_17130,N_18049);
and U19558 (N_19558,N_17108,N_16447);
and U19559 (N_19559,N_16466,N_15993);
nor U19560 (N_19560,N_17544,N_15637);
xnor U19561 (N_19561,N_17098,N_17303);
nand U19562 (N_19562,N_16351,N_17732);
nand U19563 (N_19563,N_18263,N_18148);
nand U19564 (N_19564,N_17856,N_16994);
and U19565 (N_19565,N_18189,N_17979);
nor U19566 (N_19566,N_17716,N_16873);
and U19567 (N_19567,N_16770,N_18634);
and U19568 (N_19568,N_17789,N_17873);
nand U19569 (N_19569,N_17596,N_15707);
or U19570 (N_19570,N_16348,N_17823);
nand U19571 (N_19571,N_17505,N_16655);
nand U19572 (N_19572,N_17447,N_16941);
xnor U19573 (N_19573,N_16392,N_18618);
nand U19574 (N_19574,N_15625,N_17748);
and U19575 (N_19575,N_16893,N_17465);
or U19576 (N_19576,N_16641,N_15833);
and U19577 (N_19577,N_17008,N_16842);
or U19578 (N_19578,N_18324,N_17876);
and U19579 (N_19579,N_17127,N_18393);
nor U19580 (N_19580,N_17422,N_15706);
nand U19581 (N_19581,N_16548,N_17722);
or U19582 (N_19582,N_17953,N_15742);
nor U19583 (N_19583,N_17609,N_18524);
or U19584 (N_19584,N_16093,N_16280);
or U19585 (N_19585,N_17307,N_17597);
nor U19586 (N_19586,N_17806,N_17504);
nand U19587 (N_19587,N_16182,N_17534);
nand U19588 (N_19588,N_18530,N_17563);
and U19589 (N_19589,N_17330,N_16907);
or U19590 (N_19590,N_16549,N_17614);
or U19591 (N_19591,N_17758,N_15885);
nand U19592 (N_19592,N_17068,N_17832);
nand U19593 (N_19593,N_18382,N_17934);
nor U19594 (N_19594,N_16068,N_18418);
and U19595 (N_19595,N_17697,N_17777);
nor U19596 (N_19596,N_18304,N_18014);
xnor U19597 (N_19597,N_16284,N_17051);
nor U19598 (N_19598,N_17027,N_17846);
nand U19599 (N_19599,N_16717,N_18273);
nor U19600 (N_19600,N_17619,N_15648);
or U19601 (N_19601,N_17691,N_17286);
and U19602 (N_19602,N_15784,N_17728);
nor U19603 (N_19603,N_18363,N_17987);
nor U19604 (N_19604,N_15810,N_16102);
nand U19605 (N_19605,N_17851,N_16012);
nor U19606 (N_19606,N_18120,N_16105);
nor U19607 (N_19607,N_17923,N_16928);
and U19608 (N_19608,N_16706,N_16303);
and U19609 (N_19609,N_18198,N_16418);
nor U19610 (N_19610,N_18290,N_16689);
xor U19611 (N_19611,N_17952,N_18622);
nor U19612 (N_19612,N_15882,N_18248);
nand U19613 (N_19613,N_17380,N_16471);
nand U19614 (N_19614,N_15955,N_17519);
nor U19615 (N_19615,N_16767,N_17955);
nor U19616 (N_19616,N_16784,N_17382);
or U19617 (N_19617,N_17779,N_18022);
or U19618 (N_19618,N_16150,N_18306);
nor U19619 (N_19619,N_17388,N_17560);
nor U19620 (N_19620,N_16649,N_18384);
and U19621 (N_19621,N_16612,N_17043);
and U19622 (N_19622,N_18210,N_17616);
nor U19623 (N_19623,N_17220,N_15663);
nand U19624 (N_19624,N_18179,N_17811);
nor U19625 (N_19625,N_18288,N_15933);
nor U19626 (N_19626,N_16130,N_15892);
nor U19627 (N_19627,N_15856,N_17514);
nor U19628 (N_19628,N_15661,N_16852);
nor U19629 (N_19629,N_18471,N_17225);
nand U19630 (N_19630,N_16070,N_16898);
and U19631 (N_19631,N_18348,N_16114);
nor U19632 (N_19632,N_17026,N_17034);
nor U19633 (N_19633,N_16190,N_16828);
nand U19634 (N_19634,N_17703,N_17074);
nand U19635 (N_19635,N_16537,N_16906);
and U19636 (N_19636,N_17476,N_18316);
nor U19637 (N_19637,N_17033,N_18260);
and U19638 (N_19638,N_18673,N_17132);
nand U19639 (N_19639,N_18458,N_17667);
nor U19640 (N_19640,N_15918,N_16678);
nor U19641 (N_19641,N_18411,N_16446);
and U19642 (N_19642,N_17367,N_16295);
and U19643 (N_19643,N_17111,N_18074);
or U19644 (N_19644,N_18027,N_16212);
xnor U19645 (N_19645,N_18535,N_17284);
or U19646 (N_19646,N_17919,N_17117);
nor U19647 (N_19647,N_16916,N_16107);
or U19648 (N_19648,N_18460,N_17926);
nand U19649 (N_19649,N_16745,N_17146);
and U19650 (N_19650,N_15852,N_17991);
or U19651 (N_19651,N_17084,N_17483);
or U19652 (N_19652,N_17924,N_18044);
and U19653 (N_19653,N_17708,N_16911);
nor U19654 (N_19654,N_18301,N_18506);
and U19655 (N_19655,N_16061,N_15738);
nand U19656 (N_19656,N_17294,N_16154);
and U19657 (N_19657,N_18505,N_16985);
nand U19658 (N_19658,N_15812,N_16206);
nor U19659 (N_19659,N_16054,N_16596);
nor U19660 (N_19660,N_16764,N_16275);
or U19661 (N_19661,N_17376,N_15759);
nand U19662 (N_19662,N_18426,N_18197);
nor U19663 (N_19663,N_17000,N_18154);
or U19664 (N_19664,N_15874,N_18454);
nand U19665 (N_19665,N_15782,N_15847);
nor U19666 (N_19666,N_16535,N_18665);
and U19667 (N_19667,N_17995,N_18676);
or U19668 (N_19668,N_18528,N_17097);
nor U19669 (N_19669,N_15887,N_16585);
and U19670 (N_19670,N_18091,N_15948);
nor U19671 (N_19671,N_17400,N_18653);
nor U19672 (N_19672,N_17518,N_17539);
nor U19673 (N_19673,N_16441,N_18353);
or U19674 (N_19674,N_18453,N_16001);
or U19675 (N_19675,N_18654,N_16322);
and U19676 (N_19676,N_15743,N_16859);
and U19677 (N_19677,N_17797,N_18321);
and U19678 (N_19678,N_15654,N_17183);
or U19679 (N_19679,N_16086,N_18402);
or U19680 (N_19680,N_18720,N_16205);
xor U19681 (N_19681,N_18736,N_17617);
nand U19682 (N_19682,N_17821,N_16635);
xor U19683 (N_19683,N_18553,N_18360);
and U19684 (N_19684,N_18327,N_18496);
nor U19685 (N_19685,N_17344,N_17040);
nand U19686 (N_19686,N_17089,N_18478);
nand U19687 (N_19687,N_16878,N_17364);
nor U19688 (N_19688,N_17547,N_15772);
nand U19689 (N_19689,N_17881,N_16624);
and U19690 (N_19690,N_16236,N_16023);
nand U19691 (N_19691,N_16653,N_16803);
nor U19692 (N_19692,N_16073,N_15873);
nor U19693 (N_19693,N_17365,N_17527);
nand U19694 (N_19694,N_16256,N_17671);
nand U19695 (N_19695,N_17150,N_16851);
xor U19696 (N_19696,N_16036,N_17394);
and U19697 (N_19697,N_16478,N_15921);
or U19698 (N_19698,N_16384,N_18734);
or U19699 (N_19699,N_17768,N_16243);
nor U19700 (N_19700,N_17570,N_18076);
and U19701 (N_19701,N_17094,N_17119);
or U19702 (N_19702,N_16926,N_18289);
or U19703 (N_19703,N_18469,N_17282);
or U19704 (N_19704,N_17964,N_17525);
nor U19705 (N_19705,N_15748,N_16445);
or U19706 (N_19706,N_15971,N_17420);
or U19707 (N_19707,N_18728,N_18225);
nor U19708 (N_19708,N_16473,N_18639);
or U19709 (N_19709,N_18391,N_18388);
or U19710 (N_19710,N_16603,N_17850);
xor U19711 (N_19711,N_18397,N_17838);
and U19712 (N_19712,N_17160,N_18376);
nand U19713 (N_19713,N_15889,N_16321);
and U19714 (N_19714,N_18721,N_17548);
nand U19715 (N_19715,N_17451,N_17157);
and U19716 (N_19716,N_16940,N_15969);
or U19717 (N_19717,N_16429,N_17664);
and U19718 (N_19718,N_15692,N_16983);
nor U19719 (N_19719,N_16448,N_15861);
and U19720 (N_19720,N_17638,N_16771);
or U19721 (N_19721,N_17237,N_17884);
nor U19722 (N_19722,N_18052,N_18407);
or U19723 (N_19723,N_15736,N_16818);
and U19724 (N_19724,N_15975,N_16144);
or U19725 (N_19725,N_16260,N_16354);
nor U19726 (N_19726,N_15640,N_15643);
or U19727 (N_19727,N_18163,N_15916);
nand U19728 (N_19728,N_17313,N_18429);
or U19729 (N_19729,N_18267,N_17868);
nand U19730 (N_19730,N_18275,N_18706);
nand U19731 (N_19731,N_18101,N_15678);
or U19732 (N_19732,N_16185,N_18347);
and U19733 (N_19733,N_18519,N_15788);
xor U19734 (N_19734,N_15780,N_17131);
nand U19735 (N_19735,N_17261,N_16628);
nand U19736 (N_19736,N_16197,N_16088);
or U19737 (N_19737,N_17943,N_17064);
and U19738 (N_19738,N_16199,N_15653);
xor U19739 (N_19739,N_18690,N_17184);
xnor U19740 (N_19740,N_17726,N_15755);
and U19741 (N_19741,N_17677,N_16971);
or U19742 (N_19742,N_16515,N_16760);
or U19743 (N_19743,N_17080,N_16925);
xnor U19744 (N_19744,N_17944,N_15626);
xnor U19745 (N_19745,N_17503,N_18580);
nand U19746 (N_19746,N_18435,N_16746);
or U19747 (N_19747,N_16762,N_17355);
nand U19748 (N_19748,N_17855,N_15768);
nor U19749 (N_19749,N_17970,N_18090);
and U19750 (N_19750,N_17573,N_16417);
or U19751 (N_19751,N_16122,N_18614);
and U19752 (N_19752,N_18042,N_17706);
nand U19753 (N_19753,N_16374,N_18493);
nor U19754 (N_19754,N_18691,N_16410);
or U19755 (N_19755,N_15725,N_16607);
nor U19756 (N_19756,N_18080,N_18525);
and U19757 (N_19757,N_16244,N_15951);
and U19758 (N_19758,N_17336,N_17053);
or U19759 (N_19759,N_18126,N_16613);
and U19760 (N_19760,N_16619,N_16124);
nor U19761 (N_19761,N_16389,N_16451);
nor U19762 (N_19762,N_17575,N_17302);
or U19763 (N_19763,N_17085,N_18473);
nand U19764 (N_19764,N_15803,N_18574);
and U19765 (N_19765,N_16813,N_18028);
and U19766 (N_19766,N_18082,N_16502);
nor U19767 (N_19767,N_17482,N_17231);
nand U19768 (N_19768,N_17727,N_18213);
and U19769 (N_19769,N_17810,N_15781);
and U19770 (N_19770,N_16887,N_17760);
nor U19771 (N_19771,N_16255,N_17234);
nor U19772 (N_19772,N_18079,N_17386);
or U19773 (N_19773,N_15966,N_17696);
nor U19774 (N_19774,N_17712,N_18548);
or U19775 (N_19775,N_15739,N_16900);
nor U19776 (N_19776,N_17452,N_15673);
nor U19777 (N_19777,N_16173,N_15991);
nand U19778 (N_19778,N_15985,N_17729);
or U19779 (N_19779,N_16696,N_18252);
or U19780 (N_19780,N_16915,N_18436);
or U19781 (N_19781,N_17833,N_18230);
or U19782 (N_19782,N_16869,N_17197);
nand U19783 (N_19783,N_17279,N_16228);
and U19784 (N_19784,N_17308,N_17535);
nand U19785 (N_19785,N_18491,N_16988);
xor U19786 (N_19786,N_16091,N_17122);
nor U19787 (N_19787,N_17385,N_18310);
or U19788 (N_19788,N_16896,N_17354);
xor U19789 (N_19789,N_16979,N_18626);
nor U19790 (N_19790,N_16352,N_18320);
or U19791 (N_19791,N_16831,N_17432);
or U19792 (N_19792,N_16367,N_17305);
or U19793 (N_19793,N_18621,N_16356);
or U19794 (N_19794,N_17356,N_16848);
and U19795 (N_19795,N_17246,N_17611);
and U19796 (N_19796,N_16037,N_17077);
nand U19797 (N_19797,N_17021,N_18466);
or U19798 (N_19798,N_18036,N_16433);
and U19799 (N_19799,N_17910,N_18373);
nor U19800 (N_19800,N_18139,N_18237);
or U19801 (N_19801,N_16247,N_17669);
or U19802 (N_19802,N_17263,N_15849);
or U19803 (N_19803,N_17602,N_16752);
nand U19804 (N_19804,N_18483,N_18141);
xor U19805 (N_19805,N_17288,N_18137);
nor U19806 (N_19806,N_15893,N_15688);
nand U19807 (N_19807,N_17381,N_16270);
or U19808 (N_19808,N_18403,N_17060);
nand U19809 (N_19809,N_16734,N_17212);
nor U19810 (N_19810,N_18004,N_18138);
nor U19811 (N_19811,N_17554,N_16806);
nor U19812 (N_19812,N_18637,N_16373);
and U19813 (N_19813,N_16758,N_16421);
nand U19814 (N_19814,N_16892,N_16063);
nor U19815 (N_19815,N_17610,N_15794);
and U19816 (N_19816,N_15959,N_18030);
and U19817 (N_19817,N_16156,N_15895);
nor U19818 (N_19818,N_17704,N_18020);
nor U19819 (N_19819,N_16709,N_15877);
or U19820 (N_19820,N_16330,N_17193);
nand U19821 (N_19821,N_16881,N_17078);
and U19822 (N_19822,N_15818,N_17493);
and U19823 (N_19823,N_17998,N_16544);
and U19824 (N_19824,N_18424,N_18392);
nand U19825 (N_19825,N_18377,N_16132);
or U19826 (N_19826,N_17994,N_16751);
or U19827 (N_19827,N_16291,N_15633);
and U19828 (N_19828,N_17650,N_16609);
or U19829 (N_19829,N_17942,N_16533);
and U19830 (N_19830,N_17781,N_16268);
or U19831 (N_19831,N_16264,N_17783);
nand U19832 (N_19832,N_17945,N_17166);
nand U19833 (N_19833,N_17479,N_15651);
and U19834 (N_19834,N_16226,N_15935);
nand U19835 (N_19835,N_17522,N_16249);
nor U19836 (N_19836,N_16000,N_18358);
nor U19837 (N_19837,N_16474,N_16721);
nand U19838 (N_19838,N_15696,N_16481);
or U19839 (N_19839,N_18693,N_16272);
nor U19840 (N_19840,N_16066,N_15720);
and U19841 (N_19841,N_15686,N_17010);
nand U19842 (N_19842,N_18232,N_15844);
nor U19843 (N_19843,N_17717,N_18281);
and U19844 (N_19844,N_17659,N_17285);
nor U19845 (N_19845,N_16024,N_16277);
nor U19846 (N_19846,N_18236,N_17637);
nor U19847 (N_19847,N_17259,N_18567);
nand U19848 (N_19848,N_15898,N_16316);
and U19849 (N_19849,N_17425,N_17822);
nand U19850 (N_19850,N_17600,N_18202);
nor U19851 (N_19851,N_16523,N_15786);
nand U19852 (N_19852,N_16962,N_17478);
or U19853 (N_19853,N_15746,N_16188);
nand U19854 (N_19854,N_18559,N_15878);
or U19855 (N_19855,N_18277,N_16534);
and U19856 (N_19856,N_17076,N_17341);
or U19857 (N_19857,N_17235,N_18683);
nor U19858 (N_19858,N_16225,N_17217);
or U19859 (N_19859,N_18616,N_17916);
and U19860 (N_19860,N_18749,N_16159);
and U19861 (N_19861,N_15799,N_17393);
and U19862 (N_19862,N_16580,N_18718);
or U19863 (N_19863,N_16267,N_16708);
and U19864 (N_19864,N_16694,N_17387);
nor U19865 (N_19865,N_16191,N_18006);
xnor U19866 (N_19866,N_17044,N_18620);
xnor U19867 (N_19867,N_17719,N_16440);
or U19868 (N_19868,N_17521,N_15628);
and U19869 (N_19869,N_16387,N_16727);
or U19870 (N_19870,N_17038,N_15915);
nand U19871 (N_19871,N_16749,N_18227);
nor U19872 (N_19872,N_18307,N_16516);
and U19873 (N_19873,N_17845,N_15645);
and U19874 (N_19874,N_15802,N_15814);
or U19875 (N_19875,N_15713,N_18125);
and U19876 (N_19876,N_17162,N_16289);
or U19877 (N_19877,N_17266,N_15906);
nor U19878 (N_19878,N_18087,N_17632);
nor U19879 (N_19879,N_17904,N_16406);
nor U19880 (N_19880,N_18472,N_18386);
or U19881 (N_19881,N_16127,N_16469);
xnor U19882 (N_19882,N_17767,N_17250);
or U19883 (N_19883,N_18470,N_17725);
and U19884 (N_19884,N_17176,N_16404);
nor U19885 (N_19885,N_16793,N_17705);
and U19886 (N_19886,N_15980,N_18062);
nor U19887 (N_19887,N_16335,N_17790);
nand U19888 (N_19888,N_15897,N_16136);
nand U19889 (N_19889,N_17446,N_18134);
or U19890 (N_19890,N_18178,N_17073);
or U19891 (N_19891,N_18395,N_15800);
and U19892 (N_19892,N_16031,N_17701);
xnor U19893 (N_19893,N_17321,N_16692);
nor U19894 (N_19894,N_16542,N_18400);
and U19895 (N_19895,N_17541,N_16338);
or U19896 (N_19896,N_17101,N_16671);
xnor U19897 (N_19897,N_17292,N_16904);
or U19898 (N_19898,N_15907,N_16158);
xnor U19899 (N_19899,N_16934,N_16895);
nand U19900 (N_19900,N_17456,N_15816);
or U19901 (N_19901,N_18328,N_17755);
or U19902 (N_19902,N_15726,N_18442);
and U19903 (N_19903,N_17069,N_18053);
xor U19904 (N_19904,N_16665,N_15982);
nor U19905 (N_19905,N_17634,N_16987);
nand U19906 (N_19906,N_17050,N_17103);
nand U19907 (N_19907,N_16493,N_16868);
nor U19908 (N_19908,N_18539,N_18265);
nand U19909 (N_19909,N_16902,N_18207);
nand U19910 (N_19910,N_16162,N_16871);
nor U19911 (N_19911,N_16398,N_17161);
nand U19912 (N_19912,N_18440,N_18543);
and U19913 (N_19913,N_17071,N_17572);
and U19914 (N_19914,N_15627,N_17056);
or U19915 (N_19915,N_15659,N_17769);
and U19916 (N_19916,N_15913,N_17314);
nor U19917 (N_19917,N_18261,N_18029);
or U19918 (N_19918,N_16993,N_17408);
or U19919 (N_19919,N_17358,N_16092);
nor U19920 (N_19920,N_16120,N_15761);
nand U19921 (N_19921,N_16875,N_16229);
or U19922 (N_19922,N_16930,N_15903);
and U19923 (N_19923,N_17721,N_15953);
or U19924 (N_19924,N_16630,N_16973);
nand U19925 (N_19925,N_15901,N_18143);
nor U19926 (N_19926,N_18368,N_17869);
and U19927 (N_19927,N_17167,N_18389);
nand U19928 (N_19928,N_17067,N_17323);
or U19929 (N_19929,N_18578,N_17630);
nor U19930 (N_19930,N_16560,N_17680);
nand U19931 (N_19931,N_18572,N_17255);
or U19932 (N_19932,N_16673,N_16739);
or U19933 (N_19933,N_17349,N_17836);
nor U19934 (N_19934,N_18305,N_18068);
nor U19935 (N_19935,N_18544,N_18104);
nand U19936 (N_19936,N_18329,N_18434);
and U19937 (N_19937,N_15758,N_17273);
nand U19938 (N_19938,N_17502,N_17620);
or U19939 (N_19939,N_18064,N_18191);
and U19940 (N_19940,N_16625,N_17612);
nor U19941 (N_19941,N_17513,N_17022);
nand U19942 (N_19942,N_18246,N_15950);
xnor U19943 (N_19943,N_17023,N_16339);
and U19944 (N_19944,N_16479,N_15721);
or U19945 (N_19945,N_18414,N_18658);
nand U19946 (N_19946,N_17177,N_18127);
nand U19947 (N_19947,N_16593,N_18123);
nand U19948 (N_19948,N_17139,N_17345);
nand U19949 (N_19949,N_17695,N_17936);
nor U19950 (N_19950,N_18067,N_17928);
or U19951 (N_19951,N_17238,N_15815);
or U19952 (N_19952,N_18054,N_18556);
or U19953 (N_19953,N_17931,N_17102);
nor U19954 (N_19954,N_17710,N_18730);
nor U19955 (N_19955,N_16301,N_17605);
or U19956 (N_19956,N_18563,N_16006);
nor U19957 (N_19957,N_16996,N_15938);
xnor U19958 (N_19958,N_18157,N_18420);
xor U19959 (N_19959,N_18396,N_18313);
and U19960 (N_19960,N_17410,N_17269);
or U19961 (N_19961,N_18086,N_18172);
nand U19962 (N_19962,N_15717,N_17772);
and U19963 (N_19963,N_15846,N_16395);
or U19964 (N_19964,N_18441,N_17165);
xor U19965 (N_19965,N_15704,N_16640);
xnor U19966 (N_19966,N_16200,N_17874);
xnor U19967 (N_19967,N_17764,N_17972);
nand U19968 (N_19968,N_17640,N_17120);
and U19969 (N_19969,N_16431,N_17281);
or U19970 (N_19970,N_16211,N_17123);
or U19971 (N_19971,N_18276,N_15724);
nor U19972 (N_19972,N_18605,N_18385);
nand U19973 (N_19973,N_16965,N_16032);
and U19974 (N_19974,N_15910,N_18489);
or U19975 (N_19975,N_17438,N_16657);
nand U19976 (N_19976,N_16886,N_16582);
nand U19977 (N_19977,N_18627,N_16135);
nand U19978 (N_19978,N_15983,N_18647);
nor U19979 (N_19979,N_16319,N_18175);
or U19980 (N_19980,N_16030,N_17564);
and U19981 (N_19981,N_18678,N_18518);
and U19982 (N_19982,N_18269,N_16382);
nor U19983 (N_19983,N_18115,N_16753);
or U19984 (N_19984,N_16647,N_17852);
and U19985 (N_19985,N_18140,N_16016);
and U19986 (N_19986,N_16763,N_18636);
and U19987 (N_19987,N_18511,N_16029);
nand U19988 (N_19988,N_18355,N_15762);
and U19989 (N_19989,N_16808,N_16047);
nand U19990 (N_19990,N_15999,N_15728);
or U19991 (N_19991,N_16358,N_15988);
and U19992 (N_19992,N_17985,N_17604);
and U19993 (N_19993,N_18108,N_18362);
nor U19994 (N_19994,N_18008,N_15940);
and U19995 (N_19995,N_18061,N_16816);
or U19996 (N_19996,N_17579,N_17242);
nor U19997 (N_19997,N_18270,N_17195);
or U19998 (N_19998,N_16050,N_16007);
and U19999 (N_19999,N_16465,N_16304);
and U20000 (N_20000,N_18494,N_18262);
or U20001 (N_20001,N_17315,N_18035);
or U20002 (N_20002,N_18129,N_16341);
nand U20003 (N_20003,N_16110,N_17481);
xnor U20004 (N_20004,N_15986,N_17984);
and U20005 (N_20005,N_17947,N_18040);
nor U20006 (N_20006,N_18731,N_18336);
or U20007 (N_20007,N_16477,N_18650);
nor U20008 (N_20008,N_16812,N_16077);
nor U20009 (N_20009,N_18476,N_18314);
and U20010 (N_20010,N_17920,N_15774);
nand U20011 (N_20011,N_16310,N_18603);
nand U20012 (N_20012,N_15676,N_18187);
or U20013 (N_20013,N_17956,N_17625);
or U20014 (N_20014,N_17464,N_16408);
or U20015 (N_20015,N_16576,N_15835);
or U20016 (N_20016,N_17441,N_16142);
and U20017 (N_20017,N_17862,N_16193);
or U20018 (N_20018,N_18501,N_16528);
and U20019 (N_20019,N_16819,N_18694);
or U20020 (N_20020,N_16065,N_16517);
or U20021 (N_20021,N_17583,N_17844);
nand U20022 (N_20022,N_17566,N_17240);
and U20023 (N_20023,N_18594,N_15888);
xnor U20024 (N_20024,N_16196,N_16227);
nand U20025 (N_20025,N_16572,N_17636);
nor U20026 (N_20026,N_15741,N_18009);
xor U20027 (N_20027,N_17966,N_17338);
or U20028 (N_20028,N_15750,N_17578);
and U20029 (N_20029,N_16078,N_18682);
or U20030 (N_20030,N_18174,N_17427);
nand U20031 (N_20031,N_17798,N_17398);
and U20032 (N_20032,N_17037,N_16317);
or U20033 (N_20033,N_16396,N_16008);
nor U20034 (N_20034,N_17109,N_16165);
and U20035 (N_20035,N_15977,N_18726);
and U20036 (N_20036,N_15819,N_18584);
xor U20037 (N_20037,N_17239,N_16296);
and U20038 (N_20038,N_17216,N_18534);
and U20039 (N_20039,N_16546,N_18503);
or U20040 (N_20040,N_18100,N_17188);
nand U20041 (N_20041,N_18536,N_16218);
and U20042 (N_20042,N_17375,N_18413);
xnor U20043 (N_20043,N_17976,N_17406);
nand U20044 (N_20044,N_18235,N_17230);
or U20045 (N_20045,N_17562,N_16355);
xnor U20046 (N_20046,N_18692,N_18046);
nand U20047 (N_20047,N_18051,N_16880);
and U20048 (N_20048,N_17052,N_17949);
nor U20049 (N_20049,N_17576,N_17207);
nand U20050 (N_20050,N_16698,N_16826);
xnor U20051 (N_20051,N_15790,N_15770);
and U20052 (N_20052,N_18099,N_17244);
nor U20053 (N_20053,N_16145,N_16380);
nand U20054 (N_20054,N_16004,N_16804);
nand U20055 (N_20055,N_18240,N_18128);
and U20056 (N_20056,N_16436,N_16161);
nand U20057 (N_20057,N_16467,N_17935);
nand U20058 (N_20058,N_18124,N_18666);
nor U20059 (N_20059,N_17409,N_17401);
nor U20060 (N_20060,N_18449,N_18255);
and U20061 (N_20061,N_18522,N_18162);
nor U20062 (N_20062,N_18523,N_18282);
and U20063 (N_20063,N_18370,N_16532);
or U20064 (N_20064,N_18180,N_17407);
nor U20065 (N_20065,N_17086,N_17828);
or U20066 (N_20066,N_17318,N_17803);
xnor U20067 (N_20067,N_18513,N_15827);
nand U20068 (N_20068,N_16616,N_18633);
xnor U20069 (N_20069,N_16557,N_17643);
nand U20070 (N_20070,N_16362,N_16094);
nand U20071 (N_20071,N_18331,N_15854);
and U20072 (N_20072,N_16025,N_16148);
or U20073 (N_20073,N_16098,N_17745);
nand U20074 (N_20074,N_17927,N_17202);
or U20075 (N_20075,N_16402,N_16057);
nand U20076 (N_20076,N_15928,N_17264);
xnor U20077 (N_20077,N_18427,N_18643);
and U20078 (N_20078,N_16055,N_16980);
nor U20079 (N_20079,N_16833,N_17672);
nor U20080 (N_20080,N_18107,N_16969);
or U20081 (N_20081,N_18218,N_17384);
nand U20082 (N_20082,N_17782,N_18417);
nand U20083 (N_20083,N_16590,N_16786);
nand U20084 (N_20084,N_16664,N_16857);
nor U20085 (N_20085,N_18317,N_16128);
or U20086 (N_20086,N_18532,N_16543);
nor U20087 (N_20087,N_18350,N_17835);
nand U20088 (N_20088,N_16151,N_16449);
nand U20089 (N_20089,N_18546,N_15631);
xnor U20090 (N_20090,N_16538,N_17948);
and U20091 (N_20091,N_15658,N_18224);
and U20092 (N_20092,N_15909,N_18105);
or U20093 (N_20093,N_16713,N_15825);
nor U20094 (N_20094,N_17668,N_18599);
and U20095 (N_20095,N_17004,N_18425);
and U20096 (N_20096,N_16051,N_16935);
nand U20097 (N_20097,N_17057,N_18135);
nand U20098 (N_20098,N_16232,N_15987);
nand U20099 (N_20099,N_17699,N_15879);
and U20100 (N_20100,N_15843,N_17467);
nand U20101 (N_20101,N_16862,N_18375);
xor U20102 (N_20102,N_18488,N_16986);
and U20103 (N_20103,N_17134,N_16327);
nor U20104 (N_20104,N_15939,N_17556);
nor U20105 (N_20105,N_16564,N_18593);
nor U20106 (N_20106,N_18164,N_15858);
and U20107 (N_20107,N_17079,N_16508);
nor U20108 (N_20108,N_16456,N_17200);
and U20109 (N_20109,N_17568,N_18589);
and U20110 (N_20110,N_16498,N_17889);
nor U20111 (N_20111,N_18078,N_18381);
nor U20112 (N_20112,N_17663,N_18371);
and U20113 (N_20113,N_17260,N_16865);
and U20114 (N_20114,N_16414,N_18480);
and U20115 (N_20115,N_17937,N_16571);
nor U20116 (N_20116,N_17988,N_15703);
and U20117 (N_20117,N_15681,N_17007);
nand U20118 (N_20118,N_15876,N_16656);
nor U20119 (N_20119,N_16430,N_17559);
and U20120 (N_20120,N_17657,N_15754);
and U20121 (N_20121,N_16623,N_18032);
and U20122 (N_20122,N_17489,N_16633);
nor U20123 (N_20123,N_15891,N_18144);
nor U20124 (N_20124,N_16371,N_16106);
xor U20125 (N_20125,N_18672,N_16519);
nor U20126 (N_20126,N_15662,N_18722);
nor U20127 (N_20127,N_17512,N_16305);
nor U20128 (N_20128,N_17254,N_18748);
nor U20129 (N_20129,N_18509,N_17233);
xnor U20130 (N_20130,N_17399,N_16659);
and U20131 (N_20131,N_16730,N_16977);
nand U20132 (N_20132,N_18451,N_16789);
nand U20133 (N_20133,N_15695,N_17316);
xnor U20134 (N_20134,N_16475,N_17473);
nand U20135 (N_20135,N_15629,N_17738);
and U20136 (N_20136,N_17412,N_17523);
nand U20137 (N_20137,N_16334,N_18021);
nand U20138 (N_20138,N_17938,N_17776);
and U20139 (N_20139,N_18687,N_16097);
nor U20140 (N_20140,N_18325,N_16109);
nor U20141 (N_20141,N_16563,N_17960);
nand U20142 (N_20142,N_16285,N_17770);
nand U20143 (N_20143,N_17332,N_17268);
or U20144 (N_20144,N_16326,N_16353);
nor U20145 (N_20145,N_15647,N_15697);
nand U20146 (N_20146,N_17248,N_18194);
or U20147 (N_20147,N_18145,N_16224);
and U20148 (N_20148,N_15832,N_17981);
and U20149 (N_20149,N_18279,N_17055);
nor U20150 (N_20150,N_18203,N_18256);
nand U20151 (N_20151,N_16100,N_17545);
nor U20152 (N_20152,N_17590,N_16214);
xor U20153 (N_20153,N_16271,N_18025);
and U20154 (N_20154,N_17624,N_17346);
nand U20155 (N_20155,N_17431,N_16905);
and U20156 (N_20156,N_16426,N_18285);
nand U20157 (N_20157,N_18023,N_16611);
nand U20158 (N_20158,N_16221,N_16460);
xor U20159 (N_20159,N_17603,N_17128);
xor U20160 (N_20160,N_16592,N_15880);
and U20161 (N_20161,N_16139,N_18502);
xor U20162 (N_20162,N_17480,N_16039);
nor U20163 (N_20163,N_16670,N_17170);
nand U20164 (N_20164,N_15682,N_15727);
or U20165 (N_20165,N_16020,N_16131);
nor U20166 (N_20166,N_18367,N_15989);
nand U20167 (N_20167,N_17289,N_15851);
or U20168 (N_20168,N_16536,N_15718);
or U20169 (N_20169,N_16140,N_16908);
nor U20170 (N_20170,N_18423,N_18735);
and U20171 (N_20171,N_18576,N_17793);
xor U20172 (N_20172,N_18412,N_17662);
or U20173 (N_20173,N_17299,N_17168);
and U20174 (N_20174,N_16119,N_17980);
and U20175 (N_20175,N_18341,N_15709);
nor U20176 (N_20176,N_17329,N_17353);
and U20177 (N_20177,N_17194,N_16921);
and U20178 (N_20178,N_15811,N_18557);
nand U20179 (N_20179,N_16486,N_17654);
nand U20180 (N_20180,N_18165,N_18445);
nand U20181 (N_20181,N_16432,N_17395);
nand U20182 (N_20182,N_17854,N_15639);
nand U20183 (N_20183,N_17593,N_16790);
nor U20184 (N_20184,N_18308,N_17342);
nor U20185 (N_20185,N_16526,N_18335);
xor U20186 (N_20186,N_16601,N_16155);
or U20187 (N_20187,N_16238,N_17218);
nand U20188 (N_20188,N_17794,N_16080);
nor U20189 (N_20189,N_16412,N_15702);
and U20190 (N_20190,N_17199,N_16559);
or U20191 (N_20191,N_16058,N_16219);
and U20192 (N_20192,N_18669,N_16409);
or U20193 (N_20193,N_16044,N_16759);
nor U20194 (N_20194,N_18450,N_17509);
and U20195 (N_20195,N_16113,N_16308);
nor U20196 (N_20196,N_18011,N_15970);
nor U20197 (N_20197,N_17357,N_16491);
and U20198 (N_20198,N_16507,N_16835);
and U20199 (N_20199,N_17372,N_17011);
or U20200 (N_20200,N_17417,N_17627);
and U20201 (N_20201,N_18387,N_18547);
nor U20202 (N_20202,N_16125,N_17709);
nand U20203 (N_20203,N_15638,N_17751);
nand U20204 (N_20204,N_18575,N_18733);
nand U20205 (N_20205,N_16932,N_16463);
nor U20206 (N_20206,N_17334,N_17436);
and U20207 (N_20207,N_17574,N_17135);
nand U20208 (N_20208,N_16038,N_17317);
and U20209 (N_20209,N_18507,N_16814);
or U20210 (N_20210,N_16942,N_17901);
nor U20211 (N_20211,N_16399,N_16959);
or U20212 (N_20212,N_18587,N_17774);
nor U20213 (N_20213,N_17439,N_16610);
nand U20214 (N_20214,N_15669,N_17820);
nor U20215 (N_20215,N_18315,N_15900);
nand U20216 (N_20216,N_17688,N_17270);
nand U20217 (N_20217,N_17658,N_17546);
nor U20218 (N_20218,N_16452,N_15693);
or U20219 (N_20219,N_18272,N_18719);
nand U20220 (N_20220,N_18201,N_17378);
or U20221 (N_20221,N_17753,N_18571);
and U20222 (N_20222,N_17046,N_17675);
and U20223 (N_20223,N_16910,N_17999);
nand U20224 (N_20224,N_16724,N_15679);
and U20225 (N_20225,N_17613,N_17549);
nand U20226 (N_20226,N_17741,N_17013);
xor U20227 (N_20227,N_16472,N_18679);
xor U20228 (N_20228,N_17571,N_16858);
nand U20229 (N_20229,N_16522,N_15752);
nand U20230 (N_20230,N_18231,N_18508);
and U20231 (N_20231,N_18623,N_17540);
nand U20232 (N_20232,N_17484,N_18059);
nand U20233 (N_20233,N_16849,N_17253);
and U20234 (N_20234,N_15700,N_17133);
and U20235 (N_20235,N_16187,N_16035);
xnor U20236 (N_20236,N_18715,N_16253);
or U20237 (N_20237,N_16422,N_18223);
nand U20238 (N_20238,N_18448,N_16622);
nor U20239 (N_20239,N_16257,N_17301);
or U20240 (N_20240,N_18026,N_17537);
or U20241 (N_20241,N_17377,N_16318);
nand U20242 (N_20242,N_15805,N_18568);
and U20243 (N_20243,N_17002,N_16485);
nand U20244 (N_20244,N_17428,N_18274);
nand U20245 (N_20245,N_15974,N_16210);
and U20246 (N_20246,N_16788,N_17072);
nand U20247 (N_20247,N_17490,N_17443);
nand U20248 (N_20248,N_15995,N_18297);
and U20249 (N_20249,N_17968,N_17744);
nor U20250 (N_20250,N_16391,N_15867);
and U20251 (N_20251,N_15997,N_17932);
nor U20252 (N_20252,N_18611,N_17581);
and U20253 (N_20253,N_17096,N_18725);
xnor U20254 (N_20254,N_17403,N_18430);
xnor U20255 (N_20255,N_16550,N_17933);
and U20256 (N_20256,N_16939,N_18176);
and U20257 (N_20257,N_17914,N_16177);
nor U20258 (N_20258,N_16682,N_17588);
nand U20259 (N_20259,N_16684,N_18717);
and U20260 (N_20260,N_16732,N_15863);
nor U20261 (N_20261,N_15807,N_15664);
nor U20262 (N_20262,N_16254,N_18149);
and U20263 (N_20263,N_16820,N_15729);
and U20264 (N_20264,N_17510,N_17099);
nand U20265 (N_20265,N_16081,N_15671);
xor U20266 (N_20266,N_15756,N_16438);
and U20267 (N_20267,N_18340,N_16854);
or U20268 (N_20268,N_17682,N_16661);
nor U20269 (N_20269,N_17586,N_16279);
nand U20270 (N_20270,N_16917,N_16700);
nand U20271 (N_20271,N_16824,N_16019);
nand U20272 (N_20272,N_18200,N_18170);
nand U20273 (N_20273,N_17172,N_18649);
or U20274 (N_20274,N_18745,N_18238);
or U20275 (N_20275,N_17750,N_18482);
nand U20276 (N_20276,N_17917,N_18569);
or U20277 (N_20277,N_17814,N_17434);
nor U20278 (N_20278,N_16434,N_17396);
nor U20279 (N_20279,N_18570,N_17059);
and U20280 (N_20280,N_18150,N_17496);
or U20281 (N_20281,N_16626,N_15870);
nor U20282 (N_20282,N_16681,N_18243);
nor U20283 (N_20283,N_17106,N_17860);
or U20284 (N_20284,N_18258,N_15760);
nor U20285 (N_20285,N_15884,N_16089);
or U20286 (N_20286,N_18342,N_17599);
nand U20287 (N_20287,N_15979,N_16676);
xnor U20288 (N_20288,N_17262,N_17645);
nor U20289 (N_20289,N_18512,N_16863);
nor U20290 (N_20290,N_18098,N_15655);
and U20291 (N_20291,N_17061,N_16978);
and U20292 (N_20292,N_16435,N_15883);
nand U20293 (N_20293,N_17796,N_18334);
or U20294 (N_20294,N_17017,N_17982);
or U20295 (N_20295,N_16579,N_16297);
nor U20296 (N_20296,N_17804,N_17005);
nand U20297 (N_20297,N_17178,N_16022);
nand U20298 (N_20298,N_17205,N_15813);
xnor U20299 (N_20299,N_17226,N_16531);
nand U20300 (N_20300,N_16853,N_16815);
nand U20301 (N_20301,N_15904,N_17070);
nand U20302 (N_20302,N_16918,N_18015);
or U20303 (N_20303,N_15698,N_18703);
nand U20304 (N_20304,N_16201,N_15914);
nor U20305 (N_20305,N_18713,N_18486);
and U20306 (N_20306,N_17498,N_16787);
and U20307 (N_20307,N_18520,N_16171);
and U20308 (N_20308,N_17236,N_17799);
nor U20309 (N_20309,N_18629,N_15926);
or U20310 (N_20310,N_16747,N_16266);
nand U20311 (N_20311,N_18742,N_17369);
nor U20312 (N_20312,N_17322,N_15913);
nor U20313 (N_20313,N_18488,N_16728);
nor U20314 (N_20314,N_15686,N_16511);
xnor U20315 (N_20315,N_18454,N_17543);
xnor U20316 (N_20316,N_17136,N_16446);
xnor U20317 (N_20317,N_17829,N_18298);
and U20318 (N_20318,N_18698,N_16345);
and U20319 (N_20319,N_18011,N_18052);
or U20320 (N_20320,N_16436,N_17071);
nor U20321 (N_20321,N_15840,N_16561);
or U20322 (N_20322,N_17296,N_17755);
or U20323 (N_20323,N_16038,N_17672);
xnor U20324 (N_20324,N_18351,N_16804);
nand U20325 (N_20325,N_16005,N_16849);
and U20326 (N_20326,N_18336,N_17096);
xor U20327 (N_20327,N_18106,N_17597);
nor U20328 (N_20328,N_18407,N_17946);
or U20329 (N_20329,N_17124,N_18533);
and U20330 (N_20330,N_17409,N_17562);
nand U20331 (N_20331,N_16102,N_18062);
nand U20332 (N_20332,N_17523,N_16667);
or U20333 (N_20333,N_18565,N_16946);
xor U20334 (N_20334,N_15641,N_18014);
nor U20335 (N_20335,N_17706,N_16729);
or U20336 (N_20336,N_17187,N_16108);
and U20337 (N_20337,N_18422,N_17247);
and U20338 (N_20338,N_17956,N_16834);
or U20339 (N_20339,N_16853,N_18124);
or U20340 (N_20340,N_17176,N_18646);
nor U20341 (N_20341,N_17541,N_17650);
nor U20342 (N_20342,N_16849,N_15826);
and U20343 (N_20343,N_15712,N_15752);
xnor U20344 (N_20344,N_16869,N_18412);
or U20345 (N_20345,N_17042,N_17665);
nor U20346 (N_20346,N_16923,N_17646);
and U20347 (N_20347,N_16155,N_15663);
nand U20348 (N_20348,N_16075,N_16914);
xor U20349 (N_20349,N_18163,N_15653);
xnor U20350 (N_20350,N_17620,N_17120);
or U20351 (N_20351,N_17232,N_15928);
and U20352 (N_20352,N_16814,N_17056);
nor U20353 (N_20353,N_17393,N_18191);
nor U20354 (N_20354,N_17813,N_17218);
and U20355 (N_20355,N_18494,N_17882);
and U20356 (N_20356,N_17647,N_16598);
and U20357 (N_20357,N_17262,N_16132);
and U20358 (N_20358,N_16935,N_17305);
or U20359 (N_20359,N_17676,N_18003);
or U20360 (N_20360,N_16355,N_16542);
nor U20361 (N_20361,N_18062,N_15882);
and U20362 (N_20362,N_15803,N_18476);
nor U20363 (N_20363,N_18132,N_17202);
xor U20364 (N_20364,N_15862,N_15803);
nand U20365 (N_20365,N_17374,N_18587);
or U20366 (N_20366,N_15956,N_16131);
nor U20367 (N_20367,N_16360,N_18198);
and U20368 (N_20368,N_18056,N_17163);
or U20369 (N_20369,N_15829,N_18396);
or U20370 (N_20370,N_17209,N_15691);
nand U20371 (N_20371,N_16073,N_16026);
nand U20372 (N_20372,N_17656,N_16488);
nand U20373 (N_20373,N_18554,N_18503);
xor U20374 (N_20374,N_18443,N_15998);
or U20375 (N_20375,N_16140,N_17270);
nor U20376 (N_20376,N_16744,N_17329);
or U20377 (N_20377,N_18523,N_16531);
and U20378 (N_20378,N_18380,N_17786);
nor U20379 (N_20379,N_17100,N_17449);
and U20380 (N_20380,N_16162,N_16243);
and U20381 (N_20381,N_15910,N_15841);
nor U20382 (N_20382,N_16247,N_18636);
nand U20383 (N_20383,N_16937,N_18271);
and U20384 (N_20384,N_17670,N_17336);
or U20385 (N_20385,N_18405,N_17800);
nor U20386 (N_20386,N_16716,N_16251);
or U20387 (N_20387,N_17314,N_18277);
nor U20388 (N_20388,N_16947,N_16012);
nand U20389 (N_20389,N_16890,N_18178);
and U20390 (N_20390,N_16145,N_17006);
or U20391 (N_20391,N_17873,N_17450);
nand U20392 (N_20392,N_15718,N_15731);
xnor U20393 (N_20393,N_15790,N_16726);
or U20394 (N_20394,N_16894,N_15969);
nor U20395 (N_20395,N_17174,N_18370);
or U20396 (N_20396,N_17962,N_16996);
nor U20397 (N_20397,N_16798,N_15749);
and U20398 (N_20398,N_18634,N_18323);
nand U20399 (N_20399,N_16186,N_17751);
nand U20400 (N_20400,N_18234,N_18230);
nand U20401 (N_20401,N_18719,N_15943);
nor U20402 (N_20402,N_17930,N_18457);
nand U20403 (N_20403,N_16559,N_17298);
nor U20404 (N_20404,N_15722,N_17460);
nand U20405 (N_20405,N_16224,N_17252);
and U20406 (N_20406,N_18508,N_17713);
nand U20407 (N_20407,N_18157,N_18446);
nand U20408 (N_20408,N_16890,N_15821);
and U20409 (N_20409,N_15916,N_16767);
nand U20410 (N_20410,N_18223,N_18246);
or U20411 (N_20411,N_18308,N_16094);
and U20412 (N_20412,N_18712,N_18139);
or U20413 (N_20413,N_18600,N_17578);
nand U20414 (N_20414,N_16279,N_17082);
or U20415 (N_20415,N_17014,N_16409);
or U20416 (N_20416,N_18426,N_18668);
or U20417 (N_20417,N_18703,N_16467);
nand U20418 (N_20418,N_17324,N_17134);
nor U20419 (N_20419,N_17843,N_18027);
or U20420 (N_20420,N_16135,N_16673);
or U20421 (N_20421,N_17672,N_17565);
xnor U20422 (N_20422,N_15961,N_18373);
nor U20423 (N_20423,N_17505,N_17236);
or U20424 (N_20424,N_16470,N_18450);
xor U20425 (N_20425,N_17462,N_18080);
or U20426 (N_20426,N_17988,N_17451);
or U20427 (N_20427,N_15772,N_17899);
nand U20428 (N_20428,N_15654,N_17816);
nor U20429 (N_20429,N_17678,N_15887);
nand U20430 (N_20430,N_17387,N_18727);
or U20431 (N_20431,N_17759,N_17401);
nand U20432 (N_20432,N_18236,N_16854);
or U20433 (N_20433,N_15743,N_16247);
and U20434 (N_20434,N_17428,N_16156);
and U20435 (N_20435,N_17425,N_15962);
nand U20436 (N_20436,N_16700,N_16868);
and U20437 (N_20437,N_16539,N_17279);
xor U20438 (N_20438,N_16893,N_16635);
xnor U20439 (N_20439,N_17897,N_16441);
nor U20440 (N_20440,N_17005,N_15722);
nor U20441 (N_20441,N_16050,N_16562);
nand U20442 (N_20442,N_15816,N_15890);
nand U20443 (N_20443,N_17088,N_16369);
nand U20444 (N_20444,N_18121,N_17115);
nand U20445 (N_20445,N_17286,N_18551);
or U20446 (N_20446,N_17676,N_15880);
or U20447 (N_20447,N_17712,N_17883);
or U20448 (N_20448,N_17772,N_16726);
nand U20449 (N_20449,N_17197,N_17259);
xnor U20450 (N_20450,N_16169,N_16045);
nor U20451 (N_20451,N_17765,N_16468);
or U20452 (N_20452,N_15959,N_16023);
nand U20453 (N_20453,N_16069,N_16884);
nor U20454 (N_20454,N_17955,N_16943);
or U20455 (N_20455,N_18555,N_18465);
or U20456 (N_20456,N_16475,N_16564);
and U20457 (N_20457,N_16765,N_17485);
nor U20458 (N_20458,N_17644,N_17269);
nor U20459 (N_20459,N_18114,N_16721);
or U20460 (N_20460,N_17355,N_17474);
and U20461 (N_20461,N_15931,N_18154);
nor U20462 (N_20462,N_17833,N_15823);
xnor U20463 (N_20463,N_16205,N_17586);
or U20464 (N_20464,N_17786,N_18140);
or U20465 (N_20465,N_17433,N_18649);
xnor U20466 (N_20466,N_17232,N_18410);
nor U20467 (N_20467,N_16418,N_16194);
nand U20468 (N_20468,N_16235,N_15704);
and U20469 (N_20469,N_16219,N_17225);
nor U20470 (N_20470,N_17321,N_16096);
and U20471 (N_20471,N_16880,N_18740);
nand U20472 (N_20472,N_18414,N_15915);
and U20473 (N_20473,N_18389,N_16233);
xor U20474 (N_20474,N_17181,N_16723);
nand U20475 (N_20475,N_18478,N_17617);
nor U20476 (N_20476,N_18148,N_15731);
nor U20477 (N_20477,N_16030,N_16045);
and U20478 (N_20478,N_18702,N_18401);
and U20479 (N_20479,N_16598,N_17327);
xor U20480 (N_20480,N_17713,N_18448);
nand U20481 (N_20481,N_18637,N_16009);
or U20482 (N_20482,N_17042,N_15970);
and U20483 (N_20483,N_15825,N_16744);
nor U20484 (N_20484,N_18101,N_18370);
and U20485 (N_20485,N_18621,N_16547);
nand U20486 (N_20486,N_16452,N_17420);
or U20487 (N_20487,N_17975,N_18456);
or U20488 (N_20488,N_16658,N_17395);
nand U20489 (N_20489,N_17273,N_16552);
and U20490 (N_20490,N_17124,N_16227);
and U20491 (N_20491,N_17577,N_18022);
nand U20492 (N_20492,N_15762,N_17226);
and U20493 (N_20493,N_17045,N_17856);
and U20494 (N_20494,N_18592,N_16395);
nor U20495 (N_20495,N_17615,N_17252);
and U20496 (N_20496,N_16706,N_17501);
nand U20497 (N_20497,N_16980,N_17819);
or U20498 (N_20498,N_16098,N_16944);
xor U20499 (N_20499,N_17692,N_17772);
xor U20500 (N_20500,N_16135,N_17273);
xor U20501 (N_20501,N_17893,N_16360);
nor U20502 (N_20502,N_16845,N_16526);
nor U20503 (N_20503,N_16573,N_16801);
or U20504 (N_20504,N_16134,N_17583);
and U20505 (N_20505,N_16589,N_15863);
nor U20506 (N_20506,N_17121,N_15906);
nand U20507 (N_20507,N_16282,N_18087);
or U20508 (N_20508,N_16252,N_16218);
xor U20509 (N_20509,N_17413,N_17793);
or U20510 (N_20510,N_17829,N_16359);
or U20511 (N_20511,N_16840,N_16995);
or U20512 (N_20512,N_16254,N_17672);
nand U20513 (N_20513,N_18262,N_16960);
nor U20514 (N_20514,N_17235,N_17538);
nor U20515 (N_20515,N_18374,N_16170);
nor U20516 (N_20516,N_18642,N_15695);
and U20517 (N_20517,N_16081,N_17651);
and U20518 (N_20518,N_17240,N_17421);
and U20519 (N_20519,N_18647,N_16337);
and U20520 (N_20520,N_18380,N_18264);
nor U20521 (N_20521,N_16643,N_18259);
or U20522 (N_20522,N_17699,N_17951);
or U20523 (N_20523,N_18552,N_16910);
xor U20524 (N_20524,N_15884,N_17961);
nor U20525 (N_20525,N_16978,N_16449);
nand U20526 (N_20526,N_17665,N_16084);
and U20527 (N_20527,N_16190,N_18742);
and U20528 (N_20528,N_16211,N_17996);
or U20529 (N_20529,N_16904,N_15985);
xnor U20530 (N_20530,N_18050,N_18056);
or U20531 (N_20531,N_15655,N_17338);
or U20532 (N_20532,N_16195,N_17952);
or U20533 (N_20533,N_15969,N_17631);
xnor U20534 (N_20534,N_16581,N_17985);
nand U20535 (N_20535,N_17456,N_17951);
and U20536 (N_20536,N_16382,N_18194);
or U20537 (N_20537,N_18084,N_15934);
xor U20538 (N_20538,N_18351,N_17195);
nor U20539 (N_20539,N_18380,N_16377);
or U20540 (N_20540,N_17854,N_18528);
and U20541 (N_20541,N_16199,N_17500);
nor U20542 (N_20542,N_17744,N_16492);
or U20543 (N_20543,N_17825,N_16632);
or U20544 (N_20544,N_17246,N_18643);
nor U20545 (N_20545,N_15650,N_18269);
xnor U20546 (N_20546,N_17545,N_17513);
nor U20547 (N_20547,N_16031,N_15816);
or U20548 (N_20548,N_16434,N_18217);
nor U20549 (N_20549,N_17126,N_15955);
nor U20550 (N_20550,N_18636,N_16845);
or U20551 (N_20551,N_18113,N_17423);
or U20552 (N_20552,N_17537,N_17042);
nand U20553 (N_20553,N_16633,N_18316);
and U20554 (N_20554,N_18120,N_18003);
xnor U20555 (N_20555,N_16626,N_16300);
nand U20556 (N_20556,N_16616,N_15882);
nand U20557 (N_20557,N_18605,N_17413);
nand U20558 (N_20558,N_16856,N_17328);
nor U20559 (N_20559,N_18666,N_16442);
nand U20560 (N_20560,N_16549,N_18048);
xor U20561 (N_20561,N_16318,N_17192);
nor U20562 (N_20562,N_16298,N_16831);
and U20563 (N_20563,N_16676,N_17641);
nor U20564 (N_20564,N_17577,N_16990);
or U20565 (N_20565,N_16414,N_16382);
nor U20566 (N_20566,N_15869,N_17299);
and U20567 (N_20567,N_16308,N_17027);
and U20568 (N_20568,N_16610,N_16606);
xor U20569 (N_20569,N_15645,N_15954);
or U20570 (N_20570,N_16651,N_18731);
and U20571 (N_20571,N_17323,N_16879);
nor U20572 (N_20572,N_16011,N_17960);
xnor U20573 (N_20573,N_15846,N_18141);
nor U20574 (N_20574,N_18061,N_18328);
or U20575 (N_20575,N_18416,N_17581);
nor U20576 (N_20576,N_16910,N_17549);
and U20577 (N_20577,N_17462,N_16537);
nand U20578 (N_20578,N_17489,N_16038);
or U20579 (N_20579,N_15860,N_18356);
nor U20580 (N_20580,N_18191,N_16956);
nor U20581 (N_20581,N_17859,N_18078);
nand U20582 (N_20582,N_15877,N_18147);
nand U20583 (N_20583,N_17006,N_18472);
nor U20584 (N_20584,N_15745,N_17142);
and U20585 (N_20585,N_17355,N_15968);
nor U20586 (N_20586,N_17037,N_18333);
or U20587 (N_20587,N_17211,N_18400);
nor U20588 (N_20588,N_16616,N_16410);
xor U20589 (N_20589,N_17548,N_15735);
or U20590 (N_20590,N_17680,N_15637);
nor U20591 (N_20591,N_17394,N_15784);
and U20592 (N_20592,N_18095,N_16458);
nor U20593 (N_20593,N_18353,N_16814);
xnor U20594 (N_20594,N_17131,N_16350);
xnor U20595 (N_20595,N_18054,N_18227);
nand U20596 (N_20596,N_16422,N_17983);
nand U20597 (N_20597,N_18240,N_17438);
or U20598 (N_20598,N_17927,N_17135);
nor U20599 (N_20599,N_15646,N_18727);
and U20600 (N_20600,N_17838,N_18339);
nor U20601 (N_20601,N_17211,N_17608);
or U20602 (N_20602,N_16715,N_15745);
or U20603 (N_20603,N_16881,N_17674);
nand U20604 (N_20604,N_16885,N_17495);
xor U20605 (N_20605,N_17877,N_16977);
and U20606 (N_20606,N_17963,N_16208);
and U20607 (N_20607,N_17869,N_18093);
and U20608 (N_20608,N_16124,N_18333);
and U20609 (N_20609,N_18284,N_17629);
nand U20610 (N_20610,N_16586,N_16769);
nor U20611 (N_20611,N_17571,N_17548);
nor U20612 (N_20612,N_17628,N_16216);
or U20613 (N_20613,N_17996,N_17527);
xnor U20614 (N_20614,N_16556,N_16652);
nor U20615 (N_20615,N_16474,N_17477);
nand U20616 (N_20616,N_18284,N_17330);
and U20617 (N_20617,N_16800,N_18094);
and U20618 (N_20618,N_17145,N_16924);
or U20619 (N_20619,N_16910,N_18040);
xnor U20620 (N_20620,N_15635,N_16898);
or U20621 (N_20621,N_15647,N_16498);
or U20622 (N_20622,N_18193,N_17623);
or U20623 (N_20623,N_17825,N_17844);
and U20624 (N_20624,N_16085,N_15843);
nand U20625 (N_20625,N_18384,N_17846);
and U20626 (N_20626,N_18683,N_17918);
or U20627 (N_20627,N_18298,N_17296);
xor U20628 (N_20628,N_15731,N_16268);
nand U20629 (N_20629,N_17141,N_17149);
nand U20630 (N_20630,N_16486,N_16612);
nor U20631 (N_20631,N_17911,N_16537);
or U20632 (N_20632,N_18360,N_16671);
nand U20633 (N_20633,N_17114,N_17511);
nand U20634 (N_20634,N_16347,N_17502);
nor U20635 (N_20635,N_18592,N_17979);
xor U20636 (N_20636,N_18363,N_16659);
nor U20637 (N_20637,N_18506,N_18419);
xor U20638 (N_20638,N_17098,N_16419);
nand U20639 (N_20639,N_18145,N_17126);
and U20640 (N_20640,N_17764,N_17294);
nand U20641 (N_20641,N_17765,N_16653);
nand U20642 (N_20642,N_18123,N_17745);
and U20643 (N_20643,N_17772,N_16072);
nor U20644 (N_20644,N_18374,N_17734);
nand U20645 (N_20645,N_15723,N_17823);
and U20646 (N_20646,N_17785,N_16629);
nor U20647 (N_20647,N_17383,N_17037);
or U20648 (N_20648,N_18049,N_15939);
and U20649 (N_20649,N_16151,N_16226);
or U20650 (N_20650,N_17281,N_16661);
nor U20651 (N_20651,N_18615,N_16772);
nand U20652 (N_20652,N_17355,N_17502);
or U20653 (N_20653,N_18125,N_17125);
and U20654 (N_20654,N_16335,N_16955);
and U20655 (N_20655,N_18643,N_17329);
or U20656 (N_20656,N_16817,N_17823);
xnor U20657 (N_20657,N_18548,N_16237);
or U20658 (N_20658,N_17270,N_17637);
nor U20659 (N_20659,N_16320,N_18460);
nand U20660 (N_20660,N_16462,N_18697);
or U20661 (N_20661,N_16367,N_15739);
and U20662 (N_20662,N_16010,N_16757);
nand U20663 (N_20663,N_18116,N_17422);
and U20664 (N_20664,N_15756,N_17622);
and U20665 (N_20665,N_17913,N_16980);
or U20666 (N_20666,N_17559,N_15639);
or U20667 (N_20667,N_17783,N_16137);
and U20668 (N_20668,N_18589,N_18328);
nor U20669 (N_20669,N_18326,N_16909);
nand U20670 (N_20670,N_17149,N_17780);
and U20671 (N_20671,N_18736,N_17242);
or U20672 (N_20672,N_17496,N_17902);
xor U20673 (N_20673,N_15981,N_16388);
nand U20674 (N_20674,N_16398,N_17549);
or U20675 (N_20675,N_15766,N_17561);
and U20676 (N_20676,N_18257,N_17696);
and U20677 (N_20677,N_17333,N_16931);
and U20678 (N_20678,N_17749,N_15971);
and U20679 (N_20679,N_18268,N_17591);
or U20680 (N_20680,N_18135,N_16976);
nand U20681 (N_20681,N_17590,N_16217);
nor U20682 (N_20682,N_16584,N_16961);
nor U20683 (N_20683,N_17381,N_17123);
xor U20684 (N_20684,N_17860,N_18586);
nor U20685 (N_20685,N_16657,N_16015);
and U20686 (N_20686,N_17777,N_18052);
nand U20687 (N_20687,N_16639,N_18632);
and U20688 (N_20688,N_16180,N_17654);
nand U20689 (N_20689,N_18342,N_16131);
or U20690 (N_20690,N_16293,N_17492);
nor U20691 (N_20691,N_17441,N_16674);
and U20692 (N_20692,N_16111,N_16290);
and U20693 (N_20693,N_15969,N_17962);
or U20694 (N_20694,N_16642,N_15970);
or U20695 (N_20695,N_18601,N_18511);
nand U20696 (N_20696,N_15691,N_16909);
nor U20697 (N_20697,N_17475,N_17451);
and U20698 (N_20698,N_18662,N_17257);
nand U20699 (N_20699,N_17338,N_16771);
nand U20700 (N_20700,N_17583,N_15673);
nor U20701 (N_20701,N_16263,N_15670);
and U20702 (N_20702,N_16321,N_17778);
nor U20703 (N_20703,N_16469,N_15998);
or U20704 (N_20704,N_18176,N_18186);
or U20705 (N_20705,N_16432,N_16111);
or U20706 (N_20706,N_16555,N_18678);
nor U20707 (N_20707,N_18499,N_17892);
and U20708 (N_20708,N_17442,N_17977);
nand U20709 (N_20709,N_16755,N_17143);
or U20710 (N_20710,N_16647,N_16480);
or U20711 (N_20711,N_16389,N_16782);
and U20712 (N_20712,N_16004,N_18132);
nor U20713 (N_20713,N_17494,N_17794);
nor U20714 (N_20714,N_17949,N_17321);
xor U20715 (N_20715,N_16838,N_17968);
xnor U20716 (N_20716,N_18587,N_17638);
or U20717 (N_20717,N_18565,N_16168);
nor U20718 (N_20718,N_15727,N_15785);
nor U20719 (N_20719,N_17989,N_16403);
nand U20720 (N_20720,N_17205,N_16287);
and U20721 (N_20721,N_16575,N_17589);
and U20722 (N_20722,N_17146,N_18675);
and U20723 (N_20723,N_16524,N_16343);
or U20724 (N_20724,N_15648,N_17626);
xor U20725 (N_20725,N_16281,N_18699);
or U20726 (N_20726,N_16084,N_17323);
nor U20727 (N_20727,N_18705,N_18185);
nor U20728 (N_20728,N_17615,N_16550);
nor U20729 (N_20729,N_18336,N_17876);
nor U20730 (N_20730,N_17223,N_18463);
nand U20731 (N_20731,N_16100,N_15647);
nor U20732 (N_20732,N_16888,N_17798);
nand U20733 (N_20733,N_18296,N_17420);
nor U20734 (N_20734,N_15796,N_15710);
nor U20735 (N_20735,N_18700,N_18070);
nand U20736 (N_20736,N_16667,N_16193);
and U20737 (N_20737,N_15830,N_16668);
nor U20738 (N_20738,N_18322,N_18594);
or U20739 (N_20739,N_18644,N_16498);
nor U20740 (N_20740,N_16999,N_16709);
nor U20741 (N_20741,N_16456,N_16239);
nand U20742 (N_20742,N_15992,N_15672);
and U20743 (N_20743,N_16330,N_16079);
nor U20744 (N_20744,N_16439,N_15775);
nor U20745 (N_20745,N_17745,N_17031);
xor U20746 (N_20746,N_15989,N_15818);
xnor U20747 (N_20747,N_17953,N_17901);
and U20748 (N_20748,N_16070,N_18205);
xor U20749 (N_20749,N_15761,N_17721);
xnor U20750 (N_20750,N_16484,N_17256);
nor U20751 (N_20751,N_16543,N_16076);
nand U20752 (N_20752,N_15684,N_17452);
nor U20753 (N_20753,N_17497,N_16466);
nor U20754 (N_20754,N_15658,N_18103);
xnor U20755 (N_20755,N_16256,N_18695);
nand U20756 (N_20756,N_18511,N_16374);
xor U20757 (N_20757,N_18730,N_16669);
and U20758 (N_20758,N_17769,N_17061);
nor U20759 (N_20759,N_16007,N_17584);
or U20760 (N_20760,N_17427,N_17418);
nand U20761 (N_20761,N_17090,N_17229);
nor U20762 (N_20762,N_16738,N_18472);
nor U20763 (N_20763,N_18208,N_18605);
or U20764 (N_20764,N_15688,N_16662);
nor U20765 (N_20765,N_18131,N_15665);
or U20766 (N_20766,N_15758,N_16834);
and U20767 (N_20767,N_18600,N_15989);
nor U20768 (N_20768,N_17946,N_18649);
and U20769 (N_20769,N_16624,N_16322);
and U20770 (N_20770,N_18061,N_16990);
and U20771 (N_20771,N_17429,N_17437);
xnor U20772 (N_20772,N_18591,N_16457);
or U20773 (N_20773,N_18043,N_16643);
nor U20774 (N_20774,N_17330,N_15816);
or U20775 (N_20775,N_17911,N_18286);
nand U20776 (N_20776,N_17353,N_16818);
and U20777 (N_20777,N_18728,N_18105);
or U20778 (N_20778,N_17354,N_17262);
and U20779 (N_20779,N_17995,N_17596);
xnor U20780 (N_20780,N_18150,N_15898);
nand U20781 (N_20781,N_15869,N_15858);
nor U20782 (N_20782,N_18061,N_16455);
or U20783 (N_20783,N_17998,N_16491);
nand U20784 (N_20784,N_17324,N_16983);
and U20785 (N_20785,N_16054,N_17942);
nand U20786 (N_20786,N_17688,N_16719);
or U20787 (N_20787,N_17356,N_16567);
nand U20788 (N_20788,N_17154,N_17627);
and U20789 (N_20789,N_16752,N_17878);
and U20790 (N_20790,N_16569,N_18549);
nand U20791 (N_20791,N_15814,N_18035);
nand U20792 (N_20792,N_17607,N_17979);
or U20793 (N_20793,N_15948,N_17810);
nor U20794 (N_20794,N_18455,N_17053);
and U20795 (N_20795,N_16621,N_17371);
nand U20796 (N_20796,N_17395,N_18531);
nor U20797 (N_20797,N_18502,N_17826);
and U20798 (N_20798,N_17441,N_16614);
or U20799 (N_20799,N_17090,N_17723);
nor U20800 (N_20800,N_18651,N_18027);
nor U20801 (N_20801,N_17007,N_17714);
nand U20802 (N_20802,N_17038,N_15801);
or U20803 (N_20803,N_15634,N_17872);
nor U20804 (N_20804,N_17063,N_17611);
nor U20805 (N_20805,N_18474,N_17170);
xnor U20806 (N_20806,N_18437,N_17888);
nand U20807 (N_20807,N_17284,N_17183);
nand U20808 (N_20808,N_16736,N_17248);
xor U20809 (N_20809,N_18211,N_18729);
and U20810 (N_20810,N_16222,N_18225);
xor U20811 (N_20811,N_16663,N_16127);
nand U20812 (N_20812,N_18003,N_18162);
nor U20813 (N_20813,N_17133,N_18582);
or U20814 (N_20814,N_16403,N_17551);
nand U20815 (N_20815,N_16933,N_18601);
xor U20816 (N_20816,N_16149,N_18687);
and U20817 (N_20817,N_17333,N_15708);
nand U20818 (N_20818,N_18459,N_18177);
nand U20819 (N_20819,N_16832,N_17681);
nor U20820 (N_20820,N_17881,N_17945);
and U20821 (N_20821,N_16187,N_17926);
nor U20822 (N_20822,N_18199,N_17898);
or U20823 (N_20823,N_16496,N_16848);
and U20824 (N_20824,N_15803,N_18507);
nand U20825 (N_20825,N_17139,N_17875);
nor U20826 (N_20826,N_18502,N_17310);
and U20827 (N_20827,N_18245,N_16066);
and U20828 (N_20828,N_18327,N_18373);
and U20829 (N_20829,N_18162,N_18065);
or U20830 (N_20830,N_18505,N_17514);
and U20831 (N_20831,N_18659,N_16015);
and U20832 (N_20832,N_18209,N_18364);
and U20833 (N_20833,N_17380,N_18151);
nor U20834 (N_20834,N_17576,N_18318);
nor U20835 (N_20835,N_17911,N_16118);
nand U20836 (N_20836,N_17957,N_17228);
or U20837 (N_20837,N_16671,N_17595);
nor U20838 (N_20838,N_16007,N_16833);
or U20839 (N_20839,N_17664,N_17718);
nor U20840 (N_20840,N_16977,N_17332);
and U20841 (N_20841,N_17844,N_16802);
and U20842 (N_20842,N_17774,N_17556);
nor U20843 (N_20843,N_16262,N_15675);
xor U20844 (N_20844,N_17256,N_17291);
nor U20845 (N_20845,N_15960,N_16643);
nor U20846 (N_20846,N_18330,N_17831);
nand U20847 (N_20847,N_17257,N_15848);
and U20848 (N_20848,N_18275,N_18607);
nor U20849 (N_20849,N_17010,N_16044);
nor U20850 (N_20850,N_18423,N_15967);
or U20851 (N_20851,N_16529,N_16311);
nor U20852 (N_20852,N_18147,N_15720);
and U20853 (N_20853,N_15688,N_16383);
nor U20854 (N_20854,N_16292,N_15706);
and U20855 (N_20855,N_17707,N_15865);
nor U20856 (N_20856,N_16123,N_18114);
xnor U20857 (N_20857,N_17938,N_18664);
xnor U20858 (N_20858,N_17046,N_16222);
xnor U20859 (N_20859,N_17176,N_17944);
or U20860 (N_20860,N_18697,N_15972);
nand U20861 (N_20861,N_16021,N_16874);
or U20862 (N_20862,N_16285,N_18178);
nor U20863 (N_20863,N_16240,N_17689);
nand U20864 (N_20864,N_15947,N_15976);
nand U20865 (N_20865,N_15735,N_16952);
nor U20866 (N_20866,N_15821,N_16048);
nor U20867 (N_20867,N_18102,N_15710);
nor U20868 (N_20868,N_18233,N_18423);
nor U20869 (N_20869,N_18237,N_16680);
nor U20870 (N_20870,N_18661,N_16992);
nor U20871 (N_20871,N_18359,N_16302);
xnor U20872 (N_20872,N_15775,N_16810);
and U20873 (N_20873,N_15939,N_18272);
xor U20874 (N_20874,N_17649,N_16329);
nand U20875 (N_20875,N_18174,N_17640);
and U20876 (N_20876,N_17749,N_16575);
nand U20877 (N_20877,N_16022,N_18744);
nand U20878 (N_20878,N_18427,N_18654);
or U20879 (N_20879,N_18538,N_17805);
nand U20880 (N_20880,N_17414,N_16849);
and U20881 (N_20881,N_17801,N_16378);
xnor U20882 (N_20882,N_18096,N_18029);
xnor U20883 (N_20883,N_16137,N_17642);
nor U20884 (N_20884,N_18552,N_17214);
and U20885 (N_20885,N_18574,N_18196);
nor U20886 (N_20886,N_15878,N_18175);
xor U20887 (N_20887,N_18629,N_17722);
or U20888 (N_20888,N_16846,N_16082);
nor U20889 (N_20889,N_18664,N_18304);
nor U20890 (N_20890,N_16492,N_18609);
nand U20891 (N_20891,N_15637,N_16199);
or U20892 (N_20892,N_16934,N_18113);
and U20893 (N_20893,N_16281,N_16368);
and U20894 (N_20894,N_15757,N_18544);
nand U20895 (N_20895,N_17115,N_16581);
or U20896 (N_20896,N_15703,N_17714);
nor U20897 (N_20897,N_17326,N_18622);
xnor U20898 (N_20898,N_18469,N_17806);
nor U20899 (N_20899,N_16827,N_16470);
nor U20900 (N_20900,N_18461,N_18211);
xnor U20901 (N_20901,N_17837,N_17333);
nand U20902 (N_20902,N_17234,N_17500);
nor U20903 (N_20903,N_16186,N_16546);
and U20904 (N_20904,N_16988,N_16667);
and U20905 (N_20905,N_17606,N_15635);
and U20906 (N_20906,N_16527,N_17661);
and U20907 (N_20907,N_16208,N_15832);
nand U20908 (N_20908,N_18627,N_15885);
nor U20909 (N_20909,N_17410,N_16640);
nor U20910 (N_20910,N_17196,N_16205);
or U20911 (N_20911,N_17392,N_16088);
or U20912 (N_20912,N_18375,N_18168);
or U20913 (N_20913,N_17632,N_17885);
and U20914 (N_20914,N_16799,N_16695);
nor U20915 (N_20915,N_16502,N_17933);
nor U20916 (N_20916,N_17763,N_17762);
xor U20917 (N_20917,N_18636,N_15757);
nor U20918 (N_20918,N_18233,N_16222);
and U20919 (N_20919,N_17369,N_16646);
or U20920 (N_20920,N_16201,N_16106);
and U20921 (N_20921,N_18411,N_16897);
or U20922 (N_20922,N_15680,N_18109);
and U20923 (N_20923,N_16697,N_18643);
nand U20924 (N_20924,N_18202,N_17588);
nand U20925 (N_20925,N_17212,N_16226);
and U20926 (N_20926,N_18746,N_16862);
xnor U20927 (N_20927,N_16223,N_17633);
and U20928 (N_20928,N_16046,N_15816);
or U20929 (N_20929,N_18211,N_17237);
or U20930 (N_20930,N_18207,N_16115);
nand U20931 (N_20931,N_15843,N_16452);
or U20932 (N_20932,N_18115,N_16156);
nand U20933 (N_20933,N_16089,N_16248);
or U20934 (N_20934,N_16426,N_16350);
nor U20935 (N_20935,N_17612,N_16405);
and U20936 (N_20936,N_16453,N_18349);
or U20937 (N_20937,N_15886,N_16402);
and U20938 (N_20938,N_16108,N_16704);
or U20939 (N_20939,N_18389,N_17184);
nor U20940 (N_20940,N_16482,N_17741);
nand U20941 (N_20941,N_17873,N_18269);
nand U20942 (N_20942,N_16559,N_18253);
xnor U20943 (N_20943,N_17126,N_15880);
nor U20944 (N_20944,N_15749,N_15929);
nand U20945 (N_20945,N_16546,N_16686);
nand U20946 (N_20946,N_18701,N_16999);
nand U20947 (N_20947,N_17929,N_17934);
and U20948 (N_20948,N_18686,N_15727);
and U20949 (N_20949,N_16769,N_16320);
nand U20950 (N_20950,N_17954,N_16389);
nor U20951 (N_20951,N_17120,N_16254);
or U20952 (N_20952,N_16027,N_18188);
or U20953 (N_20953,N_16413,N_17158);
nor U20954 (N_20954,N_16589,N_16926);
and U20955 (N_20955,N_17944,N_18678);
nand U20956 (N_20956,N_17892,N_18735);
or U20957 (N_20957,N_16894,N_15721);
or U20958 (N_20958,N_17819,N_16622);
or U20959 (N_20959,N_17087,N_16860);
and U20960 (N_20960,N_17861,N_17692);
or U20961 (N_20961,N_15692,N_17676);
nand U20962 (N_20962,N_17457,N_15995);
nor U20963 (N_20963,N_17193,N_16540);
and U20964 (N_20964,N_15757,N_18695);
nand U20965 (N_20965,N_16739,N_18693);
xnor U20966 (N_20966,N_17178,N_16194);
or U20967 (N_20967,N_16894,N_17095);
nor U20968 (N_20968,N_17574,N_18175);
or U20969 (N_20969,N_17257,N_15961);
nand U20970 (N_20970,N_16844,N_17651);
nor U20971 (N_20971,N_17991,N_18081);
nand U20972 (N_20972,N_16856,N_18229);
or U20973 (N_20973,N_16424,N_16921);
and U20974 (N_20974,N_18569,N_15912);
and U20975 (N_20975,N_17229,N_18604);
xor U20976 (N_20976,N_18668,N_16871);
or U20977 (N_20977,N_16517,N_16034);
nand U20978 (N_20978,N_17201,N_16375);
or U20979 (N_20979,N_16251,N_15712);
nand U20980 (N_20980,N_16415,N_16223);
and U20981 (N_20981,N_16388,N_18174);
and U20982 (N_20982,N_17121,N_16486);
nand U20983 (N_20983,N_16286,N_17010);
nor U20984 (N_20984,N_18290,N_17322);
and U20985 (N_20985,N_18057,N_17061);
nand U20986 (N_20986,N_17075,N_18397);
nor U20987 (N_20987,N_17085,N_15975);
nor U20988 (N_20988,N_16223,N_17673);
and U20989 (N_20989,N_16712,N_18457);
or U20990 (N_20990,N_17572,N_16368);
and U20991 (N_20991,N_18308,N_18084);
and U20992 (N_20992,N_15916,N_18295);
nor U20993 (N_20993,N_16607,N_17928);
nor U20994 (N_20994,N_17247,N_17028);
and U20995 (N_20995,N_18472,N_18348);
nor U20996 (N_20996,N_17417,N_16756);
nand U20997 (N_20997,N_15890,N_16901);
nand U20998 (N_20998,N_16953,N_18741);
nand U20999 (N_20999,N_17865,N_18290);
xnor U21000 (N_21000,N_16484,N_16257);
or U21001 (N_21001,N_16355,N_18365);
or U21002 (N_21002,N_17677,N_17796);
and U21003 (N_21003,N_15830,N_16375);
nand U21004 (N_21004,N_18087,N_15932);
nand U21005 (N_21005,N_18612,N_17319);
and U21006 (N_21006,N_15655,N_18427);
or U21007 (N_21007,N_18116,N_18600);
nor U21008 (N_21008,N_16659,N_18460);
nor U21009 (N_21009,N_16468,N_16846);
nand U21010 (N_21010,N_18190,N_16930);
or U21011 (N_21011,N_16502,N_16935);
nand U21012 (N_21012,N_18575,N_18519);
nand U21013 (N_21013,N_15743,N_16590);
nand U21014 (N_21014,N_17209,N_15643);
or U21015 (N_21015,N_18068,N_17351);
nor U21016 (N_21016,N_16206,N_18256);
nor U21017 (N_21017,N_17890,N_16319);
nor U21018 (N_21018,N_15952,N_18440);
or U21019 (N_21019,N_17145,N_16952);
or U21020 (N_21020,N_17322,N_16313);
and U21021 (N_21021,N_16278,N_18550);
nor U21022 (N_21022,N_15740,N_18329);
xnor U21023 (N_21023,N_18188,N_16207);
xnor U21024 (N_21024,N_17378,N_18298);
xnor U21025 (N_21025,N_17818,N_15770);
nand U21026 (N_21026,N_18286,N_16190);
and U21027 (N_21027,N_18038,N_16284);
nand U21028 (N_21028,N_17044,N_15799);
nand U21029 (N_21029,N_17711,N_16895);
and U21030 (N_21030,N_17629,N_18100);
xor U21031 (N_21031,N_17755,N_18002);
nand U21032 (N_21032,N_16531,N_16971);
nand U21033 (N_21033,N_15693,N_18061);
nand U21034 (N_21034,N_16836,N_15856);
nand U21035 (N_21035,N_18245,N_17068);
nand U21036 (N_21036,N_16943,N_17298);
or U21037 (N_21037,N_17371,N_16298);
nor U21038 (N_21038,N_17017,N_18470);
and U21039 (N_21039,N_18302,N_18359);
nor U21040 (N_21040,N_17400,N_17308);
nand U21041 (N_21041,N_15910,N_17986);
or U21042 (N_21042,N_17742,N_17340);
nor U21043 (N_21043,N_18470,N_15766);
and U21044 (N_21044,N_17412,N_18749);
or U21045 (N_21045,N_18640,N_15896);
nor U21046 (N_21046,N_17018,N_17637);
or U21047 (N_21047,N_17520,N_15876);
and U21048 (N_21048,N_16322,N_16355);
and U21049 (N_21049,N_17905,N_18406);
or U21050 (N_21050,N_17302,N_16046);
xnor U21051 (N_21051,N_16908,N_18320);
nand U21052 (N_21052,N_15972,N_17065);
or U21053 (N_21053,N_17671,N_18252);
nand U21054 (N_21054,N_16465,N_16576);
and U21055 (N_21055,N_16954,N_18635);
nor U21056 (N_21056,N_16300,N_17995);
or U21057 (N_21057,N_18498,N_17655);
and U21058 (N_21058,N_16827,N_17129);
or U21059 (N_21059,N_17663,N_17949);
or U21060 (N_21060,N_16610,N_16804);
nand U21061 (N_21061,N_17844,N_15853);
or U21062 (N_21062,N_15723,N_16576);
and U21063 (N_21063,N_16039,N_16916);
or U21064 (N_21064,N_18351,N_16332);
nor U21065 (N_21065,N_17813,N_18216);
xnor U21066 (N_21066,N_17506,N_18390);
xnor U21067 (N_21067,N_16543,N_16991);
and U21068 (N_21068,N_17689,N_15953);
nor U21069 (N_21069,N_16796,N_18495);
nor U21070 (N_21070,N_17055,N_18533);
xnor U21071 (N_21071,N_17853,N_17479);
xor U21072 (N_21072,N_17783,N_16041);
or U21073 (N_21073,N_17613,N_16979);
nor U21074 (N_21074,N_17566,N_18614);
or U21075 (N_21075,N_16707,N_15639);
nand U21076 (N_21076,N_16151,N_15839);
nand U21077 (N_21077,N_16096,N_16901);
nor U21078 (N_21078,N_17677,N_15729);
or U21079 (N_21079,N_16587,N_18414);
or U21080 (N_21080,N_18588,N_16466);
or U21081 (N_21081,N_16367,N_18241);
and U21082 (N_21082,N_18695,N_16296);
and U21083 (N_21083,N_16984,N_18294);
nand U21084 (N_21084,N_16263,N_15845);
and U21085 (N_21085,N_15973,N_18053);
or U21086 (N_21086,N_17102,N_17299);
xnor U21087 (N_21087,N_15700,N_16458);
or U21088 (N_21088,N_17165,N_18263);
and U21089 (N_21089,N_17324,N_18132);
nor U21090 (N_21090,N_18468,N_16910);
nand U21091 (N_21091,N_17168,N_18229);
xnor U21092 (N_21092,N_18182,N_16253);
and U21093 (N_21093,N_16487,N_15988);
and U21094 (N_21094,N_17497,N_16767);
or U21095 (N_21095,N_15959,N_17494);
and U21096 (N_21096,N_16203,N_18342);
nand U21097 (N_21097,N_18148,N_16372);
or U21098 (N_21098,N_17797,N_17750);
or U21099 (N_21099,N_15712,N_17867);
or U21100 (N_21100,N_16852,N_16917);
and U21101 (N_21101,N_18389,N_17657);
nand U21102 (N_21102,N_17908,N_18118);
and U21103 (N_21103,N_16113,N_17836);
or U21104 (N_21104,N_17223,N_17378);
or U21105 (N_21105,N_17923,N_15717);
nor U21106 (N_21106,N_17599,N_17582);
nand U21107 (N_21107,N_16768,N_15839);
nand U21108 (N_21108,N_17808,N_17659);
and U21109 (N_21109,N_17597,N_17805);
nor U21110 (N_21110,N_17356,N_16730);
or U21111 (N_21111,N_15689,N_17553);
nand U21112 (N_21112,N_15719,N_16088);
nor U21113 (N_21113,N_16552,N_17016);
nor U21114 (N_21114,N_16066,N_16467);
nor U21115 (N_21115,N_17750,N_15743);
or U21116 (N_21116,N_17445,N_17614);
and U21117 (N_21117,N_15627,N_16002);
and U21118 (N_21118,N_18086,N_17460);
or U21119 (N_21119,N_17377,N_18422);
or U21120 (N_21120,N_16590,N_16013);
or U21121 (N_21121,N_18122,N_16978);
and U21122 (N_21122,N_16613,N_16989);
or U21123 (N_21123,N_16554,N_17294);
and U21124 (N_21124,N_15736,N_16392);
nand U21125 (N_21125,N_16166,N_18008);
nand U21126 (N_21126,N_17391,N_18002);
nor U21127 (N_21127,N_17964,N_17691);
or U21128 (N_21128,N_16144,N_17240);
or U21129 (N_21129,N_17851,N_15811);
or U21130 (N_21130,N_15780,N_18183);
nor U21131 (N_21131,N_17839,N_16749);
or U21132 (N_21132,N_17539,N_18519);
nand U21133 (N_21133,N_18549,N_17781);
nor U21134 (N_21134,N_17914,N_16187);
and U21135 (N_21135,N_17580,N_16491);
nor U21136 (N_21136,N_17490,N_16789);
nor U21137 (N_21137,N_16347,N_16764);
nand U21138 (N_21138,N_16900,N_17194);
and U21139 (N_21139,N_17468,N_16307);
nand U21140 (N_21140,N_16381,N_16316);
nor U21141 (N_21141,N_17935,N_16787);
and U21142 (N_21142,N_17038,N_18601);
and U21143 (N_21143,N_17213,N_16187);
nor U21144 (N_21144,N_15950,N_15709);
or U21145 (N_21145,N_16386,N_15711);
xor U21146 (N_21146,N_16809,N_16118);
and U21147 (N_21147,N_18738,N_18283);
nand U21148 (N_21148,N_17218,N_17488);
nand U21149 (N_21149,N_16668,N_17586);
nand U21150 (N_21150,N_18620,N_18274);
xnor U21151 (N_21151,N_17556,N_17688);
and U21152 (N_21152,N_18716,N_16558);
or U21153 (N_21153,N_16844,N_16057);
xnor U21154 (N_21154,N_16693,N_18520);
and U21155 (N_21155,N_17459,N_18110);
and U21156 (N_21156,N_17922,N_17424);
xor U21157 (N_21157,N_18231,N_17460);
or U21158 (N_21158,N_18429,N_17243);
nand U21159 (N_21159,N_18659,N_16857);
or U21160 (N_21160,N_17799,N_16565);
and U21161 (N_21161,N_17947,N_17289);
and U21162 (N_21162,N_18215,N_18485);
or U21163 (N_21163,N_17145,N_17413);
or U21164 (N_21164,N_17385,N_17946);
and U21165 (N_21165,N_17023,N_18150);
and U21166 (N_21166,N_16915,N_17809);
or U21167 (N_21167,N_16968,N_17794);
and U21168 (N_21168,N_17139,N_15756);
nand U21169 (N_21169,N_17315,N_15766);
nand U21170 (N_21170,N_16130,N_18229);
or U21171 (N_21171,N_16110,N_16060);
nand U21172 (N_21172,N_18284,N_17276);
and U21173 (N_21173,N_17516,N_15882);
xnor U21174 (N_21174,N_18314,N_18699);
or U21175 (N_21175,N_17672,N_17471);
and U21176 (N_21176,N_16951,N_16689);
nor U21177 (N_21177,N_18117,N_15731);
and U21178 (N_21178,N_16539,N_16631);
xnor U21179 (N_21179,N_17791,N_15660);
nand U21180 (N_21180,N_16049,N_18354);
nand U21181 (N_21181,N_15919,N_18528);
and U21182 (N_21182,N_17495,N_17801);
or U21183 (N_21183,N_16627,N_18300);
or U21184 (N_21184,N_16828,N_18546);
or U21185 (N_21185,N_16657,N_15905);
xor U21186 (N_21186,N_17543,N_16754);
and U21187 (N_21187,N_17684,N_17493);
nor U21188 (N_21188,N_17335,N_16976);
or U21189 (N_21189,N_17177,N_17165);
or U21190 (N_21190,N_16676,N_17327);
nand U21191 (N_21191,N_15874,N_17731);
and U21192 (N_21192,N_18485,N_16800);
nand U21193 (N_21193,N_16651,N_18465);
or U21194 (N_21194,N_16807,N_16261);
nand U21195 (N_21195,N_17285,N_16805);
xor U21196 (N_21196,N_17770,N_17170);
or U21197 (N_21197,N_17004,N_17108);
nor U21198 (N_21198,N_18691,N_18162);
nor U21199 (N_21199,N_16929,N_17262);
nand U21200 (N_21200,N_17535,N_16886);
and U21201 (N_21201,N_16607,N_18177);
nand U21202 (N_21202,N_18451,N_17256);
and U21203 (N_21203,N_17389,N_15627);
nor U21204 (N_21204,N_18710,N_17371);
nand U21205 (N_21205,N_18368,N_18091);
xor U21206 (N_21206,N_17515,N_15901);
xnor U21207 (N_21207,N_16720,N_18497);
xor U21208 (N_21208,N_18620,N_16683);
or U21209 (N_21209,N_18158,N_15626);
or U21210 (N_21210,N_16608,N_18392);
or U21211 (N_21211,N_18616,N_17814);
or U21212 (N_21212,N_16328,N_17519);
nand U21213 (N_21213,N_17351,N_18456);
and U21214 (N_21214,N_16636,N_17713);
xnor U21215 (N_21215,N_17609,N_16007);
nand U21216 (N_21216,N_17758,N_16925);
and U21217 (N_21217,N_15948,N_17844);
or U21218 (N_21218,N_18152,N_17557);
nand U21219 (N_21219,N_16605,N_17827);
nand U21220 (N_21220,N_16929,N_16938);
or U21221 (N_21221,N_18030,N_16457);
nand U21222 (N_21222,N_17803,N_17715);
nand U21223 (N_21223,N_18489,N_18181);
nand U21224 (N_21224,N_17393,N_16814);
and U21225 (N_21225,N_18596,N_18313);
nand U21226 (N_21226,N_16958,N_17920);
nor U21227 (N_21227,N_18578,N_16104);
nand U21228 (N_21228,N_16823,N_16072);
nand U21229 (N_21229,N_15866,N_16436);
or U21230 (N_21230,N_16518,N_18712);
nor U21231 (N_21231,N_15942,N_16385);
nor U21232 (N_21232,N_18725,N_15649);
or U21233 (N_21233,N_16949,N_15749);
and U21234 (N_21234,N_16460,N_16049);
nor U21235 (N_21235,N_18517,N_17831);
and U21236 (N_21236,N_18720,N_16302);
or U21237 (N_21237,N_15725,N_17620);
or U21238 (N_21238,N_16836,N_18736);
nand U21239 (N_21239,N_17702,N_18627);
or U21240 (N_21240,N_15743,N_18267);
nor U21241 (N_21241,N_18060,N_16686);
or U21242 (N_21242,N_17136,N_17221);
nand U21243 (N_21243,N_15845,N_16633);
and U21244 (N_21244,N_18658,N_16067);
nor U21245 (N_21245,N_16751,N_18678);
or U21246 (N_21246,N_15828,N_16101);
xnor U21247 (N_21247,N_16644,N_16707);
nor U21248 (N_21248,N_18255,N_15878);
and U21249 (N_21249,N_16974,N_17099);
nand U21250 (N_21250,N_16083,N_17978);
nor U21251 (N_21251,N_16274,N_18418);
nand U21252 (N_21252,N_16187,N_18069);
or U21253 (N_21253,N_16691,N_17138);
and U21254 (N_21254,N_17009,N_16068);
nand U21255 (N_21255,N_16290,N_15983);
nand U21256 (N_21256,N_17582,N_17041);
or U21257 (N_21257,N_15889,N_17314);
nor U21258 (N_21258,N_17622,N_17694);
or U21259 (N_21259,N_16850,N_17710);
nand U21260 (N_21260,N_17238,N_17762);
nor U21261 (N_21261,N_17197,N_17740);
nand U21262 (N_21262,N_17124,N_16795);
nand U21263 (N_21263,N_17495,N_18140);
nand U21264 (N_21264,N_18268,N_17654);
nand U21265 (N_21265,N_16561,N_18135);
or U21266 (N_21266,N_18147,N_16735);
nand U21267 (N_21267,N_16038,N_15991);
and U21268 (N_21268,N_18308,N_18672);
xnor U21269 (N_21269,N_16232,N_18566);
nand U21270 (N_21270,N_17861,N_17051);
nand U21271 (N_21271,N_18196,N_16354);
xor U21272 (N_21272,N_16718,N_18734);
nand U21273 (N_21273,N_17932,N_16772);
nor U21274 (N_21274,N_17873,N_18082);
nor U21275 (N_21275,N_18675,N_17951);
or U21276 (N_21276,N_17988,N_16085);
nor U21277 (N_21277,N_17635,N_15927);
nor U21278 (N_21278,N_18405,N_16671);
nor U21279 (N_21279,N_16478,N_16215);
or U21280 (N_21280,N_16597,N_18523);
nand U21281 (N_21281,N_17901,N_18342);
or U21282 (N_21282,N_17158,N_17296);
and U21283 (N_21283,N_17276,N_17014);
or U21284 (N_21284,N_17905,N_17988);
nor U21285 (N_21285,N_17321,N_16500);
xor U21286 (N_21286,N_16177,N_15816);
nor U21287 (N_21287,N_18648,N_18617);
or U21288 (N_21288,N_18521,N_16909);
nor U21289 (N_21289,N_16209,N_17091);
or U21290 (N_21290,N_17011,N_17545);
nand U21291 (N_21291,N_17789,N_18385);
and U21292 (N_21292,N_18278,N_17207);
nand U21293 (N_21293,N_16168,N_17828);
or U21294 (N_21294,N_16743,N_17477);
and U21295 (N_21295,N_16063,N_16379);
nor U21296 (N_21296,N_15936,N_17264);
and U21297 (N_21297,N_17734,N_18202);
nor U21298 (N_21298,N_18629,N_17454);
xnor U21299 (N_21299,N_17692,N_17962);
nor U21300 (N_21300,N_16988,N_16684);
and U21301 (N_21301,N_17483,N_16454);
or U21302 (N_21302,N_16105,N_18151);
and U21303 (N_21303,N_17347,N_18369);
or U21304 (N_21304,N_18325,N_18582);
nor U21305 (N_21305,N_18732,N_18049);
nand U21306 (N_21306,N_16800,N_15929);
nor U21307 (N_21307,N_15874,N_17200);
or U21308 (N_21308,N_15957,N_16527);
nand U21309 (N_21309,N_18428,N_18427);
nor U21310 (N_21310,N_16935,N_17616);
nand U21311 (N_21311,N_15740,N_15749);
nor U21312 (N_21312,N_17675,N_17662);
nor U21313 (N_21313,N_18386,N_17790);
and U21314 (N_21314,N_16031,N_15885);
nor U21315 (N_21315,N_16416,N_18677);
nor U21316 (N_21316,N_17906,N_18140);
and U21317 (N_21317,N_16075,N_17169);
nand U21318 (N_21318,N_17147,N_15710);
nor U21319 (N_21319,N_15960,N_18209);
nand U21320 (N_21320,N_17002,N_16299);
and U21321 (N_21321,N_18292,N_17622);
or U21322 (N_21322,N_17690,N_16955);
nor U21323 (N_21323,N_15638,N_17851);
nor U21324 (N_21324,N_16441,N_15987);
and U21325 (N_21325,N_17064,N_16996);
and U21326 (N_21326,N_17211,N_15790);
nand U21327 (N_21327,N_16821,N_15931);
nand U21328 (N_21328,N_17682,N_17967);
and U21329 (N_21329,N_18107,N_18141);
and U21330 (N_21330,N_18354,N_17859);
xor U21331 (N_21331,N_16802,N_15786);
nand U21332 (N_21332,N_16694,N_17473);
or U21333 (N_21333,N_18695,N_17256);
nand U21334 (N_21334,N_18133,N_15993);
and U21335 (N_21335,N_18280,N_17032);
or U21336 (N_21336,N_18524,N_18022);
nand U21337 (N_21337,N_16885,N_18386);
and U21338 (N_21338,N_15845,N_17101);
xnor U21339 (N_21339,N_17128,N_15786);
or U21340 (N_21340,N_16863,N_17118);
nand U21341 (N_21341,N_17252,N_17537);
and U21342 (N_21342,N_15796,N_16473);
nand U21343 (N_21343,N_18668,N_17920);
and U21344 (N_21344,N_17740,N_17241);
nand U21345 (N_21345,N_16363,N_16751);
nor U21346 (N_21346,N_17448,N_18747);
and U21347 (N_21347,N_17038,N_17566);
nor U21348 (N_21348,N_16682,N_16313);
and U21349 (N_21349,N_18278,N_17242);
nand U21350 (N_21350,N_18249,N_18222);
and U21351 (N_21351,N_16035,N_15817);
nor U21352 (N_21352,N_17512,N_16907);
and U21353 (N_21353,N_16342,N_16274);
nor U21354 (N_21354,N_15738,N_18190);
nand U21355 (N_21355,N_17342,N_15971);
or U21356 (N_21356,N_18744,N_16895);
and U21357 (N_21357,N_15858,N_16417);
or U21358 (N_21358,N_15650,N_15693);
nor U21359 (N_21359,N_16474,N_18514);
and U21360 (N_21360,N_17151,N_15702);
and U21361 (N_21361,N_17717,N_18263);
or U21362 (N_21362,N_18128,N_16393);
nor U21363 (N_21363,N_16347,N_18547);
nand U21364 (N_21364,N_18223,N_16873);
or U21365 (N_21365,N_16494,N_16704);
xor U21366 (N_21366,N_17364,N_17844);
and U21367 (N_21367,N_17789,N_17173);
nor U21368 (N_21368,N_17202,N_16859);
or U21369 (N_21369,N_18374,N_17395);
or U21370 (N_21370,N_16687,N_16605);
and U21371 (N_21371,N_18330,N_17789);
or U21372 (N_21372,N_17977,N_18553);
nand U21373 (N_21373,N_16981,N_15718);
or U21374 (N_21374,N_16551,N_18171);
nand U21375 (N_21375,N_18717,N_16080);
and U21376 (N_21376,N_18576,N_15962);
or U21377 (N_21377,N_16770,N_16594);
xnor U21378 (N_21378,N_16562,N_17777);
or U21379 (N_21379,N_18264,N_16163);
xor U21380 (N_21380,N_18403,N_16167);
and U21381 (N_21381,N_17401,N_17500);
xor U21382 (N_21382,N_15941,N_18049);
nor U21383 (N_21383,N_17563,N_18015);
nor U21384 (N_21384,N_16574,N_17057);
nor U21385 (N_21385,N_16976,N_17244);
and U21386 (N_21386,N_16789,N_17302);
xor U21387 (N_21387,N_18749,N_15864);
nor U21388 (N_21388,N_15702,N_17693);
nand U21389 (N_21389,N_16998,N_18101);
or U21390 (N_21390,N_16567,N_18018);
and U21391 (N_21391,N_17467,N_17217);
nor U21392 (N_21392,N_15661,N_16552);
or U21393 (N_21393,N_18091,N_17707);
and U21394 (N_21394,N_16002,N_16867);
or U21395 (N_21395,N_17659,N_16367);
or U21396 (N_21396,N_17125,N_15936);
and U21397 (N_21397,N_18208,N_17192);
and U21398 (N_21398,N_18577,N_15690);
nand U21399 (N_21399,N_16912,N_16047);
and U21400 (N_21400,N_16713,N_18217);
nand U21401 (N_21401,N_18608,N_16035);
nor U21402 (N_21402,N_17738,N_16004);
or U21403 (N_21403,N_16126,N_16866);
or U21404 (N_21404,N_16949,N_16682);
and U21405 (N_21405,N_16638,N_16603);
nor U21406 (N_21406,N_18496,N_16027);
nand U21407 (N_21407,N_15841,N_15774);
xnor U21408 (N_21408,N_16654,N_18043);
nor U21409 (N_21409,N_16358,N_16306);
and U21410 (N_21410,N_16482,N_17843);
nor U21411 (N_21411,N_18520,N_15661);
or U21412 (N_21412,N_16050,N_16037);
nor U21413 (N_21413,N_17955,N_16486);
or U21414 (N_21414,N_16535,N_15636);
or U21415 (N_21415,N_16864,N_16624);
and U21416 (N_21416,N_17638,N_18306);
nor U21417 (N_21417,N_16347,N_17312);
or U21418 (N_21418,N_16977,N_17287);
nor U21419 (N_21419,N_16731,N_17872);
or U21420 (N_21420,N_18328,N_18333);
xor U21421 (N_21421,N_16656,N_17612);
and U21422 (N_21422,N_17587,N_17479);
nand U21423 (N_21423,N_16012,N_17373);
nor U21424 (N_21424,N_17020,N_17621);
or U21425 (N_21425,N_18110,N_18145);
and U21426 (N_21426,N_16923,N_18528);
nor U21427 (N_21427,N_18446,N_17547);
nor U21428 (N_21428,N_16600,N_17051);
and U21429 (N_21429,N_17612,N_16811);
or U21430 (N_21430,N_16050,N_15945);
and U21431 (N_21431,N_15659,N_17311);
nor U21432 (N_21432,N_16063,N_16306);
nor U21433 (N_21433,N_16613,N_18455);
or U21434 (N_21434,N_16325,N_18181);
nor U21435 (N_21435,N_17730,N_16844);
nor U21436 (N_21436,N_16113,N_16654);
or U21437 (N_21437,N_15951,N_17972);
or U21438 (N_21438,N_16919,N_17526);
or U21439 (N_21439,N_15819,N_18265);
or U21440 (N_21440,N_18180,N_16996);
nor U21441 (N_21441,N_16285,N_16655);
nand U21442 (N_21442,N_18552,N_16070);
nand U21443 (N_21443,N_18118,N_16718);
nand U21444 (N_21444,N_18653,N_17069);
nor U21445 (N_21445,N_16481,N_17901);
nand U21446 (N_21446,N_16077,N_15631);
and U21447 (N_21447,N_15792,N_15748);
nor U21448 (N_21448,N_17098,N_17862);
nor U21449 (N_21449,N_17104,N_17527);
or U21450 (N_21450,N_16251,N_18437);
nor U21451 (N_21451,N_15935,N_17755);
and U21452 (N_21452,N_17985,N_17174);
and U21453 (N_21453,N_17989,N_15939);
nand U21454 (N_21454,N_16243,N_17264);
xnor U21455 (N_21455,N_18479,N_16448);
nor U21456 (N_21456,N_18218,N_17473);
nor U21457 (N_21457,N_16165,N_17754);
nand U21458 (N_21458,N_17816,N_18713);
nor U21459 (N_21459,N_17136,N_18650);
nor U21460 (N_21460,N_16270,N_15764);
or U21461 (N_21461,N_18157,N_17620);
nor U21462 (N_21462,N_16413,N_16671);
or U21463 (N_21463,N_15903,N_18694);
and U21464 (N_21464,N_18419,N_16524);
xnor U21465 (N_21465,N_17313,N_17345);
nor U21466 (N_21466,N_16145,N_17929);
nor U21467 (N_21467,N_17697,N_18605);
nand U21468 (N_21468,N_17248,N_17592);
and U21469 (N_21469,N_16286,N_15814);
or U21470 (N_21470,N_16948,N_18047);
or U21471 (N_21471,N_18361,N_15792);
nor U21472 (N_21472,N_18391,N_16969);
or U21473 (N_21473,N_16096,N_16447);
nand U21474 (N_21474,N_17752,N_16053);
nor U21475 (N_21475,N_16801,N_16263);
and U21476 (N_21476,N_16100,N_16005);
and U21477 (N_21477,N_16303,N_18317);
and U21478 (N_21478,N_17788,N_18043);
nand U21479 (N_21479,N_18679,N_17503);
and U21480 (N_21480,N_17136,N_18524);
xor U21481 (N_21481,N_17768,N_16976);
nand U21482 (N_21482,N_18736,N_18101);
and U21483 (N_21483,N_17022,N_17699);
nand U21484 (N_21484,N_17628,N_17572);
nor U21485 (N_21485,N_16742,N_16276);
nand U21486 (N_21486,N_18550,N_15698);
or U21487 (N_21487,N_16118,N_17753);
nand U21488 (N_21488,N_17650,N_17969);
nor U21489 (N_21489,N_18268,N_16267);
nor U21490 (N_21490,N_17624,N_16801);
nand U21491 (N_21491,N_15719,N_16430);
nor U21492 (N_21492,N_18023,N_15715);
xor U21493 (N_21493,N_16865,N_16130);
nand U21494 (N_21494,N_17661,N_17156);
or U21495 (N_21495,N_17695,N_15812);
nor U21496 (N_21496,N_15825,N_18329);
and U21497 (N_21497,N_16388,N_16888);
nand U21498 (N_21498,N_18571,N_16421);
nor U21499 (N_21499,N_16019,N_16472);
nand U21500 (N_21500,N_15949,N_16899);
nand U21501 (N_21501,N_18241,N_16134);
xnor U21502 (N_21502,N_18696,N_18479);
or U21503 (N_21503,N_15846,N_17299);
nand U21504 (N_21504,N_17515,N_16726);
or U21505 (N_21505,N_17277,N_18293);
or U21506 (N_21506,N_17084,N_15678);
or U21507 (N_21507,N_18255,N_16194);
xor U21508 (N_21508,N_17236,N_15945);
nand U21509 (N_21509,N_18075,N_15685);
or U21510 (N_21510,N_17789,N_16257);
nor U21511 (N_21511,N_16117,N_17101);
or U21512 (N_21512,N_16039,N_18685);
nand U21513 (N_21513,N_15680,N_16018);
xor U21514 (N_21514,N_16837,N_17970);
nor U21515 (N_21515,N_16773,N_17890);
nor U21516 (N_21516,N_16849,N_16288);
nand U21517 (N_21517,N_17183,N_17910);
xnor U21518 (N_21518,N_18005,N_16404);
nand U21519 (N_21519,N_16548,N_17997);
or U21520 (N_21520,N_16145,N_17860);
nand U21521 (N_21521,N_18088,N_18121);
nand U21522 (N_21522,N_18672,N_18749);
and U21523 (N_21523,N_18174,N_17899);
and U21524 (N_21524,N_16511,N_16689);
nor U21525 (N_21525,N_17084,N_16902);
or U21526 (N_21526,N_18255,N_15842);
nand U21527 (N_21527,N_16095,N_18421);
xnor U21528 (N_21528,N_18439,N_16947);
nand U21529 (N_21529,N_17333,N_18728);
nor U21530 (N_21530,N_16571,N_17764);
and U21531 (N_21531,N_15686,N_16052);
or U21532 (N_21532,N_17945,N_16459);
and U21533 (N_21533,N_17326,N_18412);
and U21534 (N_21534,N_17053,N_18686);
and U21535 (N_21535,N_17109,N_18286);
nand U21536 (N_21536,N_17953,N_18631);
or U21537 (N_21537,N_16346,N_18245);
and U21538 (N_21538,N_18132,N_17291);
or U21539 (N_21539,N_18704,N_16998);
or U21540 (N_21540,N_18618,N_16440);
nor U21541 (N_21541,N_17970,N_16681);
nand U21542 (N_21542,N_16106,N_17088);
nor U21543 (N_21543,N_17310,N_17493);
and U21544 (N_21544,N_18608,N_17561);
or U21545 (N_21545,N_15873,N_16547);
or U21546 (N_21546,N_16237,N_15741);
nor U21547 (N_21547,N_17976,N_16215);
or U21548 (N_21548,N_18632,N_18183);
nor U21549 (N_21549,N_18715,N_18556);
nand U21550 (N_21550,N_18298,N_15890);
and U21551 (N_21551,N_17904,N_16632);
nand U21552 (N_21552,N_18413,N_18616);
or U21553 (N_21553,N_15664,N_15627);
and U21554 (N_21554,N_18414,N_17500);
nand U21555 (N_21555,N_17452,N_17263);
or U21556 (N_21556,N_18294,N_18325);
nand U21557 (N_21557,N_18452,N_16992);
nand U21558 (N_21558,N_18624,N_17158);
and U21559 (N_21559,N_17212,N_17140);
nand U21560 (N_21560,N_16521,N_17706);
nor U21561 (N_21561,N_16327,N_16133);
nand U21562 (N_21562,N_16669,N_18726);
and U21563 (N_21563,N_17812,N_16121);
nand U21564 (N_21564,N_16441,N_16730);
or U21565 (N_21565,N_17359,N_18051);
nand U21566 (N_21566,N_18721,N_18071);
and U21567 (N_21567,N_18641,N_18156);
nor U21568 (N_21568,N_17836,N_17004);
nor U21569 (N_21569,N_16880,N_18182);
or U21570 (N_21570,N_16597,N_17686);
nor U21571 (N_21571,N_17421,N_16381);
nor U21572 (N_21572,N_15921,N_18079);
and U21573 (N_21573,N_17324,N_16104);
or U21574 (N_21574,N_17107,N_17067);
nor U21575 (N_21575,N_17992,N_16943);
or U21576 (N_21576,N_15933,N_18118);
and U21577 (N_21577,N_16782,N_18202);
and U21578 (N_21578,N_15696,N_18182);
nor U21579 (N_21579,N_18438,N_18587);
or U21580 (N_21580,N_17258,N_15906);
and U21581 (N_21581,N_17331,N_16145);
nand U21582 (N_21582,N_16034,N_15727);
nand U21583 (N_21583,N_18253,N_18374);
and U21584 (N_21584,N_17909,N_17222);
or U21585 (N_21585,N_17881,N_15680);
xor U21586 (N_21586,N_18163,N_16702);
and U21587 (N_21587,N_17101,N_17866);
nand U21588 (N_21588,N_18272,N_17264);
nor U21589 (N_21589,N_16515,N_16471);
or U21590 (N_21590,N_15782,N_16734);
nor U21591 (N_21591,N_17047,N_16170);
nor U21592 (N_21592,N_16313,N_17681);
nor U21593 (N_21593,N_17514,N_16428);
nand U21594 (N_21594,N_16228,N_16769);
and U21595 (N_21595,N_17935,N_18041);
or U21596 (N_21596,N_16938,N_16109);
or U21597 (N_21597,N_16324,N_17439);
nand U21598 (N_21598,N_16425,N_18107);
and U21599 (N_21599,N_17044,N_16589);
xnor U21600 (N_21600,N_18515,N_18042);
and U21601 (N_21601,N_18403,N_17174);
and U21602 (N_21602,N_15866,N_17467);
and U21603 (N_21603,N_17496,N_18632);
nor U21604 (N_21604,N_16437,N_16578);
nand U21605 (N_21605,N_17855,N_17049);
xnor U21606 (N_21606,N_15960,N_16942);
and U21607 (N_21607,N_17037,N_17694);
and U21608 (N_21608,N_15749,N_16967);
and U21609 (N_21609,N_17383,N_16067);
xor U21610 (N_21610,N_16193,N_15784);
or U21611 (N_21611,N_18560,N_16019);
or U21612 (N_21612,N_16786,N_17276);
nand U21613 (N_21613,N_16664,N_15781);
and U21614 (N_21614,N_17563,N_16288);
or U21615 (N_21615,N_18421,N_17018);
nor U21616 (N_21616,N_16409,N_18190);
nand U21617 (N_21617,N_18662,N_15845);
nand U21618 (N_21618,N_17529,N_16913);
and U21619 (N_21619,N_16212,N_16275);
nand U21620 (N_21620,N_16620,N_16150);
nor U21621 (N_21621,N_18703,N_15947);
xor U21622 (N_21622,N_15895,N_16110);
and U21623 (N_21623,N_18416,N_16705);
and U21624 (N_21624,N_18475,N_16113);
nand U21625 (N_21625,N_16081,N_16919);
nor U21626 (N_21626,N_16950,N_15955);
or U21627 (N_21627,N_16880,N_16059);
nand U21628 (N_21628,N_17754,N_18210);
and U21629 (N_21629,N_18470,N_16836);
nor U21630 (N_21630,N_16801,N_15672);
or U21631 (N_21631,N_17209,N_15980);
and U21632 (N_21632,N_15693,N_17811);
nand U21633 (N_21633,N_17614,N_17876);
and U21634 (N_21634,N_17761,N_17477);
and U21635 (N_21635,N_16673,N_16528);
or U21636 (N_21636,N_15817,N_17300);
or U21637 (N_21637,N_16697,N_18479);
xnor U21638 (N_21638,N_18177,N_17364);
and U21639 (N_21639,N_17697,N_18369);
and U21640 (N_21640,N_18482,N_18032);
nand U21641 (N_21641,N_16508,N_17818);
nor U21642 (N_21642,N_16551,N_16408);
xor U21643 (N_21643,N_16724,N_18687);
nor U21644 (N_21644,N_15861,N_15669);
and U21645 (N_21645,N_16982,N_18628);
or U21646 (N_21646,N_16740,N_18494);
nor U21647 (N_21647,N_16134,N_17504);
nor U21648 (N_21648,N_17016,N_16615);
xor U21649 (N_21649,N_18605,N_17870);
nor U21650 (N_21650,N_17812,N_16189);
and U21651 (N_21651,N_17106,N_18425);
or U21652 (N_21652,N_18539,N_16629);
or U21653 (N_21653,N_18295,N_17256);
nor U21654 (N_21654,N_18337,N_17724);
or U21655 (N_21655,N_15782,N_17701);
nand U21656 (N_21656,N_18246,N_18394);
xor U21657 (N_21657,N_18739,N_17229);
xor U21658 (N_21658,N_16596,N_16546);
or U21659 (N_21659,N_17504,N_17602);
or U21660 (N_21660,N_18257,N_16366);
or U21661 (N_21661,N_18432,N_15761);
nand U21662 (N_21662,N_16116,N_16805);
nor U21663 (N_21663,N_18072,N_18317);
or U21664 (N_21664,N_17421,N_18589);
nand U21665 (N_21665,N_16662,N_17122);
or U21666 (N_21666,N_16346,N_16248);
nand U21667 (N_21667,N_16420,N_17219);
nor U21668 (N_21668,N_17668,N_16622);
and U21669 (N_21669,N_16899,N_17399);
nand U21670 (N_21670,N_16595,N_15896);
nand U21671 (N_21671,N_18065,N_16051);
nor U21672 (N_21672,N_15919,N_16863);
or U21673 (N_21673,N_16185,N_18413);
and U21674 (N_21674,N_16723,N_17559);
and U21675 (N_21675,N_17268,N_16623);
nor U21676 (N_21676,N_15876,N_17008);
and U21677 (N_21677,N_18576,N_15989);
or U21678 (N_21678,N_15794,N_16855);
and U21679 (N_21679,N_15662,N_16550);
and U21680 (N_21680,N_16178,N_16103);
nand U21681 (N_21681,N_15801,N_16263);
or U21682 (N_21682,N_18267,N_17107);
nand U21683 (N_21683,N_18707,N_16527);
nor U21684 (N_21684,N_16664,N_17723);
nor U21685 (N_21685,N_17435,N_18475);
nor U21686 (N_21686,N_16134,N_16733);
or U21687 (N_21687,N_16519,N_15914);
nand U21688 (N_21688,N_16513,N_17491);
nor U21689 (N_21689,N_18615,N_18243);
nor U21690 (N_21690,N_16310,N_17183);
or U21691 (N_21691,N_17286,N_16436);
nor U21692 (N_21692,N_17506,N_15963);
nand U21693 (N_21693,N_18495,N_17291);
or U21694 (N_21694,N_17670,N_17431);
and U21695 (N_21695,N_16969,N_17192);
nor U21696 (N_21696,N_18473,N_16477);
and U21697 (N_21697,N_15797,N_16071);
nand U21698 (N_21698,N_18063,N_18592);
and U21699 (N_21699,N_17538,N_16478);
nor U21700 (N_21700,N_16618,N_15627);
nand U21701 (N_21701,N_17640,N_16808);
nor U21702 (N_21702,N_17422,N_16143);
xnor U21703 (N_21703,N_16099,N_18563);
and U21704 (N_21704,N_18688,N_16847);
nor U21705 (N_21705,N_17522,N_16733);
xor U21706 (N_21706,N_17617,N_18505);
or U21707 (N_21707,N_16230,N_16794);
or U21708 (N_21708,N_16915,N_18743);
nor U21709 (N_21709,N_17954,N_16068);
and U21710 (N_21710,N_16151,N_16088);
and U21711 (N_21711,N_16939,N_15833);
xnor U21712 (N_21712,N_17273,N_17042);
or U21713 (N_21713,N_16252,N_18675);
and U21714 (N_21714,N_18441,N_18345);
and U21715 (N_21715,N_18556,N_18032);
or U21716 (N_21716,N_17637,N_17034);
xnor U21717 (N_21717,N_17316,N_18496);
or U21718 (N_21718,N_16082,N_15891);
nand U21719 (N_21719,N_16978,N_18123);
and U21720 (N_21720,N_16235,N_16849);
nor U21721 (N_21721,N_17250,N_18414);
nand U21722 (N_21722,N_17792,N_16229);
and U21723 (N_21723,N_15952,N_17536);
nand U21724 (N_21724,N_17876,N_17279);
nand U21725 (N_21725,N_17630,N_18425);
nor U21726 (N_21726,N_16530,N_15686);
and U21727 (N_21727,N_16693,N_18235);
and U21728 (N_21728,N_16424,N_18646);
or U21729 (N_21729,N_16056,N_16838);
nor U21730 (N_21730,N_18163,N_17873);
nand U21731 (N_21731,N_17624,N_18661);
nor U21732 (N_21732,N_17904,N_17301);
xor U21733 (N_21733,N_16330,N_17140);
xor U21734 (N_21734,N_16776,N_18248);
nor U21735 (N_21735,N_15690,N_18141);
or U21736 (N_21736,N_18290,N_17131);
nor U21737 (N_21737,N_16873,N_18490);
and U21738 (N_21738,N_16227,N_18232);
nand U21739 (N_21739,N_18616,N_17732);
and U21740 (N_21740,N_15662,N_17247);
nand U21741 (N_21741,N_17157,N_16996);
xnor U21742 (N_21742,N_16075,N_16870);
or U21743 (N_21743,N_17774,N_17156);
nor U21744 (N_21744,N_15678,N_18351);
nor U21745 (N_21745,N_16631,N_17969);
nor U21746 (N_21746,N_18651,N_18601);
nand U21747 (N_21747,N_16159,N_16172);
nand U21748 (N_21748,N_18397,N_17813);
and U21749 (N_21749,N_17352,N_17612);
or U21750 (N_21750,N_17593,N_16552);
xor U21751 (N_21751,N_16952,N_18599);
xor U21752 (N_21752,N_17526,N_18562);
and U21753 (N_21753,N_17756,N_16761);
or U21754 (N_21754,N_18222,N_18386);
nand U21755 (N_21755,N_17049,N_16900);
nor U21756 (N_21756,N_16596,N_16295);
and U21757 (N_21757,N_16818,N_16544);
or U21758 (N_21758,N_18275,N_17030);
and U21759 (N_21759,N_17658,N_15890);
xnor U21760 (N_21760,N_18122,N_16182);
or U21761 (N_21761,N_15754,N_15848);
and U21762 (N_21762,N_16778,N_17169);
nor U21763 (N_21763,N_16344,N_15950);
nor U21764 (N_21764,N_17567,N_16352);
nand U21765 (N_21765,N_17716,N_18552);
and U21766 (N_21766,N_17138,N_17747);
nor U21767 (N_21767,N_18304,N_18677);
xor U21768 (N_21768,N_18432,N_17721);
or U21769 (N_21769,N_15996,N_17083);
and U21770 (N_21770,N_16406,N_18740);
and U21771 (N_21771,N_16725,N_18330);
nor U21772 (N_21772,N_16911,N_15829);
xor U21773 (N_21773,N_16183,N_17409);
and U21774 (N_21774,N_18714,N_16924);
or U21775 (N_21775,N_18352,N_16382);
nor U21776 (N_21776,N_17432,N_17781);
xor U21777 (N_21777,N_16829,N_18042);
or U21778 (N_21778,N_18305,N_18419);
or U21779 (N_21779,N_18315,N_18500);
and U21780 (N_21780,N_15681,N_18353);
or U21781 (N_21781,N_15898,N_16774);
nand U21782 (N_21782,N_16834,N_18485);
xnor U21783 (N_21783,N_17274,N_16759);
and U21784 (N_21784,N_16932,N_17453);
and U21785 (N_21785,N_17950,N_17486);
nand U21786 (N_21786,N_17035,N_18184);
or U21787 (N_21787,N_17229,N_16885);
xnor U21788 (N_21788,N_16339,N_18290);
nand U21789 (N_21789,N_17507,N_18270);
and U21790 (N_21790,N_17990,N_15634);
or U21791 (N_21791,N_16171,N_15925);
and U21792 (N_21792,N_17843,N_17223);
or U21793 (N_21793,N_17495,N_15627);
or U21794 (N_21794,N_16258,N_17130);
nand U21795 (N_21795,N_15815,N_16753);
and U21796 (N_21796,N_17264,N_17248);
nor U21797 (N_21797,N_17397,N_16549);
and U21798 (N_21798,N_18405,N_17373);
xnor U21799 (N_21799,N_16293,N_18692);
or U21800 (N_21800,N_16360,N_17500);
or U21801 (N_21801,N_18728,N_16422);
and U21802 (N_21802,N_16843,N_18442);
and U21803 (N_21803,N_17541,N_18722);
or U21804 (N_21804,N_17549,N_17430);
and U21805 (N_21805,N_16511,N_18373);
nor U21806 (N_21806,N_17662,N_16249);
or U21807 (N_21807,N_17747,N_17650);
or U21808 (N_21808,N_18692,N_16617);
nand U21809 (N_21809,N_18386,N_17974);
nand U21810 (N_21810,N_16814,N_16876);
nand U21811 (N_21811,N_16698,N_16779);
xnor U21812 (N_21812,N_17483,N_17145);
nand U21813 (N_21813,N_17725,N_15744);
nor U21814 (N_21814,N_18022,N_16165);
nand U21815 (N_21815,N_17228,N_15883);
or U21816 (N_21816,N_18286,N_16779);
nor U21817 (N_21817,N_17712,N_16841);
nand U21818 (N_21818,N_15881,N_17138);
nor U21819 (N_21819,N_17806,N_18375);
nand U21820 (N_21820,N_16859,N_15805);
or U21821 (N_21821,N_15669,N_15807);
or U21822 (N_21822,N_18573,N_16202);
nor U21823 (N_21823,N_16498,N_18331);
and U21824 (N_21824,N_15810,N_17145);
nor U21825 (N_21825,N_16362,N_16454);
and U21826 (N_21826,N_16596,N_18254);
nand U21827 (N_21827,N_18190,N_17943);
and U21828 (N_21828,N_17455,N_18254);
nor U21829 (N_21829,N_16533,N_17964);
and U21830 (N_21830,N_18354,N_17851);
and U21831 (N_21831,N_16314,N_18590);
or U21832 (N_21832,N_16614,N_17155);
xnor U21833 (N_21833,N_17248,N_15724);
and U21834 (N_21834,N_18545,N_18151);
nor U21835 (N_21835,N_17514,N_18547);
nand U21836 (N_21836,N_17793,N_16718);
nor U21837 (N_21837,N_15861,N_16404);
and U21838 (N_21838,N_17695,N_18024);
nor U21839 (N_21839,N_15670,N_18506);
nor U21840 (N_21840,N_15759,N_17266);
and U21841 (N_21841,N_17207,N_18730);
or U21842 (N_21842,N_18741,N_17000);
nand U21843 (N_21843,N_16363,N_17193);
nor U21844 (N_21844,N_17362,N_15656);
nand U21845 (N_21845,N_15770,N_18070);
or U21846 (N_21846,N_15836,N_17897);
xor U21847 (N_21847,N_15744,N_16946);
and U21848 (N_21848,N_16359,N_18054);
nand U21849 (N_21849,N_18510,N_16548);
and U21850 (N_21850,N_16893,N_18188);
nor U21851 (N_21851,N_16169,N_17329);
and U21852 (N_21852,N_16595,N_16857);
xor U21853 (N_21853,N_16672,N_17545);
nor U21854 (N_21854,N_15776,N_16138);
or U21855 (N_21855,N_16977,N_18574);
and U21856 (N_21856,N_17935,N_15641);
nand U21857 (N_21857,N_16454,N_18009);
nand U21858 (N_21858,N_17335,N_17549);
or U21859 (N_21859,N_16103,N_17065);
nand U21860 (N_21860,N_16152,N_16052);
nand U21861 (N_21861,N_15766,N_15980);
or U21862 (N_21862,N_16938,N_18137);
nand U21863 (N_21863,N_16471,N_18191);
or U21864 (N_21864,N_16120,N_16804);
xnor U21865 (N_21865,N_16760,N_16928);
and U21866 (N_21866,N_18528,N_15874);
and U21867 (N_21867,N_16568,N_15791);
nand U21868 (N_21868,N_17701,N_16936);
or U21869 (N_21869,N_17488,N_15739);
or U21870 (N_21870,N_18525,N_15783);
or U21871 (N_21871,N_17707,N_17118);
and U21872 (N_21872,N_17034,N_16734);
or U21873 (N_21873,N_16537,N_17393);
and U21874 (N_21874,N_18205,N_18611);
or U21875 (N_21875,N_19385,N_20461);
nor U21876 (N_21876,N_18905,N_19977);
nor U21877 (N_21877,N_19414,N_21611);
nand U21878 (N_21878,N_21379,N_20096);
or U21879 (N_21879,N_19506,N_20433);
and U21880 (N_21880,N_20390,N_20725);
nor U21881 (N_21881,N_20247,N_20653);
and U21882 (N_21882,N_20799,N_21720);
xnor U21883 (N_21883,N_19469,N_20153);
nand U21884 (N_21884,N_21800,N_20526);
or U21885 (N_21885,N_21524,N_19846);
and U21886 (N_21886,N_21075,N_21277);
and U21887 (N_21887,N_20746,N_19554);
and U21888 (N_21888,N_21713,N_19794);
and U21889 (N_21889,N_21325,N_20307);
nand U21890 (N_21890,N_21013,N_20661);
and U21891 (N_21891,N_20850,N_21257);
or U21892 (N_21892,N_21061,N_19729);
or U21893 (N_21893,N_20720,N_21512);
and U21894 (N_21894,N_20992,N_21862);
nor U21895 (N_21895,N_21266,N_19395);
and U21896 (N_21896,N_21667,N_19911);
xnor U21897 (N_21897,N_19586,N_20624);
xnor U21898 (N_21898,N_21248,N_19797);
nand U21899 (N_21899,N_19090,N_20860);
or U21900 (N_21900,N_21843,N_21399);
or U21901 (N_21901,N_21112,N_19152);
and U21902 (N_21902,N_19838,N_19324);
nor U21903 (N_21903,N_21766,N_19015);
nor U21904 (N_21904,N_21556,N_21105);
or U21905 (N_21905,N_20928,N_19275);
nor U21906 (N_21906,N_20454,N_20453);
or U21907 (N_21907,N_19102,N_18967);
xnor U21908 (N_21908,N_20508,N_20649);
nand U21909 (N_21909,N_21641,N_20132);
nor U21910 (N_21910,N_19572,N_19644);
xnor U21911 (N_21911,N_21805,N_19675);
xnor U21912 (N_21912,N_20470,N_20417);
nor U21913 (N_21913,N_21161,N_19227);
and U21914 (N_21914,N_21673,N_19159);
or U21915 (N_21915,N_20945,N_21133);
and U21916 (N_21916,N_20870,N_19773);
nor U21917 (N_21917,N_20736,N_19202);
nor U21918 (N_21918,N_19490,N_19235);
or U21919 (N_21919,N_20848,N_19335);
nand U21920 (N_21920,N_20152,N_20608);
nand U21921 (N_21921,N_19585,N_19634);
nand U21922 (N_21922,N_19072,N_21077);
or U21923 (N_21923,N_20305,N_20030);
nand U21924 (N_21924,N_19618,N_19825);
nand U21925 (N_21925,N_19183,N_20936);
nand U21926 (N_21926,N_19296,N_21488);
and U21927 (N_21927,N_21559,N_21165);
nor U21928 (N_21928,N_19927,N_19390);
or U21929 (N_21929,N_20200,N_21218);
and U21930 (N_21930,N_19428,N_19824);
nor U21931 (N_21931,N_20116,N_20335);
nand U21932 (N_21932,N_20236,N_20790);
and U21933 (N_21933,N_20239,N_19532);
or U21934 (N_21934,N_20756,N_20830);
and U21935 (N_21935,N_20772,N_19473);
nor U21936 (N_21936,N_18805,N_20405);
xnor U21937 (N_21937,N_21770,N_20513);
nor U21938 (N_21938,N_21267,N_21371);
nor U21939 (N_21939,N_21547,N_20209);
nand U21940 (N_21940,N_20856,N_19737);
and U21941 (N_21941,N_19745,N_19289);
nor U21942 (N_21942,N_19454,N_18800);
nand U21943 (N_21943,N_18788,N_19643);
or U21944 (N_21944,N_20668,N_21265);
and U21945 (N_21945,N_19806,N_21116);
and U21946 (N_21946,N_19213,N_20241);
or U21947 (N_21947,N_19693,N_20806);
nand U21948 (N_21948,N_18822,N_19795);
or U21949 (N_21949,N_19995,N_19859);
nand U21950 (N_21950,N_21059,N_20038);
nand U21951 (N_21951,N_19487,N_21478);
or U21952 (N_21952,N_18773,N_21600);
or U21953 (N_21953,N_20586,N_20706);
xor U21954 (N_21954,N_19187,N_19182);
xnor U21955 (N_21955,N_20766,N_21605);
or U21956 (N_21956,N_19312,N_21167);
and U21957 (N_21957,N_19852,N_20399);
nand U21958 (N_21958,N_19816,N_19493);
and U21959 (N_21959,N_19242,N_20011);
xnor U21960 (N_21960,N_21226,N_20352);
or U21961 (N_21961,N_19793,N_21416);
nor U21962 (N_21962,N_20383,N_20646);
or U21963 (N_21963,N_19201,N_19430);
nor U21964 (N_21964,N_19880,N_19548);
and U21965 (N_21965,N_19214,N_19136);
nand U21966 (N_21966,N_18863,N_21384);
nand U21967 (N_21967,N_20047,N_18772);
or U21968 (N_21968,N_20373,N_21534);
or U21969 (N_21969,N_19318,N_20425);
nand U21970 (N_21970,N_21444,N_20398);
nand U21971 (N_21971,N_18993,N_19547);
nand U21972 (N_21972,N_20917,N_19319);
and U21973 (N_21973,N_19457,N_20146);
or U21974 (N_21974,N_21767,N_20963);
xnor U21975 (N_21975,N_21376,N_19885);
nor U21976 (N_21976,N_21680,N_21617);
nor U21977 (N_21977,N_20252,N_19293);
xor U21978 (N_21978,N_21561,N_20622);
and U21979 (N_21979,N_20026,N_19582);
or U21980 (N_21980,N_21250,N_21782);
nor U21981 (N_21981,N_20544,N_19221);
nand U21982 (N_21982,N_19328,N_21708);
nor U21983 (N_21983,N_20444,N_19360);
nand U21984 (N_21984,N_19789,N_20426);
and U21985 (N_21985,N_19787,N_20217);
and U21986 (N_21986,N_20292,N_19144);
and U21987 (N_21987,N_19354,N_21836);
and U21988 (N_21988,N_21391,N_20017);
nor U21989 (N_21989,N_19987,N_20862);
or U21990 (N_21990,N_19934,N_21866);
or U21991 (N_21991,N_19650,N_18938);
or U21992 (N_21992,N_19524,N_20614);
nand U21993 (N_21993,N_21507,N_20561);
nor U21994 (N_21994,N_20696,N_19892);
or U21995 (N_21995,N_21586,N_20016);
nor U21996 (N_21996,N_20286,N_20476);
nand U21997 (N_21997,N_19241,N_18831);
or U21998 (N_21998,N_20602,N_20967);
nor U21999 (N_21999,N_21402,N_20609);
nor U22000 (N_22000,N_20881,N_20818);
and U22001 (N_22001,N_19006,N_18755);
and U22002 (N_22002,N_19406,N_21317);
nor U22003 (N_22003,N_19267,N_20697);
and U22004 (N_22004,N_20601,N_21249);
and U22005 (N_22005,N_19263,N_21633);
nor U22006 (N_22006,N_18991,N_21349);
nor U22007 (N_22007,N_21432,N_20548);
or U22008 (N_22008,N_21870,N_21580);
and U22009 (N_22009,N_19302,N_19649);
or U22010 (N_22010,N_21850,N_20483);
nor U22011 (N_22011,N_21184,N_20698);
nand U22012 (N_22012,N_20741,N_19879);
xor U22013 (N_22013,N_19416,N_20838);
and U22014 (N_22014,N_20313,N_20515);
or U22015 (N_22015,N_19606,N_19191);
or U22016 (N_22016,N_21276,N_19812);
and U22017 (N_22017,N_19398,N_19450);
and U22018 (N_22018,N_18781,N_20348);
or U22019 (N_22019,N_19936,N_19563);
nand U22020 (N_22020,N_19233,N_20314);
xor U22021 (N_22021,N_21018,N_19978);
xnor U22022 (N_22022,N_19786,N_18780);
or U22023 (N_22023,N_21754,N_20732);
nor U22024 (N_22024,N_20186,N_19481);
and U22025 (N_22025,N_20949,N_21304);
nand U22026 (N_22026,N_20310,N_21234);
xor U22027 (N_22027,N_20176,N_20853);
xor U22028 (N_22028,N_19740,N_19162);
nand U22029 (N_22029,N_21859,N_20402);
and U22030 (N_22030,N_21025,N_21066);
and U22031 (N_22031,N_20161,N_20414);
nand U22032 (N_22032,N_21515,N_19022);
and U22033 (N_22033,N_19361,N_19268);
nor U22034 (N_22034,N_19620,N_21851);
and U22035 (N_22035,N_19001,N_21595);
nand U22036 (N_22036,N_18795,N_20377);
and U22037 (N_22037,N_21021,N_20566);
or U22038 (N_22038,N_19796,N_19903);
nor U22039 (N_22039,N_20125,N_18857);
nor U22040 (N_22040,N_19981,N_21530);
and U22041 (N_22041,N_19346,N_21132);
xor U22042 (N_22042,N_20953,N_21867);
and U22043 (N_22043,N_20671,N_20920);
nand U22044 (N_22044,N_20371,N_21287);
nand U22045 (N_22045,N_21099,N_21430);
or U22046 (N_22046,N_20784,N_19248);
or U22047 (N_22047,N_21784,N_20360);
nand U22048 (N_22048,N_19935,N_19168);
xor U22049 (N_22049,N_20839,N_21101);
and U22050 (N_22050,N_19921,N_21733);
nand U22051 (N_22051,N_19500,N_21729);
and U22052 (N_22052,N_20267,N_20112);
nand U22053 (N_22053,N_18799,N_21838);
and U22054 (N_22054,N_20676,N_19850);
nand U22055 (N_22055,N_21320,N_21811);
nor U22056 (N_22056,N_19388,N_19082);
nand U22057 (N_22057,N_21124,N_21688);
nand U22058 (N_22058,N_19783,N_20173);
and U22059 (N_22059,N_19661,N_18767);
and U22060 (N_22060,N_20948,N_20046);
xnor U22061 (N_22061,N_21721,N_19621);
nand U22062 (N_22062,N_21775,N_21139);
nor U22063 (N_22063,N_20707,N_19348);
nor U22064 (N_22064,N_21763,N_20900);
and U22065 (N_22065,N_19625,N_21477);
nand U22066 (N_22066,N_19823,N_21872);
nand U22067 (N_22067,N_19066,N_20221);
and U22068 (N_22068,N_18859,N_19768);
or U22069 (N_22069,N_20867,N_21807);
or U22070 (N_22070,N_20689,N_21318);
or U22071 (N_22071,N_21160,N_21815);
nand U22072 (N_22072,N_21189,N_19843);
nand U22073 (N_22073,N_21566,N_18880);
nor U22074 (N_22074,N_20118,N_20800);
nand U22075 (N_22075,N_21211,N_21168);
xor U22076 (N_22076,N_21195,N_21847);
and U22077 (N_22077,N_19018,N_20504);
nor U22078 (N_22078,N_21632,N_18865);
and U22079 (N_22079,N_20634,N_21187);
xor U22080 (N_22080,N_19185,N_21053);
nand U22081 (N_22081,N_19177,N_20378);
nand U22082 (N_22082,N_18881,N_19610);
nor U22083 (N_22083,N_20632,N_19065);
and U22084 (N_22084,N_19369,N_21868);
and U22085 (N_22085,N_19826,N_21464);
nor U22086 (N_22086,N_19867,N_20554);
and U22087 (N_22087,N_19148,N_21358);
and U22088 (N_22088,N_20965,N_19928);
nor U22089 (N_22089,N_20884,N_21400);
and U22090 (N_22090,N_18867,N_21239);
nor U22091 (N_22091,N_18877,N_20994);
nand U22092 (N_22092,N_19280,N_19725);
or U22093 (N_22093,N_19020,N_20281);
or U22094 (N_22094,N_21502,N_20429);
and U22095 (N_22095,N_20133,N_20809);
and U22096 (N_22096,N_20436,N_18823);
xor U22097 (N_22097,N_20082,N_19767);
and U22098 (N_22098,N_19231,N_19904);
nand U22099 (N_22099,N_20442,N_20189);
nor U22100 (N_22100,N_21609,N_20938);
xnor U22101 (N_22101,N_18783,N_21288);
nand U22102 (N_22102,N_19984,N_18873);
nand U22103 (N_22103,N_19580,N_20787);
nand U22104 (N_22104,N_19735,N_20475);
nor U22105 (N_22105,N_21303,N_21735);
and U22106 (N_22106,N_19820,N_20395);
and U22107 (N_22107,N_19688,N_19045);
nor U22108 (N_22108,N_20263,N_21179);
nand U22109 (N_22109,N_19766,N_19827);
xor U22110 (N_22110,N_19597,N_21086);
xor U22111 (N_22111,N_21216,N_20775);
and U22112 (N_22112,N_21292,N_20404);
xnor U22113 (N_22113,N_19855,N_19641);
nand U22114 (N_22114,N_19942,N_20983);
nor U22115 (N_22115,N_20690,N_19853);
nor U22116 (N_22116,N_20776,N_20160);
nor U22117 (N_22117,N_19111,N_19085);
and U22118 (N_22118,N_19042,N_21087);
nor U22119 (N_22119,N_19646,N_20647);
nor U22120 (N_22120,N_20880,N_21014);
and U22121 (N_22121,N_19590,N_19556);
and U22122 (N_22122,N_21653,N_18987);
nor U22123 (N_22123,N_20641,N_20207);
or U22124 (N_22124,N_21438,N_20912);
nand U22125 (N_22125,N_19657,N_21152);
nand U22126 (N_22126,N_19209,N_21486);
xnor U22127 (N_22127,N_20225,N_20851);
xor U22128 (N_22128,N_21163,N_18809);
and U22129 (N_22129,N_18937,N_21030);
or U22130 (N_22130,N_19502,N_19953);
or U22131 (N_22131,N_20633,N_19550);
or U22132 (N_22132,N_18752,N_20100);
and U22133 (N_22133,N_21011,N_18977);
or U22134 (N_22134,N_18888,N_19630);
or U22135 (N_22135,N_20233,N_19672);
nor U22136 (N_22136,N_21026,N_21630);
nand U22137 (N_22137,N_21448,N_19432);
xor U22138 (N_22138,N_21204,N_19551);
or U22139 (N_22139,N_19321,N_19807);
and U22140 (N_22140,N_19011,N_19100);
or U22141 (N_22141,N_19659,N_19472);
nor U22142 (N_22142,N_18784,N_20032);
nor U22143 (N_22143,N_19083,N_21006);
and U22144 (N_22144,N_20505,N_21835);
nor U22145 (N_22145,N_20878,N_21806);
and U22146 (N_22146,N_19704,N_18849);
and U22147 (N_22147,N_21857,N_18957);
or U22148 (N_22148,N_19894,N_21821);
xor U22149 (N_22149,N_19519,N_19679);
nand U22150 (N_22150,N_19165,N_19362);
nand U22151 (N_22151,N_21529,N_20447);
nand U22152 (N_22152,N_18872,N_19193);
nand U22153 (N_22153,N_21517,N_21415);
nor U22154 (N_22154,N_18952,N_21186);
nand U22155 (N_22155,N_20113,N_20055);
nor U22156 (N_22156,N_18900,N_21795);
or U22157 (N_22157,N_20908,N_20275);
nor U22158 (N_22158,N_19565,N_20175);
and U22159 (N_22159,N_21230,N_20235);
xor U22160 (N_22160,N_21315,N_21575);
nor U22161 (N_22161,N_20295,N_19763);
nand U22162 (N_22162,N_20393,N_18860);
nor U22163 (N_22163,N_21793,N_20023);
xnor U22164 (N_22164,N_21581,N_20342);
and U22165 (N_22165,N_20537,N_19663);
nor U22166 (N_22166,N_20365,N_21107);
nand U22167 (N_22167,N_20198,N_21656);
and U22168 (N_22168,N_20401,N_21064);
nor U22169 (N_22169,N_21037,N_21192);
xnor U22170 (N_22170,N_19062,N_19393);
nor U22171 (N_22171,N_21297,N_19579);
nand U22172 (N_22172,N_20083,N_19093);
nand U22173 (N_22173,N_20381,N_18970);
nand U22174 (N_22174,N_20069,N_19637);
nor U22175 (N_22175,N_20902,N_19632);
nand U22176 (N_22176,N_21626,N_18946);
and U22177 (N_22177,N_19098,N_20387);
or U22178 (N_22178,N_20128,N_21412);
xnor U22179 (N_22179,N_18759,N_19308);
and U22180 (N_22180,N_19094,N_19558);
and U22181 (N_22181,N_20539,N_20076);
or U22182 (N_22182,N_19635,N_20306);
xnor U22183 (N_22183,N_20795,N_20296);
nand U22184 (N_22184,N_20887,N_20205);
and U22185 (N_22185,N_21310,N_20397);
nand U22186 (N_22186,N_20626,N_20535);
and U22187 (N_22187,N_20150,N_20238);
and U22188 (N_22188,N_20199,N_21406);
xor U22189 (N_22189,N_20635,N_19913);
nor U22190 (N_22190,N_18886,N_21191);
nand U22191 (N_22191,N_21308,N_19128);
and U22192 (N_22192,N_21823,N_21788);
nor U22193 (N_22193,N_19864,N_19803);
or U22194 (N_22194,N_19596,N_19443);
or U22195 (N_22195,N_21732,N_19560);
and U22196 (N_22196,N_21833,N_20211);
or U22197 (N_22197,N_20322,N_21428);
and U22198 (N_22198,N_20833,N_20312);
or U22199 (N_22199,N_21646,N_19033);
nor U22200 (N_22200,N_20542,N_21748);
and U22201 (N_22201,N_19517,N_19583);
nor U22202 (N_22202,N_21584,N_20723);
and U22203 (N_22203,N_20773,N_20817);
nor U22204 (N_22204,N_19441,N_20558);
or U22205 (N_22205,N_21177,N_20557);
nand U22206 (N_22206,N_20291,N_21178);
xor U22207 (N_22207,N_19306,N_19969);
or U22208 (N_22208,N_21360,N_20328);
xor U22209 (N_22209,N_20164,N_20258);
nand U22210 (N_22210,N_20611,N_19754);
nand U22211 (N_22211,N_19199,N_20599);
nand U22212 (N_22212,N_20490,N_21055);
nand U22213 (N_22213,N_19239,N_20203);
nor U22214 (N_22214,N_19531,N_21786);
and U22215 (N_22215,N_21022,N_20813);
or U22216 (N_22216,N_20659,N_20143);
nor U22217 (N_22217,N_18948,N_20666);
nor U22218 (N_22218,N_20785,N_21343);
nand U22219 (N_22219,N_19535,N_21028);
or U22220 (N_22220,N_20280,N_21142);
nor U22221 (N_22221,N_21072,N_18861);
nand U22222 (N_22222,N_20202,N_20740);
and U22223 (N_22223,N_18840,N_21834);
and U22224 (N_22224,N_20792,N_21715);
nand U22225 (N_22225,N_18955,N_20520);
nor U22226 (N_22226,N_21692,N_21621);
and U22227 (N_22227,N_19157,N_20375);
or U22228 (N_22228,N_18838,N_21705);
nor U22229 (N_22229,N_19092,N_20568);
nor U22230 (N_22230,N_21557,N_19110);
xnor U22231 (N_22231,N_21813,N_21500);
nand U22232 (N_22232,N_20540,N_21232);
and U22233 (N_22233,N_20279,N_21274);
nand U22234 (N_22234,N_21712,N_19702);
and U22235 (N_22235,N_19989,N_19760);
nand U22236 (N_22236,N_19249,N_18813);
or U22237 (N_22237,N_19470,N_20793);
nand U22238 (N_22238,N_20008,N_20122);
or U22239 (N_22239,N_18884,N_20517);
or U22240 (N_22240,N_19409,N_20509);
nor U22241 (N_22241,N_21435,N_18899);
xnor U22242 (N_22242,N_20941,N_20685);
nor U22243 (N_22243,N_19707,N_20521);
nand U22244 (N_22244,N_19648,N_20005);
or U22245 (N_22245,N_21624,N_19782);
xnor U22246 (N_22246,N_19835,N_20054);
or U22247 (N_22247,N_19190,N_20768);
nand U22248 (N_22248,N_19815,N_18958);
or U22249 (N_22249,N_21175,N_20910);
or U22250 (N_22250,N_18908,N_20670);
or U22251 (N_22251,N_18976,N_19647);
or U22252 (N_22252,N_19125,N_21042);
nor U22253 (N_22253,N_19272,N_20935);
nand U22254 (N_22254,N_20229,N_20081);
and U22255 (N_22255,N_19628,N_19337);
nor U22256 (N_22256,N_21659,N_19276);
or U22257 (N_22257,N_18928,N_20187);
xor U22258 (N_22258,N_21518,N_19521);
or U22259 (N_22259,N_19771,N_21331);
and U22260 (N_22260,N_19357,N_20484);
nand U22261 (N_22261,N_20665,N_21468);
nor U22262 (N_22262,N_19709,N_20970);
nor U22263 (N_22263,N_21062,N_21057);
and U22264 (N_22264,N_20063,N_20019);
nor U22265 (N_22265,N_20237,N_20837);
and U22266 (N_22266,N_21678,N_20584);
xnor U22267 (N_22267,N_21660,N_18782);
and U22268 (N_22268,N_20960,N_19699);
nand U22269 (N_22269,N_20944,N_21150);
xor U22270 (N_22270,N_19330,N_18858);
and U22271 (N_22271,N_21466,N_20619);
and U22272 (N_22272,N_19949,N_19608);
nor U22273 (N_22273,N_20731,N_21046);
nor U22274 (N_22274,N_19420,N_19617);
or U22275 (N_22275,N_21212,N_21869);
or U22276 (N_22276,N_19962,N_19080);
nor U22277 (N_22277,N_20828,N_19857);
xnor U22278 (N_22278,N_20273,N_19320);
nand U22279 (N_22279,N_21840,N_20876);
nor U22280 (N_22280,N_18851,N_19207);
and U22281 (N_22281,N_18933,N_20648);
or U22282 (N_22282,N_19799,N_19000);
or U22283 (N_22283,N_18753,N_19731);
and U22284 (N_22284,N_21096,N_20257);
and U22285 (N_22285,N_18924,N_20148);
nand U22286 (N_22286,N_18964,N_20260);
and U22287 (N_22287,N_21804,N_20188);
nor U22288 (N_22288,N_19872,N_19684);
and U22289 (N_22289,N_21585,N_21153);
or U22290 (N_22290,N_21004,N_20230);
xor U22291 (N_22291,N_18918,N_19848);
and U22292 (N_22292,N_19652,N_19738);
nand U22293 (N_22293,N_19192,N_21606);
or U22294 (N_22294,N_20718,N_20391);
or U22295 (N_22295,N_18969,N_20214);
and U22296 (N_22296,N_21612,N_20170);
or U22297 (N_22297,N_19299,N_19313);
nand U22298 (N_22298,N_19683,N_20323);
xor U22299 (N_22299,N_19076,N_19455);
and U22300 (N_22300,N_18999,N_21709);
and U22301 (N_22301,N_19780,N_19129);
or U22302 (N_22302,N_18750,N_20906);
or U22303 (N_22303,N_18931,N_19339);
or U22304 (N_22304,N_20615,N_19211);
and U22305 (N_22305,N_19452,N_20162);
and U22306 (N_22306,N_20012,N_21576);
nor U22307 (N_22307,N_20448,N_19077);
or U22308 (N_22308,N_19595,N_21613);
or U22309 (N_22309,N_19744,N_19909);
and U22310 (N_22310,N_20077,N_21684);
nor U22311 (N_22311,N_21069,N_21776);
nand U22312 (N_22312,N_20159,N_19957);
nand U22313 (N_22313,N_21002,N_19200);
or U22314 (N_22314,N_21742,N_21451);
and U22315 (N_22315,N_21134,N_21221);
or U22316 (N_22316,N_21545,N_20067);
xor U22317 (N_22317,N_20049,N_19405);
nand U22318 (N_22318,N_19234,N_20645);
nand U22319 (N_22319,N_20832,N_20702);
and U22320 (N_22320,N_19252,N_20749);
and U22321 (N_22321,N_19266,N_19940);
nand U22322 (N_22322,N_20465,N_20037);
nand U22323 (N_22323,N_20982,N_20169);
and U22324 (N_22324,N_20918,N_20577);
and U22325 (N_22325,N_19607,N_21637);
and U22326 (N_22326,N_19107,N_18853);
and U22327 (N_22327,N_19273,N_19779);
nor U22328 (N_22328,N_20048,N_19651);
or U22329 (N_22329,N_21129,N_19064);
nor U22330 (N_22330,N_21662,N_21527);
or U22331 (N_22331,N_21362,N_21569);
or U22332 (N_22332,N_19967,N_19026);
and U22333 (N_22333,N_19220,N_20097);
or U22334 (N_22334,N_20673,N_21238);
and U22335 (N_22335,N_18806,N_19166);
nor U22336 (N_22336,N_21631,N_21185);
and U22337 (N_22337,N_20576,N_20743);
and U22338 (N_22338,N_21726,N_19349);
nor U22339 (N_22339,N_19530,N_20114);
and U22340 (N_22340,N_19973,N_19331);
or U22341 (N_22341,N_21299,N_20687);
nor U22342 (N_22342,N_19353,N_20123);
or U22343 (N_22343,N_19633,N_21095);
or U22344 (N_22344,N_21388,N_20873);
or U22345 (N_22345,N_19510,N_19467);
nor U22346 (N_22346,N_21407,N_20388);
or U22347 (N_22347,N_18911,N_18844);
nand U22348 (N_22348,N_19809,N_21844);
nand U22349 (N_22349,N_19374,N_19791);
or U22350 (N_22350,N_19060,N_20512);
nand U22351 (N_22351,N_19179,N_20178);
nand U22352 (N_22352,N_21141,N_18779);
or U22353 (N_22353,N_19021,N_20471);
and U22354 (N_22354,N_21452,N_19706);
xor U22355 (N_22355,N_19655,N_20350);
nand U22356 (N_22356,N_20620,N_21829);
and U22357 (N_22357,N_21526,N_21745);
or U22358 (N_22358,N_19619,N_19477);
or U22359 (N_22359,N_20823,N_21738);
or U22360 (N_22360,N_20129,N_21802);
nand U22361 (N_22361,N_21245,N_19847);
and U22362 (N_22362,N_20803,N_21118);
nand U22363 (N_22363,N_19236,N_18950);
or U22364 (N_22364,N_19176,N_19992);
nand U22365 (N_22365,N_20643,N_21675);
and U22366 (N_22366,N_20014,N_18934);
xnor U22367 (N_22367,N_21373,N_19845);
nand U22368 (N_22368,N_21643,N_19309);
or U22369 (N_22369,N_19539,N_19955);
or U22370 (N_22370,N_21206,N_20503);
or U22371 (N_22371,N_21294,N_19139);
and U22372 (N_22372,N_19424,N_20571);
and U22373 (N_22373,N_21854,N_19151);
nand U22374 (N_22374,N_19440,N_20763);
nand U22375 (N_22375,N_18871,N_19370);
xor U22376 (N_22376,N_18972,N_21397);
and U22377 (N_22377,N_21233,N_21326);
xnor U22378 (N_22378,N_21871,N_18856);
and U22379 (N_22379,N_19664,N_18814);
nor U22380 (N_22380,N_20145,N_19980);
or U22381 (N_22381,N_21340,N_20013);
or U22382 (N_22382,N_19392,N_19070);
and U22383 (N_22383,N_19351,N_19537);
nor U22384 (N_22384,N_20245,N_21849);
nand U22385 (N_22385,N_20091,N_19333);
nand U22386 (N_22386,N_21345,N_20575);
or U22387 (N_22387,N_20562,N_20142);
nor U22388 (N_22388,N_20410,N_19584);
and U22389 (N_22389,N_21555,N_19629);
and U22390 (N_22390,N_18920,N_20406);
nand U22391 (N_22391,N_21597,N_21263);
or U22392 (N_22392,N_19713,N_21483);
nand U22393 (N_22393,N_21202,N_19158);
nand U22394 (N_22394,N_21778,N_19126);
nor U22395 (N_22395,N_19216,N_18968);
nor U22396 (N_22396,N_20859,N_21682);
or U22397 (N_22397,N_19897,N_20578);
xor U22398 (N_22398,N_19422,N_21696);
or U22399 (N_22399,N_19429,N_19821);
or U22400 (N_22400,N_21032,N_21383);
or U22401 (N_22401,N_19419,N_19068);
and U22402 (N_22402,N_19923,N_21789);
nor U22403 (N_22403,N_21511,N_20255);
and U22404 (N_22404,N_21197,N_20915);
and U22405 (N_22405,N_21182,N_18876);
nor U22406 (N_22406,N_21372,N_20086);
or U22407 (N_22407,N_18763,N_19053);
or U22408 (N_22408,N_18775,N_19317);
and U22409 (N_22409,N_19479,N_18898);
and U22410 (N_22410,N_19007,N_18930);
nor U22411 (N_22411,N_21280,N_21727);
or U22412 (N_22412,N_19426,N_20212);
nor U22413 (N_22413,N_18778,N_19938);
or U22414 (N_22414,N_21572,N_21542);
nor U22415 (N_22415,N_19078,N_20553);
or U22416 (N_22416,N_21719,N_18875);
and U22417 (N_22417,N_18923,N_19051);
and U22418 (N_22418,N_19756,N_18825);
nor U22419 (N_22419,N_20977,N_20753);
or U22420 (N_22420,N_21173,N_20272);
or U22421 (N_22421,N_21366,N_19951);
nor U22422 (N_22422,N_20024,N_21476);
nor U22423 (N_22423,N_19132,N_19097);
or U22424 (N_22424,N_19952,N_21490);
nor U22425 (N_22425,N_21311,N_19063);
and U22426 (N_22426,N_21335,N_19837);
nor U22427 (N_22427,N_20226,N_20637);
xor U22428 (N_22428,N_20701,N_20065);
nor U22429 (N_22429,N_20259,N_20498);
nor U22430 (N_22430,N_19013,N_20950);
and U22431 (N_22431,N_18793,N_20863);
nand U22432 (N_22432,N_20136,N_20196);
and U22433 (N_22433,N_21493,N_19716);
nor U22434 (N_22434,N_19178,N_19545);
and U22435 (N_22435,N_21751,N_21454);
and U22436 (N_22436,N_19464,N_21669);
nor U22437 (N_22437,N_19366,N_21620);
nor U22438 (N_22438,N_19764,N_21841);
xor U22439 (N_22439,N_20814,N_21290);
xnor U22440 (N_22440,N_19552,N_21506);
nand U22441 (N_22441,N_19059,N_21339);
and U22442 (N_22442,N_20734,N_21162);
nand U22443 (N_22443,N_20499,N_19964);
or U22444 (N_22444,N_18798,N_20893);
and U22445 (N_22445,N_19528,N_21019);
nand U22446 (N_22446,N_20572,N_19592);
xor U22447 (N_22447,N_21780,N_18832);
xor U22448 (N_22448,N_19163,N_18895);
and U22449 (N_22449,N_21144,N_20421);
xor U22450 (N_22450,N_21352,N_18756);
nand U22451 (N_22451,N_20165,N_20058);
and U22452 (N_22452,N_21785,N_21654);
and U22453 (N_22453,N_19930,N_19613);
nand U22454 (N_22454,N_21200,N_20010);
xnor U22455 (N_22455,N_20684,N_20827);
or U22456 (N_22456,N_18981,N_21601);
nand U22457 (N_22457,N_21773,N_20688);
and U22458 (N_22458,N_19471,N_19839);
or U22459 (N_22459,N_19622,N_21083);
nor U22460 (N_22460,N_19084,N_19746);
nand U22461 (N_22461,N_19569,N_21111);
or U22462 (N_22462,N_20845,N_21401);
nor U22463 (N_22463,N_20998,N_19161);
or U22464 (N_22464,N_20061,N_21571);
and U22465 (N_22465,N_21540,N_19381);
or U22466 (N_22466,N_20380,N_19736);
nand U22467 (N_22467,N_19985,N_19403);
xor U22468 (N_22468,N_20075,N_20480);
or U22469 (N_22469,N_20527,N_19237);
nor U22470 (N_22470,N_21627,N_20339);
xnor U22471 (N_22471,N_21676,N_20758);
and U22472 (N_22472,N_19873,N_20979);
or U22473 (N_22473,N_18810,N_21762);
nor U22474 (N_22474,N_19439,N_21307);
xor U22475 (N_22475,N_19876,N_21718);
xnor U22476 (N_22476,N_20035,N_21092);
or U22477 (N_22477,N_21702,N_19055);
xnor U22478 (N_22478,N_19734,N_19024);
and U22479 (N_22479,N_21136,N_18816);
xor U22480 (N_22480,N_18988,N_20710);
nand U22481 (N_22481,N_19676,N_21552);
nor U22482 (N_22482,N_20709,N_18953);
and U22483 (N_22483,N_19972,N_20976);
and U22484 (N_22484,N_19282,N_20654);
or U22485 (N_22485,N_19609,N_20779);
and U22486 (N_22486,N_20904,N_20737);
nand U22487 (N_22487,N_21717,N_21409);
and U22488 (N_22488,N_19680,N_20104);
and U22489 (N_22489,N_20117,N_20786);
nand U22490 (N_22490,N_19533,N_19862);
and U22491 (N_22491,N_18975,N_18786);
nor U22492 (N_22492,N_20791,N_20427);
nor U22493 (N_22493,N_20361,N_20997);
or U22494 (N_22494,N_21741,N_19790);
nand U22495 (N_22495,N_21183,N_21009);
nand U22496 (N_22496,N_20705,N_21487);
nor U22497 (N_22497,N_19495,N_21861);
nand U22498 (N_22498,N_20595,N_21048);
nor U22499 (N_22499,N_20493,N_19461);
nor U22500 (N_22500,N_20213,N_19542);
nor U22501 (N_22501,N_19150,N_19677);
nand U22502 (N_22502,N_20455,N_20330);
and U22503 (N_22503,N_20969,N_18922);
and U22504 (N_22504,N_20463,N_21396);
nand U22505 (N_22505,N_19697,N_21359);
or U22506 (N_22506,N_19124,N_21647);
or U22507 (N_22507,N_19303,N_19260);
nor U22508 (N_22508,N_19326,N_20336);
and U22509 (N_22509,N_19698,N_20349);
nor U22510 (N_22510,N_19057,N_19931);
nor U22511 (N_22511,N_20748,N_20500);
and U22512 (N_22512,N_20411,N_21610);
nand U22513 (N_22513,N_19222,N_21458);
nor U22514 (N_22514,N_20006,N_20894);
nor U22515 (N_22515,N_20971,N_19501);
or U22516 (N_22516,N_19536,N_18939);
nor U22517 (N_22517,N_18834,N_21301);
and U22518 (N_22518,N_20254,N_19476);
nand U22519 (N_22519,N_20777,N_19588);
or U22520 (N_22520,N_20802,N_20721);
xnor U22521 (N_22521,N_19974,N_20771);
nor U22522 (N_22522,N_20501,N_19567);
and U22523 (N_22523,N_20340,N_20451);
or U22524 (N_22524,N_21091,N_20990);
or U22525 (N_22525,N_20897,N_20171);
or U22526 (N_22526,N_18926,N_20140);
nor U22527 (N_22527,N_19300,N_21272);
nor U22528 (N_22528,N_20826,N_20516);
nand U22529 (N_22529,N_19777,N_18915);
xnor U22530 (N_22530,N_21323,N_19367);
nor U22531 (N_22531,N_21003,N_19474);
and U22532 (N_22532,N_21138,N_20445);
or U22533 (N_22533,N_20929,N_19889);
nor U22534 (N_22534,N_19149,N_19329);
nor U22535 (N_22535,N_19612,N_19882);
or U22536 (N_22536,N_21724,N_18940);
and U22537 (N_22537,N_19979,N_18847);
nor U22538 (N_22538,N_21514,N_19307);
nand U22539 (N_22539,N_21089,N_20888);
nor U22540 (N_22540,N_21651,N_19181);
nand U22541 (N_22541,N_19058,N_18829);
nor U22542 (N_22542,N_21864,N_21102);
nor U22543 (N_22543,N_21264,N_21420);
and U22544 (N_22544,N_20120,N_21337);
and U22545 (N_22545,N_21753,N_21273);
nand U22546 (N_22546,N_20804,N_21342);
or U22547 (N_22547,N_19154,N_21169);
nand U22548 (N_22548,N_20264,N_20986);
nand U22549 (N_22549,N_19714,N_19770);
xnor U22550 (N_22550,N_20495,N_18949);
or U22551 (N_22551,N_21497,N_19755);
nand U22552 (N_22552,N_20570,N_18815);
xnor U22553 (N_22553,N_19954,N_21224);
or U22554 (N_22554,N_19122,N_19288);
nand U22555 (N_22555,N_21519,N_20073);
and U22556 (N_22556,N_19994,N_19250);
nand U22557 (N_22557,N_20699,N_20925);
and U22558 (N_22558,N_18760,N_20588);
nand U22559 (N_22559,N_19352,N_19513);
nand U22560 (N_22560,N_21207,N_19397);
or U22561 (N_22561,N_20244,N_19976);
nor U22562 (N_22562,N_20439,N_21758);
nand U22563 (N_22563,N_18882,N_19460);
and U22564 (N_22564,N_20222,N_19769);
and U22565 (N_22565,N_19488,N_21663);
nand U22566 (N_22566,N_20177,N_19396);
nor U22567 (N_22567,N_21067,N_21368);
and U22568 (N_22568,N_19049,N_19660);
and U22569 (N_22569,N_19627,N_20598);
nor U22570 (N_22570,N_21333,N_20890);
and U22571 (N_22571,N_21521,N_21130);
nor U22572 (N_22572,N_19877,N_19776);
xor U22573 (N_22573,N_20957,N_21357);
and U22574 (N_22574,N_20134,N_21393);
and U22575 (N_22575,N_21286,N_21856);
nor U22576 (N_22576,N_20752,N_19520);
and U22577 (N_22577,N_21598,N_21463);
and U22578 (N_22578,N_19749,N_20528);
or U22579 (N_22579,N_20473,N_19462);
nor U22580 (N_22580,N_20001,N_18866);
and U22581 (N_22581,N_18789,N_19143);
nor U22582 (N_22582,N_20385,N_21461);
nand U22583 (N_22583,N_20724,N_21036);
nand U22584 (N_22584,N_21779,N_18768);
nor U22585 (N_22585,N_21213,N_21743);
nor U22586 (N_22586,N_21208,N_19413);
and U22587 (N_22587,N_19828,N_21475);
nor U22588 (N_22588,N_18917,N_20507);
or U22589 (N_22589,N_21312,N_19712);
or U22590 (N_22590,N_21691,N_21769);
nor U22591 (N_22591,N_19640,N_20868);
nand U22592 (N_22592,N_21270,N_18912);
or U22593 (N_22593,N_20251,N_20760);
nor U22594 (N_22594,N_21243,N_19116);
nor U22595 (N_22595,N_20438,N_19708);
xnor U22596 (N_22596,N_21378,N_21604);
or U22597 (N_22597,N_21855,N_19834);
nand U22598 (N_22598,N_20959,N_21471);
nor U22599 (N_22599,N_19037,N_20491);
nand U22600 (N_22600,N_18776,N_21269);
and U22601 (N_22601,N_20821,N_19818);
nor U22602 (N_22602,N_20218,N_20921);
nor U22603 (N_22603,N_19578,N_20441);
or U22604 (N_22604,N_19902,N_20607);
nand U22605 (N_22605,N_18833,N_20329);
xnor U22606 (N_22606,N_19485,N_20108);
nor U22607 (N_22607,N_21842,N_20679);
nor U22608 (N_22608,N_20094,N_21282);
or U22609 (N_22609,N_19408,N_20234);
xor U22610 (N_22610,N_20288,N_21749);
nand U22611 (N_22611,N_19449,N_18796);
and U22612 (N_22612,N_21755,N_19591);
xnor U22613 (N_22613,N_21363,N_19244);
nand U22614 (N_22614,N_21051,N_19983);
nand U22615 (N_22615,N_19189,N_21792);
nor U22616 (N_22616,N_21482,N_19251);
and U22617 (N_22617,N_21324,N_19670);
or U22618 (N_22618,N_21166,N_19491);
or U22619 (N_22619,N_21457,N_20745);
xor U22620 (N_22620,N_19484,N_20031);
or U22621 (N_22621,N_19836,N_20716);
and U22622 (N_22622,N_21513,N_20068);
xor U22623 (N_22623,N_19998,N_20951);
nor U22624 (N_22624,N_20370,N_20742);
nor U22625 (N_22625,N_20909,N_21033);
nand U22626 (N_22626,N_20834,N_21645);
nand U22627 (N_22627,N_19691,N_21825);
nor U22628 (N_22628,N_19915,N_20765);
or U22629 (N_22629,N_19912,N_20783);
nand U22630 (N_22630,N_21445,N_20469);
or U22631 (N_22631,N_21336,N_20007);
nor U22632 (N_22632,N_19448,N_19854);
and U22633 (N_22633,N_19269,N_19830);
nor U22634 (N_22634,N_20919,N_20232);
or U22635 (N_22635,N_20372,N_19759);
nor U22636 (N_22636,N_21781,N_20124);
nor U22637 (N_22637,N_20703,N_18792);
and U22638 (N_22638,N_19840,N_20840);
and U22639 (N_22639,N_21043,N_21240);
or U22640 (N_22640,N_20911,N_19841);
and U22641 (N_22641,N_20300,N_19056);
nand U22642 (N_22642,N_20583,N_21275);
and U22643 (N_22643,N_20518,N_19028);
or U22644 (N_22644,N_21370,N_19005);
or U22645 (N_22645,N_21070,N_19871);
and U22646 (N_22646,N_20650,N_21424);
and U22647 (N_22647,N_21596,N_19336);
xor U22648 (N_22648,N_21531,N_21629);
and U22649 (N_22649,N_19345,N_20327);
xor U22650 (N_22650,N_21686,N_20754);
nand U22651 (N_22651,N_19598,N_20636);
nor U22652 (N_22652,N_18824,N_20662);
and U22653 (N_22653,N_18902,N_21744);
and U22654 (N_22654,N_21484,N_19425);
or U22655 (N_22655,N_21429,N_19226);
nand U22656 (N_22656,N_20613,N_21668);
nand U22657 (N_22657,N_21300,N_20192);
nand U22658 (N_22658,N_19965,N_19741);
and U22659 (N_22659,N_20801,N_21338);
nor U22660 (N_22660,N_18996,N_21865);
nor U22661 (N_22661,N_19858,N_21005);
nor U22662 (N_22662,N_19451,N_21453);
and U22663 (N_22663,N_21085,N_19908);
nand U22664 (N_22664,N_19412,N_21058);
xnor U22665 (N_22665,N_19039,N_19860);
nor U22666 (N_22666,N_21012,N_18998);
nand U22667 (N_22667,N_19512,N_19656);
and U22668 (N_22668,N_18901,N_19813);
nor U22669 (N_22669,N_20115,N_19174);
or U22670 (N_22670,N_19874,N_19798);
or U22671 (N_22671,N_21255,N_19762);
or U22672 (N_22672,N_18942,N_19407);
or U22673 (N_22673,N_18887,N_19486);
xnor U22674 (N_22674,N_20989,N_21774);
and U22675 (N_22675,N_19543,N_21485);
or U22676 (N_22676,N_19113,N_21685);
and U22677 (N_22677,N_21607,N_21029);
or U22678 (N_22678,N_19692,N_19559);
nand U22679 (N_22679,N_21425,N_20105);
or U22680 (N_22680,N_21683,N_18929);
and U22681 (N_22681,N_21472,N_18966);
nand U22682 (N_22682,N_19230,N_19215);
nand U22683 (N_22683,N_19261,N_18910);
xnor U22684 (N_22684,N_21830,N_19722);
nor U22685 (N_22685,N_19564,N_19208);
and U22686 (N_22686,N_19073,N_20616);
xnor U22687 (N_22687,N_19599,N_21710);
nand U22688 (N_22688,N_18843,N_18837);
or U22689 (N_22689,N_18836,N_19851);
or U22690 (N_22690,N_19228,N_20559);
xor U22691 (N_22691,N_19890,N_18994);
nand U22692 (N_22692,N_19091,N_20556);
nand U22693 (N_22693,N_19727,N_18963);
nand U22694 (N_22694,N_20905,N_18869);
nand U22695 (N_22695,N_20223,N_19946);
or U22696 (N_22696,N_20138,N_21469);
or U22697 (N_22697,N_20593,N_20119);
nand U22698 (N_22698,N_20000,N_21316);
and U22699 (N_22699,N_21707,N_20585);
nor U22700 (N_22700,N_18986,N_21223);
and U22701 (N_22701,N_20009,N_21137);
nand U22702 (N_22702,N_21344,N_18980);
or U22703 (N_22703,N_21664,N_18774);
xor U22704 (N_22704,N_19456,N_21665);
nor U22705 (N_22705,N_20759,N_18919);
xnor U22706 (N_22706,N_20738,N_20324);
and U22707 (N_22707,N_21328,N_19870);
or U22708 (N_22708,N_20550,N_20974);
nor U22709 (N_22709,N_18754,N_21494);
or U22710 (N_22710,N_21752,N_18913);
or U22711 (N_22711,N_21228,N_20822);
nor U22712 (N_22712,N_19932,N_20923);
nand U22713 (N_22713,N_19988,N_19138);
xnor U22714 (N_22714,N_21140,N_21110);
nand U22715 (N_22715,N_20297,N_18839);
nor U22716 (N_22716,N_20877,N_18835);
nor U22717 (N_22717,N_21305,N_20713);
and U22718 (N_22718,N_18794,N_21699);
or U22719 (N_22719,N_19970,N_20195);
nand U22720 (N_22720,N_20220,N_21225);
or U22721 (N_22721,N_18936,N_21302);
nand U22722 (N_22722,N_20579,N_20303);
nand U22723 (N_22723,N_19270,N_21579);
or U22724 (N_22724,N_21681,N_20675);
nand U22725 (N_22725,N_21381,N_19996);
and U22726 (N_22726,N_19197,N_19522);
nand U22727 (N_22727,N_21131,N_19040);
nand U22728 (N_22728,N_19112,N_20541);
or U22729 (N_22729,N_21151,N_20589);
nand U22730 (N_22730,N_20824,N_19861);
and U22731 (N_22731,N_19365,N_19032);
and U22732 (N_22732,N_21848,N_19096);
and U22733 (N_22733,N_19050,N_21853);
and U22734 (N_22734,N_20062,N_19682);
xor U22735 (N_22735,N_20183,N_21251);
nor U22736 (N_22736,N_18997,N_20798);
nand U22737 (N_22737,N_20651,N_20871);
and U22738 (N_22738,N_20274,N_19376);
nand U22739 (N_22739,N_19901,N_20066);
nor U22740 (N_22740,N_20376,N_21017);
nor U22741 (N_22741,N_19188,N_21480);
nand U22742 (N_22742,N_21084,N_18984);
and U22743 (N_22743,N_19038,N_20767);
nor U22744 (N_22744,N_21309,N_19990);
nor U22745 (N_22745,N_20021,N_19423);
nor U22746 (N_22746,N_20457,N_20677);
and U22747 (N_22747,N_20733,N_19748);
nor U22748 (N_22748,N_20363,N_21109);
nor U22749 (N_22749,N_19274,N_19600);
or U22750 (N_22750,N_21098,N_18827);
and U22751 (N_22751,N_21436,N_21117);
nor U22752 (N_22752,N_18896,N_19445);
or U22753 (N_22753,N_19180,N_20268);
and U22754 (N_22754,N_21289,N_20603);
or U22755 (N_22755,N_21704,N_21574);
or U22756 (N_22756,N_19603,N_18770);
nor U22757 (N_22757,N_21801,N_21209);
nor U22758 (N_22758,N_20681,N_20590);
nor U22759 (N_22759,N_21532,N_20538);
and U22760 (N_22760,N_18971,N_19997);
xor U22761 (N_22761,N_20131,N_20942);
or U22762 (N_22762,N_19343,N_21426);
or U22763 (N_22763,N_21404,N_20004);
and U22764 (N_22764,N_19480,N_19002);
nand U22765 (N_22765,N_20916,N_20631);
or U22766 (N_22766,N_20755,N_20789);
or U22767 (N_22767,N_21405,N_18909);
nand U22768 (N_22768,N_19371,N_21293);
nor U22769 (N_22769,N_19071,N_19153);
and U22770 (N_22770,N_20796,N_18846);
xnor U22771 (N_22771,N_20625,N_21268);
nand U22772 (N_22772,N_20514,N_19172);
or U22773 (N_22773,N_20722,N_19614);
nor U22774 (N_22774,N_21076,N_19743);
xnor U22775 (N_22775,N_21027,N_19146);
nor U22776 (N_22776,N_21593,N_19752);
and U22777 (N_22777,N_20883,N_19701);
or U22778 (N_22778,N_19119,N_20107);
nand U22779 (N_22779,N_21812,N_20034);
or U22780 (N_22780,N_19095,N_19415);
and U22781 (N_22781,N_20761,N_20174);
or U22782 (N_22782,N_20700,N_20256);
or U22783 (N_22783,N_21413,N_21170);
nand U22784 (N_22784,N_19099,N_20831);
nor U22785 (N_22785,N_19863,N_19304);
xnor U22786 (N_22786,N_20623,N_20629);
xnor U22787 (N_22787,N_20892,N_19265);
nand U22788 (N_22788,N_20808,N_20040);
and U22789 (N_22789,N_19822,N_21817);
or U22790 (N_22790,N_19285,N_21622);
nor U22791 (N_22791,N_19993,N_20003);
and U22792 (N_22792,N_20555,N_19377);
nand U22793 (N_22793,N_20240,N_18787);
nor U22794 (N_22794,N_21433,N_19003);
or U22795 (N_22795,N_20712,N_20400);
nor U22796 (N_22796,N_19810,N_20351);
or U22797 (N_22797,N_19438,N_21045);
or U22798 (N_22798,N_19732,N_21496);
xnor U22799 (N_22799,N_20565,N_20180);
and U22800 (N_22800,N_20937,N_21222);
or U22801 (N_22801,N_19382,N_19044);
nor U22802 (N_22802,N_19043,N_19899);
and U22803 (N_22803,N_21176,N_20769);
and U22804 (N_22804,N_20630,N_19380);
nand U22805 (N_22805,N_19418,N_20751);
nand U22806 (N_22806,N_19875,N_21462);
or U22807 (N_22807,N_21852,N_20658);
or U22808 (N_22808,N_20270,N_19605);
nand U22809 (N_22809,N_21567,N_18960);
nand U22810 (N_22810,N_19133,N_20284);
nand U22811 (N_22811,N_19718,N_20396);
nor U22812 (N_22812,N_19281,N_19373);
or U22813 (N_22813,N_21246,N_20366);
or U22814 (N_22814,N_19114,N_20283);
nand U22815 (N_22815,N_21711,N_21695);
nor U22816 (N_22816,N_20686,N_19884);
nor U22817 (N_22817,N_19792,N_18916);
nor U22818 (N_22818,N_21599,N_20204);
or U22819 (N_22819,N_20903,N_21387);
or U22820 (N_22820,N_21180,N_19717);
nor U22821 (N_22821,N_20946,N_19947);
and U22822 (N_22822,N_19503,N_19417);
nand U22823 (N_22823,N_21777,N_19103);
nor U22824 (N_22824,N_19920,N_19642);
nand U22825 (N_22825,N_21419,N_20262);
nand U22826 (N_22826,N_20510,N_21220);
or U22827 (N_22827,N_21700,N_20343);
nand U22828 (N_22828,N_20052,N_20835);
or U22829 (N_22829,N_19943,N_20456);
nor U22830 (N_22830,N_20027,N_21088);
or U22831 (N_22831,N_20985,N_20711);
nand U22832 (N_22832,N_19896,N_21049);
xnor U22833 (N_22833,N_21509,N_20139);
and U22834 (N_22834,N_19386,N_20999);
nand U22835 (N_22835,N_21874,N_21155);
nand U22836 (N_22836,N_20246,N_19218);
nand U22837 (N_22837,N_21060,N_21159);
nor U22838 (N_22838,N_19507,N_20652);
nor U22839 (N_22839,N_19014,N_21672);
and U22840 (N_22840,N_20126,N_20874);
and U22841 (N_22841,N_20392,N_20846);
nor U22842 (N_22842,N_19259,N_21505);
nand U22843 (N_22843,N_20276,N_21796);
and U22844 (N_22844,N_21608,N_19347);
or U22845 (N_22845,N_19968,N_21498);
or U22846 (N_22846,N_19387,N_21577);
xor U22847 (N_22847,N_19747,N_19088);
nor U22848 (N_22848,N_21016,N_18893);
nor U22849 (N_22849,N_19399,N_21056);
or U22850 (N_22850,N_21285,N_21123);
nor U22851 (N_22851,N_19258,N_18961);
and U22852 (N_22852,N_21768,N_21190);
nor U22853 (N_22853,N_20975,N_18852);
and U22854 (N_22854,N_20726,N_19294);
xnor U22855 (N_22855,N_21499,N_20519);
nand U22856 (N_22856,N_19298,N_20071);
nor U22857 (N_22857,N_20020,N_21615);
and U22858 (N_22858,N_19577,N_21024);
or U22859 (N_22859,N_19842,N_21543);
nand U22860 (N_22860,N_18956,N_19434);
xor U22861 (N_22861,N_19594,N_19223);
nor U22862 (N_22862,N_21443,N_21115);
xnor U22863 (N_22863,N_21592,N_20318);
nor U22864 (N_22864,N_21706,N_20266);
nand U22865 (N_22865,N_18820,N_18819);
or U22866 (N_22866,N_21757,N_19482);
or U22867 (N_22867,N_20413,N_19447);
nor U22868 (N_22868,N_18818,N_19694);
nand U22869 (N_22869,N_20956,N_18868);
nand U22870 (N_22870,N_21819,N_19238);
nand U22871 (N_22871,N_21538,N_19561);
or U22872 (N_22872,N_21473,N_21047);
nor U22873 (N_22873,N_19264,N_19905);
and U22874 (N_22874,N_21020,N_21219);
nor U22875 (N_22875,N_19856,N_21201);
xnor U22876 (N_22876,N_18890,N_21537);
or U22877 (N_22877,N_20099,N_18995);
nand U22878 (N_22878,N_21583,N_21348);
nand U22879 (N_22879,N_21196,N_18841);
and U22880 (N_22880,N_19134,N_21638);
nand U22881 (N_22881,N_20591,N_20092);
nand U22882 (N_22882,N_20452,N_21655);
or U22883 (N_22883,N_21810,N_19278);
nand U22884 (N_22884,N_21495,N_19893);
nor U22885 (N_22885,N_19497,N_21361);
and U22886 (N_22886,N_21694,N_20337);
or U22887 (N_22887,N_21623,N_19052);
nor U22888 (N_22888,N_19459,N_19696);
nor U22889 (N_22889,N_19910,N_18751);
nand U22890 (N_22890,N_21799,N_18932);
or U22891 (N_22891,N_19131,N_20669);
and U22892 (N_22892,N_20309,N_19917);
nand U22893 (N_22893,N_20374,N_21728);
and U22894 (N_22894,N_20345,N_20523);
and U22895 (N_22895,N_21602,N_21467);
nand U22896 (N_22896,N_20939,N_20958);
or U22897 (N_22897,N_21410,N_19316);
or U22898 (N_22898,N_19549,N_19108);
or U22899 (N_22899,N_21794,N_20231);
nand U22900 (N_22900,N_19120,N_19673);
nand U22901 (N_22901,N_21374,N_19478);
or U22902 (N_22902,N_19945,N_20219);
and U22903 (N_22903,N_20458,N_20151);
nor U22904 (N_22904,N_20981,N_19433);
and U22905 (N_22905,N_19626,N_21670);
and U22906 (N_22906,N_21347,N_19529);
nand U22907 (N_22907,N_19205,N_19719);
and U22908 (N_22908,N_20227,N_18757);
nand U22909 (N_22909,N_21689,N_21635);
nor U22910 (N_22910,N_21148,N_21671);
and U22911 (N_22911,N_20747,N_19332);
xnor U22912 (N_22912,N_21052,N_19217);
and U22913 (N_22913,N_21001,N_21281);
nor U22914 (N_22914,N_19730,N_19925);
and U22915 (N_22915,N_20934,N_20770);
nor U22916 (N_22916,N_18862,N_19341);
or U22917 (N_22917,N_21256,N_19156);
nand U22918 (N_22918,N_21650,N_19137);
or U22919 (N_22919,N_20354,N_20865);
nor U22920 (N_22920,N_19645,N_21603);
nand U22921 (N_22921,N_21354,N_20482);
or U22922 (N_22922,N_20101,N_19886);
nand U22923 (N_22923,N_21253,N_19287);
and U22924 (N_22924,N_21417,N_19636);
and U22925 (N_22925,N_20181,N_19173);
nand U22926 (N_22926,N_20078,N_19383);
or U22927 (N_22927,N_19898,N_19130);
or U22928 (N_22928,N_20434,N_21097);
xor U22929 (N_22929,N_21039,N_20033);
nor U22930 (N_22930,N_20836,N_20355);
nor U22931 (N_22931,N_20587,N_20952);
and U22932 (N_22932,N_19008,N_19653);
nor U22933 (N_22933,N_21356,N_21442);
xnor U22934 (N_22934,N_19681,N_18947);
and U22935 (N_22935,N_20682,N_20592);
or U22936 (N_22936,N_20022,N_18785);
xor U22937 (N_22937,N_19658,N_20708);
nand U22938 (N_22938,N_19726,N_20663);
nand U22939 (N_22939,N_20102,N_20774);
and U22940 (N_22940,N_20545,N_21369);
or U22941 (N_22941,N_20311,N_20842);
nand U22942 (N_22942,N_21826,N_18889);
and U22943 (N_22943,N_21522,N_20628);
or U22944 (N_22944,N_19802,N_19245);
and U22945 (N_22945,N_19571,N_21822);
or U22946 (N_22946,N_19442,N_20489);
and U22947 (N_22947,N_19906,N_19900);
nand U22948 (N_22948,N_20638,N_19555);
nor U22949 (N_22949,N_19687,N_21364);
or U22950 (N_22950,N_20788,N_19141);
nor U22951 (N_22951,N_21334,N_19784);
nor U22952 (N_22952,N_20604,N_18883);
or U22953 (N_22953,N_20781,N_19167);
nor U22954 (N_22954,N_21283,N_19171);
or U22955 (N_22955,N_21231,N_19690);
or U22956 (N_22956,N_21846,N_19212);
or U22957 (N_22957,N_18874,N_20466);
and U22958 (N_22958,N_19671,N_21217);
nor U22959 (N_22959,N_21698,N_20210);
or U22960 (N_22960,N_19808,N_21023);
and U22961 (N_22961,N_20966,N_19924);
and U22962 (N_22962,N_18904,N_21386);
nor U22963 (N_22963,N_21797,N_20459);
nor U22964 (N_22964,N_21143,N_21441);
nand U22965 (N_22965,N_21128,N_21422);
nand U22966 (N_22966,N_20660,N_21330);
nor U22967 (N_22967,N_19394,N_21090);
or U22968 (N_22968,N_19515,N_19624);
nand U22969 (N_22969,N_21474,N_19775);
or U22970 (N_22970,N_19453,N_21737);
or U22971 (N_22971,N_19186,N_21481);
nand U22972 (N_22972,N_20358,N_18765);
nor U22973 (N_22973,N_19389,N_20168);
or U22974 (N_22974,N_19492,N_21389);
nand U22975 (N_22975,N_20468,N_21171);
or U22976 (N_22976,N_20474,N_18897);
nand U22977 (N_22977,N_20347,N_21587);
nor U22978 (N_22978,N_21618,N_21582);
nand U22979 (N_22979,N_20933,N_21787);
nand U22980 (N_22980,N_20432,N_21820);
and U22981 (N_22981,N_21164,N_18761);
xor U22982 (N_22982,N_20430,N_21157);
nand U22983 (N_22983,N_18811,N_20678);
nor U22984 (N_22984,N_19224,N_19667);
or U22985 (N_22985,N_20386,N_21261);
nor U22986 (N_22986,N_20253,N_20610);
and U22987 (N_22987,N_19358,N_20423);
or U22988 (N_22988,N_19914,N_21418);
nor U22989 (N_22989,N_19036,N_18771);
and U22990 (N_22990,N_20191,N_19788);
nor U22991 (N_22991,N_21114,N_18979);
nor U22992 (N_22992,N_21640,N_21558);
or U22993 (N_22993,N_19372,N_21648);
nor U22994 (N_22994,N_19887,N_21278);
or U22995 (N_22995,N_21271,N_19035);
or U22996 (N_22996,N_21536,N_21353);
xor U22997 (N_22997,N_21491,N_19489);
nor U22998 (N_22998,N_21346,N_20250);
nand U22999 (N_22999,N_20762,N_19283);
nand U23000 (N_23000,N_19499,N_21355);
and U23001 (N_23001,N_20581,N_20522);
and U23002 (N_23002,N_20201,N_21181);
or U23003 (N_23003,N_21759,N_18764);
or U23004 (N_23004,N_19087,N_20524);
xor U23005 (N_23005,N_19950,N_20353);
nand U23006 (N_23006,N_21121,N_20407);
nand U23007 (N_23007,N_19662,N_21590);
and U23008 (N_23008,N_19164,N_20194);
or U23009 (N_23009,N_21332,N_20051);
and U23010 (N_23010,N_21394,N_20529);
or U23011 (N_23011,N_21465,N_21750);
or U23012 (N_23012,N_21193,N_21554);
nand U23013 (N_23013,N_19573,N_18925);
xor U23014 (N_23014,N_19801,N_19546);
and U23015 (N_23015,N_21377,N_20428);
or U23016 (N_23016,N_19356,N_21439);
nand U23017 (N_23017,N_21693,N_20379);
and U23018 (N_23018,N_19589,N_20326);
and U23019 (N_23019,N_19534,N_19883);
or U23020 (N_23020,N_18978,N_19256);
or U23021 (N_23021,N_19048,N_19866);
or U23022 (N_23022,N_18894,N_21747);
nor U23023 (N_23023,N_19384,N_20551);
xnor U23024 (N_23024,N_19029,N_18803);
and U23025 (N_23025,N_20167,N_21570);
nand U23026 (N_23026,N_20715,N_21677);
nand U23027 (N_23027,N_20460,N_21546);
xor U23028 (N_23028,N_20667,N_20228);
and U23029 (N_23029,N_20533,N_18801);
or U23030 (N_23030,N_19025,N_21565);
and U23031 (N_23031,N_21298,N_21516);
nor U23032 (N_23032,N_21734,N_21731);
nor U23033 (N_23033,N_20302,N_20158);
nand U23034 (N_23034,N_19463,N_20812);
and U23035 (N_23035,N_19054,N_19568);
nand U23036 (N_23036,N_21427,N_20672);
nor U23037 (N_23037,N_20015,N_20317);
nand U23038 (N_23038,N_19437,N_19700);
nand U23039 (N_23039,N_20750,N_19705);
or U23040 (N_23040,N_20277,N_21034);
or U23041 (N_23041,N_19325,N_19926);
nor U23042 (N_23042,N_21639,N_19031);
and U23043 (N_23043,N_19363,N_19401);
or U23044 (N_23044,N_21044,N_19527);
and U23045 (N_23045,N_20056,N_19674);
nand U23046 (N_23046,N_21081,N_21260);
or U23047 (N_23047,N_20841,N_19575);
and U23048 (N_23048,N_20025,N_19041);
nor U23049 (N_23049,N_21539,N_21687);
nand U23050 (N_23050,N_21548,N_20534);
nor U23051 (N_23051,N_20098,N_20901);
and U23052 (N_23052,N_21035,N_20972);
and U23053 (N_23053,N_20815,N_19301);
nor U23054 (N_23054,N_19009,N_19089);
nand U23055 (N_23055,N_19465,N_20440);
or U23056 (N_23056,N_20472,N_18828);
xor U23057 (N_23057,N_19991,N_20418);
nand U23058 (N_23058,N_21798,N_18864);
nor U23059 (N_23059,N_20072,N_21563);
and U23060 (N_23060,N_19868,N_21736);
nor U23061 (N_23061,N_20166,N_21119);
or U23062 (N_23062,N_19086,N_20130);
and U23063 (N_23063,N_20810,N_19315);
nand U23064 (N_23064,N_21295,N_21440);
nand U23065 (N_23065,N_21351,N_20121);
or U23066 (N_23066,N_19314,N_19939);
or U23067 (N_23067,N_19355,N_20955);
and U23068 (N_23068,N_20156,N_20891);
nand U23069 (N_23069,N_19368,N_21716);
or U23070 (N_23070,N_19436,N_21450);
nand U23071 (N_23071,N_19819,N_20844);
or U23072 (N_23072,N_21827,N_19075);
nand U23073 (N_23073,N_21319,N_21007);
and U23074 (N_23074,N_21258,N_20869);
nand U23075 (N_23075,N_21235,N_21808);
nand U23076 (N_23076,N_21227,N_20087);
and U23077 (N_23077,N_19916,N_19105);
or U23078 (N_23078,N_20879,N_20642);
and U23079 (N_23079,N_18921,N_19375);
xnor U23080 (N_23080,N_21205,N_20334);
nor U23081 (N_23081,N_20356,N_21722);
and U23082 (N_23082,N_20973,N_19229);
and U23083 (N_23083,N_20617,N_19292);
or U23084 (N_23084,N_19811,N_19421);
and U23085 (N_23085,N_20298,N_21158);
xor U23086 (N_23086,N_21690,N_20861);
nand U23087 (N_23087,N_19342,N_19468);
or U23088 (N_23088,N_19685,N_20450);
nor U23089 (N_23089,N_20409,N_19958);
and U23090 (N_23090,N_19160,N_19277);
nand U23091 (N_23091,N_19203,N_19327);
nand U23092 (N_23092,N_20088,N_20485);
nor U23093 (N_23093,N_19079,N_20315);
or U23094 (N_23094,N_21321,N_18962);
nand U23095 (N_23095,N_21156,N_20680);
and U23096 (N_23096,N_19196,N_19271);
or U23097 (N_23097,N_18808,N_20182);
or U23098 (N_23098,N_19204,N_20582);
nand U23099 (N_23099,N_21642,N_20954);
and U23100 (N_23100,N_20215,N_18812);
xnor U23101 (N_23101,N_20127,N_20567);
or U23102 (N_23102,N_21459,N_20216);
nor U23103 (N_23103,N_20487,N_20511);
xor U23104 (N_23104,N_20940,N_21244);
and U23105 (N_23105,N_21135,N_20346);
or U23106 (N_23106,N_19724,N_19106);
nand U23107 (N_23107,N_19475,N_19444);
xnor U23108 (N_23108,N_21210,N_21074);
nand U23109 (N_23109,N_20525,N_21831);
and U23110 (N_23110,N_20497,N_21528);
nor U23111 (N_23111,N_20816,N_21636);
nor U23112 (N_23112,N_20057,N_19523);
and U23113 (N_23113,N_20486,N_19284);
or U23114 (N_23114,N_21306,N_21071);
or U23115 (N_23115,N_20477,N_18903);
xor U23116 (N_23116,N_21740,N_21573);
and U23117 (N_23117,N_20847,N_21094);
and U23118 (N_23118,N_21199,N_20819);
xor U23119 (N_23119,N_20179,N_20627);
nand U23120 (N_23120,N_18791,N_19865);
and U23121 (N_23121,N_19869,N_19833);
nand U23122 (N_23122,N_19720,N_20331);
nand U23123 (N_23123,N_19340,N_18821);
and U23124 (N_23124,N_20991,N_19566);
xor U23125 (N_23125,N_20184,N_20043);
xor U23126 (N_23126,N_20424,N_18855);
nand U23127 (N_23127,N_20605,N_21791);
or U23128 (N_23128,N_21254,N_19322);
nand U23129 (N_23129,N_18943,N_20437);
nand U23130 (N_23130,N_20190,N_19206);
or U23131 (N_23131,N_20594,N_19963);
xnor U23132 (N_23132,N_19570,N_19169);
and U23133 (N_23133,N_21560,N_19253);
and U23134 (N_23134,N_20412,N_21549);
nor U23135 (N_23135,N_18797,N_21279);
and U23136 (N_23136,N_20596,N_21479);
or U23137 (N_23137,N_21284,N_19262);
and U23138 (N_23138,N_19127,N_19728);
or U23139 (N_23139,N_21146,N_19540);
nand U23140 (N_23140,N_20357,N_21723);
nand U23141 (N_23141,N_20993,N_21106);
or U23142 (N_23142,N_20294,N_19240);
or U23143 (N_23143,N_20764,N_20289);
nor U23144 (N_23144,N_19496,N_20293);
nand U23145 (N_23145,N_21104,N_20612);
and U23146 (N_23146,N_20932,N_18941);
nand U23147 (N_23147,N_19831,N_19631);
nor U23148 (N_23148,N_20039,N_21126);
or U23149 (N_23149,N_20018,N_21040);
and U23150 (N_23150,N_21503,N_19379);
xor U23151 (N_23151,N_19639,N_20962);
or U23152 (N_23152,N_20308,N_19505);
xor U23153 (N_23153,N_20155,N_19891);
and U23154 (N_23154,N_19907,N_21068);
nand U23155 (N_23155,N_21247,N_19689);
nand U23156 (N_23156,N_20208,N_20564);
nand U23157 (N_23157,N_19311,N_20805);
nor U23158 (N_23158,N_19402,N_21214);
xnor U23159 (N_23159,N_21031,N_19695);
xnor U23160 (N_23160,N_20547,N_21421);
nor U23161 (N_23161,N_19514,N_21772);
nor U23162 (N_23162,N_21375,N_21431);
or U23163 (N_23163,N_19668,N_19665);
or U23164 (N_23164,N_20924,N_21644);
xnor U23165 (N_23165,N_20560,N_20987);
and U23166 (N_23166,N_19601,N_19016);
nor U23167 (N_23167,N_21666,N_21229);
and U23168 (N_23168,N_20382,N_19971);
nand U23169 (N_23169,N_19147,N_19115);
or U23170 (N_23170,N_20265,N_19508);
xnor U23171 (N_23171,N_20416,N_20064);
nand U23172 (N_23172,N_20408,N_21215);
nand U23173 (N_23173,N_21525,N_21456);
and U23174 (N_23174,N_19785,N_21380);
and U23175 (N_23175,N_20344,N_19959);
and U23176 (N_23176,N_19703,N_19279);
nor U23177 (N_23177,N_20872,N_20811);
or U23178 (N_23178,N_19742,N_21828);
and U23179 (N_23179,N_20964,N_19750);
and U23180 (N_23180,N_20079,N_21093);
or U23181 (N_23181,N_18807,N_21589);
and U23182 (N_23182,N_19602,N_21008);
nand U23183 (N_23183,N_21510,N_19751);
nor U23184 (N_23184,N_20193,N_19525);
and U23185 (N_23185,N_19986,N_20106);
or U23186 (N_23186,N_19975,N_19638);
or U23187 (N_23187,N_21845,N_21000);
nand U23188 (N_23188,N_20913,N_19030);
and U23189 (N_23189,N_21873,N_20478);
or U23190 (N_23190,N_21080,N_19290);
and U23191 (N_23191,N_21824,N_21329);
nand U23192 (N_23192,N_21839,N_20552);
nand U23193 (N_23193,N_19257,N_19615);
and U23194 (N_23194,N_21739,N_20369);
nand U23195 (N_23195,N_19034,N_20041);
and U23196 (N_23196,N_21108,N_20889);
or U23197 (N_23197,N_19654,N_20085);
or U23198 (N_23198,N_20029,N_21147);
xnor U23199 (N_23199,N_19574,N_20304);
nand U23200 (N_23200,N_20896,N_20320);
and U23201 (N_23201,N_21814,N_19391);
and U23202 (N_23202,N_20580,N_21697);
and U23203 (N_23203,N_20197,N_21790);
xnor U23204 (N_23204,N_20243,N_21408);
and U23205 (N_23205,N_19844,N_21616);
or U23206 (N_23206,N_19944,N_19604);
xor U23207 (N_23207,N_21832,N_21127);
or U23208 (N_23208,N_20316,N_19919);
and U23209 (N_23209,N_21259,N_20403);
and U23210 (N_23210,N_20807,N_20144);
and U23211 (N_23211,N_21172,N_20907);
and U23212 (N_23212,N_19295,N_21382);
and U23213 (N_23213,N_19243,N_20389);
and U23214 (N_23214,N_21725,N_20794);
and U23215 (N_23215,N_20886,N_19761);
nand U23216 (N_23216,N_21322,N_21625);
nor U23217 (N_23217,N_21188,N_20530);
nor U23218 (N_23218,N_20730,N_19297);
xor U23219 (N_23219,N_19184,N_19982);
and U23220 (N_23220,N_19509,N_20135);
or U23221 (N_23221,N_18854,N_20858);
nand U23222 (N_23222,N_20248,N_21535);
nor U23223 (N_23223,N_21564,N_19140);
nand U23224 (N_23224,N_20462,N_19814);
and U23225 (N_23225,N_19587,N_19446);
and U23226 (N_23226,N_19027,N_18817);
nor U23227 (N_23227,N_21674,N_19123);
xnor U23228 (N_23228,N_20172,N_21313);
or U23229 (N_23229,N_19721,N_20922);
nor U23230 (N_23230,N_21341,N_18891);
nor U23231 (N_23231,N_21619,N_20597);
nor U23232 (N_23232,N_19246,N_21291);
nand U23233 (N_23233,N_20206,N_19805);
nand U23234 (N_23234,N_20074,N_19593);
nor U23235 (N_23235,N_19427,N_20546);
or U23236 (N_23236,N_20084,N_21756);
and U23237 (N_23237,N_20852,N_20341);
and U23238 (N_23238,N_18885,N_19334);
and U23239 (N_23239,N_21816,N_19305);
nor U23240 (N_23240,N_19047,N_20825);
and U23241 (N_23241,N_21446,N_18879);
xnor U23242 (N_23242,N_19323,N_20947);
or U23243 (N_23243,N_20435,N_20875);
or U23244 (N_23244,N_21803,N_20321);
nor U23245 (N_23245,N_20573,N_19338);
nand U23246 (N_23246,N_19781,N_21050);
nor U23247 (N_23247,N_19118,N_19616);
nand U23248 (N_23248,N_18758,N_18927);
xor U23249 (N_23249,N_21470,N_19948);
and U23250 (N_23250,N_21414,N_19538);
nor U23251 (N_23251,N_18906,N_20093);
nand U23252 (N_23252,N_21252,N_19458);
nand U23253 (N_23253,N_21365,N_20419);
nor U23254 (N_23254,N_20044,N_20036);
nor U23255 (N_23255,N_21437,N_18982);
nand U23256 (N_23256,N_21125,N_18935);
or U23257 (N_23257,N_20278,N_18907);
and U23258 (N_23258,N_20531,N_21658);
nand U23259 (N_23259,N_20319,N_20980);
nor U23260 (N_23260,N_20691,N_19933);
and U23261 (N_23261,N_20829,N_18989);
or U23262 (N_23262,N_19109,N_20961);
or U23263 (N_23263,N_20502,N_21236);
nand U23264 (N_23264,N_18892,N_19800);
and U23265 (N_23265,N_20359,N_19772);
and U23266 (N_23266,N_18878,N_20103);
or U23267 (N_23267,N_21550,N_18842);
nor U23268 (N_23268,N_20080,N_19774);
or U23269 (N_23269,N_20506,N_21591);
nand U23270 (N_23270,N_21562,N_21449);
xnor U23271 (N_23271,N_20431,N_20449);
nand U23272 (N_23272,N_21652,N_19739);
and U23273 (N_23273,N_19121,N_20420);
and U23274 (N_23274,N_19494,N_20060);
and U23275 (N_23275,N_20694,N_20606);
nand U23276 (N_23276,N_19888,N_21082);
nand U23277 (N_23277,N_19623,N_20443);
or U23278 (N_23278,N_20930,N_19678);
and U23279 (N_23279,N_19576,N_20683);
or U23280 (N_23280,N_20618,N_19142);
or U23281 (N_23281,N_20549,N_18762);
and U23282 (N_23282,N_21079,N_21818);
xnor U23283 (N_23283,N_21863,N_21447);
and U23284 (N_23284,N_19012,N_21679);
and U23285 (N_23285,N_20111,N_19019);
and U23286 (N_23286,N_20050,N_20563);
or U23287 (N_23287,N_20574,N_20415);
nor U23288 (N_23288,N_21403,N_21760);
nand U23289 (N_23289,N_18870,N_19895);
nor U23290 (N_23290,N_19715,N_18992);
and U23291 (N_23291,N_21038,N_19404);
and U23292 (N_23292,N_21628,N_19710);
nor U23293 (N_23293,N_19956,N_18845);
nor U23294 (N_23294,N_20995,N_18826);
and U23295 (N_23295,N_20744,N_19918);
or U23296 (N_23296,N_20927,N_21578);
and U23297 (N_23297,N_21657,N_20984);
and U23298 (N_23298,N_21100,N_21262);
or U23299 (N_23299,N_19562,N_19960);
and U23300 (N_23300,N_21041,N_21489);
or U23301 (N_23301,N_18802,N_20695);
xor U23302 (N_23302,N_19431,N_19255);
or U23303 (N_23303,N_20154,N_20394);
nor U23304 (N_23304,N_21015,N_19829);
or U23305 (N_23305,N_19937,N_19061);
nand U23306 (N_23306,N_20729,N_19004);
and U23307 (N_23307,N_20070,N_20644);
and U23308 (N_23308,N_20332,N_20714);
or U23309 (N_23309,N_19198,N_21588);
and U23310 (N_23310,N_19553,N_18985);
and U23311 (N_23311,N_20137,N_21390);
xor U23312 (N_23312,N_21241,N_19400);
nor U23313 (N_23313,N_19170,N_19435);
nor U23314 (N_23314,N_21746,N_18777);
nand U23315 (N_23315,N_20059,N_20778);
and U23316 (N_23316,N_20600,N_20727);
nand U23317 (N_23317,N_21237,N_19411);
nor U23318 (N_23318,N_19466,N_19483);
nand U23319 (N_23319,N_20536,N_19155);
and U23320 (N_23320,N_18974,N_20287);
or U23321 (N_23321,N_21113,N_19817);
nor U23322 (N_23322,N_18769,N_21078);
or U23323 (N_23323,N_20996,N_19225);
xnor U23324 (N_23324,N_20285,N_20820);
xor U23325 (N_23325,N_20914,N_20854);
nand U23326 (N_23326,N_21198,N_18965);
or U23327 (N_23327,N_20978,N_21194);
and U23328 (N_23328,N_21122,N_21398);
nand U23329 (N_23329,N_20968,N_20338);
and U23330 (N_23330,N_20532,N_19081);
nor U23331 (N_23331,N_20857,N_18766);
xor U23332 (N_23332,N_21392,N_20797);
nand U23333 (N_23333,N_20089,N_20157);
and U23334 (N_23334,N_19611,N_19023);
or U23335 (N_23335,N_19017,N_20674);
or U23336 (N_23336,N_21544,N_20757);
and U23337 (N_23337,N_20467,N_20367);
nand U23338 (N_23338,N_19219,N_19010);
xor U23339 (N_23339,N_18983,N_21568);
nand U23340 (N_23340,N_20739,N_19557);
nand U23341 (N_23341,N_18790,N_19378);
nor U23342 (N_23342,N_20147,N_20185);
and U23343 (N_23343,N_19878,N_20943);
nand U23344 (N_23344,N_19881,N_21367);
or U23345 (N_23345,N_19686,N_19666);
nand U23346 (N_23346,N_19344,N_20002);
xor U23347 (N_23347,N_19359,N_18973);
and U23348 (N_23348,N_20045,N_19669);
and U23349 (N_23349,N_20864,N_20639);
xnor U23350 (N_23350,N_19364,N_18959);
and U23351 (N_23351,N_21423,N_21504);
or U23352 (N_23352,N_19067,N_19232);
nor U23353 (N_23353,N_21703,N_19832);
and U23354 (N_23354,N_19753,N_20446);
nor U23355 (N_23355,N_20479,N_21073);
or U23356 (N_23356,N_18850,N_20719);
nand U23357 (N_23357,N_20290,N_19516);
nand U23358 (N_23358,N_19526,N_20095);
and U23359 (N_23359,N_20384,N_20657);
or U23360 (N_23360,N_20492,N_21520);
or U23361 (N_23361,N_20704,N_21120);
nor U23362 (N_23362,N_21594,N_21837);
nor U23363 (N_23363,N_19286,N_19410);
or U23364 (N_23364,N_20149,N_18944);
xnor U23365 (N_23365,N_20269,N_21661);
and U23366 (N_23366,N_21764,N_20333);
and U23367 (N_23367,N_20496,N_21063);
nor U23368 (N_23368,N_20621,N_19247);
nor U23369 (N_23369,N_19929,N_21783);
or U23370 (N_23370,N_19101,N_19723);
and U23371 (N_23371,N_19941,N_20843);
xor U23372 (N_23372,N_21858,N_21761);
nor U23373 (N_23373,N_19778,N_20271);
or U23374 (N_23374,N_21149,N_20882);
xor U23375 (N_23375,N_21649,N_20735);
nand U23376 (N_23376,N_19135,N_19117);
nand U23377 (N_23377,N_20931,N_20224);
and U23378 (N_23378,N_21054,N_20141);
or U23379 (N_23379,N_20640,N_20543);
nand U23380 (N_23380,N_19541,N_20849);
nor U23381 (N_23381,N_20926,N_21523);
and U23382 (N_23382,N_20895,N_21553);
nor U23383 (N_23383,N_21154,N_20728);
or U23384 (N_23384,N_21455,N_21145);
or U23385 (N_23385,N_21103,N_21501);
nor U23386 (N_23386,N_19074,N_19758);
or U23387 (N_23387,N_21701,N_19733);
or U23388 (N_23388,N_21508,N_20282);
and U23389 (N_23389,N_20481,N_20494);
nand U23390 (N_23390,N_21730,N_20110);
xor U23391 (N_23391,N_18945,N_20464);
nand U23392 (N_23392,N_20109,N_19498);
xor U23393 (N_23393,N_20655,N_19104);
xnor U23394 (N_23394,N_20866,N_20042);
or U23395 (N_23395,N_19175,N_21065);
or U23396 (N_23396,N_19291,N_19544);
and U23397 (N_23397,N_21010,N_19961);
xor U23398 (N_23398,N_20301,N_20028);
or U23399 (N_23399,N_21765,N_20898);
nor U23400 (N_23400,N_18990,N_20780);
and U23401 (N_23401,N_21203,N_21860);
xnor U23402 (N_23402,N_20163,N_19069);
nand U23403 (N_23403,N_21492,N_20664);
or U23404 (N_23404,N_21533,N_21327);
nand U23405 (N_23405,N_20053,N_18954);
and U23406 (N_23406,N_21242,N_21411);
and U23407 (N_23407,N_20569,N_21551);
and U23408 (N_23408,N_21296,N_19966);
nor U23409 (N_23409,N_19922,N_20717);
or U23410 (N_23410,N_20368,N_21460);
nor U23411 (N_23411,N_18951,N_20364);
nand U23412 (N_23412,N_21614,N_19511);
or U23413 (N_23413,N_20422,N_18830);
nor U23414 (N_23414,N_20488,N_20656);
and U23415 (N_23415,N_20692,N_20249);
and U23416 (N_23416,N_21771,N_20362);
nor U23417 (N_23417,N_21714,N_19046);
or U23418 (N_23418,N_19195,N_19145);
nand U23419 (N_23419,N_19310,N_20325);
or U23420 (N_23420,N_19504,N_19804);
or U23421 (N_23421,N_19765,N_19711);
or U23422 (N_23422,N_20693,N_21434);
or U23423 (N_23423,N_21395,N_20885);
or U23424 (N_23424,N_21634,N_21541);
or U23425 (N_23425,N_18848,N_21350);
xor U23426 (N_23426,N_20899,N_20242);
or U23427 (N_23427,N_21809,N_18914);
or U23428 (N_23428,N_20855,N_21174);
nand U23429 (N_23429,N_20782,N_20261);
or U23430 (N_23430,N_21385,N_19350);
or U23431 (N_23431,N_19194,N_19254);
nor U23432 (N_23432,N_18804,N_20090);
and U23433 (N_23433,N_20988,N_19849);
nand U23434 (N_23434,N_19518,N_21314);
and U23435 (N_23435,N_19581,N_20299);
nand U23436 (N_23436,N_19210,N_19757);
and U23437 (N_23437,N_19999,N_20576);
nor U23438 (N_23438,N_19407,N_21154);
xor U23439 (N_23439,N_20247,N_21744);
nor U23440 (N_23440,N_18812,N_21811);
nor U23441 (N_23441,N_21330,N_20693);
and U23442 (N_23442,N_19671,N_20441);
or U23443 (N_23443,N_21643,N_19138);
nor U23444 (N_23444,N_20302,N_19601);
xnor U23445 (N_23445,N_19448,N_19394);
and U23446 (N_23446,N_20922,N_20473);
nor U23447 (N_23447,N_21611,N_18856);
nor U23448 (N_23448,N_20548,N_19000);
nand U23449 (N_23449,N_21580,N_20130);
and U23450 (N_23450,N_18811,N_20358);
nand U23451 (N_23451,N_20937,N_21357);
or U23452 (N_23452,N_21637,N_20741);
xor U23453 (N_23453,N_21642,N_20244);
and U23454 (N_23454,N_20800,N_20060);
nor U23455 (N_23455,N_21110,N_21811);
nand U23456 (N_23456,N_20593,N_20284);
nand U23457 (N_23457,N_20681,N_19425);
and U23458 (N_23458,N_20242,N_20537);
nand U23459 (N_23459,N_20950,N_21547);
or U23460 (N_23460,N_19107,N_19644);
nand U23461 (N_23461,N_20339,N_20436);
xnor U23462 (N_23462,N_21505,N_21484);
and U23463 (N_23463,N_21778,N_20760);
xnor U23464 (N_23464,N_21711,N_19710);
nand U23465 (N_23465,N_21466,N_21434);
or U23466 (N_23466,N_20088,N_20232);
or U23467 (N_23467,N_20771,N_21770);
and U23468 (N_23468,N_19539,N_21119);
nand U23469 (N_23469,N_20261,N_20816);
or U23470 (N_23470,N_20078,N_19894);
and U23471 (N_23471,N_19044,N_20083);
nor U23472 (N_23472,N_19113,N_21574);
nand U23473 (N_23473,N_19063,N_20174);
and U23474 (N_23474,N_21308,N_21434);
nor U23475 (N_23475,N_20126,N_20692);
nand U23476 (N_23476,N_20835,N_20633);
nor U23477 (N_23477,N_19348,N_20698);
nand U23478 (N_23478,N_19446,N_19045);
nor U23479 (N_23479,N_18778,N_19410);
or U23480 (N_23480,N_19379,N_19804);
nand U23481 (N_23481,N_20000,N_19473);
or U23482 (N_23482,N_20503,N_20498);
and U23483 (N_23483,N_21611,N_19763);
and U23484 (N_23484,N_20707,N_19328);
nor U23485 (N_23485,N_18872,N_21288);
or U23486 (N_23486,N_18774,N_20635);
nor U23487 (N_23487,N_20715,N_19868);
or U23488 (N_23488,N_21624,N_19272);
nor U23489 (N_23489,N_21430,N_20112);
and U23490 (N_23490,N_19041,N_19987);
nand U23491 (N_23491,N_20574,N_19678);
and U23492 (N_23492,N_20573,N_21065);
nor U23493 (N_23493,N_19266,N_19470);
and U23494 (N_23494,N_20537,N_18954);
xnor U23495 (N_23495,N_20483,N_20997);
nand U23496 (N_23496,N_19776,N_19749);
nand U23497 (N_23497,N_19896,N_20290);
or U23498 (N_23498,N_18980,N_20371);
and U23499 (N_23499,N_21806,N_19473);
nand U23500 (N_23500,N_20528,N_20706);
and U23501 (N_23501,N_20539,N_21242);
xnor U23502 (N_23502,N_21592,N_21819);
nor U23503 (N_23503,N_18968,N_21218);
xnor U23504 (N_23504,N_20955,N_21433);
nand U23505 (N_23505,N_19083,N_19610);
nor U23506 (N_23506,N_19970,N_19344);
nor U23507 (N_23507,N_19877,N_21196);
xnor U23508 (N_23508,N_18949,N_19893);
nor U23509 (N_23509,N_20667,N_18778);
nand U23510 (N_23510,N_20193,N_19942);
nand U23511 (N_23511,N_19805,N_19383);
nand U23512 (N_23512,N_20965,N_20761);
nor U23513 (N_23513,N_20084,N_21522);
and U23514 (N_23514,N_20771,N_19350);
xor U23515 (N_23515,N_21285,N_20788);
and U23516 (N_23516,N_19490,N_20206);
nand U23517 (N_23517,N_21191,N_21425);
nand U23518 (N_23518,N_19679,N_19094);
and U23519 (N_23519,N_21846,N_21190);
and U23520 (N_23520,N_19726,N_19618);
nand U23521 (N_23521,N_20528,N_19456);
or U23522 (N_23522,N_21716,N_19193);
or U23523 (N_23523,N_21002,N_21261);
and U23524 (N_23524,N_20261,N_19479);
nor U23525 (N_23525,N_20482,N_19511);
and U23526 (N_23526,N_21247,N_20999);
and U23527 (N_23527,N_19353,N_21053);
nor U23528 (N_23528,N_20742,N_19363);
nor U23529 (N_23529,N_20625,N_18874);
or U23530 (N_23530,N_19591,N_21775);
xnor U23531 (N_23531,N_19057,N_20348);
xnor U23532 (N_23532,N_20381,N_19182);
nor U23533 (N_23533,N_21831,N_19137);
and U23534 (N_23534,N_20027,N_19029);
and U23535 (N_23535,N_20682,N_21071);
nand U23536 (N_23536,N_20080,N_20607);
nand U23537 (N_23537,N_21000,N_20562);
or U23538 (N_23538,N_21464,N_19115);
and U23539 (N_23539,N_19375,N_20873);
xor U23540 (N_23540,N_21351,N_21584);
and U23541 (N_23541,N_21286,N_19550);
or U23542 (N_23542,N_19270,N_19555);
nand U23543 (N_23543,N_19206,N_20849);
and U23544 (N_23544,N_19081,N_20523);
nand U23545 (N_23545,N_19717,N_20021);
nor U23546 (N_23546,N_21458,N_20165);
or U23547 (N_23547,N_19603,N_20224);
nor U23548 (N_23548,N_21168,N_21152);
or U23549 (N_23549,N_20726,N_19943);
nand U23550 (N_23550,N_21078,N_19138);
nand U23551 (N_23551,N_19980,N_21615);
or U23552 (N_23552,N_20921,N_20663);
or U23553 (N_23553,N_19703,N_19662);
nand U23554 (N_23554,N_20560,N_19827);
or U23555 (N_23555,N_20757,N_19330);
and U23556 (N_23556,N_20719,N_21443);
nor U23557 (N_23557,N_19005,N_19601);
nand U23558 (N_23558,N_21786,N_20815);
nand U23559 (N_23559,N_18836,N_19878);
or U23560 (N_23560,N_21082,N_19449);
xnor U23561 (N_23561,N_21322,N_21083);
nor U23562 (N_23562,N_21856,N_21705);
xnor U23563 (N_23563,N_20007,N_20433);
and U23564 (N_23564,N_20406,N_19775);
and U23565 (N_23565,N_21105,N_20373);
nor U23566 (N_23566,N_20241,N_19876);
and U23567 (N_23567,N_20639,N_20280);
xnor U23568 (N_23568,N_18940,N_19557);
nor U23569 (N_23569,N_21806,N_19584);
and U23570 (N_23570,N_19695,N_19401);
or U23571 (N_23571,N_21137,N_21060);
and U23572 (N_23572,N_19360,N_20484);
xnor U23573 (N_23573,N_19210,N_19703);
nand U23574 (N_23574,N_19191,N_21729);
and U23575 (N_23575,N_21234,N_20804);
or U23576 (N_23576,N_19119,N_19442);
nor U23577 (N_23577,N_19724,N_20857);
nand U23578 (N_23578,N_20842,N_20664);
nor U23579 (N_23579,N_20499,N_20672);
nand U23580 (N_23580,N_21481,N_20139);
or U23581 (N_23581,N_20636,N_19253);
nand U23582 (N_23582,N_19105,N_19398);
or U23583 (N_23583,N_19446,N_19659);
or U23584 (N_23584,N_19956,N_21148);
nand U23585 (N_23585,N_21490,N_21043);
nand U23586 (N_23586,N_21167,N_20368);
or U23587 (N_23587,N_21845,N_19525);
nor U23588 (N_23588,N_21790,N_20786);
xor U23589 (N_23589,N_19746,N_20294);
nor U23590 (N_23590,N_20360,N_19476);
or U23591 (N_23591,N_20557,N_19891);
nor U23592 (N_23592,N_19491,N_20651);
nor U23593 (N_23593,N_20814,N_21206);
or U23594 (N_23594,N_21659,N_19543);
nor U23595 (N_23595,N_19934,N_21258);
or U23596 (N_23596,N_20922,N_21700);
and U23597 (N_23597,N_21291,N_21262);
and U23598 (N_23598,N_20890,N_20697);
nand U23599 (N_23599,N_19553,N_19849);
nand U23600 (N_23600,N_19075,N_20141);
nand U23601 (N_23601,N_20720,N_20061);
or U23602 (N_23602,N_19660,N_20264);
xor U23603 (N_23603,N_20153,N_20852);
or U23604 (N_23604,N_19934,N_19549);
or U23605 (N_23605,N_20436,N_21308);
nand U23606 (N_23606,N_20492,N_21386);
nor U23607 (N_23607,N_20691,N_19144);
and U23608 (N_23608,N_20064,N_20846);
nand U23609 (N_23609,N_19702,N_20579);
and U23610 (N_23610,N_20716,N_20491);
or U23611 (N_23611,N_21793,N_19067);
nor U23612 (N_23612,N_21239,N_20346);
and U23613 (N_23613,N_19642,N_18957);
and U23614 (N_23614,N_19261,N_19456);
or U23615 (N_23615,N_20303,N_19778);
nand U23616 (N_23616,N_20448,N_21459);
nand U23617 (N_23617,N_21281,N_19820);
nor U23618 (N_23618,N_21488,N_20748);
nand U23619 (N_23619,N_21297,N_21724);
xnor U23620 (N_23620,N_19957,N_20428);
and U23621 (N_23621,N_20937,N_20828);
nand U23622 (N_23622,N_20913,N_20731);
or U23623 (N_23623,N_21166,N_21344);
nor U23624 (N_23624,N_20260,N_21264);
nor U23625 (N_23625,N_21500,N_19528);
or U23626 (N_23626,N_21711,N_21220);
or U23627 (N_23627,N_19070,N_21822);
or U23628 (N_23628,N_20784,N_19927);
xor U23629 (N_23629,N_20888,N_20267);
and U23630 (N_23630,N_20323,N_18863);
or U23631 (N_23631,N_19955,N_20034);
nand U23632 (N_23632,N_21702,N_19984);
xnor U23633 (N_23633,N_20529,N_21273);
nor U23634 (N_23634,N_20848,N_18898);
or U23635 (N_23635,N_20106,N_20950);
and U23636 (N_23636,N_20714,N_19468);
or U23637 (N_23637,N_19045,N_20972);
or U23638 (N_23638,N_20485,N_20274);
or U23639 (N_23639,N_19722,N_20331);
or U23640 (N_23640,N_20965,N_20716);
and U23641 (N_23641,N_20965,N_19368);
nor U23642 (N_23642,N_21414,N_19878);
nor U23643 (N_23643,N_18947,N_21256);
nor U23644 (N_23644,N_19672,N_19624);
or U23645 (N_23645,N_19099,N_20591);
nor U23646 (N_23646,N_20545,N_20116);
or U23647 (N_23647,N_19298,N_20759);
nor U23648 (N_23648,N_20095,N_20765);
nand U23649 (N_23649,N_18945,N_19492);
and U23650 (N_23650,N_18850,N_19724);
nand U23651 (N_23651,N_21411,N_19052);
and U23652 (N_23652,N_19343,N_21512);
xor U23653 (N_23653,N_19733,N_21330);
xnor U23654 (N_23654,N_20195,N_20934);
nor U23655 (N_23655,N_21245,N_20381);
and U23656 (N_23656,N_21185,N_21799);
or U23657 (N_23657,N_20173,N_21644);
nand U23658 (N_23658,N_20634,N_21833);
nor U23659 (N_23659,N_19787,N_20037);
xor U23660 (N_23660,N_20525,N_19445);
nor U23661 (N_23661,N_20281,N_20447);
and U23662 (N_23662,N_20507,N_19197);
nand U23663 (N_23663,N_21112,N_20387);
and U23664 (N_23664,N_19155,N_20559);
or U23665 (N_23665,N_21105,N_20985);
or U23666 (N_23666,N_20333,N_20027);
and U23667 (N_23667,N_19181,N_21857);
and U23668 (N_23668,N_20548,N_19060);
or U23669 (N_23669,N_20196,N_19253);
nand U23670 (N_23670,N_20214,N_21693);
and U23671 (N_23671,N_20011,N_19378);
nor U23672 (N_23672,N_19884,N_20612);
or U23673 (N_23673,N_20367,N_19013);
xor U23674 (N_23674,N_19747,N_21659);
or U23675 (N_23675,N_20040,N_20817);
xor U23676 (N_23676,N_20870,N_21700);
or U23677 (N_23677,N_18977,N_19792);
nor U23678 (N_23678,N_21264,N_20679);
nand U23679 (N_23679,N_19626,N_20013);
or U23680 (N_23680,N_19737,N_21576);
nand U23681 (N_23681,N_19159,N_20046);
nand U23682 (N_23682,N_20947,N_20061);
xor U23683 (N_23683,N_19068,N_19555);
and U23684 (N_23684,N_19066,N_19154);
nor U23685 (N_23685,N_19694,N_19987);
or U23686 (N_23686,N_20304,N_19510);
and U23687 (N_23687,N_19335,N_21016);
nand U23688 (N_23688,N_20273,N_21114);
or U23689 (N_23689,N_21496,N_19718);
nand U23690 (N_23690,N_19762,N_21838);
nand U23691 (N_23691,N_21740,N_18949);
and U23692 (N_23692,N_18988,N_21561);
or U23693 (N_23693,N_20291,N_18798);
nor U23694 (N_23694,N_19626,N_19715);
or U23695 (N_23695,N_18855,N_19689);
nor U23696 (N_23696,N_18907,N_20930);
xnor U23697 (N_23697,N_19122,N_20714);
nor U23698 (N_23698,N_20827,N_21376);
nor U23699 (N_23699,N_20597,N_19913);
nand U23700 (N_23700,N_20664,N_21755);
and U23701 (N_23701,N_20270,N_19996);
and U23702 (N_23702,N_20153,N_21737);
nand U23703 (N_23703,N_21582,N_20175);
nor U23704 (N_23704,N_19926,N_19711);
and U23705 (N_23705,N_19129,N_20823);
or U23706 (N_23706,N_19135,N_20300);
and U23707 (N_23707,N_20591,N_19339);
and U23708 (N_23708,N_21471,N_19921);
and U23709 (N_23709,N_21335,N_21400);
nor U23710 (N_23710,N_20538,N_19013);
and U23711 (N_23711,N_19535,N_19286);
or U23712 (N_23712,N_20961,N_20113);
xnor U23713 (N_23713,N_20300,N_20082);
or U23714 (N_23714,N_21313,N_20428);
and U23715 (N_23715,N_21652,N_20261);
xnor U23716 (N_23716,N_19836,N_21721);
nand U23717 (N_23717,N_19818,N_21097);
nor U23718 (N_23718,N_18890,N_19989);
nor U23719 (N_23719,N_21254,N_20832);
and U23720 (N_23720,N_21384,N_19739);
nand U23721 (N_23721,N_21031,N_20513);
or U23722 (N_23722,N_21277,N_18989);
nand U23723 (N_23723,N_19543,N_19983);
nor U23724 (N_23724,N_20737,N_20680);
nor U23725 (N_23725,N_20299,N_20328);
nand U23726 (N_23726,N_19585,N_19253);
or U23727 (N_23727,N_21858,N_21455);
nand U23728 (N_23728,N_21364,N_19684);
nand U23729 (N_23729,N_20553,N_21156);
xnor U23730 (N_23730,N_20731,N_21128);
nand U23731 (N_23731,N_21748,N_19458);
nor U23732 (N_23732,N_20771,N_21289);
nand U23733 (N_23733,N_20078,N_18838);
and U23734 (N_23734,N_18795,N_20383);
nor U23735 (N_23735,N_20792,N_21261);
nand U23736 (N_23736,N_21871,N_19759);
or U23737 (N_23737,N_19873,N_20345);
nor U23738 (N_23738,N_19689,N_21700);
or U23739 (N_23739,N_21478,N_19214);
and U23740 (N_23740,N_21519,N_20476);
nor U23741 (N_23741,N_20835,N_21342);
nand U23742 (N_23742,N_21316,N_21874);
and U23743 (N_23743,N_20976,N_20645);
nand U23744 (N_23744,N_20289,N_21209);
nand U23745 (N_23745,N_21464,N_20277);
nand U23746 (N_23746,N_20834,N_21800);
nor U23747 (N_23747,N_21871,N_21016);
xor U23748 (N_23748,N_21005,N_19955);
nand U23749 (N_23749,N_20319,N_19301);
and U23750 (N_23750,N_19497,N_21682);
nor U23751 (N_23751,N_21218,N_19096);
or U23752 (N_23752,N_21523,N_21258);
nor U23753 (N_23753,N_18899,N_19471);
and U23754 (N_23754,N_20747,N_20969);
nand U23755 (N_23755,N_19846,N_19955);
nor U23756 (N_23756,N_18937,N_21161);
and U23757 (N_23757,N_19453,N_19487);
and U23758 (N_23758,N_20580,N_19608);
nand U23759 (N_23759,N_21556,N_21747);
or U23760 (N_23760,N_20326,N_19478);
nand U23761 (N_23761,N_19332,N_19502);
xor U23762 (N_23762,N_21519,N_19544);
or U23763 (N_23763,N_21568,N_21862);
xnor U23764 (N_23764,N_19197,N_18970);
nand U23765 (N_23765,N_19752,N_21752);
nand U23766 (N_23766,N_20002,N_19089);
or U23767 (N_23767,N_21830,N_21808);
or U23768 (N_23768,N_21354,N_19275);
or U23769 (N_23769,N_19856,N_19908);
and U23770 (N_23770,N_20508,N_20873);
or U23771 (N_23771,N_20515,N_20107);
nor U23772 (N_23772,N_20841,N_21669);
and U23773 (N_23773,N_20120,N_20788);
nand U23774 (N_23774,N_19892,N_20851);
or U23775 (N_23775,N_18920,N_20307);
nand U23776 (N_23776,N_20813,N_21356);
or U23777 (N_23777,N_20661,N_19081);
nand U23778 (N_23778,N_21388,N_19133);
nor U23779 (N_23779,N_21791,N_20862);
nand U23780 (N_23780,N_20086,N_19564);
and U23781 (N_23781,N_21565,N_20913);
nor U23782 (N_23782,N_19063,N_19353);
and U23783 (N_23783,N_19681,N_21202);
nor U23784 (N_23784,N_19697,N_19988);
or U23785 (N_23785,N_18825,N_20976);
and U23786 (N_23786,N_20922,N_18752);
or U23787 (N_23787,N_20177,N_19456);
nor U23788 (N_23788,N_21776,N_19072);
nand U23789 (N_23789,N_20075,N_18954);
nor U23790 (N_23790,N_20500,N_19610);
nor U23791 (N_23791,N_19892,N_20208);
or U23792 (N_23792,N_19506,N_21148);
or U23793 (N_23793,N_21682,N_21819);
nand U23794 (N_23794,N_19790,N_19545);
and U23795 (N_23795,N_20637,N_21407);
or U23796 (N_23796,N_18947,N_21840);
xnor U23797 (N_23797,N_18780,N_21135);
or U23798 (N_23798,N_19659,N_20536);
or U23799 (N_23799,N_18873,N_20771);
nor U23800 (N_23800,N_20643,N_19048);
nand U23801 (N_23801,N_21070,N_19478);
and U23802 (N_23802,N_18760,N_19376);
or U23803 (N_23803,N_21032,N_19005);
nor U23804 (N_23804,N_21426,N_19766);
nor U23805 (N_23805,N_19642,N_18854);
xnor U23806 (N_23806,N_20467,N_20428);
xnor U23807 (N_23807,N_19318,N_19045);
xor U23808 (N_23808,N_21674,N_19909);
nor U23809 (N_23809,N_20208,N_20857);
and U23810 (N_23810,N_21210,N_18770);
xnor U23811 (N_23811,N_19798,N_19738);
and U23812 (N_23812,N_21475,N_19899);
or U23813 (N_23813,N_20410,N_19936);
and U23814 (N_23814,N_20929,N_21870);
nand U23815 (N_23815,N_21041,N_20750);
or U23816 (N_23816,N_19816,N_18882);
nor U23817 (N_23817,N_19315,N_19467);
and U23818 (N_23818,N_20949,N_21838);
nand U23819 (N_23819,N_21838,N_18945);
nor U23820 (N_23820,N_18772,N_20539);
or U23821 (N_23821,N_19255,N_20079);
xnor U23822 (N_23822,N_19517,N_21507);
or U23823 (N_23823,N_21348,N_18803);
nand U23824 (N_23824,N_18753,N_20615);
and U23825 (N_23825,N_20667,N_21511);
and U23826 (N_23826,N_20369,N_20740);
nand U23827 (N_23827,N_20482,N_20893);
nor U23828 (N_23828,N_19787,N_20425);
and U23829 (N_23829,N_20639,N_19160);
and U23830 (N_23830,N_19789,N_20970);
and U23831 (N_23831,N_20515,N_19926);
and U23832 (N_23832,N_20723,N_21461);
or U23833 (N_23833,N_19984,N_19835);
nand U23834 (N_23834,N_19918,N_20072);
nor U23835 (N_23835,N_19383,N_20998);
or U23836 (N_23836,N_21353,N_20316);
nand U23837 (N_23837,N_20810,N_21173);
nor U23838 (N_23838,N_20896,N_19479);
nor U23839 (N_23839,N_21365,N_21000);
nand U23840 (N_23840,N_19227,N_19308);
nand U23841 (N_23841,N_21762,N_21656);
and U23842 (N_23842,N_19909,N_19051);
or U23843 (N_23843,N_19640,N_19563);
xnor U23844 (N_23844,N_19261,N_20365);
nand U23845 (N_23845,N_21010,N_21739);
nor U23846 (N_23846,N_18860,N_19097);
nor U23847 (N_23847,N_20042,N_20620);
nand U23848 (N_23848,N_21031,N_18954);
and U23849 (N_23849,N_21795,N_19177);
and U23850 (N_23850,N_21423,N_21069);
or U23851 (N_23851,N_19930,N_20190);
nor U23852 (N_23852,N_21266,N_21327);
nor U23853 (N_23853,N_19737,N_19095);
and U23854 (N_23854,N_19641,N_20571);
or U23855 (N_23855,N_20619,N_19761);
or U23856 (N_23856,N_21681,N_20550);
nor U23857 (N_23857,N_20449,N_20584);
xnor U23858 (N_23858,N_19119,N_19497);
nand U23859 (N_23859,N_20843,N_20174);
nor U23860 (N_23860,N_19704,N_21391);
or U23861 (N_23861,N_20519,N_21282);
xor U23862 (N_23862,N_21870,N_19011);
nand U23863 (N_23863,N_20841,N_19133);
nor U23864 (N_23864,N_20024,N_20577);
nand U23865 (N_23865,N_18804,N_20509);
nand U23866 (N_23866,N_19382,N_21055);
or U23867 (N_23867,N_20148,N_21792);
nand U23868 (N_23868,N_21614,N_20612);
nand U23869 (N_23869,N_21477,N_20256);
and U23870 (N_23870,N_20717,N_21260);
nor U23871 (N_23871,N_21034,N_19121);
nor U23872 (N_23872,N_20028,N_19946);
or U23873 (N_23873,N_19655,N_19152);
xor U23874 (N_23874,N_21445,N_20005);
and U23875 (N_23875,N_20561,N_20317);
nor U23876 (N_23876,N_20041,N_20579);
or U23877 (N_23877,N_20320,N_19224);
and U23878 (N_23878,N_19604,N_19466);
and U23879 (N_23879,N_20962,N_18935);
nand U23880 (N_23880,N_20747,N_19646);
and U23881 (N_23881,N_19182,N_20225);
or U23882 (N_23882,N_19934,N_20776);
or U23883 (N_23883,N_20024,N_19824);
nor U23884 (N_23884,N_20772,N_20207);
nor U23885 (N_23885,N_19109,N_18804);
or U23886 (N_23886,N_21530,N_20180);
and U23887 (N_23887,N_19221,N_20307);
or U23888 (N_23888,N_20500,N_19656);
nor U23889 (N_23889,N_20051,N_21255);
nor U23890 (N_23890,N_21223,N_21862);
nand U23891 (N_23891,N_20640,N_20959);
nand U23892 (N_23892,N_19236,N_20668);
nor U23893 (N_23893,N_21070,N_19726);
and U23894 (N_23894,N_19986,N_19607);
or U23895 (N_23895,N_20596,N_19816);
and U23896 (N_23896,N_19857,N_19540);
nand U23897 (N_23897,N_20351,N_19672);
and U23898 (N_23898,N_19568,N_21782);
and U23899 (N_23899,N_21687,N_21599);
and U23900 (N_23900,N_20935,N_21233);
nand U23901 (N_23901,N_21594,N_19552);
or U23902 (N_23902,N_19258,N_18988);
and U23903 (N_23903,N_21043,N_21711);
or U23904 (N_23904,N_19505,N_19154);
nand U23905 (N_23905,N_21846,N_20437);
or U23906 (N_23906,N_19201,N_21853);
and U23907 (N_23907,N_20345,N_20748);
nand U23908 (N_23908,N_19762,N_18777);
nor U23909 (N_23909,N_21568,N_19895);
nand U23910 (N_23910,N_19767,N_19535);
nor U23911 (N_23911,N_21574,N_20003);
xnor U23912 (N_23912,N_21081,N_19604);
and U23913 (N_23913,N_21862,N_19169);
xnor U23914 (N_23914,N_20825,N_19022);
xnor U23915 (N_23915,N_19863,N_19918);
and U23916 (N_23916,N_19571,N_21747);
or U23917 (N_23917,N_18824,N_20352);
nand U23918 (N_23918,N_18962,N_21815);
nand U23919 (N_23919,N_19564,N_20920);
and U23920 (N_23920,N_21204,N_20647);
and U23921 (N_23921,N_18933,N_21637);
nand U23922 (N_23922,N_21008,N_20316);
or U23923 (N_23923,N_21840,N_20963);
nand U23924 (N_23924,N_20472,N_18949);
and U23925 (N_23925,N_21560,N_19125);
xor U23926 (N_23926,N_20048,N_21605);
or U23927 (N_23927,N_19141,N_20311);
and U23928 (N_23928,N_20261,N_19348);
nor U23929 (N_23929,N_19814,N_21424);
nand U23930 (N_23930,N_19204,N_21715);
nor U23931 (N_23931,N_19614,N_19659);
nand U23932 (N_23932,N_21034,N_20794);
or U23933 (N_23933,N_21023,N_21510);
or U23934 (N_23934,N_19232,N_20555);
nor U23935 (N_23935,N_19558,N_19663);
nand U23936 (N_23936,N_21147,N_20654);
or U23937 (N_23937,N_20564,N_19712);
nor U23938 (N_23938,N_21280,N_21041);
nand U23939 (N_23939,N_20096,N_20253);
nor U23940 (N_23940,N_20851,N_20099);
nor U23941 (N_23941,N_20148,N_19099);
and U23942 (N_23942,N_20669,N_21733);
and U23943 (N_23943,N_21674,N_20324);
nor U23944 (N_23944,N_20673,N_19443);
and U23945 (N_23945,N_21116,N_20128);
and U23946 (N_23946,N_19250,N_20646);
nor U23947 (N_23947,N_20918,N_20406);
or U23948 (N_23948,N_21099,N_21082);
nor U23949 (N_23949,N_21115,N_20459);
and U23950 (N_23950,N_19454,N_21157);
nand U23951 (N_23951,N_19128,N_20562);
nand U23952 (N_23952,N_21662,N_20290);
nand U23953 (N_23953,N_20250,N_21545);
xnor U23954 (N_23954,N_21533,N_20891);
or U23955 (N_23955,N_20172,N_18964);
nand U23956 (N_23956,N_21465,N_19754);
and U23957 (N_23957,N_21342,N_21750);
nor U23958 (N_23958,N_21012,N_19271);
nor U23959 (N_23959,N_19381,N_21839);
xor U23960 (N_23960,N_19051,N_21213);
or U23961 (N_23961,N_21382,N_20458);
or U23962 (N_23962,N_21486,N_18780);
nor U23963 (N_23963,N_18883,N_21012);
nand U23964 (N_23964,N_20078,N_20754);
xor U23965 (N_23965,N_19738,N_21746);
or U23966 (N_23966,N_21345,N_21815);
and U23967 (N_23967,N_19904,N_21712);
nand U23968 (N_23968,N_21137,N_21417);
nand U23969 (N_23969,N_21397,N_19529);
xnor U23970 (N_23970,N_20507,N_20376);
or U23971 (N_23971,N_19753,N_20139);
and U23972 (N_23972,N_18792,N_19196);
nor U23973 (N_23973,N_20394,N_20272);
and U23974 (N_23974,N_19680,N_21043);
or U23975 (N_23975,N_20045,N_20229);
or U23976 (N_23976,N_19491,N_20470);
and U23977 (N_23977,N_20454,N_18754);
nor U23978 (N_23978,N_18837,N_21530);
nor U23979 (N_23979,N_20934,N_20964);
or U23980 (N_23980,N_21794,N_19784);
nand U23981 (N_23981,N_20406,N_19818);
nand U23982 (N_23982,N_20860,N_19361);
xor U23983 (N_23983,N_21591,N_19004);
nor U23984 (N_23984,N_19968,N_20071);
nor U23985 (N_23985,N_18900,N_18956);
and U23986 (N_23986,N_19884,N_20573);
xnor U23987 (N_23987,N_20493,N_19363);
nand U23988 (N_23988,N_19631,N_19377);
or U23989 (N_23989,N_20881,N_21447);
xor U23990 (N_23990,N_20610,N_19470);
xnor U23991 (N_23991,N_19578,N_18770);
xnor U23992 (N_23992,N_19824,N_20786);
or U23993 (N_23993,N_19927,N_19972);
or U23994 (N_23994,N_19897,N_21078);
and U23995 (N_23995,N_21479,N_20414);
nor U23996 (N_23996,N_19422,N_21389);
and U23997 (N_23997,N_20204,N_20088);
and U23998 (N_23998,N_21059,N_19445);
and U23999 (N_23999,N_21859,N_21326);
nand U24000 (N_24000,N_20198,N_19080);
nand U24001 (N_24001,N_19186,N_20213);
nor U24002 (N_24002,N_20659,N_21744);
nand U24003 (N_24003,N_21641,N_20046);
nor U24004 (N_24004,N_18966,N_20038);
or U24005 (N_24005,N_19883,N_20005);
or U24006 (N_24006,N_18807,N_21159);
xor U24007 (N_24007,N_20884,N_19879);
and U24008 (N_24008,N_20341,N_20228);
nand U24009 (N_24009,N_20067,N_19417);
nor U24010 (N_24010,N_19151,N_20996);
or U24011 (N_24011,N_19908,N_19727);
nor U24012 (N_24012,N_19308,N_19870);
and U24013 (N_24013,N_20377,N_19194);
nor U24014 (N_24014,N_21528,N_19723);
and U24015 (N_24015,N_18872,N_19541);
xnor U24016 (N_24016,N_20358,N_21484);
nand U24017 (N_24017,N_20254,N_20608);
nor U24018 (N_24018,N_19085,N_18819);
and U24019 (N_24019,N_19758,N_21409);
and U24020 (N_24020,N_21657,N_18791);
and U24021 (N_24021,N_20120,N_20104);
nor U24022 (N_24022,N_21793,N_20790);
nand U24023 (N_24023,N_21840,N_19701);
nor U24024 (N_24024,N_19284,N_21108);
and U24025 (N_24025,N_19019,N_19014);
or U24026 (N_24026,N_19234,N_19460);
and U24027 (N_24027,N_20059,N_20540);
nor U24028 (N_24028,N_18885,N_21026);
nor U24029 (N_24029,N_19194,N_20957);
and U24030 (N_24030,N_20994,N_18919);
or U24031 (N_24031,N_21085,N_21031);
nand U24032 (N_24032,N_21028,N_21179);
nand U24033 (N_24033,N_20878,N_18918);
nor U24034 (N_24034,N_19208,N_19047);
and U24035 (N_24035,N_20231,N_20749);
and U24036 (N_24036,N_20473,N_20200);
xnor U24037 (N_24037,N_21295,N_20100);
or U24038 (N_24038,N_19157,N_20155);
nor U24039 (N_24039,N_20018,N_18880);
or U24040 (N_24040,N_21494,N_21832);
and U24041 (N_24041,N_21320,N_19582);
nand U24042 (N_24042,N_20491,N_20849);
xor U24043 (N_24043,N_19939,N_19181);
or U24044 (N_24044,N_21737,N_21219);
or U24045 (N_24045,N_19041,N_21785);
or U24046 (N_24046,N_19294,N_19599);
nor U24047 (N_24047,N_21331,N_19042);
nand U24048 (N_24048,N_21728,N_21236);
nand U24049 (N_24049,N_20053,N_21456);
or U24050 (N_24050,N_19277,N_19790);
or U24051 (N_24051,N_19825,N_21385);
nor U24052 (N_24052,N_19869,N_19001);
and U24053 (N_24053,N_19105,N_19301);
or U24054 (N_24054,N_19166,N_20506);
nor U24055 (N_24055,N_19203,N_19335);
or U24056 (N_24056,N_19819,N_19649);
nand U24057 (N_24057,N_21536,N_19561);
and U24058 (N_24058,N_21787,N_19035);
nor U24059 (N_24059,N_18813,N_19640);
xor U24060 (N_24060,N_20696,N_20552);
nand U24061 (N_24061,N_21855,N_21787);
or U24062 (N_24062,N_21539,N_18851);
nand U24063 (N_24063,N_20600,N_20434);
or U24064 (N_24064,N_19462,N_19643);
or U24065 (N_24065,N_19592,N_21858);
or U24066 (N_24066,N_20225,N_19549);
or U24067 (N_24067,N_21504,N_20753);
and U24068 (N_24068,N_19563,N_21311);
nand U24069 (N_24069,N_18752,N_20278);
nand U24070 (N_24070,N_19829,N_20565);
or U24071 (N_24071,N_19757,N_21093);
nand U24072 (N_24072,N_19286,N_20553);
and U24073 (N_24073,N_19135,N_21420);
nand U24074 (N_24074,N_19414,N_21862);
and U24075 (N_24075,N_20226,N_21542);
or U24076 (N_24076,N_21432,N_19998);
nor U24077 (N_24077,N_19134,N_20955);
and U24078 (N_24078,N_19329,N_21631);
nand U24079 (N_24079,N_18852,N_20622);
nand U24080 (N_24080,N_20119,N_19071);
nor U24081 (N_24081,N_19532,N_20068);
and U24082 (N_24082,N_21294,N_19189);
and U24083 (N_24083,N_20757,N_20019);
or U24084 (N_24084,N_20652,N_21024);
nor U24085 (N_24085,N_19797,N_20917);
and U24086 (N_24086,N_20536,N_19313);
and U24087 (N_24087,N_21149,N_19056);
xor U24088 (N_24088,N_20688,N_21866);
or U24089 (N_24089,N_21696,N_21715);
and U24090 (N_24090,N_18851,N_19541);
and U24091 (N_24091,N_19398,N_19731);
or U24092 (N_24092,N_19180,N_19320);
and U24093 (N_24093,N_20933,N_19544);
or U24094 (N_24094,N_20466,N_19636);
nand U24095 (N_24095,N_19755,N_19856);
nor U24096 (N_24096,N_18886,N_19127);
and U24097 (N_24097,N_19979,N_20512);
nor U24098 (N_24098,N_20069,N_19597);
and U24099 (N_24099,N_19189,N_19963);
nor U24100 (N_24100,N_19363,N_20285);
nand U24101 (N_24101,N_19090,N_20000);
nor U24102 (N_24102,N_21821,N_21574);
nor U24103 (N_24103,N_18960,N_20783);
or U24104 (N_24104,N_20531,N_20155);
or U24105 (N_24105,N_21508,N_19438);
and U24106 (N_24106,N_21537,N_21868);
nor U24107 (N_24107,N_21377,N_19139);
or U24108 (N_24108,N_21492,N_20304);
and U24109 (N_24109,N_21797,N_19850);
nor U24110 (N_24110,N_19926,N_19769);
nand U24111 (N_24111,N_20515,N_19671);
nor U24112 (N_24112,N_20497,N_20634);
xnor U24113 (N_24113,N_20274,N_19093);
nand U24114 (N_24114,N_20731,N_19682);
or U24115 (N_24115,N_20136,N_20705);
xor U24116 (N_24116,N_19422,N_20022);
nor U24117 (N_24117,N_18753,N_20119);
or U24118 (N_24118,N_20603,N_20324);
or U24119 (N_24119,N_18960,N_19975);
nand U24120 (N_24120,N_19070,N_20556);
nor U24121 (N_24121,N_20886,N_18974);
nand U24122 (N_24122,N_21322,N_19050);
and U24123 (N_24123,N_20353,N_21771);
or U24124 (N_24124,N_18992,N_21178);
or U24125 (N_24125,N_20472,N_18889);
nand U24126 (N_24126,N_20380,N_19744);
nor U24127 (N_24127,N_21351,N_19962);
nor U24128 (N_24128,N_19443,N_19426);
and U24129 (N_24129,N_20254,N_21726);
and U24130 (N_24130,N_21660,N_21087);
xor U24131 (N_24131,N_21236,N_18964);
nand U24132 (N_24132,N_19996,N_21195);
nand U24133 (N_24133,N_19030,N_19750);
and U24134 (N_24134,N_18839,N_19285);
nor U24135 (N_24135,N_19769,N_19993);
nand U24136 (N_24136,N_18928,N_21137);
or U24137 (N_24137,N_20950,N_21031);
nand U24138 (N_24138,N_19775,N_21544);
nand U24139 (N_24139,N_19655,N_20062);
nor U24140 (N_24140,N_19001,N_19861);
and U24141 (N_24141,N_20063,N_18832);
or U24142 (N_24142,N_21575,N_20615);
or U24143 (N_24143,N_18845,N_19524);
nor U24144 (N_24144,N_21166,N_20272);
nor U24145 (N_24145,N_21625,N_20059);
xnor U24146 (N_24146,N_19568,N_20425);
nand U24147 (N_24147,N_21583,N_19153);
and U24148 (N_24148,N_18803,N_20274);
or U24149 (N_24149,N_21409,N_20247);
or U24150 (N_24150,N_19816,N_20423);
or U24151 (N_24151,N_19588,N_19897);
nor U24152 (N_24152,N_21239,N_19345);
nand U24153 (N_24153,N_21840,N_21435);
and U24154 (N_24154,N_20584,N_20474);
nand U24155 (N_24155,N_20487,N_21258);
nor U24156 (N_24156,N_21221,N_19145);
or U24157 (N_24157,N_19666,N_20586);
xor U24158 (N_24158,N_20309,N_19942);
nand U24159 (N_24159,N_21836,N_20474);
nand U24160 (N_24160,N_21064,N_20410);
xor U24161 (N_24161,N_20408,N_19718);
and U24162 (N_24162,N_21831,N_19024);
nand U24163 (N_24163,N_19433,N_20072);
and U24164 (N_24164,N_20204,N_19878);
and U24165 (N_24165,N_19110,N_20791);
nor U24166 (N_24166,N_20045,N_21183);
nand U24167 (N_24167,N_20574,N_21683);
and U24168 (N_24168,N_21808,N_20084);
nand U24169 (N_24169,N_19613,N_19124);
xnor U24170 (N_24170,N_19376,N_19605);
and U24171 (N_24171,N_19334,N_21612);
or U24172 (N_24172,N_19032,N_20228);
nand U24173 (N_24173,N_21688,N_20803);
nand U24174 (N_24174,N_21770,N_21362);
or U24175 (N_24175,N_19580,N_21233);
and U24176 (N_24176,N_19676,N_20527);
nor U24177 (N_24177,N_21249,N_20832);
xnor U24178 (N_24178,N_20924,N_19464);
and U24179 (N_24179,N_19928,N_19926);
and U24180 (N_24180,N_20742,N_21206);
and U24181 (N_24181,N_19973,N_21105);
nor U24182 (N_24182,N_19284,N_20183);
nor U24183 (N_24183,N_20515,N_21450);
and U24184 (N_24184,N_19815,N_20927);
or U24185 (N_24185,N_19131,N_21233);
or U24186 (N_24186,N_19473,N_21187);
nor U24187 (N_24187,N_21019,N_20622);
nor U24188 (N_24188,N_21155,N_19269);
xor U24189 (N_24189,N_21346,N_20642);
nand U24190 (N_24190,N_20966,N_20796);
or U24191 (N_24191,N_20657,N_21089);
or U24192 (N_24192,N_19120,N_20415);
and U24193 (N_24193,N_20815,N_19035);
nand U24194 (N_24194,N_20419,N_21392);
nor U24195 (N_24195,N_19977,N_19425);
and U24196 (N_24196,N_21718,N_19587);
nand U24197 (N_24197,N_18887,N_20353);
xnor U24198 (N_24198,N_18940,N_21083);
nor U24199 (N_24199,N_19322,N_20076);
nand U24200 (N_24200,N_18939,N_19699);
nand U24201 (N_24201,N_19896,N_20446);
nand U24202 (N_24202,N_21517,N_19452);
and U24203 (N_24203,N_20120,N_21599);
nor U24204 (N_24204,N_20288,N_21796);
or U24205 (N_24205,N_21200,N_19652);
nand U24206 (N_24206,N_21213,N_20350);
nand U24207 (N_24207,N_21399,N_19386);
nand U24208 (N_24208,N_19628,N_19698);
nand U24209 (N_24209,N_20539,N_21318);
or U24210 (N_24210,N_19482,N_21738);
nor U24211 (N_24211,N_19282,N_20257);
nand U24212 (N_24212,N_19547,N_20780);
and U24213 (N_24213,N_19186,N_21515);
or U24214 (N_24214,N_20843,N_21243);
nor U24215 (N_24215,N_20127,N_20653);
and U24216 (N_24216,N_21000,N_20585);
nand U24217 (N_24217,N_21552,N_20014);
xor U24218 (N_24218,N_18857,N_18995);
or U24219 (N_24219,N_21333,N_21789);
or U24220 (N_24220,N_19602,N_19984);
nand U24221 (N_24221,N_20616,N_21640);
and U24222 (N_24222,N_20608,N_19952);
and U24223 (N_24223,N_19817,N_20684);
or U24224 (N_24224,N_19130,N_18818);
or U24225 (N_24225,N_19122,N_20826);
nor U24226 (N_24226,N_20157,N_19994);
and U24227 (N_24227,N_19818,N_19882);
nand U24228 (N_24228,N_19515,N_21480);
and U24229 (N_24229,N_19347,N_20460);
nand U24230 (N_24230,N_18986,N_19575);
nand U24231 (N_24231,N_19510,N_21661);
or U24232 (N_24232,N_18827,N_21549);
nand U24233 (N_24233,N_21277,N_21596);
or U24234 (N_24234,N_19653,N_18768);
or U24235 (N_24235,N_19879,N_18795);
and U24236 (N_24236,N_20767,N_21561);
or U24237 (N_24237,N_21427,N_19285);
nor U24238 (N_24238,N_19595,N_20779);
or U24239 (N_24239,N_21549,N_21324);
or U24240 (N_24240,N_19464,N_20538);
or U24241 (N_24241,N_20936,N_19988);
nand U24242 (N_24242,N_19667,N_18937);
nand U24243 (N_24243,N_18955,N_19080);
nor U24244 (N_24244,N_19852,N_19834);
nor U24245 (N_24245,N_19430,N_21818);
nand U24246 (N_24246,N_19719,N_19673);
nand U24247 (N_24247,N_19953,N_18795);
or U24248 (N_24248,N_20856,N_18809);
nand U24249 (N_24249,N_21867,N_20933);
and U24250 (N_24250,N_19878,N_20578);
xnor U24251 (N_24251,N_20051,N_19448);
nand U24252 (N_24252,N_20105,N_20370);
nor U24253 (N_24253,N_21661,N_19030);
or U24254 (N_24254,N_21438,N_21109);
xor U24255 (N_24255,N_21612,N_19308);
nor U24256 (N_24256,N_21356,N_20823);
and U24257 (N_24257,N_19113,N_20367);
nor U24258 (N_24258,N_18958,N_21298);
nor U24259 (N_24259,N_20927,N_19107);
and U24260 (N_24260,N_21786,N_19169);
and U24261 (N_24261,N_20336,N_18790);
nor U24262 (N_24262,N_19240,N_19547);
or U24263 (N_24263,N_20756,N_19211);
nor U24264 (N_24264,N_20406,N_21284);
nor U24265 (N_24265,N_20849,N_19982);
nand U24266 (N_24266,N_21070,N_21453);
nor U24267 (N_24267,N_21658,N_19604);
nor U24268 (N_24268,N_20384,N_20943);
and U24269 (N_24269,N_18838,N_19732);
or U24270 (N_24270,N_19348,N_21048);
and U24271 (N_24271,N_20056,N_19358);
xor U24272 (N_24272,N_21190,N_21723);
nand U24273 (N_24273,N_21446,N_19184);
and U24274 (N_24274,N_21628,N_21076);
nor U24275 (N_24275,N_21542,N_20498);
nand U24276 (N_24276,N_19486,N_20715);
nand U24277 (N_24277,N_19431,N_21334);
nor U24278 (N_24278,N_19741,N_19125);
or U24279 (N_24279,N_19103,N_20228);
and U24280 (N_24280,N_19376,N_18977);
or U24281 (N_24281,N_21186,N_18991);
or U24282 (N_24282,N_19894,N_20184);
nand U24283 (N_24283,N_21808,N_19097);
nand U24284 (N_24284,N_21236,N_21520);
xnor U24285 (N_24285,N_18869,N_21801);
or U24286 (N_24286,N_21112,N_19395);
and U24287 (N_24287,N_19248,N_20823);
nor U24288 (N_24288,N_19396,N_21609);
nor U24289 (N_24289,N_20467,N_20271);
and U24290 (N_24290,N_19554,N_20372);
xor U24291 (N_24291,N_18918,N_21378);
nand U24292 (N_24292,N_21210,N_18805);
xnor U24293 (N_24293,N_20749,N_21298);
or U24294 (N_24294,N_21037,N_19967);
nor U24295 (N_24295,N_20119,N_19568);
xor U24296 (N_24296,N_20913,N_19670);
nor U24297 (N_24297,N_21327,N_21679);
nand U24298 (N_24298,N_20544,N_19337);
nand U24299 (N_24299,N_19197,N_20536);
or U24300 (N_24300,N_18954,N_19424);
and U24301 (N_24301,N_18796,N_19257);
xnor U24302 (N_24302,N_21387,N_19885);
nor U24303 (N_24303,N_19486,N_21629);
nand U24304 (N_24304,N_20947,N_21503);
and U24305 (N_24305,N_19881,N_20520);
nor U24306 (N_24306,N_20711,N_20032);
and U24307 (N_24307,N_21074,N_20877);
nand U24308 (N_24308,N_21297,N_21261);
or U24309 (N_24309,N_21586,N_20680);
or U24310 (N_24310,N_20282,N_18971);
or U24311 (N_24311,N_20075,N_21429);
nor U24312 (N_24312,N_21009,N_20002);
or U24313 (N_24313,N_19627,N_20640);
nand U24314 (N_24314,N_19121,N_20680);
xor U24315 (N_24315,N_18997,N_18778);
nor U24316 (N_24316,N_19711,N_20939);
nand U24317 (N_24317,N_19080,N_21640);
nand U24318 (N_24318,N_21045,N_19833);
nor U24319 (N_24319,N_21280,N_21187);
and U24320 (N_24320,N_19226,N_19305);
and U24321 (N_24321,N_20629,N_19347);
and U24322 (N_24322,N_21749,N_19197);
nor U24323 (N_24323,N_20529,N_20683);
xor U24324 (N_24324,N_20477,N_19169);
nand U24325 (N_24325,N_21022,N_18888);
and U24326 (N_24326,N_20019,N_19931);
or U24327 (N_24327,N_21266,N_21386);
nor U24328 (N_24328,N_21147,N_19346);
or U24329 (N_24329,N_19820,N_19770);
xnor U24330 (N_24330,N_21603,N_18936);
nor U24331 (N_24331,N_21614,N_21105);
and U24332 (N_24332,N_19048,N_18939);
nor U24333 (N_24333,N_19754,N_20831);
xor U24334 (N_24334,N_18988,N_20097);
nand U24335 (N_24335,N_21337,N_20255);
and U24336 (N_24336,N_19178,N_21401);
nand U24337 (N_24337,N_18831,N_20316);
nand U24338 (N_24338,N_21127,N_19163);
nor U24339 (N_24339,N_19634,N_20241);
nor U24340 (N_24340,N_19453,N_20017);
xnor U24341 (N_24341,N_21094,N_19186);
nand U24342 (N_24342,N_19498,N_20520);
and U24343 (N_24343,N_21316,N_19884);
and U24344 (N_24344,N_19515,N_21856);
and U24345 (N_24345,N_18995,N_19780);
xnor U24346 (N_24346,N_20114,N_19855);
nand U24347 (N_24347,N_18848,N_19184);
xor U24348 (N_24348,N_19502,N_19896);
nor U24349 (N_24349,N_20438,N_20197);
nand U24350 (N_24350,N_19808,N_20466);
nor U24351 (N_24351,N_19444,N_18963);
or U24352 (N_24352,N_21542,N_19536);
nor U24353 (N_24353,N_19095,N_19564);
nor U24354 (N_24354,N_21130,N_20579);
nand U24355 (N_24355,N_20786,N_20211);
or U24356 (N_24356,N_19176,N_21448);
nor U24357 (N_24357,N_19383,N_20412);
and U24358 (N_24358,N_20110,N_19053);
or U24359 (N_24359,N_20933,N_21455);
nand U24360 (N_24360,N_19635,N_18885);
nand U24361 (N_24361,N_19643,N_19113);
nor U24362 (N_24362,N_21509,N_19834);
nor U24363 (N_24363,N_20626,N_21328);
nor U24364 (N_24364,N_19124,N_19787);
nand U24365 (N_24365,N_19254,N_20696);
xor U24366 (N_24366,N_19581,N_21563);
nor U24367 (N_24367,N_20105,N_20490);
and U24368 (N_24368,N_18921,N_20836);
nor U24369 (N_24369,N_20557,N_21757);
and U24370 (N_24370,N_19850,N_20985);
and U24371 (N_24371,N_20475,N_20623);
and U24372 (N_24372,N_21337,N_21500);
nand U24373 (N_24373,N_20028,N_20668);
or U24374 (N_24374,N_19734,N_19308);
nand U24375 (N_24375,N_20810,N_20925);
nand U24376 (N_24376,N_19680,N_20728);
or U24377 (N_24377,N_20559,N_19608);
nor U24378 (N_24378,N_19129,N_19907);
xor U24379 (N_24379,N_19578,N_20389);
xnor U24380 (N_24380,N_19951,N_19706);
and U24381 (N_24381,N_20990,N_20723);
nand U24382 (N_24382,N_20694,N_21613);
and U24383 (N_24383,N_20789,N_21531);
and U24384 (N_24384,N_20218,N_19346);
nand U24385 (N_24385,N_19490,N_20455);
nor U24386 (N_24386,N_20310,N_20649);
nor U24387 (N_24387,N_21627,N_21352);
nor U24388 (N_24388,N_19519,N_19776);
xnor U24389 (N_24389,N_20906,N_18795);
nand U24390 (N_24390,N_21359,N_20886);
or U24391 (N_24391,N_20367,N_19855);
xor U24392 (N_24392,N_19416,N_19031);
or U24393 (N_24393,N_20414,N_20608);
nand U24394 (N_24394,N_20835,N_20125);
nor U24395 (N_24395,N_20494,N_20111);
nand U24396 (N_24396,N_19779,N_18823);
nand U24397 (N_24397,N_19981,N_21574);
nor U24398 (N_24398,N_19740,N_20299);
and U24399 (N_24399,N_20292,N_21283);
or U24400 (N_24400,N_20829,N_21156);
nor U24401 (N_24401,N_19721,N_20700);
and U24402 (N_24402,N_20503,N_20655);
or U24403 (N_24403,N_21745,N_19541);
and U24404 (N_24404,N_21396,N_20378);
or U24405 (N_24405,N_21350,N_21637);
nand U24406 (N_24406,N_19967,N_20379);
and U24407 (N_24407,N_20936,N_19238);
and U24408 (N_24408,N_19377,N_20264);
nor U24409 (N_24409,N_21211,N_20598);
and U24410 (N_24410,N_21306,N_20305);
nor U24411 (N_24411,N_19170,N_18751);
and U24412 (N_24412,N_19731,N_21728);
nor U24413 (N_24413,N_21599,N_21291);
xnor U24414 (N_24414,N_20615,N_21778);
and U24415 (N_24415,N_19134,N_20611);
nor U24416 (N_24416,N_21215,N_20441);
or U24417 (N_24417,N_20298,N_21604);
nor U24418 (N_24418,N_21496,N_21358);
nor U24419 (N_24419,N_20231,N_19539);
nor U24420 (N_24420,N_19078,N_20381);
and U24421 (N_24421,N_19143,N_20864);
and U24422 (N_24422,N_21799,N_21472);
nor U24423 (N_24423,N_19643,N_21080);
nor U24424 (N_24424,N_19122,N_20493);
nor U24425 (N_24425,N_19786,N_20369);
nand U24426 (N_24426,N_20924,N_20100);
xor U24427 (N_24427,N_18761,N_19287);
nor U24428 (N_24428,N_20533,N_19357);
nor U24429 (N_24429,N_18996,N_21800);
and U24430 (N_24430,N_20716,N_19306);
nand U24431 (N_24431,N_21158,N_19162);
nand U24432 (N_24432,N_19215,N_19083);
nand U24433 (N_24433,N_18774,N_20760);
or U24434 (N_24434,N_21554,N_18979);
and U24435 (N_24435,N_19160,N_19987);
nor U24436 (N_24436,N_20704,N_21043);
and U24437 (N_24437,N_18897,N_18904);
nor U24438 (N_24438,N_21867,N_18786);
nand U24439 (N_24439,N_19645,N_19390);
nand U24440 (N_24440,N_21638,N_20169);
and U24441 (N_24441,N_21090,N_19433);
and U24442 (N_24442,N_21705,N_19458);
nand U24443 (N_24443,N_20320,N_21704);
or U24444 (N_24444,N_20583,N_20856);
or U24445 (N_24445,N_19001,N_19556);
xnor U24446 (N_24446,N_20473,N_19692);
nand U24447 (N_24447,N_20648,N_21226);
nor U24448 (N_24448,N_18831,N_20107);
and U24449 (N_24449,N_19420,N_21831);
or U24450 (N_24450,N_21707,N_19291);
xnor U24451 (N_24451,N_21152,N_20072);
nand U24452 (N_24452,N_20287,N_18759);
or U24453 (N_24453,N_19254,N_20501);
or U24454 (N_24454,N_19605,N_20204);
and U24455 (N_24455,N_21402,N_20633);
xor U24456 (N_24456,N_19224,N_20352);
nor U24457 (N_24457,N_20663,N_20237);
nor U24458 (N_24458,N_19605,N_18975);
nand U24459 (N_24459,N_21512,N_19030);
and U24460 (N_24460,N_21357,N_19347);
nand U24461 (N_24461,N_20530,N_21008);
and U24462 (N_24462,N_20309,N_20033);
or U24463 (N_24463,N_20481,N_20733);
and U24464 (N_24464,N_21871,N_20227);
nand U24465 (N_24465,N_21317,N_18777);
and U24466 (N_24466,N_20041,N_21058);
nor U24467 (N_24467,N_18976,N_20628);
nand U24468 (N_24468,N_18985,N_20895);
xnor U24469 (N_24469,N_20337,N_18907);
and U24470 (N_24470,N_21507,N_19141);
or U24471 (N_24471,N_19351,N_19739);
and U24472 (N_24472,N_20417,N_18844);
xor U24473 (N_24473,N_21617,N_18975);
nor U24474 (N_24474,N_19041,N_21258);
xnor U24475 (N_24475,N_20490,N_21416);
nor U24476 (N_24476,N_21090,N_19715);
nand U24477 (N_24477,N_18964,N_19886);
or U24478 (N_24478,N_19142,N_19318);
nor U24479 (N_24479,N_20340,N_21425);
or U24480 (N_24480,N_19311,N_19691);
nor U24481 (N_24481,N_18897,N_19769);
xnor U24482 (N_24482,N_20757,N_20006);
and U24483 (N_24483,N_19292,N_19390);
or U24484 (N_24484,N_19466,N_20092);
and U24485 (N_24485,N_18945,N_20675);
and U24486 (N_24486,N_20742,N_19218);
nand U24487 (N_24487,N_19878,N_21261);
or U24488 (N_24488,N_20372,N_21305);
nand U24489 (N_24489,N_20973,N_21267);
nor U24490 (N_24490,N_19242,N_21331);
or U24491 (N_24491,N_19737,N_21797);
and U24492 (N_24492,N_21403,N_21343);
nand U24493 (N_24493,N_19195,N_21529);
nand U24494 (N_24494,N_21237,N_19676);
and U24495 (N_24495,N_21147,N_21655);
xnor U24496 (N_24496,N_19971,N_20737);
nor U24497 (N_24497,N_19314,N_19628);
or U24498 (N_24498,N_19704,N_21509);
or U24499 (N_24499,N_20097,N_19888);
and U24500 (N_24500,N_20027,N_19760);
nor U24501 (N_24501,N_19788,N_19913);
and U24502 (N_24502,N_21818,N_19376);
and U24503 (N_24503,N_19562,N_18791);
and U24504 (N_24504,N_19447,N_21345);
nand U24505 (N_24505,N_20076,N_18811);
xor U24506 (N_24506,N_21620,N_19276);
nor U24507 (N_24507,N_19566,N_19599);
and U24508 (N_24508,N_21474,N_20722);
and U24509 (N_24509,N_19427,N_21123);
or U24510 (N_24510,N_19712,N_20674);
nand U24511 (N_24511,N_20076,N_19156);
or U24512 (N_24512,N_18813,N_21017);
and U24513 (N_24513,N_20603,N_20970);
nor U24514 (N_24514,N_20600,N_18866);
nor U24515 (N_24515,N_19980,N_20394);
or U24516 (N_24516,N_20060,N_21814);
nand U24517 (N_24517,N_19926,N_21808);
xor U24518 (N_24518,N_18800,N_19638);
and U24519 (N_24519,N_21041,N_19868);
nand U24520 (N_24520,N_21696,N_19795);
nand U24521 (N_24521,N_18772,N_20241);
xnor U24522 (N_24522,N_20753,N_20119);
xor U24523 (N_24523,N_20823,N_20972);
or U24524 (N_24524,N_19730,N_19678);
nor U24525 (N_24525,N_21047,N_20625);
nor U24526 (N_24526,N_20870,N_19505);
nor U24527 (N_24527,N_21043,N_20062);
or U24528 (N_24528,N_20317,N_21285);
nand U24529 (N_24529,N_18888,N_21338);
nand U24530 (N_24530,N_21113,N_19188);
nand U24531 (N_24531,N_20817,N_19579);
nand U24532 (N_24532,N_20361,N_21197);
nand U24533 (N_24533,N_18987,N_21502);
or U24534 (N_24534,N_20817,N_19469);
or U24535 (N_24535,N_19747,N_21609);
and U24536 (N_24536,N_20593,N_19286);
nand U24537 (N_24537,N_20001,N_20671);
nor U24538 (N_24538,N_21592,N_19231);
nand U24539 (N_24539,N_18854,N_19409);
xnor U24540 (N_24540,N_18766,N_21442);
xnor U24541 (N_24541,N_21763,N_21644);
nand U24542 (N_24542,N_21305,N_19614);
nand U24543 (N_24543,N_19645,N_19159);
nand U24544 (N_24544,N_21129,N_20528);
and U24545 (N_24545,N_21030,N_21787);
xor U24546 (N_24546,N_20065,N_18962);
or U24547 (N_24547,N_21002,N_19569);
xnor U24548 (N_24548,N_19793,N_20441);
xnor U24549 (N_24549,N_19434,N_20059);
nor U24550 (N_24550,N_21172,N_19278);
or U24551 (N_24551,N_20897,N_20531);
nand U24552 (N_24552,N_20330,N_20089);
nor U24553 (N_24553,N_19155,N_21860);
and U24554 (N_24554,N_19284,N_18943);
nand U24555 (N_24555,N_18995,N_19025);
and U24556 (N_24556,N_19984,N_19970);
nand U24557 (N_24557,N_21128,N_19491);
nand U24558 (N_24558,N_21783,N_19739);
nand U24559 (N_24559,N_19022,N_20089);
nor U24560 (N_24560,N_20682,N_21192);
nor U24561 (N_24561,N_21334,N_19250);
xnor U24562 (N_24562,N_18808,N_20888);
and U24563 (N_24563,N_21296,N_20820);
nor U24564 (N_24564,N_21314,N_21551);
and U24565 (N_24565,N_20720,N_21533);
nand U24566 (N_24566,N_19289,N_20687);
nand U24567 (N_24567,N_19189,N_21419);
and U24568 (N_24568,N_21852,N_21479);
and U24569 (N_24569,N_19044,N_20029);
xnor U24570 (N_24570,N_19797,N_20741);
nand U24571 (N_24571,N_21661,N_20192);
or U24572 (N_24572,N_20839,N_20603);
nor U24573 (N_24573,N_20224,N_19706);
or U24574 (N_24574,N_21318,N_21606);
or U24575 (N_24575,N_19171,N_19823);
nand U24576 (N_24576,N_20435,N_20965);
nand U24577 (N_24577,N_21739,N_19310);
or U24578 (N_24578,N_21000,N_20558);
nand U24579 (N_24579,N_19849,N_21588);
and U24580 (N_24580,N_20421,N_20087);
and U24581 (N_24581,N_21149,N_20332);
nor U24582 (N_24582,N_21571,N_21794);
nor U24583 (N_24583,N_20912,N_19014);
or U24584 (N_24584,N_20679,N_20569);
nor U24585 (N_24585,N_19323,N_19049);
or U24586 (N_24586,N_19348,N_20710);
nor U24587 (N_24587,N_21813,N_21160);
nor U24588 (N_24588,N_21505,N_21654);
nand U24589 (N_24589,N_20419,N_20631);
and U24590 (N_24590,N_19343,N_19057);
xor U24591 (N_24591,N_19211,N_19806);
nand U24592 (N_24592,N_19108,N_19316);
nand U24593 (N_24593,N_19927,N_21162);
nor U24594 (N_24594,N_18961,N_20199);
nor U24595 (N_24595,N_21454,N_19538);
xor U24596 (N_24596,N_21785,N_21811);
or U24597 (N_24597,N_19011,N_21274);
xnor U24598 (N_24598,N_19837,N_19170);
and U24599 (N_24599,N_19459,N_19000);
nand U24600 (N_24600,N_21128,N_18916);
or U24601 (N_24601,N_20747,N_21117);
nor U24602 (N_24602,N_21853,N_20322);
and U24603 (N_24603,N_19696,N_21609);
and U24604 (N_24604,N_19902,N_20523);
and U24605 (N_24605,N_19662,N_20565);
and U24606 (N_24606,N_21824,N_20346);
nand U24607 (N_24607,N_21086,N_19890);
and U24608 (N_24608,N_21487,N_20461);
and U24609 (N_24609,N_21392,N_21160);
and U24610 (N_24610,N_21752,N_19584);
nor U24611 (N_24611,N_20676,N_18870);
nand U24612 (N_24612,N_19814,N_19557);
and U24613 (N_24613,N_19038,N_19908);
nor U24614 (N_24614,N_19500,N_21265);
xnor U24615 (N_24615,N_20840,N_21593);
and U24616 (N_24616,N_18889,N_21097);
nand U24617 (N_24617,N_19140,N_21668);
and U24618 (N_24618,N_19612,N_19061);
or U24619 (N_24619,N_19603,N_21341);
xnor U24620 (N_24620,N_20379,N_18752);
nand U24621 (N_24621,N_19719,N_20387);
xnor U24622 (N_24622,N_21185,N_21389);
or U24623 (N_24623,N_20231,N_20932);
nor U24624 (N_24624,N_21147,N_18955);
xnor U24625 (N_24625,N_20673,N_20392);
or U24626 (N_24626,N_19366,N_21834);
nor U24627 (N_24627,N_21536,N_20289);
nand U24628 (N_24628,N_20315,N_19177);
nor U24629 (N_24629,N_21764,N_21202);
or U24630 (N_24630,N_19102,N_20018);
and U24631 (N_24631,N_21562,N_20928);
nor U24632 (N_24632,N_20812,N_21355);
or U24633 (N_24633,N_19119,N_21163);
nand U24634 (N_24634,N_21804,N_21381);
nand U24635 (N_24635,N_19095,N_20535);
or U24636 (N_24636,N_19043,N_20888);
and U24637 (N_24637,N_20269,N_20024);
and U24638 (N_24638,N_21289,N_20214);
nor U24639 (N_24639,N_20520,N_20009);
or U24640 (N_24640,N_20824,N_20850);
nor U24641 (N_24641,N_20911,N_21235);
xor U24642 (N_24642,N_19178,N_21120);
or U24643 (N_24643,N_21439,N_20202);
nand U24644 (N_24644,N_20425,N_18824);
nand U24645 (N_24645,N_19801,N_21790);
or U24646 (N_24646,N_19178,N_21508);
nor U24647 (N_24647,N_21805,N_19341);
nand U24648 (N_24648,N_21160,N_18931);
or U24649 (N_24649,N_20981,N_20425);
and U24650 (N_24650,N_19376,N_20302);
or U24651 (N_24651,N_21144,N_21376);
or U24652 (N_24652,N_21514,N_21261);
or U24653 (N_24653,N_20966,N_21409);
nor U24654 (N_24654,N_19386,N_21452);
nor U24655 (N_24655,N_18763,N_19268);
or U24656 (N_24656,N_21550,N_20623);
or U24657 (N_24657,N_21342,N_21371);
and U24658 (N_24658,N_18841,N_19778);
nand U24659 (N_24659,N_21790,N_19472);
nor U24660 (N_24660,N_20723,N_19971);
nor U24661 (N_24661,N_20915,N_20773);
nor U24662 (N_24662,N_19347,N_19064);
xor U24663 (N_24663,N_21381,N_19718);
nand U24664 (N_24664,N_20843,N_20521);
nor U24665 (N_24665,N_21530,N_19425);
or U24666 (N_24666,N_20136,N_20657);
or U24667 (N_24667,N_19362,N_21573);
and U24668 (N_24668,N_21410,N_21671);
or U24669 (N_24669,N_21091,N_18765);
or U24670 (N_24670,N_20267,N_21533);
xnor U24671 (N_24671,N_20541,N_20801);
nor U24672 (N_24672,N_18951,N_21743);
and U24673 (N_24673,N_21631,N_20262);
nand U24674 (N_24674,N_21455,N_20880);
nor U24675 (N_24675,N_20037,N_21159);
nand U24676 (N_24676,N_21854,N_20954);
nand U24677 (N_24677,N_19409,N_18971);
nor U24678 (N_24678,N_21244,N_19713);
and U24679 (N_24679,N_19054,N_19067);
nor U24680 (N_24680,N_20889,N_20583);
nand U24681 (N_24681,N_19552,N_19412);
xnor U24682 (N_24682,N_19265,N_20483);
or U24683 (N_24683,N_21020,N_21631);
and U24684 (N_24684,N_21650,N_19396);
or U24685 (N_24685,N_21848,N_20669);
nand U24686 (N_24686,N_19843,N_18818);
or U24687 (N_24687,N_21211,N_21195);
and U24688 (N_24688,N_20758,N_20164);
nor U24689 (N_24689,N_20418,N_21436);
and U24690 (N_24690,N_20000,N_21536);
nor U24691 (N_24691,N_20250,N_20470);
nand U24692 (N_24692,N_21071,N_20164);
nand U24693 (N_24693,N_21079,N_21305);
nand U24694 (N_24694,N_20809,N_21091);
or U24695 (N_24695,N_20397,N_21514);
and U24696 (N_24696,N_21613,N_21140);
nand U24697 (N_24697,N_19132,N_19697);
nor U24698 (N_24698,N_21254,N_21381);
xor U24699 (N_24699,N_21393,N_18809);
nand U24700 (N_24700,N_21298,N_19182);
nor U24701 (N_24701,N_20942,N_19876);
and U24702 (N_24702,N_19030,N_20244);
nand U24703 (N_24703,N_19715,N_19790);
and U24704 (N_24704,N_20208,N_21603);
and U24705 (N_24705,N_19703,N_21354);
nor U24706 (N_24706,N_21621,N_21198);
nor U24707 (N_24707,N_20779,N_19924);
nor U24708 (N_24708,N_21322,N_20634);
nand U24709 (N_24709,N_19462,N_21678);
nor U24710 (N_24710,N_19059,N_21391);
and U24711 (N_24711,N_20987,N_18975);
or U24712 (N_24712,N_18752,N_21764);
nand U24713 (N_24713,N_21167,N_20008);
and U24714 (N_24714,N_21755,N_19150);
nor U24715 (N_24715,N_18860,N_19320);
and U24716 (N_24716,N_21741,N_18877);
nor U24717 (N_24717,N_21349,N_20716);
nand U24718 (N_24718,N_18861,N_19923);
nand U24719 (N_24719,N_18763,N_21410);
nand U24720 (N_24720,N_21450,N_21060);
nand U24721 (N_24721,N_21493,N_20812);
or U24722 (N_24722,N_19850,N_18808);
nor U24723 (N_24723,N_20343,N_19494);
or U24724 (N_24724,N_19760,N_21638);
xnor U24725 (N_24725,N_20181,N_21203);
or U24726 (N_24726,N_20033,N_19351);
and U24727 (N_24727,N_20208,N_19719);
nor U24728 (N_24728,N_20529,N_19897);
xnor U24729 (N_24729,N_21642,N_20075);
and U24730 (N_24730,N_21801,N_19243);
nor U24731 (N_24731,N_20656,N_21739);
nor U24732 (N_24732,N_21122,N_20224);
and U24733 (N_24733,N_20496,N_21201);
or U24734 (N_24734,N_19153,N_19638);
nand U24735 (N_24735,N_20464,N_18860);
nor U24736 (N_24736,N_18959,N_20633);
nand U24737 (N_24737,N_20994,N_19093);
and U24738 (N_24738,N_19568,N_21832);
and U24739 (N_24739,N_19351,N_19034);
nand U24740 (N_24740,N_19200,N_19849);
or U24741 (N_24741,N_19311,N_20045);
and U24742 (N_24742,N_20439,N_19776);
xnor U24743 (N_24743,N_19522,N_19327);
nand U24744 (N_24744,N_19596,N_19964);
nand U24745 (N_24745,N_21698,N_20694);
nand U24746 (N_24746,N_21387,N_20240);
and U24747 (N_24747,N_21547,N_19599);
and U24748 (N_24748,N_21187,N_21005);
nor U24749 (N_24749,N_21461,N_19144);
nor U24750 (N_24750,N_20641,N_18830);
xor U24751 (N_24751,N_19142,N_19680);
nor U24752 (N_24752,N_18891,N_21044);
nand U24753 (N_24753,N_20313,N_20828);
nand U24754 (N_24754,N_21715,N_20488);
or U24755 (N_24755,N_18765,N_21754);
and U24756 (N_24756,N_20451,N_21178);
xor U24757 (N_24757,N_19296,N_19760);
nand U24758 (N_24758,N_18824,N_20693);
xor U24759 (N_24759,N_20555,N_20989);
nor U24760 (N_24760,N_20958,N_21002);
and U24761 (N_24761,N_19455,N_19923);
nor U24762 (N_24762,N_20407,N_21718);
and U24763 (N_24763,N_20508,N_21208);
or U24764 (N_24764,N_19418,N_21013);
or U24765 (N_24765,N_19443,N_18758);
and U24766 (N_24766,N_21597,N_19194);
and U24767 (N_24767,N_20629,N_21719);
nor U24768 (N_24768,N_21542,N_20030);
and U24769 (N_24769,N_19153,N_20947);
and U24770 (N_24770,N_19845,N_19821);
and U24771 (N_24771,N_20582,N_19731);
xor U24772 (N_24772,N_19501,N_20813);
xnor U24773 (N_24773,N_21327,N_20727);
and U24774 (N_24774,N_20465,N_21315);
xor U24775 (N_24775,N_19251,N_19966);
nand U24776 (N_24776,N_20355,N_20645);
and U24777 (N_24777,N_21177,N_20664);
or U24778 (N_24778,N_20931,N_21536);
nor U24779 (N_24779,N_18855,N_19845);
nor U24780 (N_24780,N_20263,N_19303);
and U24781 (N_24781,N_19392,N_20972);
or U24782 (N_24782,N_20768,N_21596);
or U24783 (N_24783,N_20575,N_21647);
xnor U24784 (N_24784,N_19855,N_20608);
nor U24785 (N_24785,N_21429,N_21109);
xor U24786 (N_24786,N_19797,N_19410);
or U24787 (N_24787,N_18769,N_20642);
and U24788 (N_24788,N_19411,N_19266);
or U24789 (N_24789,N_21296,N_19129);
and U24790 (N_24790,N_18876,N_21002);
or U24791 (N_24791,N_19749,N_21790);
nor U24792 (N_24792,N_20091,N_20527);
nor U24793 (N_24793,N_19946,N_18867);
xnor U24794 (N_24794,N_20571,N_19299);
nand U24795 (N_24795,N_19764,N_20756);
or U24796 (N_24796,N_21221,N_20939);
or U24797 (N_24797,N_20121,N_20357);
nor U24798 (N_24798,N_21056,N_21004);
nand U24799 (N_24799,N_20566,N_20189);
nand U24800 (N_24800,N_20120,N_21407);
nor U24801 (N_24801,N_18988,N_21575);
or U24802 (N_24802,N_19966,N_20645);
nor U24803 (N_24803,N_19478,N_20962);
nor U24804 (N_24804,N_20287,N_21862);
xor U24805 (N_24805,N_20957,N_19097);
or U24806 (N_24806,N_19656,N_19854);
xnor U24807 (N_24807,N_18972,N_19024);
xnor U24808 (N_24808,N_18844,N_19238);
nand U24809 (N_24809,N_20513,N_20787);
and U24810 (N_24810,N_20601,N_19382);
or U24811 (N_24811,N_20220,N_21290);
nand U24812 (N_24812,N_19253,N_19318);
nand U24813 (N_24813,N_20654,N_18969);
nand U24814 (N_24814,N_20979,N_19613);
or U24815 (N_24815,N_19653,N_20792);
xor U24816 (N_24816,N_19235,N_19160);
nand U24817 (N_24817,N_19476,N_20156);
nand U24818 (N_24818,N_21616,N_21618);
or U24819 (N_24819,N_20640,N_19507);
nand U24820 (N_24820,N_19494,N_19231);
nand U24821 (N_24821,N_19453,N_19224);
and U24822 (N_24822,N_19108,N_21866);
xnor U24823 (N_24823,N_21540,N_20900);
and U24824 (N_24824,N_21552,N_21174);
nand U24825 (N_24825,N_18998,N_19505);
and U24826 (N_24826,N_20605,N_19863);
nand U24827 (N_24827,N_18983,N_20557);
nand U24828 (N_24828,N_18894,N_19460);
nor U24829 (N_24829,N_19508,N_20994);
and U24830 (N_24830,N_20180,N_19853);
and U24831 (N_24831,N_19821,N_18892);
xor U24832 (N_24832,N_19590,N_20962);
nand U24833 (N_24833,N_19367,N_21561);
nand U24834 (N_24834,N_21569,N_21552);
nand U24835 (N_24835,N_21231,N_20662);
xor U24836 (N_24836,N_20524,N_21042);
nand U24837 (N_24837,N_20954,N_21153);
and U24838 (N_24838,N_21695,N_20116);
nor U24839 (N_24839,N_19351,N_21628);
xor U24840 (N_24840,N_20998,N_20580);
and U24841 (N_24841,N_21206,N_18807);
or U24842 (N_24842,N_19928,N_19473);
nand U24843 (N_24843,N_21039,N_19357);
nor U24844 (N_24844,N_20061,N_21223);
and U24845 (N_24845,N_21321,N_19650);
and U24846 (N_24846,N_20654,N_19431);
or U24847 (N_24847,N_21670,N_21277);
nand U24848 (N_24848,N_19688,N_21578);
nor U24849 (N_24849,N_21162,N_21168);
nor U24850 (N_24850,N_21145,N_21300);
or U24851 (N_24851,N_19454,N_21051);
nor U24852 (N_24852,N_19422,N_20917);
or U24853 (N_24853,N_21259,N_20466);
xnor U24854 (N_24854,N_19381,N_20442);
nand U24855 (N_24855,N_21421,N_20404);
nand U24856 (N_24856,N_21293,N_20708);
or U24857 (N_24857,N_19447,N_20211);
or U24858 (N_24858,N_21294,N_19257);
and U24859 (N_24859,N_21565,N_20162);
or U24860 (N_24860,N_20795,N_21274);
and U24861 (N_24861,N_20984,N_19288);
or U24862 (N_24862,N_21054,N_21283);
nand U24863 (N_24863,N_20594,N_21383);
or U24864 (N_24864,N_19410,N_18906);
nor U24865 (N_24865,N_21533,N_19104);
and U24866 (N_24866,N_19752,N_20249);
nand U24867 (N_24867,N_19265,N_21203);
or U24868 (N_24868,N_19847,N_21336);
nor U24869 (N_24869,N_20981,N_19882);
nor U24870 (N_24870,N_19737,N_20559);
nor U24871 (N_24871,N_21388,N_21536);
xnor U24872 (N_24872,N_19793,N_21252);
and U24873 (N_24873,N_21073,N_19752);
nand U24874 (N_24874,N_19290,N_19226);
nand U24875 (N_24875,N_21002,N_19206);
or U24876 (N_24876,N_19794,N_19314);
nor U24877 (N_24877,N_20845,N_19089);
or U24878 (N_24878,N_20602,N_20494);
xnor U24879 (N_24879,N_18865,N_19043);
nand U24880 (N_24880,N_19824,N_20600);
nand U24881 (N_24881,N_19515,N_21568);
nor U24882 (N_24882,N_21609,N_21572);
or U24883 (N_24883,N_19020,N_20717);
nor U24884 (N_24884,N_20452,N_19137);
and U24885 (N_24885,N_20850,N_20699);
or U24886 (N_24886,N_21063,N_20349);
xor U24887 (N_24887,N_20410,N_19128);
xnor U24888 (N_24888,N_21373,N_19516);
nor U24889 (N_24889,N_20067,N_21751);
nor U24890 (N_24890,N_20908,N_19735);
and U24891 (N_24891,N_19725,N_21517);
nand U24892 (N_24892,N_19787,N_21781);
nand U24893 (N_24893,N_20122,N_20533);
nand U24894 (N_24894,N_18836,N_21618);
and U24895 (N_24895,N_19088,N_20939);
and U24896 (N_24896,N_20559,N_20777);
xnor U24897 (N_24897,N_21829,N_19336);
or U24898 (N_24898,N_20876,N_19637);
and U24899 (N_24899,N_19470,N_19523);
nand U24900 (N_24900,N_19591,N_21400);
and U24901 (N_24901,N_19030,N_19930);
nand U24902 (N_24902,N_20397,N_20122);
nand U24903 (N_24903,N_21191,N_20177);
xnor U24904 (N_24904,N_19062,N_19894);
nor U24905 (N_24905,N_20528,N_20274);
nor U24906 (N_24906,N_20531,N_20951);
nor U24907 (N_24907,N_19586,N_19280);
nor U24908 (N_24908,N_19736,N_18883);
nor U24909 (N_24909,N_21469,N_19435);
and U24910 (N_24910,N_19749,N_20434);
nand U24911 (N_24911,N_19209,N_19032);
and U24912 (N_24912,N_19969,N_19727);
nand U24913 (N_24913,N_20097,N_20659);
nor U24914 (N_24914,N_20312,N_21476);
and U24915 (N_24915,N_20111,N_20400);
nand U24916 (N_24916,N_21523,N_19555);
and U24917 (N_24917,N_20387,N_18943);
nor U24918 (N_24918,N_19606,N_20169);
and U24919 (N_24919,N_19041,N_19009);
or U24920 (N_24920,N_19632,N_21481);
and U24921 (N_24921,N_18898,N_21674);
nand U24922 (N_24922,N_18825,N_20311);
nand U24923 (N_24923,N_20963,N_20322);
and U24924 (N_24924,N_20686,N_20046);
and U24925 (N_24925,N_20997,N_21534);
or U24926 (N_24926,N_20551,N_20464);
nand U24927 (N_24927,N_20071,N_19212);
and U24928 (N_24928,N_20907,N_19526);
and U24929 (N_24929,N_19630,N_21501);
or U24930 (N_24930,N_18948,N_21604);
and U24931 (N_24931,N_21415,N_19041);
nor U24932 (N_24932,N_20575,N_19002);
or U24933 (N_24933,N_21348,N_21604);
and U24934 (N_24934,N_20667,N_21131);
nand U24935 (N_24935,N_20645,N_19103);
xnor U24936 (N_24936,N_21385,N_19853);
nor U24937 (N_24937,N_18831,N_20359);
and U24938 (N_24938,N_21751,N_20456);
and U24939 (N_24939,N_20135,N_20938);
nor U24940 (N_24940,N_19912,N_21511);
nor U24941 (N_24941,N_19986,N_19585);
and U24942 (N_24942,N_21557,N_21809);
nand U24943 (N_24943,N_18893,N_19178);
and U24944 (N_24944,N_19073,N_19793);
or U24945 (N_24945,N_21345,N_19624);
or U24946 (N_24946,N_20691,N_19758);
and U24947 (N_24947,N_19682,N_19157);
nand U24948 (N_24948,N_20255,N_19842);
nor U24949 (N_24949,N_20862,N_19696);
nor U24950 (N_24950,N_21181,N_21037);
or U24951 (N_24951,N_21561,N_20571);
and U24952 (N_24952,N_21104,N_19091);
and U24953 (N_24953,N_21414,N_21236);
nand U24954 (N_24954,N_19547,N_19587);
and U24955 (N_24955,N_21023,N_19778);
and U24956 (N_24956,N_18757,N_21483);
xnor U24957 (N_24957,N_20913,N_21748);
and U24958 (N_24958,N_19859,N_20147);
or U24959 (N_24959,N_19338,N_18864);
nor U24960 (N_24960,N_19449,N_19605);
nor U24961 (N_24961,N_20115,N_19830);
or U24962 (N_24962,N_19373,N_19064);
and U24963 (N_24963,N_21677,N_20193);
nor U24964 (N_24964,N_21701,N_20999);
or U24965 (N_24965,N_20083,N_20746);
or U24966 (N_24966,N_21814,N_19840);
nand U24967 (N_24967,N_19413,N_18927);
nand U24968 (N_24968,N_18757,N_19364);
nor U24969 (N_24969,N_21789,N_19195);
nor U24970 (N_24970,N_20287,N_20541);
nor U24971 (N_24971,N_21791,N_19179);
nor U24972 (N_24972,N_20353,N_19658);
or U24973 (N_24973,N_18934,N_19445);
nor U24974 (N_24974,N_20458,N_20649);
nor U24975 (N_24975,N_20204,N_20702);
nand U24976 (N_24976,N_19529,N_19494);
or U24977 (N_24977,N_20738,N_20579);
nor U24978 (N_24978,N_19081,N_19963);
nand U24979 (N_24979,N_20109,N_20477);
nand U24980 (N_24980,N_20903,N_19740);
nand U24981 (N_24981,N_20628,N_21073);
nand U24982 (N_24982,N_19243,N_19132);
nand U24983 (N_24983,N_20101,N_19422);
nand U24984 (N_24984,N_19437,N_18923);
and U24985 (N_24985,N_20731,N_19246);
and U24986 (N_24986,N_20729,N_20111);
xor U24987 (N_24987,N_21582,N_21324);
or U24988 (N_24988,N_19972,N_21304);
or U24989 (N_24989,N_20988,N_19553);
or U24990 (N_24990,N_19486,N_20581);
nand U24991 (N_24991,N_21131,N_19556);
nor U24992 (N_24992,N_20153,N_21710);
or U24993 (N_24993,N_18806,N_19214);
or U24994 (N_24994,N_19750,N_19796);
nor U24995 (N_24995,N_21623,N_19292);
xor U24996 (N_24996,N_20047,N_18763);
or U24997 (N_24997,N_19000,N_21536);
or U24998 (N_24998,N_19493,N_19100);
nand U24999 (N_24999,N_20043,N_21547);
xnor UO_0 (O_0,N_24320,N_23114);
or UO_1 (O_1,N_22327,N_24068);
and UO_2 (O_2,N_23126,N_23997);
nor UO_3 (O_3,N_24926,N_24568);
xnor UO_4 (O_4,N_22686,N_24486);
or UO_5 (O_5,N_24507,N_24716);
and UO_6 (O_6,N_22492,N_23320);
nand UO_7 (O_7,N_24178,N_23674);
xor UO_8 (O_8,N_23771,N_23491);
xnor UO_9 (O_9,N_24375,N_24441);
nand UO_10 (O_10,N_24688,N_24429);
or UO_11 (O_11,N_22651,N_23575);
and UO_12 (O_12,N_24682,N_24808);
nand UO_13 (O_13,N_24487,N_22553);
and UO_14 (O_14,N_23365,N_24756);
nor UO_15 (O_15,N_23151,N_22920);
nand UO_16 (O_16,N_23901,N_23883);
or UO_17 (O_17,N_22352,N_24280);
and UO_18 (O_18,N_23594,N_24657);
nor UO_19 (O_19,N_22406,N_24311);
nand UO_20 (O_20,N_22059,N_24386);
nand UO_21 (O_21,N_22106,N_23058);
and UO_22 (O_22,N_23744,N_23010);
nand UO_23 (O_23,N_22608,N_21940);
xor UO_24 (O_24,N_24780,N_22743);
nor UO_25 (O_25,N_23557,N_22120);
and UO_26 (O_26,N_23445,N_22110);
and UO_27 (O_27,N_22595,N_24952);
and UO_28 (O_28,N_22262,N_23696);
nor UO_29 (O_29,N_23641,N_21989);
nor UO_30 (O_30,N_24293,N_24318);
xor UO_31 (O_31,N_22171,N_23726);
and UO_32 (O_32,N_23900,N_21988);
xor UO_33 (O_33,N_23029,N_22502);
nand UO_34 (O_34,N_24356,N_22934);
and UO_35 (O_35,N_22832,N_24860);
or UO_36 (O_36,N_23977,N_24238);
or UO_37 (O_37,N_24433,N_22444);
nor UO_38 (O_38,N_24382,N_23429);
nand UO_39 (O_39,N_24829,N_24329);
nor UO_40 (O_40,N_22831,N_22551);
and UO_41 (O_41,N_24976,N_22792);
xor UO_42 (O_42,N_24466,N_22081);
nor UO_43 (O_43,N_24727,N_22716);
or UO_44 (O_44,N_24287,N_24800);
or UO_45 (O_45,N_23005,N_24425);
or UO_46 (O_46,N_24518,N_24701);
nor UO_47 (O_47,N_23720,N_22529);
or UO_48 (O_48,N_22732,N_22390);
and UO_49 (O_49,N_22637,N_23070);
or UO_50 (O_50,N_24485,N_24809);
or UO_51 (O_51,N_24685,N_23030);
and UO_52 (O_52,N_24286,N_24640);
nor UO_53 (O_53,N_22225,N_22190);
or UO_54 (O_54,N_23555,N_22523);
xnor UO_55 (O_55,N_23342,N_22034);
nor UO_56 (O_56,N_22538,N_21879);
or UO_57 (O_57,N_23886,N_22535);
nand UO_58 (O_58,N_21890,N_24457);
nor UO_59 (O_59,N_22069,N_22270);
and UO_60 (O_60,N_22905,N_24134);
and UO_61 (O_61,N_24531,N_23716);
nor UO_62 (O_62,N_24530,N_24438);
nand UO_63 (O_63,N_23207,N_21927);
nor UO_64 (O_64,N_21950,N_24924);
nand UO_65 (O_65,N_23566,N_24624);
nor UO_66 (O_66,N_22672,N_22654);
or UO_67 (O_67,N_23194,N_24172);
or UO_68 (O_68,N_23522,N_24129);
nor UO_69 (O_69,N_23602,N_23556);
nor UO_70 (O_70,N_24615,N_22849);
and UO_71 (O_71,N_23586,N_23948);
and UO_72 (O_72,N_24360,N_24533);
or UO_73 (O_73,N_21992,N_24902);
xnor UO_74 (O_74,N_22450,N_23062);
and UO_75 (O_75,N_23650,N_23091);
and UO_76 (O_76,N_24559,N_23806);
nor UO_77 (O_77,N_22917,N_22240);
and UO_78 (O_78,N_24519,N_22884);
nor UO_79 (O_79,N_22058,N_22638);
nand UO_80 (O_80,N_23262,N_24960);
nor UO_81 (O_81,N_23847,N_23971);
and UO_82 (O_82,N_24529,N_22969);
nand UO_83 (O_83,N_24736,N_24005);
and UO_84 (O_84,N_22900,N_23042);
nor UO_85 (O_85,N_21931,N_24231);
nand UO_86 (O_86,N_23895,N_23468);
nand UO_87 (O_87,N_24648,N_23316);
nor UO_88 (O_88,N_22130,N_23982);
nand UO_89 (O_89,N_24414,N_24986);
or UO_90 (O_90,N_22630,N_24089);
nor UO_91 (O_91,N_24334,N_23874);
and UO_92 (O_92,N_24883,N_21974);
and UO_93 (O_93,N_23577,N_23307);
nand UO_94 (O_94,N_21990,N_22203);
nor UO_95 (O_95,N_23408,N_23434);
nor UO_96 (O_96,N_24228,N_23687);
nand UO_97 (O_97,N_23795,N_24097);
nand UO_98 (O_98,N_24171,N_24206);
nand UO_99 (O_99,N_23609,N_24107);
or UO_100 (O_100,N_22016,N_23372);
or UO_101 (O_101,N_22495,N_23222);
or UO_102 (O_102,N_24775,N_22956);
nor UO_103 (O_103,N_22873,N_23564);
nor UO_104 (O_104,N_22250,N_24575);
nand UO_105 (O_105,N_22620,N_23815);
nor UO_106 (O_106,N_24475,N_24418);
and UO_107 (O_107,N_22824,N_23155);
and UO_108 (O_108,N_22966,N_24948);
and UO_109 (O_109,N_21893,N_24950);
or UO_110 (O_110,N_23084,N_23177);
or UO_111 (O_111,N_22937,N_23006);
nor UO_112 (O_112,N_24762,N_23255);
nor UO_113 (O_113,N_23184,N_21942);
xor UO_114 (O_114,N_22558,N_24304);
nand UO_115 (O_115,N_22435,N_24778);
nor UO_116 (O_116,N_24901,N_23119);
nand UO_117 (O_117,N_21972,N_23373);
and UO_118 (O_118,N_23117,N_22978);
nor UO_119 (O_119,N_24539,N_22091);
and UO_120 (O_120,N_22636,N_24261);
nor UO_121 (O_121,N_23394,N_22709);
nand UO_122 (O_122,N_24580,N_24381);
xnor UO_123 (O_123,N_22441,N_23103);
or UO_124 (O_124,N_24627,N_23406);
nor UO_125 (O_125,N_24750,N_23921);
or UO_126 (O_126,N_23607,N_24361);
or UO_127 (O_127,N_23427,N_24050);
and UO_128 (O_128,N_24151,N_24871);
xor UO_129 (O_129,N_24608,N_22283);
and UO_130 (O_130,N_22547,N_22744);
xor UO_131 (O_131,N_22028,N_23656);
nand UO_132 (O_132,N_23987,N_24257);
or UO_133 (O_133,N_24879,N_23509);
or UO_134 (O_134,N_21943,N_23894);
or UO_135 (O_135,N_24018,N_24020);
nand UO_136 (O_136,N_24385,N_24120);
and UO_137 (O_137,N_24613,N_23519);
nor UO_138 (O_138,N_22735,N_21935);
and UO_139 (O_139,N_23423,N_24663);
nor UO_140 (O_140,N_24152,N_22417);
xnor UO_141 (O_141,N_23024,N_24600);
nor UO_142 (O_142,N_22197,N_22606);
and UO_143 (O_143,N_23187,N_22570);
nor UO_144 (O_144,N_22546,N_24073);
nor UO_145 (O_145,N_24093,N_22384);
xor UO_146 (O_146,N_24678,N_22481);
nor UO_147 (O_147,N_23672,N_24269);
nand UO_148 (O_148,N_22919,N_24392);
nand UO_149 (O_149,N_24255,N_23623);
nor UO_150 (O_150,N_24470,N_24511);
nor UO_151 (O_151,N_23147,N_23714);
nor UO_152 (O_152,N_22680,N_22316);
or UO_153 (O_153,N_22658,N_23397);
and UO_154 (O_154,N_24143,N_23466);
and UO_155 (O_155,N_23392,N_24747);
nand UO_156 (O_156,N_24467,N_23165);
or UO_157 (O_157,N_23610,N_22685);
nor UO_158 (O_158,N_24870,N_23381);
or UO_159 (O_159,N_22005,N_24934);
nand UO_160 (O_160,N_22101,N_23475);
and UO_161 (O_161,N_23769,N_22914);
nor UO_162 (O_162,N_22756,N_21999);
nand UO_163 (O_163,N_24612,N_23549);
nand UO_164 (O_164,N_21899,N_22819);
nand UO_165 (O_165,N_22255,N_24781);
nor UO_166 (O_166,N_22191,N_24201);
nor UO_167 (O_167,N_22200,N_23315);
or UO_168 (O_168,N_21977,N_24291);
nand UO_169 (O_169,N_23620,N_22548);
and UO_170 (O_170,N_23888,N_22902);
xor UO_171 (O_171,N_23951,N_22291);
and UO_172 (O_172,N_22017,N_22345);
or UO_173 (O_173,N_22883,N_23374);
and UO_174 (O_174,N_21930,N_21877);
nand UO_175 (O_175,N_23628,N_23118);
and UO_176 (O_176,N_24430,N_24204);
and UO_177 (O_177,N_22749,N_23388);
or UO_178 (O_178,N_22252,N_22333);
nor UO_179 (O_179,N_22602,N_22415);
nor UO_180 (O_180,N_23679,N_23698);
and UO_181 (O_181,N_22152,N_23780);
and UO_182 (O_182,N_23823,N_23668);
and UO_183 (O_183,N_22768,N_22555);
or UO_184 (O_184,N_24935,N_22635);
and UO_185 (O_185,N_24319,N_24294);
nor UO_186 (O_186,N_22413,N_24521);
and UO_187 (O_187,N_22282,N_23966);
nand UO_188 (O_188,N_22108,N_23304);
and UO_189 (O_189,N_23197,N_22587);
and UO_190 (O_190,N_24340,N_23776);
or UO_191 (O_191,N_24570,N_23428);
or UO_192 (O_192,N_24308,N_22426);
nor UO_193 (O_193,N_22031,N_23565);
nor UO_194 (O_194,N_23879,N_22961);
or UO_195 (O_195,N_23133,N_22713);
or UO_196 (O_196,N_22276,N_24621);
or UO_197 (O_197,N_23738,N_24740);
and UO_198 (O_198,N_22738,N_23600);
and UO_199 (O_199,N_24564,N_24514);
nor UO_200 (O_200,N_24633,N_24119);
or UO_201 (O_201,N_23759,N_22012);
nand UO_202 (O_202,N_23527,N_24397);
and UO_203 (O_203,N_23431,N_22051);
and UO_204 (O_204,N_22964,N_22950);
nor UO_205 (O_205,N_21906,N_24919);
or UO_206 (O_206,N_23282,N_22092);
or UO_207 (O_207,N_22463,N_24281);
nand UO_208 (O_208,N_24289,N_22422);
and UO_209 (O_209,N_23673,N_23975);
and UO_210 (O_210,N_22099,N_24165);
nor UO_211 (O_211,N_23905,N_22418);
nor UO_212 (O_212,N_22607,N_23560);
nand UO_213 (O_213,N_22246,N_22509);
or UO_214 (O_214,N_22701,N_22077);
xnor UO_215 (O_215,N_24796,N_23188);
or UO_216 (O_216,N_22731,N_22598);
and UO_217 (O_217,N_23362,N_24015);
nor UO_218 (O_218,N_22863,N_22391);
nand UO_219 (O_219,N_24041,N_24807);
or UO_220 (O_220,N_23956,N_21966);
or UO_221 (O_221,N_24225,N_23449);
and UO_222 (O_222,N_23723,N_24783);
nand UO_223 (O_223,N_22922,N_24732);
nor UO_224 (O_224,N_24148,N_23200);
or UO_225 (O_225,N_22036,N_24984);
or UO_226 (O_226,N_24370,N_22531);
and UO_227 (O_227,N_23477,N_23409);
or UO_228 (O_228,N_23020,N_22464);
and UO_229 (O_229,N_22898,N_23183);
nand UO_230 (O_230,N_24694,N_24272);
nor UO_231 (O_231,N_22584,N_22767);
and UO_232 (O_232,N_22334,N_24478);
nand UO_233 (O_233,N_24704,N_24208);
nor UO_234 (O_234,N_22088,N_24906);
nor UO_235 (O_235,N_23023,N_21944);
or UO_236 (O_236,N_23680,N_22449);
or UO_237 (O_237,N_23358,N_23414);
xnor UO_238 (O_238,N_24819,N_23099);
and UO_239 (O_239,N_22520,N_24757);
nand UO_240 (O_240,N_22820,N_23772);
and UO_241 (O_241,N_21991,N_24468);
nand UO_242 (O_242,N_22998,N_22562);
nand UO_243 (O_243,N_24066,N_24927);
or UO_244 (O_244,N_22440,N_23225);
xor UO_245 (O_245,N_23938,N_21937);
nand UO_246 (O_246,N_23887,N_22826);
or UO_247 (O_247,N_22168,N_21916);
nor UO_248 (O_248,N_24354,N_23713);
and UO_249 (O_249,N_22526,N_22396);
nand UO_250 (O_250,N_24472,N_22879);
and UO_251 (O_251,N_23068,N_22503);
nor UO_252 (O_252,N_24275,N_22321);
xnor UO_253 (O_253,N_22420,N_24210);
nand UO_254 (O_254,N_23047,N_21882);
or UO_255 (O_255,N_24122,N_22882);
or UO_256 (O_256,N_24597,N_22003);
and UO_257 (O_257,N_22625,N_24974);
nor UO_258 (O_258,N_22999,N_24173);
xnor UO_259 (O_259,N_23435,N_24273);
or UO_260 (O_260,N_23180,N_22699);
nand UO_261 (O_261,N_23532,N_23606);
or UO_262 (O_262,N_22881,N_22466);
and UO_263 (O_263,N_23367,N_23923);
nor UO_264 (O_264,N_23537,N_22315);
nor UO_265 (O_265,N_24798,N_22907);
and UO_266 (O_266,N_23860,N_23101);
nand UO_267 (O_267,N_22867,N_22967);
or UO_268 (O_268,N_23318,N_23974);
and UO_269 (O_269,N_22568,N_24290);
nand UO_270 (O_270,N_22377,N_23290);
nor UO_271 (O_271,N_23278,N_22303);
nand UO_272 (O_272,N_23181,N_23123);
nand UO_273 (O_273,N_23174,N_24708);
nand UO_274 (O_274,N_23520,N_23078);
or UO_275 (O_275,N_24136,N_24040);
nand UO_276 (O_276,N_24916,N_22522);
nand UO_277 (O_277,N_23533,N_24956);
nand UO_278 (O_278,N_24142,N_24056);
nor UO_279 (O_279,N_23846,N_23833);
nand UO_280 (O_280,N_22830,N_22461);
nor UO_281 (O_281,N_24953,N_24345);
xnor UO_282 (O_282,N_23075,N_24734);
nor UO_283 (O_283,N_22670,N_23809);
nor UO_284 (O_284,N_24052,N_23785);
and UO_285 (O_285,N_24981,N_23962);
nor UO_286 (O_286,N_22847,N_24044);
nor UO_287 (O_287,N_22762,N_22215);
nor UO_288 (O_288,N_24153,N_24834);
nor UO_289 (O_289,N_23357,N_24712);
xnor UO_290 (O_290,N_24551,N_22206);
nand UO_291 (O_291,N_24652,N_22434);
or UO_292 (O_292,N_22056,N_22096);
and UO_293 (O_293,N_22633,N_24185);
nor UO_294 (O_294,N_22985,N_24247);
and UO_295 (O_295,N_24479,N_22126);
or UO_296 (O_296,N_22893,N_22361);
xnor UO_297 (O_297,N_23762,N_22545);
or UO_298 (O_298,N_24801,N_24113);
nor UO_299 (O_299,N_24510,N_24315);
nand UO_300 (O_300,N_22770,N_23892);
xnor UO_301 (O_301,N_22747,N_23515);
nand UO_302 (O_302,N_22267,N_24667);
nand UO_303 (O_303,N_23060,N_22726);
nor UO_304 (O_304,N_23044,N_22593);
nand UO_305 (O_305,N_24218,N_24332);
or UO_306 (O_306,N_22404,N_22410);
nand UO_307 (O_307,N_22165,N_24335);
xnor UO_308 (O_308,N_22187,N_22453);
nand UO_309 (O_309,N_24166,N_24163);
nand UO_310 (O_310,N_23239,N_24488);
or UO_311 (O_311,N_23399,N_22612);
or UO_312 (O_312,N_22136,N_23404);
and UO_313 (O_313,N_23994,N_23274);
or UO_314 (O_314,N_23360,N_24966);
nor UO_315 (O_315,N_23271,N_23678);
or UO_316 (O_316,N_24673,N_22247);
xor UO_317 (O_317,N_24967,N_24146);
nor UO_318 (O_318,N_24671,N_23067);
nand UO_319 (O_319,N_22336,N_22387);
and UO_320 (O_320,N_24080,N_24058);
and UO_321 (O_321,N_22231,N_24130);
nand UO_322 (O_322,N_24482,N_22354);
nor UO_323 (O_323,N_22093,N_24101);
nand UO_324 (O_324,N_22155,N_22667);
nor UO_325 (O_325,N_22254,N_23032);
and UO_326 (O_326,N_22540,N_24545);
nor UO_327 (O_327,N_24106,N_24534);
nand UO_328 (O_328,N_23243,N_23967);
nor UO_329 (O_329,N_23579,N_24816);
nand UO_330 (O_330,N_24090,N_23462);
nor UO_331 (O_331,N_24229,N_22477);
and UO_332 (O_332,N_23418,N_24234);
or UO_333 (O_333,N_21915,N_22666);
xnor UO_334 (O_334,N_23637,N_21921);
or UO_335 (O_335,N_23295,N_22242);
and UO_336 (O_336,N_22712,N_23261);
and UO_337 (O_337,N_23548,N_22367);
xnor UO_338 (O_338,N_24636,N_22379);
nand UO_339 (O_339,N_24585,N_22925);
nand UO_340 (O_340,N_22552,N_21983);
or UO_341 (O_341,N_23983,N_21936);
nand UO_342 (O_342,N_22312,N_22624);
and UO_343 (O_343,N_24592,N_23450);
and UO_344 (O_344,N_24104,N_24951);
nor UO_345 (O_345,N_22166,N_22261);
nand UO_346 (O_346,N_23709,N_23784);
or UO_347 (O_347,N_22933,N_22341);
nand UO_348 (O_348,N_22549,N_24037);
or UO_349 (O_349,N_22196,N_23878);
or UO_350 (O_350,N_22629,N_22072);
xor UO_351 (O_351,N_23211,N_22765);
nand UO_352 (O_352,N_23161,N_23265);
nor UO_353 (O_353,N_24616,N_23990);
and UO_354 (O_354,N_22193,N_23742);
nor UO_355 (O_355,N_24968,N_21909);
nand UO_356 (O_356,N_22090,N_23233);
or UO_357 (O_357,N_23986,N_21958);
or UO_358 (O_358,N_23416,N_24284);
or UO_359 (O_359,N_23138,N_22446);
or UO_360 (O_360,N_23333,N_22219);
and UO_361 (O_361,N_24765,N_24782);
or UO_362 (O_362,N_21963,N_24372);
and UO_363 (O_363,N_22118,N_21896);
nand UO_364 (O_364,N_21982,N_23253);
nand UO_365 (O_365,N_23480,N_22338);
or UO_366 (O_366,N_23733,N_23734);
nand UO_367 (O_367,N_24285,N_22433);
nand UO_368 (O_368,N_23494,N_23632);
or UO_369 (O_369,N_22484,N_24619);
and UO_370 (O_370,N_22340,N_22289);
nand UO_371 (O_371,N_23715,N_23837);
and UO_372 (O_372,N_23787,N_22786);
and UO_373 (O_373,N_23467,N_23814);
nand UO_374 (O_374,N_23242,N_22386);
or UO_375 (O_375,N_24296,N_22438);
nand UO_376 (O_376,N_23389,N_22063);
and UO_377 (O_377,N_23684,N_22696);
and UO_378 (O_378,N_24063,N_22890);
and UO_379 (O_379,N_23803,N_24846);
nand UO_380 (O_380,N_23033,N_24353);
or UO_381 (O_381,N_24847,N_24242);
and UO_382 (O_382,N_23595,N_24591);
nor UO_383 (O_383,N_23972,N_24443);
nor UO_384 (O_384,N_24745,N_24057);
xnor UO_385 (O_385,N_22271,N_22483);
xnor UO_386 (O_386,N_22482,N_23230);
and UO_387 (O_387,N_22370,N_22577);
and UO_388 (O_388,N_23286,N_22251);
or UO_389 (O_389,N_24722,N_24117);
xnor UO_390 (O_390,N_24450,N_22565);
nor UO_391 (O_391,N_21919,N_23935);
nand UO_392 (O_392,N_22711,N_24799);
or UO_393 (O_393,N_22928,N_23019);
nand UO_394 (O_394,N_23245,N_22124);
nand UO_395 (O_395,N_22833,N_23598);
nand UO_396 (O_396,N_21967,N_22989);
nand UO_397 (O_397,N_23090,N_23248);
or UO_398 (O_398,N_23897,N_22698);
or UO_399 (O_399,N_22724,N_22997);
nor UO_400 (O_400,N_23306,N_24092);
nand UO_401 (O_401,N_24715,N_22360);
nor UO_402 (O_402,N_24046,N_24759);
and UO_403 (O_403,N_22897,N_24920);
or UO_404 (O_404,N_23920,N_24604);
xnor UO_405 (O_405,N_22733,N_24094);
xnor UO_406 (O_406,N_23591,N_22605);
nor UO_407 (O_407,N_23953,N_24776);
nor UO_408 (O_408,N_22994,N_22513);
xor UO_409 (O_409,N_23731,N_24011);
or UO_410 (O_410,N_23796,N_24905);
and UO_411 (O_411,N_24825,N_23336);
and UO_412 (O_412,N_23385,N_24223);
or UO_413 (O_413,N_22432,N_24202);
nor UO_414 (O_414,N_22052,N_24035);
nor UO_415 (O_415,N_22653,N_24049);
nand UO_416 (O_416,N_23283,N_23876);
and UO_417 (O_417,N_24900,N_22821);
nor UO_418 (O_418,N_22279,N_21895);
nand UO_419 (O_419,N_22049,N_24831);
nor UO_420 (O_420,N_23223,N_23139);
nor UO_421 (O_421,N_24666,N_22032);
and UO_422 (O_422,N_24265,N_23137);
and UO_423 (O_423,N_22769,N_22145);
or UO_424 (O_424,N_23364,N_22201);
nor UO_425 (O_425,N_23175,N_24216);
xor UO_426 (O_426,N_22401,N_22086);
nand UO_427 (O_427,N_22763,N_23670);
or UO_428 (O_428,N_23189,N_22889);
and UO_429 (O_429,N_23804,N_23736);
nand UO_430 (O_430,N_23236,N_23947);
nor UO_431 (O_431,N_23378,N_23182);
or UO_432 (O_432,N_23718,N_24492);
and UO_433 (O_433,N_24581,N_24112);
or UO_434 (O_434,N_22601,N_23021);
or UO_435 (O_435,N_24793,N_22977);
or UO_436 (O_436,N_23774,N_23391);
nand UO_437 (O_437,N_24251,N_21981);
and UO_438 (O_438,N_24700,N_23880);
nor UO_439 (O_439,N_22924,N_24271);
and UO_440 (O_440,N_23361,N_23917);
and UO_441 (O_441,N_22597,N_22947);
and UO_442 (O_442,N_22425,N_22868);
or UO_443 (O_443,N_24863,N_22729);
and UO_444 (O_444,N_24654,N_22913);
nand UO_445 (O_445,N_24249,N_22437);
xnor UO_446 (O_446,N_22773,N_24548);
and UO_447 (O_447,N_22573,N_24882);
or UO_448 (O_448,N_22885,N_22467);
nor UO_449 (O_449,N_22603,N_24552);
nor UO_450 (O_450,N_23842,N_22147);
nor UO_451 (O_451,N_23825,N_24802);
nand UO_452 (O_452,N_22673,N_24890);
or UO_453 (O_453,N_23095,N_21978);
or UO_454 (O_454,N_22815,N_24741);
nand UO_455 (O_455,N_23981,N_24380);
nand UO_456 (O_456,N_23257,N_23636);
or UO_457 (O_457,N_24422,N_23116);
and UO_458 (O_458,N_23241,N_22588);
xnor UO_459 (O_459,N_23011,N_24729);
or UO_460 (O_460,N_22641,N_23927);
nor UO_461 (O_461,N_22809,N_24689);
and UO_462 (O_462,N_22870,N_24724);
xor UO_463 (O_463,N_24274,N_22869);
xnor UO_464 (O_464,N_22395,N_22304);
or UO_465 (O_465,N_22501,N_23324);
nand UO_466 (O_466,N_23799,N_23944);
and UO_467 (O_467,N_22243,N_23677);
nand UO_468 (O_468,N_22296,N_24990);
and UO_469 (O_469,N_24582,N_24810);
and UO_470 (O_470,N_24696,N_22544);
or UO_471 (O_471,N_23178,N_22143);
or UO_472 (O_472,N_23703,N_24213);
nor UO_473 (O_473,N_23642,N_23370);
nor UO_474 (O_474,N_24124,N_24197);
nor UO_475 (O_475,N_22311,N_22648);
xnor UO_476 (O_476,N_22154,N_23700);
or UO_477 (O_477,N_22486,N_21960);
nand UO_478 (O_478,N_22277,N_24432);
or UO_479 (O_479,N_23193,N_22113);
nor UO_480 (O_480,N_24408,N_23576);
nand UO_481 (O_481,N_22002,N_24188);
nand UO_482 (O_482,N_23767,N_24358);
and UO_483 (O_483,N_24840,N_24140);
and UO_484 (O_484,N_23952,N_22493);
or UO_485 (O_485,N_23755,N_24896);
or UO_486 (O_486,N_23828,N_23702);
nand UO_487 (O_487,N_22491,N_22179);
or UO_488 (O_488,N_24494,N_24084);
and UO_489 (O_489,N_24645,N_22471);
nand UO_490 (O_490,N_23162,N_24096);
nor UO_491 (O_491,N_22455,N_23959);
or UO_492 (O_492,N_24602,N_23108);
and UO_493 (O_493,N_22211,N_22656);
and UO_494 (O_494,N_23810,N_22026);
nand UO_495 (O_495,N_24025,N_22524);
or UO_496 (O_496,N_22518,N_23201);
or UO_497 (O_497,N_22006,N_23176);
or UO_498 (O_498,N_22351,N_24791);
nand UO_499 (O_499,N_24365,N_23789);
and UO_500 (O_500,N_23940,N_23158);
nand UO_501 (O_501,N_24664,N_23422);
and UO_502 (O_502,N_23481,N_23907);
and UO_503 (O_503,N_24342,N_24181);
nand UO_504 (O_504,N_24283,N_24909);
nand UO_505 (O_505,N_22910,N_23072);
nor UO_506 (O_506,N_23297,N_24127);
nand UO_507 (O_507,N_22827,N_24668);
nor UO_508 (O_508,N_22681,N_21946);
and UO_509 (O_509,N_23043,N_23496);
and UO_510 (O_510,N_23215,N_23778);
nand UO_511 (O_511,N_23048,N_24062);
or UO_512 (O_512,N_24209,N_23603);
nor UO_513 (O_513,N_23226,N_23942);
nor UO_514 (O_514,N_22375,N_22102);
or UO_515 (O_515,N_24702,N_24626);
and UO_516 (O_516,N_23824,N_22170);
nand UO_517 (O_517,N_23505,N_24452);
or UO_518 (O_518,N_23275,N_23053);
and UO_519 (O_519,N_24632,N_24064);
nor UO_520 (O_520,N_23054,N_24784);
nand UO_521 (O_521,N_22087,N_22644);
or UO_522 (O_522,N_24417,N_23224);
nand UO_523 (O_523,N_22628,N_23764);
nand UO_524 (O_524,N_24407,N_22594);
nor UO_525 (O_525,N_23440,N_21975);
and UO_526 (O_526,N_24509,N_22398);
nor UO_527 (O_527,N_23074,N_22427);
and UO_528 (O_528,N_23685,N_22462);
nor UO_529 (O_529,N_22314,N_24447);
xnor UO_530 (O_530,N_23745,N_24998);
nand UO_531 (O_531,N_23658,N_22064);
and UO_532 (O_532,N_23746,N_23873);
and UO_533 (O_533,N_22475,N_24503);
nor UO_534 (O_534,N_24607,N_24637);
nand UO_535 (O_535,N_24861,N_23782);
nand UO_536 (O_536,N_23471,N_23902);
nor UO_537 (O_537,N_23479,N_24159);
or UO_538 (O_538,N_23489,N_22162);
nand UO_539 (O_539,N_24126,N_22151);
and UO_540 (O_540,N_23150,N_23322);
and UO_541 (O_541,N_24149,N_22766);
xor UO_542 (O_542,N_24614,N_22675);
nand UO_543 (O_543,N_22098,N_22188);
nor UO_544 (O_544,N_23238,N_21993);
xor UO_545 (O_545,N_22137,N_23688);
or UO_546 (O_546,N_22355,N_22926);
nand UO_547 (O_547,N_22488,N_22851);
and UO_548 (O_548,N_24520,N_22621);
or UO_549 (O_549,N_22543,N_24961);
nor UO_550 (O_550,N_24815,N_23862);
nand UO_551 (O_551,N_23559,N_22572);
or UO_552 (O_552,N_22973,N_22579);
and UO_553 (O_553,N_23601,N_22507);
nand UO_554 (O_554,N_22397,N_22062);
xor UO_555 (O_555,N_22429,N_23722);
nand UO_556 (O_556,N_23424,N_23928);
nand UO_557 (O_557,N_24977,N_23300);
xor UO_558 (O_558,N_23848,N_24496);
nor UO_559 (O_559,N_23506,N_23046);
or UO_560 (O_560,N_22615,N_22041);
xor UO_561 (O_561,N_22400,N_24811);
nor UO_562 (O_562,N_24313,N_23793);
and UO_563 (O_563,N_24434,N_22986);
and UO_564 (O_564,N_22984,N_22452);
nand UO_565 (O_565,N_22646,N_22874);
nor UO_566 (O_566,N_23403,N_22478);
or UO_567 (O_567,N_23508,N_24212);
nand UO_568 (O_568,N_23497,N_22592);
or UO_569 (O_569,N_23196,N_23237);
or UO_570 (O_570,N_22614,N_23683);
xnor UO_571 (O_571,N_24331,N_23206);
nor UO_572 (O_572,N_22053,N_24017);
nor UO_573 (O_573,N_24133,N_22676);
and UO_574 (O_574,N_24598,N_23384);
nor UO_575 (O_575,N_24138,N_22076);
nand UO_576 (O_576,N_23984,N_21891);
nor UO_577 (O_577,N_23277,N_22094);
xor UO_578 (O_578,N_24118,N_21907);
or UO_579 (O_579,N_24705,N_23546);
nand UO_580 (O_580,N_22385,N_22078);
nand UO_581 (O_581,N_22025,N_22419);
or UO_582 (O_582,N_22185,N_24396);
nand UO_583 (O_583,N_22199,N_24205);
xnor UO_584 (O_584,N_21998,N_22600);
and UO_585 (O_585,N_22734,N_24350);
nor UO_586 (O_586,N_22887,N_24219);
nand UO_587 (O_587,N_22177,N_24609);
or UO_588 (O_588,N_22319,N_24341);
xor UO_589 (O_589,N_23573,N_24856);
and UO_590 (O_590,N_22133,N_22044);
and UO_591 (O_591,N_24258,N_22105);
and UO_592 (O_592,N_23686,N_23589);
or UO_593 (O_593,N_24282,N_24584);
nand UO_594 (O_594,N_22784,N_24681);
or UO_595 (O_595,N_23350,N_23844);
nand UO_596 (O_596,N_22290,N_23587);
and UO_597 (O_597,N_24036,N_24562);
nor UO_598 (O_598,N_22694,N_24932);
xnor UO_599 (O_599,N_24670,N_22660);
or UO_600 (O_600,N_22264,N_22877);
xor UO_601 (O_601,N_24899,N_23380);
or UO_602 (O_602,N_24435,N_22865);
nor UO_603 (O_603,N_23049,N_22232);
or UO_604 (O_604,N_23819,N_22953);
nor UO_605 (O_605,N_23386,N_24939);
nor UO_606 (O_606,N_24406,N_24072);
and UO_607 (O_607,N_24471,N_24262);
nand UO_608 (O_608,N_24110,N_23875);
and UO_609 (O_609,N_22123,N_21973);
nor UO_610 (O_610,N_24309,N_23478);
or UO_611 (O_611,N_21923,N_24491);
nand UO_612 (O_612,N_23014,N_23453);
and UO_613 (O_613,N_22497,N_21996);
and UO_614 (O_614,N_24818,N_23701);
nor UO_615 (O_615,N_22782,N_24211);
xor UO_616 (O_616,N_22708,N_22226);
nand UO_617 (O_617,N_23798,N_24842);
and UO_618 (O_618,N_24038,N_23638);
nor UO_619 (O_619,N_24426,N_22888);
nand UO_620 (O_620,N_23344,N_24944);
or UO_621 (O_621,N_24307,N_23045);
or UO_622 (O_622,N_23061,N_22172);
and UO_623 (O_623,N_22359,N_23347);
and UO_624 (O_624,N_24082,N_24179);
nand UO_625 (O_625,N_23335,N_22829);
or UO_626 (O_626,N_24594,N_24484);
or UO_627 (O_627,N_22741,N_24189);
nor UO_628 (O_628,N_22499,N_22574);
or UO_629 (O_629,N_21976,N_24737);
nor UO_630 (O_630,N_22918,N_22479);
nand UO_631 (O_631,N_24363,N_23616);
nor UO_632 (O_632,N_22008,N_21885);
or UO_633 (O_633,N_24973,N_24191);
and UO_634 (O_634,N_24317,N_23662);
nor UO_635 (O_635,N_22046,N_24982);
nand UO_636 (O_636,N_24469,N_23963);
or UO_637 (O_637,N_23353,N_23488);
xnor UO_638 (O_638,N_24075,N_24725);
nand UO_639 (O_639,N_22816,N_22693);
nand UO_640 (O_640,N_22647,N_24412);
nor UO_641 (O_641,N_23872,N_24889);
nand UO_642 (O_642,N_24735,N_22856);
or UO_643 (O_643,N_22284,N_24256);
and UO_644 (O_644,N_24941,N_24227);
nand UO_645 (O_645,N_22828,N_23882);
nand UO_646 (O_646,N_23486,N_23783);
or UO_647 (O_647,N_24310,N_24013);
or UO_648 (O_648,N_22822,N_21880);
and UO_649 (O_649,N_21965,N_24965);
nor UO_650 (O_650,N_23076,N_22468);
nor UO_651 (O_651,N_24643,N_23558);
nand UO_652 (O_652,N_22683,N_24473);
nand UO_653 (O_653,N_23111,N_24733);
or UO_654 (O_654,N_22752,N_23132);
nor UO_655 (O_655,N_22343,N_24314);
nor UO_656 (O_656,N_24221,N_22198);
nor UO_657 (O_657,N_22227,N_22212);
or UO_658 (O_658,N_24603,N_24912);
and UO_659 (O_659,N_22504,N_23411);
or UO_660 (O_660,N_22084,N_22119);
or UO_661 (O_661,N_24498,N_24622);
or UO_662 (O_662,N_22642,N_23654);
and UO_663 (O_663,N_22300,N_23507);
xor UO_664 (O_664,N_22718,N_22542);
nor UO_665 (O_665,N_22104,N_21949);
and UO_666 (O_666,N_22760,N_22717);
nand UO_667 (O_667,N_23811,N_23395);
nand UO_668 (O_668,N_23913,N_24675);
nor UO_669 (O_669,N_22428,N_22082);
and UO_670 (O_670,N_24768,N_22811);
and UO_671 (O_671,N_24413,N_24516);
or UO_672 (O_672,N_24877,N_24769);
and UO_673 (O_673,N_22498,N_23841);
nor UO_674 (O_674,N_22127,N_22023);
or UO_675 (O_675,N_23708,N_22010);
or UO_676 (O_676,N_23136,N_22347);
nand UO_677 (O_677,N_23393,N_23249);
nor UO_678 (O_678,N_24388,N_24794);
and UO_679 (O_679,N_24194,N_24145);
nand UO_680 (O_680,N_23109,N_24949);
and UO_681 (O_681,N_23288,N_23869);
or UO_682 (O_682,N_24144,N_22412);
and UO_683 (O_683,N_24557,N_22472);
nor UO_684 (O_684,N_23992,N_22901);
and UO_685 (O_685,N_23169,N_24088);
or UO_686 (O_686,N_24170,N_23791);
nand UO_687 (O_687,N_24558,N_24907);
and UO_688 (O_688,N_23457,N_23135);
nand UO_689 (O_689,N_24709,N_22313);
nor UO_690 (O_690,N_22834,N_23419);
or UO_691 (O_691,N_22164,N_22358);
or UO_692 (O_692,N_22328,N_23797);
and UO_693 (O_693,N_22727,N_24822);
xor UO_694 (O_694,N_24911,N_24087);
or UO_695 (O_695,N_22457,N_22442);
nand UO_696 (O_696,N_24480,N_22720);
nor UO_697 (O_697,N_23018,N_23889);
nor UO_698 (O_698,N_23263,N_23217);
and UO_699 (O_699,N_24665,N_24395);
nand UO_700 (O_700,N_22135,N_22704);
nand UO_701 (O_701,N_23834,N_24806);
and UO_702 (O_702,N_23034,N_22561);
and UO_703 (O_703,N_22039,N_24158);
nand UO_704 (O_704,N_22537,N_22494);
nor UO_705 (O_705,N_24489,N_23382);
nand UO_706 (O_706,N_24996,N_23443);
and UO_707 (O_707,N_22510,N_23216);
and UO_708 (O_708,N_24695,N_22256);
and UO_709 (O_709,N_22301,N_23433);
nor UO_710 (O_710,N_22590,N_23960);
xor UO_711 (O_711,N_24493,N_23965);
nor UO_712 (O_712,N_24364,N_24904);
nor UO_713 (O_713,N_22702,N_22714);
or UO_714 (O_714,N_24537,N_22260);
or UO_715 (O_715,N_24536,N_24753);
nor UO_716 (O_716,N_22393,N_22035);
or UO_717 (O_717,N_22456,N_24542);
nand UO_718 (O_718,N_22536,N_23941);
and UO_719 (O_719,N_23037,N_24766);
or UO_720 (O_720,N_22268,N_22715);
or UO_721 (O_721,N_24692,N_22554);
nand UO_722 (O_722,N_23055,N_24620);
or UO_723 (O_723,N_23432,N_22976);
nor UO_724 (O_724,N_24102,N_24937);
and UO_725 (O_725,N_22599,N_24362);
xor UO_726 (O_726,N_21917,N_23001);
and UO_727 (O_727,N_24872,N_22297);
and UO_728 (O_728,N_22018,N_23071);
or UO_729 (O_729,N_24698,N_22661);
xnor UO_730 (O_730,N_24687,N_23870);
nor UO_731 (O_731,N_22631,N_22965);
nor UO_732 (O_732,N_23857,N_22719);
nor UO_733 (O_733,N_23583,N_24086);
xnor UO_734 (O_734,N_22394,N_23534);
and UO_735 (O_735,N_22436,N_24481);
nor UO_736 (O_736,N_22189,N_23113);
or UO_737 (O_737,N_24394,N_22758);
and UO_738 (O_738,N_24634,N_23752);
nand UO_739 (O_739,N_24121,N_21911);
nor UO_740 (O_740,N_23845,N_22020);
nor UO_741 (O_741,N_23321,N_23328);
nor UO_742 (O_742,N_23028,N_22923);
xnor UO_743 (O_743,N_22376,N_21951);
and UO_744 (O_744,N_24987,N_24175);
or UO_745 (O_745,N_24728,N_23203);
nor UO_746 (O_746,N_23822,N_23852);
or UO_747 (O_747,N_22318,N_23149);
and UO_748 (O_748,N_22679,N_24074);
and UO_749 (O_749,N_23473,N_21971);
and UO_750 (O_750,N_24804,N_22810);
or UO_751 (O_751,N_22447,N_23725);
nand UO_752 (O_752,N_23648,N_24099);
and UO_753 (O_753,N_23554,N_23871);
and UO_754 (O_754,N_22596,N_24738);
or UO_755 (O_755,N_24572,N_22611);
nor UO_756 (O_756,N_22141,N_22662);
or UO_757 (O_757,N_24014,N_24114);
and UO_758 (O_758,N_21954,N_23843);
or UO_759 (O_759,N_24655,N_24962);
and UO_760 (O_760,N_24244,N_21952);
and UO_761 (O_761,N_22623,N_22295);
nor UO_762 (O_762,N_23025,N_24680);
xnor UO_763 (O_763,N_23013,N_23402);
and UO_764 (O_764,N_23653,N_24797);
xor UO_765 (O_765,N_23081,N_22700);
nand UO_766 (O_766,N_24546,N_23596);
and UO_767 (O_767,N_24260,N_23168);
nand UO_768 (O_768,N_24858,N_22349);
or UO_769 (O_769,N_22775,N_22936);
nand UO_770 (O_770,N_24502,N_24526);
and UO_771 (O_771,N_24416,N_24590);
nor UO_772 (O_772,N_23663,N_23830);
nor UO_773 (O_773,N_22216,N_22959);
and UO_774 (O_774,N_23210,N_23931);
nand UO_775 (O_775,N_22737,N_23707);
nand UO_776 (O_776,N_21897,N_24182);
nand UO_777 (O_777,N_23664,N_23608);
nand UO_778 (O_778,N_24411,N_22532);
or UO_779 (O_779,N_24055,N_23737);
and UO_780 (O_780,N_23140,N_23832);
nand UO_781 (O_781,N_23387,N_24440);
nor UO_782 (O_782,N_24891,N_23400);
nand UO_783 (O_783,N_22309,N_23995);
nand UO_784 (O_784,N_23893,N_24187);
nor UO_785 (O_785,N_24085,N_22695);
and UO_786 (O_786,N_22241,N_23890);
and UO_787 (O_787,N_22273,N_22306);
or UO_788 (O_788,N_22280,N_22980);
xor UO_789 (O_789,N_24544,N_22539);
and UO_790 (O_790,N_24830,N_23343);
nor UO_791 (O_791,N_24852,N_24268);
or UO_792 (O_792,N_24374,N_23096);
nand UO_793 (O_793,N_22789,N_24659);
nor UO_794 (O_794,N_23643,N_23510);
and UO_795 (O_795,N_23925,N_23268);
nand UO_796 (O_796,N_23777,N_24000);
nand UO_797 (O_797,N_24348,N_22740);
or UO_798 (O_798,N_23317,N_22233);
and UO_799 (O_799,N_22244,N_22904);
nor UO_800 (O_800,N_24326,N_22777);
nor UO_801 (O_801,N_24979,N_24790);
xor UO_802 (O_802,N_23968,N_24969);
nor UO_803 (O_803,N_22380,N_24541);
and UO_804 (O_804,N_23906,N_22929);
xor UO_805 (O_805,N_24109,N_24660);
and UO_806 (O_806,N_22872,N_22911);
xnor UO_807 (O_807,N_24042,N_24312);
and UO_808 (O_808,N_21914,N_23521);
nor UO_809 (O_809,N_22817,N_23773);
or UO_810 (O_810,N_22951,N_22048);
or UO_811 (O_811,N_23186,N_23273);
and UO_812 (O_812,N_22121,N_23854);
xnor UO_813 (O_813,N_22236,N_22886);
xnor UO_814 (O_814,N_24839,N_22589);
nor UO_815 (O_815,N_23689,N_23454);
nand UO_816 (O_816,N_22941,N_24644);
nand UO_817 (O_817,N_23826,N_24403);
or UO_818 (O_818,N_23250,N_24917);
nand UO_819 (O_819,N_23504,N_22991);
nand UO_820 (O_820,N_23969,N_24803);
nand UO_821 (O_821,N_24565,N_23000);
and UO_822 (O_822,N_24091,N_22876);
xnor UO_823 (O_823,N_24183,N_22783);
nand UO_824 (O_824,N_23671,N_21945);
or UO_825 (O_825,N_22399,N_23881);
nor UO_826 (O_826,N_24453,N_22298);
nor UO_827 (O_827,N_22995,N_23909);
nor UO_828 (O_828,N_22040,N_24001);
and UO_829 (O_829,N_24147,N_24864);
nand UO_830 (O_830,N_24618,N_24538);
nor UO_831 (O_831,N_22971,N_22960);
or UO_832 (O_832,N_23763,N_23345);
or UO_833 (O_833,N_22272,N_24220);
and UO_834 (O_834,N_23775,N_24103);
nand UO_835 (O_835,N_24235,N_22689);
nand UO_836 (O_836,N_24885,N_24054);
xor UO_837 (O_837,N_23259,N_23430);
or UO_838 (O_838,N_23341,N_24589);
and UO_839 (O_839,N_24161,N_23989);
nor UO_840 (O_840,N_22981,N_24065);
nor UO_841 (O_841,N_24193,N_22181);
and UO_842 (O_842,N_22797,N_23164);
and UO_843 (O_843,N_22663,N_23246);
nor UO_844 (O_844,N_23690,N_23661);
or UO_845 (O_845,N_22987,N_23166);
xnor UO_846 (O_846,N_23652,N_23185);
and UO_847 (O_847,N_22047,N_23121);
nand UO_848 (O_848,N_23308,N_24628);
nand UO_849 (O_849,N_22892,N_22448);
and UO_850 (O_850,N_23334,N_24302);
nand UO_851 (O_851,N_22652,N_23130);
or UO_852 (O_852,N_22916,N_22055);
nor UO_853 (O_853,N_24669,N_23066);
nand UO_854 (O_854,N_24125,N_21908);
nor UO_855 (O_855,N_22129,N_23209);
nand UO_856 (O_856,N_21995,N_23523);
nand UO_857 (O_857,N_22812,N_24910);
or UO_858 (O_858,N_24878,N_23812);
nand UO_859 (O_859,N_23437,N_23979);
nand UO_860 (O_860,N_22511,N_23195);
xor UO_861 (O_861,N_23853,N_22331);
and UO_862 (O_862,N_23314,N_24959);
nor UO_863 (O_863,N_22940,N_22787);
nor UO_864 (O_864,N_23651,N_22000);
or UO_865 (O_865,N_23980,N_22581);
xor UO_866 (O_866,N_22935,N_22411);
nor UO_867 (O_867,N_23535,N_22210);
nor UO_868 (O_868,N_22075,N_22061);
or UO_869 (O_869,N_23998,N_22571);
and UO_870 (O_870,N_23553,N_24032);
nand UO_871 (O_871,N_23635,N_24656);
nor UO_872 (O_872,N_22723,N_22408);
nor UO_873 (O_873,N_24448,N_23160);
and UO_874 (O_874,N_22664,N_22403);
nor UO_875 (O_875,N_24264,N_22167);
or UO_876 (O_876,N_22962,N_24276);
or UO_877 (O_877,N_22906,N_21953);
or UO_878 (O_878,N_23363,N_24343);
or UO_879 (O_879,N_23484,N_24813);
or UO_880 (O_880,N_24303,N_23719);
xnor UO_881 (O_881,N_24501,N_22205);
and UO_882 (O_882,N_23582,N_23916);
nand UO_883 (O_883,N_23291,N_24828);
nor UO_884 (O_884,N_23086,N_22294);
xnor UO_885 (O_885,N_24483,N_23490);
or UO_886 (O_886,N_22015,N_24869);
or UO_887 (O_887,N_24321,N_23022);
nor UO_888 (O_888,N_23142,N_23613);
and UO_889 (O_889,N_23866,N_23908);
nor UO_890 (O_890,N_23885,N_23572);
nor UO_891 (O_891,N_22586,N_22423);
nor UO_892 (O_892,N_24746,N_23483);
xnor UO_893 (O_893,N_22163,N_23501);
and UO_894 (O_894,N_22153,N_22684);
or UO_895 (O_895,N_23540,N_23247);
nor UO_896 (O_896,N_23128,N_24824);
xnor UO_897 (O_897,N_24936,N_24154);
xor UO_898 (O_898,N_24777,N_24195);
xnor UO_899 (O_899,N_23080,N_22138);
or UO_900 (O_900,N_24499,N_23127);
nand UO_901 (O_901,N_24773,N_23040);
or UO_902 (O_902,N_21912,N_24751);
nor UO_903 (O_903,N_23524,N_23821);
or UO_904 (O_904,N_22908,N_23303);
nor UO_905 (O_905,N_24230,N_24377);
nor UO_906 (O_906,N_23134,N_23611);
and UO_907 (O_907,N_22416,N_23721);
nand UO_908 (O_908,N_22778,N_23401);
and UO_909 (O_909,N_23950,N_24137);
nand UO_910 (O_910,N_23097,N_24421);
nor UO_911 (O_911,N_23412,N_23499);
or UO_912 (O_912,N_24886,N_22424);
nand UO_913 (O_913,N_23163,N_23781);
and UO_914 (O_914,N_21941,N_23699);
or UO_915 (O_915,N_22183,N_22871);
nor UO_916 (O_916,N_22125,N_24449);
nor UO_917 (O_917,N_24192,N_22274);
xnor UO_918 (O_918,N_23599,N_24295);
nand UO_919 (O_919,N_24259,N_23790);
nand UO_920 (O_920,N_23538,N_22500);
nand UO_921 (O_921,N_22074,N_23622);
nor UO_922 (O_922,N_22921,N_23220);
nor UO_923 (O_923,N_22258,N_23213);
or UO_924 (O_924,N_24355,N_24779);
and UO_925 (O_925,N_23368,N_22459);
and UO_926 (O_926,N_23173,N_23630);
nand UO_927 (O_927,N_24324,N_23009);
or UO_928 (O_928,N_22691,N_24366);
nand UO_929 (O_929,N_24462,N_22128);
nor UO_930 (O_930,N_24744,N_24921);
nand UO_931 (O_931,N_23912,N_22071);
and UO_932 (O_932,N_23858,N_22317);
nand UO_933 (O_933,N_21997,N_23511);
and UO_934 (O_934,N_23415,N_24131);
nor UO_935 (O_935,N_24903,N_24288);
nor UO_936 (O_936,N_24686,N_23697);
and UO_937 (O_937,N_23516,N_24894);
and UO_938 (O_938,N_24930,N_22852);
and UO_939 (O_939,N_24378,N_23659);
and UO_940 (O_940,N_23083,N_23351);
nor UO_941 (O_941,N_23667,N_24989);
and UO_942 (O_942,N_23094,N_23279);
and UO_943 (O_943,N_22903,N_23218);
or UO_944 (O_944,N_21934,N_22583);
nor UO_945 (O_945,N_22582,N_24415);
and UO_946 (O_946,N_23146,N_22307);
nand UO_947 (O_947,N_22218,N_24061);
or UO_948 (O_948,N_24697,N_24027);
and UO_949 (O_949,N_24409,N_22618);
or UO_950 (O_950,N_22982,N_23088);
or UO_951 (O_951,N_22818,N_23884);
and UO_952 (O_952,N_23961,N_21938);
xnor UO_953 (O_953,N_23645,N_23235);
or UO_954 (O_954,N_24186,N_22037);
or UO_955 (O_955,N_22649,N_23619);
xnor UO_956 (O_956,N_23451,N_22958);
xnor UO_957 (O_957,N_23861,N_23838);
nand UO_958 (O_958,N_24292,N_23272);
nand UO_959 (O_959,N_22793,N_21968);
nand UO_960 (O_960,N_21922,N_22122);
nor UO_961 (O_961,N_24155,N_24004);
or UO_962 (O_962,N_23937,N_23605);
nand UO_963 (O_963,N_23472,N_22293);
xor UO_964 (O_964,N_22173,N_22038);
nand UO_965 (O_965,N_24459,N_22363);
nand UO_966 (O_966,N_24748,N_23800);
nand UO_967 (O_967,N_24384,N_24316);
and UO_968 (O_968,N_22474,N_23199);
xor UO_969 (O_969,N_23313,N_24820);
nand UO_970 (O_970,N_24029,N_23682);
and UO_971 (O_971,N_22208,N_23390);
nor UO_972 (O_972,N_24543,N_22014);
or UO_973 (O_973,N_22857,N_23758);
or UO_974 (O_974,N_23750,N_23089);
nor UO_975 (O_975,N_24711,N_24076);
and UO_976 (O_976,N_23770,N_24008);
nand UO_977 (O_977,N_23330,N_23801);
and UO_978 (O_978,N_24770,N_21947);
nand UO_979 (O_979,N_22530,N_24009);
nor UO_980 (O_980,N_24931,N_24047);
or UO_981 (O_981,N_24942,N_23031);
nand UO_982 (O_982,N_23904,N_22146);
and UO_983 (O_983,N_24012,N_24105);
nand UO_984 (O_984,N_23461,N_22392);
nand UO_985 (O_985,N_23212,N_23442);
and UO_986 (O_986,N_23669,N_24788);
and UO_987 (O_987,N_24252,N_24508);
nor UO_988 (O_988,N_22895,N_22186);
xor UO_989 (O_989,N_23996,N_21955);
and UO_990 (O_990,N_23298,N_22107);
nand UO_991 (O_991,N_23369,N_24506);
and UO_992 (O_992,N_24250,N_23748);
xnor UO_993 (O_993,N_24972,N_24881);
and UO_994 (O_994,N_22519,N_24955);
or UO_995 (O_995,N_24460,N_24873);
and UO_996 (O_996,N_23476,N_22325);
nand UO_997 (O_997,N_22932,N_21905);
nand UO_998 (O_998,N_24003,N_23943);
and UO_999 (O_999,N_23529,N_23482);
nor UO_1000 (O_1000,N_22238,N_24593);
or UO_1001 (O_1001,N_23855,N_23079);
and UO_1002 (O_1002,N_24868,N_23337);
or UO_1003 (O_1003,N_22665,N_24928);
or UO_1004 (O_1004,N_24792,N_22067);
or UO_1005 (O_1005,N_22324,N_22160);
nor UO_1006 (O_1006,N_23375,N_23756);
nor UO_1007 (O_1007,N_24983,N_23693);
or UO_1008 (O_1008,N_22374,N_22808);
xor UO_1009 (O_1009,N_21894,N_24504);
xor UO_1010 (O_1010,N_24610,N_24730);
and UO_1011 (O_1011,N_23541,N_23851);
nand UO_1012 (O_1012,N_23260,N_24336);
or UO_1013 (O_1013,N_22993,N_22184);
and UO_1014 (O_1014,N_24635,N_23050);
and UO_1015 (O_1015,N_21888,N_22100);
xor UO_1016 (O_1016,N_23309,N_22021);
or UO_1017 (O_1017,N_21920,N_23007);
nor UO_1018 (O_1018,N_22813,N_24207);
nor UO_1019 (O_1019,N_23085,N_22066);
xnor UO_1020 (O_1020,N_23891,N_24532);
and UO_1021 (O_1021,N_22176,N_24141);
xor UO_1022 (O_1022,N_23536,N_24938);
nor UO_1023 (O_1023,N_23057,N_22169);
nand UO_1024 (O_1024,N_24028,N_22687);
nand UO_1025 (O_1025,N_22364,N_24100);
nor UO_1026 (O_1026,N_24446,N_22332);
nand UO_1027 (O_1027,N_24837,N_24970);
and UO_1028 (O_1028,N_23712,N_22791);
nor UO_1029 (O_1029,N_22470,N_24240);
or UO_1030 (O_1030,N_24821,N_22801);
xnor UO_1031 (O_1031,N_23421,N_23131);
nor UO_1032 (O_1032,N_24946,N_24455);
or UO_1033 (O_1033,N_24742,N_21994);
nand UO_1034 (O_1034,N_24016,N_23547);
nor UO_1035 (O_1035,N_21962,N_23999);
nand UO_1036 (O_1036,N_24199,N_22095);
xor UO_1037 (O_1037,N_23728,N_23976);
nand UO_1038 (O_1038,N_22515,N_23093);
and UO_1039 (O_1039,N_22855,N_22772);
nor UO_1040 (O_1040,N_24649,N_24992);
xnor UO_1041 (O_1041,N_24555,N_24423);
nand UO_1042 (O_1042,N_24232,N_22838);
and UO_1043 (O_1043,N_23204,N_23646);
nand UO_1044 (O_1044,N_22677,N_24787);
or UO_1045 (O_1045,N_23593,N_23439);
nand UO_1046 (O_1046,N_23145,N_23528);
or UO_1047 (O_1047,N_23463,N_23949);
nand UO_1048 (O_1048,N_24629,N_22938);
or UO_1049 (O_1049,N_22541,N_23751);
or UO_1050 (O_1050,N_24445,N_23383);
or UO_1051 (O_1051,N_23706,N_23377);
or UO_1052 (O_1052,N_22841,N_22278);
xnor UO_1053 (O_1053,N_24749,N_22912);
nand UO_1054 (O_1054,N_24752,N_21875);
xnor UO_1055 (O_1055,N_23899,N_24914);
nor UO_1056 (O_1056,N_23526,N_22706);
nand UO_1057 (O_1057,N_21984,N_23198);
or UO_1058 (O_1058,N_23170,N_23410);
nand UO_1059 (O_1059,N_23639,N_24344);
nor UO_1060 (O_1060,N_23063,N_23561);
nor UO_1061 (O_1061,N_23460,N_22657);
and UO_1062 (O_1062,N_24512,N_23740);
nand UO_1063 (O_1063,N_22846,N_23003);
nand UO_1064 (O_1064,N_23802,N_22943);
and UO_1065 (O_1065,N_23311,N_22326);
and UO_1066 (O_1066,N_23059,N_23514);
or UO_1067 (O_1067,N_21913,N_22609);
nand UO_1068 (O_1068,N_24006,N_24071);
xor UO_1069 (O_1069,N_24337,N_22806);
and UO_1070 (O_1070,N_24855,N_23323);
or UO_1071 (O_1071,N_24024,N_22825);
or UO_1072 (O_1072,N_23788,N_22083);
and UO_1073 (O_1073,N_24527,N_21980);
nor UO_1074 (O_1074,N_22944,N_23939);
or UO_1075 (O_1075,N_24940,N_23786);
nor UO_1076 (O_1076,N_22156,N_21901);
and UO_1077 (O_1077,N_23666,N_24373);
nand UO_1078 (O_1078,N_21979,N_22054);
nor UO_1079 (O_1079,N_22460,N_22954);
nand UO_1080 (O_1080,N_23585,N_22175);
and UO_1081 (O_1081,N_24045,N_22323);
and UO_1082 (O_1082,N_23970,N_22330);
nor UO_1083 (O_1083,N_21939,N_23144);
xnor UO_1084 (O_1084,N_23299,N_24995);
nor UO_1085 (O_1085,N_24719,N_22213);
nand UO_1086 (O_1086,N_23266,N_23954);
and UO_1087 (O_1087,N_24444,N_24349);
and UO_1088 (O_1088,N_24599,N_22550);
and UO_1089 (O_1089,N_22992,N_24167);
nand UO_1090 (O_1090,N_24908,N_24933);
nor UO_1091 (O_1091,N_24835,N_21933);
or UO_1092 (O_1092,N_23550,N_22073);
nor UO_1093 (O_1093,N_22286,N_24476);
and UO_1094 (O_1094,N_23064,N_23747);
nand UO_1095 (O_1095,N_23436,N_23827);
nor UO_1096 (O_1096,N_23154,N_22207);
or UO_1097 (O_1097,N_21878,N_22975);
or UO_1098 (O_1098,N_22443,N_23676);
or UO_1099 (O_1099,N_24156,N_24053);
nand UO_1100 (O_1100,N_22650,N_23459);
nand UO_1101 (O_1101,N_23569,N_22748);
nand UO_1102 (O_1102,N_22144,N_22445);
nand UO_1103 (O_1103,N_23936,N_23396);
nor UO_1104 (O_1104,N_24964,N_24458);
or UO_1105 (O_1105,N_23517,N_24707);
nor UO_1106 (O_1106,N_22131,N_23692);
xnor UO_1107 (O_1107,N_23179,N_22655);
xnor UO_1108 (O_1108,N_22496,N_22739);
and UO_1109 (O_1109,N_22180,N_22346);
and UO_1110 (O_1110,N_24997,N_23794);
and UO_1111 (O_1111,N_24246,N_24322);
or UO_1112 (O_1112,N_24497,N_23525);
or UO_1113 (O_1113,N_22007,N_24383);
and UO_1114 (O_1114,N_22626,N_22234);
nand UO_1115 (O_1115,N_22753,N_24650);
xor UO_1116 (O_1116,N_21900,N_24241);
and UO_1117 (O_1117,N_23329,N_24164);
or UO_1118 (O_1118,N_23768,N_22983);
and UO_1119 (O_1119,N_22622,N_24405);
or UO_1120 (O_1120,N_22150,N_23092);
or UO_1121 (O_1121,N_24339,N_24651);
or UO_1122 (O_1122,N_22795,N_23649);
or UO_1123 (O_1123,N_24710,N_22974);
xnor UO_1124 (O_1124,N_22506,N_22678);
and UO_1125 (O_1125,N_22682,N_23426);
and UO_1126 (O_1126,N_23694,N_22781);
nor UO_1127 (O_1127,N_23629,N_22476);
nor UO_1128 (O_1128,N_23634,N_24030);
xor UO_1129 (O_1129,N_22204,N_24647);
nor UO_1130 (O_1130,N_24892,N_23441);
and UO_1131 (O_1131,N_24693,N_24505);
nand UO_1132 (O_1132,N_24376,N_23287);
nand UO_1133 (O_1133,N_24333,N_24601);
or UO_1134 (O_1134,N_23946,N_23816);
nand UO_1135 (O_1135,N_21957,N_23352);
or UO_1136 (O_1136,N_24880,N_23711);
and UO_1137 (O_1137,N_23340,N_24826);
and UO_1138 (O_1138,N_23107,N_22454);
and UO_1139 (O_1139,N_24352,N_22366);
nor UO_1140 (O_1140,N_23205,N_22955);
xnor UO_1141 (O_1141,N_23129,N_23371);
and UO_1142 (O_1142,N_23792,N_24684);
and UO_1143 (O_1143,N_21876,N_24897);
nor UO_1144 (O_1144,N_24298,N_23627);
nand UO_1145 (O_1145,N_23190,N_22564);
or UO_1146 (O_1146,N_23957,N_24929);
xor UO_1147 (O_1147,N_23542,N_21926);
or UO_1148 (O_1148,N_22968,N_23267);
nand UO_1149 (O_1149,N_23221,N_22839);
xor UO_1150 (O_1150,N_23849,N_24895);
or UO_1151 (O_1151,N_23354,N_23765);
nand UO_1152 (O_1152,N_21929,N_23192);
xnor UO_1153 (O_1153,N_23818,N_22117);
nand UO_1154 (O_1154,N_22742,N_24706);
or UO_1155 (O_1155,N_23753,N_22305);
nor UO_1156 (O_1156,N_23580,N_22899);
nand UO_1157 (O_1157,N_24245,N_22891);
nor UO_1158 (O_1158,N_23552,N_23695);
or UO_1159 (O_1159,N_22383,N_22533);
and UO_1160 (O_1160,N_21961,N_23592);
nand UO_1161 (O_1161,N_24817,N_23531);
and UO_1162 (O_1162,N_24957,N_24424);
or UO_1163 (O_1163,N_24190,N_24301);
and UO_1164 (O_1164,N_23405,N_22414);
or UO_1165 (O_1165,N_24224,N_22643);
or UO_1166 (O_1166,N_22373,N_22728);
nor UO_1167 (O_1167,N_24679,N_23156);
nand UO_1168 (O_1168,N_23813,N_24862);
or UO_1169 (O_1169,N_21956,N_22859);
and UO_1170 (O_1170,N_22329,N_23016);
nor UO_1171 (O_1171,N_23570,N_24330);
or UO_1172 (O_1172,N_24236,N_23835);
and UO_1173 (O_1173,N_23251,N_24069);
nand UO_1174 (O_1174,N_24583,N_22927);
nand UO_1175 (O_1175,N_22616,N_24958);
nor UO_1176 (O_1176,N_22751,N_24263);
nand UO_1177 (O_1177,N_22972,N_24767);
nor UO_1178 (O_1178,N_24605,N_22746);
nand UO_1179 (O_1179,N_22112,N_21928);
nand UO_1180 (O_1180,N_23675,N_23125);
and UO_1181 (O_1181,N_24764,N_23305);
and UO_1182 (O_1182,N_24070,N_23618);
nand UO_1183 (O_1183,N_24022,N_24399);
xnor UO_1184 (O_1184,N_23681,N_22362);
nand UO_1185 (O_1185,N_23705,N_23425);
or UO_1186 (O_1186,N_24132,N_22514);
or UO_1187 (O_1187,N_23153,N_22217);
xnor UO_1188 (O_1188,N_22909,N_24789);
or UO_1189 (O_1189,N_24699,N_22337);
nand UO_1190 (O_1190,N_23614,N_24067);
nor UO_1191 (O_1191,N_23284,N_22949);
nand UO_1192 (O_1192,N_23444,N_24359);
nand UO_1193 (O_1193,N_21985,N_24866);
or UO_1194 (O_1194,N_22029,N_24162);
nor UO_1195 (O_1195,N_22024,N_22837);
or UO_1196 (O_1196,N_22710,N_22861);
xnor UO_1197 (O_1197,N_22421,N_23027);
and UO_1198 (O_1198,N_24439,N_24874);
nand UO_1199 (O_1199,N_23991,N_21918);
nand UO_1200 (O_1200,N_22705,N_24177);
nand UO_1201 (O_1201,N_23438,N_23285);
and UO_1202 (O_1202,N_24019,N_23710);
nor UO_1203 (O_1203,N_24277,N_24404);
nor UO_1204 (O_1204,N_24867,N_24690);
xor UO_1205 (O_1205,N_22310,N_23100);
and UO_1206 (O_1206,N_22703,N_22613);
and UO_1207 (O_1207,N_24595,N_24007);
nand UO_1208 (O_1208,N_24812,N_22344);
or UO_1209 (O_1209,N_23487,N_24999);
or UO_1210 (O_1210,N_23301,N_22848);
nand UO_1211 (O_1211,N_24524,N_24623);
or UO_1212 (O_1212,N_21898,N_24827);
xnor UO_1213 (O_1213,N_22774,N_23929);
nand UO_1214 (O_1214,N_24174,N_21881);
and UO_1215 (O_1215,N_24915,N_23584);
nor UO_1216 (O_1216,N_22785,N_22505);
nand UO_1217 (O_1217,N_24427,N_22799);
xor UO_1218 (O_1218,N_23294,N_23911);
or UO_1219 (O_1219,N_23464,N_24168);
xor UO_1220 (O_1220,N_24661,N_24980);
nand UO_1221 (O_1221,N_24954,N_24390);
and UO_1222 (O_1222,N_24419,N_21969);
nand UO_1223 (O_1223,N_24617,N_24556);
xor UO_1224 (O_1224,N_22223,N_24606);
nor UO_1225 (O_1225,N_23417,N_23512);
nand UO_1226 (O_1226,N_24034,N_22803);
xnor UO_1227 (O_1227,N_22730,N_23831);
xnor UO_1228 (O_1228,N_22407,N_22619);
nor UO_1229 (O_1229,N_24500,N_24023);
nor UO_1230 (O_1230,N_23456,N_23633);
or UO_1231 (O_1231,N_24683,N_23229);
nand UO_1232 (O_1232,N_22116,N_22807);
nor UO_1233 (O_1233,N_23735,N_22802);
nor UO_1234 (O_1234,N_24833,N_24203);
nand UO_1235 (O_1235,N_24876,N_24465);
nand UO_1236 (O_1236,N_24368,N_24233);
or UO_1237 (O_1237,N_24078,N_23898);
xor UO_1238 (O_1238,N_24758,N_24157);
or UO_1239 (O_1239,N_24123,N_23973);
nand UO_1240 (O_1240,N_24115,N_23012);
nand UO_1241 (O_1241,N_23015,N_22451);
nand UO_1242 (O_1242,N_23896,N_24577);
nand UO_1243 (O_1243,N_22527,N_23839);
nor UO_1244 (O_1244,N_22381,N_24253);
nor UO_1245 (O_1245,N_23148,N_24836);
nor UO_1246 (O_1246,N_24677,N_22139);
xor UO_1247 (O_1247,N_22591,N_22065);
and UO_1248 (O_1248,N_22896,N_23864);
nor UO_1249 (O_1249,N_23115,N_24838);
nor UO_1250 (O_1250,N_23106,N_23448);
and UO_1251 (O_1251,N_24853,N_24714);
nand UO_1252 (O_1252,N_24180,N_22800);
and UO_1253 (O_1253,N_22485,N_22804);
nand UO_1254 (O_1254,N_23761,N_23493);
or UO_1255 (O_1255,N_22796,N_22322);
nor UO_1256 (O_1256,N_23829,N_23052);
xor UO_1257 (O_1257,N_24898,N_22013);
nor UO_1258 (O_1258,N_24398,N_23513);
nand UO_1259 (O_1259,N_24464,N_24513);
and UO_1260 (O_1260,N_24428,N_22220);
xor UO_1261 (O_1261,N_23214,N_22079);
xnor UO_1262 (O_1262,N_24726,N_22805);
nor UO_1263 (O_1263,N_22952,N_22405);
or UO_1264 (O_1264,N_23159,N_24128);
nor UO_1265 (O_1265,N_24596,N_24226);
nor UO_1266 (O_1266,N_22878,N_24278);
or UO_1267 (O_1267,N_23727,N_22563);
or UO_1268 (O_1268,N_24327,N_22697);
nand UO_1269 (O_1269,N_24048,N_24567);
xnor UO_1270 (O_1270,N_22257,N_22788);
or UO_1271 (O_1271,N_24760,N_23657);
or UO_1272 (O_1272,N_23124,N_22287);
nor UO_1273 (O_1273,N_24588,N_24561);
nand UO_1274 (O_1274,N_24774,N_24642);
or UO_1275 (O_1275,N_24095,N_24963);
nand UO_1276 (O_1276,N_24461,N_23563);
and UO_1277 (O_1277,N_24865,N_22875);
and UO_1278 (O_1278,N_23914,N_23458);
nand UO_1279 (O_1279,N_22996,N_24351);
nor UO_1280 (O_1280,N_23820,N_24731);
and UO_1281 (O_1281,N_24574,N_23105);
xnor UO_1282 (O_1282,N_22835,N_24991);
nor UO_1283 (O_1283,N_22263,N_24051);
nand UO_1284 (O_1284,N_24560,N_24723);
and UO_1285 (O_1285,N_22578,N_21903);
or UO_1286 (O_1286,N_23539,N_23919);
and UO_1287 (O_1287,N_23231,N_23219);
nand UO_1288 (O_1288,N_23232,N_24578);
nand UO_1289 (O_1289,N_22559,N_23269);
nand UO_1290 (O_1290,N_21948,N_22779);
or UO_1291 (O_1291,N_24477,N_23102);
or UO_1292 (O_1292,N_22736,N_24843);
and UO_1293 (O_1293,N_22866,N_23302);
nor UO_1294 (O_1294,N_23945,N_23625);
xnor UO_1295 (O_1295,N_24653,N_24641);
xnor UO_1296 (O_1296,N_22060,N_22576);
and UO_1297 (O_1297,N_21932,N_22245);
xor UO_1298 (O_1298,N_23655,N_24717);
nor UO_1299 (O_1299,N_24703,N_24184);
xor UO_1300 (O_1300,N_24713,N_24755);
and UO_1301 (O_1301,N_24357,N_24611);
nand UO_1302 (O_1302,N_23626,N_24918);
nor UO_1303 (O_1303,N_23452,N_22224);
or UO_1304 (O_1304,N_23597,N_21889);
or UO_1305 (O_1305,N_22202,N_24338);
xor UO_1306 (O_1306,N_22850,N_24279);
nor UO_1307 (O_1307,N_24243,N_23581);
and UO_1308 (O_1308,N_23955,N_24658);
nor UO_1309 (O_1309,N_22103,N_22161);
xnor UO_1310 (O_1310,N_24267,N_22158);
nor UO_1311 (O_1311,N_24436,N_24347);
nor UO_1312 (O_1312,N_23455,N_22378);
or UO_1313 (O_1313,N_23503,N_23757);
nor UO_1314 (O_1314,N_22221,N_23339);
or UO_1315 (O_1315,N_22109,N_22754);
xnor UO_1316 (O_1316,N_22668,N_21884);
and UO_1317 (O_1317,N_23141,N_24237);
nand UO_1318 (O_1318,N_23065,N_23933);
nor UO_1319 (O_1319,N_23485,N_24300);
nor UO_1320 (O_1320,N_23571,N_23624);
and UO_1321 (O_1321,N_22365,N_23808);
and UO_1322 (O_1322,N_22690,N_23252);
nor UO_1323 (O_1323,N_24495,N_22302);
and UO_1324 (O_1324,N_22970,N_23915);
nand UO_1325 (O_1325,N_23958,N_22230);
nand UO_1326 (O_1326,N_24079,N_23604);
or UO_1327 (O_1327,N_24563,N_22845);
or UO_1328 (O_1328,N_23087,N_24887);
or UO_1329 (O_1329,N_24043,N_22864);
nand UO_1330 (O_1330,N_23817,N_22585);
nor UO_1331 (O_1331,N_24010,N_23545);
xor UO_1332 (O_1332,N_24522,N_23359);
and UO_1333 (O_1333,N_22858,N_23202);
nor UO_1334 (O_1334,N_22516,N_24402);
nand UO_1335 (O_1335,N_22308,N_22115);
or UO_1336 (O_1336,N_22942,N_22853);
nand UO_1337 (O_1337,N_22534,N_23338);
nand UO_1338 (O_1338,N_23924,N_24587);
nand UO_1339 (O_1339,N_22292,N_22148);
nor UO_1340 (O_1340,N_24988,N_22480);
and UO_1341 (O_1341,N_23228,N_24638);
nor UO_1342 (O_1342,N_24410,N_22033);
xnor UO_1343 (O_1343,N_23588,N_22159);
and UO_1344 (O_1344,N_23356,N_24474);
nand UO_1345 (O_1345,N_24305,N_22759);
nor UO_1346 (O_1346,N_24554,N_23413);
and UO_1347 (O_1347,N_22521,N_23104);
nor UO_1348 (O_1348,N_23749,N_22990);
or UO_1349 (O_1349,N_22823,N_23741);
nand UO_1350 (O_1350,N_23152,N_22894);
nor UO_1351 (O_1351,N_24859,N_24754);
or UO_1352 (O_1352,N_24108,N_23567);
xnor UO_1353 (O_1353,N_22402,N_24884);
and UO_1354 (O_1354,N_24761,N_24662);
and UO_1355 (O_1355,N_22157,N_24923);
nor UO_1356 (O_1356,N_24985,N_23474);
xor UO_1357 (O_1357,N_24306,N_21924);
nor UO_1358 (O_1358,N_22632,N_22027);
nor UO_1359 (O_1359,N_22222,N_22068);
nor UO_1360 (O_1360,N_23617,N_23863);
or UO_1361 (O_1361,N_22931,N_23993);
or UO_1362 (O_1362,N_24848,N_22750);
xor UO_1363 (O_1363,N_24672,N_23562);
and UO_1364 (O_1364,N_23039,N_24523);
and UO_1365 (O_1365,N_23760,N_23568);
nand UO_1366 (O_1366,N_23469,N_24060);
and UO_1367 (O_1367,N_24586,N_22659);
nand UO_1368 (O_1368,N_22178,N_22057);
nand UO_1369 (O_1369,N_23877,N_24111);
nor UO_1370 (O_1370,N_23244,N_24786);
nand UO_1371 (O_1371,N_22580,N_24569);
xnor UO_1372 (O_1372,N_22627,N_22814);
xor UO_1373 (O_1373,N_23332,N_24254);
nor UO_1374 (O_1374,N_24625,N_24718);
and UO_1375 (O_1375,N_24002,N_24785);
nor UO_1376 (O_1376,N_22097,N_22764);
nor UO_1377 (O_1377,N_22508,N_23665);
nor UO_1378 (O_1378,N_23502,N_23836);
or UO_1379 (O_1379,N_23926,N_22566);
and UO_1380 (O_1380,N_23932,N_24200);
nor UO_1381 (O_1381,N_22945,N_23660);
nor UO_1382 (O_1382,N_24371,N_23167);
and UO_1383 (O_1383,N_24832,N_22745);
nand UO_1384 (O_1384,N_22339,N_23327);
and UO_1385 (O_1385,N_24922,N_24739);
and UO_1386 (O_1386,N_22356,N_21910);
or UO_1387 (O_1387,N_22528,N_22880);
and UO_1388 (O_1388,N_22368,N_24297);
nand UO_1389 (O_1389,N_23856,N_23805);
nor UO_1390 (O_1390,N_24841,N_24490);
or UO_1391 (O_1391,N_22842,N_24266);
nand UO_1392 (O_1392,N_22085,N_22009);
xor UO_1393 (O_1393,N_23704,N_22132);
and UO_1394 (O_1394,N_23112,N_22050);
and UO_1395 (O_1395,N_24215,N_23739);
or UO_1396 (O_1396,N_22771,N_22557);
or UO_1397 (O_1397,N_23446,N_22320);
nand UO_1398 (O_1398,N_24875,N_24328);
xnor UO_1399 (O_1399,N_22042,N_23551);
or UO_1400 (O_1400,N_22070,N_24169);
nor UO_1401 (O_1401,N_23910,N_24993);
or UO_1402 (O_1402,N_22721,N_24823);
nor UO_1403 (O_1403,N_24571,N_23495);
nor UO_1404 (O_1404,N_24576,N_24540);
and UO_1405 (O_1405,N_22487,N_23056);
nor UO_1406 (O_1406,N_23331,N_22430);
nor UO_1407 (O_1407,N_24400,N_24971);
or UO_1408 (O_1408,N_24646,N_22755);
or UO_1409 (O_1409,N_22043,N_23868);
nor UO_1410 (O_1410,N_22019,N_23840);
xor UO_1411 (O_1411,N_24369,N_23376);
and UO_1412 (O_1412,N_24222,N_22840);
xor UO_1413 (O_1413,N_24854,N_22357);
and UO_1414 (O_1414,N_23004,N_24631);
or UO_1415 (O_1415,N_24674,N_22192);
nor UO_1416 (O_1416,N_23082,N_23865);
and UO_1417 (O_1417,N_22140,N_23264);
or UO_1418 (O_1418,N_23008,N_24239);
and UO_1419 (O_1419,N_24454,N_23254);
nand UO_1420 (O_1420,N_24031,N_23276);
nor UO_1421 (O_1421,N_22239,N_23281);
nor UO_1422 (O_1422,N_22469,N_24844);
nand UO_1423 (O_1423,N_23110,N_23631);
or UO_1424 (O_1424,N_22946,N_23270);
or UO_1425 (O_1425,N_22275,N_23988);
or UO_1426 (O_1426,N_21925,N_23543);
nand UO_1427 (O_1427,N_24217,N_22228);
or UO_1428 (O_1428,N_24387,N_24525);
nand UO_1429 (O_1429,N_23492,N_23398);
xor UO_1430 (O_1430,N_22948,N_24437);
nand UO_1431 (O_1431,N_23026,N_23051);
or UO_1432 (O_1432,N_23754,N_24026);
and UO_1433 (O_1433,N_23280,N_22266);
xnor UO_1434 (O_1434,N_22111,N_22979);
and UO_1435 (O_1435,N_22134,N_24456);
nor UO_1436 (O_1436,N_23470,N_22862);
xor UO_1437 (O_1437,N_23348,N_24059);
or UO_1438 (O_1438,N_22844,N_22640);
or UO_1439 (O_1439,N_22353,N_22335);
or UO_1440 (O_1440,N_23191,N_22722);
and UO_1441 (O_1441,N_23036,N_23407);
nor UO_1442 (O_1442,N_24573,N_23644);
and UO_1443 (O_1443,N_22299,N_22265);
nor UO_1444 (O_1444,N_24323,N_23208);
and UO_1445 (O_1445,N_24553,N_23544);
and UO_1446 (O_1446,N_22645,N_22490);
or UO_1447 (O_1447,N_24814,N_22350);
xor UO_1448 (O_1448,N_24566,N_24763);
nor UO_1449 (O_1449,N_23122,N_23069);
and UO_1450 (O_1450,N_24391,N_22248);
xnor UO_1451 (O_1451,N_24116,N_23859);
or UO_1452 (O_1452,N_22517,N_22229);
nand UO_1453 (O_1453,N_24517,N_22214);
and UO_1454 (O_1454,N_22639,N_22371);
nor UO_1455 (O_1455,N_22556,N_23227);
nand UO_1456 (O_1456,N_24947,N_23325);
nor UO_1457 (O_1457,N_23867,N_24150);
nor UO_1458 (O_1458,N_23590,N_22195);
nor UO_1459 (O_1459,N_23143,N_24098);
nand UO_1460 (O_1460,N_24857,N_24039);
or UO_1461 (O_1461,N_24943,N_22114);
or UO_1462 (O_1462,N_24535,N_24721);
or UO_1463 (O_1463,N_22512,N_23098);
and UO_1464 (O_1464,N_23171,N_21964);
nor UO_1465 (O_1465,N_23289,N_23729);
nand UO_1466 (O_1466,N_24299,N_21904);
and UO_1467 (O_1467,N_22259,N_22707);
nor UO_1468 (O_1468,N_24913,N_24639);
nand UO_1469 (O_1469,N_23172,N_22045);
nand UO_1470 (O_1470,N_23578,N_22915);
nand UO_1471 (O_1471,N_24795,N_24139);
nand UO_1472 (O_1472,N_23766,N_22790);
or UO_1473 (O_1473,N_23964,N_24676);
nor UO_1474 (O_1474,N_23349,N_22458);
and UO_1475 (O_1475,N_21987,N_23647);
xor UO_1476 (O_1476,N_23017,N_24805);
nand UO_1477 (O_1477,N_24547,N_24893);
nor UO_1478 (O_1478,N_23234,N_22575);
and UO_1479 (O_1479,N_23038,N_23465);
nand UO_1480 (O_1480,N_22669,N_21886);
and UO_1481 (O_1481,N_22860,N_23732);
nor UO_1482 (O_1482,N_22569,N_22209);
or UO_1483 (O_1483,N_24549,N_23934);
nor UO_1484 (O_1484,N_22671,N_22843);
nand UO_1485 (O_1485,N_22560,N_24081);
nor UO_1486 (O_1486,N_24176,N_24451);
and UO_1487 (O_1487,N_21892,N_21902);
nand UO_1488 (O_1488,N_24630,N_24845);
and UO_1489 (O_1489,N_24850,N_23292);
nor UO_1490 (O_1490,N_23612,N_24743);
xor UO_1491 (O_1491,N_22473,N_22182);
or UO_1492 (O_1492,N_24420,N_22617);
or UO_1493 (O_1493,N_23312,N_22567);
nand UO_1494 (O_1494,N_24888,N_23296);
or UO_1495 (O_1495,N_22688,N_23918);
or UO_1496 (O_1496,N_22674,N_22142);
xnor UO_1497 (O_1497,N_24160,N_22389);
and UO_1498 (O_1498,N_22235,N_22957);
nor UO_1499 (O_1499,N_23903,N_24994);
xnor UO_1500 (O_1500,N_23420,N_21883);
nor UO_1501 (O_1501,N_22930,N_24021);
xnor UO_1502 (O_1502,N_24135,N_24720);
nor UO_1503 (O_1503,N_24431,N_24528);
nand UO_1504 (O_1504,N_23978,N_24196);
and UO_1505 (O_1505,N_22249,N_23319);
or UO_1506 (O_1506,N_22489,N_21986);
or UO_1507 (O_1507,N_24771,N_24515);
nor UO_1508 (O_1508,N_22253,N_24691);
or UO_1509 (O_1509,N_22174,N_23073);
xnor UO_1510 (O_1510,N_22080,N_24579);
nor UO_1511 (O_1511,N_23779,N_24033);
or UO_1512 (O_1512,N_23717,N_22194);
nor UO_1513 (O_1513,N_23498,N_22022);
or UO_1514 (O_1514,N_21887,N_21970);
xor UO_1515 (O_1515,N_23240,N_23002);
or UO_1516 (O_1516,N_22269,N_22794);
and UO_1517 (O_1517,N_23355,N_24978);
and UO_1518 (O_1518,N_23310,N_24077);
and UO_1519 (O_1519,N_24248,N_22761);
or UO_1520 (O_1520,N_23447,N_22798);
nand UO_1521 (O_1521,N_23743,N_22692);
or UO_1522 (O_1522,N_23077,N_23293);
nand UO_1523 (O_1523,N_22285,N_23326);
nor UO_1524 (O_1524,N_23615,N_22431);
or UO_1525 (O_1525,N_23041,N_22089);
or UO_1526 (O_1526,N_24849,N_22963);
or UO_1527 (O_1527,N_24442,N_24851);
nand UO_1528 (O_1528,N_24975,N_22382);
nand UO_1529 (O_1529,N_24367,N_23258);
nand UO_1530 (O_1530,N_23621,N_22988);
xor UO_1531 (O_1531,N_24772,N_22465);
nor UO_1532 (O_1532,N_23530,N_22388);
or UO_1533 (O_1533,N_22525,N_23574);
xnor UO_1534 (O_1534,N_22854,N_23120);
or UO_1535 (O_1535,N_23724,N_24198);
nand UO_1536 (O_1536,N_23930,N_22011);
nand UO_1537 (O_1537,N_24463,N_24550);
or UO_1538 (O_1538,N_22281,N_22342);
nor UO_1539 (O_1539,N_24389,N_22634);
nand UO_1540 (O_1540,N_22776,N_22237);
nor UO_1541 (O_1541,N_24346,N_23985);
or UO_1542 (O_1542,N_23850,N_23035);
or UO_1543 (O_1543,N_23346,N_22348);
or UO_1544 (O_1544,N_22757,N_23518);
and UO_1545 (O_1545,N_22001,N_22836);
or UO_1546 (O_1546,N_23366,N_22439);
nand UO_1547 (O_1547,N_24945,N_22725);
xnor UO_1548 (O_1548,N_22149,N_22780);
or UO_1549 (O_1549,N_24214,N_24325);
and UO_1550 (O_1550,N_24379,N_24270);
nor UO_1551 (O_1551,N_24083,N_23640);
or UO_1552 (O_1552,N_22939,N_23379);
or UO_1553 (O_1553,N_23157,N_22372);
nor UO_1554 (O_1554,N_21959,N_23691);
nand UO_1555 (O_1555,N_22610,N_22369);
or UO_1556 (O_1556,N_23807,N_24393);
nand UO_1557 (O_1557,N_22288,N_22030);
or UO_1558 (O_1558,N_22409,N_24401);
nor UO_1559 (O_1559,N_24925,N_23256);
nand UO_1560 (O_1560,N_23500,N_23922);
and UO_1561 (O_1561,N_22004,N_22604);
and UO_1562 (O_1562,N_23730,N_24814);
or UO_1563 (O_1563,N_22463,N_24901);
or UO_1564 (O_1564,N_23166,N_23331);
nor UO_1565 (O_1565,N_23161,N_24689);
or UO_1566 (O_1566,N_24283,N_22735);
nand UO_1567 (O_1567,N_23360,N_24942);
nand UO_1568 (O_1568,N_23469,N_24744);
nor UO_1569 (O_1569,N_23382,N_24621);
and UO_1570 (O_1570,N_24295,N_24703);
nor UO_1571 (O_1571,N_24093,N_22254);
or UO_1572 (O_1572,N_22317,N_23708);
xor UO_1573 (O_1573,N_22569,N_22384);
nor UO_1574 (O_1574,N_22536,N_24468);
and UO_1575 (O_1575,N_23553,N_23473);
xnor UO_1576 (O_1576,N_23608,N_23523);
nand UO_1577 (O_1577,N_23082,N_23125);
nor UO_1578 (O_1578,N_22892,N_23782);
and UO_1579 (O_1579,N_23456,N_24071);
or UO_1580 (O_1580,N_23132,N_22722);
or UO_1581 (O_1581,N_22681,N_24982);
and UO_1582 (O_1582,N_22622,N_22457);
and UO_1583 (O_1583,N_21972,N_24502);
and UO_1584 (O_1584,N_22513,N_23628);
and UO_1585 (O_1585,N_24980,N_22178);
or UO_1586 (O_1586,N_24340,N_22972);
and UO_1587 (O_1587,N_22695,N_24242);
nand UO_1588 (O_1588,N_22485,N_24673);
nor UO_1589 (O_1589,N_22941,N_23262);
nand UO_1590 (O_1590,N_22119,N_24593);
nor UO_1591 (O_1591,N_24126,N_22142);
and UO_1592 (O_1592,N_24552,N_23174);
nand UO_1593 (O_1593,N_22553,N_24050);
nand UO_1594 (O_1594,N_24274,N_22006);
or UO_1595 (O_1595,N_24536,N_22485);
and UO_1596 (O_1596,N_23425,N_23356);
nand UO_1597 (O_1597,N_23954,N_22785);
xnor UO_1598 (O_1598,N_22675,N_24890);
or UO_1599 (O_1599,N_24981,N_23643);
nor UO_1600 (O_1600,N_22349,N_22986);
nand UO_1601 (O_1601,N_22518,N_23428);
and UO_1602 (O_1602,N_22210,N_24872);
and UO_1603 (O_1603,N_24716,N_22930);
or UO_1604 (O_1604,N_24715,N_24919);
nand UO_1605 (O_1605,N_24681,N_24162);
nor UO_1606 (O_1606,N_22468,N_23276);
and UO_1607 (O_1607,N_24926,N_24172);
and UO_1608 (O_1608,N_23841,N_23002);
xor UO_1609 (O_1609,N_22111,N_23992);
and UO_1610 (O_1610,N_22726,N_24422);
nor UO_1611 (O_1611,N_22030,N_23035);
xor UO_1612 (O_1612,N_22331,N_21960);
nand UO_1613 (O_1613,N_24277,N_23071);
nor UO_1614 (O_1614,N_23835,N_24769);
or UO_1615 (O_1615,N_23818,N_21992);
and UO_1616 (O_1616,N_22735,N_22348);
nand UO_1617 (O_1617,N_22552,N_23604);
nor UO_1618 (O_1618,N_22825,N_22654);
and UO_1619 (O_1619,N_24412,N_23626);
nand UO_1620 (O_1620,N_23324,N_24022);
nor UO_1621 (O_1621,N_22690,N_23772);
and UO_1622 (O_1622,N_22008,N_24174);
or UO_1623 (O_1623,N_22044,N_24838);
and UO_1624 (O_1624,N_24621,N_22994);
or UO_1625 (O_1625,N_23936,N_22044);
or UO_1626 (O_1626,N_24940,N_24317);
xnor UO_1627 (O_1627,N_22680,N_24442);
and UO_1628 (O_1628,N_23507,N_22291);
and UO_1629 (O_1629,N_23371,N_23322);
or UO_1630 (O_1630,N_24720,N_23790);
nor UO_1631 (O_1631,N_23404,N_23557);
nor UO_1632 (O_1632,N_24393,N_24933);
nand UO_1633 (O_1633,N_23432,N_22315);
and UO_1634 (O_1634,N_24906,N_21975);
nand UO_1635 (O_1635,N_22543,N_23939);
xor UO_1636 (O_1636,N_23788,N_23856);
and UO_1637 (O_1637,N_23996,N_22363);
nor UO_1638 (O_1638,N_24872,N_22105);
or UO_1639 (O_1639,N_24908,N_23434);
nor UO_1640 (O_1640,N_23832,N_22379);
nor UO_1641 (O_1641,N_23731,N_23276);
nor UO_1642 (O_1642,N_24502,N_24373);
nor UO_1643 (O_1643,N_22654,N_24762);
nor UO_1644 (O_1644,N_24656,N_24740);
or UO_1645 (O_1645,N_23257,N_22708);
and UO_1646 (O_1646,N_24872,N_24345);
xor UO_1647 (O_1647,N_22830,N_22563);
and UO_1648 (O_1648,N_23769,N_24019);
or UO_1649 (O_1649,N_23867,N_24871);
and UO_1650 (O_1650,N_22747,N_22599);
or UO_1651 (O_1651,N_24991,N_24678);
and UO_1652 (O_1652,N_24351,N_22537);
nand UO_1653 (O_1653,N_22191,N_22363);
or UO_1654 (O_1654,N_22920,N_23058);
nand UO_1655 (O_1655,N_22349,N_24723);
nor UO_1656 (O_1656,N_22551,N_22412);
nand UO_1657 (O_1657,N_22496,N_22505);
nand UO_1658 (O_1658,N_22280,N_24215);
nor UO_1659 (O_1659,N_22193,N_22119);
nor UO_1660 (O_1660,N_22014,N_22396);
or UO_1661 (O_1661,N_24431,N_24988);
or UO_1662 (O_1662,N_23819,N_24265);
nor UO_1663 (O_1663,N_23350,N_22270);
nor UO_1664 (O_1664,N_23974,N_22056);
nand UO_1665 (O_1665,N_21982,N_23145);
xnor UO_1666 (O_1666,N_23553,N_23378);
or UO_1667 (O_1667,N_23524,N_24290);
or UO_1668 (O_1668,N_24524,N_23546);
xnor UO_1669 (O_1669,N_22871,N_24497);
or UO_1670 (O_1670,N_24780,N_21876);
or UO_1671 (O_1671,N_22689,N_21933);
nor UO_1672 (O_1672,N_23632,N_24407);
nand UO_1673 (O_1673,N_22511,N_23076);
and UO_1674 (O_1674,N_21966,N_22850);
nand UO_1675 (O_1675,N_22967,N_22417);
nand UO_1676 (O_1676,N_24780,N_23514);
or UO_1677 (O_1677,N_23137,N_24480);
nor UO_1678 (O_1678,N_22816,N_22218);
nor UO_1679 (O_1679,N_23066,N_24403);
or UO_1680 (O_1680,N_23678,N_21959);
or UO_1681 (O_1681,N_22123,N_23372);
or UO_1682 (O_1682,N_23506,N_22169);
nor UO_1683 (O_1683,N_22009,N_22074);
or UO_1684 (O_1684,N_24621,N_23327);
nor UO_1685 (O_1685,N_23313,N_22341);
or UO_1686 (O_1686,N_24672,N_24076);
nor UO_1687 (O_1687,N_22107,N_23221);
and UO_1688 (O_1688,N_23250,N_23400);
nand UO_1689 (O_1689,N_24284,N_22406);
nand UO_1690 (O_1690,N_24505,N_24181);
nor UO_1691 (O_1691,N_23668,N_22994);
or UO_1692 (O_1692,N_23918,N_22013);
and UO_1693 (O_1693,N_24380,N_23847);
xor UO_1694 (O_1694,N_24117,N_24441);
or UO_1695 (O_1695,N_24097,N_24638);
nand UO_1696 (O_1696,N_22915,N_24462);
or UO_1697 (O_1697,N_22036,N_23726);
xnor UO_1698 (O_1698,N_24683,N_22810);
nor UO_1699 (O_1699,N_23819,N_23223);
and UO_1700 (O_1700,N_23523,N_24052);
nor UO_1701 (O_1701,N_23113,N_22767);
or UO_1702 (O_1702,N_24253,N_24789);
and UO_1703 (O_1703,N_22486,N_23051);
and UO_1704 (O_1704,N_24079,N_24796);
and UO_1705 (O_1705,N_22632,N_23802);
nand UO_1706 (O_1706,N_23142,N_24785);
nor UO_1707 (O_1707,N_23766,N_22665);
nand UO_1708 (O_1708,N_23899,N_24164);
and UO_1709 (O_1709,N_23373,N_22117);
and UO_1710 (O_1710,N_22084,N_24861);
nand UO_1711 (O_1711,N_23154,N_24539);
xnor UO_1712 (O_1712,N_22007,N_21971);
nand UO_1713 (O_1713,N_23925,N_23482);
nand UO_1714 (O_1714,N_23640,N_22337);
nand UO_1715 (O_1715,N_22227,N_22211);
nand UO_1716 (O_1716,N_22594,N_24174);
or UO_1717 (O_1717,N_23057,N_23307);
or UO_1718 (O_1718,N_24500,N_22423);
or UO_1719 (O_1719,N_22334,N_22743);
nand UO_1720 (O_1720,N_24311,N_22303);
and UO_1721 (O_1721,N_24826,N_24789);
and UO_1722 (O_1722,N_22558,N_23515);
or UO_1723 (O_1723,N_24505,N_23531);
and UO_1724 (O_1724,N_22228,N_22732);
nand UO_1725 (O_1725,N_22295,N_24616);
nand UO_1726 (O_1726,N_23847,N_22985);
nor UO_1727 (O_1727,N_21933,N_23509);
nor UO_1728 (O_1728,N_22216,N_22325);
nor UO_1729 (O_1729,N_23209,N_23842);
or UO_1730 (O_1730,N_24014,N_24023);
nand UO_1731 (O_1731,N_23059,N_24472);
and UO_1732 (O_1732,N_24090,N_23414);
and UO_1733 (O_1733,N_23734,N_22515);
or UO_1734 (O_1734,N_22785,N_23054);
or UO_1735 (O_1735,N_22739,N_23013);
xor UO_1736 (O_1736,N_22401,N_24415);
and UO_1737 (O_1737,N_24166,N_24005);
or UO_1738 (O_1738,N_22216,N_24466);
nand UO_1739 (O_1739,N_22286,N_23920);
nand UO_1740 (O_1740,N_22629,N_24293);
and UO_1741 (O_1741,N_23619,N_24665);
and UO_1742 (O_1742,N_21906,N_24259);
nand UO_1743 (O_1743,N_22929,N_24804);
or UO_1744 (O_1744,N_24162,N_24748);
or UO_1745 (O_1745,N_24265,N_22782);
or UO_1746 (O_1746,N_21924,N_22712);
and UO_1747 (O_1747,N_23616,N_24791);
nand UO_1748 (O_1748,N_22280,N_24666);
nor UO_1749 (O_1749,N_24180,N_24571);
nand UO_1750 (O_1750,N_23816,N_23657);
nor UO_1751 (O_1751,N_22333,N_23388);
xor UO_1752 (O_1752,N_23156,N_23040);
and UO_1753 (O_1753,N_23549,N_24731);
nand UO_1754 (O_1754,N_23153,N_23240);
nand UO_1755 (O_1755,N_22998,N_23123);
nor UO_1756 (O_1756,N_23662,N_22348);
or UO_1757 (O_1757,N_23624,N_23887);
nor UO_1758 (O_1758,N_22147,N_22699);
nor UO_1759 (O_1759,N_22086,N_24341);
nor UO_1760 (O_1760,N_23023,N_22270);
or UO_1761 (O_1761,N_22056,N_24031);
and UO_1762 (O_1762,N_23035,N_23426);
or UO_1763 (O_1763,N_24896,N_22869);
nand UO_1764 (O_1764,N_22937,N_22103);
nor UO_1765 (O_1765,N_22361,N_23716);
or UO_1766 (O_1766,N_24154,N_23800);
nand UO_1767 (O_1767,N_23795,N_22734);
nand UO_1768 (O_1768,N_24019,N_24451);
xor UO_1769 (O_1769,N_22383,N_24573);
nor UO_1770 (O_1770,N_22174,N_24656);
or UO_1771 (O_1771,N_24548,N_23484);
and UO_1772 (O_1772,N_24940,N_23805);
and UO_1773 (O_1773,N_22011,N_23609);
and UO_1774 (O_1774,N_24909,N_24310);
nor UO_1775 (O_1775,N_22192,N_22142);
or UO_1776 (O_1776,N_23962,N_22979);
nand UO_1777 (O_1777,N_24207,N_23741);
nor UO_1778 (O_1778,N_24321,N_22063);
nor UO_1779 (O_1779,N_23844,N_22436);
or UO_1780 (O_1780,N_24319,N_24456);
nor UO_1781 (O_1781,N_22048,N_23935);
or UO_1782 (O_1782,N_24130,N_23043);
and UO_1783 (O_1783,N_23856,N_22307);
nand UO_1784 (O_1784,N_23885,N_23107);
nand UO_1785 (O_1785,N_22933,N_23107);
xnor UO_1786 (O_1786,N_24345,N_24009);
nand UO_1787 (O_1787,N_24817,N_22297);
nand UO_1788 (O_1788,N_24952,N_23664);
or UO_1789 (O_1789,N_23655,N_23877);
nor UO_1790 (O_1790,N_23846,N_24404);
and UO_1791 (O_1791,N_23552,N_23790);
nand UO_1792 (O_1792,N_23671,N_24607);
or UO_1793 (O_1793,N_24937,N_22514);
or UO_1794 (O_1794,N_24241,N_23990);
xor UO_1795 (O_1795,N_22240,N_24047);
and UO_1796 (O_1796,N_22569,N_24368);
and UO_1797 (O_1797,N_24783,N_22204);
nand UO_1798 (O_1798,N_22821,N_24414);
nand UO_1799 (O_1799,N_23321,N_24314);
or UO_1800 (O_1800,N_22963,N_22766);
or UO_1801 (O_1801,N_22315,N_24600);
nor UO_1802 (O_1802,N_21939,N_24052);
nand UO_1803 (O_1803,N_23360,N_23125);
nand UO_1804 (O_1804,N_23864,N_22953);
or UO_1805 (O_1805,N_22740,N_22719);
or UO_1806 (O_1806,N_23511,N_22085);
nor UO_1807 (O_1807,N_22515,N_24059);
or UO_1808 (O_1808,N_24717,N_24953);
and UO_1809 (O_1809,N_22296,N_24599);
nor UO_1810 (O_1810,N_23522,N_23210);
xor UO_1811 (O_1811,N_24112,N_22347);
xnor UO_1812 (O_1812,N_22465,N_24277);
nor UO_1813 (O_1813,N_21922,N_23847);
xor UO_1814 (O_1814,N_22954,N_24652);
nor UO_1815 (O_1815,N_23499,N_22835);
or UO_1816 (O_1816,N_24357,N_24643);
nand UO_1817 (O_1817,N_23540,N_22990);
nor UO_1818 (O_1818,N_22677,N_23560);
or UO_1819 (O_1819,N_23507,N_24487);
and UO_1820 (O_1820,N_22585,N_24832);
nand UO_1821 (O_1821,N_22837,N_22838);
nand UO_1822 (O_1822,N_22430,N_23609);
nor UO_1823 (O_1823,N_22362,N_23742);
and UO_1824 (O_1824,N_24679,N_22745);
nor UO_1825 (O_1825,N_23395,N_24748);
and UO_1826 (O_1826,N_23195,N_24541);
and UO_1827 (O_1827,N_22565,N_24223);
and UO_1828 (O_1828,N_21950,N_24376);
or UO_1829 (O_1829,N_23923,N_24422);
or UO_1830 (O_1830,N_22614,N_22635);
and UO_1831 (O_1831,N_23349,N_22512);
xnor UO_1832 (O_1832,N_23138,N_24791);
nor UO_1833 (O_1833,N_22476,N_24904);
or UO_1834 (O_1834,N_22167,N_24352);
or UO_1835 (O_1835,N_23373,N_24857);
nor UO_1836 (O_1836,N_23941,N_23902);
or UO_1837 (O_1837,N_22482,N_22298);
or UO_1838 (O_1838,N_22661,N_24021);
nand UO_1839 (O_1839,N_24818,N_24993);
xnor UO_1840 (O_1840,N_23350,N_22932);
nor UO_1841 (O_1841,N_24097,N_24123);
xnor UO_1842 (O_1842,N_23240,N_21921);
nor UO_1843 (O_1843,N_23982,N_23229);
and UO_1844 (O_1844,N_24661,N_22024);
nand UO_1845 (O_1845,N_24123,N_23606);
and UO_1846 (O_1846,N_24312,N_23788);
nand UO_1847 (O_1847,N_22101,N_23732);
nor UO_1848 (O_1848,N_24354,N_22890);
nand UO_1849 (O_1849,N_23913,N_24387);
and UO_1850 (O_1850,N_24886,N_24378);
and UO_1851 (O_1851,N_22914,N_22705);
nand UO_1852 (O_1852,N_22228,N_24192);
xor UO_1853 (O_1853,N_23247,N_22886);
nor UO_1854 (O_1854,N_23906,N_23457);
nand UO_1855 (O_1855,N_23247,N_23900);
xnor UO_1856 (O_1856,N_23711,N_22712);
or UO_1857 (O_1857,N_22260,N_23165);
or UO_1858 (O_1858,N_24825,N_22154);
and UO_1859 (O_1859,N_24417,N_23908);
and UO_1860 (O_1860,N_22531,N_24318);
xor UO_1861 (O_1861,N_22652,N_22496);
nor UO_1862 (O_1862,N_23781,N_24341);
nor UO_1863 (O_1863,N_24207,N_22701);
nand UO_1864 (O_1864,N_23784,N_21940);
xnor UO_1865 (O_1865,N_23820,N_24124);
and UO_1866 (O_1866,N_22051,N_22821);
nor UO_1867 (O_1867,N_24076,N_23351);
and UO_1868 (O_1868,N_21905,N_23582);
nand UO_1869 (O_1869,N_24211,N_24895);
or UO_1870 (O_1870,N_24138,N_22524);
and UO_1871 (O_1871,N_22457,N_22290);
nand UO_1872 (O_1872,N_23135,N_23605);
nand UO_1873 (O_1873,N_24291,N_24756);
nor UO_1874 (O_1874,N_24765,N_23097);
nor UO_1875 (O_1875,N_24724,N_22284);
xnor UO_1876 (O_1876,N_23485,N_22939);
and UO_1877 (O_1877,N_23742,N_22694);
nor UO_1878 (O_1878,N_22244,N_23961);
nor UO_1879 (O_1879,N_23498,N_24842);
xnor UO_1880 (O_1880,N_24766,N_23986);
nand UO_1881 (O_1881,N_22395,N_21886);
nor UO_1882 (O_1882,N_24301,N_22530);
or UO_1883 (O_1883,N_22920,N_23280);
nor UO_1884 (O_1884,N_24590,N_23717);
nand UO_1885 (O_1885,N_23295,N_22266);
or UO_1886 (O_1886,N_23389,N_23398);
or UO_1887 (O_1887,N_23319,N_22448);
and UO_1888 (O_1888,N_24494,N_23294);
nor UO_1889 (O_1889,N_23961,N_24774);
nand UO_1890 (O_1890,N_23043,N_22068);
and UO_1891 (O_1891,N_23663,N_22858);
or UO_1892 (O_1892,N_22981,N_22037);
xor UO_1893 (O_1893,N_21915,N_24486);
xnor UO_1894 (O_1894,N_23930,N_23908);
and UO_1895 (O_1895,N_22980,N_22510);
or UO_1896 (O_1896,N_22828,N_24838);
nand UO_1897 (O_1897,N_22155,N_24114);
and UO_1898 (O_1898,N_22670,N_24880);
nand UO_1899 (O_1899,N_23867,N_24496);
or UO_1900 (O_1900,N_24744,N_24157);
or UO_1901 (O_1901,N_23887,N_22926);
and UO_1902 (O_1902,N_22390,N_22156);
nand UO_1903 (O_1903,N_22901,N_23408);
and UO_1904 (O_1904,N_22035,N_23949);
xor UO_1905 (O_1905,N_23349,N_23417);
nand UO_1906 (O_1906,N_23537,N_22368);
nor UO_1907 (O_1907,N_22068,N_22968);
or UO_1908 (O_1908,N_22211,N_21920);
nand UO_1909 (O_1909,N_24339,N_23830);
nand UO_1910 (O_1910,N_22414,N_22596);
or UO_1911 (O_1911,N_23050,N_24820);
nand UO_1912 (O_1912,N_24313,N_22517);
nor UO_1913 (O_1913,N_22753,N_23718);
or UO_1914 (O_1914,N_24556,N_22147);
nand UO_1915 (O_1915,N_22957,N_23755);
nand UO_1916 (O_1916,N_21921,N_23189);
nor UO_1917 (O_1917,N_24230,N_23596);
or UO_1918 (O_1918,N_23888,N_23314);
nor UO_1919 (O_1919,N_22816,N_24883);
and UO_1920 (O_1920,N_22857,N_22470);
nor UO_1921 (O_1921,N_24248,N_22973);
or UO_1922 (O_1922,N_23948,N_23512);
or UO_1923 (O_1923,N_22226,N_23668);
nand UO_1924 (O_1924,N_22364,N_23330);
nand UO_1925 (O_1925,N_22475,N_22506);
nor UO_1926 (O_1926,N_23266,N_24411);
nand UO_1927 (O_1927,N_22204,N_23188);
or UO_1928 (O_1928,N_22210,N_23774);
xor UO_1929 (O_1929,N_24319,N_21897);
and UO_1930 (O_1930,N_23772,N_22516);
or UO_1931 (O_1931,N_23672,N_23403);
and UO_1932 (O_1932,N_22727,N_23367);
nand UO_1933 (O_1933,N_24322,N_22235);
nor UO_1934 (O_1934,N_23386,N_24982);
nand UO_1935 (O_1935,N_24722,N_22428);
nor UO_1936 (O_1936,N_24908,N_24712);
and UO_1937 (O_1937,N_24230,N_23246);
or UO_1938 (O_1938,N_24515,N_22318);
and UO_1939 (O_1939,N_22454,N_24740);
nor UO_1940 (O_1940,N_23129,N_24689);
or UO_1941 (O_1941,N_23359,N_21981);
nand UO_1942 (O_1942,N_22928,N_24387);
nand UO_1943 (O_1943,N_24273,N_22868);
nor UO_1944 (O_1944,N_24692,N_24959);
or UO_1945 (O_1945,N_24049,N_23898);
nand UO_1946 (O_1946,N_24393,N_24545);
or UO_1947 (O_1947,N_23336,N_24347);
nand UO_1948 (O_1948,N_23645,N_22982);
and UO_1949 (O_1949,N_21979,N_23048);
or UO_1950 (O_1950,N_23325,N_22951);
nor UO_1951 (O_1951,N_24778,N_23725);
or UO_1952 (O_1952,N_23473,N_22347);
or UO_1953 (O_1953,N_22841,N_23180);
nand UO_1954 (O_1954,N_24606,N_23122);
nand UO_1955 (O_1955,N_23507,N_24185);
or UO_1956 (O_1956,N_22144,N_22045);
xor UO_1957 (O_1957,N_24168,N_23297);
or UO_1958 (O_1958,N_22520,N_22264);
and UO_1959 (O_1959,N_24288,N_22392);
and UO_1960 (O_1960,N_24313,N_22126);
nor UO_1961 (O_1961,N_23754,N_22861);
nand UO_1962 (O_1962,N_24170,N_24851);
and UO_1963 (O_1963,N_24479,N_21935);
nor UO_1964 (O_1964,N_22566,N_21979);
and UO_1965 (O_1965,N_22601,N_23946);
and UO_1966 (O_1966,N_24199,N_24360);
nand UO_1967 (O_1967,N_23009,N_23897);
nand UO_1968 (O_1968,N_23373,N_24884);
xnor UO_1969 (O_1969,N_23934,N_22873);
and UO_1970 (O_1970,N_22620,N_23720);
and UO_1971 (O_1971,N_23542,N_21944);
nand UO_1972 (O_1972,N_23293,N_23042);
and UO_1973 (O_1973,N_23779,N_23204);
or UO_1974 (O_1974,N_24539,N_23000);
or UO_1975 (O_1975,N_23014,N_24309);
nand UO_1976 (O_1976,N_22553,N_22790);
nor UO_1977 (O_1977,N_24322,N_22686);
nor UO_1978 (O_1978,N_24892,N_22532);
nor UO_1979 (O_1979,N_22845,N_23716);
nor UO_1980 (O_1980,N_24961,N_24824);
xor UO_1981 (O_1981,N_23425,N_22392);
nor UO_1982 (O_1982,N_24242,N_23093);
nor UO_1983 (O_1983,N_22859,N_23904);
nor UO_1984 (O_1984,N_24029,N_22821);
nand UO_1985 (O_1985,N_22241,N_23730);
nand UO_1986 (O_1986,N_22695,N_23422);
or UO_1987 (O_1987,N_22110,N_22659);
or UO_1988 (O_1988,N_23690,N_23208);
or UO_1989 (O_1989,N_22831,N_23517);
and UO_1990 (O_1990,N_24052,N_22103);
and UO_1991 (O_1991,N_24728,N_24514);
or UO_1992 (O_1992,N_24097,N_22901);
nand UO_1993 (O_1993,N_22500,N_22701);
and UO_1994 (O_1994,N_22480,N_23016);
and UO_1995 (O_1995,N_24771,N_23881);
and UO_1996 (O_1996,N_22282,N_23741);
nand UO_1997 (O_1997,N_24214,N_22531);
nand UO_1998 (O_1998,N_21966,N_22918);
and UO_1999 (O_1999,N_22521,N_24115);
and UO_2000 (O_2000,N_23033,N_23067);
nor UO_2001 (O_2001,N_23137,N_24489);
nor UO_2002 (O_2002,N_24647,N_24478);
and UO_2003 (O_2003,N_22321,N_22870);
nand UO_2004 (O_2004,N_23315,N_22450);
and UO_2005 (O_2005,N_22020,N_23420);
nor UO_2006 (O_2006,N_22967,N_22605);
and UO_2007 (O_2007,N_23142,N_23959);
or UO_2008 (O_2008,N_22063,N_23490);
nor UO_2009 (O_2009,N_23202,N_23920);
or UO_2010 (O_2010,N_22364,N_24849);
nand UO_2011 (O_2011,N_23808,N_24149);
or UO_2012 (O_2012,N_24270,N_24723);
and UO_2013 (O_2013,N_22537,N_23481);
nor UO_2014 (O_2014,N_22763,N_24477);
or UO_2015 (O_2015,N_24441,N_23344);
and UO_2016 (O_2016,N_24468,N_24625);
nand UO_2017 (O_2017,N_24213,N_22030);
nor UO_2018 (O_2018,N_23935,N_24824);
or UO_2019 (O_2019,N_23632,N_24747);
or UO_2020 (O_2020,N_23841,N_22208);
and UO_2021 (O_2021,N_23207,N_24321);
or UO_2022 (O_2022,N_24537,N_24143);
nor UO_2023 (O_2023,N_23214,N_22951);
or UO_2024 (O_2024,N_24757,N_24295);
and UO_2025 (O_2025,N_22678,N_23072);
and UO_2026 (O_2026,N_22888,N_24984);
nand UO_2027 (O_2027,N_22613,N_23575);
or UO_2028 (O_2028,N_22708,N_22921);
and UO_2029 (O_2029,N_23968,N_22069);
nor UO_2030 (O_2030,N_22707,N_22818);
nor UO_2031 (O_2031,N_23143,N_22134);
and UO_2032 (O_2032,N_23139,N_24383);
nand UO_2033 (O_2033,N_23325,N_24948);
and UO_2034 (O_2034,N_22420,N_21896);
and UO_2035 (O_2035,N_23431,N_24920);
xnor UO_2036 (O_2036,N_23947,N_22336);
or UO_2037 (O_2037,N_24225,N_24303);
nor UO_2038 (O_2038,N_22510,N_22837);
and UO_2039 (O_2039,N_23409,N_24269);
or UO_2040 (O_2040,N_23561,N_23927);
and UO_2041 (O_2041,N_24439,N_22418);
nand UO_2042 (O_2042,N_24768,N_23948);
and UO_2043 (O_2043,N_21904,N_24804);
nor UO_2044 (O_2044,N_24475,N_22947);
nor UO_2045 (O_2045,N_24886,N_23081);
and UO_2046 (O_2046,N_22527,N_23605);
nand UO_2047 (O_2047,N_23769,N_24848);
xnor UO_2048 (O_2048,N_23697,N_22588);
or UO_2049 (O_2049,N_24527,N_23018);
nor UO_2050 (O_2050,N_22839,N_24333);
and UO_2051 (O_2051,N_22268,N_23716);
or UO_2052 (O_2052,N_24691,N_24906);
or UO_2053 (O_2053,N_22644,N_22132);
or UO_2054 (O_2054,N_22760,N_24266);
nand UO_2055 (O_2055,N_24892,N_23368);
and UO_2056 (O_2056,N_23326,N_24012);
and UO_2057 (O_2057,N_22543,N_24298);
or UO_2058 (O_2058,N_23202,N_22316);
or UO_2059 (O_2059,N_24426,N_24449);
or UO_2060 (O_2060,N_24845,N_22889);
and UO_2061 (O_2061,N_23415,N_22435);
nand UO_2062 (O_2062,N_24225,N_23470);
and UO_2063 (O_2063,N_24289,N_23396);
or UO_2064 (O_2064,N_24231,N_23527);
nand UO_2065 (O_2065,N_24727,N_23896);
xor UO_2066 (O_2066,N_22762,N_23204);
and UO_2067 (O_2067,N_22978,N_24958);
nor UO_2068 (O_2068,N_24181,N_24964);
xor UO_2069 (O_2069,N_23547,N_24062);
nor UO_2070 (O_2070,N_22673,N_23639);
nor UO_2071 (O_2071,N_24975,N_22453);
and UO_2072 (O_2072,N_22708,N_24447);
nor UO_2073 (O_2073,N_22142,N_22437);
nand UO_2074 (O_2074,N_22921,N_22217);
and UO_2075 (O_2075,N_23684,N_21936);
and UO_2076 (O_2076,N_22312,N_21918);
and UO_2077 (O_2077,N_23822,N_23296);
and UO_2078 (O_2078,N_23780,N_22660);
nor UO_2079 (O_2079,N_23308,N_22976);
or UO_2080 (O_2080,N_24587,N_23786);
nor UO_2081 (O_2081,N_24229,N_24053);
and UO_2082 (O_2082,N_22296,N_22001);
and UO_2083 (O_2083,N_22968,N_24414);
and UO_2084 (O_2084,N_22965,N_23610);
and UO_2085 (O_2085,N_24227,N_23568);
nand UO_2086 (O_2086,N_24168,N_24976);
xor UO_2087 (O_2087,N_23340,N_22536);
nand UO_2088 (O_2088,N_23120,N_22478);
and UO_2089 (O_2089,N_22902,N_21962);
xor UO_2090 (O_2090,N_22859,N_22121);
nor UO_2091 (O_2091,N_23579,N_23694);
and UO_2092 (O_2092,N_23041,N_24766);
nor UO_2093 (O_2093,N_21964,N_23544);
and UO_2094 (O_2094,N_22060,N_24084);
xnor UO_2095 (O_2095,N_22781,N_24204);
nor UO_2096 (O_2096,N_22566,N_22397);
nor UO_2097 (O_2097,N_23305,N_24032);
nand UO_2098 (O_2098,N_22862,N_23301);
nand UO_2099 (O_2099,N_22541,N_22236);
nor UO_2100 (O_2100,N_22630,N_23533);
nor UO_2101 (O_2101,N_24960,N_24473);
or UO_2102 (O_2102,N_24410,N_23141);
and UO_2103 (O_2103,N_23664,N_24147);
nand UO_2104 (O_2104,N_22159,N_24137);
or UO_2105 (O_2105,N_23827,N_22281);
nand UO_2106 (O_2106,N_24686,N_24627);
and UO_2107 (O_2107,N_22964,N_22102);
nand UO_2108 (O_2108,N_22910,N_23490);
nand UO_2109 (O_2109,N_22479,N_24343);
and UO_2110 (O_2110,N_24382,N_23110);
and UO_2111 (O_2111,N_22502,N_23368);
or UO_2112 (O_2112,N_23326,N_22473);
nor UO_2113 (O_2113,N_22999,N_24775);
nor UO_2114 (O_2114,N_23615,N_23372);
nand UO_2115 (O_2115,N_23992,N_22509);
nand UO_2116 (O_2116,N_22452,N_23360);
nand UO_2117 (O_2117,N_22827,N_22344);
and UO_2118 (O_2118,N_24125,N_23539);
and UO_2119 (O_2119,N_23960,N_23389);
nor UO_2120 (O_2120,N_24614,N_23289);
xnor UO_2121 (O_2121,N_23415,N_24677);
nor UO_2122 (O_2122,N_22083,N_24637);
or UO_2123 (O_2123,N_23551,N_22026);
or UO_2124 (O_2124,N_24972,N_24795);
xor UO_2125 (O_2125,N_22574,N_22471);
nor UO_2126 (O_2126,N_24621,N_22405);
and UO_2127 (O_2127,N_24535,N_23770);
xor UO_2128 (O_2128,N_22011,N_24549);
or UO_2129 (O_2129,N_24784,N_22580);
nand UO_2130 (O_2130,N_23240,N_23231);
or UO_2131 (O_2131,N_24032,N_23660);
and UO_2132 (O_2132,N_24050,N_24748);
and UO_2133 (O_2133,N_23827,N_24911);
xnor UO_2134 (O_2134,N_24713,N_23522);
nand UO_2135 (O_2135,N_22284,N_23763);
or UO_2136 (O_2136,N_24632,N_22832);
nor UO_2137 (O_2137,N_22392,N_21953);
or UO_2138 (O_2138,N_24665,N_22687);
or UO_2139 (O_2139,N_21945,N_24379);
nor UO_2140 (O_2140,N_22875,N_24661);
and UO_2141 (O_2141,N_24362,N_22126);
xnor UO_2142 (O_2142,N_23053,N_22775);
nor UO_2143 (O_2143,N_24220,N_22320);
and UO_2144 (O_2144,N_23950,N_23040);
and UO_2145 (O_2145,N_22815,N_23991);
and UO_2146 (O_2146,N_22246,N_23560);
and UO_2147 (O_2147,N_22773,N_22549);
or UO_2148 (O_2148,N_22017,N_23578);
and UO_2149 (O_2149,N_23532,N_22866);
nand UO_2150 (O_2150,N_22742,N_24130);
nor UO_2151 (O_2151,N_23344,N_21915);
and UO_2152 (O_2152,N_24018,N_24817);
or UO_2153 (O_2153,N_24273,N_23958);
nand UO_2154 (O_2154,N_24558,N_22474);
nand UO_2155 (O_2155,N_22074,N_22952);
and UO_2156 (O_2156,N_22200,N_22664);
or UO_2157 (O_2157,N_24136,N_24799);
or UO_2158 (O_2158,N_22375,N_22447);
or UO_2159 (O_2159,N_23425,N_24252);
or UO_2160 (O_2160,N_22349,N_22822);
and UO_2161 (O_2161,N_22101,N_23229);
nand UO_2162 (O_2162,N_24591,N_24543);
nand UO_2163 (O_2163,N_23365,N_22519);
and UO_2164 (O_2164,N_23464,N_23295);
nor UO_2165 (O_2165,N_21925,N_24303);
nand UO_2166 (O_2166,N_22265,N_24351);
nor UO_2167 (O_2167,N_22365,N_24346);
nand UO_2168 (O_2168,N_23631,N_23245);
nor UO_2169 (O_2169,N_23109,N_22646);
and UO_2170 (O_2170,N_23075,N_22192);
and UO_2171 (O_2171,N_24864,N_24547);
nor UO_2172 (O_2172,N_23134,N_24596);
nand UO_2173 (O_2173,N_23645,N_23615);
or UO_2174 (O_2174,N_22609,N_23697);
or UO_2175 (O_2175,N_23072,N_22835);
and UO_2176 (O_2176,N_22748,N_24134);
and UO_2177 (O_2177,N_22647,N_22969);
nand UO_2178 (O_2178,N_24979,N_24414);
nand UO_2179 (O_2179,N_23830,N_24175);
or UO_2180 (O_2180,N_21933,N_22064);
nor UO_2181 (O_2181,N_21940,N_22744);
and UO_2182 (O_2182,N_23804,N_24873);
and UO_2183 (O_2183,N_22217,N_24186);
or UO_2184 (O_2184,N_23177,N_24737);
or UO_2185 (O_2185,N_24427,N_24989);
nand UO_2186 (O_2186,N_22843,N_23389);
nor UO_2187 (O_2187,N_24679,N_22420);
xnor UO_2188 (O_2188,N_24903,N_24917);
nand UO_2189 (O_2189,N_22826,N_23239);
nor UO_2190 (O_2190,N_22229,N_23268);
or UO_2191 (O_2191,N_23005,N_22230);
nand UO_2192 (O_2192,N_22016,N_24322);
or UO_2193 (O_2193,N_21921,N_22990);
xor UO_2194 (O_2194,N_24821,N_21881);
or UO_2195 (O_2195,N_22198,N_24223);
and UO_2196 (O_2196,N_22303,N_23167);
and UO_2197 (O_2197,N_23438,N_22527);
nor UO_2198 (O_2198,N_23695,N_23048);
nor UO_2199 (O_2199,N_24957,N_24915);
or UO_2200 (O_2200,N_24238,N_24263);
and UO_2201 (O_2201,N_22959,N_22552);
nand UO_2202 (O_2202,N_24591,N_23472);
and UO_2203 (O_2203,N_22922,N_22484);
xor UO_2204 (O_2204,N_22253,N_23226);
nand UO_2205 (O_2205,N_22945,N_22583);
nor UO_2206 (O_2206,N_22151,N_22736);
nand UO_2207 (O_2207,N_23307,N_22656);
nor UO_2208 (O_2208,N_23864,N_23273);
nor UO_2209 (O_2209,N_24736,N_24060);
or UO_2210 (O_2210,N_22906,N_22660);
and UO_2211 (O_2211,N_22935,N_24876);
nor UO_2212 (O_2212,N_22437,N_22294);
nand UO_2213 (O_2213,N_22177,N_24904);
or UO_2214 (O_2214,N_23698,N_24875);
and UO_2215 (O_2215,N_22573,N_23965);
xor UO_2216 (O_2216,N_22259,N_22192);
or UO_2217 (O_2217,N_23823,N_21912);
or UO_2218 (O_2218,N_23735,N_24869);
xor UO_2219 (O_2219,N_23470,N_23924);
or UO_2220 (O_2220,N_22121,N_22080);
and UO_2221 (O_2221,N_21957,N_24163);
nor UO_2222 (O_2222,N_24497,N_22919);
or UO_2223 (O_2223,N_22200,N_24713);
nor UO_2224 (O_2224,N_23333,N_23892);
xnor UO_2225 (O_2225,N_24191,N_24375);
and UO_2226 (O_2226,N_23914,N_22192);
and UO_2227 (O_2227,N_22989,N_23982);
nand UO_2228 (O_2228,N_24157,N_23741);
or UO_2229 (O_2229,N_23750,N_23715);
and UO_2230 (O_2230,N_24506,N_23122);
nand UO_2231 (O_2231,N_24411,N_22787);
xor UO_2232 (O_2232,N_22646,N_24084);
or UO_2233 (O_2233,N_24430,N_23434);
and UO_2234 (O_2234,N_22683,N_23915);
and UO_2235 (O_2235,N_24413,N_21904);
nor UO_2236 (O_2236,N_22466,N_22786);
and UO_2237 (O_2237,N_24205,N_23570);
or UO_2238 (O_2238,N_23612,N_24247);
or UO_2239 (O_2239,N_24657,N_24292);
nor UO_2240 (O_2240,N_23563,N_23235);
nand UO_2241 (O_2241,N_24978,N_22123);
or UO_2242 (O_2242,N_24897,N_24056);
nand UO_2243 (O_2243,N_24329,N_23924);
or UO_2244 (O_2244,N_21998,N_24285);
nor UO_2245 (O_2245,N_24095,N_23902);
nor UO_2246 (O_2246,N_22692,N_24078);
nand UO_2247 (O_2247,N_22949,N_22262);
and UO_2248 (O_2248,N_24076,N_22641);
or UO_2249 (O_2249,N_24128,N_23490);
nand UO_2250 (O_2250,N_22336,N_24979);
nor UO_2251 (O_2251,N_24166,N_24083);
nand UO_2252 (O_2252,N_23907,N_22822);
xor UO_2253 (O_2253,N_24839,N_24713);
or UO_2254 (O_2254,N_22259,N_23061);
nand UO_2255 (O_2255,N_23798,N_23261);
nand UO_2256 (O_2256,N_22399,N_24277);
and UO_2257 (O_2257,N_24332,N_22305);
nand UO_2258 (O_2258,N_24051,N_23988);
nor UO_2259 (O_2259,N_22246,N_24337);
or UO_2260 (O_2260,N_24531,N_23100);
or UO_2261 (O_2261,N_22926,N_22276);
nor UO_2262 (O_2262,N_23308,N_22050);
nand UO_2263 (O_2263,N_23817,N_22612);
or UO_2264 (O_2264,N_23034,N_24258);
nand UO_2265 (O_2265,N_24103,N_23758);
and UO_2266 (O_2266,N_24022,N_22956);
and UO_2267 (O_2267,N_23557,N_21898);
or UO_2268 (O_2268,N_23729,N_22178);
or UO_2269 (O_2269,N_22071,N_22494);
nor UO_2270 (O_2270,N_23257,N_22105);
nor UO_2271 (O_2271,N_23755,N_22106);
nand UO_2272 (O_2272,N_23738,N_22617);
nor UO_2273 (O_2273,N_23798,N_22829);
nor UO_2274 (O_2274,N_23865,N_23196);
xor UO_2275 (O_2275,N_23046,N_23779);
nand UO_2276 (O_2276,N_24323,N_23166);
xor UO_2277 (O_2277,N_23007,N_21925);
nor UO_2278 (O_2278,N_23815,N_23250);
and UO_2279 (O_2279,N_24927,N_24233);
and UO_2280 (O_2280,N_24116,N_23912);
xnor UO_2281 (O_2281,N_24324,N_23071);
nand UO_2282 (O_2282,N_23919,N_22175);
nand UO_2283 (O_2283,N_22850,N_24083);
or UO_2284 (O_2284,N_22617,N_24190);
or UO_2285 (O_2285,N_22992,N_23001);
xor UO_2286 (O_2286,N_24794,N_24973);
or UO_2287 (O_2287,N_24212,N_23879);
and UO_2288 (O_2288,N_24007,N_23457);
nor UO_2289 (O_2289,N_24882,N_24684);
nand UO_2290 (O_2290,N_23615,N_24839);
or UO_2291 (O_2291,N_23550,N_24457);
xnor UO_2292 (O_2292,N_21917,N_24675);
or UO_2293 (O_2293,N_22788,N_22023);
nor UO_2294 (O_2294,N_23218,N_24774);
nand UO_2295 (O_2295,N_24403,N_24830);
nand UO_2296 (O_2296,N_22344,N_24193);
nor UO_2297 (O_2297,N_22917,N_24061);
or UO_2298 (O_2298,N_23236,N_22494);
nor UO_2299 (O_2299,N_24515,N_24210);
nor UO_2300 (O_2300,N_24336,N_22981);
or UO_2301 (O_2301,N_23538,N_22290);
nand UO_2302 (O_2302,N_23182,N_23136);
nor UO_2303 (O_2303,N_22054,N_24497);
and UO_2304 (O_2304,N_23931,N_22519);
or UO_2305 (O_2305,N_24945,N_24737);
or UO_2306 (O_2306,N_22218,N_22425);
or UO_2307 (O_2307,N_23988,N_24824);
nand UO_2308 (O_2308,N_21959,N_24978);
and UO_2309 (O_2309,N_23938,N_23285);
and UO_2310 (O_2310,N_24747,N_24046);
nor UO_2311 (O_2311,N_23958,N_22333);
xor UO_2312 (O_2312,N_23809,N_22860);
nor UO_2313 (O_2313,N_22798,N_22409);
nor UO_2314 (O_2314,N_23989,N_23625);
xnor UO_2315 (O_2315,N_24214,N_23288);
xor UO_2316 (O_2316,N_24707,N_23172);
and UO_2317 (O_2317,N_23682,N_22318);
nor UO_2318 (O_2318,N_22529,N_24418);
and UO_2319 (O_2319,N_21916,N_24549);
nand UO_2320 (O_2320,N_22672,N_24812);
nor UO_2321 (O_2321,N_24825,N_22436);
or UO_2322 (O_2322,N_24083,N_22420);
and UO_2323 (O_2323,N_23028,N_21897);
xor UO_2324 (O_2324,N_22386,N_23544);
nand UO_2325 (O_2325,N_23645,N_22847);
nand UO_2326 (O_2326,N_24238,N_24622);
and UO_2327 (O_2327,N_23514,N_22137);
nor UO_2328 (O_2328,N_24773,N_23960);
nor UO_2329 (O_2329,N_23044,N_22645);
or UO_2330 (O_2330,N_22705,N_21879);
nand UO_2331 (O_2331,N_22899,N_24988);
xor UO_2332 (O_2332,N_22482,N_23751);
nor UO_2333 (O_2333,N_23850,N_22544);
xor UO_2334 (O_2334,N_24656,N_23607);
nor UO_2335 (O_2335,N_24316,N_23521);
and UO_2336 (O_2336,N_22019,N_22890);
xor UO_2337 (O_2337,N_24559,N_23406);
nand UO_2338 (O_2338,N_24318,N_22681);
nor UO_2339 (O_2339,N_23885,N_24185);
and UO_2340 (O_2340,N_24048,N_23794);
nor UO_2341 (O_2341,N_22989,N_24334);
nor UO_2342 (O_2342,N_24789,N_23022);
or UO_2343 (O_2343,N_23844,N_23028);
nor UO_2344 (O_2344,N_22681,N_23320);
nand UO_2345 (O_2345,N_24500,N_23108);
nand UO_2346 (O_2346,N_23017,N_22648);
and UO_2347 (O_2347,N_23462,N_23837);
nand UO_2348 (O_2348,N_23120,N_24138);
or UO_2349 (O_2349,N_24358,N_23020);
nor UO_2350 (O_2350,N_24520,N_23678);
xnor UO_2351 (O_2351,N_24034,N_24023);
or UO_2352 (O_2352,N_23974,N_24973);
xnor UO_2353 (O_2353,N_22746,N_22034);
nand UO_2354 (O_2354,N_22033,N_24816);
or UO_2355 (O_2355,N_24456,N_24704);
or UO_2356 (O_2356,N_22518,N_22015);
and UO_2357 (O_2357,N_21958,N_23173);
nand UO_2358 (O_2358,N_21914,N_23308);
or UO_2359 (O_2359,N_23269,N_24250);
and UO_2360 (O_2360,N_24780,N_24870);
and UO_2361 (O_2361,N_24279,N_24432);
nor UO_2362 (O_2362,N_22075,N_24495);
and UO_2363 (O_2363,N_24048,N_23379);
nor UO_2364 (O_2364,N_21922,N_22281);
nor UO_2365 (O_2365,N_23417,N_23765);
nor UO_2366 (O_2366,N_22048,N_23175);
and UO_2367 (O_2367,N_22005,N_21970);
nor UO_2368 (O_2368,N_24815,N_23911);
xnor UO_2369 (O_2369,N_22167,N_24372);
nor UO_2370 (O_2370,N_22271,N_22308);
nor UO_2371 (O_2371,N_22202,N_23740);
nor UO_2372 (O_2372,N_22335,N_24189);
or UO_2373 (O_2373,N_23277,N_24933);
xnor UO_2374 (O_2374,N_23993,N_23577);
nand UO_2375 (O_2375,N_23142,N_23270);
or UO_2376 (O_2376,N_22148,N_23762);
nand UO_2377 (O_2377,N_22820,N_22123);
or UO_2378 (O_2378,N_23237,N_22105);
xor UO_2379 (O_2379,N_23597,N_22031);
or UO_2380 (O_2380,N_23920,N_23500);
or UO_2381 (O_2381,N_22234,N_23146);
or UO_2382 (O_2382,N_23170,N_24236);
nand UO_2383 (O_2383,N_22843,N_22801);
or UO_2384 (O_2384,N_23788,N_23451);
or UO_2385 (O_2385,N_23124,N_24949);
or UO_2386 (O_2386,N_23612,N_24577);
or UO_2387 (O_2387,N_24289,N_23540);
or UO_2388 (O_2388,N_21902,N_23810);
or UO_2389 (O_2389,N_23362,N_22979);
and UO_2390 (O_2390,N_24723,N_22967);
nor UO_2391 (O_2391,N_23531,N_23277);
nand UO_2392 (O_2392,N_24713,N_22875);
or UO_2393 (O_2393,N_23442,N_22325);
nand UO_2394 (O_2394,N_22909,N_24914);
xnor UO_2395 (O_2395,N_23867,N_22725);
nor UO_2396 (O_2396,N_23450,N_24255);
or UO_2397 (O_2397,N_21956,N_23664);
nor UO_2398 (O_2398,N_23890,N_24056);
xor UO_2399 (O_2399,N_24635,N_24557);
xor UO_2400 (O_2400,N_23227,N_22241);
nand UO_2401 (O_2401,N_22956,N_24420);
nor UO_2402 (O_2402,N_23866,N_23689);
nor UO_2403 (O_2403,N_22885,N_22575);
and UO_2404 (O_2404,N_23012,N_21901);
xor UO_2405 (O_2405,N_22909,N_24572);
nand UO_2406 (O_2406,N_23484,N_22087);
nor UO_2407 (O_2407,N_22198,N_23535);
xnor UO_2408 (O_2408,N_24024,N_24159);
or UO_2409 (O_2409,N_23488,N_24695);
nand UO_2410 (O_2410,N_23889,N_24519);
nor UO_2411 (O_2411,N_23699,N_22716);
or UO_2412 (O_2412,N_22051,N_24475);
and UO_2413 (O_2413,N_23006,N_22166);
nand UO_2414 (O_2414,N_24820,N_22585);
or UO_2415 (O_2415,N_23768,N_24651);
nor UO_2416 (O_2416,N_22025,N_23724);
and UO_2417 (O_2417,N_24664,N_23613);
or UO_2418 (O_2418,N_23695,N_23435);
and UO_2419 (O_2419,N_24377,N_23909);
nand UO_2420 (O_2420,N_24958,N_24141);
xor UO_2421 (O_2421,N_22071,N_24294);
and UO_2422 (O_2422,N_22847,N_23331);
nand UO_2423 (O_2423,N_22177,N_23502);
and UO_2424 (O_2424,N_22423,N_22041);
nand UO_2425 (O_2425,N_22572,N_22036);
or UO_2426 (O_2426,N_24330,N_22948);
nor UO_2427 (O_2427,N_23389,N_23743);
and UO_2428 (O_2428,N_23456,N_24121);
and UO_2429 (O_2429,N_23078,N_23697);
xnor UO_2430 (O_2430,N_24708,N_23436);
or UO_2431 (O_2431,N_24833,N_22612);
and UO_2432 (O_2432,N_23660,N_23976);
and UO_2433 (O_2433,N_24539,N_21888);
and UO_2434 (O_2434,N_24554,N_23878);
or UO_2435 (O_2435,N_23317,N_23151);
nor UO_2436 (O_2436,N_23177,N_23203);
nand UO_2437 (O_2437,N_23077,N_23764);
nor UO_2438 (O_2438,N_24884,N_24485);
and UO_2439 (O_2439,N_22577,N_23905);
and UO_2440 (O_2440,N_24872,N_22431);
nand UO_2441 (O_2441,N_24095,N_22316);
nand UO_2442 (O_2442,N_24201,N_22253);
and UO_2443 (O_2443,N_21947,N_23997);
or UO_2444 (O_2444,N_24954,N_22759);
and UO_2445 (O_2445,N_22331,N_24605);
nand UO_2446 (O_2446,N_23281,N_23645);
nand UO_2447 (O_2447,N_24543,N_24111);
nand UO_2448 (O_2448,N_24584,N_21989);
or UO_2449 (O_2449,N_24878,N_21998);
nor UO_2450 (O_2450,N_23092,N_24794);
or UO_2451 (O_2451,N_24621,N_22240);
and UO_2452 (O_2452,N_21964,N_23402);
nor UO_2453 (O_2453,N_24844,N_24428);
or UO_2454 (O_2454,N_24830,N_23217);
nand UO_2455 (O_2455,N_22034,N_23320);
nand UO_2456 (O_2456,N_23001,N_22112);
or UO_2457 (O_2457,N_24122,N_22709);
nor UO_2458 (O_2458,N_21980,N_24569);
nor UO_2459 (O_2459,N_22551,N_21947);
nand UO_2460 (O_2460,N_24410,N_22425);
nor UO_2461 (O_2461,N_22526,N_22042);
nor UO_2462 (O_2462,N_22523,N_22644);
or UO_2463 (O_2463,N_23985,N_23748);
xnor UO_2464 (O_2464,N_23386,N_23454);
nand UO_2465 (O_2465,N_23407,N_23030);
or UO_2466 (O_2466,N_24244,N_23735);
or UO_2467 (O_2467,N_24755,N_23215);
nand UO_2468 (O_2468,N_24764,N_21883);
nor UO_2469 (O_2469,N_22935,N_22521);
and UO_2470 (O_2470,N_24013,N_21932);
nor UO_2471 (O_2471,N_22651,N_23063);
nand UO_2472 (O_2472,N_24987,N_23702);
nor UO_2473 (O_2473,N_23072,N_22154);
nor UO_2474 (O_2474,N_22955,N_23605);
nor UO_2475 (O_2475,N_23760,N_24847);
xor UO_2476 (O_2476,N_22618,N_24041);
and UO_2477 (O_2477,N_22610,N_22043);
and UO_2478 (O_2478,N_23974,N_23345);
nand UO_2479 (O_2479,N_23127,N_23561);
nand UO_2480 (O_2480,N_21969,N_24326);
and UO_2481 (O_2481,N_23214,N_22436);
or UO_2482 (O_2482,N_22382,N_24255);
xnor UO_2483 (O_2483,N_24978,N_23320);
and UO_2484 (O_2484,N_23688,N_23706);
nand UO_2485 (O_2485,N_23022,N_21893);
nor UO_2486 (O_2486,N_21928,N_23334);
or UO_2487 (O_2487,N_24362,N_22180);
nand UO_2488 (O_2488,N_23726,N_22025);
xnor UO_2489 (O_2489,N_24934,N_22368);
nand UO_2490 (O_2490,N_24415,N_24262);
and UO_2491 (O_2491,N_22751,N_24219);
xnor UO_2492 (O_2492,N_22352,N_23974);
nand UO_2493 (O_2493,N_22540,N_24041);
nand UO_2494 (O_2494,N_21888,N_22833);
nand UO_2495 (O_2495,N_23867,N_24926);
nor UO_2496 (O_2496,N_22861,N_22840);
or UO_2497 (O_2497,N_23543,N_22603);
xnor UO_2498 (O_2498,N_23540,N_24512);
and UO_2499 (O_2499,N_22198,N_22281);
or UO_2500 (O_2500,N_24938,N_23736);
or UO_2501 (O_2501,N_23971,N_23067);
or UO_2502 (O_2502,N_22075,N_22801);
nand UO_2503 (O_2503,N_24401,N_22037);
xor UO_2504 (O_2504,N_24193,N_23947);
nand UO_2505 (O_2505,N_22775,N_23301);
nor UO_2506 (O_2506,N_24733,N_22272);
nor UO_2507 (O_2507,N_24774,N_23660);
nor UO_2508 (O_2508,N_24628,N_23239);
xnor UO_2509 (O_2509,N_23810,N_23126);
nor UO_2510 (O_2510,N_23116,N_24863);
nand UO_2511 (O_2511,N_22812,N_22699);
and UO_2512 (O_2512,N_24269,N_22987);
nand UO_2513 (O_2513,N_23189,N_22419);
or UO_2514 (O_2514,N_23946,N_22177);
or UO_2515 (O_2515,N_22181,N_22236);
and UO_2516 (O_2516,N_22715,N_22138);
xnor UO_2517 (O_2517,N_24604,N_21916);
or UO_2518 (O_2518,N_22391,N_22953);
or UO_2519 (O_2519,N_22185,N_23511);
and UO_2520 (O_2520,N_23458,N_23156);
nand UO_2521 (O_2521,N_23789,N_23498);
or UO_2522 (O_2522,N_24337,N_22181);
or UO_2523 (O_2523,N_22917,N_24381);
or UO_2524 (O_2524,N_24824,N_23356);
and UO_2525 (O_2525,N_21988,N_22772);
or UO_2526 (O_2526,N_24598,N_24323);
nor UO_2527 (O_2527,N_23350,N_22725);
xor UO_2528 (O_2528,N_23429,N_24778);
nand UO_2529 (O_2529,N_21945,N_22535);
and UO_2530 (O_2530,N_24274,N_22282);
nor UO_2531 (O_2531,N_24078,N_21983);
nor UO_2532 (O_2532,N_22280,N_22664);
and UO_2533 (O_2533,N_23975,N_23938);
xor UO_2534 (O_2534,N_24230,N_23302);
or UO_2535 (O_2535,N_24721,N_22279);
xnor UO_2536 (O_2536,N_24448,N_24781);
and UO_2537 (O_2537,N_21894,N_23404);
and UO_2538 (O_2538,N_22719,N_24811);
nand UO_2539 (O_2539,N_22541,N_21908);
or UO_2540 (O_2540,N_22689,N_23341);
nor UO_2541 (O_2541,N_24738,N_22484);
nand UO_2542 (O_2542,N_24997,N_23416);
or UO_2543 (O_2543,N_24294,N_23737);
and UO_2544 (O_2544,N_24072,N_24505);
and UO_2545 (O_2545,N_23020,N_24177);
xor UO_2546 (O_2546,N_22185,N_23260);
nand UO_2547 (O_2547,N_23463,N_22655);
and UO_2548 (O_2548,N_24407,N_23065);
nor UO_2549 (O_2549,N_23487,N_23999);
nor UO_2550 (O_2550,N_24674,N_23698);
and UO_2551 (O_2551,N_22739,N_23676);
or UO_2552 (O_2552,N_22224,N_23663);
xor UO_2553 (O_2553,N_24795,N_21980);
nand UO_2554 (O_2554,N_22088,N_22528);
xor UO_2555 (O_2555,N_23447,N_22035);
and UO_2556 (O_2556,N_23474,N_24791);
or UO_2557 (O_2557,N_21895,N_22642);
and UO_2558 (O_2558,N_22473,N_23035);
nor UO_2559 (O_2559,N_24343,N_22588);
nand UO_2560 (O_2560,N_23268,N_22332);
and UO_2561 (O_2561,N_24179,N_24577);
nor UO_2562 (O_2562,N_24561,N_24346);
xnor UO_2563 (O_2563,N_24543,N_23156);
or UO_2564 (O_2564,N_24105,N_24403);
nor UO_2565 (O_2565,N_23236,N_24674);
nand UO_2566 (O_2566,N_21990,N_23317);
xnor UO_2567 (O_2567,N_22193,N_23987);
xnor UO_2568 (O_2568,N_22407,N_21900);
or UO_2569 (O_2569,N_22827,N_23319);
nor UO_2570 (O_2570,N_23904,N_24263);
nand UO_2571 (O_2571,N_22481,N_23939);
nor UO_2572 (O_2572,N_23788,N_23139);
xor UO_2573 (O_2573,N_23486,N_22568);
or UO_2574 (O_2574,N_23761,N_24483);
or UO_2575 (O_2575,N_23812,N_24841);
nor UO_2576 (O_2576,N_24629,N_24935);
nor UO_2577 (O_2577,N_23674,N_23112);
nand UO_2578 (O_2578,N_23965,N_24530);
nor UO_2579 (O_2579,N_24945,N_23533);
and UO_2580 (O_2580,N_23360,N_23682);
nand UO_2581 (O_2581,N_24283,N_24814);
nand UO_2582 (O_2582,N_24281,N_22779);
nand UO_2583 (O_2583,N_24117,N_24491);
nor UO_2584 (O_2584,N_22417,N_24709);
nor UO_2585 (O_2585,N_24529,N_24865);
and UO_2586 (O_2586,N_22139,N_22495);
nor UO_2587 (O_2587,N_23213,N_24774);
nor UO_2588 (O_2588,N_22442,N_23349);
nor UO_2589 (O_2589,N_23197,N_22024);
or UO_2590 (O_2590,N_22999,N_23571);
nand UO_2591 (O_2591,N_22691,N_24444);
and UO_2592 (O_2592,N_23466,N_22969);
or UO_2593 (O_2593,N_23566,N_22548);
and UO_2594 (O_2594,N_22080,N_23720);
xnor UO_2595 (O_2595,N_23711,N_23540);
nor UO_2596 (O_2596,N_24527,N_22966);
nand UO_2597 (O_2597,N_22995,N_24201);
nand UO_2598 (O_2598,N_22708,N_22141);
xor UO_2599 (O_2599,N_23905,N_24138);
nand UO_2600 (O_2600,N_22132,N_23484);
xor UO_2601 (O_2601,N_24660,N_22137);
nand UO_2602 (O_2602,N_24514,N_24885);
nand UO_2603 (O_2603,N_22575,N_23992);
xor UO_2604 (O_2604,N_24891,N_24792);
and UO_2605 (O_2605,N_23443,N_24249);
or UO_2606 (O_2606,N_23022,N_23008);
nor UO_2607 (O_2607,N_24609,N_24913);
and UO_2608 (O_2608,N_22646,N_23484);
nor UO_2609 (O_2609,N_24375,N_22872);
and UO_2610 (O_2610,N_23481,N_24238);
or UO_2611 (O_2611,N_22832,N_24115);
nand UO_2612 (O_2612,N_22469,N_24239);
or UO_2613 (O_2613,N_23386,N_22045);
or UO_2614 (O_2614,N_24388,N_23824);
and UO_2615 (O_2615,N_23905,N_22900);
xnor UO_2616 (O_2616,N_22009,N_23686);
or UO_2617 (O_2617,N_22500,N_23304);
or UO_2618 (O_2618,N_22103,N_23437);
nand UO_2619 (O_2619,N_24837,N_22984);
or UO_2620 (O_2620,N_22085,N_22655);
and UO_2621 (O_2621,N_24718,N_23639);
xor UO_2622 (O_2622,N_22476,N_22208);
nand UO_2623 (O_2623,N_24306,N_24686);
nand UO_2624 (O_2624,N_22310,N_22089);
nand UO_2625 (O_2625,N_23717,N_22035);
or UO_2626 (O_2626,N_22810,N_24983);
and UO_2627 (O_2627,N_22357,N_24978);
nor UO_2628 (O_2628,N_23166,N_24327);
nand UO_2629 (O_2629,N_24100,N_22122);
or UO_2630 (O_2630,N_24567,N_22813);
xor UO_2631 (O_2631,N_22067,N_24014);
nor UO_2632 (O_2632,N_22376,N_23826);
or UO_2633 (O_2633,N_22176,N_22200);
and UO_2634 (O_2634,N_22836,N_23042);
or UO_2635 (O_2635,N_23943,N_24271);
and UO_2636 (O_2636,N_21885,N_24946);
nor UO_2637 (O_2637,N_22626,N_23545);
and UO_2638 (O_2638,N_23796,N_22401);
nand UO_2639 (O_2639,N_21911,N_22137);
nor UO_2640 (O_2640,N_22757,N_23457);
and UO_2641 (O_2641,N_24601,N_23501);
nor UO_2642 (O_2642,N_22643,N_23326);
nand UO_2643 (O_2643,N_23017,N_22529);
nor UO_2644 (O_2644,N_22242,N_24208);
nand UO_2645 (O_2645,N_23811,N_23226);
or UO_2646 (O_2646,N_23568,N_24545);
xnor UO_2647 (O_2647,N_22564,N_22930);
nor UO_2648 (O_2648,N_23277,N_23057);
and UO_2649 (O_2649,N_24003,N_22408);
or UO_2650 (O_2650,N_23445,N_22668);
and UO_2651 (O_2651,N_21993,N_23033);
nor UO_2652 (O_2652,N_22775,N_22188);
or UO_2653 (O_2653,N_23049,N_22246);
or UO_2654 (O_2654,N_24660,N_24869);
nor UO_2655 (O_2655,N_23543,N_22097);
and UO_2656 (O_2656,N_22228,N_24342);
and UO_2657 (O_2657,N_22560,N_23006);
nand UO_2658 (O_2658,N_22561,N_22404);
or UO_2659 (O_2659,N_21908,N_22073);
nor UO_2660 (O_2660,N_23027,N_23856);
nor UO_2661 (O_2661,N_21929,N_22076);
nand UO_2662 (O_2662,N_23199,N_23098);
nor UO_2663 (O_2663,N_22351,N_24879);
xor UO_2664 (O_2664,N_22518,N_24820);
xor UO_2665 (O_2665,N_22563,N_24746);
nor UO_2666 (O_2666,N_24678,N_22903);
and UO_2667 (O_2667,N_22151,N_22177);
or UO_2668 (O_2668,N_24107,N_22308);
or UO_2669 (O_2669,N_22033,N_22659);
nand UO_2670 (O_2670,N_22624,N_22732);
or UO_2671 (O_2671,N_24674,N_24806);
and UO_2672 (O_2672,N_24790,N_22864);
nor UO_2673 (O_2673,N_24457,N_23391);
and UO_2674 (O_2674,N_21956,N_23596);
and UO_2675 (O_2675,N_24226,N_23788);
nand UO_2676 (O_2676,N_23325,N_21927);
or UO_2677 (O_2677,N_24779,N_23889);
or UO_2678 (O_2678,N_21917,N_24740);
or UO_2679 (O_2679,N_24890,N_24907);
nand UO_2680 (O_2680,N_23346,N_24363);
nor UO_2681 (O_2681,N_24464,N_24086);
nor UO_2682 (O_2682,N_24383,N_22367);
xnor UO_2683 (O_2683,N_22507,N_22274);
and UO_2684 (O_2684,N_23200,N_23047);
nor UO_2685 (O_2685,N_24483,N_24097);
nor UO_2686 (O_2686,N_21915,N_23732);
nand UO_2687 (O_2687,N_23258,N_24742);
xor UO_2688 (O_2688,N_22595,N_23831);
or UO_2689 (O_2689,N_24566,N_24786);
nand UO_2690 (O_2690,N_23162,N_24426);
nand UO_2691 (O_2691,N_23144,N_23465);
nor UO_2692 (O_2692,N_24197,N_23887);
nand UO_2693 (O_2693,N_22062,N_23290);
xor UO_2694 (O_2694,N_24572,N_24482);
nand UO_2695 (O_2695,N_23202,N_24286);
and UO_2696 (O_2696,N_23852,N_23271);
nand UO_2697 (O_2697,N_23629,N_24944);
xnor UO_2698 (O_2698,N_22809,N_24390);
and UO_2699 (O_2699,N_23817,N_22082);
and UO_2700 (O_2700,N_24291,N_22281);
or UO_2701 (O_2701,N_22935,N_24635);
nand UO_2702 (O_2702,N_21898,N_23099);
nor UO_2703 (O_2703,N_24879,N_22214);
xor UO_2704 (O_2704,N_21910,N_22350);
or UO_2705 (O_2705,N_24462,N_24271);
and UO_2706 (O_2706,N_23661,N_22342);
and UO_2707 (O_2707,N_24211,N_24423);
or UO_2708 (O_2708,N_23572,N_22803);
and UO_2709 (O_2709,N_22885,N_22481);
or UO_2710 (O_2710,N_22424,N_22525);
xnor UO_2711 (O_2711,N_24845,N_24268);
nand UO_2712 (O_2712,N_23582,N_21934);
xor UO_2713 (O_2713,N_23613,N_22098);
and UO_2714 (O_2714,N_23066,N_23198);
or UO_2715 (O_2715,N_24969,N_24987);
nor UO_2716 (O_2716,N_23432,N_23672);
or UO_2717 (O_2717,N_24424,N_24103);
nor UO_2718 (O_2718,N_24316,N_21947);
or UO_2719 (O_2719,N_24909,N_24732);
nor UO_2720 (O_2720,N_24103,N_24979);
or UO_2721 (O_2721,N_22628,N_22232);
nand UO_2722 (O_2722,N_24896,N_22584);
or UO_2723 (O_2723,N_24065,N_23207);
nor UO_2724 (O_2724,N_24075,N_24467);
xnor UO_2725 (O_2725,N_22714,N_24484);
nand UO_2726 (O_2726,N_23902,N_24654);
and UO_2727 (O_2727,N_23764,N_22947);
and UO_2728 (O_2728,N_24559,N_22078);
and UO_2729 (O_2729,N_24629,N_23720);
or UO_2730 (O_2730,N_24677,N_24121);
nand UO_2731 (O_2731,N_23061,N_23229);
or UO_2732 (O_2732,N_22366,N_22042);
xnor UO_2733 (O_2733,N_23226,N_22620);
and UO_2734 (O_2734,N_22157,N_22547);
or UO_2735 (O_2735,N_24946,N_24415);
or UO_2736 (O_2736,N_24504,N_24112);
xor UO_2737 (O_2737,N_22489,N_24505);
and UO_2738 (O_2738,N_23953,N_24386);
or UO_2739 (O_2739,N_23776,N_22435);
nor UO_2740 (O_2740,N_23875,N_22454);
or UO_2741 (O_2741,N_24726,N_22510);
and UO_2742 (O_2742,N_24315,N_24301);
xor UO_2743 (O_2743,N_24722,N_22402);
and UO_2744 (O_2744,N_23071,N_22408);
or UO_2745 (O_2745,N_24231,N_22704);
or UO_2746 (O_2746,N_23372,N_22876);
and UO_2747 (O_2747,N_24490,N_23108);
nand UO_2748 (O_2748,N_22163,N_23469);
nor UO_2749 (O_2749,N_24437,N_22582);
and UO_2750 (O_2750,N_22460,N_24276);
xor UO_2751 (O_2751,N_22734,N_22951);
and UO_2752 (O_2752,N_24741,N_24935);
nand UO_2753 (O_2753,N_23456,N_23365);
nand UO_2754 (O_2754,N_24109,N_22976);
nand UO_2755 (O_2755,N_21957,N_22735);
nor UO_2756 (O_2756,N_24555,N_22459);
and UO_2757 (O_2757,N_23272,N_22111);
nand UO_2758 (O_2758,N_22912,N_23865);
nand UO_2759 (O_2759,N_24817,N_24369);
and UO_2760 (O_2760,N_22751,N_22743);
nand UO_2761 (O_2761,N_22104,N_23735);
nor UO_2762 (O_2762,N_22797,N_24607);
xor UO_2763 (O_2763,N_24989,N_22351);
nand UO_2764 (O_2764,N_24203,N_22715);
nor UO_2765 (O_2765,N_22276,N_24846);
or UO_2766 (O_2766,N_22609,N_24707);
nand UO_2767 (O_2767,N_22447,N_23364);
nor UO_2768 (O_2768,N_22814,N_24371);
nand UO_2769 (O_2769,N_22194,N_24814);
and UO_2770 (O_2770,N_23018,N_24083);
nand UO_2771 (O_2771,N_23531,N_23986);
nand UO_2772 (O_2772,N_24336,N_22437);
nand UO_2773 (O_2773,N_23432,N_21998);
nor UO_2774 (O_2774,N_23276,N_22636);
and UO_2775 (O_2775,N_22036,N_24139);
nand UO_2776 (O_2776,N_21896,N_22026);
and UO_2777 (O_2777,N_22014,N_22517);
nor UO_2778 (O_2778,N_21995,N_23153);
nor UO_2779 (O_2779,N_23447,N_22451);
and UO_2780 (O_2780,N_22099,N_22649);
nand UO_2781 (O_2781,N_23965,N_24971);
nor UO_2782 (O_2782,N_23185,N_21894);
nand UO_2783 (O_2783,N_23644,N_21917);
nor UO_2784 (O_2784,N_24088,N_24646);
or UO_2785 (O_2785,N_22481,N_22596);
xor UO_2786 (O_2786,N_22953,N_24176);
or UO_2787 (O_2787,N_22108,N_24171);
nor UO_2788 (O_2788,N_22316,N_22350);
nand UO_2789 (O_2789,N_23631,N_22479);
and UO_2790 (O_2790,N_22997,N_23909);
nor UO_2791 (O_2791,N_22806,N_23403);
or UO_2792 (O_2792,N_23531,N_23406);
or UO_2793 (O_2793,N_24006,N_22035);
nand UO_2794 (O_2794,N_22271,N_24155);
nor UO_2795 (O_2795,N_23684,N_24887);
xor UO_2796 (O_2796,N_24649,N_24105);
nor UO_2797 (O_2797,N_23225,N_24840);
nor UO_2798 (O_2798,N_23011,N_22884);
and UO_2799 (O_2799,N_22309,N_23223);
or UO_2800 (O_2800,N_22168,N_23082);
nor UO_2801 (O_2801,N_24141,N_22910);
or UO_2802 (O_2802,N_22032,N_22978);
nor UO_2803 (O_2803,N_23638,N_23324);
nor UO_2804 (O_2804,N_22972,N_24787);
xor UO_2805 (O_2805,N_21965,N_24722);
nand UO_2806 (O_2806,N_23550,N_23428);
or UO_2807 (O_2807,N_23706,N_22788);
and UO_2808 (O_2808,N_22118,N_22001);
or UO_2809 (O_2809,N_24297,N_22464);
nand UO_2810 (O_2810,N_22285,N_23232);
and UO_2811 (O_2811,N_24465,N_23766);
nor UO_2812 (O_2812,N_22457,N_23969);
nand UO_2813 (O_2813,N_24869,N_24117);
and UO_2814 (O_2814,N_23795,N_22127);
and UO_2815 (O_2815,N_24938,N_24682);
nor UO_2816 (O_2816,N_24365,N_23599);
and UO_2817 (O_2817,N_23621,N_23450);
nor UO_2818 (O_2818,N_22840,N_24886);
and UO_2819 (O_2819,N_23976,N_21914);
nand UO_2820 (O_2820,N_24349,N_24916);
nand UO_2821 (O_2821,N_22415,N_22236);
and UO_2822 (O_2822,N_22995,N_22316);
nor UO_2823 (O_2823,N_24601,N_24732);
nand UO_2824 (O_2824,N_24552,N_21886);
or UO_2825 (O_2825,N_24764,N_22048);
nand UO_2826 (O_2826,N_24582,N_24288);
xor UO_2827 (O_2827,N_22742,N_23426);
nor UO_2828 (O_2828,N_22570,N_23894);
nor UO_2829 (O_2829,N_23074,N_24210);
nand UO_2830 (O_2830,N_22675,N_22866);
nor UO_2831 (O_2831,N_23967,N_24988);
nand UO_2832 (O_2832,N_24026,N_23760);
nand UO_2833 (O_2833,N_23145,N_24737);
or UO_2834 (O_2834,N_22227,N_22667);
nor UO_2835 (O_2835,N_22420,N_23074);
nor UO_2836 (O_2836,N_24263,N_23885);
nand UO_2837 (O_2837,N_23754,N_23583);
and UO_2838 (O_2838,N_24191,N_22056);
and UO_2839 (O_2839,N_23013,N_23709);
xor UO_2840 (O_2840,N_24392,N_22668);
nor UO_2841 (O_2841,N_23573,N_23746);
xor UO_2842 (O_2842,N_24083,N_23758);
or UO_2843 (O_2843,N_22783,N_22637);
or UO_2844 (O_2844,N_24144,N_24541);
and UO_2845 (O_2845,N_23723,N_22336);
nand UO_2846 (O_2846,N_23774,N_24783);
or UO_2847 (O_2847,N_22703,N_24456);
nor UO_2848 (O_2848,N_24612,N_23526);
nor UO_2849 (O_2849,N_23686,N_24619);
xor UO_2850 (O_2850,N_22225,N_22334);
and UO_2851 (O_2851,N_22386,N_23603);
nor UO_2852 (O_2852,N_22095,N_22765);
nor UO_2853 (O_2853,N_24750,N_23422);
nor UO_2854 (O_2854,N_22436,N_23828);
nor UO_2855 (O_2855,N_23740,N_23469);
nand UO_2856 (O_2856,N_22373,N_23984);
nand UO_2857 (O_2857,N_24991,N_23282);
and UO_2858 (O_2858,N_23139,N_23252);
xor UO_2859 (O_2859,N_22117,N_23522);
and UO_2860 (O_2860,N_22336,N_24661);
and UO_2861 (O_2861,N_23764,N_22518);
or UO_2862 (O_2862,N_24436,N_22331);
or UO_2863 (O_2863,N_23211,N_23386);
or UO_2864 (O_2864,N_24257,N_23490);
xor UO_2865 (O_2865,N_24873,N_24381);
and UO_2866 (O_2866,N_22406,N_24918);
xnor UO_2867 (O_2867,N_23766,N_23267);
and UO_2868 (O_2868,N_23184,N_22144);
or UO_2869 (O_2869,N_22016,N_23090);
nor UO_2870 (O_2870,N_23005,N_24805);
nor UO_2871 (O_2871,N_23467,N_22703);
and UO_2872 (O_2872,N_24692,N_24837);
or UO_2873 (O_2873,N_22034,N_24480);
or UO_2874 (O_2874,N_22649,N_24553);
nor UO_2875 (O_2875,N_22979,N_22534);
nand UO_2876 (O_2876,N_24614,N_22478);
nand UO_2877 (O_2877,N_24682,N_22585);
xnor UO_2878 (O_2878,N_24058,N_21997);
or UO_2879 (O_2879,N_22588,N_22536);
xnor UO_2880 (O_2880,N_23350,N_22316);
nor UO_2881 (O_2881,N_24489,N_24162);
or UO_2882 (O_2882,N_24702,N_23406);
nor UO_2883 (O_2883,N_23419,N_23614);
and UO_2884 (O_2884,N_22040,N_23877);
nor UO_2885 (O_2885,N_22103,N_24453);
nand UO_2886 (O_2886,N_24129,N_24889);
nand UO_2887 (O_2887,N_24993,N_22104);
nor UO_2888 (O_2888,N_24948,N_24289);
and UO_2889 (O_2889,N_24514,N_23054);
nand UO_2890 (O_2890,N_22045,N_24993);
or UO_2891 (O_2891,N_23956,N_24988);
xor UO_2892 (O_2892,N_24518,N_24614);
nand UO_2893 (O_2893,N_22642,N_23684);
and UO_2894 (O_2894,N_23301,N_22062);
nor UO_2895 (O_2895,N_22403,N_22280);
nor UO_2896 (O_2896,N_23853,N_24249);
nor UO_2897 (O_2897,N_24569,N_24033);
or UO_2898 (O_2898,N_22577,N_22527);
and UO_2899 (O_2899,N_24648,N_21877);
nand UO_2900 (O_2900,N_22373,N_24882);
and UO_2901 (O_2901,N_23503,N_22552);
nor UO_2902 (O_2902,N_21898,N_24382);
xor UO_2903 (O_2903,N_24179,N_23139);
nand UO_2904 (O_2904,N_22164,N_23306);
or UO_2905 (O_2905,N_22371,N_22230);
and UO_2906 (O_2906,N_24663,N_23892);
and UO_2907 (O_2907,N_22443,N_23223);
nor UO_2908 (O_2908,N_22248,N_23059);
and UO_2909 (O_2909,N_24184,N_22250);
nand UO_2910 (O_2910,N_24471,N_22570);
nand UO_2911 (O_2911,N_23137,N_24693);
nor UO_2912 (O_2912,N_22151,N_22998);
nand UO_2913 (O_2913,N_23951,N_22632);
or UO_2914 (O_2914,N_23669,N_22769);
and UO_2915 (O_2915,N_23781,N_22581);
and UO_2916 (O_2916,N_22423,N_24109);
nand UO_2917 (O_2917,N_23947,N_23598);
xnor UO_2918 (O_2918,N_22048,N_24282);
and UO_2919 (O_2919,N_23793,N_22527);
nand UO_2920 (O_2920,N_23038,N_23903);
or UO_2921 (O_2921,N_23498,N_23233);
nand UO_2922 (O_2922,N_24230,N_23734);
nand UO_2923 (O_2923,N_23576,N_23590);
or UO_2924 (O_2924,N_22313,N_24451);
and UO_2925 (O_2925,N_24021,N_24741);
and UO_2926 (O_2926,N_23672,N_22590);
nor UO_2927 (O_2927,N_23187,N_22043);
and UO_2928 (O_2928,N_24116,N_24703);
and UO_2929 (O_2929,N_23548,N_24229);
xnor UO_2930 (O_2930,N_23746,N_22856);
and UO_2931 (O_2931,N_23941,N_24627);
nand UO_2932 (O_2932,N_24023,N_22855);
and UO_2933 (O_2933,N_24181,N_24268);
nor UO_2934 (O_2934,N_23185,N_23246);
nand UO_2935 (O_2935,N_22018,N_23676);
nor UO_2936 (O_2936,N_23824,N_24896);
nor UO_2937 (O_2937,N_23106,N_23126);
and UO_2938 (O_2938,N_23796,N_22086);
nor UO_2939 (O_2939,N_24685,N_24441);
nand UO_2940 (O_2940,N_24521,N_21980);
or UO_2941 (O_2941,N_22138,N_23662);
nand UO_2942 (O_2942,N_22150,N_22767);
nand UO_2943 (O_2943,N_23138,N_24733);
nor UO_2944 (O_2944,N_23410,N_21967);
or UO_2945 (O_2945,N_22533,N_24098);
nand UO_2946 (O_2946,N_22078,N_24814);
nor UO_2947 (O_2947,N_24785,N_23105);
or UO_2948 (O_2948,N_22989,N_23183);
nand UO_2949 (O_2949,N_24375,N_23755);
nor UO_2950 (O_2950,N_21889,N_22285);
and UO_2951 (O_2951,N_23254,N_23380);
nor UO_2952 (O_2952,N_23246,N_22758);
or UO_2953 (O_2953,N_22228,N_24685);
nor UO_2954 (O_2954,N_21983,N_23552);
and UO_2955 (O_2955,N_23867,N_23045);
and UO_2956 (O_2956,N_24933,N_22982);
or UO_2957 (O_2957,N_22955,N_24442);
nor UO_2958 (O_2958,N_22114,N_22045);
nor UO_2959 (O_2959,N_22709,N_22936);
xor UO_2960 (O_2960,N_23290,N_23099);
and UO_2961 (O_2961,N_22193,N_21951);
nand UO_2962 (O_2962,N_22241,N_21943);
and UO_2963 (O_2963,N_22969,N_23924);
nand UO_2964 (O_2964,N_22346,N_24006);
nand UO_2965 (O_2965,N_23825,N_24352);
and UO_2966 (O_2966,N_24270,N_22484);
and UO_2967 (O_2967,N_24319,N_23147);
and UO_2968 (O_2968,N_24437,N_23131);
nor UO_2969 (O_2969,N_24275,N_23667);
or UO_2970 (O_2970,N_23683,N_22627);
and UO_2971 (O_2971,N_23766,N_23342);
xnor UO_2972 (O_2972,N_24993,N_23751);
and UO_2973 (O_2973,N_23127,N_22790);
and UO_2974 (O_2974,N_24175,N_22692);
nor UO_2975 (O_2975,N_24602,N_22971);
and UO_2976 (O_2976,N_23753,N_22775);
and UO_2977 (O_2977,N_22313,N_24475);
and UO_2978 (O_2978,N_23478,N_22808);
or UO_2979 (O_2979,N_23409,N_23674);
nor UO_2980 (O_2980,N_24942,N_22512);
and UO_2981 (O_2981,N_22788,N_24507);
nor UO_2982 (O_2982,N_24055,N_22889);
and UO_2983 (O_2983,N_23017,N_22242);
xor UO_2984 (O_2984,N_24130,N_22114);
xnor UO_2985 (O_2985,N_23947,N_22998);
and UO_2986 (O_2986,N_24837,N_23837);
xnor UO_2987 (O_2987,N_23297,N_23273);
nor UO_2988 (O_2988,N_24085,N_22151);
nor UO_2989 (O_2989,N_24216,N_24140);
and UO_2990 (O_2990,N_23061,N_23667);
xor UO_2991 (O_2991,N_24197,N_22341);
and UO_2992 (O_2992,N_21896,N_22671);
nor UO_2993 (O_2993,N_22779,N_24942);
or UO_2994 (O_2994,N_22879,N_24929);
and UO_2995 (O_2995,N_22600,N_23220);
and UO_2996 (O_2996,N_24562,N_24660);
and UO_2997 (O_2997,N_22304,N_24501);
and UO_2998 (O_2998,N_24327,N_23117);
and UO_2999 (O_2999,N_24033,N_23322);
endmodule