module basic_1500_15000_2000_120_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_612,In_1161);
xor U1 (N_1,In_780,In_658);
xor U2 (N_2,In_1427,In_1139);
xor U3 (N_3,In_944,In_820);
or U4 (N_4,In_1119,In_359);
xnor U5 (N_5,In_33,In_815);
and U6 (N_6,In_760,In_867);
nand U7 (N_7,In_273,In_446);
or U8 (N_8,In_902,In_769);
nand U9 (N_9,In_739,In_1127);
and U10 (N_10,In_877,In_159);
xor U11 (N_11,In_244,In_556);
or U12 (N_12,In_1415,In_1066);
nor U13 (N_13,In_215,In_1272);
xor U14 (N_14,In_371,In_714);
and U15 (N_15,In_781,In_202);
and U16 (N_16,In_126,In_532);
xnor U17 (N_17,In_675,In_942);
and U18 (N_18,In_1038,In_285);
or U19 (N_19,In_919,In_239);
xor U20 (N_20,In_205,In_542);
xnor U21 (N_21,In_1394,In_649);
xnor U22 (N_22,In_292,In_1336);
and U23 (N_23,In_3,In_1190);
xor U24 (N_24,In_138,In_331);
nor U25 (N_25,In_1383,In_1247);
nand U26 (N_26,In_1406,In_523);
and U27 (N_27,In_416,In_408);
or U28 (N_28,In_601,In_551);
xor U29 (N_29,In_1124,In_834);
and U30 (N_30,In_892,In_741);
xnor U31 (N_31,In_364,In_878);
xor U32 (N_32,In_317,In_924);
or U33 (N_33,In_1085,In_754);
nand U34 (N_34,In_1377,In_825);
xor U35 (N_35,In_1293,In_483);
or U36 (N_36,In_797,In_955);
and U37 (N_37,In_170,In_271);
nand U38 (N_38,In_1051,In_132);
nor U39 (N_39,In_558,In_861);
nand U40 (N_40,In_354,In_162);
and U41 (N_41,In_241,In_787);
or U42 (N_42,In_397,In_898);
xnor U43 (N_43,In_534,In_1153);
nor U44 (N_44,In_1009,In_435);
nand U45 (N_45,In_1226,In_913);
nor U46 (N_46,In_802,In_581);
xnor U47 (N_47,In_335,In_607);
or U48 (N_48,In_1180,In_1351);
and U49 (N_49,In_1441,In_488);
nand U50 (N_50,In_885,In_835);
nor U51 (N_51,In_1388,In_1392);
xnor U52 (N_52,In_939,In_1007);
and U53 (N_53,In_1491,In_169);
xnor U54 (N_54,In_310,In_24);
or U55 (N_55,In_712,In_1474);
nand U56 (N_56,In_1454,In_1116);
or U57 (N_57,In_938,In_383);
or U58 (N_58,In_1154,In_590);
xnor U59 (N_59,In_1198,In_1283);
and U60 (N_60,In_710,In_544);
and U61 (N_61,In_728,In_738);
and U62 (N_62,In_194,In_398);
and U63 (N_63,In_909,In_1270);
xnor U64 (N_64,In_676,In_584);
xor U65 (N_65,In_396,In_1481);
or U66 (N_66,In_69,In_429);
or U67 (N_67,In_485,In_887);
and U68 (N_68,In_1475,In_507);
or U69 (N_69,In_744,In_1445);
nor U70 (N_70,In_286,In_618);
and U71 (N_71,In_390,In_1488);
xnor U72 (N_72,In_980,In_60);
or U73 (N_73,In_452,In_831);
xor U74 (N_74,In_325,In_360);
nand U75 (N_75,In_236,In_1160);
or U76 (N_76,In_1387,In_954);
nand U77 (N_77,In_1232,In_756);
nand U78 (N_78,In_56,In_962);
nand U79 (N_79,In_685,In_260);
or U80 (N_80,In_621,In_920);
nand U81 (N_81,In_414,In_168);
nand U82 (N_82,In_573,In_1109);
and U83 (N_83,In_255,In_245);
nor U84 (N_84,In_845,In_234);
xnor U85 (N_85,In_425,In_71);
nor U86 (N_86,In_1442,In_1296);
nor U87 (N_87,In_1027,In_1311);
nor U88 (N_88,In_571,In_1013);
and U89 (N_89,In_131,In_1255);
nor U90 (N_90,In_1337,In_119);
nand U91 (N_91,In_596,In_998);
nand U92 (N_92,In_1464,In_953);
and U93 (N_93,In_283,In_1142);
or U94 (N_94,In_631,In_536);
or U95 (N_95,In_546,In_748);
nor U96 (N_96,In_970,In_1050);
nand U97 (N_97,In_883,In_904);
nand U98 (N_98,In_86,In_1405);
nor U99 (N_99,In_718,In_231);
or U100 (N_100,In_874,In_143);
and U101 (N_101,In_1147,In_1469);
or U102 (N_102,In_145,In_48);
xor U103 (N_103,In_1301,In_716);
nand U104 (N_104,In_243,In_193);
and U105 (N_105,In_495,In_1400);
nand U106 (N_106,In_1067,In_54);
xor U107 (N_107,In_1094,In_1416);
xor U108 (N_108,In_931,In_1429);
or U109 (N_109,In_1058,In_430);
and U110 (N_110,In_448,In_295);
xor U111 (N_111,In_721,In_1450);
xor U112 (N_112,In_1318,In_380);
xor U113 (N_113,In_1288,In_413);
or U114 (N_114,In_735,In_513);
nor U115 (N_115,In_966,In_1365);
nand U116 (N_116,In_696,In_1290);
nand U117 (N_117,In_727,In_646);
nand U118 (N_118,In_777,In_1184);
nor U119 (N_119,In_1167,In_1343);
and U120 (N_120,In_404,In_1494);
and U121 (N_121,In_1054,In_855);
and U122 (N_122,In_1156,In_580);
xor U123 (N_123,In_180,In_148);
nand U124 (N_124,In_1059,In_625);
xor U125 (N_125,In_809,In_1499);
or U126 (N_126,In_102,In_740);
xor U127 (N_127,In_31,N_25);
or U128 (N_128,In_183,In_1462);
or U129 (N_129,In_1074,N_21);
or U130 (N_130,In_1209,In_43);
nand U131 (N_131,In_1331,In_147);
nor U132 (N_132,In_703,In_936);
nor U133 (N_133,In_784,In_237);
and U134 (N_134,In_116,In_1271);
or U135 (N_135,In_345,In_1277);
nor U136 (N_136,In_896,In_274);
and U137 (N_137,In_402,In_1287);
and U138 (N_138,In_788,In_491);
or U139 (N_139,In_1137,In_313);
or U140 (N_140,In_14,N_23);
nand U141 (N_141,N_38,In_562);
and U142 (N_142,In_349,N_15);
xnor U143 (N_143,In_582,In_606);
nand U144 (N_144,N_31,In_643);
nand U145 (N_145,In_689,In_1436);
nor U146 (N_146,In_1261,In_1123);
xnor U147 (N_147,In_254,In_269);
xnor U148 (N_148,In_1303,In_932);
nor U149 (N_149,In_806,In_732);
and U150 (N_150,In_419,In_1157);
nand U151 (N_151,In_620,In_474);
and U152 (N_152,In_1477,In_1448);
xor U153 (N_153,In_945,In_709);
nor U154 (N_154,In_1332,In_1289);
and U155 (N_155,N_57,In_753);
or U156 (N_156,In_1170,In_400);
xor U157 (N_157,In_299,In_1186);
and U158 (N_158,In_1122,In_1078);
nand U159 (N_159,In_961,In_458);
or U160 (N_160,In_699,In_711);
nand U161 (N_161,In_336,In_795);
nand U162 (N_162,In_27,In_905);
nor U163 (N_163,In_1250,In_475);
and U164 (N_164,In_177,In_1158);
or U165 (N_165,In_541,In_1313);
nand U166 (N_166,In_768,In_440);
or U167 (N_167,In_41,In_1231);
xnor U168 (N_168,In_92,In_506);
or U169 (N_169,In_94,In_752);
or U170 (N_170,In_1487,In_978);
or U171 (N_171,In_1108,In_557);
or U172 (N_172,In_1335,In_468);
nor U173 (N_173,In_910,In_505);
nand U174 (N_174,In_736,N_105);
or U175 (N_175,In_73,In_288);
xnor U176 (N_176,In_1071,In_698);
or U177 (N_177,In_785,In_251);
nand U178 (N_178,In_512,In_1079);
nand U179 (N_179,In_1222,N_113);
or U180 (N_180,N_51,In_1361);
or U181 (N_181,In_516,In_278);
xnor U182 (N_182,In_770,N_30);
nand U183 (N_183,In_662,In_589);
nand U184 (N_184,N_29,In_280);
nor U185 (N_185,In_370,In_918);
xor U186 (N_186,In_720,In_1200);
xor U187 (N_187,In_833,In_303);
nor U188 (N_188,In_87,In_302);
nand U189 (N_189,In_20,In_935);
nand U190 (N_190,In_958,In_1446);
xnor U191 (N_191,In_1463,In_1461);
and U192 (N_192,N_91,In_713);
and U193 (N_193,In_977,In_1049);
and U194 (N_194,In_384,In_894);
and U195 (N_195,In_45,In_1372);
and U196 (N_196,In_1113,In_1149);
xor U197 (N_197,In_640,In_233);
nor U198 (N_198,In_1017,N_110);
nor U199 (N_199,N_102,N_59);
xor U200 (N_200,In_337,In_1401);
or U201 (N_201,N_32,In_628);
or U202 (N_202,In_778,In_1326);
nor U203 (N_203,In_708,N_13);
or U204 (N_204,In_1245,In_122);
or U205 (N_205,In_882,In_1181);
nor U206 (N_206,In_250,In_441);
nor U207 (N_207,In_249,In_213);
or U208 (N_208,In_53,In_263);
and U209 (N_209,In_749,N_27);
and U210 (N_210,In_1333,In_1279);
nor U211 (N_211,In_873,In_839);
xor U212 (N_212,In_117,In_659);
and U213 (N_213,In_912,In_563);
or U214 (N_214,In_1213,In_329);
and U215 (N_215,In_232,In_914);
or U216 (N_216,N_83,In_1177);
and U217 (N_217,In_1323,N_89);
or U218 (N_218,In_1374,In_1025);
and U219 (N_219,In_1032,In_750);
nor U220 (N_220,N_55,In_201);
nand U221 (N_221,In_1064,In_1422);
xor U222 (N_222,In_1362,N_98);
nand U223 (N_223,In_454,In_1080);
and U224 (N_224,In_547,In_890);
nand U225 (N_225,In_1233,In_805);
and U226 (N_226,In_1444,In_341);
nand U227 (N_227,N_36,In_1479);
xnor U228 (N_228,In_927,In_90);
nor U229 (N_229,In_995,In_683);
or U230 (N_230,In_1035,In_819);
nand U231 (N_231,In_410,N_56);
nor U232 (N_232,N_11,In_1033);
nor U233 (N_233,In_976,In_372);
nor U234 (N_234,In_949,N_22);
xnor U235 (N_235,N_74,In_991);
and U236 (N_236,In_219,In_1482);
nand U237 (N_237,N_104,In_543);
and U238 (N_238,In_1391,In_993);
nor U239 (N_239,N_5,In_210);
nand U240 (N_240,In_465,In_1098);
or U241 (N_241,In_992,In_1175);
nand U242 (N_242,In_864,In_476);
nor U243 (N_243,In_997,In_141);
xnor U244 (N_244,N_17,In_681);
nor U245 (N_245,In_1280,In_235);
xor U246 (N_246,In_17,In_665);
xor U247 (N_247,In_1041,In_479);
nand U248 (N_248,N_120,N_69);
nor U249 (N_249,In_636,In_179);
or U250 (N_250,In_262,In_137);
or U251 (N_251,In_511,In_1138);
nand U252 (N_252,In_1497,In_83);
xor U253 (N_253,In_828,In_520);
nand U254 (N_254,In_42,In_836);
or U255 (N_255,N_49,In_106);
and U256 (N_256,N_47,In_674);
xor U257 (N_257,In_967,In_1001);
nand U258 (N_258,In_0,In_308);
and U259 (N_259,In_1456,In_774);
nor U260 (N_260,In_1355,In_1126);
nand U261 (N_261,N_12,In_161);
and U262 (N_262,In_776,In_1384);
or U263 (N_263,In_1130,In_1129);
and U264 (N_264,In_1100,In_591);
nand U265 (N_265,In_841,In_1015);
xnor U266 (N_266,In_652,In_1110);
or U267 (N_267,In_1172,In_804);
nor U268 (N_268,In_144,In_587);
nor U269 (N_269,In_1452,In_943);
nand U270 (N_270,In_1063,In_859);
xnor U271 (N_271,In_810,In_605);
and U272 (N_272,In_737,In_1403);
nand U273 (N_273,In_690,In_97);
and U274 (N_274,In_1371,In_952);
nand U275 (N_275,In_1389,N_43);
nand U276 (N_276,In_352,In_579);
or U277 (N_277,In_478,In_1225);
and U278 (N_278,In_844,In_217);
nand U279 (N_279,In_218,In_1024);
nor U280 (N_280,In_617,In_807);
nor U281 (N_281,N_172,In_996);
nand U282 (N_282,N_230,N_72);
xnor U283 (N_283,In_525,In_188);
or U284 (N_284,In_394,In_1254);
xnor U285 (N_285,In_1359,In_379);
and U286 (N_286,In_610,In_100);
xnor U287 (N_287,In_880,In_930);
xor U288 (N_288,In_816,In_779);
nand U289 (N_289,In_694,In_1239);
nor U290 (N_290,In_228,In_627);
or U291 (N_291,In_1458,In_1368);
nand U292 (N_292,In_172,In_1349);
and U293 (N_293,In_875,In_1473);
xor U294 (N_294,In_985,In_1274);
or U295 (N_295,N_184,In_136);
nor U296 (N_296,In_548,In_1029);
xnor U297 (N_297,In_268,In_36);
or U298 (N_298,In_990,In_950);
xnor U299 (N_299,N_222,In_82);
and U300 (N_300,In_751,In_705);
and U301 (N_301,In_1056,In_850);
xnor U302 (N_302,In_1259,In_1484);
nand U303 (N_303,In_129,In_1055);
xnor U304 (N_304,In_1246,In_486);
nand U305 (N_305,N_175,In_1089);
nand U306 (N_306,In_956,In_704);
or U307 (N_307,In_406,In_1021);
xnor U308 (N_308,In_1470,N_177);
and U309 (N_309,In_515,In_164);
xnor U310 (N_310,In_18,In_553);
or U311 (N_311,In_1026,In_963);
xor U312 (N_312,In_1457,In_629);
nor U313 (N_313,In_570,In_790);
or U314 (N_314,In_1447,In_267);
nand U315 (N_315,N_204,In_490);
or U316 (N_316,In_473,N_48);
nand U317 (N_317,In_858,In_1189);
or U318 (N_318,N_130,N_199);
xor U319 (N_319,In_1424,In_1218);
nor U320 (N_320,In_1165,In_1162);
nor U321 (N_321,In_1312,In_1081);
or U322 (N_322,In_293,In_765);
nand U323 (N_323,N_241,N_92);
xnor U324 (N_324,In_901,In_971);
nor U325 (N_325,N_81,In_615);
nand U326 (N_326,N_60,In_1060);
xnor U327 (N_327,In_12,In_870);
nor U328 (N_328,In_1144,N_195);
xnor U329 (N_329,N_167,In_98);
nor U330 (N_330,In_456,In_1214);
nor U331 (N_331,In_363,In_879);
xor U332 (N_332,In_578,N_224);
and U333 (N_333,In_1199,In_261);
xor U334 (N_334,In_1315,In_1155);
nor U335 (N_335,In_598,In_847);
xnor U336 (N_336,In_554,In_789);
nor U337 (N_337,In_142,In_975);
xnor U338 (N_338,In_1438,In_895);
xor U339 (N_339,N_14,In_1466);
and U340 (N_340,In_450,In_811);
nand U341 (N_341,In_343,In_660);
and U342 (N_342,In_1182,In_1227);
nand U343 (N_343,In_1370,In_96);
or U344 (N_344,In_871,In_89);
nor U345 (N_345,In_731,In_1028);
nand U346 (N_346,N_214,In_772);
xnor U347 (N_347,In_127,In_560);
nand U348 (N_348,In_1097,In_114);
nor U349 (N_349,In_916,In_111);
nor U350 (N_350,In_801,In_1252);
nand U351 (N_351,In_291,In_1096);
nand U352 (N_352,In_632,In_214);
and U353 (N_353,In_13,In_1224);
or U354 (N_354,In_1215,In_298);
nor U355 (N_355,In_10,In_821);
nor U356 (N_356,N_111,In_614);
xor U357 (N_357,N_196,N_157);
nor U358 (N_358,In_1114,N_67);
and U359 (N_359,In_1393,In_595);
or U360 (N_360,In_823,In_284);
and U361 (N_361,In_891,In_366);
nand U362 (N_362,N_93,In_968);
and U363 (N_363,In_128,In_6);
nand U364 (N_364,N_203,In_51);
or U365 (N_365,In_687,N_193);
nor U366 (N_366,N_53,In_1240);
nand U367 (N_367,In_1188,N_154);
or U368 (N_368,In_593,In_677);
nor U369 (N_369,N_220,N_8);
nand U370 (N_370,In_1476,In_107);
nand U371 (N_371,In_64,In_1248);
nand U372 (N_372,In_1256,In_761);
and U373 (N_373,N_227,In_318);
nand U374 (N_374,N_164,In_600);
nand U375 (N_375,In_1203,In_32);
and U376 (N_376,In_763,N_202);
and U377 (N_377,In_1451,N_165);
nand U378 (N_378,N_304,In_477);
and U379 (N_379,N_46,In_758);
nand U380 (N_380,N_235,In_586);
or U381 (N_381,N_66,In_1273);
or U382 (N_382,In_1070,In_424);
xnor U383 (N_383,N_269,In_158);
or U384 (N_384,In_434,In_866);
and U385 (N_385,In_814,N_95);
nor U386 (N_386,In_767,N_245);
nand U387 (N_387,N_160,N_151);
nand U388 (N_388,In_851,In_986);
xor U389 (N_389,In_266,N_233);
nor U390 (N_390,In_1228,In_799);
and U391 (N_391,In_247,N_284);
nor U392 (N_392,N_19,In_258);
nor U393 (N_393,In_340,In_399);
or U394 (N_394,In_602,In_622);
xnor U395 (N_395,In_1202,In_984);
nand U396 (N_396,In_59,In_613);
xnor U397 (N_397,In_226,In_1434);
nor U398 (N_398,N_6,N_64);
nand U399 (N_399,N_140,In_1143);
nor U400 (N_400,In_1428,N_87);
or U401 (N_401,N_79,In_462);
or U402 (N_402,In_361,In_393);
nand U403 (N_403,In_881,N_124);
and U404 (N_404,In_746,In_29);
and U405 (N_405,In_668,N_285);
xor U406 (N_406,In_7,N_86);
nand U407 (N_407,In_496,In_467);
nor U408 (N_408,In_178,In_190);
or U409 (N_409,In_46,In_420);
and U410 (N_410,In_470,N_180);
and U411 (N_411,In_661,In_623);
nor U412 (N_412,In_74,In_1052);
and U413 (N_413,N_322,In_1235);
nand U414 (N_414,In_552,In_1297);
xnor U415 (N_415,In_1151,In_911);
nor U416 (N_416,N_237,In_925);
xor U417 (N_417,N_297,In_1364);
nand U418 (N_418,In_585,N_20);
or U419 (N_419,In_1347,In_466);
or U420 (N_420,N_145,In_577);
nor U421 (N_421,In_843,N_296);
nor U422 (N_422,N_82,In_155);
xnor U423 (N_423,In_389,In_9);
and U424 (N_424,In_65,In_530);
or U425 (N_425,In_1490,In_50);
or U426 (N_426,In_1241,In_837);
nor U427 (N_427,In_294,In_353);
xor U428 (N_428,In_522,N_213);
nor U429 (N_429,N_242,In_1093);
nor U430 (N_430,In_88,In_1354);
nand U431 (N_431,In_1201,In_907);
and U432 (N_432,In_742,In_1005);
or U433 (N_433,N_374,N_182);
nor U434 (N_434,In_1402,In_745);
or U435 (N_435,N_90,N_147);
or U436 (N_436,In_707,In_422);
nand U437 (N_437,In_1091,In_679);
and U438 (N_438,In_1133,N_240);
nand U439 (N_439,In_594,In_762);
or U440 (N_440,In_1229,In_1284);
nor U441 (N_441,In_1220,In_238);
or U442 (N_442,In_521,In_1195);
and U443 (N_443,In_264,N_362);
xor U444 (N_444,N_314,In_133);
and U445 (N_445,N_4,In_830);
xnor U446 (N_446,In_401,In_109);
and U447 (N_447,In_1106,N_298);
nor U448 (N_448,N_279,N_207);
and U449 (N_449,In_1178,In_203);
and U450 (N_450,In_937,In_906);
nand U451 (N_451,In_1016,In_198);
xor U452 (N_452,In_1327,In_1291);
or U453 (N_453,In_225,In_437);
nand U454 (N_454,In_574,In_1414);
nor U455 (N_455,In_1219,N_281);
xnor U456 (N_456,In_1304,In_733);
nor U457 (N_457,N_58,In_1329);
and U458 (N_458,In_1238,In_1125);
and U459 (N_459,In_988,In_1338);
or U460 (N_460,In_1410,N_189);
or U461 (N_461,N_171,In_663);
or U462 (N_462,In_1281,In_824);
nand U463 (N_463,In_800,In_757);
nand U464 (N_464,In_344,In_603);
xor U465 (N_465,In_1031,In_860);
nor U466 (N_466,In_1194,N_10);
nand U467 (N_467,In_1294,In_1350);
xnor U468 (N_468,In_1236,N_112);
nor U469 (N_469,In_68,N_370);
nand U470 (N_470,In_1367,In_1046);
xnor U471 (N_471,N_187,In_619);
xor U472 (N_472,In_1265,N_192);
xor U473 (N_473,In_852,In_469);
and U474 (N_474,In_154,N_268);
nand U475 (N_475,In_1423,In_427);
and U476 (N_476,In_1258,In_356);
xnor U477 (N_477,N_320,In_840);
or U478 (N_478,In_583,In_480);
and U479 (N_479,In_436,N_366);
and U480 (N_480,In_52,In_1196);
nor U481 (N_481,In_514,In_616);
and U482 (N_482,N_149,In_156);
or U483 (N_483,In_1169,In_1431);
and U484 (N_484,In_79,In_108);
nor U485 (N_485,In_832,N_153);
and U486 (N_486,N_333,In_1437);
or U487 (N_487,In_28,In_626);
nand U488 (N_488,In_940,In_431);
nand U489 (N_489,In_888,In_281);
and U490 (N_490,N_287,In_853);
nor U491 (N_491,In_375,In_826);
nand U492 (N_492,In_112,In_113);
nor U493 (N_493,N_138,N_355);
nor U494 (N_494,In_152,In_301);
xnor U495 (N_495,In_1012,In_987);
xnor U496 (N_496,N_198,N_339);
or U497 (N_497,N_253,In_350);
nor U498 (N_498,In_1084,In_793);
nor U499 (N_499,In_1208,In_1320);
or U500 (N_500,N_419,In_248);
or U501 (N_501,N_219,N_103);
nand U502 (N_502,N_422,N_341);
xnor U503 (N_503,N_398,In_378);
or U504 (N_504,In_726,N_427);
xnor U505 (N_505,In_44,N_452);
and U506 (N_506,In_734,N_469);
and U507 (N_507,In_1449,N_238);
and U508 (N_508,In_682,N_343);
and U509 (N_509,N_479,N_33);
xor U510 (N_510,N_247,N_276);
nand U511 (N_511,In_415,N_373);
xnor U512 (N_512,In_123,In_1360);
xor U513 (N_513,In_481,N_496);
nand U514 (N_514,In_1045,In_857);
nand U515 (N_515,In_518,In_808);
xnor U516 (N_516,In_418,N_179);
nand U517 (N_517,In_498,In_639);
nand U518 (N_518,N_289,In_886);
nor U519 (N_519,N_170,In_207);
nand U520 (N_520,In_199,In_501);
and U521 (N_521,In_550,N_412);
or U522 (N_522,In_1382,In_564);
and U523 (N_523,N_383,In_1292);
nor U524 (N_524,In_391,In_319);
nand U525 (N_525,N_337,In_270);
and U526 (N_526,N_463,N_116);
and U527 (N_527,In_1211,N_354);
xnor U528 (N_528,N_100,In_1485);
xnor U529 (N_529,In_1206,In_764);
xor U530 (N_530,In_1483,N_232);
xor U531 (N_531,N_215,N_88);
nor U532 (N_532,In_1379,In_272);
and U533 (N_533,In_320,In_208);
or U534 (N_534,N_303,N_386);
nand U535 (N_535,In_638,N_234);
and U536 (N_536,In_1341,N_377);
nor U537 (N_537,N_143,N_384);
nor U538 (N_538,N_399,N_126);
or U539 (N_539,N_37,N_217);
nor U540 (N_540,In_1102,In_1430);
and U541 (N_541,In_1348,In_1166);
nor U542 (N_542,N_371,N_302);
nand U543 (N_543,In_47,N_329);
or U544 (N_544,N_379,N_150);
xnor U545 (N_545,N_125,In_759);
nor U546 (N_546,In_1205,In_539);
nor U547 (N_547,In_307,N_437);
xor U548 (N_548,N_161,In_1319);
nor U549 (N_549,N_440,N_300);
xor U550 (N_550,In_279,N_259);
and U551 (N_551,In_812,In_1316);
and U552 (N_552,In_540,N_325);
nor U553 (N_553,N_471,In_381);
or U554 (N_554,N_292,In_1408);
nand U555 (N_555,N_223,In_326);
nor U556 (N_556,In_1465,In_1176);
nor U557 (N_557,In_256,In_535);
xnor U558 (N_558,In_1285,In_667);
nand U559 (N_559,N_257,N_2);
nand U560 (N_560,In_803,In_332);
nor U561 (N_561,N_488,In_212);
or U562 (N_562,In_528,In_1065);
nor U563 (N_563,N_128,N_50);
and U564 (N_564,In_1468,In_1471);
xnor U565 (N_565,In_999,N_96);
and U566 (N_566,In_941,In_903);
xnor U567 (N_567,In_1134,In_634);
xnor U568 (N_568,N_243,In_1099);
and U569 (N_569,In_829,N_353);
xnor U570 (N_570,N_394,In_1253);
xnor U571 (N_571,N_75,In_222);
nand U572 (N_572,N_401,In_934);
nand U573 (N_573,N_406,N_486);
nor U574 (N_574,N_291,In_1421);
nor U575 (N_575,In_1191,In_1040);
or U576 (N_576,In_672,In_77);
nor U577 (N_577,In_1230,N_97);
nor U578 (N_578,N_40,In_884);
or U579 (N_579,In_445,In_75);
nor U580 (N_580,In_1036,In_489);
or U581 (N_581,N_260,In_1302);
nand U582 (N_582,In_182,N_244);
or U583 (N_583,In_1118,N_123);
xnor U584 (N_584,N_470,N_148);
nor U585 (N_585,In_1039,In_1420);
xor U586 (N_586,In_463,In_537);
and U587 (N_587,In_641,In_1419);
or U588 (N_588,In_103,In_355);
and U589 (N_589,In_187,N_158);
nand U590 (N_590,N_361,In_524);
xor U591 (N_591,N_218,In_305);
nor U592 (N_592,N_262,In_181);
nor U593 (N_593,In_339,In_1216);
nand U594 (N_594,N_136,In_1417);
nor U595 (N_595,In_277,In_1378);
nand U596 (N_596,In_730,N_344);
nand U597 (N_597,In_1014,N_381);
or U598 (N_598,In_863,In_872);
nor U599 (N_599,N_326,N_462);
xor U600 (N_600,In_1363,In_457);
or U601 (N_601,In_917,In_11);
xnor U602 (N_602,N_425,In_1244);
and U603 (N_603,In_798,In_1295);
xor U604 (N_604,In_4,In_1148);
xnor U605 (N_605,In_959,N_282);
and U606 (N_606,In_115,N_107);
nor U607 (N_607,N_474,In_865);
nor U608 (N_608,In_351,In_146);
or U609 (N_609,In_1305,N_80);
and U610 (N_610,In_817,In_242);
or U611 (N_611,N_417,In_472);
and U612 (N_612,In_206,N_142);
and U613 (N_613,In_333,N_449);
or U614 (N_614,In_1440,N_205);
nand U615 (N_615,In_1425,N_335);
nand U616 (N_616,In_722,N_174);
nor U617 (N_617,N_71,N_489);
or U618 (N_618,In_922,N_178);
and U619 (N_619,N_334,In_695);
nor U620 (N_620,N_327,N_340);
nor U621 (N_621,In_120,In_1433);
nor U622 (N_622,In_650,N_348);
and U623 (N_623,In_948,In_933);
nor U624 (N_624,N_299,In_392);
nand U625 (N_625,In_1264,In_189);
and U626 (N_626,N_68,In_321);
xor U627 (N_627,N_85,N_332);
nor U628 (N_628,N_593,N_457);
nand U629 (N_629,In_1047,In_57);
nand U630 (N_630,In_311,N_318);
nand U631 (N_631,In_499,N_512);
xnor U632 (N_632,N_408,N_211);
nor U633 (N_633,In_1489,In_1112);
or U634 (N_634,In_644,N_342);
or U635 (N_635,In_1375,N_616);
nand U636 (N_636,In_220,N_517);
nor U637 (N_637,N_579,N_129);
nor U638 (N_638,In_1187,In_697);
nand U639 (N_639,In_230,In_1115);
xnor U640 (N_640,In_1242,In_645);
or U641 (N_641,N_94,N_364);
nor U642 (N_642,In_656,In_1486);
nor U643 (N_643,In_604,In_637);
or U644 (N_644,In_1042,In_118);
nor U645 (N_645,In_1478,In_276);
nor U646 (N_646,N_532,In_1019);
xor U647 (N_647,N_494,N_585);
or U648 (N_648,N_275,N_589);
nor U649 (N_649,In_1111,N_16);
xor U650 (N_650,N_530,N_559);
and U651 (N_651,In_565,N_133);
nor U652 (N_652,In_1263,N_317);
xor U653 (N_653,N_439,In_484);
and U654 (N_654,In_76,In_259);
nand U655 (N_655,In_786,In_951);
or U656 (N_656,In_38,In_1069);
nor U657 (N_657,In_1498,In_671);
or U658 (N_658,N_545,N_375);
and U659 (N_659,In_185,N_294);
and U660 (N_660,N_212,N_248);
nand U661 (N_661,N_468,N_441);
nand U662 (N_662,In_1426,N_426);
or U663 (N_663,In_139,In_1369);
xor U664 (N_664,In_503,In_854);
and U665 (N_665,In_982,N_435);
xor U666 (N_666,In_994,N_546);
and U667 (N_667,In_167,N_272);
nand U668 (N_668,N_249,In_149);
and U669 (N_669,N_507,In_1467);
nand U670 (N_670,N_542,N_273);
nand U671 (N_671,N_239,N_429);
nor U672 (N_672,In_5,In_1366);
xnor U673 (N_673,In_1243,In_1358);
nor U674 (N_674,In_1010,N_256);
xor U675 (N_675,In_1076,N_519);
nor U676 (N_676,In_1011,In_1310);
xnor U677 (N_677,In_265,In_85);
and U678 (N_678,In_1455,In_1171);
nor U679 (N_679,N_152,N_573);
nor U680 (N_680,N_388,N_135);
nor U681 (N_681,In_40,In_504);
nand U682 (N_682,N_622,N_310);
xnor U683 (N_683,N_413,In_531);
or U684 (N_684,In_449,N_623);
and U685 (N_685,N_430,In_386);
and U686 (N_686,N_534,N_78);
nand U687 (N_687,N_448,In_1146);
xnor U688 (N_688,N_250,In_529);
and U689 (N_689,N_506,N_359);
nor U690 (N_690,In_1037,In_1459);
xnor U691 (N_691,N_606,N_528);
nor U692 (N_692,In_946,In_1345);
nand U693 (N_693,In_494,In_66);
xnor U694 (N_694,In_1168,In_290);
and U695 (N_695,In_567,In_130);
nor U696 (N_696,In_1339,In_176);
and U697 (N_697,N_34,In_755);
nand U698 (N_698,In_1298,In_428);
or U699 (N_699,N_24,In_300);
xor U700 (N_700,In_1004,N_264);
xor U701 (N_701,N_159,N_403);
nand U702 (N_702,N_395,In_701);
nand U703 (N_703,In_838,N_587);
or U704 (N_704,In_192,In_1340);
nand U705 (N_705,N_600,N_183);
xor U706 (N_706,In_224,N_500);
or U707 (N_707,N_563,In_915);
nand U708 (N_708,In_282,N_531);
or U709 (N_709,In_334,N_351);
or U710 (N_710,In_566,N_290);
nand U711 (N_711,N_0,N_511);
or U712 (N_712,N_186,In_1460);
nand U713 (N_713,N_544,N_131);
nand U714 (N_714,In_1306,N_524);
nand U715 (N_715,In_93,N_378);
or U716 (N_716,In_1003,In_1300);
nand U717 (N_717,In_1043,N_502);
xor U718 (N_718,In_827,N_580);
and U719 (N_719,N_434,In_597);
and U720 (N_720,In_330,N_328);
and U721 (N_721,In_1179,In_1356);
xor U722 (N_722,N_108,In_287);
nand U723 (N_723,In_1087,In_304);
and U724 (N_724,N_387,In_67);
nor U725 (N_725,N_321,N_495);
nor U726 (N_726,N_543,In_1237);
xor U727 (N_727,In_1409,N_491);
xor U728 (N_728,N_409,N_541);
xnor U729 (N_729,In_1083,N_132);
nand U730 (N_730,N_231,In_559);
nor U731 (N_731,N_330,In_412);
nand U732 (N_732,In_165,In_1048);
xnor U733 (N_733,N_581,N_267);
nor U734 (N_734,In_965,In_1092);
and U735 (N_735,In_312,N_614);
or U736 (N_736,In_1346,N_229);
nor U737 (N_737,N_173,N_410);
xor U738 (N_738,N_41,N_389);
nand U739 (N_739,In_22,In_1121);
xnor U740 (N_740,In_72,N_608);
and U741 (N_741,In_314,In_1260);
xnor U742 (N_742,In_1185,N_492);
nand U743 (N_743,In_869,In_862);
and U744 (N_744,In_1269,N_122);
nor U745 (N_745,In_101,N_367);
xnor U746 (N_746,In_411,N_609);
or U747 (N_747,N_521,In_1381);
and U748 (N_748,In_1145,In_191);
xor U749 (N_749,N_121,N_604);
nand U750 (N_750,In_1385,N_52);
nand U751 (N_751,N_691,In_519);
or U752 (N_752,In_725,In_724);
xor U753 (N_753,N_445,N_251);
or U754 (N_754,N_637,In_1307);
or U755 (N_755,N_450,In_1018);
nand U756 (N_756,In_921,N_571);
nand U757 (N_757,N_438,N_312);
xnor U758 (N_758,In_421,N_65);
xnor U759 (N_759,N_447,N_115);
and U760 (N_760,N_558,In_773);
nor U761 (N_761,In_1197,N_687);
nand U762 (N_762,In_609,In_91);
and U763 (N_763,In_388,In_373);
and U764 (N_764,N_619,In_70);
nor U765 (N_765,In_497,N_526);
and U766 (N_766,In_124,In_791);
or U767 (N_767,N_336,N_513);
or U768 (N_768,In_691,In_324);
xnor U769 (N_769,In_1131,In_253);
or U770 (N_770,N_7,N_363);
xor U771 (N_771,In_747,N_188);
or U772 (N_772,In_84,N_631);
xor U773 (N_773,N_590,In_670);
xor U774 (N_774,In_702,N_660);
and U775 (N_775,In_204,N_548);
or U776 (N_776,N_642,N_659);
nand U777 (N_777,In_459,N_576);
xnor U778 (N_778,In_1407,In_200);
nor U779 (N_779,In_1480,In_1321);
or U780 (N_780,In_849,In_80);
nand U781 (N_781,N_635,N_725);
nand U782 (N_782,N_301,N_311);
or U783 (N_783,In_1282,N_533);
and U784 (N_784,In_608,N_501);
nand U785 (N_785,N_677,N_191);
and U786 (N_786,In_771,N_482);
or U787 (N_787,In_1136,N_681);
and U788 (N_788,In_1373,In_216);
nand U789 (N_789,N_671,N_700);
xnor U790 (N_790,N_368,In_947);
or U791 (N_791,In_323,N_498);
nand U792 (N_792,In_58,N_689);
or U793 (N_793,N_701,N_433);
nand U794 (N_794,N_101,N_520);
and U795 (N_795,In_796,N_358);
or U796 (N_796,In_1223,In_1443);
and U797 (N_797,In_376,N_114);
nand U798 (N_798,In_153,N_737);
nor U799 (N_799,N_560,In_1251);
or U800 (N_800,N_416,In_160);
xor U801 (N_801,N_627,In_289);
or U802 (N_802,N_638,N_306);
nor U803 (N_803,N_391,N_607);
xnor U804 (N_804,N_666,N_216);
or U805 (N_805,In_327,In_960);
nand U806 (N_806,In_526,N_602);
nor U807 (N_807,In_897,In_1173);
nor U808 (N_808,In_409,N_538);
xnor U809 (N_809,N_644,In_1413);
nand U810 (N_810,In_818,In_1163);
nand U811 (N_811,N_567,N_263);
xor U812 (N_812,N_688,In_171);
xnor U813 (N_813,In_240,N_663);
nor U814 (N_814,In_647,In_792);
or U815 (N_815,In_923,N_568);
nor U816 (N_816,N_628,N_345);
nor U817 (N_817,N_346,N_246);
or U818 (N_818,In_492,In_1020);
and U819 (N_819,In_633,N_713);
nor U820 (N_820,In_1128,N_586);
or U821 (N_821,N_683,In_443);
nand U822 (N_822,N_293,N_45);
nand U823 (N_823,N_295,N_485);
nor U824 (N_824,In_432,N_547);
and U825 (N_825,N_679,In_195);
nand U826 (N_826,In_527,N_432);
and U827 (N_827,In_686,In_166);
nand U828 (N_828,N_396,In_669);
and U829 (N_829,N_655,N_451);
xor U830 (N_830,In_983,N_286);
nand U831 (N_831,N_424,N_732);
or U832 (N_832,N_331,In_348);
and U833 (N_833,In_1386,In_635);
xnor U834 (N_834,N_658,In_926);
nor U835 (N_835,N_119,In_1324);
xor U836 (N_836,N_540,In_1204);
and U837 (N_837,N_583,In_599);
and U838 (N_838,In_1453,In_723);
nand U839 (N_839,In_455,N_649);
xnor U840 (N_840,N_698,In_385);
and U841 (N_841,N_380,N_514);
and U842 (N_842,In_99,N_473);
nor U843 (N_843,In_23,N_552);
or U844 (N_844,N_106,In_1061);
xnor U845 (N_845,N_747,N_453);
and U846 (N_846,N_708,N_421);
nand U847 (N_847,N_601,N_551);
xnor U848 (N_848,N_536,N_621);
or U849 (N_849,In_8,N_305);
xnor U850 (N_850,In_630,In_196);
nor U851 (N_851,N_1,In_648);
and U852 (N_852,In_1266,N_618);
and U853 (N_853,N_39,N_400);
nor U854 (N_854,In_362,In_1152);
or U855 (N_855,In_26,In_453);
nor U856 (N_856,N_557,N_748);
or U857 (N_857,In_1062,In_717);
xor U858 (N_858,N_228,N_487);
and U859 (N_859,In_655,N_407);
and U860 (N_860,In_973,In_63);
nor U861 (N_861,N_484,N_455);
nand U862 (N_862,N_503,In_684);
or U863 (N_863,N_316,N_645);
and U864 (N_864,In_592,N_744);
nand U865 (N_865,In_1495,N_712);
nand U866 (N_866,N_307,In_688);
nand U867 (N_867,In_1353,In_1101);
or U868 (N_868,In_1380,N_73);
and U869 (N_869,N_475,N_261);
and U870 (N_870,N_226,In_15);
nand U871 (N_871,N_525,N_443);
and U872 (N_872,In_229,N_582);
nand U873 (N_873,N_592,In_1117);
and U874 (N_874,N_704,N_431);
nand U875 (N_875,N_554,N_861);
xnor U876 (N_876,In_221,N_594);
and U877 (N_877,N_869,N_796);
and U878 (N_878,In_555,N_778);
or U879 (N_879,N_781,N_674);
or U880 (N_880,N_662,In_1086);
xnor U881 (N_881,N_18,N_564);
and U882 (N_882,N_117,In_1212);
xnor U883 (N_883,In_1325,N_629);
nor U884 (N_884,N_770,N_680);
xnor U885 (N_885,In_775,N_813);
xor U886 (N_886,N_118,N_369);
or U887 (N_887,N_814,N_783);
or U888 (N_888,In_21,In_368);
nor U889 (N_889,In_105,N_352);
nand U890 (N_890,In_508,N_739);
xnor U891 (N_891,N_868,In_868);
nor U892 (N_892,N_442,N_772);
or U893 (N_893,N_35,In_61);
nand U894 (N_894,In_1344,In_1314);
and U895 (N_895,N_633,N_848);
xor U896 (N_896,N_717,N_753);
nand U897 (N_897,N_319,In_464);
nor U898 (N_898,N_865,In_700);
and U899 (N_899,N_740,In_794);
or U900 (N_900,N_497,In_471);
nor U901 (N_901,In_1404,N_365);
and U902 (N_902,N_699,In_1002);
nor U903 (N_903,N_867,N_873);
or U904 (N_904,In_1210,N_376);
nor U905 (N_905,N_789,In_876);
nand U906 (N_906,N_411,N_574);
xnor U907 (N_907,N_709,In_1334);
nor U908 (N_908,N_745,In_673);
xnor U909 (N_909,N_743,N_347);
nand U910 (N_910,N_795,N_860);
xor U911 (N_911,N_181,In_246);
or U912 (N_912,N_610,In_39);
and U913 (N_913,In_1278,N_812);
nor U914 (N_914,In_900,N_695);
nand U915 (N_915,N_518,N_837);
nand U916 (N_916,In_309,In_49);
or U917 (N_917,N_707,In_227);
nor U918 (N_918,In_338,N_436);
and U919 (N_919,In_461,In_150);
xnor U920 (N_920,In_1088,In_439);
xnor U921 (N_921,N_620,N_799);
nand U922 (N_922,In_533,In_125);
nor U923 (N_923,In_569,In_928);
xor U924 (N_924,N_596,In_19);
and U925 (N_925,In_517,N_784);
xor U926 (N_926,N_849,N_270);
nand U927 (N_927,In_666,N_62);
or U928 (N_928,N_810,In_315);
or U929 (N_929,In_407,N_338);
xor U930 (N_930,N_750,In_1342);
nor U931 (N_931,N_779,In_929);
nand U932 (N_932,In_642,N_832);
nand U933 (N_933,In_1174,In_1183);
nor U934 (N_934,N_672,N_800);
or U935 (N_935,In_322,In_1023);
or U936 (N_936,In_1309,N_749);
nor U937 (N_937,N_850,In_140);
nand U938 (N_938,N_357,N_639);
nand U939 (N_939,In_157,N_209);
xnor U940 (N_940,N_856,N_817);
xor U941 (N_941,N_350,N_838);
nor U942 (N_942,In_1141,N_141);
nand U943 (N_943,N_575,N_458);
and U944 (N_944,In_1030,N_527);
nand U945 (N_945,In_715,N_402);
nor U946 (N_946,N_842,In_1034);
or U947 (N_947,In_1418,N_405);
or U948 (N_948,In_1286,N_791);
nor U949 (N_949,In_316,In_134);
nand U950 (N_950,N_761,In_893);
and U951 (N_951,N_640,N_798);
xor U952 (N_952,N_803,N_323);
and U953 (N_953,In_55,N_818);
and U954 (N_954,N_561,In_358);
and U955 (N_955,In_969,N_28);
and U956 (N_956,In_1,N_390);
nand U957 (N_957,N_522,In_1120);
xor U958 (N_958,N_265,N_420);
xor U959 (N_959,N_721,N_591);
nor U960 (N_960,In_1193,N_308);
xor U961 (N_961,In_1328,N_767);
and U962 (N_962,In_1399,In_197);
nor U963 (N_963,In_423,In_743);
nor U964 (N_964,In_822,N_769);
xor U965 (N_965,N_309,N_650);
and U966 (N_966,N_555,In_211);
nor U967 (N_967,In_1077,N_288);
or U968 (N_968,In_972,N_742);
xnor U969 (N_969,N_70,N_428);
or U970 (N_970,N_210,In_1432);
nor U971 (N_971,N_509,In_1396);
nor U972 (N_972,In_382,In_848);
and U973 (N_973,N_692,N_752);
nand U974 (N_974,In_95,N_356);
nand U975 (N_975,In_444,In_842);
xnor U976 (N_976,In_611,N_611);
or U977 (N_977,N_615,N_139);
nor U978 (N_978,N_197,N_827);
xnor U979 (N_979,In_500,In_460);
nand U980 (N_980,In_395,N_858);
nor U981 (N_981,N_613,N_483);
xor U982 (N_982,In_173,N_176);
and U983 (N_983,N_846,N_565);
nor U984 (N_984,N_252,N_647);
nor U985 (N_985,N_572,N_870);
or U986 (N_986,In_447,In_163);
nor U987 (N_987,N_185,In_783);
and U988 (N_988,N_382,N_780);
nor U989 (N_989,N_626,In_62);
nor U990 (N_990,N_459,In_1276);
xnor U991 (N_991,N_313,N_166);
or U992 (N_992,N_874,N_194);
nor U993 (N_993,N_535,N_236);
and U994 (N_994,N_277,N_617);
or U995 (N_995,N_834,In_1357);
xor U996 (N_996,In_1090,N_505);
or U997 (N_997,N_751,N_757);
or U998 (N_998,In_989,In_1150);
or U999 (N_999,N_819,N_661);
nor U1000 (N_1000,N_808,N_756);
xor U1001 (N_1001,N_144,N_254);
nand U1002 (N_1002,N_902,In_1397);
nand U1003 (N_1003,N_634,N_667);
nand U1004 (N_1004,N_678,In_664);
or U1005 (N_1005,In_135,N_941);
xnor U1006 (N_1006,N_738,N_948);
xor U1007 (N_1007,N_632,N_797);
xnor U1008 (N_1008,N_910,N_372);
or U1009 (N_1009,In_549,N_146);
xor U1010 (N_1010,In_889,In_981);
or U1011 (N_1011,In_575,N_971);
or U1012 (N_1012,N_771,In_1249);
nand U1013 (N_1013,N_630,N_969);
nor U1014 (N_1014,N_516,N_765);
xor U1015 (N_1015,N_599,N_929);
and U1016 (N_1016,In_1057,N_714);
nor U1017 (N_1017,In_296,In_1257);
and U1018 (N_1018,In_121,N_914);
xor U1019 (N_1019,N_982,In_2);
or U1020 (N_1020,N_225,In_1164);
nand U1021 (N_1021,In_1412,N_888);
and U1022 (N_1022,N_99,N_776);
or U1023 (N_1023,N_879,N_786);
xor U1024 (N_1024,N_964,N_831);
or U1025 (N_1025,N_731,N_959);
or U1026 (N_1026,In_252,N_675);
and U1027 (N_1027,N_863,In_846);
or U1028 (N_1028,N_127,N_283);
xor U1029 (N_1029,N_917,N_905);
and U1030 (N_1030,N_840,N_957);
nor U1031 (N_1031,N_966,N_852);
and U1032 (N_1032,N_939,N_673);
nand U1033 (N_1033,N_156,In_1234);
and U1034 (N_1034,N_668,N_996);
xor U1035 (N_1035,In_1322,N_807);
nand U1036 (N_1036,N_423,N_539);
nand U1037 (N_1037,In_693,N_711);
xnor U1038 (N_1038,N_465,N_624);
nor U1039 (N_1039,N_898,N_537);
nor U1040 (N_1040,N_9,N_792);
xnor U1041 (N_1041,In_438,In_572);
and U1042 (N_1042,N_880,In_1390);
and U1043 (N_1043,N_651,N_901);
and U1044 (N_1044,N_862,N_762);
or U1045 (N_1045,N_991,N_360);
xnor U1046 (N_1046,N_774,In_1192);
and U1047 (N_1047,N_790,N_973);
or U1048 (N_1048,In_654,N_999);
or U1049 (N_1049,N_493,In_1492);
xor U1050 (N_1050,N_515,N_954);
nand U1051 (N_1051,N_990,N_923);
nand U1052 (N_1052,N_918,N_903);
nand U1053 (N_1053,N_933,N_900);
xnor U1054 (N_1054,N_899,N_913);
and U1055 (N_1055,N_643,N_706);
xnor U1056 (N_1056,In_1107,In_706);
and U1057 (N_1057,In_346,N_764);
nand U1058 (N_1058,N_919,N_788);
or U1059 (N_1059,N_490,N_461);
nand U1060 (N_1060,In_493,N_993);
nor U1061 (N_1061,N_773,N_851);
nand U1062 (N_1062,N_956,N_464);
or U1063 (N_1063,N_978,N_255);
nor U1064 (N_1064,N_975,In_417);
xnor U1065 (N_1065,N_895,In_1008);
nand U1066 (N_1066,N_570,In_1000);
nand U1067 (N_1067,In_377,In_104);
xor U1068 (N_1068,In_1376,N_904);
nor U1069 (N_1069,N_777,N_909);
xor U1070 (N_1070,In_502,In_342);
nor U1071 (N_1071,In_151,N_648);
nor U1072 (N_1072,In_1135,In_184);
and U1073 (N_1073,In_357,N_997);
xnor U1074 (N_1074,N_972,In_257);
xnor U1075 (N_1075,N_577,N_657);
nor U1076 (N_1076,N_718,N_726);
or U1077 (N_1077,In_1140,N_735);
xor U1078 (N_1078,In_1398,N_603);
xnor U1079 (N_1079,N_829,In_509);
xor U1080 (N_1080,N_988,N_896);
and U1081 (N_1081,N_578,N_598);
xnor U1082 (N_1082,N_208,N_877);
nor U1083 (N_1083,N_987,N_883);
xor U1084 (N_1084,In_78,N_924);
nor U1085 (N_1085,N_754,N_927);
or U1086 (N_1086,N_758,N_864);
xor U1087 (N_1087,N_550,N_801);
and U1088 (N_1088,N_477,In_680);
and U1089 (N_1089,N_857,In_1352);
nand U1090 (N_1090,N_26,N_926);
nor U1091 (N_1091,N_835,N_705);
nor U1092 (N_1092,In_1439,In_367);
nor U1093 (N_1093,N_221,N_885);
nand U1094 (N_1094,N_947,N_682);
xor U1095 (N_1095,In_856,N_670);
nand U1096 (N_1096,N_595,N_654);
xor U1097 (N_1097,In_1095,N_976);
nand U1098 (N_1098,N_190,In_81);
xnor U1099 (N_1099,N_392,N_523);
and U1100 (N_1100,N_845,N_816);
nand U1101 (N_1101,In_1053,In_766);
or U1102 (N_1102,In_908,N_84);
nor U1103 (N_1103,N_953,N_921);
xnor U1104 (N_1104,N_943,N_815);
xnor U1105 (N_1105,N_958,N_979);
or U1106 (N_1106,N_824,N_893);
nand U1107 (N_1107,N_809,N_562);
or U1108 (N_1108,In_1072,N_936);
nor U1109 (N_1109,N_952,N_349);
or U1110 (N_1110,N_951,N_727);
xor U1111 (N_1111,N_984,In_957);
nand U1112 (N_1112,In_403,N_508);
nand U1113 (N_1113,In_576,In_25);
nand U1114 (N_1114,N_641,N_274);
nor U1115 (N_1115,N_76,N_805);
and U1116 (N_1116,N_878,N_266);
and U1117 (N_1117,N_793,In_365);
or U1118 (N_1118,N_734,In_1082);
xor U1119 (N_1119,N_970,N_890);
nand U1120 (N_1120,N_931,N_855);
nand U1121 (N_1121,N_324,In_1073);
nor U1122 (N_1122,N_859,N_168);
or U1123 (N_1123,In_16,N_703);
nand U1124 (N_1124,In_1262,In_624);
or U1125 (N_1125,N_887,N_1055);
nand U1126 (N_1126,N_625,N_605);
or U1127 (N_1127,N_998,N_1075);
or U1128 (N_1128,N_1090,N_258);
xnor U1129 (N_1129,N_928,N_1068);
and U1130 (N_1130,N_992,In_1308);
and U1131 (N_1131,N_1029,N_822);
nand U1132 (N_1132,N_720,N_1020);
xnor U1133 (N_1133,N_823,In_35);
and U1134 (N_1134,N_1094,N_804);
nor U1135 (N_1135,N_529,N_697);
nand U1136 (N_1136,In_387,In_1103);
and U1137 (N_1137,N_588,In_174);
xor U1138 (N_1138,N_944,N_1017);
nand U1139 (N_1139,N_315,N_397);
nand U1140 (N_1140,N_955,N_1058);
xnor U1141 (N_1141,N_1043,N_162);
xnor U1142 (N_1142,N_684,N_907);
xor U1143 (N_1143,N_646,N_866);
nor U1144 (N_1144,N_980,N_1087);
xor U1145 (N_1145,N_930,In_729);
nand U1146 (N_1146,N_1082,In_899);
nand U1147 (N_1147,In_651,In_1330);
or U1148 (N_1148,In_1299,N_1023);
and U1149 (N_1149,N_871,N_1019);
nand U1150 (N_1150,N_994,In_347);
nand U1151 (N_1151,N_1105,N_960);
xnor U1152 (N_1152,N_1070,N_665);
nand U1153 (N_1153,In_561,N_690);
nor U1154 (N_1154,N_911,N_1121);
and U1155 (N_1155,N_710,N_724);
and U1156 (N_1156,N_686,N_1064);
and U1157 (N_1157,N_1048,N_995);
nand U1158 (N_1158,In_405,N_1106);
and U1159 (N_1159,N_932,N_1050);
nand U1160 (N_1160,N_1080,In_1207);
nand U1161 (N_1161,N_1030,N_1014);
xor U1162 (N_1162,N_1040,N_1027);
or U1163 (N_1163,N_768,N_280);
nor U1164 (N_1164,N_1083,N_1053);
and U1165 (N_1165,N_715,N_1051);
nand U1166 (N_1166,N_460,In_1268);
nor U1167 (N_1167,N_478,N_967);
and U1168 (N_1168,In_297,N_61);
and U1169 (N_1169,N_1114,N_1028);
nor U1170 (N_1170,N_1099,N_843);
and U1171 (N_1171,N_418,In_1132);
nand U1172 (N_1172,N_1092,N_636);
nor U1173 (N_1173,N_1041,N_1011);
and U1174 (N_1174,N_1012,In_1395);
xnor U1175 (N_1175,N_787,In_275);
xnor U1176 (N_1176,N_949,N_481);
or U1177 (N_1177,In_1104,In_1217);
or U1178 (N_1178,N_1010,In_209);
and U1179 (N_1179,N_1031,In_538);
nand U1180 (N_1180,N_1108,N_1085);
nor U1181 (N_1181,N_1061,N_1066);
xnor U1182 (N_1182,N_763,N_556);
and U1183 (N_1183,N_977,In_1105);
nor U1184 (N_1184,N_584,N_986);
nand U1185 (N_1185,N_1037,N_1021);
xor U1186 (N_1186,N_1084,N_1044);
nand U1187 (N_1187,N_825,N_882);
and U1188 (N_1188,N_1104,N_847);
nand U1189 (N_1189,In_1068,N_612);
or U1190 (N_1190,In_1275,N_746);
nor U1191 (N_1191,N_1096,N_794);
or U1192 (N_1192,N_1078,N_811);
or U1193 (N_1193,In_1006,N_504);
xor U1194 (N_1194,In_482,N_1091);
or U1195 (N_1195,N_922,N_897);
and U1196 (N_1196,N_1042,N_730);
xor U1197 (N_1197,N_1086,N_1047);
nand U1198 (N_1198,N_456,In_1472);
xor U1199 (N_1199,In_1493,N_985);
nor U1200 (N_1200,In_1411,N_1002);
and U1201 (N_1201,N_881,N_1118);
xor U1202 (N_1202,N_962,N_1013);
nand U1203 (N_1203,In_433,N_946);
or U1204 (N_1204,N_466,N_1074);
or U1205 (N_1205,N_472,In_34);
xnor U1206 (N_1206,In_186,N_886);
xnor U1207 (N_1207,N_1117,N_1122);
nand U1208 (N_1208,N_1008,N_820);
or U1209 (N_1209,N_1006,N_741);
nor U1210 (N_1210,N_664,N_1034);
xor U1211 (N_1211,N_569,N_652);
nor U1212 (N_1212,N_937,N_826);
nand U1213 (N_1213,N_42,In_426);
nand U1214 (N_1214,N_653,N_908);
nand U1215 (N_1215,In_30,N_1124);
nand U1216 (N_1216,N_1001,N_669);
nor U1217 (N_1217,N_1073,N_785);
nand U1218 (N_1218,N_1000,N_1054);
and U1219 (N_1219,N_467,N_963);
nand U1220 (N_1220,N_989,N_676);
nor U1221 (N_1221,N_875,In_223);
nand U1222 (N_1222,In_1317,N_1113);
and U1223 (N_1223,In_719,N_782);
and U1224 (N_1224,In_568,In_110);
and U1225 (N_1225,In_369,N_1004);
or U1226 (N_1226,N_1093,In_678);
nand U1227 (N_1227,In_1267,N_1052);
or U1228 (N_1228,N_1123,In_545);
or U1229 (N_1229,N_802,N_1089);
nand U1230 (N_1230,N_1079,N_833);
nand U1231 (N_1231,In_1044,N_1100);
and U1232 (N_1232,N_476,N_1063);
nor U1233 (N_1233,In_328,N_722);
and U1234 (N_1234,In_374,N_1072);
or U1235 (N_1235,N_1067,N_981);
nor U1236 (N_1236,N_1069,N_1024);
or U1237 (N_1237,N_1077,In_964);
and U1238 (N_1238,N_1049,N_385);
and U1239 (N_1239,N_1076,N_716);
xor U1240 (N_1240,In_37,N_889);
or U1241 (N_1241,N_1038,N_1045);
xor U1242 (N_1242,N_915,In_692);
xnor U1243 (N_1243,N_566,N_841);
xnor U1244 (N_1244,N_728,N_1065);
nor U1245 (N_1245,N_836,N_1103);
or U1246 (N_1246,N_775,N_1060);
nand U1247 (N_1247,N_925,N_844);
or U1248 (N_1248,N_1025,N_912);
or U1249 (N_1249,N_894,N_968);
nor U1250 (N_1250,N_965,N_1137);
nand U1251 (N_1251,N_206,N_1232);
or U1252 (N_1252,N_1172,N_1156);
nand U1253 (N_1253,N_480,N_1214);
xnor U1254 (N_1254,In_1496,In_442);
or U1255 (N_1255,N_1005,N_1225);
or U1256 (N_1256,N_1224,N_1120);
and U1257 (N_1257,N_1217,N_1178);
and U1258 (N_1258,N_1227,N_940);
nand U1259 (N_1259,N_454,N_1159);
nor U1260 (N_1260,N_1180,N_1187);
nor U1261 (N_1261,N_1242,N_1155);
or U1262 (N_1262,N_1109,N_872);
or U1263 (N_1263,N_1240,N_733);
xor U1264 (N_1264,N_1228,In_974);
nand U1265 (N_1265,N_1184,N_755);
and U1266 (N_1266,N_1164,N_1160);
nand U1267 (N_1267,N_44,N_1152);
and U1268 (N_1268,N_1098,N_1143);
and U1269 (N_1269,N_1195,N_974);
and U1270 (N_1270,N_1125,N_1165);
or U1271 (N_1271,N_1233,N_1131);
nor U1272 (N_1272,N_1059,N_1204);
nor U1273 (N_1273,In_979,N_1241);
nand U1274 (N_1274,N_1230,N_1111);
or U1275 (N_1275,N_1150,N_884);
and U1276 (N_1276,N_759,N_892);
and U1277 (N_1277,N_961,In_653);
or U1278 (N_1278,N_1141,N_1088);
xor U1279 (N_1279,N_766,N_1161);
nor U1280 (N_1280,N_1062,N_1200);
and U1281 (N_1281,N_1036,In_510);
or U1282 (N_1282,N_1209,N_1162);
xor U1283 (N_1283,N_1144,N_1212);
xnor U1284 (N_1284,N_1033,N_278);
nand U1285 (N_1285,N_1147,N_1221);
nand U1286 (N_1286,N_1127,N_1208);
nand U1287 (N_1287,N_1193,In_588);
xnor U1288 (N_1288,N_414,N_1151);
nor U1289 (N_1289,N_1138,N_821);
xor U1290 (N_1290,N_1003,N_1201);
nor U1291 (N_1291,N_839,N_876);
nand U1292 (N_1292,N_1133,N_1173);
and U1293 (N_1293,N_1149,N_1186);
xnor U1294 (N_1294,N_1198,N_1231);
nor U1295 (N_1295,In_782,N_719);
nand U1296 (N_1296,N_444,N_1207);
and U1297 (N_1297,N_1203,N_1007);
and U1298 (N_1298,N_3,N_702);
or U1299 (N_1299,N_656,N_983);
or U1300 (N_1300,N_1057,N_1192);
nor U1301 (N_1301,N_1166,N_1039);
and U1302 (N_1302,N_1163,N_1026);
and U1303 (N_1303,N_1206,N_1119);
nand U1304 (N_1304,N_1148,N_1247);
nor U1305 (N_1305,N_1095,N_510);
and U1306 (N_1306,In_1022,In_1221);
nand U1307 (N_1307,N_1115,N_201);
nand U1308 (N_1308,N_1239,N_1130);
nand U1309 (N_1309,N_1210,N_1226);
and U1310 (N_1310,N_1181,N_1154);
or U1311 (N_1311,N_1216,N_446);
and U1312 (N_1312,In_487,N_1035);
and U1313 (N_1313,N_853,N_1188);
or U1314 (N_1314,N_1213,N_1220);
nor U1315 (N_1315,N_1249,N_1135);
nand U1316 (N_1316,In_306,N_1171);
and U1317 (N_1317,N_1190,N_1248);
or U1318 (N_1318,N_685,N_830);
or U1319 (N_1319,N_854,N_1128);
or U1320 (N_1320,N_1146,N_271);
or U1321 (N_1321,N_1245,N_1046);
nor U1322 (N_1322,N_935,N_942);
xor U1323 (N_1323,N_1129,N_1246);
nand U1324 (N_1324,N_404,N_597);
xor U1325 (N_1325,N_200,N_1022);
and U1326 (N_1326,N_696,N_828);
xor U1327 (N_1327,In_1075,N_1177);
nor U1328 (N_1328,N_169,N_1015);
nor U1329 (N_1329,N_393,N_1158);
nor U1330 (N_1330,N_499,N_1153);
nor U1331 (N_1331,N_1142,N_693);
xnor U1332 (N_1332,N_1179,N_1139);
nand U1333 (N_1333,N_1205,N_723);
xnor U1334 (N_1334,N_945,N_694);
nor U1335 (N_1335,N_1116,N_1244);
nand U1336 (N_1336,In_813,N_1071);
nand U1337 (N_1337,N_934,N_1032);
nand U1338 (N_1338,N_1194,N_1140);
xor U1339 (N_1339,N_1134,N_1219);
nor U1340 (N_1340,N_1218,N_950);
nand U1341 (N_1341,N_109,N_415);
nand U1342 (N_1342,N_54,N_920);
nand U1343 (N_1343,N_1234,N_1056);
or U1344 (N_1344,N_1211,N_1189);
xor U1345 (N_1345,N_1238,In_175);
xor U1346 (N_1346,N_1175,N_1112);
or U1347 (N_1347,N_1235,N_1183);
and U1348 (N_1348,N_137,N_1222);
nor U1349 (N_1349,N_1174,N_1236);
nor U1350 (N_1350,N_163,N_134);
and U1351 (N_1351,N_1169,N_155);
nand U1352 (N_1352,N_1237,N_1243);
nor U1353 (N_1353,N_1107,N_1182);
nand U1354 (N_1354,N_1199,N_1110);
xor U1355 (N_1355,N_1168,N_891);
xnor U1356 (N_1356,N_1223,N_1009);
xor U1357 (N_1357,N_1126,N_760);
nor U1358 (N_1358,N_1185,N_1196);
xnor U1359 (N_1359,N_906,N_1229);
nor U1360 (N_1360,N_1197,N_1157);
nor U1361 (N_1361,N_1101,N_1170);
xor U1362 (N_1362,N_1145,N_806);
xnor U1363 (N_1363,N_1097,N_729);
or U1364 (N_1364,N_736,N_1215);
and U1365 (N_1365,N_77,N_1191);
and U1366 (N_1366,In_1159,N_916);
nand U1367 (N_1367,N_1136,N_1016);
or U1368 (N_1368,N_63,In_1435);
nor U1369 (N_1369,N_1202,N_1176);
or U1370 (N_1370,N_549,N_1081);
nor U1371 (N_1371,N_1167,N_938);
nor U1372 (N_1372,In_451,N_553);
or U1373 (N_1373,N_1132,N_1102);
nand U1374 (N_1374,In_657,N_1018);
xnor U1375 (N_1375,N_1314,N_1290);
or U1376 (N_1376,N_1251,N_1301);
or U1377 (N_1377,N_1258,N_1260);
nor U1378 (N_1378,N_1341,N_1266);
xor U1379 (N_1379,N_1317,N_1313);
and U1380 (N_1380,N_1287,N_1362);
nor U1381 (N_1381,N_1322,N_1330);
nand U1382 (N_1382,N_1271,N_1368);
or U1383 (N_1383,N_1336,N_1295);
or U1384 (N_1384,N_1340,N_1324);
or U1385 (N_1385,N_1250,N_1361);
nand U1386 (N_1386,N_1355,N_1357);
xnor U1387 (N_1387,N_1373,N_1310);
xor U1388 (N_1388,N_1289,N_1252);
xnor U1389 (N_1389,N_1305,N_1363);
nor U1390 (N_1390,N_1291,N_1306);
and U1391 (N_1391,N_1293,N_1263);
nand U1392 (N_1392,N_1369,N_1300);
and U1393 (N_1393,N_1273,N_1269);
xnor U1394 (N_1394,N_1356,N_1344);
nand U1395 (N_1395,N_1337,N_1288);
or U1396 (N_1396,N_1339,N_1277);
or U1397 (N_1397,N_1284,N_1304);
nand U1398 (N_1398,N_1358,N_1346);
or U1399 (N_1399,N_1272,N_1267);
nand U1400 (N_1400,N_1285,N_1281);
nor U1401 (N_1401,N_1335,N_1255);
xor U1402 (N_1402,N_1275,N_1351);
nor U1403 (N_1403,N_1366,N_1360);
nand U1404 (N_1404,N_1352,N_1350);
and U1405 (N_1405,N_1326,N_1307);
xor U1406 (N_1406,N_1321,N_1354);
and U1407 (N_1407,N_1270,N_1365);
nand U1408 (N_1408,N_1256,N_1332);
or U1409 (N_1409,N_1253,N_1342);
or U1410 (N_1410,N_1283,N_1348);
or U1411 (N_1411,N_1282,N_1264);
xnor U1412 (N_1412,N_1334,N_1359);
or U1413 (N_1413,N_1353,N_1372);
or U1414 (N_1414,N_1308,N_1328);
xor U1415 (N_1415,N_1349,N_1338);
nor U1416 (N_1416,N_1323,N_1364);
nand U1417 (N_1417,N_1261,N_1371);
and U1418 (N_1418,N_1311,N_1312);
nor U1419 (N_1419,N_1319,N_1367);
and U1420 (N_1420,N_1297,N_1278);
nor U1421 (N_1421,N_1296,N_1265);
nor U1422 (N_1422,N_1294,N_1327);
xnor U1423 (N_1423,N_1318,N_1333);
and U1424 (N_1424,N_1370,N_1262);
xnor U1425 (N_1425,N_1316,N_1302);
or U1426 (N_1426,N_1320,N_1257);
xor U1427 (N_1427,N_1280,N_1309);
and U1428 (N_1428,N_1259,N_1343);
and U1429 (N_1429,N_1298,N_1329);
nor U1430 (N_1430,N_1347,N_1274);
nor U1431 (N_1431,N_1292,N_1299);
xor U1432 (N_1432,N_1279,N_1315);
nand U1433 (N_1433,N_1331,N_1268);
nand U1434 (N_1434,N_1325,N_1286);
nor U1435 (N_1435,N_1345,N_1374);
or U1436 (N_1436,N_1303,N_1276);
nand U1437 (N_1437,N_1254,N_1266);
nor U1438 (N_1438,N_1285,N_1261);
xnor U1439 (N_1439,N_1260,N_1256);
xor U1440 (N_1440,N_1332,N_1262);
nand U1441 (N_1441,N_1255,N_1276);
or U1442 (N_1442,N_1356,N_1318);
nand U1443 (N_1443,N_1359,N_1297);
or U1444 (N_1444,N_1362,N_1288);
nand U1445 (N_1445,N_1340,N_1317);
xnor U1446 (N_1446,N_1301,N_1297);
and U1447 (N_1447,N_1338,N_1322);
and U1448 (N_1448,N_1353,N_1336);
nand U1449 (N_1449,N_1263,N_1336);
and U1450 (N_1450,N_1255,N_1313);
nor U1451 (N_1451,N_1354,N_1348);
nand U1452 (N_1452,N_1266,N_1256);
and U1453 (N_1453,N_1303,N_1350);
and U1454 (N_1454,N_1303,N_1353);
xor U1455 (N_1455,N_1351,N_1326);
and U1456 (N_1456,N_1360,N_1277);
nor U1457 (N_1457,N_1289,N_1301);
and U1458 (N_1458,N_1285,N_1335);
and U1459 (N_1459,N_1312,N_1268);
nand U1460 (N_1460,N_1273,N_1354);
or U1461 (N_1461,N_1314,N_1288);
nand U1462 (N_1462,N_1268,N_1328);
or U1463 (N_1463,N_1353,N_1300);
nor U1464 (N_1464,N_1288,N_1342);
and U1465 (N_1465,N_1347,N_1301);
and U1466 (N_1466,N_1281,N_1365);
or U1467 (N_1467,N_1266,N_1292);
and U1468 (N_1468,N_1367,N_1304);
nor U1469 (N_1469,N_1279,N_1282);
nor U1470 (N_1470,N_1268,N_1360);
nor U1471 (N_1471,N_1339,N_1303);
nand U1472 (N_1472,N_1350,N_1322);
or U1473 (N_1473,N_1270,N_1250);
nor U1474 (N_1474,N_1293,N_1266);
nor U1475 (N_1475,N_1349,N_1329);
and U1476 (N_1476,N_1317,N_1311);
or U1477 (N_1477,N_1282,N_1353);
and U1478 (N_1478,N_1275,N_1346);
or U1479 (N_1479,N_1347,N_1288);
nor U1480 (N_1480,N_1267,N_1359);
and U1481 (N_1481,N_1301,N_1258);
nor U1482 (N_1482,N_1283,N_1274);
or U1483 (N_1483,N_1297,N_1286);
nand U1484 (N_1484,N_1263,N_1353);
xor U1485 (N_1485,N_1327,N_1363);
nor U1486 (N_1486,N_1311,N_1290);
xnor U1487 (N_1487,N_1301,N_1332);
xnor U1488 (N_1488,N_1357,N_1294);
and U1489 (N_1489,N_1350,N_1282);
and U1490 (N_1490,N_1261,N_1361);
nand U1491 (N_1491,N_1364,N_1328);
nand U1492 (N_1492,N_1344,N_1278);
xnor U1493 (N_1493,N_1264,N_1343);
nor U1494 (N_1494,N_1357,N_1273);
nor U1495 (N_1495,N_1295,N_1283);
nor U1496 (N_1496,N_1307,N_1289);
xor U1497 (N_1497,N_1257,N_1271);
nand U1498 (N_1498,N_1356,N_1371);
or U1499 (N_1499,N_1374,N_1335);
xnor U1500 (N_1500,N_1404,N_1435);
or U1501 (N_1501,N_1499,N_1440);
nand U1502 (N_1502,N_1421,N_1429);
and U1503 (N_1503,N_1385,N_1476);
and U1504 (N_1504,N_1459,N_1383);
or U1505 (N_1505,N_1452,N_1494);
and U1506 (N_1506,N_1451,N_1464);
or U1507 (N_1507,N_1434,N_1406);
nand U1508 (N_1508,N_1405,N_1481);
xor U1509 (N_1509,N_1461,N_1477);
or U1510 (N_1510,N_1387,N_1415);
and U1511 (N_1511,N_1399,N_1475);
nand U1512 (N_1512,N_1381,N_1472);
or U1513 (N_1513,N_1417,N_1473);
xnor U1514 (N_1514,N_1482,N_1426);
nand U1515 (N_1515,N_1409,N_1431);
and U1516 (N_1516,N_1388,N_1444);
nor U1517 (N_1517,N_1397,N_1398);
or U1518 (N_1518,N_1389,N_1490);
or U1519 (N_1519,N_1391,N_1375);
and U1520 (N_1520,N_1438,N_1402);
nand U1521 (N_1521,N_1420,N_1376);
xnor U1522 (N_1522,N_1423,N_1463);
xnor U1523 (N_1523,N_1489,N_1449);
or U1524 (N_1524,N_1395,N_1380);
xnor U1525 (N_1525,N_1474,N_1418);
and U1526 (N_1526,N_1419,N_1469);
xnor U1527 (N_1527,N_1446,N_1487);
xnor U1528 (N_1528,N_1460,N_1400);
or U1529 (N_1529,N_1416,N_1479);
or U1530 (N_1530,N_1448,N_1379);
xnor U1531 (N_1531,N_1447,N_1491);
xor U1532 (N_1532,N_1443,N_1483);
nor U1533 (N_1533,N_1401,N_1478);
nor U1534 (N_1534,N_1467,N_1394);
nand U1535 (N_1535,N_1378,N_1462);
nor U1536 (N_1536,N_1377,N_1488);
nand U1537 (N_1537,N_1485,N_1410);
nor U1538 (N_1538,N_1384,N_1386);
nand U1539 (N_1539,N_1442,N_1437);
or U1540 (N_1540,N_1439,N_1496);
or U1541 (N_1541,N_1393,N_1430);
nor U1542 (N_1542,N_1484,N_1411);
nand U1543 (N_1543,N_1392,N_1468);
or U1544 (N_1544,N_1441,N_1454);
or U1545 (N_1545,N_1436,N_1413);
nor U1546 (N_1546,N_1453,N_1407);
and U1547 (N_1547,N_1465,N_1382);
xor U1548 (N_1548,N_1412,N_1433);
and U1549 (N_1549,N_1471,N_1456);
and U1550 (N_1550,N_1408,N_1396);
and U1551 (N_1551,N_1428,N_1470);
xor U1552 (N_1552,N_1390,N_1498);
or U1553 (N_1553,N_1450,N_1492);
nand U1554 (N_1554,N_1455,N_1457);
nand U1555 (N_1555,N_1458,N_1403);
and U1556 (N_1556,N_1480,N_1493);
or U1557 (N_1557,N_1422,N_1427);
nand U1558 (N_1558,N_1432,N_1497);
xnor U1559 (N_1559,N_1445,N_1425);
xor U1560 (N_1560,N_1414,N_1486);
or U1561 (N_1561,N_1424,N_1466);
xnor U1562 (N_1562,N_1495,N_1385);
nand U1563 (N_1563,N_1380,N_1496);
and U1564 (N_1564,N_1419,N_1375);
xor U1565 (N_1565,N_1423,N_1398);
and U1566 (N_1566,N_1452,N_1489);
and U1567 (N_1567,N_1399,N_1404);
or U1568 (N_1568,N_1435,N_1430);
and U1569 (N_1569,N_1375,N_1386);
or U1570 (N_1570,N_1398,N_1411);
xor U1571 (N_1571,N_1394,N_1465);
nand U1572 (N_1572,N_1499,N_1485);
or U1573 (N_1573,N_1434,N_1492);
xor U1574 (N_1574,N_1392,N_1485);
xor U1575 (N_1575,N_1423,N_1417);
and U1576 (N_1576,N_1475,N_1388);
and U1577 (N_1577,N_1457,N_1448);
nand U1578 (N_1578,N_1441,N_1472);
and U1579 (N_1579,N_1405,N_1382);
nand U1580 (N_1580,N_1404,N_1391);
xnor U1581 (N_1581,N_1473,N_1389);
nand U1582 (N_1582,N_1404,N_1437);
nand U1583 (N_1583,N_1462,N_1456);
and U1584 (N_1584,N_1444,N_1396);
or U1585 (N_1585,N_1493,N_1410);
nand U1586 (N_1586,N_1416,N_1459);
and U1587 (N_1587,N_1403,N_1478);
and U1588 (N_1588,N_1480,N_1485);
nand U1589 (N_1589,N_1453,N_1414);
xnor U1590 (N_1590,N_1471,N_1484);
or U1591 (N_1591,N_1440,N_1426);
xnor U1592 (N_1592,N_1482,N_1461);
and U1593 (N_1593,N_1435,N_1386);
nor U1594 (N_1594,N_1410,N_1384);
nor U1595 (N_1595,N_1441,N_1395);
xnor U1596 (N_1596,N_1463,N_1413);
nor U1597 (N_1597,N_1393,N_1464);
or U1598 (N_1598,N_1420,N_1435);
nor U1599 (N_1599,N_1494,N_1417);
and U1600 (N_1600,N_1474,N_1416);
and U1601 (N_1601,N_1486,N_1450);
or U1602 (N_1602,N_1465,N_1412);
nor U1603 (N_1603,N_1447,N_1478);
and U1604 (N_1604,N_1406,N_1449);
nor U1605 (N_1605,N_1400,N_1496);
or U1606 (N_1606,N_1484,N_1439);
xnor U1607 (N_1607,N_1472,N_1404);
nand U1608 (N_1608,N_1494,N_1469);
xor U1609 (N_1609,N_1400,N_1375);
and U1610 (N_1610,N_1453,N_1419);
or U1611 (N_1611,N_1458,N_1425);
nor U1612 (N_1612,N_1381,N_1486);
nor U1613 (N_1613,N_1384,N_1480);
xor U1614 (N_1614,N_1401,N_1485);
or U1615 (N_1615,N_1445,N_1415);
nor U1616 (N_1616,N_1454,N_1492);
or U1617 (N_1617,N_1457,N_1386);
or U1618 (N_1618,N_1485,N_1455);
nor U1619 (N_1619,N_1457,N_1379);
nand U1620 (N_1620,N_1448,N_1402);
nand U1621 (N_1621,N_1425,N_1396);
nand U1622 (N_1622,N_1443,N_1385);
xor U1623 (N_1623,N_1394,N_1488);
nand U1624 (N_1624,N_1458,N_1422);
nand U1625 (N_1625,N_1500,N_1543);
nand U1626 (N_1626,N_1524,N_1506);
nand U1627 (N_1627,N_1502,N_1539);
and U1628 (N_1628,N_1589,N_1578);
or U1629 (N_1629,N_1536,N_1556);
or U1630 (N_1630,N_1549,N_1602);
nor U1631 (N_1631,N_1504,N_1604);
and U1632 (N_1632,N_1587,N_1620);
or U1633 (N_1633,N_1547,N_1530);
nand U1634 (N_1634,N_1513,N_1515);
xor U1635 (N_1635,N_1619,N_1510);
nand U1636 (N_1636,N_1550,N_1548);
xor U1637 (N_1637,N_1605,N_1512);
and U1638 (N_1638,N_1600,N_1566);
and U1639 (N_1639,N_1580,N_1579);
nand U1640 (N_1640,N_1565,N_1557);
xnor U1641 (N_1641,N_1526,N_1518);
nand U1642 (N_1642,N_1595,N_1607);
and U1643 (N_1643,N_1535,N_1583);
or U1644 (N_1644,N_1603,N_1614);
and U1645 (N_1645,N_1599,N_1581);
xnor U1646 (N_1646,N_1597,N_1590);
or U1647 (N_1647,N_1501,N_1591);
or U1648 (N_1648,N_1570,N_1517);
and U1649 (N_1649,N_1527,N_1559);
and U1650 (N_1650,N_1552,N_1584);
nor U1651 (N_1651,N_1577,N_1511);
or U1652 (N_1652,N_1521,N_1563);
or U1653 (N_1653,N_1612,N_1516);
and U1654 (N_1654,N_1594,N_1574);
xor U1655 (N_1655,N_1528,N_1615);
or U1656 (N_1656,N_1613,N_1610);
nor U1657 (N_1657,N_1542,N_1534);
nand U1658 (N_1658,N_1598,N_1553);
nand U1659 (N_1659,N_1609,N_1537);
or U1660 (N_1660,N_1541,N_1617);
xnor U1661 (N_1661,N_1573,N_1571);
and U1662 (N_1662,N_1585,N_1569);
and U1663 (N_1663,N_1520,N_1608);
nor U1664 (N_1664,N_1564,N_1514);
nor U1665 (N_1665,N_1588,N_1544);
nor U1666 (N_1666,N_1561,N_1558);
nand U1667 (N_1667,N_1616,N_1508);
xor U1668 (N_1668,N_1505,N_1555);
nor U1669 (N_1669,N_1601,N_1575);
or U1670 (N_1670,N_1560,N_1531);
xnor U1671 (N_1671,N_1586,N_1519);
nor U1672 (N_1672,N_1545,N_1532);
or U1673 (N_1673,N_1624,N_1606);
nand U1674 (N_1674,N_1592,N_1509);
or U1675 (N_1675,N_1568,N_1503);
or U1676 (N_1676,N_1533,N_1622);
xor U1677 (N_1677,N_1593,N_1522);
or U1678 (N_1678,N_1618,N_1562);
xor U1679 (N_1679,N_1540,N_1611);
or U1680 (N_1680,N_1567,N_1551);
and U1681 (N_1681,N_1572,N_1523);
xnor U1682 (N_1682,N_1546,N_1507);
xor U1683 (N_1683,N_1554,N_1576);
or U1684 (N_1684,N_1596,N_1538);
nor U1685 (N_1685,N_1621,N_1582);
nand U1686 (N_1686,N_1623,N_1529);
xor U1687 (N_1687,N_1525,N_1544);
or U1688 (N_1688,N_1540,N_1518);
xor U1689 (N_1689,N_1567,N_1531);
nor U1690 (N_1690,N_1581,N_1547);
nand U1691 (N_1691,N_1515,N_1578);
xnor U1692 (N_1692,N_1585,N_1525);
nand U1693 (N_1693,N_1584,N_1542);
nand U1694 (N_1694,N_1540,N_1562);
nand U1695 (N_1695,N_1502,N_1596);
and U1696 (N_1696,N_1552,N_1619);
nor U1697 (N_1697,N_1614,N_1619);
nand U1698 (N_1698,N_1579,N_1607);
and U1699 (N_1699,N_1552,N_1603);
or U1700 (N_1700,N_1593,N_1534);
or U1701 (N_1701,N_1502,N_1517);
nor U1702 (N_1702,N_1520,N_1515);
and U1703 (N_1703,N_1608,N_1551);
or U1704 (N_1704,N_1623,N_1614);
xnor U1705 (N_1705,N_1603,N_1543);
xnor U1706 (N_1706,N_1622,N_1526);
and U1707 (N_1707,N_1581,N_1574);
xnor U1708 (N_1708,N_1586,N_1526);
and U1709 (N_1709,N_1504,N_1568);
nor U1710 (N_1710,N_1591,N_1507);
or U1711 (N_1711,N_1608,N_1581);
and U1712 (N_1712,N_1540,N_1598);
nand U1713 (N_1713,N_1541,N_1608);
and U1714 (N_1714,N_1555,N_1534);
nand U1715 (N_1715,N_1529,N_1613);
nor U1716 (N_1716,N_1508,N_1563);
and U1717 (N_1717,N_1614,N_1515);
nand U1718 (N_1718,N_1583,N_1569);
or U1719 (N_1719,N_1583,N_1529);
or U1720 (N_1720,N_1591,N_1553);
nand U1721 (N_1721,N_1524,N_1549);
and U1722 (N_1722,N_1589,N_1558);
nand U1723 (N_1723,N_1546,N_1591);
nor U1724 (N_1724,N_1515,N_1548);
nand U1725 (N_1725,N_1619,N_1610);
nand U1726 (N_1726,N_1622,N_1507);
or U1727 (N_1727,N_1564,N_1531);
nor U1728 (N_1728,N_1550,N_1604);
nor U1729 (N_1729,N_1583,N_1505);
xor U1730 (N_1730,N_1561,N_1552);
or U1731 (N_1731,N_1596,N_1566);
or U1732 (N_1732,N_1609,N_1585);
and U1733 (N_1733,N_1574,N_1588);
nor U1734 (N_1734,N_1624,N_1534);
and U1735 (N_1735,N_1612,N_1518);
or U1736 (N_1736,N_1523,N_1510);
or U1737 (N_1737,N_1500,N_1541);
nor U1738 (N_1738,N_1612,N_1527);
nor U1739 (N_1739,N_1561,N_1555);
nor U1740 (N_1740,N_1509,N_1516);
xor U1741 (N_1741,N_1622,N_1590);
or U1742 (N_1742,N_1548,N_1595);
and U1743 (N_1743,N_1605,N_1619);
nand U1744 (N_1744,N_1506,N_1501);
and U1745 (N_1745,N_1576,N_1569);
or U1746 (N_1746,N_1595,N_1589);
xor U1747 (N_1747,N_1600,N_1539);
and U1748 (N_1748,N_1531,N_1528);
nor U1749 (N_1749,N_1579,N_1624);
or U1750 (N_1750,N_1654,N_1658);
and U1751 (N_1751,N_1647,N_1635);
and U1752 (N_1752,N_1703,N_1721);
nand U1753 (N_1753,N_1699,N_1695);
nand U1754 (N_1754,N_1670,N_1636);
or U1755 (N_1755,N_1637,N_1710);
and U1756 (N_1756,N_1681,N_1645);
xor U1757 (N_1757,N_1687,N_1631);
or U1758 (N_1758,N_1718,N_1702);
xnor U1759 (N_1759,N_1665,N_1685);
xor U1760 (N_1760,N_1648,N_1630);
nand U1761 (N_1761,N_1692,N_1732);
nand U1762 (N_1762,N_1736,N_1734);
nand U1763 (N_1763,N_1727,N_1694);
nand U1764 (N_1764,N_1634,N_1707);
and U1765 (N_1765,N_1684,N_1726);
or U1766 (N_1766,N_1678,N_1671);
xor U1767 (N_1767,N_1741,N_1642);
nor U1768 (N_1768,N_1659,N_1646);
or U1769 (N_1769,N_1705,N_1704);
and U1770 (N_1770,N_1673,N_1632);
and U1771 (N_1771,N_1663,N_1728);
nand U1772 (N_1772,N_1643,N_1679);
nand U1773 (N_1773,N_1698,N_1650);
nor U1774 (N_1774,N_1667,N_1666);
and U1775 (N_1775,N_1745,N_1733);
or U1776 (N_1776,N_1655,N_1723);
and U1777 (N_1777,N_1700,N_1706);
or U1778 (N_1778,N_1696,N_1625);
nand U1779 (N_1779,N_1713,N_1656);
or U1780 (N_1780,N_1664,N_1724);
or U1781 (N_1781,N_1709,N_1649);
nor U1782 (N_1782,N_1715,N_1627);
nor U1783 (N_1783,N_1740,N_1653);
nand U1784 (N_1784,N_1638,N_1693);
or U1785 (N_1785,N_1746,N_1725);
nand U1786 (N_1786,N_1662,N_1714);
or U1787 (N_1787,N_1735,N_1719);
and U1788 (N_1788,N_1629,N_1668);
xnor U1789 (N_1789,N_1747,N_1744);
nand U1790 (N_1790,N_1651,N_1657);
xor U1791 (N_1791,N_1691,N_1628);
and U1792 (N_1792,N_1738,N_1730);
or U1793 (N_1793,N_1672,N_1712);
nor U1794 (N_1794,N_1748,N_1644);
and U1795 (N_1795,N_1689,N_1669);
nor U1796 (N_1796,N_1697,N_1660);
and U1797 (N_1797,N_1717,N_1640);
xor U1798 (N_1798,N_1682,N_1677);
or U1799 (N_1799,N_1626,N_1641);
nand U1800 (N_1800,N_1729,N_1674);
nor U1801 (N_1801,N_1675,N_1639);
nor U1802 (N_1802,N_1742,N_1676);
or U1803 (N_1803,N_1690,N_1711);
and U1804 (N_1804,N_1686,N_1652);
or U1805 (N_1805,N_1683,N_1749);
nor U1806 (N_1806,N_1720,N_1708);
nand U1807 (N_1807,N_1722,N_1737);
and U1808 (N_1808,N_1743,N_1701);
and U1809 (N_1809,N_1661,N_1716);
nor U1810 (N_1810,N_1680,N_1731);
nand U1811 (N_1811,N_1688,N_1633);
xnor U1812 (N_1812,N_1739,N_1635);
and U1813 (N_1813,N_1745,N_1741);
and U1814 (N_1814,N_1666,N_1726);
xnor U1815 (N_1815,N_1636,N_1745);
xor U1816 (N_1816,N_1658,N_1650);
and U1817 (N_1817,N_1720,N_1745);
nor U1818 (N_1818,N_1748,N_1719);
xor U1819 (N_1819,N_1632,N_1694);
nand U1820 (N_1820,N_1671,N_1688);
and U1821 (N_1821,N_1731,N_1702);
nor U1822 (N_1822,N_1645,N_1676);
nand U1823 (N_1823,N_1708,N_1683);
nand U1824 (N_1824,N_1731,N_1740);
nor U1825 (N_1825,N_1668,N_1709);
and U1826 (N_1826,N_1697,N_1670);
nand U1827 (N_1827,N_1721,N_1661);
nand U1828 (N_1828,N_1749,N_1719);
nor U1829 (N_1829,N_1636,N_1736);
and U1830 (N_1830,N_1625,N_1652);
xor U1831 (N_1831,N_1731,N_1715);
or U1832 (N_1832,N_1705,N_1727);
or U1833 (N_1833,N_1643,N_1690);
nor U1834 (N_1834,N_1734,N_1691);
or U1835 (N_1835,N_1667,N_1716);
xnor U1836 (N_1836,N_1728,N_1707);
nor U1837 (N_1837,N_1684,N_1625);
nand U1838 (N_1838,N_1748,N_1639);
xnor U1839 (N_1839,N_1730,N_1652);
or U1840 (N_1840,N_1721,N_1630);
or U1841 (N_1841,N_1710,N_1719);
nand U1842 (N_1842,N_1680,N_1692);
or U1843 (N_1843,N_1744,N_1651);
xnor U1844 (N_1844,N_1690,N_1640);
or U1845 (N_1845,N_1647,N_1650);
and U1846 (N_1846,N_1652,N_1737);
nor U1847 (N_1847,N_1693,N_1659);
xor U1848 (N_1848,N_1641,N_1740);
xor U1849 (N_1849,N_1625,N_1632);
nor U1850 (N_1850,N_1721,N_1729);
nor U1851 (N_1851,N_1669,N_1726);
nor U1852 (N_1852,N_1673,N_1701);
nand U1853 (N_1853,N_1749,N_1627);
xor U1854 (N_1854,N_1720,N_1716);
nor U1855 (N_1855,N_1722,N_1683);
and U1856 (N_1856,N_1653,N_1716);
or U1857 (N_1857,N_1695,N_1749);
nand U1858 (N_1858,N_1706,N_1696);
nor U1859 (N_1859,N_1699,N_1627);
nor U1860 (N_1860,N_1693,N_1725);
nand U1861 (N_1861,N_1732,N_1678);
xnor U1862 (N_1862,N_1728,N_1730);
or U1863 (N_1863,N_1636,N_1629);
or U1864 (N_1864,N_1663,N_1681);
nand U1865 (N_1865,N_1733,N_1692);
xor U1866 (N_1866,N_1717,N_1678);
or U1867 (N_1867,N_1736,N_1730);
nor U1868 (N_1868,N_1741,N_1701);
xor U1869 (N_1869,N_1665,N_1651);
nor U1870 (N_1870,N_1746,N_1650);
and U1871 (N_1871,N_1745,N_1663);
nor U1872 (N_1872,N_1713,N_1714);
and U1873 (N_1873,N_1662,N_1694);
or U1874 (N_1874,N_1705,N_1745);
or U1875 (N_1875,N_1830,N_1869);
and U1876 (N_1876,N_1751,N_1765);
or U1877 (N_1877,N_1782,N_1847);
nand U1878 (N_1878,N_1865,N_1760);
nand U1879 (N_1879,N_1810,N_1799);
or U1880 (N_1880,N_1779,N_1833);
or U1881 (N_1881,N_1796,N_1805);
or U1882 (N_1882,N_1825,N_1866);
and U1883 (N_1883,N_1831,N_1789);
nand U1884 (N_1884,N_1856,N_1823);
nor U1885 (N_1885,N_1843,N_1758);
or U1886 (N_1886,N_1838,N_1834);
or U1887 (N_1887,N_1874,N_1812);
nor U1888 (N_1888,N_1794,N_1761);
or U1889 (N_1889,N_1815,N_1802);
nor U1890 (N_1890,N_1801,N_1762);
or U1891 (N_1891,N_1839,N_1787);
and U1892 (N_1892,N_1840,N_1793);
nor U1893 (N_1893,N_1767,N_1819);
and U1894 (N_1894,N_1848,N_1868);
or U1895 (N_1895,N_1862,N_1807);
or U1896 (N_1896,N_1826,N_1818);
nor U1897 (N_1897,N_1870,N_1808);
and U1898 (N_1898,N_1858,N_1770);
and U1899 (N_1899,N_1871,N_1853);
nor U1900 (N_1900,N_1849,N_1776);
or U1901 (N_1901,N_1841,N_1809);
and U1902 (N_1902,N_1851,N_1777);
xnor U1903 (N_1903,N_1864,N_1790);
or U1904 (N_1904,N_1757,N_1814);
nand U1905 (N_1905,N_1752,N_1828);
and U1906 (N_1906,N_1832,N_1791);
nand U1907 (N_1907,N_1768,N_1804);
or U1908 (N_1908,N_1854,N_1803);
nand U1909 (N_1909,N_1764,N_1795);
nand U1910 (N_1910,N_1785,N_1786);
nor U1911 (N_1911,N_1873,N_1763);
or U1912 (N_1912,N_1775,N_1829);
nor U1913 (N_1913,N_1778,N_1771);
xnor U1914 (N_1914,N_1850,N_1855);
or U1915 (N_1915,N_1846,N_1759);
nand U1916 (N_1916,N_1822,N_1813);
nand U1917 (N_1917,N_1769,N_1750);
nand U1918 (N_1918,N_1788,N_1844);
xnor U1919 (N_1919,N_1772,N_1753);
or U1920 (N_1920,N_1859,N_1792);
and U1921 (N_1921,N_1800,N_1811);
or U1922 (N_1922,N_1766,N_1852);
nand U1923 (N_1923,N_1842,N_1816);
or U1924 (N_1924,N_1827,N_1845);
and U1925 (N_1925,N_1784,N_1835);
and U1926 (N_1926,N_1867,N_1797);
and U1927 (N_1927,N_1754,N_1817);
xor U1928 (N_1928,N_1824,N_1872);
or U1929 (N_1929,N_1774,N_1781);
or U1930 (N_1930,N_1806,N_1798);
or U1931 (N_1931,N_1780,N_1836);
and U1932 (N_1932,N_1773,N_1756);
xor U1933 (N_1933,N_1821,N_1860);
and U1934 (N_1934,N_1837,N_1783);
nor U1935 (N_1935,N_1861,N_1863);
and U1936 (N_1936,N_1857,N_1820);
or U1937 (N_1937,N_1755,N_1805);
and U1938 (N_1938,N_1769,N_1854);
and U1939 (N_1939,N_1804,N_1773);
or U1940 (N_1940,N_1786,N_1873);
xnor U1941 (N_1941,N_1767,N_1803);
or U1942 (N_1942,N_1828,N_1855);
xnor U1943 (N_1943,N_1795,N_1866);
nor U1944 (N_1944,N_1865,N_1832);
nand U1945 (N_1945,N_1769,N_1788);
or U1946 (N_1946,N_1861,N_1810);
xor U1947 (N_1947,N_1853,N_1765);
or U1948 (N_1948,N_1865,N_1786);
nand U1949 (N_1949,N_1846,N_1795);
or U1950 (N_1950,N_1830,N_1808);
and U1951 (N_1951,N_1849,N_1786);
nor U1952 (N_1952,N_1820,N_1804);
xnor U1953 (N_1953,N_1786,N_1819);
and U1954 (N_1954,N_1791,N_1765);
xor U1955 (N_1955,N_1785,N_1766);
nand U1956 (N_1956,N_1757,N_1817);
nand U1957 (N_1957,N_1846,N_1780);
nand U1958 (N_1958,N_1798,N_1791);
nor U1959 (N_1959,N_1756,N_1779);
xnor U1960 (N_1960,N_1754,N_1794);
or U1961 (N_1961,N_1761,N_1802);
and U1962 (N_1962,N_1834,N_1773);
xor U1963 (N_1963,N_1830,N_1819);
and U1964 (N_1964,N_1759,N_1868);
nor U1965 (N_1965,N_1863,N_1832);
nor U1966 (N_1966,N_1826,N_1834);
nor U1967 (N_1967,N_1839,N_1772);
nor U1968 (N_1968,N_1869,N_1866);
nor U1969 (N_1969,N_1799,N_1831);
and U1970 (N_1970,N_1767,N_1810);
or U1971 (N_1971,N_1838,N_1754);
nand U1972 (N_1972,N_1828,N_1771);
nand U1973 (N_1973,N_1808,N_1860);
xor U1974 (N_1974,N_1806,N_1791);
nand U1975 (N_1975,N_1774,N_1822);
and U1976 (N_1976,N_1753,N_1805);
nand U1977 (N_1977,N_1818,N_1849);
and U1978 (N_1978,N_1761,N_1756);
or U1979 (N_1979,N_1762,N_1779);
or U1980 (N_1980,N_1838,N_1866);
nand U1981 (N_1981,N_1754,N_1789);
and U1982 (N_1982,N_1835,N_1774);
xnor U1983 (N_1983,N_1837,N_1864);
or U1984 (N_1984,N_1821,N_1816);
and U1985 (N_1985,N_1762,N_1792);
or U1986 (N_1986,N_1778,N_1847);
and U1987 (N_1987,N_1861,N_1829);
or U1988 (N_1988,N_1761,N_1790);
or U1989 (N_1989,N_1823,N_1855);
xor U1990 (N_1990,N_1808,N_1837);
and U1991 (N_1991,N_1802,N_1841);
xor U1992 (N_1992,N_1856,N_1783);
or U1993 (N_1993,N_1869,N_1782);
xor U1994 (N_1994,N_1832,N_1803);
and U1995 (N_1995,N_1809,N_1839);
and U1996 (N_1996,N_1763,N_1791);
or U1997 (N_1997,N_1804,N_1774);
nand U1998 (N_1998,N_1821,N_1862);
or U1999 (N_1999,N_1766,N_1761);
nand U2000 (N_2000,N_1923,N_1892);
or U2001 (N_2001,N_1905,N_1972);
nand U2002 (N_2002,N_1925,N_1979);
or U2003 (N_2003,N_1949,N_1968);
and U2004 (N_2004,N_1882,N_1919);
and U2005 (N_2005,N_1921,N_1898);
and U2006 (N_2006,N_1963,N_1960);
nand U2007 (N_2007,N_1899,N_1989);
or U2008 (N_2008,N_1961,N_1910);
nor U2009 (N_2009,N_1952,N_1916);
and U2010 (N_2010,N_1928,N_1965);
nand U2011 (N_2011,N_1911,N_1931);
or U2012 (N_2012,N_1980,N_1981);
nand U2013 (N_2013,N_1937,N_1966);
or U2014 (N_2014,N_1995,N_1954);
xor U2015 (N_2015,N_1973,N_1987);
nor U2016 (N_2016,N_1897,N_1984);
or U2017 (N_2017,N_1948,N_1967);
xnor U2018 (N_2018,N_1985,N_1906);
nor U2019 (N_2019,N_1976,N_1942);
and U2020 (N_2020,N_1909,N_1876);
nand U2021 (N_2021,N_1932,N_1939);
xor U2022 (N_2022,N_1951,N_1901);
xnor U2023 (N_2023,N_1946,N_1917);
or U2024 (N_2024,N_1885,N_1881);
and U2025 (N_2025,N_1969,N_1924);
or U2026 (N_2026,N_1978,N_1999);
xor U2027 (N_2027,N_1922,N_1996);
or U2028 (N_2028,N_1986,N_1927);
nand U2029 (N_2029,N_1904,N_1880);
xor U2030 (N_2030,N_1988,N_1920);
nand U2031 (N_2031,N_1982,N_1902);
nor U2032 (N_2032,N_1955,N_1957);
and U2033 (N_2033,N_1940,N_1935);
xnor U2034 (N_2034,N_1947,N_1887);
or U2035 (N_2035,N_1893,N_1894);
nand U2036 (N_2036,N_1992,N_1958);
xor U2037 (N_2037,N_1945,N_1883);
xor U2038 (N_2038,N_1900,N_1977);
nand U2039 (N_2039,N_1878,N_1914);
nand U2040 (N_2040,N_1929,N_1918);
nor U2041 (N_2041,N_1962,N_1936);
nor U2042 (N_2042,N_1884,N_1944);
or U2043 (N_2043,N_1912,N_1933);
or U2044 (N_2044,N_1938,N_1879);
xor U2045 (N_2045,N_1950,N_1998);
xor U2046 (N_2046,N_1964,N_1975);
xnor U2047 (N_2047,N_1956,N_1959);
nand U2048 (N_2048,N_1970,N_1994);
xnor U2049 (N_2049,N_1943,N_1934);
or U2050 (N_2050,N_1875,N_1915);
and U2051 (N_2051,N_1990,N_1907);
and U2052 (N_2052,N_1941,N_1983);
or U2053 (N_2053,N_1908,N_1971);
nor U2054 (N_2054,N_1903,N_1895);
or U2055 (N_2055,N_1877,N_1913);
nand U2056 (N_2056,N_1997,N_1993);
or U2057 (N_2057,N_1974,N_1886);
and U2058 (N_2058,N_1930,N_1991);
nor U2059 (N_2059,N_1888,N_1953);
nor U2060 (N_2060,N_1891,N_1896);
or U2061 (N_2061,N_1889,N_1890);
and U2062 (N_2062,N_1926,N_1973);
nand U2063 (N_2063,N_1884,N_1962);
nand U2064 (N_2064,N_1963,N_1997);
nand U2065 (N_2065,N_1908,N_1898);
nor U2066 (N_2066,N_1966,N_1931);
or U2067 (N_2067,N_1885,N_1957);
nor U2068 (N_2068,N_1903,N_1884);
nor U2069 (N_2069,N_1960,N_1920);
nor U2070 (N_2070,N_1920,N_1971);
nand U2071 (N_2071,N_1959,N_1996);
or U2072 (N_2072,N_1975,N_1915);
nand U2073 (N_2073,N_1890,N_1881);
nor U2074 (N_2074,N_1979,N_1927);
nand U2075 (N_2075,N_1956,N_1882);
xor U2076 (N_2076,N_1888,N_1956);
nor U2077 (N_2077,N_1926,N_1888);
or U2078 (N_2078,N_1944,N_1995);
or U2079 (N_2079,N_1919,N_1910);
or U2080 (N_2080,N_1940,N_1979);
nor U2081 (N_2081,N_1960,N_1990);
or U2082 (N_2082,N_1892,N_1985);
xnor U2083 (N_2083,N_1945,N_1939);
xor U2084 (N_2084,N_1919,N_1988);
or U2085 (N_2085,N_1915,N_1906);
nand U2086 (N_2086,N_1933,N_1922);
xnor U2087 (N_2087,N_1909,N_1935);
nand U2088 (N_2088,N_1913,N_1891);
and U2089 (N_2089,N_1892,N_1887);
or U2090 (N_2090,N_1901,N_1937);
xor U2091 (N_2091,N_1878,N_1950);
or U2092 (N_2092,N_1884,N_1987);
xnor U2093 (N_2093,N_1886,N_1896);
nor U2094 (N_2094,N_1891,N_1952);
xor U2095 (N_2095,N_1997,N_1920);
and U2096 (N_2096,N_1977,N_1953);
or U2097 (N_2097,N_1892,N_1917);
or U2098 (N_2098,N_1902,N_1893);
xor U2099 (N_2099,N_1898,N_1983);
or U2100 (N_2100,N_1909,N_1896);
and U2101 (N_2101,N_1998,N_1963);
nand U2102 (N_2102,N_1887,N_1898);
xor U2103 (N_2103,N_1914,N_1949);
nor U2104 (N_2104,N_1900,N_1927);
nand U2105 (N_2105,N_1980,N_1889);
and U2106 (N_2106,N_1946,N_1903);
or U2107 (N_2107,N_1981,N_1991);
or U2108 (N_2108,N_1991,N_1994);
or U2109 (N_2109,N_1940,N_1942);
nor U2110 (N_2110,N_1911,N_1881);
nor U2111 (N_2111,N_1905,N_1875);
xor U2112 (N_2112,N_1977,N_1979);
or U2113 (N_2113,N_1913,N_1914);
and U2114 (N_2114,N_1986,N_1890);
and U2115 (N_2115,N_1921,N_1990);
nor U2116 (N_2116,N_1981,N_1882);
and U2117 (N_2117,N_1877,N_1957);
or U2118 (N_2118,N_1883,N_1886);
nand U2119 (N_2119,N_1922,N_1925);
or U2120 (N_2120,N_1915,N_1953);
nor U2121 (N_2121,N_1905,N_1961);
nor U2122 (N_2122,N_1894,N_1955);
nor U2123 (N_2123,N_1887,N_1971);
or U2124 (N_2124,N_1924,N_1894);
nor U2125 (N_2125,N_2038,N_2107);
xor U2126 (N_2126,N_2015,N_2094);
nor U2127 (N_2127,N_2085,N_2005);
and U2128 (N_2128,N_2003,N_2102);
and U2129 (N_2129,N_2020,N_2012);
nand U2130 (N_2130,N_2081,N_2087);
or U2131 (N_2131,N_2034,N_2070);
xor U2132 (N_2132,N_2100,N_2104);
nand U2133 (N_2133,N_2018,N_2069);
xor U2134 (N_2134,N_2097,N_2121);
or U2135 (N_2135,N_2058,N_2096);
and U2136 (N_2136,N_2082,N_2116);
and U2137 (N_2137,N_2063,N_2090);
xnor U2138 (N_2138,N_2047,N_2077);
nand U2139 (N_2139,N_2055,N_2074);
nand U2140 (N_2140,N_2083,N_2039);
nand U2141 (N_2141,N_2093,N_2050);
nor U2142 (N_2142,N_2109,N_2006);
nand U2143 (N_2143,N_2098,N_2073);
nand U2144 (N_2144,N_2072,N_2029);
or U2145 (N_2145,N_2078,N_2008);
or U2146 (N_2146,N_2103,N_2106);
xnor U2147 (N_2147,N_2004,N_2000);
or U2148 (N_2148,N_2124,N_2042);
nor U2149 (N_2149,N_2043,N_2092);
nor U2150 (N_2150,N_2007,N_2037);
nor U2151 (N_2151,N_2028,N_2060);
or U2152 (N_2152,N_2067,N_2009);
and U2153 (N_2153,N_2064,N_2076);
xnor U2154 (N_2154,N_2075,N_2026);
or U2155 (N_2155,N_2071,N_2032);
nand U2156 (N_2156,N_2084,N_2051);
or U2157 (N_2157,N_2019,N_2017);
nand U2158 (N_2158,N_2059,N_2024);
nand U2159 (N_2159,N_2010,N_2086);
nand U2160 (N_2160,N_2068,N_2120);
or U2161 (N_2161,N_2117,N_2035);
nor U2162 (N_2162,N_2088,N_2011);
nand U2163 (N_2163,N_2123,N_2095);
xnor U2164 (N_2164,N_2065,N_2001);
or U2165 (N_2165,N_2030,N_2080);
nor U2166 (N_2166,N_2114,N_2033);
and U2167 (N_2167,N_2118,N_2048);
or U2168 (N_2168,N_2036,N_2112);
and U2169 (N_2169,N_2111,N_2023);
nand U2170 (N_2170,N_2105,N_2027);
and U2171 (N_2171,N_2049,N_2099);
xnor U2172 (N_2172,N_2040,N_2041);
and U2173 (N_2173,N_2045,N_2119);
or U2174 (N_2174,N_2053,N_2057);
or U2175 (N_2175,N_2115,N_2054);
nand U2176 (N_2176,N_2101,N_2113);
and U2177 (N_2177,N_2014,N_2122);
xnor U2178 (N_2178,N_2052,N_2056);
nor U2179 (N_2179,N_2031,N_2002);
nor U2180 (N_2180,N_2016,N_2091);
nor U2181 (N_2181,N_2079,N_2021);
and U2182 (N_2182,N_2046,N_2066);
nor U2183 (N_2183,N_2110,N_2062);
or U2184 (N_2184,N_2022,N_2108);
xnor U2185 (N_2185,N_2089,N_2044);
xor U2186 (N_2186,N_2025,N_2013);
and U2187 (N_2187,N_2061,N_2069);
nor U2188 (N_2188,N_2122,N_2073);
or U2189 (N_2189,N_2085,N_2026);
nand U2190 (N_2190,N_2077,N_2119);
nand U2191 (N_2191,N_2111,N_2084);
xnor U2192 (N_2192,N_2057,N_2076);
xor U2193 (N_2193,N_2072,N_2033);
or U2194 (N_2194,N_2081,N_2023);
nand U2195 (N_2195,N_2028,N_2093);
nor U2196 (N_2196,N_2076,N_2018);
and U2197 (N_2197,N_2000,N_2092);
and U2198 (N_2198,N_2035,N_2020);
xnor U2199 (N_2199,N_2046,N_2104);
nor U2200 (N_2200,N_2066,N_2013);
or U2201 (N_2201,N_2110,N_2074);
or U2202 (N_2202,N_2020,N_2018);
and U2203 (N_2203,N_2074,N_2005);
xor U2204 (N_2204,N_2110,N_2037);
or U2205 (N_2205,N_2115,N_2057);
nor U2206 (N_2206,N_2102,N_2067);
nor U2207 (N_2207,N_2011,N_2118);
xor U2208 (N_2208,N_2095,N_2087);
nand U2209 (N_2209,N_2034,N_2124);
and U2210 (N_2210,N_2089,N_2024);
or U2211 (N_2211,N_2089,N_2058);
xor U2212 (N_2212,N_2033,N_2100);
xnor U2213 (N_2213,N_2114,N_2049);
nor U2214 (N_2214,N_2053,N_2033);
nor U2215 (N_2215,N_2119,N_2034);
nor U2216 (N_2216,N_2016,N_2099);
nand U2217 (N_2217,N_2051,N_2085);
nand U2218 (N_2218,N_2078,N_2098);
nand U2219 (N_2219,N_2113,N_2104);
and U2220 (N_2220,N_2100,N_2026);
and U2221 (N_2221,N_2030,N_2014);
nor U2222 (N_2222,N_2083,N_2000);
xor U2223 (N_2223,N_2037,N_2089);
or U2224 (N_2224,N_2109,N_2000);
xnor U2225 (N_2225,N_2116,N_2121);
or U2226 (N_2226,N_2076,N_2104);
and U2227 (N_2227,N_2099,N_2088);
nor U2228 (N_2228,N_2098,N_2086);
and U2229 (N_2229,N_2072,N_2109);
xor U2230 (N_2230,N_2101,N_2114);
and U2231 (N_2231,N_2007,N_2027);
or U2232 (N_2232,N_2006,N_2072);
xor U2233 (N_2233,N_2078,N_2025);
nand U2234 (N_2234,N_2102,N_2116);
or U2235 (N_2235,N_2018,N_2046);
and U2236 (N_2236,N_2011,N_2113);
nor U2237 (N_2237,N_2090,N_2088);
or U2238 (N_2238,N_2113,N_2034);
nor U2239 (N_2239,N_2090,N_2104);
xnor U2240 (N_2240,N_2112,N_2122);
nand U2241 (N_2241,N_2095,N_2024);
or U2242 (N_2242,N_2070,N_2114);
or U2243 (N_2243,N_2043,N_2101);
nor U2244 (N_2244,N_2025,N_2109);
nor U2245 (N_2245,N_2109,N_2067);
nor U2246 (N_2246,N_2049,N_2044);
and U2247 (N_2247,N_2000,N_2079);
nor U2248 (N_2248,N_2085,N_2006);
nor U2249 (N_2249,N_2123,N_2053);
or U2250 (N_2250,N_2229,N_2232);
nand U2251 (N_2251,N_2233,N_2218);
nand U2252 (N_2252,N_2231,N_2138);
nor U2253 (N_2253,N_2167,N_2128);
or U2254 (N_2254,N_2130,N_2145);
xor U2255 (N_2255,N_2153,N_2149);
and U2256 (N_2256,N_2155,N_2202);
and U2257 (N_2257,N_2188,N_2141);
and U2258 (N_2258,N_2144,N_2239);
nand U2259 (N_2259,N_2224,N_2127);
nor U2260 (N_2260,N_2236,N_2154);
xor U2261 (N_2261,N_2192,N_2173);
or U2262 (N_2262,N_2193,N_2184);
nor U2263 (N_2263,N_2205,N_2219);
and U2264 (N_2264,N_2196,N_2163);
and U2265 (N_2265,N_2133,N_2198);
xor U2266 (N_2266,N_2142,N_2201);
or U2267 (N_2267,N_2182,N_2179);
and U2268 (N_2268,N_2131,N_2180);
and U2269 (N_2269,N_2209,N_2217);
and U2270 (N_2270,N_2165,N_2151);
and U2271 (N_2271,N_2140,N_2164);
xor U2272 (N_2272,N_2194,N_2222);
or U2273 (N_2273,N_2207,N_2204);
nor U2274 (N_2274,N_2146,N_2132);
nand U2275 (N_2275,N_2230,N_2187);
nand U2276 (N_2276,N_2223,N_2220);
xor U2277 (N_2277,N_2249,N_2214);
nor U2278 (N_2278,N_2147,N_2190);
xnor U2279 (N_2279,N_2195,N_2212);
and U2280 (N_2280,N_2243,N_2197);
and U2281 (N_2281,N_2169,N_2150);
xor U2282 (N_2282,N_2148,N_2170);
and U2283 (N_2283,N_2215,N_2175);
or U2284 (N_2284,N_2136,N_2172);
nand U2285 (N_2285,N_2189,N_2159);
nor U2286 (N_2286,N_2237,N_2227);
nand U2287 (N_2287,N_2241,N_2174);
or U2288 (N_2288,N_2221,N_2246);
xor U2289 (N_2289,N_2247,N_2199);
and U2290 (N_2290,N_2208,N_2211);
xnor U2291 (N_2291,N_2152,N_2139);
xnor U2292 (N_2292,N_2157,N_2186);
nand U2293 (N_2293,N_2178,N_2183);
or U2294 (N_2294,N_2158,N_2235);
and U2295 (N_2295,N_2129,N_2171);
nand U2296 (N_2296,N_2137,N_2203);
or U2297 (N_2297,N_2200,N_2191);
and U2298 (N_2298,N_2242,N_2160);
nand U2299 (N_2299,N_2228,N_2216);
and U2300 (N_2300,N_2156,N_2177);
or U2301 (N_2301,N_2176,N_2238);
or U2302 (N_2302,N_2161,N_2143);
and U2303 (N_2303,N_2240,N_2134);
or U2304 (N_2304,N_2126,N_2185);
nand U2305 (N_2305,N_2248,N_2226);
xnor U2306 (N_2306,N_2210,N_2166);
nand U2307 (N_2307,N_2206,N_2245);
xnor U2308 (N_2308,N_2125,N_2225);
xor U2309 (N_2309,N_2168,N_2213);
and U2310 (N_2310,N_2162,N_2135);
or U2311 (N_2311,N_2234,N_2244);
nor U2312 (N_2312,N_2181,N_2227);
nand U2313 (N_2313,N_2197,N_2178);
and U2314 (N_2314,N_2199,N_2190);
or U2315 (N_2315,N_2237,N_2137);
and U2316 (N_2316,N_2161,N_2148);
xnor U2317 (N_2317,N_2205,N_2206);
or U2318 (N_2318,N_2196,N_2170);
or U2319 (N_2319,N_2247,N_2245);
xnor U2320 (N_2320,N_2169,N_2226);
xnor U2321 (N_2321,N_2231,N_2219);
nand U2322 (N_2322,N_2233,N_2198);
or U2323 (N_2323,N_2149,N_2147);
or U2324 (N_2324,N_2224,N_2167);
or U2325 (N_2325,N_2221,N_2200);
nor U2326 (N_2326,N_2216,N_2199);
or U2327 (N_2327,N_2214,N_2132);
nand U2328 (N_2328,N_2178,N_2173);
xnor U2329 (N_2329,N_2155,N_2153);
and U2330 (N_2330,N_2223,N_2196);
nand U2331 (N_2331,N_2218,N_2229);
nand U2332 (N_2332,N_2228,N_2167);
xor U2333 (N_2333,N_2221,N_2154);
nor U2334 (N_2334,N_2225,N_2163);
and U2335 (N_2335,N_2249,N_2156);
and U2336 (N_2336,N_2191,N_2240);
and U2337 (N_2337,N_2153,N_2151);
or U2338 (N_2338,N_2151,N_2148);
nand U2339 (N_2339,N_2134,N_2130);
or U2340 (N_2340,N_2138,N_2130);
or U2341 (N_2341,N_2153,N_2176);
xor U2342 (N_2342,N_2240,N_2232);
nand U2343 (N_2343,N_2172,N_2232);
or U2344 (N_2344,N_2126,N_2229);
or U2345 (N_2345,N_2238,N_2224);
nor U2346 (N_2346,N_2183,N_2228);
or U2347 (N_2347,N_2249,N_2142);
nor U2348 (N_2348,N_2155,N_2189);
nand U2349 (N_2349,N_2154,N_2162);
or U2350 (N_2350,N_2214,N_2156);
nand U2351 (N_2351,N_2170,N_2167);
nor U2352 (N_2352,N_2163,N_2235);
or U2353 (N_2353,N_2133,N_2202);
and U2354 (N_2354,N_2187,N_2238);
and U2355 (N_2355,N_2125,N_2169);
or U2356 (N_2356,N_2190,N_2226);
nor U2357 (N_2357,N_2221,N_2209);
nand U2358 (N_2358,N_2200,N_2224);
xor U2359 (N_2359,N_2188,N_2201);
nand U2360 (N_2360,N_2175,N_2151);
nor U2361 (N_2361,N_2201,N_2179);
or U2362 (N_2362,N_2127,N_2222);
xor U2363 (N_2363,N_2176,N_2128);
nor U2364 (N_2364,N_2142,N_2171);
or U2365 (N_2365,N_2183,N_2148);
and U2366 (N_2366,N_2167,N_2147);
nand U2367 (N_2367,N_2139,N_2151);
nand U2368 (N_2368,N_2211,N_2189);
or U2369 (N_2369,N_2148,N_2186);
and U2370 (N_2370,N_2206,N_2204);
xnor U2371 (N_2371,N_2132,N_2133);
or U2372 (N_2372,N_2205,N_2161);
nor U2373 (N_2373,N_2219,N_2154);
nand U2374 (N_2374,N_2129,N_2167);
and U2375 (N_2375,N_2254,N_2252);
xnor U2376 (N_2376,N_2322,N_2257);
and U2377 (N_2377,N_2284,N_2253);
and U2378 (N_2378,N_2273,N_2350);
nand U2379 (N_2379,N_2367,N_2277);
xor U2380 (N_2380,N_2255,N_2270);
xor U2381 (N_2381,N_2360,N_2371);
xor U2382 (N_2382,N_2356,N_2261);
xnor U2383 (N_2383,N_2309,N_2288);
or U2384 (N_2384,N_2313,N_2324);
nor U2385 (N_2385,N_2279,N_2352);
nand U2386 (N_2386,N_2302,N_2272);
and U2387 (N_2387,N_2365,N_2264);
nor U2388 (N_2388,N_2323,N_2334);
nor U2389 (N_2389,N_2280,N_2336);
xnor U2390 (N_2390,N_2266,N_2312);
or U2391 (N_2391,N_2263,N_2287);
or U2392 (N_2392,N_2256,N_2316);
xnor U2393 (N_2393,N_2301,N_2291);
or U2394 (N_2394,N_2359,N_2320);
nor U2395 (N_2395,N_2298,N_2321);
nor U2396 (N_2396,N_2317,N_2271);
xor U2397 (N_2397,N_2300,N_2297);
and U2398 (N_2398,N_2346,N_2315);
xor U2399 (N_2399,N_2258,N_2357);
nor U2400 (N_2400,N_2276,N_2342);
or U2401 (N_2401,N_2260,N_2274);
xnor U2402 (N_2402,N_2325,N_2289);
or U2403 (N_2403,N_2267,N_2310);
nand U2404 (N_2404,N_2327,N_2281);
nand U2405 (N_2405,N_2348,N_2335);
or U2406 (N_2406,N_2283,N_2293);
nand U2407 (N_2407,N_2250,N_2340);
nand U2408 (N_2408,N_2311,N_2296);
and U2409 (N_2409,N_2354,N_2286);
or U2410 (N_2410,N_2307,N_2339);
nand U2411 (N_2411,N_2366,N_2308);
nand U2412 (N_2412,N_2251,N_2328);
and U2413 (N_2413,N_2268,N_2330);
nor U2414 (N_2414,N_2294,N_2373);
and U2415 (N_2415,N_2299,N_2347);
nor U2416 (N_2416,N_2275,N_2319);
and U2417 (N_2417,N_2370,N_2349);
and U2418 (N_2418,N_2304,N_2331);
and U2419 (N_2419,N_2333,N_2332);
nor U2420 (N_2420,N_2343,N_2338);
nor U2421 (N_2421,N_2326,N_2290);
and U2422 (N_2422,N_2303,N_2372);
nand U2423 (N_2423,N_2278,N_2329);
xnor U2424 (N_2424,N_2318,N_2314);
nor U2425 (N_2425,N_2358,N_2265);
nand U2426 (N_2426,N_2292,N_2295);
or U2427 (N_2427,N_2306,N_2361);
and U2428 (N_2428,N_2374,N_2259);
and U2429 (N_2429,N_2351,N_2285);
nor U2430 (N_2430,N_2364,N_2363);
or U2431 (N_2431,N_2262,N_2369);
and U2432 (N_2432,N_2269,N_2282);
or U2433 (N_2433,N_2305,N_2355);
or U2434 (N_2434,N_2344,N_2341);
nand U2435 (N_2435,N_2362,N_2345);
or U2436 (N_2436,N_2368,N_2353);
nor U2437 (N_2437,N_2337,N_2351);
and U2438 (N_2438,N_2287,N_2314);
or U2439 (N_2439,N_2301,N_2363);
xnor U2440 (N_2440,N_2370,N_2311);
xnor U2441 (N_2441,N_2304,N_2253);
nand U2442 (N_2442,N_2260,N_2345);
and U2443 (N_2443,N_2306,N_2264);
xor U2444 (N_2444,N_2284,N_2341);
and U2445 (N_2445,N_2346,N_2328);
and U2446 (N_2446,N_2334,N_2299);
and U2447 (N_2447,N_2329,N_2369);
or U2448 (N_2448,N_2366,N_2315);
nand U2449 (N_2449,N_2341,N_2368);
nor U2450 (N_2450,N_2293,N_2367);
nor U2451 (N_2451,N_2335,N_2362);
nand U2452 (N_2452,N_2358,N_2311);
nand U2453 (N_2453,N_2305,N_2329);
or U2454 (N_2454,N_2257,N_2337);
nand U2455 (N_2455,N_2317,N_2261);
and U2456 (N_2456,N_2294,N_2323);
or U2457 (N_2457,N_2335,N_2257);
xor U2458 (N_2458,N_2269,N_2295);
nand U2459 (N_2459,N_2335,N_2291);
nand U2460 (N_2460,N_2352,N_2363);
xor U2461 (N_2461,N_2277,N_2268);
and U2462 (N_2462,N_2265,N_2350);
xor U2463 (N_2463,N_2287,N_2366);
or U2464 (N_2464,N_2357,N_2333);
and U2465 (N_2465,N_2320,N_2251);
nand U2466 (N_2466,N_2316,N_2359);
nor U2467 (N_2467,N_2340,N_2300);
and U2468 (N_2468,N_2289,N_2266);
nor U2469 (N_2469,N_2269,N_2337);
and U2470 (N_2470,N_2298,N_2355);
and U2471 (N_2471,N_2268,N_2310);
xnor U2472 (N_2472,N_2307,N_2326);
nor U2473 (N_2473,N_2363,N_2309);
xnor U2474 (N_2474,N_2251,N_2354);
nor U2475 (N_2475,N_2268,N_2287);
nor U2476 (N_2476,N_2282,N_2369);
or U2477 (N_2477,N_2307,N_2341);
and U2478 (N_2478,N_2304,N_2308);
nor U2479 (N_2479,N_2309,N_2304);
or U2480 (N_2480,N_2297,N_2272);
xor U2481 (N_2481,N_2316,N_2302);
nor U2482 (N_2482,N_2360,N_2257);
or U2483 (N_2483,N_2355,N_2352);
or U2484 (N_2484,N_2319,N_2370);
xor U2485 (N_2485,N_2338,N_2354);
xor U2486 (N_2486,N_2328,N_2351);
nand U2487 (N_2487,N_2340,N_2333);
and U2488 (N_2488,N_2337,N_2258);
and U2489 (N_2489,N_2252,N_2266);
and U2490 (N_2490,N_2340,N_2285);
xnor U2491 (N_2491,N_2348,N_2353);
and U2492 (N_2492,N_2334,N_2271);
nand U2493 (N_2493,N_2308,N_2370);
xnor U2494 (N_2494,N_2328,N_2275);
xnor U2495 (N_2495,N_2352,N_2268);
or U2496 (N_2496,N_2277,N_2355);
or U2497 (N_2497,N_2265,N_2258);
nand U2498 (N_2498,N_2277,N_2279);
and U2499 (N_2499,N_2294,N_2276);
and U2500 (N_2500,N_2439,N_2408);
nand U2501 (N_2501,N_2447,N_2380);
xnor U2502 (N_2502,N_2490,N_2438);
or U2503 (N_2503,N_2395,N_2496);
xor U2504 (N_2504,N_2389,N_2468);
nor U2505 (N_2505,N_2497,N_2430);
nor U2506 (N_2506,N_2426,N_2428);
or U2507 (N_2507,N_2472,N_2471);
nand U2508 (N_2508,N_2383,N_2425);
nor U2509 (N_2509,N_2416,N_2449);
nand U2510 (N_2510,N_2381,N_2494);
nand U2511 (N_2511,N_2410,N_2463);
or U2512 (N_2512,N_2467,N_2495);
nor U2513 (N_2513,N_2435,N_2406);
and U2514 (N_2514,N_2485,N_2484);
and U2515 (N_2515,N_2407,N_2459);
and U2516 (N_2516,N_2479,N_2436);
xnor U2517 (N_2517,N_2441,N_2415);
nor U2518 (N_2518,N_2431,N_2394);
nor U2519 (N_2519,N_2391,N_2448);
nand U2520 (N_2520,N_2477,N_2433);
xor U2521 (N_2521,N_2424,N_2390);
nor U2522 (N_2522,N_2385,N_2491);
or U2523 (N_2523,N_2453,N_2401);
xor U2524 (N_2524,N_2451,N_2392);
nor U2525 (N_2525,N_2411,N_2469);
or U2526 (N_2526,N_2404,N_2414);
or U2527 (N_2527,N_2418,N_2375);
nor U2528 (N_2528,N_2455,N_2452);
nand U2529 (N_2529,N_2420,N_2386);
and U2530 (N_2530,N_2481,N_2444);
and U2531 (N_2531,N_2443,N_2461);
nor U2532 (N_2532,N_2437,N_2387);
nor U2533 (N_2533,N_2454,N_2400);
nand U2534 (N_2534,N_2384,N_2475);
or U2535 (N_2535,N_2417,N_2402);
nor U2536 (N_2536,N_2399,N_2434);
and U2537 (N_2537,N_2480,N_2377);
or U2538 (N_2538,N_2450,N_2470);
xnor U2539 (N_2539,N_2409,N_2421);
nor U2540 (N_2540,N_2466,N_2440);
nor U2541 (N_2541,N_2379,N_2464);
and U2542 (N_2542,N_2465,N_2458);
nor U2543 (N_2543,N_2442,N_2422);
xnor U2544 (N_2544,N_2405,N_2446);
nor U2545 (N_2545,N_2493,N_2398);
and U2546 (N_2546,N_2488,N_2393);
xnor U2547 (N_2547,N_2492,N_2427);
or U2548 (N_2548,N_2487,N_2498);
nand U2549 (N_2549,N_2445,N_2396);
nand U2550 (N_2550,N_2419,N_2397);
or U2551 (N_2551,N_2382,N_2423);
xnor U2552 (N_2552,N_2378,N_2462);
xor U2553 (N_2553,N_2412,N_2489);
or U2554 (N_2554,N_2413,N_2473);
xor U2555 (N_2555,N_2499,N_2483);
xor U2556 (N_2556,N_2429,N_2460);
or U2557 (N_2557,N_2478,N_2403);
nand U2558 (N_2558,N_2457,N_2474);
and U2559 (N_2559,N_2432,N_2476);
and U2560 (N_2560,N_2486,N_2376);
and U2561 (N_2561,N_2388,N_2456);
xnor U2562 (N_2562,N_2482,N_2489);
and U2563 (N_2563,N_2401,N_2436);
xor U2564 (N_2564,N_2464,N_2421);
nor U2565 (N_2565,N_2436,N_2447);
and U2566 (N_2566,N_2485,N_2414);
nand U2567 (N_2567,N_2432,N_2483);
nand U2568 (N_2568,N_2395,N_2484);
nand U2569 (N_2569,N_2492,N_2441);
or U2570 (N_2570,N_2470,N_2376);
xnor U2571 (N_2571,N_2393,N_2403);
nand U2572 (N_2572,N_2384,N_2499);
xor U2573 (N_2573,N_2465,N_2469);
xor U2574 (N_2574,N_2418,N_2483);
nor U2575 (N_2575,N_2405,N_2418);
or U2576 (N_2576,N_2450,N_2483);
xnor U2577 (N_2577,N_2414,N_2410);
and U2578 (N_2578,N_2418,N_2479);
nor U2579 (N_2579,N_2432,N_2489);
nor U2580 (N_2580,N_2393,N_2435);
and U2581 (N_2581,N_2459,N_2446);
nand U2582 (N_2582,N_2425,N_2386);
and U2583 (N_2583,N_2459,N_2449);
nor U2584 (N_2584,N_2402,N_2465);
or U2585 (N_2585,N_2469,N_2454);
and U2586 (N_2586,N_2414,N_2397);
and U2587 (N_2587,N_2385,N_2468);
or U2588 (N_2588,N_2386,N_2399);
xor U2589 (N_2589,N_2470,N_2463);
xor U2590 (N_2590,N_2400,N_2434);
nand U2591 (N_2591,N_2412,N_2454);
or U2592 (N_2592,N_2388,N_2444);
or U2593 (N_2593,N_2455,N_2389);
nand U2594 (N_2594,N_2465,N_2438);
nor U2595 (N_2595,N_2475,N_2389);
or U2596 (N_2596,N_2431,N_2473);
nor U2597 (N_2597,N_2398,N_2475);
nor U2598 (N_2598,N_2472,N_2498);
nor U2599 (N_2599,N_2495,N_2414);
xnor U2600 (N_2600,N_2390,N_2403);
nand U2601 (N_2601,N_2425,N_2436);
nand U2602 (N_2602,N_2417,N_2478);
nor U2603 (N_2603,N_2480,N_2393);
or U2604 (N_2604,N_2434,N_2416);
xnor U2605 (N_2605,N_2497,N_2471);
and U2606 (N_2606,N_2427,N_2423);
xor U2607 (N_2607,N_2471,N_2376);
and U2608 (N_2608,N_2453,N_2482);
or U2609 (N_2609,N_2390,N_2444);
or U2610 (N_2610,N_2413,N_2492);
xor U2611 (N_2611,N_2421,N_2398);
xnor U2612 (N_2612,N_2395,N_2399);
and U2613 (N_2613,N_2435,N_2475);
or U2614 (N_2614,N_2388,N_2379);
and U2615 (N_2615,N_2460,N_2481);
nor U2616 (N_2616,N_2400,N_2433);
nand U2617 (N_2617,N_2446,N_2401);
nor U2618 (N_2618,N_2402,N_2481);
or U2619 (N_2619,N_2441,N_2411);
and U2620 (N_2620,N_2442,N_2431);
or U2621 (N_2621,N_2493,N_2443);
or U2622 (N_2622,N_2415,N_2485);
xor U2623 (N_2623,N_2417,N_2414);
xnor U2624 (N_2624,N_2404,N_2376);
nand U2625 (N_2625,N_2543,N_2563);
xnor U2626 (N_2626,N_2613,N_2533);
nand U2627 (N_2627,N_2589,N_2513);
or U2628 (N_2628,N_2588,N_2506);
xnor U2629 (N_2629,N_2548,N_2527);
or U2630 (N_2630,N_2587,N_2584);
nor U2631 (N_2631,N_2599,N_2518);
xor U2632 (N_2632,N_2524,N_2593);
or U2633 (N_2633,N_2609,N_2585);
or U2634 (N_2634,N_2586,N_2536);
xor U2635 (N_2635,N_2614,N_2620);
or U2636 (N_2636,N_2608,N_2534);
nand U2637 (N_2637,N_2551,N_2594);
or U2638 (N_2638,N_2601,N_2550);
xnor U2639 (N_2639,N_2544,N_2610);
or U2640 (N_2640,N_2616,N_2532);
and U2641 (N_2641,N_2528,N_2503);
nand U2642 (N_2642,N_2570,N_2545);
and U2643 (N_2643,N_2529,N_2603);
nand U2644 (N_2644,N_2549,N_2615);
or U2645 (N_2645,N_2520,N_2501);
or U2646 (N_2646,N_2623,N_2619);
and U2647 (N_2647,N_2574,N_2592);
and U2648 (N_2648,N_2602,N_2515);
xnor U2649 (N_2649,N_2617,N_2531);
xnor U2650 (N_2650,N_2547,N_2541);
nand U2651 (N_2651,N_2517,N_2582);
nor U2652 (N_2652,N_2578,N_2604);
xnor U2653 (N_2653,N_2576,N_2596);
xor U2654 (N_2654,N_2552,N_2612);
nand U2655 (N_2655,N_2502,N_2580);
or U2656 (N_2656,N_2561,N_2510);
or U2657 (N_2657,N_2571,N_2525);
xnor U2658 (N_2658,N_2572,N_2542);
and U2659 (N_2659,N_2507,N_2575);
or U2660 (N_2660,N_2560,N_2516);
xor U2661 (N_2661,N_2591,N_2569);
nand U2662 (N_2662,N_2505,N_2624);
xor U2663 (N_2663,N_2562,N_2538);
and U2664 (N_2664,N_2553,N_2621);
nor U2665 (N_2665,N_2522,N_2607);
and U2666 (N_2666,N_2537,N_2508);
and U2667 (N_2667,N_2546,N_2558);
or U2668 (N_2668,N_2514,N_2600);
or U2669 (N_2669,N_2597,N_2581);
nor U2670 (N_2670,N_2598,N_2521);
nor U2671 (N_2671,N_2500,N_2618);
nor U2672 (N_2672,N_2565,N_2568);
nand U2673 (N_2673,N_2554,N_2611);
and U2674 (N_2674,N_2595,N_2605);
and U2675 (N_2675,N_2564,N_2606);
nand U2676 (N_2676,N_2566,N_2583);
or U2677 (N_2677,N_2523,N_2511);
nor U2678 (N_2678,N_2590,N_2556);
and U2679 (N_2679,N_2509,N_2577);
nand U2680 (N_2680,N_2530,N_2535);
or U2681 (N_2681,N_2559,N_2622);
or U2682 (N_2682,N_2512,N_2504);
nor U2683 (N_2683,N_2526,N_2579);
nand U2684 (N_2684,N_2573,N_2555);
and U2685 (N_2685,N_2567,N_2557);
xor U2686 (N_2686,N_2539,N_2540);
xor U2687 (N_2687,N_2519,N_2553);
nand U2688 (N_2688,N_2541,N_2606);
and U2689 (N_2689,N_2506,N_2510);
or U2690 (N_2690,N_2532,N_2540);
or U2691 (N_2691,N_2563,N_2557);
nor U2692 (N_2692,N_2516,N_2607);
and U2693 (N_2693,N_2530,N_2542);
or U2694 (N_2694,N_2594,N_2520);
and U2695 (N_2695,N_2555,N_2602);
or U2696 (N_2696,N_2515,N_2547);
xor U2697 (N_2697,N_2518,N_2602);
xnor U2698 (N_2698,N_2592,N_2590);
nor U2699 (N_2699,N_2619,N_2579);
nor U2700 (N_2700,N_2500,N_2565);
and U2701 (N_2701,N_2531,N_2563);
and U2702 (N_2702,N_2552,N_2595);
and U2703 (N_2703,N_2540,N_2522);
nor U2704 (N_2704,N_2559,N_2551);
and U2705 (N_2705,N_2521,N_2546);
and U2706 (N_2706,N_2505,N_2598);
or U2707 (N_2707,N_2604,N_2590);
and U2708 (N_2708,N_2517,N_2548);
nor U2709 (N_2709,N_2574,N_2589);
nand U2710 (N_2710,N_2533,N_2615);
nand U2711 (N_2711,N_2540,N_2619);
nand U2712 (N_2712,N_2566,N_2568);
or U2713 (N_2713,N_2560,N_2556);
nor U2714 (N_2714,N_2502,N_2531);
or U2715 (N_2715,N_2616,N_2618);
and U2716 (N_2716,N_2568,N_2603);
nand U2717 (N_2717,N_2522,N_2527);
or U2718 (N_2718,N_2525,N_2504);
xnor U2719 (N_2719,N_2568,N_2538);
nor U2720 (N_2720,N_2590,N_2500);
xor U2721 (N_2721,N_2524,N_2614);
nand U2722 (N_2722,N_2500,N_2572);
xor U2723 (N_2723,N_2529,N_2534);
nand U2724 (N_2724,N_2560,N_2593);
and U2725 (N_2725,N_2577,N_2541);
xnor U2726 (N_2726,N_2552,N_2602);
nor U2727 (N_2727,N_2560,N_2566);
nand U2728 (N_2728,N_2538,N_2563);
nor U2729 (N_2729,N_2525,N_2542);
nand U2730 (N_2730,N_2516,N_2550);
and U2731 (N_2731,N_2592,N_2529);
or U2732 (N_2732,N_2523,N_2562);
nand U2733 (N_2733,N_2551,N_2513);
nor U2734 (N_2734,N_2542,N_2597);
nand U2735 (N_2735,N_2547,N_2509);
nand U2736 (N_2736,N_2519,N_2532);
or U2737 (N_2737,N_2565,N_2556);
nand U2738 (N_2738,N_2578,N_2555);
and U2739 (N_2739,N_2514,N_2507);
xor U2740 (N_2740,N_2586,N_2572);
nor U2741 (N_2741,N_2557,N_2549);
nor U2742 (N_2742,N_2566,N_2623);
nand U2743 (N_2743,N_2623,N_2583);
nor U2744 (N_2744,N_2603,N_2544);
nand U2745 (N_2745,N_2605,N_2601);
or U2746 (N_2746,N_2595,N_2569);
xnor U2747 (N_2747,N_2530,N_2559);
or U2748 (N_2748,N_2614,N_2530);
nand U2749 (N_2749,N_2557,N_2613);
xor U2750 (N_2750,N_2678,N_2676);
xnor U2751 (N_2751,N_2709,N_2726);
and U2752 (N_2752,N_2644,N_2720);
and U2753 (N_2753,N_2730,N_2652);
nor U2754 (N_2754,N_2645,N_2684);
xor U2755 (N_2755,N_2663,N_2685);
nand U2756 (N_2756,N_2653,N_2735);
nor U2757 (N_2757,N_2675,N_2748);
or U2758 (N_2758,N_2740,N_2744);
or U2759 (N_2759,N_2641,N_2650);
nor U2760 (N_2760,N_2712,N_2629);
or U2761 (N_2761,N_2706,N_2746);
and U2762 (N_2762,N_2673,N_2669);
and U2763 (N_2763,N_2634,N_2711);
and U2764 (N_2764,N_2661,N_2693);
and U2765 (N_2765,N_2638,N_2691);
or U2766 (N_2766,N_2695,N_2659);
or U2767 (N_2767,N_2640,N_2725);
nor U2768 (N_2768,N_2665,N_2660);
and U2769 (N_2769,N_2636,N_2738);
and U2770 (N_2770,N_2626,N_2639);
and U2771 (N_2771,N_2716,N_2700);
nand U2772 (N_2772,N_2657,N_2646);
xnor U2773 (N_2773,N_2731,N_2666);
nand U2774 (N_2774,N_2713,N_2707);
nor U2775 (N_2775,N_2719,N_2747);
xnor U2776 (N_2776,N_2701,N_2642);
xnor U2777 (N_2777,N_2687,N_2633);
xnor U2778 (N_2778,N_2728,N_2743);
and U2779 (N_2779,N_2635,N_2699);
xor U2780 (N_2780,N_2689,N_2702);
nor U2781 (N_2781,N_2690,N_2734);
or U2782 (N_2782,N_2704,N_2741);
nand U2783 (N_2783,N_2627,N_2697);
xor U2784 (N_2784,N_2667,N_2727);
and U2785 (N_2785,N_2737,N_2654);
nand U2786 (N_2786,N_2670,N_2625);
nor U2787 (N_2787,N_2630,N_2723);
xnor U2788 (N_2788,N_2749,N_2643);
xnor U2789 (N_2789,N_2742,N_2722);
or U2790 (N_2790,N_2677,N_2739);
nor U2791 (N_2791,N_2717,N_2688);
nor U2792 (N_2792,N_2703,N_2705);
xnor U2793 (N_2793,N_2718,N_2637);
nor U2794 (N_2794,N_2710,N_2721);
xor U2795 (N_2795,N_2674,N_2745);
or U2796 (N_2796,N_2628,N_2647);
xor U2797 (N_2797,N_2672,N_2671);
xnor U2798 (N_2798,N_2649,N_2708);
or U2799 (N_2799,N_2651,N_2662);
and U2800 (N_2800,N_2683,N_2632);
xnor U2801 (N_2801,N_2736,N_2682);
xor U2802 (N_2802,N_2696,N_2664);
nor U2803 (N_2803,N_2733,N_2631);
nand U2804 (N_2804,N_2679,N_2656);
and U2805 (N_2805,N_2686,N_2715);
and U2806 (N_2806,N_2729,N_2668);
and U2807 (N_2807,N_2698,N_2655);
nand U2808 (N_2808,N_2658,N_2714);
or U2809 (N_2809,N_2692,N_2694);
nand U2810 (N_2810,N_2724,N_2680);
xnor U2811 (N_2811,N_2648,N_2732);
or U2812 (N_2812,N_2681,N_2625);
nand U2813 (N_2813,N_2642,N_2740);
or U2814 (N_2814,N_2637,N_2669);
xnor U2815 (N_2815,N_2647,N_2691);
nor U2816 (N_2816,N_2635,N_2718);
xor U2817 (N_2817,N_2682,N_2737);
or U2818 (N_2818,N_2698,N_2660);
and U2819 (N_2819,N_2740,N_2634);
xor U2820 (N_2820,N_2706,N_2718);
nand U2821 (N_2821,N_2705,N_2653);
or U2822 (N_2822,N_2681,N_2635);
and U2823 (N_2823,N_2659,N_2630);
nand U2824 (N_2824,N_2630,N_2722);
nor U2825 (N_2825,N_2650,N_2634);
nand U2826 (N_2826,N_2656,N_2711);
or U2827 (N_2827,N_2642,N_2628);
nor U2828 (N_2828,N_2633,N_2704);
nand U2829 (N_2829,N_2715,N_2719);
xor U2830 (N_2830,N_2690,N_2730);
nor U2831 (N_2831,N_2648,N_2680);
nand U2832 (N_2832,N_2706,N_2710);
nor U2833 (N_2833,N_2633,N_2745);
xnor U2834 (N_2834,N_2642,N_2688);
nor U2835 (N_2835,N_2669,N_2671);
nand U2836 (N_2836,N_2655,N_2651);
and U2837 (N_2837,N_2690,N_2696);
nor U2838 (N_2838,N_2722,N_2710);
nand U2839 (N_2839,N_2703,N_2625);
and U2840 (N_2840,N_2684,N_2704);
and U2841 (N_2841,N_2702,N_2672);
nor U2842 (N_2842,N_2686,N_2713);
or U2843 (N_2843,N_2745,N_2643);
xor U2844 (N_2844,N_2650,N_2677);
nor U2845 (N_2845,N_2667,N_2740);
and U2846 (N_2846,N_2682,N_2688);
or U2847 (N_2847,N_2747,N_2679);
nor U2848 (N_2848,N_2687,N_2694);
or U2849 (N_2849,N_2684,N_2717);
xnor U2850 (N_2850,N_2699,N_2681);
and U2851 (N_2851,N_2693,N_2672);
nor U2852 (N_2852,N_2721,N_2706);
or U2853 (N_2853,N_2626,N_2718);
and U2854 (N_2854,N_2638,N_2653);
nor U2855 (N_2855,N_2736,N_2724);
nand U2856 (N_2856,N_2646,N_2633);
and U2857 (N_2857,N_2635,N_2678);
and U2858 (N_2858,N_2705,N_2744);
xnor U2859 (N_2859,N_2712,N_2739);
and U2860 (N_2860,N_2742,N_2668);
nor U2861 (N_2861,N_2727,N_2689);
or U2862 (N_2862,N_2695,N_2735);
or U2863 (N_2863,N_2655,N_2740);
xor U2864 (N_2864,N_2716,N_2680);
or U2865 (N_2865,N_2666,N_2712);
nand U2866 (N_2866,N_2670,N_2662);
nor U2867 (N_2867,N_2715,N_2664);
or U2868 (N_2868,N_2730,N_2638);
nor U2869 (N_2869,N_2717,N_2719);
nor U2870 (N_2870,N_2667,N_2657);
xnor U2871 (N_2871,N_2686,N_2726);
nand U2872 (N_2872,N_2637,N_2678);
or U2873 (N_2873,N_2629,N_2654);
nand U2874 (N_2874,N_2735,N_2737);
nand U2875 (N_2875,N_2831,N_2757);
nor U2876 (N_2876,N_2782,N_2838);
nand U2877 (N_2877,N_2816,N_2864);
nand U2878 (N_2878,N_2760,N_2813);
nand U2879 (N_2879,N_2872,N_2859);
or U2880 (N_2880,N_2826,N_2833);
and U2881 (N_2881,N_2874,N_2800);
nor U2882 (N_2882,N_2828,N_2865);
and U2883 (N_2883,N_2769,N_2799);
nand U2884 (N_2884,N_2750,N_2784);
nor U2885 (N_2885,N_2790,N_2755);
or U2886 (N_2886,N_2855,N_2804);
or U2887 (N_2887,N_2763,N_2817);
and U2888 (N_2888,N_2815,N_2762);
or U2889 (N_2889,N_2824,N_2845);
or U2890 (N_2890,N_2780,N_2772);
nor U2891 (N_2891,N_2779,N_2798);
xor U2892 (N_2892,N_2837,N_2751);
and U2893 (N_2893,N_2811,N_2848);
and U2894 (N_2894,N_2842,N_2856);
xnor U2895 (N_2895,N_2778,N_2850);
nand U2896 (N_2896,N_2777,N_2793);
or U2897 (N_2897,N_2805,N_2767);
nand U2898 (N_2898,N_2832,N_2776);
nand U2899 (N_2899,N_2808,N_2871);
nand U2900 (N_2900,N_2787,N_2812);
xnor U2901 (N_2901,N_2797,N_2774);
and U2902 (N_2902,N_2814,N_2775);
or U2903 (N_2903,N_2771,N_2795);
nand U2904 (N_2904,N_2766,N_2768);
xor U2905 (N_2905,N_2868,N_2796);
and U2906 (N_2906,N_2792,N_2830);
or U2907 (N_2907,N_2841,N_2756);
and U2908 (N_2908,N_2773,N_2840);
and U2909 (N_2909,N_2809,N_2835);
nand U2910 (N_2910,N_2758,N_2844);
nand U2911 (N_2911,N_2802,N_2788);
nand U2912 (N_2912,N_2851,N_2807);
nor U2913 (N_2913,N_2858,N_2754);
nand U2914 (N_2914,N_2854,N_2862);
or U2915 (N_2915,N_2786,N_2801);
nor U2916 (N_2916,N_2819,N_2794);
nor U2917 (N_2917,N_2829,N_2820);
xnor U2918 (N_2918,N_2839,N_2827);
xnor U2919 (N_2919,N_2823,N_2810);
or U2920 (N_2920,N_2765,N_2759);
nor U2921 (N_2921,N_2860,N_2770);
nor U2922 (N_2922,N_2822,N_2870);
and U2923 (N_2923,N_2857,N_2764);
xor U2924 (N_2924,N_2869,N_2861);
nand U2925 (N_2925,N_2825,N_2846);
or U2926 (N_2926,N_2753,N_2821);
and U2927 (N_2927,N_2785,N_2836);
nand U2928 (N_2928,N_2852,N_2847);
xor U2929 (N_2929,N_2818,N_2863);
nand U2930 (N_2930,N_2806,N_2834);
nand U2931 (N_2931,N_2803,N_2791);
or U2932 (N_2932,N_2761,N_2843);
and U2933 (N_2933,N_2789,N_2866);
nor U2934 (N_2934,N_2849,N_2752);
nor U2935 (N_2935,N_2781,N_2783);
xor U2936 (N_2936,N_2873,N_2853);
xor U2937 (N_2937,N_2867,N_2861);
nand U2938 (N_2938,N_2867,N_2856);
xor U2939 (N_2939,N_2830,N_2801);
xnor U2940 (N_2940,N_2845,N_2794);
nand U2941 (N_2941,N_2855,N_2801);
or U2942 (N_2942,N_2769,N_2863);
or U2943 (N_2943,N_2811,N_2852);
nand U2944 (N_2944,N_2821,N_2750);
or U2945 (N_2945,N_2823,N_2781);
nand U2946 (N_2946,N_2780,N_2801);
and U2947 (N_2947,N_2859,N_2763);
or U2948 (N_2948,N_2784,N_2815);
or U2949 (N_2949,N_2867,N_2824);
or U2950 (N_2950,N_2843,N_2874);
and U2951 (N_2951,N_2826,N_2769);
nand U2952 (N_2952,N_2771,N_2789);
nand U2953 (N_2953,N_2844,N_2776);
and U2954 (N_2954,N_2852,N_2791);
nand U2955 (N_2955,N_2795,N_2756);
and U2956 (N_2956,N_2780,N_2765);
or U2957 (N_2957,N_2871,N_2820);
or U2958 (N_2958,N_2799,N_2814);
xnor U2959 (N_2959,N_2808,N_2831);
and U2960 (N_2960,N_2862,N_2824);
or U2961 (N_2961,N_2825,N_2845);
xor U2962 (N_2962,N_2815,N_2750);
and U2963 (N_2963,N_2766,N_2829);
xor U2964 (N_2964,N_2766,N_2796);
and U2965 (N_2965,N_2837,N_2852);
or U2966 (N_2966,N_2854,N_2847);
and U2967 (N_2967,N_2797,N_2816);
xor U2968 (N_2968,N_2848,N_2776);
xor U2969 (N_2969,N_2802,N_2844);
nor U2970 (N_2970,N_2768,N_2822);
or U2971 (N_2971,N_2754,N_2795);
nor U2972 (N_2972,N_2785,N_2777);
and U2973 (N_2973,N_2850,N_2870);
nand U2974 (N_2974,N_2827,N_2801);
or U2975 (N_2975,N_2819,N_2806);
nand U2976 (N_2976,N_2807,N_2798);
or U2977 (N_2977,N_2811,N_2828);
nor U2978 (N_2978,N_2842,N_2751);
and U2979 (N_2979,N_2763,N_2815);
nor U2980 (N_2980,N_2773,N_2756);
nand U2981 (N_2981,N_2826,N_2871);
or U2982 (N_2982,N_2815,N_2814);
or U2983 (N_2983,N_2864,N_2835);
and U2984 (N_2984,N_2754,N_2847);
nor U2985 (N_2985,N_2812,N_2813);
and U2986 (N_2986,N_2834,N_2788);
or U2987 (N_2987,N_2776,N_2829);
nor U2988 (N_2988,N_2830,N_2853);
xnor U2989 (N_2989,N_2782,N_2874);
xnor U2990 (N_2990,N_2848,N_2784);
nand U2991 (N_2991,N_2840,N_2760);
and U2992 (N_2992,N_2850,N_2805);
nand U2993 (N_2993,N_2796,N_2851);
xor U2994 (N_2994,N_2870,N_2806);
and U2995 (N_2995,N_2831,N_2806);
nand U2996 (N_2996,N_2840,N_2786);
and U2997 (N_2997,N_2757,N_2860);
and U2998 (N_2998,N_2767,N_2871);
xor U2999 (N_2999,N_2764,N_2807);
or U3000 (N_3000,N_2892,N_2997);
or U3001 (N_3001,N_2917,N_2896);
nor U3002 (N_3002,N_2991,N_2891);
nand U3003 (N_3003,N_2921,N_2918);
nor U3004 (N_3004,N_2937,N_2899);
or U3005 (N_3005,N_2898,N_2967);
and U3006 (N_3006,N_2875,N_2876);
nand U3007 (N_3007,N_2999,N_2959);
and U3008 (N_3008,N_2882,N_2878);
and U3009 (N_3009,N_2877,N_2982);
nor U3010 (N_3010,N_2912,N_2950);
nand U3011 (N_3011,N_2890,N_2975);
xor U3012 (N_3012,N_2985,N_2961);
xnor U3013 (N_3013,N_2998,N_2910);
and U3014 (N_3014,N_2993,N_2879);
and U3015 (N_3015,N_2954,N_2940);
or U3016 (N_3016,N_2971,N_2949);
and U3017 (N_3017,N_2939,N_2972);
or U3018 (N_3018,N_2907,N_2911);
or U3019 (N_3019,N_2955,N_2938);
nand U3020 (N_3020,N_2984,N_2893);
or U3021 (N_3021,N_2969,N_2909);
xor U3022 (N_3022,N_2958,N_2887);
nor U3023 (N_3023,N_2953,N_2885);
nor U3024 (N_3024,N_2988,N_2915);
nor U3025 (N_3025,N_2995,N_2884);
nand U3026 (N_3026,N_2904,N_2978);
and U3027 (N_3027,N_2943,N_2928);
or U3028 (N_3028,N_2895,N_2990);
xor U3029 (N_3029,N_2880,N_2960);
nand U3030 (N_3030,N_2916,N_2944);
and U3031 (N_3031,N_2962,N_2930);
and U3032 (N_3032,N_2996,N_2946);
nor U3033 (N_3033,N_2957,N_2966);
nor U3034 (N_3034,N_2901,N_2926);
xor U3035 (N_3035,N_2888,N_2968);
or U3036 (N_3036,N_2900,N_2963);
and U3037 (N_3037,N_2986,N_2932);
xor U3038 (N_3038,N_2886,N_2894);
and U3039 (N_3039,N_2977,N_2934);
nor U3040 (N_3040,N_2948,N_2994);
or U3041 (N_3041,N_2914,N_2906);
nand U3042 (N_3042,N_2925,N_2951);
nor U3043 (N_3043,N_2987,N_2942);
or U3044 (N_3044,N_2945,N_2883);
and U3045 (N_3045,N_2933,N_2931);
and U3046 (N_3046,N_2920,N_2923);
or U3047 (N_3047,N_2980,N_2889);
xnor U3048 (N_3048,N_2924,N_2956);
xor U3049 (N_3049,N_2974,N_2970);
nor U3050 (N_3050,N_2952,N_2941);
and U3051 (N_3051,N_2964,N_2947);
and U3052 (N_3052,N_2903,N_2913);
and U3053 (N_3053,N_2935,N_2922);
and U3054 (N_3054,N_2908,N_2992);
nor U3055 (N_3055,N_2976,N_2983);
xor U3056 (N_3056,N_2905,N_2919);
xor U3057 (N_3057,N_2897,N_2979);
or U3058 (N_3058,N_2973,N_2936);
nor U3059 (N_3059,N_2981,N_2927);
nor U3060 (N_3060,N_2989,N_2881);
xor U3061 (N_3061,N_2929,N_2902);
and U3062 (N_3062,N_2965,N_2879);
or U3063 (N_3063,N_2945,N_2908);
nand U3064 (N_3064,N_2932,N_2994);
xnor U3065 (N_3065,N_2946,N_2969);
or U3066 (N_3066,N_2891,N_2964);
and U3067 (N_3067,N_2966,N_2953);
nand U3068 (N_3068,N_2901,N_2976);
nand U3069 (N_3069,N_2998,N_2956);
xnor U3070 (N_3070,N_2983,N_2919);
xnor U3071 (N_3071,N_2879,N_2892);
or U3072 (N_3072,N_2932,N_2910);
xor U3073 (N_3073,N_2959,N_2920);
and U3074 (N_3074,N_2929,N_2913);
or U3075 (N_3075,N_2938,N_2897);
and U3076 (N_3076,N_2986,N_2889);
or U3077 (N_3077,N_2929,N_2983);
nand U3078 (N_3078,N_2922,N_2912);
nand U3079 (N_3079,N_2986,N_2881);
or U3080 (N_3080,N_2997,N_2898);
and U3081 (N_3081,N_2887,N_2876);
or U3082 (N_3082,N_2978,N_2898);
nor U3083 (N_3083,N_2968,N_2944);
nand U3084 (N_3084,N_2946,N_2989);
and U3085 (N_3085,N_2880,N_2887);
nor U3086 (N_3086,N_2996,N_2941);
or U3087 (N_3087,N_2969,N_2902);
or U3088 (N_3088,N_2898,N_2927);
nand U3089 (N_3089,N_2908,N_2980);
nor U3090 (N_3090,N_2953,N_2880);
and U3091 (N_3091,N_2958,N_2919);
and U3092 (N_3092,N_2959,N_2876);
xnor U3093 (N_3093,N_2957,N_2947);
nor U3094 (N_3094,N_2896,N_2930);
or U3095 (N_3095,N_2969,N_2949);
or U3096 (N_3096,N_2949,N_2931);
and U3097 (N_3097,N_2918,N_2992);
and U3098 (N_3098,N_2898,N_2928);
and U3099 (N_3099,N_2899,N_2942);
nor U3100 (N_3100,N_2929,N_2948);
and U3101 (N_3101,N_2960,N_2945);
and U3102 (N_3102,N_2958,N_2895);
xor U3103 (N_3103,N_2916,N_2903);
nor U3104 (N_3104,N_2889,N_2963);
nand U3105 (N_3105,N_2990,N_2979);
xor U3106 (N_3106,N_2905,N_2930);
nand U3107 (N_3107,N_2929,N_2926);
and U3108 (N_3108,N_2948,N_2925);
nor U3109 (N_3109,N_2984,N_2949);
and U3110 (N_3110,N_2883,N_2895);
xor U3111 (N_3111,N_2947,N_2962);
nor U3112 (N_3112,N_2919,N_2956);
nand U3113 (N_3113,N_2875,N_2994);
nor U3114 (N_3114,N_2904,N_2964);
xor U3115 (N_3115,N_2940,N_2899);
or U3116 (N_3116,N_2999,N_2894);
and U3117 (N_3117,N_2972,N_2953);
and U3118 (N_3118,N_2985,N_2966);
nor U3119 (N_3119,N_2956,N_2954);
or U3120 (N_3120,N_2939,N_2962);
nor U3121 (N_3121,N_2953,N_2991);
nor U3122 (N_3122,N_2953,N_2896);
nor U3123 (N_3123,N_2887,N_2899);
and U3124 (N_3124,N_2947,N_2921);
or U3125 (N_3125,N_3086,N_3012);
or U3126 (N_3126,N_3024,N_3082);
nand U3127 (N_3127,N_3075,N_3107);
and U3128 (N_3128,N_3043,N_3027);
or U3129 (N_3129,N_3115,N_3039);
or U3130 (N_3130,N_3041,N_3080);
xor U3131 (N_3131,N_3083,N_3035);
and U3132 (N_3132,N_3100,N_3023);
or U3133 (N_3133,N_3051,N_3111);
or U3134 (N_3134,N_3077,N_3009);
nor U3135 (N_3135,N_3014,N_3010);
and U3136 (N_3136,N_3029,N_3050);
and U3137 (N_3137,N_3017,N_3076);
xor U3138 (N_3138,N_3070,N_3113);
nor U3139 (N_3139,N_3072,N_3047);
and U3140 (N_3140,N_3019,N_3096);
xnor U3141 (N_3141,N_3015,N_3011);
or U3142 (N_3142,N_3102,N_3025);
nand U3143 (N_3143,N_3109,N_3042);
or U3144 (N_3144,N_3053,N_3104);
xnor U3145 (N_3145,N_3001,N_3002);
and U3146 (N_3146,N_3000,N_3006);
or U3147 (N_3147,N_3062,N_3037);
nor U3148 (N_3148,N_3094,N_3044);
nand U3149 (N_3149,N_3112,N_3033);
xor U3150 (N_3150,N_3088,N_3048);
or U3151 (N_3151,N_3065,N_3097);
nor U3152 (N_3152,N_3060,N_3058);
xor U3153 (N_3153,N_3118,N_3038);
or U3154 (N_3154,N_3028,N_3067);
and U3155 (N_3155,N_3055,N_3124);
nor U3156 (N_3156,N_3101,N_3008);
xnor U3157 (N_3157,N_3061,N_3056);
or U3158 (N_3158,N_3030,N_3081);
nand U3159 (N_3159,N_3117,N_3103);
nand U3160 (N_3160,N_3049,N_3022);
nand U3161 (N_3161,N_3040,N_3007);
nor U3162 (N_3162,N_3016,N_3123);
nor U3163 (N_3163,N_3046,N_3093);
xnor U3164 (N_3164,N_3071,N_3106);
or U3165 (N_3165,N_3021,N_3066);
nor U3166 (N_3166,N_3026,N_3089);
and U3167 (N_3167,N_3045,N_3069);
nor U3168 (N_3168,N_3078,N_3090);
nor U3169 (N_3169,N_3087,N_3074);
nand U3170 (N_3170,N_3036,N_3110);
nand U3171 (N_3171,N_3108,N_3003);
or U3172 (N_3172,N_3098,N_3005);
nor U3173 (N_3173,N_3095,N_3120);
or U3174 (N_3174,N_3079,N_3092);
and U3175 (N_3175,N_3116,N_3032);
and U3176 (N_3176,N_3052,N_3091);
nand U3177 (N_3177,N_3114,N_3057);
nor U3178 (N_3178,N_3084,N_3013);
and U3179 (N_3179,N_3018,N_3034);
nor U3180 (N_3180,N_3099,N_3105);
xor U3181 (N_3181,N_3004,N_3059);
nand U3182 (N_3182,N_3085,N_3064);
nor U3183 (N_3183,N_3031,N_3121);
and U3184 (N_3184,N_3119,N_3122);
nor U3185 (N_3185,N_3063,N_3054);
xor U3186 (N_3186,N_3020,N_3068);
xnor U3187 (N_3187,N_3073,N_3050);
or U3188 (N_3188,N_3103,N_3105);
xnor U3189 (N_3189,N_3044,N_3026);
or U3190 (N_3190,N_3037,N_3013);
nand U3191 (N_3191,N_3086,N_3101);
nor U3192 (N_3192,N_3103,N_3096);
or U3193 (N_3193,N_3111,N_3050);
xnor U3194 (N_3194,N_3110,N_3075);
xnor U3195 (N_3195,N_3061,N_3062);
xnor U3196 (N_3196,N_3097,N_3018);
xnor U3197 (N_3197,N_3017,N_3106);
nand U3198 (N_3198,N_3037,N_3020);
or U3199 (N_3199,N_3065,N_3062);
or U3200 (N_3200,N_3084,N_3067);
or U3201 (N_3201,N_3043,N_3050);
or U3202 (N_3202,N_3025,N_3108);
nor U3203 (N_3203,N_3089,N_3122);
or U3204 (N_3204,N_3079,N_3027);
xnor U3205 (N_3205,N_3113,N_3012);
or U3206 (N_3206,N_3086,N_3095);
and U3207 (N_3207,N_3062,N_3049);
nand U3208 (N_3208,N_3011,N_3012);
and U3209 (N_3209,N_3084,N_3033);
nor U3210 (N_3210,N_3029,N_3079);
nand U3211 (N_3211,N_3106,N_3062);
and U3212 (N_3212,N_3000,N_3015);
nand U3213 (N_3213,N_3090,N_3020);
xor U3214 (N_3214,N_3014,N_3069);
xor U3215 (N_3215,N_3061,N_3047);
xor U3216 (N_3216,N_3006,N_3041);
or U3217 (N_3217,N_3080,N_3102);
nor U3218 (N_3218,N_3094,N_3085);
nor U3219 (N_3219,N_3034,N_3067);
or U3220 (N_3220,N_3088,N_3031);
xor U3221 (N_3221,N_3100,N_3071);
and U3222 (N_3222,N_3099,N_3038);
and U3223 (N_3223,N_3097,N_3112);
xor U3224 (N_3224,N_3074,N_3039);
xnor U3225 (N_3225,N_3058,N_3009);
and U3226 (N_3226,N_3035,N_3059);
nor U3227 (N_3227,N_3064,N_3034);
or U3228 (N_3228,N_3036,N_3082);
nand U3229 (N_3229,N_3065,N_3107);
and U3230 (N_3230,N_3074,N_3023);
or U3231 (N_3231,N_3015,N_3124);
nor U3232 (N_3232,N_3077,N_3119);
and U3233 (N_3233,N_3029,N_3098);
xor U3234 (N_3234,N_3120,N_3054);
nand U3235 (N_3235,N_3038,N_3074);
nand U3236 (N_3236,N_3084,N_3110);
nand U3237 (N_3237,N_3104,N_3102);
xor U3238 (N_3238,N_3083,N_3026);
nand U3239 (N_3239,N_3111,N_3102);
xnor U3240 (N_3240,N_3116,N_3012);
nor U3241 (N_3241,N_3024,N_3030);
and U3242 (N_3242,N_3012,N_3064);
xnor U3243 (N_3243,N_3115,N_3017);
or U3244 (N_3244,N_3023,N_3091);
nor U3245 (N_3245,N_3122,N_3080);
or U3246 (N_3246,N_3041,N_3073);
nand U3247 (N_3247,N_3069,N_3040);
nor U3248 (N_3248,N_3076,N_3092);
nand U3249 (N_3249,N_3063,N_3017);
xnor U3250 (N_3250,N_3159,N_3172);
nand U3251 (N_3251,N_3177,N_3187);
and U3252 (N_3252,N_3248,N_3232);
or U3253 (N_3253,N_3174,N_3161);
and U3254 (N_3254,N_3238,N_3203);
and U3255 (N_3255,N_3202,N_3144);
or U3256 (N_3256,N_3240,N_3222);
or U3257 (N_3257,N_3169,N_3227);
nor U3258 (N_3258,N_3181,N_3244);
nand U3259 (N_3259,N_3197,N_3148);
and U3260 (N_3260,N_3241,N_3193);
xnor U3261 (N_3261,N_3237,N_3182);
and U3262 (N_3262,N_3180,N_3143);
and U3263 (N_3263,N_3206,N_3243);
xnor U3264 (N_3264,N_3175,N_3171);
nor U3265 (N_3265,N_3200,N_3249);
nand U3266 (N_3266,N_3208,N_3163);
and U3267 (N_3267,N_3166,N_3225);
nor U3268 (N_3268,N_3155,N_3145);
or U3269 (N_3269,N_3167,N_3191);
nor U3270 (N_3270,N_3242,N_3195);
nand U3271 (N_3271,N_3160,N_3224);
nand U3272 (N_3272,N_3186,N_3216);
or U3273 (N_3273,N_3127,N_3136);
and U3274 (N_3274,N_3233,N_3135);
nor U3275 (N_3275,N_3134,N_3150);
xnor U3276 (N_3276,N_3185,N_3207);
nor U3277 (N_3277,N_3176,N_3140);
xnor U3278 (N_3278,N_3178,N_3146);
and U3279 (N_3279,N_3183,N_3162);
xnor U3280 (N_3280,N_3139,N_3215);
or U3281 (N_3281,N_3219,N_3211);
xnor U3282 (N_3282,N_3198,N_3130);
or U3283 (N_3283,N_3129,N_3151);
nor U3284 (N_3284,N_3190,N_3126);
nand U3285 (N_3285,N_3137,N_3131);
xnor U3286 (N_3286,N_3170,N_3141);
nor U3287 (N_3287,N_3205,N_3223);
nand U3288 (N_3288,N_3165,N_3231);
nor U3289 (N_3289,N_3184,N_3210);
and U3290 (N_3290,N_3218,N_3152);
or U3291 (N_3291,N_3194,N_3246);
nor U3292 (N_3292,N_3201,N_3221);
xor U3293 (N_3293,N_3236,N_3247);
or U3294 (N_3294,N_3153,N_3128);
and U3295 (N_3295,N_3204,N_3196);
xnor U3296 (N_3296,N_3228,N_3212);
nand U3297 (N_3297,N_3230,N_3179);
nand U3298 (N_3298,N_3125,N_3188);
or U3299 (N_3299,N_3213,N_3217);
or U3300 (N_3300,N_3142,N_3189);
nor U3301 (N_3301,N_3235,N_3192);
nand U3302 (N_3302,N_3154,N_3199);
xnor U3303 (N_3303,N_3164,N_3220);
nor U3304 (N_3304,N_3226,N_3229);
or U3305 (N_3305,N_3138,N_3209);
nor U3306 (N_3306,N_3157,N_3245);
and U3307 (N_3307,N_3173,N_3133);
and U3308 (N_3308,N_3156,N_3149);
or U3309 (N_3309,N_3168,N_3234);
nand U3310 (N_3310,N_3239,N_3147);
nand U3311 (N_3311,N_3214,N_3132);
nor U3312 (N_3312,N_3158,N_3139);
and U3313 (N_3313,N_3220,N_3135);
and U3314 (N_3314,N_3178,N_3150);
and U3315 (N_3315,N_3228,N_3129);
or U3316 (N_3316,N_3186,N_3203);
or U3317 (N_3317,N_3249,N_3196);
nand U3318 (N_3318,N_3131,N_3194);
or U3319 (N_3319,N_3189,N_3126);
nor U3320 (N_3320,N_3128,N_3203);
xnor U3321 (N_3321,N_3157,N_3242);
nand U3322 (N_3322,N_3194,N_3160);
nor U3323 (N_3323,N_3221,N_3199);
or U3324 (N_3324,N_3223,N_3225);
or U3325 (N_3325,N_3231,N_3211);
nand U3326 (N_3326,N_3206,N_3152);
or U3327 (N_3327,N_3185,N_3214);
xor U3328 (N_3328,N_3160,N_3211);
or U3329 (N_3329,N_3169,N_3127);
xnor U3330 (N_3330,N_3150,N_3228);
nand U3331 (N_3331,N_3125,N_3202);
nand U3332 (N_3332,N_3245,N_3199);
and U3333 (N_3333,N_3238,N_3157);
nand U3334 (N_3334,N_3129,N_3131);
nor U3335 (N_3335,N_3136,N_3154);
nand U3336 (N_3336,N_3147,N_3229);
and U3337 (N_3337,N_3225,N_3142);
xor U3338 (N_3338,N_3230,N_3212);
or U3339 (N_3339,N_3217,N_3214);
nor U3340 (N_3340,N_3170,N_3201);
nor U3341 (N_3341,N_3214,N_3134);
nor U3342 (N_3342,N_3164,N_3245);
or U3343 (N_3343,N_3146,N_3160);
or U3344 (N_3344,N_3213,N_3241);
nor U3345 (N_3345,N_3190,N_3169);
xnor U3346 (N_3346,N_3187,N_3194);
and U3347 (N_3347,N_3247,N_3144);
and U3348 (N_3348,N_3191,N_3187);
or U3349 (N_3349,N_3193,N_3136);
and U3350 (N_3350,N_3146,N_3129);
and U3351 (N_3351,N_3226,N_3131);
nor U3352 (N_3352,N_3143,N_3230);
nand U3353 (N_3353,N_3212,N_3174);
xor U3354 (N_3354,N_3249,N_3248);
and U3355 (N_3355,N_3204,N_3127);
nor U3356 (N_3356,N_3143,N_3156);
nand U3357 (N_3357,N_3140,N_3175);
nor U3358 (N_3358,N_3207,N_3125);
xnor U3359 (N_3359,N_3141,N_3199);
xnor U3360 (N_3360,N_3217,N_3181);
xor U3361 (N_3361,N_3206,N_3192);
nand U3362 (N_3362,N_3223,N_3125);
nor U3363 (N_3363,N_3178,N_3241);
xnor U3364 (N_3364,N_3157,N_3138);
xor U3365 (N_3365,N_3172,N_3137);
xnor U3366 (N_3366,N_3145,N_3218);
nand U3367 (N_3367,N_3128,N_3168);
and U3368 (N_3368,N_3190,N_3179);
nand U3369 (N_3369,N_3149,N_3215);
nand U3370 (N_3370,N_3220,N_3181);
nor U3371 (N_3371,N_3242,N_3133);
or U3372 (N_3372,N_3210,N_3162);
or U3373 (N_3373,N_3167,N_3169);
nand U3374 (N_3374,N_3142,N_3140);
or U3375 (N_3375,N_3352,N_3288);
nand U3376 (N_3376,N_3369,N_3319);
xor U3377 (N_3377,N_3254,N_3356);
xnor U3378 (N_3378,N_3342,N_3373);
or U3379 (N_3379,N_3338,N_3370);
xnor U3380 (N_3380,N_3297,N_3348);
nand U3381 (N_3381,N_3295,N_3326);
or U3382 (N_3382,N_3306,N_3327);
xnor U3383 (N_3383,N_3349,N_3325);
and U3384 (N_3384,N_3262,N_3331);
and U3385 (N_3385,N_3362,N_3263);
nand U3386 (N_3386,N_3276,N_3293);
and U3387 (N_3387,N_3323,N_3301);
or U3388 (N_3388,N_3258,N_3272);
and U3389 (N_3389,N_3266,N_3360);
xor U3390 (N_3390,N_3343,N_3279);
or U3391 (N_3391,N_3336,N_3332);
or U3392 (N_3392,N_3282,N_3318);
xor U3393 (N_3393,N_3269,N_3291);
or U3394 (N_3394,N_3265,N_3341);
or U3395 (N_3395,N_3366,N_3310);
nand U3396 (N_3396,N_3251,N_3355);
or U3397 (N_3397,N_3294,N_3328);
xor U3398 (N_3398,N_3273,N_3344);
and U3399 (N_3399,N_3299,N_3371);
nor U3400 (N_3400,N_3340,N_3312);
nand U3401 (N_3401,N_3302,N_3309);
nor U3402 (N_3402,N_3361,N_3322);
and U3403 (N_3403,N_3284,N_3281);
nand U3404 (N_3404,N_3314,N_3256);
nor U3405 (N_3405,N_3353,N_3285);
nor U3406 (N_3406,N_3365,N_3320);
nand U3407 (N_3407,N_3252,N_3317);
nand U3408 (N_3408,N_3283,N_3303);
and U3409 (N_3409,N_3290,N_3267);
and U3410 (N_3410,N_3358,N_3307);
nor U3411 (N_3411,N_3354,N_3337);
xnor U3412 (N_3412,N_3300,N_3333);
xor U3413 (N_3413,N_3261,N_3286);
nor U3414 (N_3414,N_3334,N_3270);
nor U3415 (N_3415,N_3330,N_3374);
or U3416 (N_3416,N_3316,N_3304);
nand U3417 (N_3417,N_3367,N_3324);
nor U3418 (N_3418,N_3305,N_3308);
or U3419 (N_3419,N_3274,N_3257);
and U3420 (N_3420,N_3298,N_3347);
xor U3421 (N_3421,N_3264,N_3345);
nand U3422 (N_3422,N_3315,N_3271);
nand U3423 (N_3423,N_3357,N_3280);
nand U3424 (N_3424,N_3255,N_3260);
nor U3425 (N_3425,N_3268,N_3350);
xor U3426 (N_3426,N_3296,N_3313);
xor U3427 (N_3427,N_3329,N_3292);
and U3428 (N_3428,N_3351,N_3368);
and U3429 (N_3429,N_3311,N_3287);
and U3430 (N_3430,N_3335,N_3278);
and U3431 (N_3431,N_3364,N_3275);
and U3432 (N_3432,N_3259,N_3277);
and U3433 (N_3433,N_3250,N_3253);
and U3434 (N_3434,N_3346,N_3321);
nand U3435 (N_3435,N_3359,N_3372);
nor U3436 (N_3436,N_3363,N_3339);
nor U3437 (N_3437,N_3289,N_3328);
nand U3438 (N_3438,N_3314,N_3305);
or U3439 (N_3439,N_3348,N_3290);
nand U3440 (N_3440,N_3301,N_3277);
nor U3441 (N_3441,N_3326,N_3322);
nor U3442 (N_3442,N_3326,N_3351);
or U3443 (N_3443,N_3305,N_3335);
nand U3444 (N_3444,N_3298,N_3305);
nor U3445 (N_3445,N_3328,N_3315);
and U3446 (N_3446,N_3341,N_3266);
nand U3447 (N_3447,N_3252,N_3307);
and U3448 (N_3448,N_3332,N_3300);
nand U3449 (N_3449,N_3292,N_3320);
nand U3450 (N_3450,N_3307,N_3373);
and U3451 (N_3451,N_3372,N_3365);
xnor U3452 (N_3452,N_3276,N_3306);
nor U3453 (N_3453,N_3273,N_3362);
or U3454 (N_3454,N_3271,N_3302);
xnor U3455 (N_3455,N_3253,N_3289);
or U3456 (N_3456,N_3302,N_3272);
nor U3457 (N_3457,N_3265,N_3358);
nand U3458 (N_3458,N_3284,N_3315);
nor U3459 (N_3459,N_3266,N_3265);
nand U3460 (N_3460,N_3322,N_3332);
and U3461 (N_3461,N_3273,N_3269);
nor U3462 (N_3462,N_3270,N_3305);
or U3463 (N_3463,N_3359,N_3374);
nor U3464 (N_3464,N_3299,N_3359);
nor U3465 (N_3465,N_3272,N_3352);
nor U3466 (N_3466,N_3355,N_3260);
and U3467 (N_3467,N_3330,N_3323);
nor U3468 (N_3468,N_3299,N_3368);
nor U3469 (N_3469,N_3358,N_3309);
and U3470 (N_3470,N_3289,N_3354);
or U3471 (N_3471,N_3252,N_3326);
nand U3472 (N_3472,N_3295,N_3300);
nor U3473 (N_3473,N_3315,N_3281);
nand U3474 (N_3474,N_3286,N_3354);
nand U3475 (N_3475,N_3254,N_3262);
and U3476 (N_3476,N_3297,N_3271);
and U3477 (N_3477,N_3289,N_3286);
or U3478 (N_3478,N_3277,N_3273);
xor U3479 (N_3479,N_3265,N_3259);
and U3480 (N_3480,N_3321,N_3326);
or U3481 (N_3481,N_3309,N_3368);
nor U3482 (N_3482,N_3250,N_3314);
xor U3483 (N_3483,N_3320,N_3339);
or U3484 (N_3484,N_3344,N_3263);
or U3485 (N_3485,N_3255,N_3291);
and U3486 (N_3486,N_3356,N_3288);
nor U3487 (N_3487,N_3302,N_3316);
or U3488 (N_3488,N_3356,N_3281);
xnor U3489 (N_3489,N_3285,N_3348);
nor U3490 (N_3490,N_3291,N_3359);
nor U3491 (N_3491,N_3307,N_3308);
nor U3492 (N_3492,N_3295,N_3252);
nor U3493 (N_3493,N_3297,N_3329);
nand U3494 (N_3494,N_3276,N_3321);
or U3495 (N_3495,N_3325,N_3305);
nor U3496 (N_3496,N_3255,N_3264);
nand U3497 (N_3497,N_3313,N_3310);
xnor U3498 (N_3498,N_3368,N_3372);
nand U3499 (N_3499,N_3283,N_3349);
xor U3500 (N_3500,N_3437,N_3492);
nor U3501 (N_3501,N_3440,N_3409);
nor U3502 (N_3502,N_3491,N_3399);
nor U3503 (N_3503,N_3468,N_3490);
nand U3504 (N_3504,N_3484,N_3417);
or U3505 (N_3505,N_3442,N_3434);
nor U3506 (N_3506,N_3480,N_3385);
nor U3507 (N_3507,N_3404,N_3498);
or U3508 (N_3508,N_3470,N_3455);
nor U3509 (N_3509,N_3378,N_3405);
nand U3510 (N_3510,N_3389,N_3446);
xnor U3511 (N_3511,N_3392,N_3375);
and U3512 (N_3512,N_3493,N_3412);
and U3513 (N_3513,N_3471,N_3431);
nand U3514 (N_3514,N_3406,N_3384);
or U3515 (N_3515,N_3423,N_3380);
nand U3516 (N_3516,N_3487,N_3407);
nand U3517 (N_3517,N_3459,N_3425);
nand U3518 (N_3518,N_3450,N_3388);
and U3519 (N_3519,N_3411,N_3383);
xnor U3520 (N_3520,N_3394,N_3447);
and U3521 (N_3521,N_3415,N_3466);
nand U3522 (N_3522,N_3419,N_3410);
and U3523 (N_3523,N_3427,N_3441);
and U3524 (N_3524,N_3390,N_3432);
nand U3525 (N_3525,N_3454,N_3452);
xor U3526 (N_3526,N_3472,N_3489);
nor U3527 (N_3527,N_3496,N_3474);
xnor U3528 (N_3528,N_3396,N_3398);
nor U3529 (N_3529,N_3403,N_3485);
xor U3530 (N_3530,N_3397,N_3462);
and U3531 (N_3531,N_3444,N_3475);
xnor U3532 (N_3532,N_3435,N_3458);
or U3533 (N_3533,N_3488,N_3426);
or U3534 (N_3534,N_3486,N_3457);
or U3535 (N_3535,N_3387,N_3408);
xnor U3536 (N_3536,N_3386,N_3393);
and U3537 (N_3537,N_3478,N_3422);
or U3538 (N_3538,N_3479,N_3449);
or U3539 (N_3539,N_3461,N_3456);
nand U3540 (N_3540,N_3420,N_3428);
nand U3541 (N_3541,N_3418,N_3443);
nor U3542 (N_3542,N_3453,N_3413);
xor U3543 (N_3543,N_3433,N_3483);
and U3544 (N_3544,N_3451,N_3379);
and U3545 (N_3545,N_3382,N_3414);
or U3546 (N_3546,N_3381,N_3469);
xor U3547 (N_3547,N_3429,N_3445);
and U3548 (N_3548,N_3430,N_3402);
nand U3549 (N_3549,N_3497,N_3436);
xnor U3550 (N_3550,N_3424,N_3463);
nor U3551 (N_3551,N_3421,N_3416);
nand U3552 (N_3552,N_3395,N_3439);
nor U3553 (N_3553,N_3464,N_3401);
or U3554 (N_3554,N_3476,N_3376);
nor U3555 (N_3555,N_3377,N_3477);
xor U3556 (N_3556,N_3400,N_3499);
nor U3557 (N_3557,N_3448,N_3460);
or U3558 (N_3558,N_3438,N_3391);
nor U3559 (N_3559,N_3473,N_3495);
or U3560 (N_3560,N_3467,N_3482);
or U3561 (N_3561,N_3465,N_3481);
and U3562 (N_3562,N_3494,N_3395);
and U3563 (N_3563,N_3485,N_3399);
xnor U3564 (N_3564,N_3437,N_3473);
xor U3565 (N_3565,N_3412,N_3391);
or U3566 (N_3566,N_3498,N_3490);
or U3567 (N_3567,N_3438,N_3383);
nand U3568 (N_3568,N_3454,N_3480);
and U3569 (N_3569,N_3433,N_3391);
or U3570 (N_3570,N_3393,N_3424);
or U3571 (N_3571,N_3480,N_3400);
nor U3572 (N_3572,N_3393,N_3475);
and U3573 (N_3573,N_3413,N_3465);
and U3574 (N_3574,N_3478,N_3398);
xnor U3575 (N_3575,N_3404,N_3476);
xnor U3576 (N_3576,N_3387,N_3482);
xor U3577 (N_3577,N_3422,N_3448);
or U3578 (N_3578,N_3454,N_3402);
or U3579 (N_3579,N_3446,N_3413);
or U3580 (N_3580,N_3377,N_3408);
nor U3581 (N_3581,N_3384,N_3434);
xnor U3582 (N_3582,N_3465,N_3496);
or U3583 (N_3583,N_3438,N_3416);
and U3584 (N_3584,N_3482,N_3494);
or U3585 (N_3585,N_3486,N_3440);
xor U3586 (N_3586,N_3453,N_3481);
or U3587 (N_3587,N_3391,N_3451);
and U3588 (N_3588,N_3399,N_3493);
nand U3589 (N_3589,N_3440,N_3495);
xnor U3590 (N_3590,N_3433,N_3437);
xor U3591 (N_3591,N_3449,N_3375);
and U3592 (N_3592,N_3486,N_3472);
nand U3593 (N_3593,N_3470,N_3392);
nand U3594 (N_3594,N_3415,N_3481);
nand U3595 (N_3595,N_3474,N_3479);
nor U3596 (N_3596,N_3453,N_3472);
and U3597 (N_3597,N_3413,N_3474);
nor U3598 (N_3598,N_3379,N_3487);
xor U3599 (N_3599,N_3459,N_3439);
nand U3600 (N_3600,N_3410,N_3402);
and U3601 (N_3601,N_3382,N_3418);
nand U3602 (N_3602,N_3485,N_3458);
xor U3603 (N_3603,N_3380,N_3470);
xor U3604 (N_3604,N_3407,N_3422);
nand U3605 (N_3605,N_3434,N_3476);
nor U3606 (N_3606,N_3497,N_3441);
nor U3607 (N_3607,N_3408,N_3446);
nand U3608 (N_3608,N_3434,N_3474);
xor U3609 (N_3609,N_3450,N_3408);
nand U3610 (N_3610,N_3494,N_3375);
or U3611 (N_3611,N_3446,N_3387);
and U3612 (N_3612,N_3488,N_3385);
nand U3613 (N_3613,N_3496,N_3414);
nand U3614 (N_3614,N_3436,N_3402);
xor U3615 (N_3615,N_3450,N_3465);
nor U3616 (N_3616,N_3405,N_3402);
nand U3617 (N_3617,N_3390,N_3386);
and U3618 (N_3618,N_3379,N_3480);
and U3619 (N_3619,N_3375,N_3381);
nand U3620 (N_3620,N_3438,N_3425);
nor U3621 (N_3621,N_3430,N_3472);
xnor U3622 (N_3622,N_3417,N_3495);
nor U3623 (N_3623,N_3454,N_3434);
nand U3624 (N_3624,N_3418,N_3470);
or U3625 (N_3625,N_3585,N_3508);
and U3626 (N_3626,N_3504,N_3612);
nand U3627 (N_3627,N_3507,N_3544);
nand U3628 (N_3628,N_3588,N_3606);
nor U3629 (N_3629,N_3522,N_3571);
and U3630 (N_3630,N_3514,N_3624);
xor U3631 (N_3631,N_3564,N_3524);
xor U3632 (N_3632,N_3583,N_3569);
nor U3633 (N_3633,N_3578,N_3611);
xnor U3634 (N_3634,N_3515,N_3609);
nand U3635 (N_3635,N_3566,N_3584);
xnor U3636 (N_3636,N_3586,N_3505);
nor U3637 (N_3637,N_3556,N_3502);
nor U3638 (N_3638,N_3558,N_3528);
nand U3639 (N_3639,N_3577,N_3595);
nor U3640 (N_3640,N_3517,N_3562);
and U3641 (N_3641,N_3597,N_3533);
nor U3642 (N_3642,N_3621,N_3529);
and U3643 (N_3643,N_3518,N_3538);
or U3644 (N_3644,N_3548,N_3525);
nor U3645 (N_3645,N_3570,N_3536);
nand U3646 (N_3646,N_3531,N_3557);
nand U3647 (N_3647,N_3589,N_3563);
or U3648 (N_3648,N_3527,N_3547);
and U3649 (N_3649,N_3576,N_3540);
xor U3650 (N_3650,N_3537,N_3512);
or U3651 (N_3651,N_3523,N_3591);
and U3652 (N_3652,N_3510,N_3511);
and U3653 (N_3653,N_3506,N_3616);
or U3654 (N_3654,N_3509,N_3605);
xor U3655 (N_3655,N_3532,N_3620);
nor U3656 (N_3656,N_3610,N_3559);
or U3657 (N_3657,N_3553,N_3615);
and U3658 (N_3658,N_3534,N_3541);
nor U3659 (N_3659,N_3618,N_3582);
xnor U3660 (N_3660,N_3617,N_3560);
xnor U3661 (N_3661,N_3604,N_3550);
and U3662 (N_3662,N_3600,N_3543);
or U3663 (N_3663,N_3542,N_3594);
nand U3664 (N_3664,N_3608,N_3539);
xnor U3665 (N_3665,N_3574,N_3521);
nand U3666 (N_3666,N_3554,N_3619);
or U3667 (N_3667,N_3551,N_3503);
nand U3668 (N_3668,N_3580,N_3519);
nor U3669 (N_3669,N_3561,N_3613);
nand U3670 (N_3670,N_3603,N_3520);
xnor U3671 (N_3671,N_3602,N_3552);
or U3672 (N_3672,N_3530,N_3607);
nor U3673 (N_3673,N_3568,N_3599);
nor U3674 (N_3674,N_3567,N_3555);
xor U3675 (N_3675,N_3593,N_3535);
nor U3676 (N_3676,N_3601,N_3596);
xnor U3677 (N_3677,N_3526,N_3572);
or U3678 (N_3678,N_3622,N_3565);
and U3679 (N_3679,N_3501,N_3581);
xor U3680 (N_3680,N_3549,N_3575);
and U3681 (N_3681,N_3516,N_3592);
and U3682 (N_3682,N_3579,N_3587);
and U3683 (N_3683,N_3573,N_3545);
and U3684 (N_3684,N_3500,N_3614);
or U3685 (N_3685,N_3590,N_3598);
xor U3686 (N_3686,N_3513,N_3623);
nand U3687 (N_3687,N_3546,N_3548);
nand U3688 (N_3688,N_3521,N_3591);
xnor U3689 (N_3689,N_3588,N_3508);
and U3690 (N_3690,N_3581,N_3535);
nor U3691 (N_3691,N_3602,N_3620);
or U3692 (N_3692,N_3593,N_3607);
nand U3693 (N_3693,N_3566,N_3535);
xor U3694 (N_3694,N_3546,N_3519);
xor U3695 (N_3695,N_3589,N_3537);
and U3696 (N_3696,N_3545,N_3515);
or U3697 (N_3697,N_3617,N_3522);
and U3698 (N_3698,N_3576,N_3559);
nand U3699 (N_3699,N_3610,N_3616);
nand U3700 (N_3700,N_3582,N_3614);
or U3701 (N_3701,N_3584,N_3561);
nand U3702 (N_3702,N_3590,N_3602);
and U3703 (N_3703,N_3581,N_3599);
nand U3704 (N_3704,N_3613,N_3576);
nor U3705 (N_3705,N_3525,N_3604);
xor U3706 (N_3706,N_3568,N_3532);
nand U3707 (N_3707,N_3609,N_3518);
nor U3708 (N_3708,N_3564,N_3609);
nor U3709 (N_3709,N_3587,N_3517);
nand U3710 (N_3710,N_3507,N_3554);
and U3711 (N_3711,N_3570,N_3554);
xnor U3712 (N_3712,N_3554,N_3603);
nand U3713 (N_3713,N_3554,N_3545);
xor U3714 (N_3714,N_3620,N_3552);
or U3715 (N_3715,N_3574,N_3538);
nor U3716 (N_3716,N_3553,N_3623);
or U3717 (N_3717,N_3561,N_3585);
xnor U3718 (N_3718,N_3549,N_3574);
xnor U3719 (N_3719,N_3529,N_3619);
or U3720 (N_3720,N_3532,N_3621);
and U3721 (N_3721,N_3565,N_3591);
nor U3722 (N_3722,N_3591,N_3588);
and U3723 (N_3723,N_3567,N_3553);
or U3724 (N_3724,N_3543,N_3560);
or U3725 (N_3725,N_3530,N_3508);
or U3726 (N_3726,N_3565,N_3612);
or U3727 (N_3727,N_3540,N_3541);
nand U3728 (N_3728,N_3595,N_3603);
and U3729 (N_3729,N_3519,N_3518);
and U3730 (N_3730,N_3501,N_3603);
nand U3731 (N_3731,N_3543,N_3522);
nor U3732 (N_3732,N_3516,N_3590);
xnor U3733 (N_3733,N_3562,N_3546);
nor U3734 (N_3734,N_3555,N_3545);
nor U3735 (N_3735,N_3524,N_3565);
or U3736 (N_3736,N_3559,N_3584);
and U3737 (N_3737,N_3504,N_3598);
or U3738 (N_3738,N_3514,N_3540);
or U3739 (N_3739,N_3579,N_3511);
xnor U3740 (N_3740,N_3623,N_3527);
xnor U3741 (N_3741,N_3512,N_3569);
and U3742 (N_3742,N_3514,N_3596);
nand U3743 (N_3743,N_3563,N_3566);
and U3744 (N_3744,N_3571,N_3601);
nor U3745 (N_3745,N_3531,N_3524);
nor U3746 (N_3746,N_3565,N_3590);
or U3747 (N_3747,N_3543,N_3552);
or U3748 (N_3748,N_3514,N_3567);
nand U3749 (N_3749,N_3588,N_3550);
nand U3750 (N_3750,N_3722,N_3682);
and U3751 (N_3751,N_3673,N_3735);
nand U3752 (N_3752,N_3630,N_3732);
or U3753 (N_3753,N_3632,N_3647);
or U3754 (N_3754,N_3748,N_3678);
and U3755 (N_3755,N_3692,N_3643);
nor U3756 (N_3756,N_3651,N_3664);
nor U3757 (N_3757,N_3729,N_3702);
xnor U3758 (N_3758,N_3652,N_3745);
nand U3759 (N_3759,N_3705,N_3718);
xor U3760 (N_3760,N_3638,N_3716);
nand U3761 (N_3761,N_3672,N_3710);
or U3762 (N_3762,N_3645,N_3746);
and U3763 (N_3763,N_3628,N_3720);
nor U3764 (N_3764,N_3626,N_3677);
nor U3765 (N_3765,N_3644,N_3742);
xnor U3766 (N_3766,N_3679,N_3658);
and U3767 (N_3767,N_3688,N_3649);
xor U3768 (N_3768,N_3723,N_3631);
nand U3769 (N_3769,N_3695,N_3687);
nor U3770 (N_3770,N_3736,N_3667);
nor U3771 (N_3771,N_3733,N_3635);
nand U3772 (N_3772,N_3731,N_3668);
and U3773 (N_3773,N_3685,N_3641);
and U3774 (N_3774,N_3627,N_3656);
or U3775 (N_3775,N_3717,N_3640);
xor U3776 (N_3776,N_3740,N_3708);
xnor U3777 (N_3777,N_3657,N_3648);
nor U3778 (N_3778,N_3694,N_3703);
and U3779 (N_3779,N_3689,N_3725);
and U3780 (N_3780,N_3669,N_3650);
nand U3781 (N_3781,N_3721,N_3642);
xnor U3782 (N_3782,N_3699,N_3715);
nand U3783 (N_3783,N_3634,N_3693);
nand U3784 (N_3784,N_3730,N_3696);
and U3785 (N_3785,N_3691,N_3655);
and U3786 (N_3786,N_3719,N_3654);
or U3787 (N_3787,N_3646,N_3671);
nand U3788 (N_3788,N_3663,N_3724);
nor U3789 (N_3789,N_3726,N_3674);
or U3790 (N_3790,N_3625,N_3690);
and U3791 (N_3791,N_3701,N_3637);
xnor U3792 (N_3792,N_3749,N_3709);
and U3793 (N_3793,N_3633,N_3706);
xor U3794 (N_3794,N_3660,N_3697);
and U3795 (N_3795,N_3704,N_3683);
xor U3796 (N_3796,N_3739,N_3676);
xor U3797 (N_3797,N_3707,N_3662);
xnor U3798 (N_3798,N_3659,N_3653);
nor U3799 (N_3799,N_3713,N_3747);
nor U3800 (N_3800,N_3734,N_3738);
nor U3801 (N_3801,N_3629,N_3741);
or U3802 (N_3802,N_3727,N_3670);
xor U3803 (N_3803,N_3686,N_3743);
or U3804 (N_3804,N_3681,N_3666);
xor U3805 (N_3805,N_3698,N_3661);
xor U3806 (N_3806,N_3665,N_3744);
and U3807 (N_3807,N_3712,N_3684);
or U3808 (N_3808,N_3639,N_3711);
and U3809 (N_3809,N_3636,N_3714);
nor U3810 (N_3810,N_3728,N_3700);
or U3811 (N_3811,N_3737,N_3675);
nor U3812 (N_3812,N_3680,N_3638);
nor U3813 (N_3813,N_3733,N_3712);
and U3814 (N_3814,N_3705,N_3716);
nand U3815 (N_3815,N_3732,N_3745);
nand U3816 (N_3816,N_3747,N_3704);
and U3817 (N_3817,N_3724,N_3667);
and U3818 (N_3818,N_3658,N_3666);
xnor U3819 (N_3819,N_3726,N_3709);
nand U3820 (N_3820,N_3703,N_3708);
nor U3821 (N_3821,N_3724,N_3638);
nand U3822 (N_3822,N_3722,N_3693);
nor U3823 (N_3823,N_3746,N_3690);
xor U3824 (N_3824,N_3720,N_3666);
nand U3825 (N_3825,N_3739,N_3748);
nand U3826 (N_3826,N_3649,N_3712);
or U3827 (N_3827,N_3707,N_3719);
nor U3828 (N_3828,N_3635,N_3716);
or U3829 (N_3829,N_3721,N_3691);
nor U3830 (N_3830,N_3625,N_3639);
or U3831 (N_3831,N_3749,N_3635);
xnor U3832 (N_3832,N_3746,N_3724);
and U3833 (N_3833,N_3649,N_3708);
nand U3834 (N_3834,N_3736,N_3637);
nor U3835 (N_3835,N_3673,N_3748);
xnor U3836 (N_3836,N_3674,N_3634);
nand U3837 (N_3837,N_3705,N_3661);
xor U3838 (N_3838,N_3693,N_3745);
xnor U3839 (N_3839,N_3633,N_3692);
nor U3840 (N_3840,N_3667,N_3673);
nand U3841 (N_3841,N_3695,N_3699);
and U3842 (N_3842,N_3706,N_3656);
or U3843 (N_3843,N_3746,N_3657);
or U3844 (N_3844,N_3667,N_3735);
nand U3845 (N_3845,N_3630,N_3725);
nor U3846 (N_3846,N_3658,N_3730);
and U3847 (N_3847,N_3702,N_3725);
or U3848 (N_3848,N_3628,N_3635);
xor U3849 (N_3849,N_3632,N_3697);
nand U3850 (N_3850,N_3745,N_3701);
or U3851 (N_3851,N_3625,N_3640);
and U3852 (N_3852,N_3738,N_3675);
nor U3853 (N_3853,N_3725,N_3707);
and U3854 (N_3854,N_3749,N_3626);
nor U3855 (N_3855,N_3667,N_3630);
or U3856 (N_3856,N_3633,N_3652);
or U3857 (N_3857,N_3641,N_3658);
nor U3858 (N_3858,N_3660,N_3673);
or U3859 (N_3859,N_3668,N_3724);
nor U3860 (N_3860,N_3702,N_3718);
xnor U3861 (N_3861,N_3679,N_3747);
nor U3862 (N_3862,N_3721,N_3628);
or U3863 (N_3863,N_3696,N_3684);
nor U3864 (N_3864,N_3651,N_3744);
or U3865 (N_3865,N_3659,N_3727);
xnor U3866 (N_3866,N_3742,N_3650);
and U3867 (N_3867,N_3707,N_3657);
nand U3868 (N_3868,N_3734,N_3659);
xnor U3869 (N_3869,N_3685,N_3678);
xor U3870 (N_3870,N_3719,N_3743);
xor U3871 (N_3871,N_3626,N_3703);
xor U3872 (N_3872,N_3650,N_3625);
or U3873 (N_3873,N_3650,N_3677);
nor U3874 (N_3874,N_3682,N_3738);
xnor U3875 (N_3875,N_3772,N_3823);
xor U3876 (N_3876,N_3782,N_3786);
nand U3877 (N_3877,N_3790,N_3807);
nor U3878 (N_3878,N_3803,N_3766);
and U3879 (N_3879,N_3794,N_3835);
nand U3880 (N_3880,N_3762,N_3833);
nor U3881 (N_3881,N_3764,N_3850);
and U3882 (N_3882,N_3795,N_3813);
and U3883 (N_3883,N_3778,N_3815);
or U3884 (N_3884,N_3817,N_3758);
and U3885 (N_3885,N_3808,N_3780);
xnor U3886 (N_3886,N_3754,N_3822);
and U3887 (N_3887,N_3865,N_3828);
xnor U3888 (N_3888,N_3806,N_3771);
and U3889 (N_3889,N_3791,N_3799);
xor U3890 (N_3890,N_3751,N_3770);
nor U3891 (N_3891,N_3842,N_3852);
and U3892 (N_3892,N_3767,N_3805);
nand U3893 (N_3893,N_3841,N_3783);
nor U3894 (N_3894,N_3866,N_3812);
xor U3895 (N_3895,N_3818,N_3831);
or U3896 (N_3896,N_3847,N_3798);
xnor U3897 (N_3897,N_3752,N_3863);
nor U3898 (N_3898,N_3784,N_3868);
xor U3899 (N_3899,N_3819,N_3838);
nand U3900 (N_3900,N_3855,N_3853);
and U3901 (N_3901,N_3873,N_3800);
and U3902 (N_3902,N_3756,N_3824);
or U3903 (N_3903,N_3827,N_3834);
xor U3904 (N_3904,N_3769,N_3792);
nor U3905 (N_3905,N_3843,N_3781);
nand U3906 (N_3906,N_3848,N_3775);
xor U3907 (N_3907,N_3845,N_3862);
or U3908 (N_3908,N_3765,N_3832);
or U3909 (N_3909,N_3776,N_3854);
xor U3910 (N_3910,N_3797,N_3802);
and U3911 (N_3911,N_3851,N_3859);
and U3912 (N_3912,N_3788,N_3761);
or U3913 (N_3913,N_3759,N_3793);
nand U3914 (N_3914,N_3849,N_3816);
xnor U3915 (N_3915,N_3872,N_3753);
nor U3916 (N_3916,N_3857,N_3874);
nor U3917 (N_3917,N_3839,N_3763);
and U3918 (N_3918,N_3844,N_3864);
nor U3919 (N_3919,N_3773,N_3830);
nor U3920 (N_3920,N_3768,N_3809);
nand U3921 (N_3921,N_3760,N_3826);
nor U3922 (N_3922,N_3814,N_3810);
nand U3923 (N_3923,N_3846,N_3821);
nand U3924 (N_3924,N_3801,N_3840);
xor U3925 (N_3925,N_3858,N_3867);
and U3926 (N_3926,N_3804,N_3861);
or U3927 (N_3927,N_3871,N_3869);
and U3928 (N_3928,N_3789,N_3750);
and U3929 (N_3929,N_3856,N_3820);
xor U3930 (N_3930,N_3755,N_3829);
xnor U3931 (N_3931,N_3836,N_3796);
xor U3932 (N_3932,N_3774,N_3837);
nor U3933 (N_3933,N_3787,N_3785);
or U3934 (N_3934,N_3757,N_3779);
xnor U3935 (N_3935,N_3860,N_3777);
xor U3936 (N_3936,N_3825,N_3870);
or U3937 (N_3937,N_3811,N_3844);
nor U3938 (N_3938,N_3769,N_3763);
xor U3939 (N_3939,N_3763,N_3804);
and U3940 (N_3940,N_3840,N_3873);
or U3941 (N_3941,N_3833,N_3785);
xnor U3942 (N_3942,N_3859,N_3832);
and U3943 (N_3943,N_3824,N_3784);
nand U3944 (N_3944,N_3789,N_3862);
or U3945 (N_3945,N_3868,N_3833);
and U3946 (N_3946,N_3802,N_3841);
xor U3947 (N_3947,N_3870,N_3783);
nand U3948 (N_3948,N_3872,N_3783);
or U3949 (N_3949,N_3872,N_3805);
nor U3950 (N_3950,N_3752,N_3798);
or U3951 (N_3951,N_3780,N_3870);
and U3952 (N_3952,N_3783,N_3795);
nor U3953 (N_3953,N_3771,N_3809);
nor U3954 (N_3954,N_3864,N_3754);
nand U3955 (N_3955,N_3812,N_3843);
xor U3956 (N_3956,N_3769,N_3840);
or U3957 (N_3957,N_3831,N_3852);
or U3958 (N_3958,N_3820,N_3762);
xnor U3959 (N_3959,N_3856,N_3847);
nand U3960 (N_3960,N_3800,N_3844);
nor U3961 (N_3961,N_3829,N_3763);
and U3962 (N_3962,N_3847,N_3809);
nand U3963 (N_3963,N_3842,N_3869);
nand U3964 (N_3964,N_3859,N_3845);
xnor U3965 (N_3965,N_3790,N_3751);
nor U3966 (N_3966,N_3840,N_3863);
nor U3967 (N_3967,N_3815,N_3873);
nor U3968 (N_3968,N_3773,N_3823);
nand U3969 (N_3969,N_3814,N_3871);
nand U3970 (N_3970,N_3825,N_3759);
xnor U3971 (N_3971,N_3868,N_3768);
or U3972 (N_3972,N_3828,N_3840);
xor U3973 (N_3973,N_3821,N_3775);
or U3974 (N_3974,N_3812,N_3750);
nand U3975 (N_3975,N_3778,N_3840);
and U3976 (N_3976,N_3859,N_3771);
nor U3977 (N_3977,N_3754,N_3871);
and U3978 (N_3978,N_3811,N_3787);
or U3979 (N_3979,N_3761,N_3757);
nor U3980 (N_3980,N_3756,N_3780);
and U3981 (N_3981,N_3832,N_3789);
nor U3982 (N_3982,N_3837,N_3751);
nand U3983 (N_3983,N_3820,N_3778);
xnor U3984 (N_3984,N_3804,N_3873);
xor U3985 (N_3985,N_3763,N_3796);
and U3986 (N_3986,N_3777,N_3838);
and U3987 (N_3987,N_3791,N_3860);
xor U3988 (N_3988,N_3752,N_3848);
or U3989 (N_3989,N_3774,N_3796);
or U3990 (N_3990,N_3790,N_3840);
nand U3991 (N_3991,N_3826,N_3802);
nor U3992 (N_3992,N_3795,N_3771);
nand U3993 (N_3993,N_3813,N_3843);
or U3994 (N_3994,N_3791,N_3778);
and U3995 (N_3995,N_3821,N_3770);
nand U3996 (N_3996,N_3860,N_3826);
nor U3997 (N_3997,N_3809,N_3796);
xnor U3998 (N_3998,N_3775,N_3862);
xor U3999 (N_3999,N_3789,N_3852);
and U4000 (N_4000,N_3916,N_3957);
xnor U4001 (N_4001,N_3934,N_3925);
or U4002 (N_4002,N_3912,N_3914);
nand U4003 (N_4003,N_3913,N_3950);
and U4004 (N_4004,N_3878,N_3894);
nand U4005 (N_4005,N_3980,N_3963);
and U4006 (N_4006,N_3910,N_3884);
nor U4007 (N_4007,N_3926,N_3973);
nand U4008 (N_4008,N_3952,N_3997);
xor U4009 (N_4009,N_3995,N_3918);
xor U4010 (N_4010,N_3919,N_3983);
nor U4011 (N_4011,N_3906,N_3885);
and U4012 (N_4012,N_3887,N_3880);
and U4013 (N_4013,N_3961,N_3978);
and U4014 (N_4014,N_3943,N_3982);
and U4015 (N_4015,N_3991,N_3984);
and U4016 (N_4016,N_3897,N_3960);
nor U4017 (N_4017,N_3882,N_3956);
or U4018 (N_4018,N_3921,N_3881);
or U4019 (N_4019,N_3979,N_3972);
and U4020 (N_4020,N_3992,N_3904);
and U4021 (N_4021,N_3905,N_3927);
xor U4022 (N_4022,N_3876,N_3917);
nor U4023 (N_4023,N_3999,N_3923);
nand U4024 (N_4024,N_3964,N_3922);
xnor U4025 (N_4025,N_3928,N_3998);
and U4026 (N_4026,N_3948,N_3937);
xor U4027 (N_4027,N_3955,N_3965);
xor U4028 (N_4028,N_3933,N_3886);
and U4029 (N_4029,N_3875,N_3987);
nor U4030 (N_4030,N_3970,N_3889);
nand U4031 (N_4031,N_3936,N_3951);
nand U4032 (N_4032,N_3935,N_3968);
nor U4033 (N_4033,N_3931,N_3958);
and U4034 (N_4034,N_3888,N_3895);
xor U4035 (N_4035,N_3945,N_3915);
or U4036 (N_4036,N_3911,N_3908);
xor U4037 (N_4037,N_3975,N_3932);
and U4038 (N_4038,N_3907,N_3990);
nor U4039 (N_4039,N_3896,N_3971);
nand U4040 (N_4040,N_3976,N_3967);
or U4041 (N_4041,N_3946,N_3909);
and U4042 (N_4042,N_3901,N_3898);
xnor U4043 (N_4043,N_3944,N_3994);
or U4044 (N_4044,N_3890,N_3977);
nand U4045 (N_4045,N_3940,N_3949);
nor U4046 (N_4046,N_3899,N_3993);
nand U4047 (N_4047,N_3941,N_3877);
or U4048 (N_4048,N_3930,N_3953);
nor U4049 (N_4049,N_3893,N_3989);
xor U4050 (N_4050,N_3892,N_3900);
nand U4051 (N_4051,N_3938,N_3985);
and U4052 (N_4052,N_3986,N_3902);
or U4053 (N_4053,N_3939,N_3920);
xnor U4054 (N_4054,N_3959,N_3947);
nand U4055 (N_4055,N_3981,N_3891);
xnor U4056 (N_4056,N_3883,N_3974);
nor U4057 (N_4057,N_3942,N_3966);
and U4058 (N_4058,N_3988,N_3954);
xnor U4059 (N_4059,N_3924,N_3996);
and U4060 (N_4060,N_3962,N_3969);
xnor U4061 (N_4061,N_3903,N_3929);
nand U4062 (N_4062,N_3879,N_3967);
and U4063 (N_4063,N_3957,N_3946);
nand U4064 (N_4064,N_3993,N_3936);
xnor U4065 (N_4065,N_3899,N_3955);
nor U4066 (N_4066,N_3915,N_3927);
and U4067 (N_4067,N_3910,N_3958);
and U4068 (N_4068,N_3946,N_3908);
or U4069 (N_4069,N_3991,N_3897);
and U4070 (N_4070,N_3977,N_3887);
nor U4071 (N_4071,N_3944,N_3945);
xor U4072 (N_4072,N_3928,N_3959);
or U4073 (N_4073,N_3996,N_3985);
xnor U4074 (N_4074,N_3925,N_3969);
xnor U4075 (N_4075,N_3953,N_3997);
and U4076 (N_4076,N_3926,N_3949);
nor U4077 (N_4077,N_3889,N_3913);
nor U4078 (N_4078,N_3995,N_3898);
and U4079 (N_4079,N_3951,N_3935);
xor U4080 (N_4080,N_3949,N_3921);
xnor U4081 (N_4081,N_3981,N_3968);
nor U4082 (N_4082,N_3927,N_3876);
and U4083 (N_4083,N_3927,N_3932);
and U4084 (N_4084,N_3963,N_3961);
and U4085 (N_4085,N_3950,N_3988);
nor U4086 (N_4086,N_3944,N_3931);
xnor U4087 (N_4087,N_3912,N_3995);
and U4088 (N_4088,N_3962,N_3898);
and U4089 (N_4089,N_3908,N_3962);
xnor U4090 (N_4090,N_3889,N_3909);
and U4091 (N_4091,N_3976,N_3990);
nor U4092 (N_4092,N_3981,N_3907);
and U4093 (N_4093,N_3883,N_3929);
nand U4094 (N_4094,N_3894,N_3991);
or U4095 (N_4095,N_3943,N_3894);
or U4096 (N_4096,N_3913,N_3914);
and U4097 (N_4097,N_3936,N_3883);
nor U4098 (N_4098,N_3914,N_3976);
and U4099 (N_4099,N_3982,N_3985);
nand U4100 (N_4100,N_3935,N_3903);
xor U4101 (N_4101,N_3979,N_3907);
and U4102 (N_4102,N_3910,N_3875);
or U4103 (N_4103,N_3882,N_3889);
and U4104 (N_4104,N_3930,N_3983);
or U4105 (N_4105,N_3941,N_3988);
and U4106 (N_4106,N_3997,N_3876);
xnor U4107 (N_4107,N_3910,N_3931);
xor U4108 (N_4108,N_3880,N_3879);
nor U4109 (N_4109,N_3954,N_3961);
nor U4110 (N_4110,N_3971,N_3897);
or U4111 (N_4111,N_3959,N_3919);
and U4112 (N_4112,N_3934,N_3882);
nor U4113 (N_4113,N_3959,N_3878);
or U4114 (N_4114,N_3894,N_3950);
xnor U4115 (N_4115,N_3969,N_3900);
nor U4116 (N_4116,N_3907,N_3943);
nand U4117 (N_4117,N_3879,N_3878);
xnor U4118 (N_4118,N_3952,N_3950);
nor U4119 (N_4119,N_3921,N_3896);
xnor U4120 (N_4120,N_3933,N_3944);
or U4121 (N_4121,N_3889,N_3893);
nand U4122 (N_4122,N_3939,N_3972);
and U4123 (N_4123,N_3946,N_3944);
nor U4124 (N_4124,N_3915,N_3953);
xnor U4125 (N_4125,N_4070,N_4094);
nand U4126 (N_4126,N_4001,N_4048);
or U4127 (N_4127,N_4020,N_4009);
nor U4128 (N_4128,N_4111,N_4008);
xor U4129 (N_4129,N_4074,N_4011);
xor U4130 (N_4130,N_4116,N_4023);
nand U4131 (N_4131,N_4079,N_4067);
or U4132 (N_4132,N_4026,N_4017);
nor U4133 (N_4133,N_4100,N_4113);
nand U4134 (N_4134,N_4005,N_4080);
or U4135 (N_4135,N_4066,N_4027);
or U4136 (N_4136,N_4015,N_4082);
nor U4137 (N_4137,N_4053,N_4041);
nand U4138 (N_4138,N_4084,N_4090);
xor U4139 (N_4139,N_4002,N_4035);
xor U4140 (N_4140,N_4089,N_4103);
xnor U4141 (N_4141,N_4006,N_4092);
nor U4142 (N_4142,N_4122,N_4019);
and U4143 (N_4143,N_4059,N_4106);
nand U4144 (N_4144,N_4110,N_4016);
or U4145 (N_4145,N_4083,N_4121);
nand U4146 (N_4146,N_4037,N_4050);
and U4147 (N_4147,N_4112,N_4018);
nor U4148 (N_4148,N_4104,N_4031);
nor U4149 (N_4149,N_4007,N_4075);
nand U4150 (N_4150,N_4087,N_4021);
nand U4151 (N_4151,N_4049,N_4096);
and U4152 (N_4152,N_4065,N_4085);
or U4153 (N_4153,N_4118,N_4057);
and U4154 (N_4154,N_4119,N_4101);
nand U4155 (N_4155,N_4025,N_4120);
and U4156 (N_4156,N_4117,N_4062);
nor U4157 (N_4157,N_4044,N_4098);
xnor U4158 (N_4158,N_4069,N_4077);
xnor U4159 (N_4159,N_4014,N_4081);
or U4160 (N_4160,N_4004,N_4073);
xnor U4161 (N_4161,N_4013,N_4054);
xor U4162 (N_4162,N_4105,N_4097);
nor U4163 (N_4163,N_4043,N_4078);
or U4164 (N_4164,N_4072,N_4115);
or U4165 (N_4165,N_4028,N_4099);
or U4166 (N_4166,N_4109,N_4036);
and U4167 (N_4167,N_4114,N_4051);
or U4168 (N_4168,N_4039,N_4012);
nand U4169 (N_4169,N_4095,N_4055);
nand U4170 (N_4170,N_4088,N_4093);
nor U4171 (N_4171,N_4030,N_4124);
or U4172 (N_4172,N_4010,N_4024);
or U4173 (N_4173,N_4040,N_4064);
nand U4174 (N_4174,N_4032,N_4063);
or U4175 (N_4175,N_4034,N_4058);
nor U4176 (N_4176,N_4102,N_4033);
and U4177 (N_4177,N_4091,N_4029);
or U4178 (N_4178,N_4076,N_4045);
or U4179 (N_4179,N_4046,N_4038);
or U4180 (N_4180,N_4107,N_4022);
or U4181 (N_4181,N_4123,N_4068);
xnor U4182 (N_4182,N_4047,N_4061);
or U4183 (N_4183,N_4086,N_4060);
nand U4184 (N_4184,N_4056,N_4003);
nand U4185 (N_4185,N_4108,N_4042);
or U4186 (N_4186,N_4052,N_4071);
xor U4187 (N_4187,N_4000,N_4036);
xnor U4188 (N_4188,N_4069,N_4076);
and U4189 (N_4189,N_4034,N_4089);
xnor U4190 (N_4190,N_4070,N_4083);
nand U4191 (N_4191,N_4046,N_4015);
and U4192 (N_4192,N_4049,N_4120);
or U4193 (N_4193,N_4084,N_4068);
xnor U4194 (N_4194,N_4124,N_4004);
xnor U4195 (N_4195,N_4082,N_4039);
or U4196 (N_4196,N_4048,N_4070);
nor U4197 (N_4197,N_4085,N_4076);
xnor U4198 (N_4198,N_4018,N_4019);
nor U4199 (N_4199,N_4102,N_4003);
nand U4200 (N_4200,N_4019,N_4059);
nand U4201 (N_4201,N_4066,N_4032);
and U4202 (N_4202,N_4113,N_4029);
xor U4203 (N_4203,N_4024,N_4013);
xnor U4204 (N_4204,N_4059,N_4098);
nand U4205 (N_4205,N_4047,N_4064);
nor U4206 (N_4206,N_4124,N_4106);
xnor U4207 (N_4207,N_4024,N_4039);
and U4208 (N_4208,N_4031,N_4035);
or U4209 (N_4209,N_4039,N_4095);
nor U4210 (N_4210,N_4111,N_4115);
nor U4211 (N_4211,N_4021,N_4052);
and U4212 (N_4212,N_4030,N_4036);
and U4213 (N_4213,N_4100,N_4089);
nand U4214 (N_4214,N_4081,N_4030);
or U4215 (N_4215,N_4093,N_4001);
and U4216 (N_4216,N_4092,N_4097);
nor U4217 (N_4217,N_4048,N_4047);
nor U4218 (N_4218,N_4048,N_4068);
nor U4219 (N_4219,N_4063,N_4018);
nor U4220 (N_4220,N_4021,N_4064);
nand U4221 (N_4221,N_4029,N_4100);
nor U4222 (N_4222,N_4014,N_4121);
xnor U4223 (N_4223,N_4091,N_4046);
xnor U4224 (N_4224,N_4085,N_4009);
and U4225 (N_4225,N_4108,N_4004);
and U4226 (N_4226,N_4034,N_4110);
nor U4227 (N_4227,N_4069,N_4114);
nor U4228 (N_4228,N_4071,N_4042);
nand U4229 (N_4229,N_4099,N_4054);
and U4230 (N_4230,N_4089,N_4010);
xnor U4231 (N_4231,N_4084,N_4000);
or U4232 (N_4232,N_4006,N_4015);
nand U4233 (N_4233,N_4003,N_4075);
or U4234 (N_4234,N_4077,N_4073);
nor U4235 (N_4235,N_4011,N_4024);
or U4236 (N_4236,N_4071,N_4018);
and U4237 (N_4237,N_4103,N_4019);
and U4238 (N_4238,N_4087,N_4102);
nor U4239 (N_4239,N_4033,N_4098);
nor U4240 (N_4240,N_4096,N_4107);
xnor U4241 (N_4241,N_4076,N_4034);
and U4242 (N_4242,N_4008,N_4013);
nand U4243 (N_4243,N_4019,N_4110);
nor U4244 (N_4244,N_4022,N_4027);
or U4245 (N_4245,N_4022,N_4030);
or U4246 (N_4246,N_4071,N_4082);
nand U4247 (N_4247,N_4110,N_4077);
xnor U4248 (N_4248,N_4068,N_4049);
nand U4249 (N_4249,N_4047,N_4037);
nor U4250 (N_4250,N_4195,N_4207);
or U4251 (N_4251,N_4171,N_4185);
xnor U4252 (N_4252,N_4176,N_4153);
xnor U4253 (N_4253,N_4236,N_4149);
and U4254 (N_4254,N_4199,N_4213);
nor U4255 (N_4255,N_4206,N_4156);
and U4256 (N_4256,N_4175,N_4217);
or U4257 (N_4257,N_4205,N_4165);
xor U4258 (N_4258,N_4196,N_4132);
and U4259 (N_4259,N_4216,N_4241);
nor U4260 (N_4260,N_4233,N_4220);
nor U4261 (N_4261,N_4145,N_4188);
or U4262 (N_4262,N_4146,N_4133);
or U4263 (N_4263,N_4224,N_4139);
or U4264 (N_4264,N_4209,N_4142);
nor U4265 (N_4265,N_4163,N_4203);
or U4266 (N_4266,N_4226,N_4125);
and U4267 (N_4267,N_4210,N_4239);
and U4268 (N_4268,N_4235,N_4174);
nor U4269 (N_4269,N_4228,N_4137);
and U4270 (N_4270,N_4212,N_4246);
or U4271 (N_4271,N_4186,N_4223);
xnor U4272 (N_4272,N_4249,N_4243);
nor U4273 (N_4273,N_4225,N_4141);
nor U4274 (N_4274,N_4166,N_4184);
xnor U4275 (N_4275,N_4127,N_4214);
xor U4276 (N_4276,N_4178,N_4157);
or U4277 (N_4277,N_4218,N_4221);
xnor U4278 (N_4278,N_4169,N_4242);
or U4279 (N_4279,N_4179,N_4136);
nand U4280 (N_4280,N_4183,N_4192);
or U4281 (N_4281,N_4182,N_4234);
nor U4282 (N_4282,N_4131,N_4126);
nand U4283 (N_4283,N_4151,N_4211);
and U4284 (N_4284,N_4180,N_4201);
or U4285 (N_4285,N_4154,N_4130);
or U4286 (N_4286,N_4244,N_4194);
and U4287 (N_4287,N_4170,N_4162);
or U4288 (N_4288,N_4144,N_4152);
xnor U4289 (N_4289,N_4173,N_4231);
xnor U4290 (N_4290,N_4238,N_4219);
and U4291 (N_4291,N_4177,N_4167);
or U4292 (N_4292,N_4159,N_4197);
xor U4293 (N_4293,N_4143,N_4147);
or U4294 (N_4294,N_4248,N_4227);
nor U4295 (N_4295,N_4138,N_4155);
and U4296 (N_4296,N_4128,N_4187);
or U4297 (N_4297,N_4240,N_4204);
xnor U4298 (N_4298,N_4245,N_4208);
and U4299 (N_4299,N_4164,N_4172);
and U4300 (N_4300,N_4160,N_4148);
xor U4301 (N_4301,N_4190,N_4140);
xnor U4302 (N_4302,N_4198,N_4168);
xor U4303 (N_4303,N_4202,N_4230);
nor U4304 (N_4304,N_4129,N_4247);
and U4305 (N_4305,N_4158,N_4232);
xnor U4306 (N_4306,N_4200,N_4191);
and U4307 (N_4307,N_4229,N_4150);
nor U4308 (N_4308,N_4237,N_4161);
nand U4309 (N_4309,N_4193,N_4222);
nor U4310 (N_4310,N_4135,N_4189);
or U4311 (N_4311,N_4215,N_4181);
nor U4312 (N_4312,N_4134,N_4176);
nand U4313 (N_4313,N_4220,N_4234);
nor U4314 (N_4314,N_4131,N_4135);
or U4315 (N_4315,N_4204,N_4141);
xor U4316 (N_4316,N_4163,N_4204);
or U4317 (N_4317,N_4165,N_4228);
nor U4318 (N_4318,N_4198,N_4138);
nand U4319 (N_4319,N_4194,N_4211);
or U4320 (N_4320,N_4137,N_4161);
and U4321 (N_4321,N_4146,N_4215);
xnor U4322 (N_4322,N_4221,N_4162);
nand U4323 (N_4323,N_4148,N_4242);
or U4324 (N_4324,N_4237,N_4126);
xnor U4325 (N_4325,N_4191,N_4219);
nand U4326 (N_4326,N_4166,N_4199);
or U4327 (N_4327,N_4234,N_4140);
nor U4328 (N_4328,N_4241,N_4177);
or U4329 (N_4329,N_4233,N_4168);
xnor U4330 (N_4330,N_4150,N_4194);
and U4331 (N_4331,N_4199,N_4209);
or U4332 (N_4332,N_4201,N_4231);
or U4333 (N_4333,N_4209,N_4231);
nand U4334 (N_4334,N_4196,N_4168);
or U4335 (N_4335,N_4184,N_4169);
or U4336 (N_4336,N_4219,N_4144);
or U4337 (N_4337,N_4248,N_4190);
nand U4338 (N_4338,N_4202,N_4205);
and U4339 (N_4339,N_4136,N_4172);
or U4340 (N_4340,N_4173,N_4175);
nand U4341 (N_4341,N_4194,N_4151);
nand U4342 (N_4342,N_4233,N_4131);
and U4343 (N_4343,N_4211,N_4228);
xnor U4344 (N_4344,N_4130,N_4147);
xor U4345 (N_4345,N_4177,N_4208);
nor U4346 (N_4346,N_4188,N_4245);
nand U4347 (N_4347,N_4130,N_4193);
nand U4348 (N_4348,N_4225,N_4217);
and U4349 (N_4349,N_4164,N_4187);
and U4350 (N_4350,N_4215,N_4170);
nand U4351 (N_4351,N_4218,N_4219);
nand U4352 (N_4352,N_4238,N_4204);
nand U4353 (N_4353,N_4246,N_4151);
nor U4354 (N_4354,N_4217,N_4185);
nor U4355 (N_4355,N_4220,N_4158);
nor U4356 (N_4356,N_4192,N_4164);
nor U4357 (N_4357,N_4200,N_4236);
nor U4358 (N_4358,N_4228,N_4172);
xor U4359 (N_4359,N_4207,N_4231);
and U4360 (N_4360,N_4202,N_4195);
nand U4361 (N_4361,N_4128,N_4213);
or U4362 (N_4362,N_4204,N_4154);
nor U4363 (N_4363,N_4140,N_4145);
xnor U4364 (N_4364,N_4126,N_4193);
xnor U4365 (N_4365,N_4222,N_4192);
nor U4366 (N_4366,N_4184,N_4218);
or U4367 (N_4367,N_4172,N_4160);
nor U4368 (N_4368,N_4235,N_4128);
xnor U4369 (N_4369,N_4170,N_4235);
nand U4370 (N_4370,N_4198,N_4230);
or U4371 (N_4371,N_4249,N_4158);
nor U4372 (N_4372,N_4217,N_4241);
xnor U4373 (N_4373,N_4136,N_4241);
nor U4374 (N_4374,N_4233,N_4234);
nand U4375 (N_4375,N_4254,N_4315);
xor U4376 (N_4376,N_4357,N_4300);
xor U4377 (N_4377,N_4335,N_4253);
xnor U4378 (N_4378,N_4287,N_4266);
nor U4379 (N_4379,N_4255,N_4288);
and U4380 (N_4380,N_4317,N_4278);
and U4381 (N_4381,N_4274,N_4333);
and U4382 (N_4382,N_4330,N_4318);
or U4383 (N_4383,N_4269,N_4296);
or U4384 (N_4384,N_4314,N_4334);
nor U4385 (N_4385,N_4348,N_4354);
nand U4386 (N_4386,N_4309,N_4292);
and U4387 (N_4387,N_4262,N_4367);
xor U4388 (N_4388,N_4361,N_4359);
or U4389 (N_4389,N_4371,N_4310);
nor U4390 (N_4390,N_4299,N_4305);
nor U4391 (N_4391,N_4280,N_4328);
or U4392 (N_4392,N_4323,N_4308);
or U4393 (N_4393,N_4325,N_4268);
and U4394 (N_4394,N_4290,N_4322);
nand U4395 (N_4395,N_4257,N_4342);
and U4396 (N_4396,N_4295,N_4327);
xnor U4397 (N_4397,N_4250,N_4332);
and U4398 (N_4398,N_4284,N_4291);
xor U4399 (N_4399,N_4350,N_4276);
xnor U4400 (N_4400,N_4265,N_4336);
and U4401 (N_4401,N_4301,N_4352);
nor U4402 (N_4402,N_4273,N_4283);
or U4403 (N_4403,N_4364,N_4331);
nand U4404 (N_4404,N_4343,N_4261);
or U4405 (N_4405,N_4259,N_4281);
or U4406 (N_4406,N_4360,N_4271);
xnor U4407 (N_4407,N_4277,N_4286);
nor U4408 (N_4408,N_4298,N_4251);
xnor U4409 (N_4409,N_4306,N_4362);
and U4410 (N_4410,N_4329,N_4264);
and U4411 (N_4411,N_4289,N_4339);
nor U4412 (N_4412,N_4370,N_4372);
or U4413 (N_4413,N_4363,N_4349);
or U4414 (N_4414,N_4369,N_4356);
or U4415 (N_4415,N_4307,N_4252);
and U4416 (N_4416,N_4321,N_4319);
and U4417 (N_4417,N_4282,N_4355);
and U4418 (N_4418,N_4366,N_4345);
nand U4419 (N_4419,N_4358,N_4303);
nand U4420 (N_4420,N_4270,N_4341);
xnor U4421 (N_4421,N_4258,N_4316);
and U4422 (N_4422,N_4294,N_4340);
or U4423 (N_4423,N_4347,N_4346);
xnor U4424 (N_4424,N_4373,N_4353);
xor U4425 (N_4425,N_4326,N_4324);
or U4426 (N_4426,N_4293,N_4302);
and U4427 (N_4427,N_4285,N_4267);
nor U4428 (N_4428,N_4374,N_4337);
nand U4429 (N_4429,N_4279,N_4312);
nand U4430 (N_4430,N_4297,N_4344);
nor U4431 (N_4431,N_4275,N_4311);
nand U4432 (N_4432,N_4313,N_4338);
or U4433 (N_4433,N_4256,N_4263);
nand U4434 (N_4434,N_4351,N_4365);
xor U4435 (N_4435,N_4260,N_4272);
nor U4436 (N_4436,N_4304,N_4320);
xnor U4437 (N_4437,N_4368,N_4254);
or U4438 (N_4438,N_4286,N_4316);
nor U4439 (N_4439,N_4333,N_4325);
or U4440 (N_4440,N_4283,N_4353);
nand U4441 (N_4441,N_4259,N_4279);
nor U4442 (N_4442,N_4266,N_4315);
or U4443 (N_4443,N_4355,N_4258);
or U4444 (N_4444,N_4303,N_4315);
nand U4445 (N_4445,N_4326,N_4288);
and U4446 (N_4446,N_4286,N_4318);
nand U4447 (N_4447,N_4323,N_4351);
and U4448 (N_4448,N_4283,N_4358);
nand U4449 (N_4449,N_4257,N_4300);
nand U4450 (N_4450,N_4314,N_4338);
and U4451 (N_4451,N_4373,N_4257);
nor U4452 (N_4452,N_4283,N_4335);
xnor U4453 (N_4453,N_4277,N_4329);
or U4454 (N_4454,N_4353,N_4293);
nor U4455 (N_4455,N_4267,N_4339);
and U4456 (N_4456,N_4308,N_4325);
and U4457 (N_4457,N_4285,N_4286);
nor U4458 (N_4458,N_4346,N_4373);
and U4459 (N_4459,N_4340,N_4275);
and U4460 (N_4460,N_4287,N_4252);
and U4461 (N_4461,N_4355,N_4257);
nor U4462 (N_4462,N_4354,N_4251);
or U4463 (N_4463,N_4283,N_4339);
nor U4464 (N_4464,N_4311,N_4276);
nor U4465 (N_4465,N_4287,N_4316);
or U4466 (N_4466,N_4364,N_4324);
nand U4467 (N_4467,N_4273,N_4324);
nand U4468 (N_4468,N_4368,N_4317);
nor U4469 (N_4469,N_4276,N_4269);
or U4470 (N_4470,N_4327,N_4276);
nor U4471 (N_4471,N_4282,N_4285);
xor U4472 (N_4472,N_4281,N_4291);
or U4473 (N_4473,N_4347,N_4357);
xnor U4474 (N_4474,N_4271,N_4290);
and U4475 (N_4475,N_4285,N_4305);
nor U4476 (N_4476,N_4311,N_4329);
and U4477 (N_4477,N_4317,N_4346);
nand U4478 (N_4478,N_4356,N_4265);
nand U4479 (N_4479,N_4352,N_4364);
nand U4480 (N_4480,N_4278,N_4281);
and U4481 (N_4481,N_4312,N_4276);
or U4482 (N_4482,N_4340,N_4281);
nor U4483 (N_4483,N_4320,N_4314);
nor U4484 (N_4484,N_4358,N_4350);
nand U4485 (N_4485,N_4267,N_4336);
nor U4486 (N_4486,N_4307,N_4318);
nor U4487 (N_4487,N_4336,N_4295);
nand U4488 (N_4488,N_4253,N_4274);
nand U4489 (N_4489,N_4308,N_4283);
xnor U4490 (N_4490,N_4366,N_4288);
xnor U4491 (N_4491,N_4372,N_4362);
nand U4492 (N_4492,N_4253,N_4329);
xnor U4493 (N_4493,N_4270,N_4307);
xnor U4494 (N_4494,N_4351,N_4315);
xor U4495 (N_4495,N_4320,N_4324);
or U4496 (N_4496,N_4259,N_4289);
nor U4497 (N_4497,N_4324,N_4343);
xnor U4498 (N_4498,N_4313,N_4303);
xor U4499 (N_4499,N_4306,N_4276);
xnor U4500 (N_4500,N_4481,N_4435);
and U4501 (N_4501,N_4387,N_4498);
and U4502 (N_4502,N_4385,N_4479);
nand U4503 (N_4503,N_4375,N_4493);
xor U4504 (N_4504,N_4419,N_4461);
nor U4505 (N_4505,N_4394,N_4488);
or U4506 (N_4506,N_4464,N_4476);
or U4507 (N_4507,N_4441,N_4451);
xor U4508 (N_4508,N_4492,N_4449);
or U4509 (N_4509,N_4499,N_4421);
nand U4510 (N_4510,N_4485,N_4408);
nand U4511 (N_4511,N_4480,N_4411);
xnor U4512 (N_4512,N_4380,N_4457);
nand U4513 (N_4513,N_4425,N_4437);
and U4514 (N_4514,N_4433,N_4459);
and U4515 (N_4515,N_4398,N_4439);
nor U4516 (N_4516,N_4392,N_4454);
nand U4517 (N_4517,N_4400,N_4412);
nor U4518 (N_4518,N_4414,N_4404);
nor U4519 (N_4519,N_4410,N_4403);
xnor U4520 (N_4520,N_4395,N_4469);
nand U4521 (N_4521,N_4381,N_4473);
nand U4522 (N_4522,N_4489,N_4470);
nor U4523 (N_4523,N_4407,N_4379);
xor U4524 (N_4524,N_4429,N_4482);
nor U4525 (N_4525,N_4401,N_4452);
xnor U4526 (N_4526,N_4450,N_4495);
nand U4527 (N_4527,N_4426,N_4418);
or U4528 (N_4528,N_4382,N_4444);
nor U4529 (N_4529,N_4467,N_4468);
and U4530 (N_4530,N_4458,N_4428);
or U4531 (N_4531,N_4424,N_4465);
or U4532 (N_4532,N_4466,N_4446);
xor U4533 (N_4533,N_4384,N_4402);
and U4534 (N_4534,N_4383,N_4443);
or U4535 (N_4535,N_4472,N_4456);
nand U4536 (N_4536,N_4455,N_4486);
nand U4537 (N_4537,N_4494,N_4422);
xnor U4538 (N_4538,N_4420,N_4390);
nand U4539 (N_4539,N_4491,N_4445);
nand U4540 (N_4540,N_4490,N_4416);
nor U4541 (N_4541,N_4460,N_4487);
nand U4542 (N_4542,N_4447,N_4438);
nand U4543 (N_4543,N_4396,N_4409);
xnor U4544 (N_4544,N_4397,N_4497);
nor U4545 (N_4545,N_4415,N_4477);
or U4546 (N_4546,N_4484,N_4431);
nand U4547 (N_4547,N_4434,N_4378);
xor U4548 (N_4548,N_4388,N_4389);
nor U4549 (N_4549,N_4474,N_4436);
nand U4550 (N_4550,N_4442,N_4496);
xor U4551 (N_4551,N_4478,N_4417);
nor U4552 (N_4552,N_4448,N_4386);
nor U4553 (N_4553,N_4393,N_4376);
xor U4554 (N_4554,N_4399,N_4440);
and U4555 (N_4555,N_4377,N_4471);
and U4556 (N_4556,N_4423,N_4430);
or U4557 (N_4557,N_4453,N_4406);
nor U4558 (N_4558,N_4391,N_4483);
nor U4559 (N_4559,N_4463,N_4413);
and U4560 (N_4560,N_4427,N_4462);
and U4561 (N_4561,N_4432,N_4475);
nand U4562 (N_4562,N_4405,N_4377);
nor U4563 (N_4563,N_4464,N_4411);
xnor U4564 (N_4564,N_4466,N_4397);
and U4565 (N_4565,N_4392,N_4409);
nor U4566 (N_4566,N_4399,N_4497);
xor U4567 (N_4567,N_4483,N_4405);
nand U4568 (N_4568,N_4427,N_4485);
or U4569 (N_4569,N_4483,N_4401);
xnor U4570 (N_4570,N_4433,N_4423);
nand U4571 (N_4571,N_4392,N_4438);
nor U4572 (N_4572,N_4425,N_4467);
or U4573 (N_4573,N_4420,N_4378);
xnor U4574 (N_4574,N_4379,N_4405);
nor U4575 (N_4575,N_4465,N_4381);
nand U4576 (N_4576,N_4435,N_4411);
and U4577 (N_4577,N_4385,N_4391);
and U4578 (N_4578,N_4487,N_4480);
nand U4579 (N_4579,N_4383,N_4468);
xor U4580 (N_4580,N_4379,N_4450);
nor U4581 (N_4581,N_4406,N_4482);
nand U4582 (N_4582,N_4416,N_4482);
or U4583 (N_4583,N_4436,N_4415);
or U4584 (N_4584,N_4498,N_4453);
xnor U4585 (N_4585,N_4456,N_4388);
and U4586 (N_4586,N_4475,N_4461);
or U4587 (N_4587,N_4394,N_4442);
and U4588 (N_4588,N_4375,N_4453);
nor U4589 (N_4589,N_4486,N_4464);
nand U4590 (N_4590,N_4433,N_4387);
and U4591 (N_4591,N_4427,N_4395);
nor U4592 (N_4592,N_4403,N_4377);
nor U4593 (N_4593,N_4393,N_4437);
or U4594 (N_4594,N_4464,N_4406);
nor U4595 (N_4595,N_4476,N_4454);
or U4596 (N_4596,N_4430,N_4471);
or U4597 (N_4597,N_4453,N_4379);
xor U4598 (N_4598,N_4487,N_4404);
xnor U4599 (N_4599,N_4401,N_4455);
nand U4600 (N_4600,N_4454,N_4492);
xnor U4601 (N_4601,N_4423,N_4402);
and U4602 (N_4602,N_4456,N_4447);
and U4603 (N_4603,N_4471,N_4404);
or U4604 (N_4604,N_4449,N_4465);
nand U4605 (N_4605,N_4462,N_4431);
nor U4606 (N_4606,N_4462,N_4467);
xor U4607 (N_4607,N_4416,N_4498);
nor U4608 (N_4608,N_4465,N_4401);
nor U4609 (N_4609,N_4427,N_4428);
xnor U4610 (N_4610,N_4435,N_4472);
or U4611 (N_4611,N_4394,N_4425);
xor U4612 (N_4612,N_4497,N_4396);
and U4613 (N_4613,N_4447,N_4424);
and U4614 (N_4614,N_4447,N_4406);
nand U4615 (N_4615,N_4454,N_4439);
and U4616 (N_4616,N_4451,N_4448);
nor U4617 (N_4617,N_4444,N_4452);
nor U4618 (N_4618,N_4491,N_4412);
and U4619 (N_4619,N_4487,N_4398);
nand U4620 (N_4620,N_4498,N_4478);
nand U4621 (N_4621,N_4444,N_4446);
xnor U4622 (N_4622,N_4446,N_4469);
or U4623 (N_4623,N_4383,N_4397);
nand U4624 (N_4624,N_4495,N_4412);
and U4625 (N_4625,N_4537,N_4503);
or U4626 (N_4626,N_4608,N_4588);
xnor U4627 (N_4627,N_4547,N_4622);
and U4628 (N_4628,N_4513,N_4580);
and U4629 (N_4629,N_4614,N_4523);
and U4630 (N_4630,N_4516,N_4551);
xor U4631 (N_4631,N_4526,N_4619);
xor U4632 (N_4632,N_4609,N_4500);
xor U4633 (N_4633,N_4606,N_4535);
nor U4634 (N_4634,N_4557,N_4563);
nand U4635 (N_4635,N_4529,N_4542);
or U4636 (N_4636,N_4617,N_4599);
xor U4637 (N_4637,N_4543,N_4561);
nand U4638 (N_4638,N_4607,N_4618);
and U4639 (N_4639,N_4527,N_4518);
nor U4640 (N_4640,N_4530,N_4534);
xor U4641 (N_4641,N_4584,N_4512);
nand U4642 (N_4642,N_4568,N_4601);
or U4643 (N_4643,N_4511,N_4560);
xor U4644 (N_4644,N_4579,N_4524);
nand U4645 (N_4645,N_4623,N_4552);
nor U4646 (N_4646,N_4578,N_4509);
xnor U4647 (N_4647,N_4525,N_4536);
xor U4648 (N_4648,N_4541,N_4502);
nor U4649 (N_4649,N_4507,N_4575);
xor U4650 (N_4650,N_4531,N_4573);
or U4651 (N_4651,N_4559,N_4596);
nor U4652 (N_4652,N_4532,N_4592);
xnor U4653 (N_4653,N_4571,N_4594);
xor U4654 (N_4654,N_4554,N_4510);
nand U4655 (N_4655,N_4528,N_4585);
and U4656 (N_4656,N_4612,N_4611);
nor U4657 (N_4657,N_4549,N_4598);
or U4658 (N_4658,N_4519,N_4548);
xor U4659 (N_4659,N_4506,N_4514);
xnor U4660 (N_4660,N_4550,N_4610);
or U4661 (N_4661,N_4553,N_4583);
xor U4662 (N_4662,N_4522,N_4605);
nor U4663 (N_4663,N_4546,N_4538);
nor U4664 (N_4664,N_4615,N_4517);
or U4665 (N_4665,N_4555,N_4570);
nand U4666 (N_4666,N_4545,N_4582);
nand U4667 (N_4667,N_4591,N_4587);
xnor U4668 (N_4668,N_4616,N_4564);
or U4669 (N_4669,N_4613,N_4581);
and U4670 (N_4670,N_4597,N_4566);
nand U4671 (N_4671,N_4586,N_4589);
xor U4672 (N_4672,N_4602,N_4501);
nor U4673 (N_4673,N_4590,N_4558);
nand U4674 (N_4674,N_4562,N_4593);
and U4675 (N_4675,N_4621,N_4520);
nor U4676 (N_4676,N_4556,N_4595);
or U4677 (N_4677,N_4540,N_4504);
or U4678 (N_4678,N_4544,N_4567);
or U4679 (N_4679,N_4620,N_4565);
nor U4680 (N_4680,N_4515,N_4624);
nand U4681 (N_4681,N_4600,N_4508);
or U4682 (N_4682,N_4577,N_4574);
and U4683 (N_4683,N_4604,N_4521);
nand U4684 (N_4684,N_4572,N_4533);
or U4685 (N_4685,N_4576,N_4603);
or U4686 (N_4686,N_4539,N_4505);
xor U4687 (N_4687,N_4569,N_4606);
nand U4688 (N_4688,N_4621,N_4548);
and U4689 (N_4689,N_4510,N_4525);
or U4690 (N_4690,N_4554,N_4574);
xnor U4691 (N_4691,N_4607,N_4566);
nand U4692 (N_4692,N_4533,N_4510);
xor U4693 (N_4693,N_4561,N_4530);
nand U4694 (N_4694,N_4537,N_4540);
and U4695 (N_4695,N_4603,N_4617);
nand U4696 (N_4696,N_4549,N_4548);
nor U4697 (N_4697,N_4562,N_4511);
and U4698 (N_4698,N_4616,N_4596);
or U4699 (N_4699,N_4553,N_4621);
nor U4700 (N_4700,N_4548,N_4606);
xor U4701 (N_4701,N_4602,N_4591);
nor U4702 (N_4702,N_4545,N_4604);
nand U4703 (N_4703,N_4545,N_4500);
nand U4704 (N_4704,N_4559,N_4552);
nand U4705 (N_4705,N_4565,N_4530);
nand U4706 (N_4706,N_4605,N_4543);
nand U4707 (N_4707,N_4589,N_4516);
and U4708 (N_4708,N_4518,N_4548);
or U4709 (N_4709,N_4573,N_4533);
nand U4710 (N_4710,N_4614,N_4584);
or U4711 (N_4711,N_4547,N_4519);
nand U4712 (N_4712,N_4590,N_4556);
and U4713 (N_4713,N_4568,N_4504);
nand U4714 (N_4714,N_4600,N_4547);
nand U4715 (N_4715,N_4574,N_4558);
and U4716 (N_4716,N_4599,N_4551);
nor U4717 (N_4717,N_4545,N_4588);
or U4718 (N_4718,N_4602,N_4624);
nand U4719 (N_4719,N_4588,N_4556);
nand U4720 (N_4720,N_4530,N_4501);
or U4721 (N_4721,N_4526,N_4544);
or U4722 (N_4722,N_4531,N_4552);
or U4723 (N_4723,N_4585,N_4600);
nor U4724 (N_4724,N_4613,N_4520);
nand U4725 (N_4725,N_4554,N_4585);
nand U4726 (N_4726,N_4591,N_4517);
and U4727 (N_4727,N_4610,N_4549);
nor U4728 (N_4728,N_4602,N_4577);
and U4729 (N_4729,N_4518,N_4530);
nor U4730 (N_4730,N_4551,N_4545);
nor U4731 (N_4731,N_4586,N_4517);
nor U4732 (N_4732,N_4562,N_4573);
nor U4733 (N_4733,N_4615,N_4584);
nor U4734 (N_4734,N_4544,N_4530);
xor U4735 (N_4735,N_4514,N_4608);
or U4736 (N_4736,N_4524,N_4506);
or U4737 (N_4737,N_4553,N_4578);
or U4738 (N_4738,N_4528,N_4601);
nor U4739 (N_4739,N_4550,N_4526);
nand U4740 (N_4740,N_4534,N_4620);
and U4741 (N_4741,N_4534,N_4566);
xor U4742 (N_4742,N_4503,N_4578);
xnor U4743 (N_4743,N_4515,N_4551);
or U4744 (N_4744,N_4592,N_4549);
or U4745 (N_4745,N_4515,N_4531);
or U4746 (N_4746,N_4534,N_4554);
nand U4747 (N_4747,N_4557,N_4621);
xor U4748 (N_4748,N_4521,N_4583);
xor U4749 (N_4749,N_4517,N_4609);
and U4750 (N_4750,N_4665,N_4690);
nor U4751 (N_4751,N_4710,N_4731);
nor U4752 (N_4752,N_4711,N_4681);
nand U4753 (N_4753,N_4655,N_4680);
xor U4754 (N_4754,N_4704,N_4669);
xor U4755 (N_4755,N_4633,N_4627);
or U4756 (N_4756,N_4642,N_4726);
xnor U4757 (N_4757,N_4639,N_4738);
xor U4758 (N_4758,N_4654,N_4729);
and U4759 (N_4759,N_4641,N_4716);
nand U4760 (N_4760,N_4628,N_4705);
xnor U4761 (N_4761,N_4743,N_4713);
nand U4762 (N_4762,N_4663,N_4652);
nand U4763 (N_4763,N_4649,N_4679);
and U4764 (N_4764,N_4703,N_4643);
and U4765 (N_4765,N_4675,N_4694);
nand U4766 (N_4766,N_4749,N_4644);
and U4767 (N_4767,N_4676,N_4709);
or U4768 (N_4768,N_4725,N_4719);
xnor U4769 (N_4769,N_4683,N_4692);
xor U4770 (N_4770,N_4689,N_4706);
nand U4771 (N_4771,N_4741,N_4670);
xnor U4772 (N_4772,N_4691,N_4634);
and U4773 (N_4773,N_4727,N_4721);
and U4774 (N_4774,N_4688,N_4724);
and U4775 (N_4775,N_4648,N_4678);
xnor U4776 (N_4776,N_4632,N_4728);
and U4777 (N_4777,N_4640,N_4699);
or U4778 (N_4778,N_4739,N_4717);
xor U4779 (N_4779,N_4636,N_4733);
nor U4780 (N_4780,N_4684,N_4714);
and U4781 (N_4781,N_4745,N_4646);
or U4782 (N_4782,N_4748,N_4723);
or U4783 (N_4783,N_4664,N_4650);
or U4784 (N_4784,N_4737,N_4707);
and U4785 (N_4785,N_4645,N_4647);
xor U4786 (N_4786,N_4682,N_4629);
nor U4787 (N_4787,N_4700,N_4658);
nor U4788 (N_4788,N_4674,N_4697);
and U4789 (N_4789,N_4740,N_4630);
and U4790 (N_4790,N_4672,N_4736);
or U4791 (N_4791,N_4747,N_4659);
nor U4792 (N_4792,N_4730,N_4671);
or U4793 (N_4793,N_4720,N_4744);
and U4794 (N_4794,N_4746,N_4661);
xnor U4795 (N_4795,N_4626,N_4637);
nand U4796 (N_4796,N_4677,N_4734);
nor U4797 (N_4797,N_4651,N_4668);
xnor U4798 (N_4798,N_4708,N_4722);
xor U4799 (N_4799,N_4735,N_4718);
xor U4800 (N_4800,N_4660,N_4635);
nor U4801 (N_4801,N_4696,N_4687);
nor U4802 (N_4802,N_4732,N_4653);
or U4803 (N_4803,N_4673,N_4656);
nand U4804 (N_4804,N_4715,N_4695);
nor U4805 (N_4805,N_4693,N_4686);
or U4806 (N_4806,N_4702,N_4657);
nor U4807 (N_4807,N_4712,N_4685);
or U4808 (N_4808,N_4625,N_4742);
nor U4809 (N_4809,N_4638,N_4662);
and U4810 (N_4810,N_4701,N_4631);
or U4811 (N_4811,N_4666,N_4667);
nor U4812 (N_4812,N_4698,N_4681);
or U4813 (N_4813,N_4636,N_4748);
and U4814 (N_4814,N_4705,N_4731);
xnor U4815 (N_4815,N_4666,N_4626);
and U4816 (N_4816,N_4641,N_4726);
xnor U4817 (N_4817,N_4697,N_4734);
or U4818 (N_4818,N_4660,N_4646);
or U4819 (N_4819,N_4699,N_4673);
nand U4820 (N_4820,N_4706,N_4694);
nand U4821 (N_4821,N_4672,N_4701);
nor U4822 (N_4822,N_4678,N_4685);
nand U4823 (N_4823,N_4711,N_4727);
xor U4824 (N_4824,N_4697,N_4741);
and U4825 (N_4825,N_4651,N_4730);
or U4826 (N_4826,N_4649,N_4737);
xor U4827 (N_4827,N_4709,N_4705);
nand U4828 (N_4828,N_4682,N_4677);
and U4829 (N_4829,N_4626,N_4628);
or U4830 (N_4830,N_4664,N_4660);
nor U4831 (N_4831,N_4656,N_4683);
or U4832 (N_4832,N_4748,N_4635);
nor U4833 (N_4833,N_4653,N_4661);
and U4834 (N_4834,N_4715,N_4687);
xnor U4835 (N_4835,N_4733,N_4630);
or U4836 (N_4836,N_4739,N_4746);
nand U4837 (N_4837,N_4698,N_4649);
nand U4838 (N_4838,N_4654,N_4738);
xor U4839 (N_4839,N_4660,N_4713);
nor U4840 (N_4840,N_4689,N_4742);
nor U4841 (N_4841,N_4627,N_4674);
or U4842 (N_4842,N_4625,N_4666);
xor U4843 (N_4843,N_4700,N_4652);
or U4844 (N_4844,N_4749,N_4680);
nand U4845 (N_4845,N_4703,N_4744);
and U4846 (N_4846,N_4673,N_4667);
nor U4847 (N_4847,N_4724,N_4685);
nand U4848 (N_4848,N_4684,N_4660);
or U4849 (N_4849,N_4728,N_4670);
nand U4850 (N_4850,N_4691,N_4747);
and U4851 (N_4851,N_4733,N_4704);
or U4852 (N_4852,N_4699,N_4718);
and U4853 (N_4853,N_4690,N_4719);
and U4854 (N_4854,N_4647,N_4693);
nand U4855 (N_4855,N_4673,N_4657);
or U4856 (N_4856,N_4661,N_4628);
and U4857 (N_4857,N_4628,N_4715);
nand U4858 (N_4858,N_4692,N_4713);
nor U4859 (N_4859,N_4721,N_4677);
nand U4860 (N_4860,N_4708,N_4723);
or U4861 (N_4861,N_4687,N_4718);
or U4862 (N_4862,N_4671,N_4659);
and U4863 (N_4863,N_4700,N_4644);
or U4864 (N_4864,N_4693,N_4710);
xnor U4865 (N_4865,N_4714,N_4708);
and U4866 (N_4866,N_4727,N_4733);
nand U4867 (N_4867,N_4749,N_4653);
nand U4868 (N_4868,N_4694,N_4698);
nand U4869 (N_4869,N_4688,N_4749);
and U4870 (N_4870,N_4686,N_4656);
and U4871 (N_4871,N_4650,N_4677);
nor U4872 (N_4872,N_4715,N_4733);
xnor U4873 (N_4873,N_4654,N_4741);
and U4874 (N_4874,N_4638,N_4708);
nor U4875 (N_4875,N_4834,N_4755);
nand U4876 (N_4876,N_4832,N_4859);
xnor U4877 (N_4877,N_4781,N_4823);
nand U4878 (N_4878,N_4821,N_4815);
nor U4879 (N_4879,N_4836,N_4854);
xor U4880 (N_4880,N_4845,N_4774);
or U4881 (N_4881,N_4853,N_4765);
nor U4882 (N_4882,N_4791,N_4752);
nor U4883 (N_4883,N_4828,N_4852);
xnor U4884 (N_4884,N_4761,N_4770);
xnor U4885 (N_4885,N_4767,N_4809);
or U4886 (N_4886,N_4757,N_4870);
and U4887 (N_4887,N_4831,N_4863);
and U4888 (N_4888,N_4826,N_4797);
and U4889 (N_4889,N_4819,N_4833);
and U4890 (N_4890,N_4799,N_4754);
nand U4891 (N_4891,N_4825,N_4776);
nor U4892 (N_4892,N_4849,N_4868);
nand U4893 (N_4893,N_4778,N_4785);
or U4894 (N_4894,N_4793,N_4783);
or U4895 (N_4895,N_4795,N_4871);
nand U4896 (N_4896,N_4794,N_4822);
nand U4897 (N_4897,N_4788,N_4777);
or U4898 (N_4898,N_4803,N_4843);
nor U4899 (N_4899,N_4760,N_4846);
nor U4900 (N_4900,N_4782,N_4808);
and U4901 (N_4901,N_4844,N_4762);
and U4902 (N_4902,N_4772,N_4806);
nand U4903 (N_4903,N_4759,N_4848);
or U4904 (N_4904,N_4779,N_4872);
nand U4905 (N_4905,N_4802,N_4796);
and U4906 (N_4906,N_4768,N_4764);
and U4907 (N_4907,N_4824,N_4798);
nand U4908 (N_4908,N_4784,N_4839);
and U4909 (N_4909,N_4751,N_4813);
nand U4910 (N_4910,N_4753,N_4850);
and U4911 (N_4911,N_4769,N_4865);
nand U4912 (N_4912,N_4812,N_4835);
xnor U4913 (N_4913,N_4756,N_4867);
or U4914 (N_4914,N_4862,N_4866);
nor U4915 (N_4915,N_4807,N_4847);
nor U4916 (N_4916,N_4804,N_4855);
and U4917 (N_4917,N_4869,N_4800);
nor U4918 (N_4918,N_4874,N_4829);
and U4919 (N_4919,N_4780,N_4873);
and U4920 (N_4920,N_4750,N_4858);
xnor U4921 (N_4921,N_4786,N_4860);
nor U4922 (N_4922,N_4842,N_4830);
xnor U4923 (N_4923,N_4851,N_4790);
and U4924 (N_4924,N_4775,N_4810);
nor U4925 (N_4925,N_4837,N_4827);
or U4926 (N_4926,N_4787,N_4841);
nor U4927 (N_4927,N_4818,N_4771);
nor U4928 (N_4928,N_4805,N_4817);
or U4929 (N_4929,N_4864,N_4816);
or U4930 (N_4930,N_4856,N_4792);
or U4931 (N_4931,N_4857,N_4801);
nor U4932 (N_4932,N_4773,N_4811);
and U4933 (N_4933,N_4838,N_4861);
nand U4934 (N_4934,N_4758,N_4766);
or U4935 (N_4935,N_4789,N_4820);
or U4936 (N_4936,N_4840,N_4814);
and U4937 (N_4937,N_4763,N_4829);
and U4938 (N_4938,N_4770,N_4823);
xnor U4939 (N_4939,N_4832,N_4760);
nor U4940 (N_4940,N_4796,N_4779);
nand U4941 (N_4941,N_4832,N_4873);
nand U4942 (N_4942,N_4767,N_4849);
nand U4943 (N_4943,N_4816,N_4752);
xor U4944 (N_4944,N_4814,N_4772);
nor U4945 (N_4945,N_4836,N_4825);
and U4946 (N_4946,N_4830,N_4859);
nand U4947 (N_4947,N_4751,N_4856);
xor U4948 (N_4948,N_4848,N_4802);
nor U4949 (N_4949,N_4759,N_4835);
nand U4950 (N_4950,N_4806,N_4770);
xnor U4951 (N_4951,N_4854,N_4781);
or U4952 (N_4952,N_4805,N_4789);
and U4953 (N_4953,N_4840,N_4804);
nor U4954 (N_4954,N_4792,N_4805);
or U4955 (N_4955,N_4865,N_4815);
or U4956 (N_4956,N_4831,N_4854);
xor U4957 (N_4957,N_4825,N_4868);
or U4958 (N_4958,N_4778,N_4821);
or U4959 (N_4959,N_4789,N_4845);
or U4960 (N_4960,N_4765,N_4857);
nor U4961 (N_4961,N_4769,N_4801);
or U4962 (N_4962,N_4808,N_4760);
and U4963 (N_4963,N_4820,N_4769);
and U4964 (N_4964,N_4792,N_4844);
or U4965 (N_4965,N_4756,N_4821);
nand U4966 (N_4966,N_4827,N_4847);
xor U4967 (N_4967,N_4837,N_4771);
xor U4968 (N_4968,N_4859,N_4854);
nand U4969 (N_4969,N_4858,N_4792);
xnor U4970 (N_4970,N_4802,N_4821);
nand U4971 (N_4971,N_4762,N_4829);
xnor U4972 (N_4972,N_4811,N_4872);
or U4973 (N_4973,N_4817,N_4832);
nor U4974 (N_4974,N_4794,N_4865);
nand U4975 (N_4975,N_4773,N_4761);
nand U4976 (N_4976,N_4766,N_4873);
and U4977 (N_4977,N_4839,N_4855);
or U4978 (N_4978,N_4811,N_4843);
nand U4979 (N_4979,N_4791,N_4869);
and U4980 (N_4980,N_4828,N_4815);
and U4981 (N_4981,N_4825,N_4786);
nor U4982 (N_4982,N_4873,N_4803);
or U4983 (N_4983,N_4797,N_4812);
or U4984 (N_4984,N_4756,N_4751);
nor U4985 (N_4985,N_4815,N_4764);
xor U4986 (N_4986,N_4844,N_4786);
and U4987 (N_4987,N_4765,N_4872);
xnor U4988 (N_4988,N_4816,N_4870);
or U4989 (N_4989,N_4751,N_4770);
xor U4990 (N_4990,N_4822,N_4764);
or U4991 (N_4991,N_4829,N_4821);
and U4992 (N_4992,N_4816,N_4823);
nand U4993 (N_4993,N_4763,N_4845);
xor U4994 (N_4994,N_4826,N_4789);
nor U4995 (N_4995,N_4757,N_4838);
nand U4996 (N_4996,N_4841,N_4799);
and U4997 (N_4997,N_4865,N_4751);
xnor U4998 (N_4998,N_4815,N_4830);
nand U4999 (N_4999,N_4827,N_4815);
nor U5000 (N_5000,N_4999,N_4876);
and U5001 (N_5001,N_4901,N_4981);
nor U5002 (N_5002,N_4878,N_4911);
nand U5003 (N_5003,N_4883,N_4924);
and U5004 (N_5004,N_4907,N_4952);
xnor U5005 (N_5005,N_4906,N_4925);
and U5006 (N_5006,N_4880,N_4899);
nor U5007 (N_5007,N_4900,N_4948);
nor U5008 (N_5008,N_4969,N_4976);
xnor U5009 (N_5009,N_4955,N_4930);
nor U5010 (N_5010,N_4931,N_4973);
nor U5011 (N_5011,N_4892,N_4914);
xnor U5012 (N_5012,N_4893,N_4912);
nor U5013 (N_5013,N_4963,N_4934);
and U5014 (N_5014,N_4958,N_4923);
xor U5015 (N_5015,N_4921,N_4903);
xnor U5016 (N_5016,N_4884,N_4894);
and U5017 (N_5017,N_4954,N_4940);
or U5018 (N_5018,N_4928,N_4950);
nand U5019 (N_5019,N_4896,N_4909);
nand U5020 (N_5020,N_4971,N_4974);
nand U5021 (N_5021,N_4986,N_4965);
and U5022 (N_5022,N_4951,N_4937);
nand U5023 (N_5023,N_4939,N_4943);
or U5024 (N_5024,N_4945,N_4875);
or U5025 (N_5025,N_4961,N_4984);
or U5026 (N_5026,N_4978,N_4929);
nand U5027 (N_5027,N_4985,N_4990);
nor U5028 (N_5028,N_4881,N_4895);
or U5029 (N_5029,N_4993,N_4916);
and U5030 (N_5030,N_4982,N_4942);
nand U5031 (N_5031,N_4913,N_4977);
and U5032 (N_5032,N_4962,N_4975);
nor U5033 (N_5033,N_4988,N_4917);
nor U5034 (N_5034,N_4989,N_4996);
nor U5035 (N_5035,N_4890,N_4898);
or U5036 (N_5036,N_4936,N_4991);
nor U5037 (N_5037,N_4922,N_4918);
and U5038 (N_5038,N_4979,N_4947);
nand U5039 (N_5039,N_4926,N_4987);
xnor U5040 (N_5040,N_4966,N_4964);
and U5041 (N_5041,N_4944,N_4932);
or U5042 (N_5042,N_4953,N_4967);
nor U5043 (N_5043,N_4920,N_4905);
or U5044 (N_5044,N_4902,N_4915);
xnor U5045 (N_5045,N_4910,N_4949);
and U5046 (N_5046,N_4970,N_4957);
nand U5047 (N_5047,N_4887,N_4941);
or U5048 (N_5048,N_4919,N_4946);
or U5049 (N_5049,N_4968,N_4956);
and U5050 (N_5050,N_4904,N_4897);
and U5051 (N_5051,N_4935,N_4972);
xnor U5052 (N_5052,N_4885,N_4927);
nand U5053 (N_5053,N_4960,N_4980);
or U5054 (N_5054,N_4889,N_4891);
nand U5055 (N_5055,N_4877,N_4959);
nor U5056 (N_5056,N_4882,N_4879);
xor U5057 (N_5057,N_4886,N_4998);
nor U5058 (N_5058,N_4938,N_4992);
xor U5059 (N_5059,N_4994,N_4995);
nor U5060 (N_5060,N_4908,N_4888);
nor U5061 (N_5061,N_4997,N_4933);
and U5062 (N_5062,N_4983,N_4937);
nand U5063 (N_5063,N_4907,N_4956);
or U5064 (N_5064,N_4989,N_4920);
xor U5065 (N_5065,N_4904,N_4990);
nand U5066 (N_5066,N_4987,N_4948);
nand U5067 (N_5067,N_4922,N_4924);
and U5068 (N_5068,N_4930,N_4899);
xnor U5069 (N_5069,N_4896,N_4990);
nor U5070 (N_5070,N_4969,N_4881);
nor U5071 (N_5071,N_4938,N_4908);
nor U5072 (N_5072,N_4894,N_4901);
nand U5073 (N_5073,N_4878,N_4945);
nor U5074 (N_5074,N_4906,N_4930);
or U5075 (N_5075,N_4994,N_4914);
nor U5076 (N_5076,N_4945,N_4967);
or U5077 (N_5077,N_4983,N_4945);
and U5078 (N_5078,N_4924,N_4963);
nor U5079 (N_5079,N_4904,N_4934);
and U5080 (N_5080,N_4922,N_4956);
or U5081 (N_5081,N_4977,N_4936);
or U5082 (N_5082,N_4903,N_4973);
or U5083 (N_5083,N_4876,N_4996);
nand U5084 (N_5084,N_4884,N_4989);
nand U5085 (N_5085,N_4955,N_4912);
and U5086 (N_5086,N_4985,N_4964);
and U5087 (N_5087,N_4892,N_4915);
or U5088 (N_5088,N_4889,N_4965);
nand U5089 (N_5089,N_4906,N_4945);
and U5090 (N_5090,N_4902,N_4973);
or U5091 (N_5091,N_4972,N_4967);
and U5092 (N_5092,N_4960,N_4940);
xor U5093 (N_5093,N_4986,N_4994);
xor U5094 (N_5094,N_4984,N_4972);
xor U5095 (N_5095,N_4906,N_4948);
xor U5096 (N_5096,N_4969,N_4944);
or U5097 (N_5097,N_4906,N_4972);
nor U5098 (N_5098,N_4949,N_4897);
and U5099 (N_5099,N_4899,N_4949);
or U5100 (N_5100,N_4971,N_4924);
nor U5101 (N_5101,N_4943,N_4896);
nand U5102 (N_5102,N_4904,N_4937);
or U5103 (N_5103,N_4882,N_4938);
or U5104 (N_5104,N_4968,N_4946);
nand U5105 (N_5105,N_4934,N_4984);
or U5106 (N_5106,N_4965,N_4899);
nand U5107 (N_5107,N_4930,N_4968);
xnor U5108 (N_5108,N_4900,N_4895);
nand U5109 (N_5109,N_4892,N_4972);
nand U5110 (N_5110,N_4900,N_4886);
nor U5111 (N_5111,N_4897,N_4890);
nand U5112 (N_5112,N_4925,N_4966);
xor U5113 (N_5113,N_4920,N_4928);
nor U5114 (N_5114,N_4980,N_4982);
nor U5115 (N_5115,N_4946,N_4983);
nand U5116 (N_5116,N_4886,N_4921);
xnor U5117 (N_5117,N_4979,N_4963);
and U5118 (N_5118,N_4904,N_4885);
nand U5119 (N_5119,N_4984,N_4936);
or U5120 (N_5120,N_4964,N_4916);
nor U5121 (N_5121,N_4975,N_4891);
or U5122 (N_5122,N_4944,N_4965);
xnor U5123 (N_5123,N_4904,N_4973);
xor U5124 (N_5124,N_4947,N_4935);
nor U5125 (N_5125,N_5093,N_5108);
or U5126 (N_5126,N_5115,N_5096);
nor U5127 (N_5127,N_5111,N_5122);
and U5128 (N_5128,N_5101,N_5049);
xor U5129 (N_5129,N_5120,N_5019);
or U5130 (N_5130,N_5103,N_5034);
nand U5131 (N_5131,N_5086,N_5112);
xor U5132 (N_5132,N_5063,N_5087);
or U5133 (N_5133,N_5100,N_5121);
nor U5134 (N_5134,N_5033,N_5051);
xor U5135 (N_5135,N_5014,N_5055);
and U5136 (N_5136,N_5045,N_5094);
or U5137 (N_5137,N_5095,N_5009);
nor U5138 (N_5138,N_5021,N_5071);
xnor U5139 (N_5139,N_5075,N_5065);
nor U5140 (N_5140,N_5124,N_5032);
nor U5141 (N_5141,N_5010,N_5068);
nand U5142 (N_5142,N_5040,N_5016);
or U5143 (N_5143,N_5073,N_5056);
or U5144 (N_5144,N_5052,N_5057);
xor U5145 (N_5145,N_5046,N_5035);
or U5146 (N_5146,N_5050,N_5001);
nand U5147 (N_5147,N_5080,N_5054);
or U5148 (N_5148,N_5053,N_5003);
nor U5149 (N_5149,N_5077,N_5030);
xor U5150 (N_5150,N_5058,N_5067);
nor U5151 (N_5151,N_5072,N_5039);
nor U5152 (N_5152,N_5041,N_5031);
and U5153 (N_5153,N_5059,N_5081);
or U5154 (N_5154,N_5047,N_5011);
xor U5155 (N_5155,N_5066,N_5015);
nand U5156 (N_5156,N_5109,N_5038);
or U5157 (N_5157,N_5018,N_5069);
or U5158 (N_5158,N_5074,N_5123);
or U5159 (N_5159,N_5102,N_5091);
xor U5160 (N_5160,N_5061,N_5006);
nor U5161 (N_5161,N_5099,N_5078);
nand U5162 (N_5162,N_5007,N_5062);
nor U5163 (N_5163,N_5114,N_5117);
or U5164 (N_5164,N_5106,N_5024);
and U5165 (N_5165,N_5089,N_5098);
xnor U5166 (N_5166,N_5097,N_5043);
and U5167 (N_5167,N_5064,N_5060);
nand U5168 (N_5168,N_5036,N_5012);
and U5169 (N_5169,N_5013,N_5044);
and U5170 (N_5170,N_5105,N_5116);
nand U5171 (N_5171,N_5027,N_5008);
nand U5172 (N_5172,N_5000,N_5076);
or U5173 (N_5173,N_5029,N_5104);
or U5174 (N_5174,N_5025,N_5026);
nor U5175 (N_5175,N_5005,N_5002);
nand U5176 (N_5176,N_5023,N_5004);
nand U5177 (N_5177,N_5092,N_5079);
and U5178 (N_5178,N_5085,N_5110);
nor U5179 (N_5179,N_5118,N_5028);
and U5180 (N_5180,N_5017,N_5088);
nor U5181 (N_5181,N_5090,N_5037);
nor U5182 (N_5182,N_5022,N_5107);
and U5183 (N_5183,N_5020,N_5083);
or U5184 (N_5184,N_5070,N_5048);
or U5185 (N_5185,N_5119,N_5042);
xor U5186 (N_5186,N_5113,N_5084);
nand U5187 (N_5187,N_5082,N_5100);
nand U5188 (N_5188,N_5024,N_5002);
or U5189 (N_5189,N_5104,N_5074);
nor U5190 (N_5190,N_5091,N_5036);
and U5191 (N_5191,N_5119,N_5016);
or U5192 (N_5192,N_5025,N_5051);
xnor U5193 (N_5193,N_5026,N_5091);
nand U5194 (N_5194,N_5084,N_5014);
or U5195 (N_5195,N_5116,N_5043);
and U5196 (N_5196,N_5086,N_5022);
nand U5197 (N_5197,N_5100,N_5007);
or U5198 (N_5198,N_5084,N_5095);
nor U5199 (N_5199,N_5019,N_5001);
nand U5200 (N_5200,N_5122,N_5035);
and U5201 (N_5201,N_5009,N_5103);
nor U5202 (N_5202,N_5034,N_5004);
and U5203 (N_5203,N_5075,N_5063);
nand U5204 (N_5204,N_5085,N_5064);
and U5205 (N_5205,N_5073,N_5069);
and U5206 (N_5206,N_5119,N_5009);
nand U5207 (N_5207,N_5062,N_5027);
xor U5208 (N_5208,N_5031,N_5036);
nor U5209 (N_5209,N_5036,N_5010);
nor U5210 (N_5210,N_5010,N_5091);
and U5211 (N_5211,N_5066,N_5060);
xor U5212 (N_5212,N_5082,N_5034);
and U5213 (N_5213,N_5113,N_5056);
nor U5214 (N_5214,N_5053,N_5085);
or U5215 (N_5215,N_5061,N_5069);
nor U5216 (N_5216,N_5086,N_5091);
nor U5217 (N_5217,N_5111,N_5059);
xor U5218 (N_5218,N_5057,N_5006);
and U5219 (N_5219,N_5072,N_5118);
xor U5220 (N_5220,N_5087,N_5029);
xor U5221 (N_5221,N_5013,N_5043);
nand U5222 (N_5222,N_5052,N_5058);
and U5223 (N_5223,N_5052,N_5124);
xor U5224 (N_5224,N_5009,N_5110);
nand U5225 (N_5225,N_5019,N_5121);
nand U5226 (N_5226,N_5018,N_5012);
or U5227 (N_5227,N_5121,N_5043);
nand U5228 (N_5228,N_5078,N_5051);
and U5229 (N_5229,N_5090,N_5103);
xor U5230 (N_5230,N_5022,N_5121);
nand U5231 (N_5231,N_5053,N_5097);
and U5232 (N_5232,N_5088,N_5015);
or U5233 (N_5233,N_5119,N_5103);
or U5234 (N_5234,N_5056,N_5094);
xor U5235 (N_5235,N_5023,N_5027);
nand U5236 (N_5236,N_5043,N_5090);
nand U5237 (N_5237,N_5083,N_5057);
xnor U5238 (N_5238,N_5050,N_5038);
nand U5239 (N_5239,N_5084,N_5013);
and U5240 (N_5240,N_5063,N_5085);
xnor U5241 (N_5241,N_5034,N_5056);
nand U5242 (N_5242,N_5089,N_5004);
nand U5243 (N_5243,N_5059,N_5042);
nor U5244 (N_5244,N_5050,N_5004);
nand U5245 (N_5245,N_5090,N_5002);
nor U5246 (N_5246,N_5100,N_5117);
or U5247 (N_5247,N_5046,N_5026);
nand U5248 (N_5248,N_5045,N_5116);
or U5249 (N_5249,N_5062,N_5054);
and U5250 (N_5250,N_5130,N_5149);
or U5251 (N_5251,N_5236,N_5156);
nor U5252 (N_5252,N_5197,N_5131);
xor U5253 (N_5253,N_5135,N_5166);
and U5254 (N_5254,N_5221,N_5219);
nand U5255 (N_5255,N_5225,N_5184);
xnor U5256 (N_5256,N_5194,N_5158);
and U5257 (N_5257,N_5224,N_5195);
and U5258 (N_5258,N_5142,N_5244);
or U5259 (N_5259,N_5128,N_5230);
or U5260 (N_5260,N_5243,N_5211);
or U5261 (N_5261,N_5154,N_5126);
nor U5262 (N_5262,N_5191,N_5233);
nand U5263 (N_5263,N_5145,N_5138);
nor U5264 (N_5264,N_5231,N_5240);
and U5265 (N_5265,N_5201,N_5165);
or U5266 (N_5266,N_5205,N_5207);
or U5267 (N_5267,N_5190,N_5210);
nor U5268 (N_5268,N_5146,N_5151);
and U5269 (N_5269,N_5204,N_5183);
and U5270 (N_5270,N_5241,N_5143);
nor U5271 (N_5271,N_5159,N_5189);
xnor U5272 (N_5272,N_5152,N_5167);
nor U5273 (N_5273,N_5169,N_5200);
nand U5274 (N_5274,N_5223,N_5177);
and U5275 (N_5275,N_5247,N_5139);
xnor U5276 (N_5276,N_5181,N_5133);
nand U5277 (N_5277,N_5192,N_5215);
nor U5278 (N_5278,N_5127,N_5237);
and U5279 (N_5279,N_5188,N_5157);
or U5280 (N_5280,N_5208,N_5162);
or U5281 (N_5281,N_5137,N_5140);
and U5282 (N_5282,N_5220,N_5185);
nand U5283 (N_5283,N_5228,N_5175);
or U5284 (N_5284,N_5144,N_5213);
or U5285 (N_5285,N_5249,N_5172);
and U5286 (N_5286,N_5209,N_5217);
nand U5287 (N_5287,N_5239,N_5176);
nand U5288 (N_5288,N_5168,N_5198);
xor U5289 (N_5289,N_5235,N_5203);
nand U5290 (N_5290,N_5182,N_5163);
and U5291 (N_5291,N_5141,N_5155);
or U5292 (N_5292,N_5199,N_5147);
xor U5293 (N_5293,N_5212,N_5148);
and U5294 (N_5294,N_5193,N_5178);
nor U5295 (N_5295,N_5222,N_5227);
or U5296 (N_5296,N_5173,N_5248);
nand U5297 (N_5297,N_5164,N_5214);
or U5298 (N_5298,N_5187,N_5180);
xor U5299 (N_5299,N_5174,N_5136);
or U5300 (N_5300,N_5161,N_5171);
xor U5301 (N_5301,N_5246,N_5170);
xor U5302 (N_5302,N_5160,N_5242);
xnor U5303 (N_5303,N_5226,N_5229);
and U5304 (N_5304,N_5132,N_5232);
and U5305 (N_5305,N_5238,N_5129);
nand U5306 (N_5306,N_5179,N_5234);
or U5307 (N_5307,N_5125,N_5206);
nand U5308 (N_5308,N_5150,N_5186);
or U5309 (N_5309,N_5153,N_5216);
and U5310 (N_5310,N_5218,N_5202);
nor U5311 (N_5311,N_5245,N_5196);
and U5312 (N_5312,N_5134,N_5125);
nor U5313 (N_5313,N_5209,N_5238);
xor U5314 (N_5314,N_5195,N_5182);
nand U5315 (N_5315,N_5243,N_5181);
xnor U5316 (N_5316,N_5182,N_5161);
xor U5317 (N_5317,N_5144,N_5161);
and U5318 (N_5318,N_5184,N_5168);
nor U5319 (N_5319,N_5155,N_5184);
and U5320 (N_5320,N_5240,N_5223);
xnor U5321 (N_5321,N_5231,N_5155);
nor U5322 (N_5322,N_5146,N_5156);
xor U5323 (N_5323,N_5176,N_5215);
or U5324 (N_5324,N_5181,N_5226);
or U5325 (N_5325,N_5246,N_5202);
xnor U5326 (N_5326,N_5203,N_5144);
or U5327 (N_5327,N_5178,N_5191);
nand U5328 (N_5328,N_5139,N_5233);
and U5329 (N_5329,N_5215,N_5222);
nor U5330 (N_5330,N_5146,N_5175);
or U5331 (N_5331,N_5161,N_5157);
or U5332 (N_5332,N_5189,N_5237);
or U5333 (N_5333,N_5215,N_5239);
or U5334 (N_5334,N_5179,N_5232);
nor U5335 (N_5335,N_5130,N_5153);
nor U5336 (N_5336,N_5217,N_5185);
xor U5337 (N_5337,N_5153,N_5179);
nor U5338 (N_5338,N_5218,N_5138);
nand U5339 (N_5339,N_5206,N_5211);
or U5340 (N_5340,N_5217,N_5238);
nor U5341 (N_5341,N_5212,N_5196);
nand U5342 (N_5342,N_5215,N_5146);
nor U5343 (N_5343,N_5146,N_5130);
nand U5344 (N_5344,N_5218,N_5154);
and U5345 (N_5345,N_5242,N_5229);
or U5346 (N_5346,N_5234,N_5139);
and U5347 (N_5347,N_5249,N_5139);
nor U5348 (N_5348,N_5211,N_5196);
nand U5349 (N_5349,N_5172,N_5222);
nand U5350 (N_5350,N_5233,N_5169);
or U5351 (N_5351,N_5150,N_5171);
nand U5352 (N_5352,N_5212,N_5143);
xnor U5353 (N_5353,N_5160,N_5177);
xnor U5354 (N_5354,N_5204,N_5227);
nand U5355 (N_5355,N_5144,N_5168);
xnor U5356 (N_5356,N_5177,N_5153);
nor U5357 (N_5357,N_5218,N_5166);
nor U5358 (N_5358,N_5157,N_5182);
nor U5359 (N_5359,N_5203,N_5200);
or U5360 (N_5360,N_5166,N_5212);
nand U5361 (N_5361,N_5128,N_5137);
or U5362 (N_5362,N_5178,N_5194);
or U5363 (N_5363,N_5217,N_5210);
and U5364 (N_5364,N_5139,N_5212);
or U5365 (N_5365,N_5201,N_5157);
and U5366 (N_5366,N_5238,N_5176);
xor U5367 (N_5367,N_5140,N_5154);
or U5368 (N_5368,N_5137,N_5245);
and U5369 (N_5369,N_5184,N_5169);
or U5370 (N_5370,N_5240,N_5160);
nand U5371 (N_5371,N_5182,N_5138);
nand U5372 (N_5372,N_5174,N_5221);
nand U5373 (N_5373,N_5234,N_5162);
or U5374 (N_5374,N_5249,N_5215);
nand U5375 (N_5375,N_5344,N_5331);
or U5376 (N_5376,N_5343,N_5324);
xor U5377 (N_5377,N_5284,N_5290);
or U5378 (N_5378,N_5318,N_5306);
and U5379 (N_5379,N_5313,N_5312);
or U5380 (N_5380,N_5311,N_5326);
nand U5381 (N_5381,N_5280,N_5370);
or U5382 (N_5382,N_5329,N_5320);
xnor U5383 (N_5383,N_5265,N_5350);
nor U5384 (N_5384,N_5319,N_5362);
and U5385 (N_5385,N_5347,N_5295);
nor U5386 (N_5386,N_5337,N_5367);
and U5387 (N_5387,N_5307,N_5283);
and U5388 (N_5388,N_5271,N_5264);
and U5389 (N_5389,N_5273,N_5372);
or U5390 (N_5390,N_5261,N_5304);
or U5391 (N_5391,N_5276,N_5349);
nor U5392 (N_5392,N_5346,N_5341);
nand U5393 (N_5393,N_5285,N_5345);
and U5394 (N_5394,N_5374,N_5291);
or U5395 (N_5395,N_5321,N_5289);
xor U5396 (N_5396,N_5263,N_5302);
xor U5397 (N_5397,N_5373,N_5352);
nand U5398 (N_5398,N_5257,N_5323);
or U5399 (N_5399,N_5277,N_5369);
and U5400 (N_5400,N_5260,N_5348);
or U5401 (N_5401,N_5332,N_5254);
or U5402 (N_5402,N_5328,N_5357);
xor U5403 (N_5403,N_5355,N_5255);
nor U5404 (N_5404,N_5286,N_5269);
nor U5405 (N_5405,N_5365,N_5335);
and U5406 (N_5406,N_5292,N_5330);
and U5407 (N_5407,N_5259,N_5268);
nand U5408 (N_5408,N_5278,N_5342);
and U5409 (N_5409,N_5303,N_5363);
or U5410 (N_5410,N_5360,N_5305);
xnor U5411 (N_5411,N_5325,N_5275);
xnor U5412 (N_5412,N_5256,N_5250);
nand U5413 (N_5413,N_5359,N_5339);
and U5414 (N_5414,N_5356,N_5266);
xnor U5415 (N_5415,N_5270,N_5300);
or U5416 (N_5416,N_5267,N_5334);
and U5417 (N_5417,N_5252,N_5340);
or U5418 (N_5418,N_5327,N_5301);
or U5419 (N_5419,N_5358,N_5294);
and U5420 (N_5420,N_5366,N_5258);
and U5421 (N_5421,N_5314,N_5279);
nor U5422 (N_5422,N_5287,N_5351);
or U5423 (N_5423,N_5333,N_5297);
or U5424 (N_5424,N_5299,N_5272);
xnor U5425 (N_5425,N_5293,N_5322);
nor U5426 (N_5426,N_5371,N_5336);
nor U5427 (N_5427,N_5288,N_5282);
or U5428 (N_5428,N_5316,N_5368);
xor U5429 (N_5429,N_5317,N_5251);
xor U5430 (N_5430,N_5354,N_5281);
and U5431 (N_5431,N_5274,N_5310);
and U5432 (N_5432,N_5338,N_5361);
nor U5433 (N_5433,N_5315,N_5309);
xnor U5434 (N_5434,N_5308,N_5296);
xor U5435 (N_5435,N_5353,N_5262);
or U5436 (N_5436,N_5298,N_5253);
or U5437 (N_5437,N_5364,N_5259);
or U5438 (N_5438,N_5254,N_5299);
xnor U5439 (N_5439,N_5359,N_5332);
nand U5440 (N_5440,N_5275,N_5256);
xor U5441 (N_5441,N_5305,N_5266);
or U5442 (N_5442,N_5333,N_5306);
or U5443 (N_5443,N_5325,N_5293);
xnor U5444 (N_5444,N_5280,N_5312);
and U5445 (N_5445,N_5275,N_5257);
nor U5446 (N_5446,N_5265,N_5332);
or U5447 (N_5447,N_5286,N_5290);
or U5448 (N_5448,N_5351,N_5329);
and U5449 (N_5449,N_5317,N_5310);
nor U5450 (N_5450,N_5360,N_5288);
or U5451 (N_5451,N_5352,N_5346);
and U5452 (N_5452,N_5370,N_5339);
and U5453 (N_5453,N_5306,N_5348);
xor U5454 (N_5454,N_5353,N_5260);
nand U5455 (N_5455,N_5250,N_5284);
and U5456 (N_5456,N_5326,N_5372);
nand U5457 (N_5457,N_5258,N_5361);
nand U5458 (N_5458,N_5334,N_5345);
nand U5459 (N_5459,N_5268,N_5284);
nor U5460 (N_5460,N_5297,N_5304);
or U5461 (N_5461,N_5333,N_5311);
nand U5462 (N_5462,N_5320,N_5265);
xor U5463 (N_5463,N_5257,N_5350);
nor U5464 (N_5464,N_5325,N_5368);
and U5465 (N_5465,N_5305,N_5302);
and U5466 (N_5466,N_5352,N_5347);
nor U5467 (N_5467,N_5284,N_5296);
nand U5468 (N_5468,N_5314,N_5366);
xor U5469 (N_5469,N_5297,N_5337);
or U5470 (N_5470,N_5319,N_5282);
nand U5471 (N_5471,N_5250,N_5337);
xor U5472 (N_5472,N_5277,N_5307);
and U5473 (N_5473,N_5363,N_5260);
nand U5474 (N_5474,N_5337,N_5300);
or U5475 (N_5475,N_5251,N_5258);
xnor U5476 (N_5476,N_5256,N_5373);
or U5477 (N_5477,N_5277,N_5301);
or U5478 (N_5478,N_5292,N_5312);
and U5479 (N_5479,N_5365,N_5366);
nor U5480 (N_5480,N_5322,N_5251);
xor U5481 (N_5481,N_5274,N_5296);
or U5482 (N_5482,N_5330,N_5315);
or U5483 (N_5483,N_5279,N_5339);
or U5484 (N_5484,N_5273,N_5323);
xor U5485 (N_5485,N_5285,N_5317);
or U5486 (N_5486,N_5319,N_5299);
nor U5487 (N_5487,N_5345,N_5344);
nor U5488 (N_5488,N_5363,N_5329);
nand U5489 (N_5489,N_5314,N_5328);
nand U5490 (N_5490,N_5266,N_5296);
xor U5491 (N_5491,N_5278,N_5355);
and U5492 (N_5492,N_5291,N_5330);
and U5493 (N_5493,N_5361,N_5256);
xnor U5494 (N_5494,N_5338,N_5329);
nor U5495 (N_5495,N_5257,N_5349);
and U5496 (N_5496,N_5324,N_5264);
and U5497 (N_5497,N_5282,N_5312);
xor U5498 (N_5498,N_5335,N_5315);
and U5499 (N_5499,N_5299,N_5270);
and U5500 (N_5500,N_5425,N_5382);
nand U5501 (N_5501,N_5427,N_5496);
xor U5502 (N_5502,N_5412,N_5422);
and U5503 (N_5503,N_5376,N_5469);
or U5504 (N_5504,N_5430,N_5477);
nand U5505 (N_5505,N_5386,N_5457);
nor U5506 (N_5506,N_5399,N_5415);
and U5507 (N_5507,N_5476,N_5464);
or U5508 (N_5508,N_5470,N_5418);
xor U5509 (N_5509,N_5447,N_5421);
or U5510 (N_5510,N_5424,N_5486);
nor U5511 (N_5511,N_5456,N_5479);
nand U5512 (N_5512,N_5380,N_5393);
or U5513 (N_5513,N_5448,N_5450);
xnor U5514 (N_5514,N_5449,N_5442);
nor U5515 (N_5515,N_5391,N_5383);
or U5516 (N_5516,N_5451,N_5419);
or U5517 (N_5517,N_5499,N_5400);
or U5518 (N_5518,N_5410,N_5394);
or U5519 (N_5519,N_5481,N_5387);
nor U5520 (N_5520,N_5417,N_5453);
nand U5521 (N_5521,N_5379,N_5426);
nand U5522 (N_5522,N_5406,N_5388);
or U5523 (N_5523,N_5443,N_5460);
nand U5524 (N_5524,N_5401,N_5475);
xnor U5525 (N_5525,N_5395,N_5491);
nor U5526 (N_5526,N_5402,N_5471);
or U5527 (N_5527,N_5459,N_5467);
xor U5528 (N_5528,N_5468,N_5483);
xnor U5529 (N_5529,N_5434,N_5461);
and U5530 (N_5530,N_5408,N_5473);
or U5531 (N_5531,N_5493,N_5390);
nor U5532 (N_5532,N_5466,N_5455);
nand U5533 (N_5533,N_5431,N_5396);
nand U5534 (N_5534,N_5414,N_5433);
or U5535 (N_5535,N_5381,N_5484);
nand U5536 (N_5536,N_5403,N_5435);
and U5537 (N_5537,N_5398,N_5472);
nand U5538 (N_5538,N_5497,N_5438);
nand U5539 (N_5539,N_5404,N_5392);
nor U5540 (N_5540,N_5432,N_5428);
or U5541 (N_5541,N_5441,N_5405);
and U5542 (N_5542,N_5492,N_5384);
and U5543 (N_5543,N_5490,N_5482);
nor U5544 (N_5544,N_5411,N_5462);
xnor U5545 (N_5545,N_5389,N_5487);
nand U5546 (N_5546,N_5420,N_5440);
or U5547 (N_5547,N_5423,N_5429);
or U5548 (N_5548,N_5378,N_5494);
nand U5549 (N_5549,N_5445,N_5488);
xor U5550 (N_5550,N_5480,N_5436);
nand U5551 (N_5551,N_5375,N_5495);
and U5552 (N_5552,N_5413,N_5458);
xnor U5553 (N_5553,N_5498,N_5409);
nand U5554 (N_5554,N_5437,N_5444);
nand U5555 (N_5555,N_5446,N_5478);
nor U5556 (N_5556,N_5377,N_5416);
xnor U5557 (N_5557,N_5397,N_5463);
xor U5558 (N_5558,N_5452,N_5385);
nor U5559 (N_5559,N_5485,N_5454);
xnor U5560 (N_5560,N_5489,N_5474);
nor U5561 (N_5561,N_5439,N_5465);
nand U5562 (N_5562,N_5407,N_5419);
and U5563 (N_5563,N_5464,N_5473);
nand U5564 (N_5564,N_5402,N_5497);
nor U5565 (N_5565,N_5471,N_5447);
and U5566 (N_5566,N_5486,N_5384);
and U5567 (N_5567,N_5498,N_5411);
and U5568 (N_5568,N_5474,N_5443);
or U5569 (N_5569,N_5488,N_5474);
nand U5570 (N_5570,N_5436,N_5422);
nand U5571 (N_5571,N_5451,N_5473);
xor U5572 (N_5572,N_5382,N_5426);
or U5573 (N_5573,N_5415,N_5375);
nor U5574 (N_5574,N_5497,N_5410);
xor U5575 (N_5575,N_5498,N_5453);
nor U5576 (N_5576,N_5441,N_5436);
xor U5577 (N_5577,N_5484,N_5494);
nor U5578 (N_5578,N_5391,N_5454);
xnor U5579 (N_5579,N_5396,N_5424);
and U5580 (N_5580,N_5405,N_5466);
and U5581 (N_5581,N_5461,N_5429);
xnor U5582 (N_5582,N_5381,N_5414);
xor U5583 (N_5583,N_5379,N_5475);
xnor U5584 (N_5584,N_5392,N_5379);
nor U5585 (N_5585,N_5382,N_5385);
or U5586 (N_5586,N_5489,N_5496);
and U5587 (N_5587,N_5407,N_5447);
xor U5588 (N_5588,N_5447,N_5415);
nor U5589 (N_5589,N_5400,N_5439);
and U5590 (N_5590,N_5435,N_5409);
xnor U5591 (N_5591,N_5402,N_5478);
or U5592 (N_5592,N_5407,N_5460);
and U5593 (N_5593,N_5456,N_5465);
and U5594 (N_5594,N_5470,N_5433);
xor U5595 (N_5595,N_5477,N_5390);
xnor U5596 (N_5596,N_5389,N_5438);
xnor U5597 (N_5597,N_5489,N_5402);
nor U5598 (N_5598,N_5408,N_5446);
or U5599 (N_5599,N_5426,N_5400);
xor U5600 (N_5600,N_5385,N_5466);
or U5601 (N_5601,N_5454,N_5418);
or U5602 (N_5602,N_5471,N_5496);
nand U5603 (N_5603,N_5393,N_5394);
and U5604 (N_5604,N_5495,N_5488);
and U5605 (N_5605,N_5422,N_5448);
xnor U5606 (N_5606,N_5439,N_5475);
nand U5607 (N_5607,N_5413,N_5397);
nand U5608 (N_5608,N_5493,N_5489);
nand U5609 (N_5609,N_5430,N_5388);
or U5610 (N_5610,N_5430,N_5406);
nand U5611 (N_5611,N_5438,N_5382);
xnor U5612 (N_5612,N_5393,N_5385);
and U5613 (N_5613,N_5472,N_5480);
nand U5614 (N_5614,N_5385,N_5433);
and U5615 (N_5615,N_5442,N_5384);
nand U5616 (N_5616,N_5453,N_5390);
nand U5617 (N_5617,N_5429,N_5399);
nand U5618 (N_5618,N_5451,N_5402);
xor U5619 (N_5619,N_5472,N_5450);
or U5620 (N_5620,N_5440,N_5488);
nor U5621 (N_5621,N_5408,N_5485);
nand U5622 (N_5622,N_5435,N_5443);
or U5623 (N_5623,N_5486,N_5471);
nand U5624 (N_5624,N_5491,N_5408);
xor U5625 (N_5625,N_5502,N_5562);
nand U5626 (N_5626,N_5588,N_5544);
nand U5627 (N_5627,N_5511,N_5507);
or U5628 (N_5628,N_5537,N_5579);
nor U5629 (N_5629,N_5587,N_5596);
nor U5630 (N_5630,N_5549,N_5560);
and U5631 (N_5631,N_5548,N_5582);
nand U5632 (N_5632,N_5584,N_5590);
nand U5633 (N_5633,N_5514,N_5608);
xor U5634 (N_5634,N_5555,N_5536);
nand U5635 (N_5635,N_5541,N_5601);
nor U5636 (N_5636,N_5612,N_5615);
nand U5637 (N_5637,N_5605,N_5546);
nand U5638 (N_5638,N_5517,N_5570);
and U5639 (N_5639,N_5504,N_5581);
xor U5640 (N_5640,N_5550,N_5532);
nor U5641 (N_5641,N_5573,N_5571);
and U5642 (N_5642,N_5547,N_5586);
or U5643 (N_5643,N_5564,N_5540);
and U5644 (N_5644,N_5597,N_5523);
xor U5645 (N_5645,N_5613,N_5561);
or U5646 (N_5646,N_5500,N_5574);
xor U5647 (N_5647,N_5526,N_5553);
nor U5648 (N_5648,N_5521,N_5524);
nor U5649 (N_5649,N_5538,N_5614);
and U5650 (N_5650,N_5528,N_5611);
xor U5651 (N_5651,N_5505,N_5531);
nor U5652 (N_5652,N_5558,N_5515);
and U5653 (N_5653,N_5604,N_5616);
nor U5654 (N_5654,N_5545,N_5533);
or U5655 (N_5655,N_5535,N_5572);
and U5656 (N_5656,N_5525,N_5591);
and U5657 (N_5657,N_5583,N_5509);
and U5658 (N_5658,N_5522,N_5618);
nor U5659 (N_5659,N_5576,N_5617);
nor U5660 (N_5660,N_5543,N_5603);
or U5661 (N_5661,N_5580,N_5539);
xnor U5662 (N_5662,N_5551,N_5624);
xnor U5663 (N_5663,N_5503,N_5520);
xor U5664 (N_5664,N_5620,N_5534);
nor U5665 (N_5665,N_5585,N_5610);
or U5666 (N_5666,N_5518,N_5563);
or U5667 (N_5667,N_5552,N_5508);
or U5668 (N_5668,N_5606,N_5513);
xnor U5669 (N_5669,N_5565,N_5578);
and U5670 (N_5670,N_5512,N_5593);
nand U5671 (N_5671,N_5556,N_5609);
xor U5672 (N_5672,N_5530,N_5510);
xor U5673 (N_5673,N_5557,N_5516);
xor U5674 (N_5674,N_5600,N_5567);
nor U5675 (N_5675,N_5559,N_5592);
nand U5676 (N_5676,N_5566,N_5607);
nor U5677 (N_5677,N_5595,N_5589);
xnor U5678 (N_5678,N_5542,N_5619);
nor U5679 (N_5679,N_5602,N_5599);
nand U5680 (N_5680,N_5506,N_5623);
nor U5681 (N_5681,N_5501,N_5577);
or U5682 (N_5682,N_5527,N_5554);
and U5683 (N_5683,N_5569,N_5622);
or U5684 (N_5684,N_5568,N_5594);
nand U5685 (N_5685,N_5519,N_5529);
xor U5686 (N_5686,N_5575,N_5598);
nor U5687 (N_5687,N_5621,N_5514);
nor U5688 (N_5688,N_5523,N_5602);
nand U5689 (N_5689,N_5560,N_5525);
nor U5690 (N_5690,N_5527,N_5571);
nor U5691 (N_5691,N_5623,N_5621);
nand U5692 (N_5692,N_5613,N_5518);
nand U5693 (N_5693,N_5587,N_5579);
nand U5694 (N_5694,N_5560,N_5511);
nand U5695 (N_5695,N_5505,N_5546);
nor U5696 (N_5696,N_5564,N_5517);
nor U5697 (N_5697,N_5571,N_5594);
xor U5698 (N_5698,N_5514,N_5604);
and U5699 (N_5699,N_5586,N_5600);
xor U5700 (N_5700,N_5596,N_5552);
xnor U5701 (N_5701,N_5611,N_5568);
nor U5702 (N_5702,N_5502,N_5601);
nand U5703 (N_5703,N_5502,N_5505);
nand U5704 (N_5704,N_5624,N_5622);
or U5705 (N_5705,N_5547,N_5601);
or U5706 (N_5706,N_5622,N_5503);
or U5707 (N_5707,N_5608,N_5549);
nand U5708 (N_5708,N_5571,N_5598);
nor U5709 (N_5709,N_5624,N_5616);
xor U5710 (N_5710,N_5553,N_5540);
and U5711 (N_5711,N_5550,N_5582);
xnor U5712 (N_5712,N_5569,N_5520);
and U5713 (N_5713,N_5592,N_5552);
xor U5714 (N_5714,N_5512,N_5531);
and U5715 (N_5715,N_5535,N_5576);
nor U5716 (N_5716,N_5550,N_5540);
or U5717 (N_5717,N_5554,N_5543);
or U5718 (N_5718,N_5614,N_5606);
nor U5719 (N_5719,N_5565,N_5603);
nand U5720 (N_5720,N_5601,N_5575);
xor U5721 (N_5721,N_5530,N_5516);
nor U5722 (N_5722,N_5590,N_5567);
nand U5723 (N_5723,N_5536,N_5593);
nor U5724 (N_5724,N_5515,N_5500);
and U5725 (N_5725,N_5560,N_5613);
or U5726 (N_5726,N_5577,N_5603);
nand U5727 (N_5727,N_5534,N_5538);
xor U5728 (N_5728,N_5604,N_5598);
nand U5729 (N_5729,N_5568,N_5582);
xnor U5730 (N_5730,N_5551,N_5536);
nor U5731 (N_5731,N_5575,N_5539);
and U5732 (N_5732,N_5562,N_5552);
nand U5733 (N_5733,N_5605,N_5583);
and U5734 (N_5734,N_5616,N_5552);
xnor U5735 (N_5735,N_5578,N_5505);
xnor U5736 (N_5736,N_5612,N_5549);
nor U5737 (N_5737,N_5540,N_5591);
or U5738 (N_5738,N_5609,N_5620);
or U5739 (N_5739,N_5571,N_5540);
or U5740 (N_5740,N_5617,N_5505);
and U5741 (N_5741,N_5513,N_5505);
xor U5742 (N_5742,N_5604,N_5610);
nor U5743 (N_5743,N_5525,N_5563);
and U5744 (N_5744,N_5506,N_5577);
and U5745 (N_5745,N_5601,N_5576);
or U5746 (N_5746,N_5509,N_5554);
or U5747 (N_5747,N_5557,N_5585);
nor U5748 (N_5748,N_5543,N_5526);
or U5749 (N_5749,N_5512,N_5615);
and U5750 (N_5750,N_5724,N_5711);
nor U5751 (N_5751,N_5641,N_5697);
nand U5752 (N_5752,N_5680,N_5664);
xor U5753 (N_5753,N_5638,N_5744);
xnor U5754 (N_5754,N_5700,N_5642);
or U5755 (N_5755,N_5651,N_5745);
nand U5756 (N_5756,N_5632,N_5736);
xnor U5757 (N_5757,N_5729,N_5705);
xor U5758 (N_5758,N_5639,N_5643);
or U5759 (N_5759,N_5675,N_5673);
or U5760 (N_5760,N_5668,N_5683);
nand U5761 (N_5761,N_5626,N_5704);
and U5762 (N_5762,N_5715,N_5650);
and U5763 (N_5763,N_5699,N_5656);
nor U5764 (N_5764,N_5660,N_5701);
nor U5765 (N_5765,N_5671,N_5702);
nor U5766 (N_5766,N_5672,N_5659);
nor U5767 (N_5767,N_5730,N_5722);
xor U5768 (N_5768,N_5630,N_5713);
or U5769 (N_5769,N_5691,N_5709);
or U5770 (N_5770,N_5644,N_5688);
nor U5771 (N_5771,N_5686,N_5634);
nand U5772 (N_5772,N_5703,N_5637);
nand U5773 (N_5773,N_5749,N_5734);
nand U5774 (N_5774,N_5678,N_5652);
xor U5775 (N_5775,N_5716,N_5738);
nor U5776 (N_5776,N_5708,N_5714);
and U5777 (N_5777,N_5698,N_5733);
or U5778 (N_5778,N_5646,N_5658);
nor U5779 (N_5779,N_5710,N_5625);
and U5780 (N_5780,N_5747,N_5666);
nor U5781 (N_5781,N_5640,N_5720);
xor U5782 (N_5782,N_5627,N_5689);
nand U5783 (N_5783,N_5676,N_5655);
nor U5784 (N_5784,N_5739,N_5731);
and U5785 (N_5785,N_5670,N_5679);
or U5786 (N_5786,N_5693,N_5721);
nand U5787 (N_5787,N_5740,N_5706);
or U5788 (N_5788,N_5694,N_5647);
xor U5789 (N_5789,N_5674,N_5717);
or U5790 (N_5790,N_5685,N_5661);
nand U5791 (N_5791,N_5696,N_5727);
nand U5792 (N_5792,N_5737,N_5636);
or U5793 (N_5793,N_5682,N_5635);
or U5794 (N_5794,N_5665,N_5663);
and U5795 (N_5795,N_5648,N_5631);
nor U5796 (N_5796,N_5748,N_5645);
nand U5797 (N_5797,N_5633,N_5677);
nor U5798 (N_5798,N_5657,N_5725);
xor U5799 (N_5799,N_5695,N_5732);
or U5800 (N_5800,N_5723,N_5728);
xnor U5801 (N_5801,N_5649,N_5743);
and U5802 (N_5802,N_5681,N_5684);
and U5803 (N_5803,N_5741,N_5746);
xor U5804 (N_5804,N_5629,N_5718);
and U5805 (N_5805,N_5719,N_5690);
nor U5806 (N_5806,N_5726,N_5692);
and U5807 (N_5807,N_5662,N_5628);
xnor U5808 (N_5808,N_5735,N_5667);
nor U5809 (N_5809,N_5687,N_5707);
and U5810 (N_5810,N_5712,N_5669);
nor U5811 (N_5811,N_5653,N_5654);
or U5812 (N_5812,N_5742,N_5722);
and U5813 (N_5813,N_5646,N_5626);
xnor U5814 (N_5814,N_5659,N_5688);
nor U5815 (N_5815,N_5669,N_5653);
xor U5816 (N_5816,N_5701,N_5744);
and U5817 (N_5817,N_5728,N_5706);
and U5818 (N_5818,N_5692,N_5738);
and U5819 (N_5819,N_5628,N_5663);
nand U5820 (N_5820,N_5644,N_5734);
nor U5821 (N_5821,N_5655,N_5703);
and U5822 (N_5822,N_5637,N_5700);
nor U5823 (N_5823,N_5631,N_5666);
nand U5824 (N_5824,N_5720,N_5656);
and U5825 (N_5825,N_5710,N_5725);
or U5826 (N_5826,N_5666,N_5626);
nor U5827 (N_5827,N_5740,N_5631);
and U5828 (N_5828,N_5725,N_5730);
xor U5829 (N_5829,N_5673,N_5637);
nand U5830 (N_5830,N_5727,N_5748);
nor U5831 (N_5831,N_5700,N_5657);
xor U5832 (N_5832,N_5700,N_5639);
and U5833 (N_5833,N_5734,N_5729);
nor U5834 (N_5834,N_5645,N_5639);
xor U5835 (N_5835,N_5651,N_5749);
xnor U5836 (N_5836,N_5721,N_5639);
and U5837 (N_5837,N_5700,N_5660);
or U5838 (N_5838,N_5695,N_5636);
xnor U5839 (N_5839,N_5729,N_5627);
xor U5840 (N_5840,N_5715,N_5651);
or U5841 (N_5841,N_5671,N_5632);
or U5842 (N_5842,N_5747,N_5667);
xor U5843 (N_5843,N_5719,N_5724);
nand U5844 (N_5844,N_5695,N_5722);
and U5845 (N_5845,N_5657,N_5729);
xor U5846 (N_5846,N_5678,N_5698);
nor U5847 (N_5847,N_5699,N_5632);
nor U5848 (N_5848,N_5711,N_5638);
nand U5849 (N_5849,N_5663,N_5649);
nand U5850 (N_5850,N_5709,N_5648);
or U5851 (N_5851,N_5694,N_5730);
and U5852 (N_5852,N_5693,N_5669);
nand U5853 (N_5853,N_5676,N_5741);
nor U5854 (N_5854,N_5729,N_5712);
nand U5855 (N_5855,N_5694,N_5635);
nand U5856 (N_5856,N_5664,N_5660);
and U5857 (N_5857,N_5721,N_5673);
nor U5858 (N_5858,N_5697,N_5637);
nor U5859 (N_5859,N_5632,N_5661);
nor U5860 (N_5860,N_5719,N_5699);
or U5861 (N_5861,N_5740,N_5634);
nand U5862 (N_5862,N_5688,N_5748);
nand U5863 (N_5863,N_5643,N_5648);
xor U5864 (N_5864,N_5702,N_5639);
xnor U5865 (N_5865,N_5729,N_5666);
and U5866 (N_5866,N_5682,N_5667);
xor U5867 (N_5867,N_5679,N_5745);
and U5868 (N_5868,N_5698,N_5686);
nand U5869 (N_5869,N_5739,N_5704);
nor U5870 (N_5870,N_5736,N_5684);
xor U5871 (N_5871,N_5715,N_5744);
nand U5872 (N_5872,N_5633,N_5645);
and U5873 (N_5873,N_5696,N_5688);
and U5874 (N_5874,N_5688,N_5702);
xnor U5875 (N_5875,N_5837,N_5842);
xor U5876 (N_5876,N_5833,N_5818);
xor U5877 (N_5877,N_5873,N_5785);
or U5878 (N_5878,N_5872,N_5825);
xnor U5879 (N_5879,N_5808,N_5801);
nand U5880 (N_5880,N_5769,N_5786);
or U5881 (N_5881,N_5753,N_5826);
nor U5882 (N_5882,N_5772,N_5838);
or U5883 (N_5883,N_5779,N_5869);
xnor U5884 (N_5884,N_5821,N_5843);
and U5885 (N_5885,N_5800,N_5788);
nor U5886 (N_5886,N_5844,N_5806);
xor U5887 (N_5887,N_5804,N_5827);
and U5888 (N_5888,N_5755,N_5812);
and U5889 (N_5889,N_5834,N_5797);
and U5890 (N_5890,N_5773,N_5813);
nand U5891 (N_5891,N_5784,N_5836);
nor U5892 (N_5892,N_5858,N_5864);
and U5893 (N_5893,N_5771,N_5765);
nand U5894 (N_5894,N_5874,N_5865);
and U5895 (N_5895,N_5829,N_5761);
nor U5896 (N_5896,N_5811,N_5856);
nor U5897 (N_5897,N_5831,N_5850);
or U5898 (N_5898,N_5814,N_5840);
or U5899 (N_5899,N_5789,N_5790);
or U5900 (N_5900,N_5764,N_5857);
and U5901 (N_5901,N_5867,N_5863);
nand U5902 (N_5902,N_5762,N_5862);
xnor U5903 (N_5903,N_5841,N_5766);
and U5904 (N_5904,N_5763,N_5820);
xnor U5905 (N_5905,N_5871,N_5830);
nand U5906 (N_5906,N_5798,N_5822);
xnor U5907 (N_5907,N_5866,N_5832);
or U5908 (N_5908,N_5824,N_5802);
xor U5909 (N_5909,N_5810,N_5839);
and U5910 (N_5910,N_5855,N_5848);
and U5911 (N_5911,N_5754,N_5854);
nand U5912 (N_5912,N_5845,N_5851);
and U5913 (N_5913,N_5815,N_5809);
xor U5914 (N_5914,N_5777,N_5787);
and U5915 (N_5915,N_5782,N_5860);
nand U5916 (N_5916,N_5805,N_5795);
xnor U5917 (N_5917,N_5853,N_5783);
or U5918 (N_5918,N_5803,N_5852);
or U5919 (N_5919,N_5796,N_5776);
xnor U5920 (N_5920,N_5849,N_5868);
nor U5921 (N_5921,N_5835,N_5757);
and U5922 (N_5922,N_5770,N_5751);
and U5923 (N_5923,N_5870,N_5793);
or U5924 (N_5924,N_5861,N_5760);
and U5925 (N_5925,N_5767,N_5817);
or U5926 (N_5926,N_5828,N_5859);
or U5927 (N_5927,N_5775,N_5756);
xor U5928 (N_5928,N_5847,N_5792);
nand U5929 (N_5929,N_5823,N_5819);
nor U5930 (N_5930,N_5750,N_5794);
or U5931 (N_5931,N_5791,N_5781);
xnor U5932 (N_5932,N_5778,N_5752);
nor U5933 (N_5933,N_5799,N_5807);
xor U5934 (N_5934,N_5759,N_5816);
xnor U5935 (N_5935,N_5768,N_5758);
or U5936 (N_5936,N_5846,N_5774);
nor U5937 (N_5937,N_5780,N_5859);
and U5938 (N_5938,N_5766,N_5829);
or U5939 (N_5939,N_5773,N_5867);
nor U5940 (N_5940,N_5840,N_5860);
nand U5941 (N_5941,N_5798,N_5850);
nor U5942 (N_5942,N_5810,N_5856);
or U5943 (N_5943,N_5865,N_5778);
nor U5944 (N_5944,N_5770,N_5791);
nor U5945 (N_5945,N_5801,N_5829);
and U5946 (N_5946,N_5828,N_5762);
xor U5947 (N_5947,N_5787,N_5833);
and U5948 (N_5948,N_5814,N_5750);
nand U5949 (N_5949,N_5869,N_5781);
or U5950 (N_5950,N_5861,N_5852);
or U5951 (N_5951,N_5830,N_5800);
nor U5952 (N_5952,N_5848,N_5838);
nand U5953 (N_5953,N_5806,N_5803);
nor U5954 (N_5954,N_5856,N_5784);
and U5955 (N_5955,N_5809,N_5849);
and U5956 (N_5956,N_5871,N_5760);
xnor U5957 (N_5957,N_5797,N_5795);
xor U5958 (N_5958,N_5812,N_5771);
nand U5959 (N_5959,N_5807,N_5837);
and U5960 (N_5960,N_5864,N_5783);
nand U5961 (N_5961,N_5847,N_5828);
xor U5962 (N_5962,N_5845,N_5796);
and U5963 (N_5963,N_5823,N_5818);
and U5964 (N_5964,N_5821,N_5824);
xnor U5965 (N_5965,N_5847,N_5848);
nor U5966 (N_5966,N_5761,N_5752);
and U5967 (N_5967,N_5843,N_5818);
xnor U5968 (N_5968,N_5827,N_5767);
nand U5969 (N_5969,N_5873,N_5799);
nor U5970 (N_5970,N_5843,N_5782);
or U5971 (N_5971,N_5855,N_5769);
nor U5972 (N_5972,N_5801,N_5820);
nand U5973 (N_5973,N_5822,N_5751);
and U5974 (N_5974,N_5825,N_5855);
xnor U5975 (N_5975,N_5853,N_5776);
xnor U5976 (N_5976,N_5867,N_5866);
or U5977 (N_5977,N_5845,N_5819);
nor U5978 (N_5978,N_5796,N_5819);
or U5979 (N_5979,N_5865,N_5856);
xor U5980 (N_5980,N_5800,N_5815);
and U5981 (N_5981,N_5814,N_5862);
or U5982 (N_5982,N_5781,N_5853);
or U5983 (N_5983,N_5781,N_5772);
nor U5984 (N_5984,N_5861,N_5757);
or U5985 (N_5985,N_5787,N_5857);
nor U5986 (N_5986,N_5820,N_5773);
nor U5987 (N_5987,N_5839,N_5851);
nor U5988 (N_5988,N_5796,N_5805);
or U5989 (N_5989,N_5839,N_5836);
and U5990 (N_5990,N_5868,N_5870);
and U5991 (N_5991,N_5784,N_5806);
xnor U5992 (N_5992,N_5762,N_5798);
nand U5993 (N_5993,N_5771,N_5850);
nor U5994 (N_5994,N_5797,N_5839);
nor U5995 (N_5995,N_5764,N_5751);
nor U5996 (N_5996,N_5759,N_5754);
or U5997 (N_5997,N_5772,N_5757);
nor U5998 (N_5998,N_5810,N_5796);
xor U5999 (N_5999,N_5785,N_5791);
or U6000 (N_6000,N_5957,N_5945);
nor U6001 (N_6001,N_5978,N_5938);
nand U6002 (N_6002,N_5972,N_5890);
nand U6003 (N_6003,N_5966,N_5924);
and U6004 (N_6004,N_5923,N_5956);
and U6005 (N_6005,N_5991,N_5949);
nand U6006 (N_6006,N_5886,N_5941);
or U6007 (N_6007,N_5975,N_5946);
nor U6008 (N_6008,N_5982,N_5951);
nor U6009 (N_6009,N_5963,N_5934);
nand U6010 (N_6010,N_5900,N_5967);
xnor U6011 (N_6011,N_5944,N_5903);
nor U6012 (N_6012,N_5904,N_5898);
or U6013 (N_6013,N_5976,N_5888);
or U6014 (N_6014,N_5910,N_5895);
or U6015 (N_6015,N_5969,N_5893);
nor U6016 (N_6016,N_5960,N_5881);
xor U6017 (N_6017,N_5998,N_5914);
nor U6018 (N_6018,N_5902,N_5954);
nand U6019 (N_6019,N_5926,N_5961);
nor U6020 (N_6020,N_5891,N_5927);
nand U6021 (N_6021,N_5911,N_5933);
and U6022 (N_6022,N_5880,N_5901);
nand U6023 (N_6023,N_5896,N_5912);
xor U6024 (N_6024,N_5964,N_5878);
xnor U6025 (N_6025,N_5915,N_5905);
nor U6026 (N_6026,N_5875,N_5970);
or U6027 (N_6027,N_5980,N_5962);
or U6028 (N_6028,N_5936,N_5977);
xor U6029 (N_6029,N_5948,N_5879);
and U6030 (N_6030,N_5920,N_5928);
nand U6031 (N_6031,N_5882,N_5918);
nand U6032 (N_6032,N_5994,N_5993);
xnor U6033 (N_6033,N_5953,N_5917);
nand U6034 (N_6034,N_5939,N_5885);
and U6035 (N_6035,N_5990,N_5986);
nor U6036 (N_6036,N_5997,N_5894);
nor U6037 (N_6037,N_5947,N_5943);
nor U6038 (N_6038,N_5930,N_5908);
and U6039 (N_6039,N_5892,N_5884);
nand U6040 (N_6040,N_5989,N_5952);
nand U6041 (N_6041,N_5965,N_5995);
xnor U6042 (N_6042,N_5979,N_5897);
xor U6043 (N_6043,N_5935,N_5883);
or U6044 (N_6044,N_5973,N_5968);
nand U6045 (N_6045,N_5906,N_5974);
nand U6046 (N_6046,N_5983,N_5988);
nand U6047 (N_6047,N_5984,N_5950);
and U6048 (N_6048,N_5940,N_5959);
xor U6049 (N_6049,N_5971,N_5999);
xor U6050 (N_6050,N_5876,N_5922);
xor U6051 (N_6051,N_5981,N_5985);
and U6052 (N_6052,N_5889,N_5916);
and U6053 (N_6053,N_5887,N_5925);
nor U6054 (N_6054,N_5958,N_5931);
and U6055 (N_6055,N_5955,N_5913);
or U6056 (N_6056,N_5996,N_5907);
nand U6057 (N_6057,N_5932,N_5987);
and U6058 (N_6058,N_5929,N_5921);
nor U6059 (N_6059,N_5877,N_5992);
nand U6060 (N_6060,N_5937,N_5899);
or U6061 (N_6061,N_5942,N_5909);
nand U6062 (N_6062,N_5919,N_5965);
nand U6063 (N_6063,N_5919,N_5937);
nor U6064 (N_6064,N_5959,N_5932);
nor U6065 (N_6065,N_5879,N_5901);
nand U6066 (N_6066,N_5981,N_5980);
nand U6067 (N_6067,N_5877,N_5890);
nor U6068 (N_6068,N_5877,N_5994);
xnor U6069 (N_6069,N_5881,N_5981);
and U6070 (N_6070,N_5938,N_5888);
and U6071 (N_6071,N_5921,N_5901);
nand U6072 (N_6072,N_5964,N_5975);
xor U6073 (N_6073,N_5985,N_5902);
nor U6074 (N_6074,N_5933,N_5944);
and U6075 (N_6075,N_5939,N_5964);
and U6076 (N_6076,N_5957,N_5960);
xnor U6077 (N_6077,N_5919,N_5908);
nand U6078 (N_6078,N_5892,N_5979);
xnor U6079 (N_6079,N_5953,N_5876);
nor U6080 (N_6080,N_5886,N_5899);
and U6081 (N_6081,N_5905,N_5909);
or U6082 (N_6082,N_5946,N_5956);
or U6083 (N_6083,N_5989,N_5942);
and U6084 (N_6084,N_5952,N_5976);
or U6085 (N_6085,N_5968,N_5889);
nand U6086 (N_6086,N_5929,N_5957);
and U6087 (N_6087,N_5990,N_5910);
nand U6088 (N_6088,N_5905,N_5977);
xor U6089 (N_6089,N_5923,N_5898);
xnor U6090 (N_6090,N_5935,N_5972);
or U6091 (N_6091,N_5919,N_5954);
nor U6092 (N_6092,N_5903,N_5879);
xor U6093 (N_6093,N_5931,N_5936);
nor U6094 (N_6094,N_5932,N_5999);
and U6095 (N_6095,N_5904,N_5933);
or U6096 (N_6096,N_5939,N_5989);
and U6097 (N_6097,N_5991,N_5955);
or U6098 (N_6098,N_5882,N_5940);
or U6099 (N_6099,N_5910,N_5947);
or U6100 (N_6100,N_5927,N_5905);
nand U6101 (N_6101,N_5897,N_5939);
and U6102 (N_6102,N_5951,N_5899);
or U6103 (N_6103,N_5946,N_5968);
or U6104 (N_6104,N_5981,N_5984);
and U6105 (N_6105,N_5935,N_5939);
nor U6106 (N_6106,N_5876,N_5929);
nor U6107 (N_6107,N_5898,N_5900);
nor U6108 (N_6108,N_5934,N_5902);
or U6109 (N_6109,N_5908,N_5974);
and U6110 (N_6110,N_5947,N_5920);
nor U6111 (N_6111,N_5995,N_5940);
xor U6112 (N_6112,N_5976,N_5921);
and U6113 (N_6113,N_5954,N_5892);
or U6114 (N_6114,N_5932,N_5920);
nor U6115 (N_6115,N_5880,N_5878);
xnor U6116 (N_6116,N_5931,N_5916);
xnor U6117 (N_6117,N_5913,N_5928);
nand U6118 (N_6118,N_5942,N_5968);
or U6119 (N_6119,N_5963,N_5950);
and U6120 (N_6120,N_5962,N_5922);
nand U6121 (N_6121,N_5916,N_5970);
nor U6122 (N_6122,N_5945,N_5894);
or U6123 (N_6123,N_5893,N_5959);
or U6124 (N_6124,N_5902,N_5992);
xnor U6125 (N_6125,N_6116,N_6091);
and U6126 (N_6126,N_6001,N_6021);
or U6127 (N_6127,N_6039,N_6065);
nand U6128 (N_6128,N_6010,N_6105);
xnor U6129 (N_6129,N_6083,N_6085);
and U6130 (N_6130,N_6030,N_6038);
or U6131 (N_6131,N_6117,N_6017);
nor U6132 (N_6132,N_6054,N_6058);
nand U6133 (N_6133,N_6029,N_6004);
nor U6134 (N_6134,N_6063,N_6108);
nor U6135 (N_6135,N_6112,N_6095);
xor U6136 (N_6136,N_6056,N_6073);
and U6137 (N_6137,N_6013,N_6086);
and U6138 (N_6138,N_6032,N_6118);
nand U6139 (N_6139,N_6031,N_6080);
or U6140 (N_6140,N_6051,N_6075);
nor U6141 (N_6141,N_6099,N_6040);
nand U6142 (N_6142,N_6092,N_6077);
nor U6143 (N_6143,N_6067,N_6103);
or U6144 (N_6144,N_6050,N_6047);
and U6145 (N_6145,N_6101,N_6074);
nor U6146 (N_6146,N_6033,N_6023);
nand U6147 (N_6147,N_6113,N_6008);
nand U6148 (N_6148,N_6096,N_6070);
or U6149 (N_6149,N_6007,N_6082);
or U6150 (N_6150,N_6025,N_6093);
and U6151 (N_6151,N_6079,N_6006);
or U6152 (N_6152,N_6104,N_6015);
xnor U6153 (N_6153,N_6053,N_6024);
nand U6154 (N_6154,N_6061,N_6057);
and U6155 (N_6155,N_6016,N_6100);
xnor U6156 (N_6156,N_6120,N_6005);
or U6157 (N_6157,N_6114,N_6036);
and U6158 (N_6158,N_6109,N_6028);
xor U6159 (N_6159,N_6052,N_6018);
and U6160 (N_6160,N_6042,N_6000);
xor U6161 (N_6161,N_6123,N_6002);
nand U6162 (N_6162,N_6022,N_6048);
or U6163 (N_6163,N_6045,N_6026);
or U6164 (N_6164,N_6071,N_6044);
xor U6165 (N_6165,N_6019,N_6110);
nor U6166 (N_6166,N_6027,N_6102);
xnor U6167 (N_6167,N_6098,N_6059);
and U6168 (N_6168,N_6090,N_6078);
nand U6169 (N_6169,N_6011,N_6068);
or U6170 (N_6170,N_6062,N_6119);
nand U6171 (N_6171,N_6124,N_6049);
or U6172 (N_6172,N_6122,N_6020);
nand U6173 (N_6173,N_6014,N_6107);
and U6174 (N_6174,N_6060,N_6003);
nand U6175 (N_6175,N_6111,N_6076);
and U6176 (N_6176,N_6121,N_6012);
and U6177 (N_6177,N_6066,N_6089);
nand U6178 (N_6178,N_6115,N_6037);
nor U6179 (N_6179,N_6064,N_6097);
xnor U6180 (N_6180,N_6094,N_6081);
xnor U6181 (N_6181,N_6087,N_6035);
and U6182 (N_6182,N_6088,N_6106);
xor U6183 (N_6183,N_6055,N_6069);
xnor U6184 (N_6184,N_6041,N_6072);
or U6185 (N_6185,N_6043,N_6046);
nor U6186 (N_6186,N_6084,N_6009);
nor U6187 (N_6187,N_6034,N_6077);
nand U6188 (N_6188,N_6058,N_6068);
xnor U6189 (N_6189,N_6052,N_6093);
and U6190 (N_6190,N_6057,N_6051);
xnor U6191 (N_6191,N_6121,N_6114);
or U6192 (N_6192,N_6028,N_6043);
nor U6193 (N_6193,N_6057,N_6059);
nand U6194 (N_6194,N_6035,N_6027);
and U6195 (N_6195,N_6019,N_6000);
nor U6196 (N_6196,N_6057,N_6010);
nand U6197 (N_6197,N_6096,N_6024);
xor U6198 (N_6198,N_6067,N_6056);
xor U6199 (N_6199,N_6100,N_6056);
and U6200 (N_6200,N_6078,N_6035);
xor U6201 (N_6201,N_6076,N_6117);
and U6202 (N_6202,N_6003,N_6096);
nor U6203 (N_6203,N_6079,N_6106);
and U6204 (N_6204,N_6118,N_6002);
or U6205 (N_6205,N_6059,N_6079);
xnor U6206 (N_6206,N_6109,N_6124);
nand U6207 (N_6207,N_6008,N_6087);
and U6208 (N_6208,N_6101,N_6000);
nand U6209 (N_6209,N_6118,N_6030);
nor U6210 (N_6210,N_6093,N_6062);
xnor U6211 (N_6211,N_6002,N_6043);
or U6212 (N_6212,N_6003,N_6029);
and U6213 (N_6213,N_6060,N_6121);
xnor U6214 (N_6214,N_6103,N_6027);
nand U6215 (N_6215,N_6063,N_6034);
xor U6216 (N_6216,N_6050,N_6057);
and U6217 (N_6217,N_6062,N_6103);
and U6218 (N_6218,N_6000,N_6122);
nand U6219 (N_6219,N_6083,N_6123);
nor U6220 (N_6220,N_6006,N_6112);
or U6221 (N_6221,N_6066,N_6076);
and U6222 (N_6222,N_6015,N_6080);
or U6223 (N_6223,N_6071,N_6042);
and U6224 (N_6224,N_6054,N_6099);
xor U6225 (N_6225,N_6016,N_6036);
or U6226 (N_6226,N_6030,N_6089);
and U6227 (N_6227,N_6123,N_6089);
nand U6228 (N_6228,N_6070,N_6010);
or U6229 (N_6229,N_6063,N_6114);
nor U6230 (N_6230,N_6017,N_6075);
or U6231 (N_6231,N_6033,N_6053);
xnor U6232 (N_6232,N_6015,N_6074);
or U6233 (N_6233,N_6082,N_6109);
nand U6234 (N_6234,N_6005,N_6033);
nand U6235 (N_6235,N_6047,N_6027);
and U6236 (N_6236,N_6090,N_6111);
or U6237 (N_6237,N_6119,N_6034);
and U6238 (N_6238,N_6074,N_6005);
and U6239 (N_6239,N_6098,N_6013);
nand U6240 (N_6240,N_6006,N_6073);
xor U6241 (N_6241,N_6086,N_6123);
and U6242 (N_6242,N_6099,N_6056);
xor U6243 (N_6243,N_6043,N_6104);
and U6244 (N_6244,N_6075,N_6037);
or U6245 (N_6245,N_6088,N_6000);
xor U6246 (N_6246,N_6060,N_6040);
or U6247 (N_6247,N_6113,N_6069);
or U6248 (N_6248,N_6114,N_6101);
nor U6249 (N_6249,N_6017,N_6095);
xnor U6250 (N_6250,N_6228,N_6191);
or U6251 (N_6251,N_6237,N_6210);
nor U6252 (N_6252,N_6131,N_6202);
and U6253 (N_6253,N_6212,N_6248);
nor U6254 (N_6254,N_6141,N_6140);
xnor U6255 (N_6255,N_6243,N_6132);
or U6256 (N_6256,N_6157,N_6133);
xor U6257 (N_6257,N_6199,N_6227);
nor U6258 (N_6258,N_6139,N_6196);
nand U6259 (N_6259,N_6229,N_6171);
or U6260 (N_6260,N_6176,N_6205);
or U6261 (N_6261,N_6137,N_6226);
nand U6262 (N_6262,N_6236,N_6180);
xnor U6263 (N_6263,N_6167,N_6249);
xor U6264 (N_6264,N_6242,N_6129);
xor U6265 (N_6265,N_6239,N_6198);
or U6266 (N_6266,N_6145,N_6233);
or U6267 (N_6267,N_6216,N_6184);
nor U6268 (N_6268,N_6207,N_6183);
nand U6269 (N_6269,N_6221,N_6142);
nor U6270 (N_6270,N_6177,N_6219);
nor U6271 (N_6271,N_6159,N_6154);
or U6272 (N_6272,N_6163,N_6128);
nor U6273 (N_6273,N_6220,N_6200);
nand U6274 (N_6274,N_6218,N_6160);
nor U6275 (N_6275,N_6185,N_6195);
xnor U6276 (N_6276,N_6204,N_6156);
nand U6277 (N_6277,N_6193,N_6188);
or U6278 (N_6278,N_6223,N_6147);
and U6279 (N_6279,N_6224,N_6169);
or U6280 (N_6280,N_6225,N_6206);
nand U6281 (N_6281,N_6194,N_6125);
or U6282 (N_6282,N_6179,N_6162);
or U6283 (N_6283,N_6155,N_6208);
or U6284 (N_6284,N_6197,N_6209);
nor U6285 (N_6285,N_6135,N_6247);
nand U6286 (N_6286,N_6232,N_6241);
nand U6287 (N_6287,N_6222,N_6148);
nand U6288 (N_6288,N_6138,N_6245);
or U6289 (N_6289,N_6126,N_6130);
xnor U6290 (N_6290,N_6201,N_6234);
xnor U6291 (N_6291,N_6238,N_6165);
and U6292 (N_6292,N_6240,N_6144);
nand U6293 (N_6293,N_6164,N_6143);
and U6294 (N_6294,N_6181,N_6244);
nand U6295 (N_6295,N_6146,N_6149);
nand U6296 (N_6296,N_6215,N_6152);
or U6297 (N_6297,N_6186,N_6235);
nand U6298 (N_6298,N_6182,N_6189);
nor U6299 (N_6299,N_6136,N_6217);
nor U6300 (N_6300,N_6213,N_6187);
nand U6301 (N_6301,N_6178,N_6172);
nor U6302 (N_6302,N_6175,N_6168);
and U6303 (N_6303,N_6203,N_6158);
xnor U6304 (N_6304,N_6190,N_6150);
nand U6305 (N_6305,N_6231,N_6166);
and U6306 (N_6306,N_6211,N_6151);
or U6307 (N_6307,N_6174,N_6214);
nand U6308 (N_6308,N_6192,N_6173);
or U6309 (N_6309,N_6134,N_6127);
nor U6310 (N_6310,N_6161,N_6246);
nor U6311 (N_6311,N_6170,N_6153);
nand U6312 (N_6312,N_6230,N_6134);
or U6313 (N_6313,N_6152,N_6162);
and U6314 (N_6314,N_6167,N_6201);
nand U6315 (N_6315,N_6172,N_6145);
xor U6316 (N_6316,N_6129,N_6244);
and U6317 (N_6317,N_6167,N_6213);
and U6318 (N_6318,N_6198,N_6244);
xnor U6319 (N_6319,N_6227,N_6228);
and U6320 (N_6320,N_6126,N_6141);
xor U6321 (N_6321,N_6180,N_6202);
xnor U6322 (N_6322,N_6200,N_6236);
xor U6323 (N_6323,N_6166,N_6153);
or U6324 (N_6324,N_6227,N_6151);
nor U6325 (N_6325,N_6179,N_6205);
or U6326 (N_6326,N_6236,N_6167);
nor U6327 (N_6327,N_6160,N_6224);
xnor U6328 (N_6328,N_6210,N_6195);
or U6329 (N_6329,N_6137,N_6218);
or U6330 (N_6330,N_6141,N_6197);
nand U6331 (N_6331,N_6249,N_6182);
nand U6332 (N_6332,N_6234,N_6184);
nor U6333 (N_6333,N_6154,N_6139);
nand U6334 (N_6334,N_6190,N_6163);
nand U6335 (N_6335,N_6220,N_6208);
nand U6336 (N_6336,N_6151,N_6236);
and U6337 (N_6337,N_6132,N_6236);
nand U6338 (N_6338,N_6195,N_6177);
nor U6339 (N_6339,N_6137,N_6205);
or U6340 (N_6340,N_6246,N_6138);
xnor U6341 (N_6341,N_6170,N_6235);
or U6342 (N_6342,N_6140,N_6213);
nand U6343 (N_6343,N_6237,N_6230);
xnor U6344 (N_6344,N_6136,N_6200);
nand U6345 (N_6345,N_6160,N_6211);
xor U6346 (N_6346,N_6217,N_6125);
or U6347 (N_6347,N_6241,N_6205);
or U6348 (N_6348,N_6227,N_6174);
and U6349 (N_6349,N_6207,N_6205);
nor U6350 (N_6350,N_6222,N_6216);
xor U6351 (N_6351,N_6226,N_6223);
or U6352 (N_6352,N_6208,N_6197);
or U6353 (N_6353,N_6162,N_6142);
nor U6354 (N_6354,N_6134,N_6217);
and U6355 (N_6355,N_6144,N_6210);
nand U6356 (N_6356,N_6241,N_6131);
nor U6357 (N_6357,N_6134,N_6169);
nor U6358 (N_6358,N_6206,N_6158);
nor U6359 (N_6359,N_6241,N_6196);
nand U6360 (N_6360,N_6241,N_6214);
nand U6361 (N_6361,N_6198,N_6162);
or U6362 (N_6362,N_6137,N_6156);
nand U6363 (N_6363,N_6189,N_6146);
or U6364 (N_6364,N_6175,N_6152);
nor U6365 (N_6365,N_6136,N_6221);
or U6366 (N_6366,N_6219,N_6207);
nand U6367 (N_6367,N_6244,N_6206);
xor U6368 (N_6368,N_6249,N_6233);
and U6369 (N_6369,N_6185,N_6240);
or U6370 (N_6370,N_6138,N_6134);
xor U6371 (N_6371,N_6151,N_6174);
nand U6372 (N_6372,N_6181,N_6225);
or U6373 (N_6373,N_6228,N_6241);
nor U6374 (N_6374,N_6197,N_6158);
nand U6375 (N_6375,N_6295,N_6353);
nor U6376 (N_6376,N_6273,N_6326);
or U6377 (N_6377,N_6362,N_6320);
xor U6378 (N_6378,N_6276,N_6342);
or U6379 (N_6379,N_6297,N_6265);
or U6380 (N_6380,N_6256,N_6327);
nor U6381 (N_6381,N_6329,N_6251);
nand U6382 (N_6382,N_6345,N_6308);
xnor U6383 (N_6383,N_6344,N_6277);
and U6384 (N_6384,N_6284,N_6321);
nor U6385 (N_6385,N_6361,N_6260);
or U6386 (N_6386,N_6313,N_6339);
nor U6387 (N_6387,N_6351,N_6301);
and U6388 (N_6388,N_6266,N_6303);
nor U6389 (N_6389,N_6330,N_6271);
xnor U6390 (N_6390,N_6356,N_6358);
nor U6391 (N_6391,N_6348,N_6275);
nand U6392 (N_6392,N_6310,N_6258);
and U6393 (N_6393,N_6322,N_6281);
nand U6394 (N_6394,N_6305,N_6364);
or U6395 (N_6395,N_6370,N_6328);
and U6396 (N_6396,N_6357,N_6352);
and U6397 (N_6397,N_6367,N_6324);
xnor U6398 (N_6398,N_6331,N_6286);
xor U6399 (N_6399,N_6355,N_6254);
or U6400 (N_6400,N_6278,N_6270);
and U6401 (N_6401,N_6341,N_6253);
nor U6402 (N_6402,N_6261,N_6274);
and U6403 (N_6403,N_6334,N_6257);
nand U6404 (N_6404,N_6306,N_6293);
and U6405 (N_6405,N_6255,N_6309);
or U6406 (N_6406,N_6343,N_6285);
and U6407 (N_6407,N_6250,N_6314);
and U6408 (N_6408,N_6298,N_6282);
nor U6409 (N_6409,N_6349,N_6268);
or U6410 (N_6410,N_6325,N_6264);
or U6411 (N_6411,N_6299,N_6263);
or U6412 (N_6412,N_6290,N_6279);
or U6413 (N_6413,N_6307,N_6346);
nor U6414 (N_6414,N_6374,N_6323);
or U6415 (N_6415,N_6287,N_6368);
nand U6416 (N_6416,N_6291,N_6302);
xnor U6417 (N_6417,N_6336,N_6366);
nand U6418 (N_6418,N_6338,N_6288);
or U6419 (N_6419,N_6340,N_6335);
or U6420 (N_6420,N_6252,N_6354);
nand U6421 (N_6421,N_6304,N_6360);
and U6422 (N_6422,N_6259,N_6317);
nor U6423 (N_6423,N_6269,N_6371);
and U6424 (N_6424,N_6267,N_6332);
xnor U6425 (N_6425,N_6372,N_6272);
xnor U6426 (N_6426,N_6262,N_6311);
xnor U6427 (N_6427,N_6292,N_6283);
and U6428 (N_6428,N_6333,N_6363);
xor U6429 (N_6429,N_6350,N_6319);
nor U6430 (N_6430,N_6318,N_6300);
xnor U6431 (N_6431,N_6289,N_6280);
or U6432 (N_6432,N_6337,N_6347);
xnor U6433 (N_6433,N_6373,N_6365);
nor U6434 (N_6434,N_6312,N_6315);
nor U6435 (N_6435,N_6359,N_6316);
xor U6436 (N_6436,N_6296,N_6369);
and U6437 (N_6437,N_6294,N_6305);
and U6438 (N_6438,N_6324,N_6295);
or U6439 (N_6439,N_6288,N_6293);
and U6440 (N_6440,N_6342,N_6324);
nor U6441 (N_6441,N_6291,N_6365);
and U6442 (N_6442,N_6331,N_6275);
nor U6443 (N_6443,N_6370,N_6297);
and U6444 (N_6444,N_6339,N_6253);
or U6445 (N_6445,N_6314,N_6289);
nand U6446 (N_6446,N_6264,N_6282);
and U6447 (N_6447,N_6354,N_6345);
nand U6448 (N_6448,N_6287,N_6276);
nand U6449 (N_6449,N_6303,N_6317);
nand U6450 (N_6450,N_6368,N_6289);
nand U6451 (N_6451,N_6261,N_6319);
xor U6452 (N_6452,N_6295,N_6367);
nand U6453 (N_6453,N_6300,N_6290);
nor U6454 (N_6454,N_6255,N_6362);
nand U6455 (N_6455,N_6260,N_6307);
nor U6456 (N_6456,N_6265,N_6273);
nor U6457 (N_6457,N_6272,N_6359);
nand U6458 (N_6458,N_6347,N_6327);
nor U6459 (N_6459,N_6293,N_6284);
nor U6460 (N_6460,N_6288,N_6280);
nand U6461 (N_6461,N_6271,N_6295);
nand U6462 (N_6462,N_6284,N_6357);
nand U6463 (N_6463,N_6359,N_6270);
nor U6464 (N_6464,N_6258,N_6287);
nand U6465 (N_6465,N_6339,N_6282);
nor U6466 (N_6466,N_6333,N_6319);
and U6467 (N_6467,N_6284,N_6277);
nand U6468 (N_6468,N_6308,N_6250);
and U6469 (N_6469,N_6370,N_6306);
nor U6470 (N_6470,N_6259,N_6364);
and U6471 (N_6471,N_6284,N_6256);
nor U6472 (N_6472,N_6344,N_6279);
or U6473 (N_6473,N_6295,N_6371);
or U6474 (N_6474,N_6371,N_6350);
and U6475 (N_6475,N_6301,N_6270);
nor U6476 (N_6476,N_6351,N_6293);
xor U6477 (N_6477,N_6305,N_6349);
nand U6478 (N_6478,N_6336,N_6302);
and U6479 (N_6479,N_6333,N_6347);
nor U6480 (N_6480,N_6330,N_6374);
nand U6481 (N_6481,N_6342,N_6336);
and U6482 (N_6482,N_6312,N_6348);
nor U6483 (N_6483,N_6264,N_6346);
nor U6484 (N_6484,N_6354,N_6326);
nand U6485 (N_6485,N_6318,N_6275);
nand U6486 (N_6486,N_6347,N_6289);
nand U6487 (N_6487,N_6308,N_6365);
nor U6488 (N_6488,N_6304,N_6332);
nor U6489 (N_6489,N_6331,N_6258);
nor U6490 (N_6490,N_6356,N_6301);
xnor U6491 (N_6491,N_6262,N_6317);
and U6492 (N_6492,N_6306,N_6368);
nand U6493 (N_6493,N_6282,N_6349);
nand U6494 (N_6494,N_6325,N_6323);
and U6495 (N_6495,N_6319,N_6316);
and U6496 (N_6496,N_6345,N_6342);
xor U6497 (N_6497,N_6309,N_6360);
xnor U6498 (N_6498,N_6253,N_6271);
xor U6499 (N_6499,N_6290,N_6313);
nor U6500 (N_6500,N_6450,N_6471);
or U6501 (N_6501,N_6492,N_6482);
and U6502 (N_6502,N_6378,N_6414);
and U6503 (N_6503,N_6388,N_6498);
and U6504 (N_6504,N_6481,N_6427);
and U6505 (N_6505,N_6486,N_6434);
or U6506 (N_6506,N_6406,N_6380);
nand U6507 (N_6507,N_6474,N_6497);
xor U6508 (N_6508,N_6392,N_6453);
xor U6509 (N_6509,N_6396,N_6475);
nor U6510 (N_6510,N_6393,N_6459);
nand U6511 (N_6511,N_6466,N_6424);
and U6512 (N_6512,N_6465,N_6455);
nand U6513 (N_6513,N_6439,N_6401);
nor U6514 (N_6514,N_6404,N_6399);
and U6515 (N_6515,N_6488,N_6448);
xnor U6516 (N_6516,N_6377,N_6461);
nand U6517 (N_6517,N_6470,N_6469);
nor U6518 (N_6518,N_6467,N_6418);
nand U6519 (N_6519,N_6426,N_6412);
or U6520 (N_6520,N_6435,N_6460);
xnor U6521 (N_6521,N_6385,N_6383);
nand U6522 (N_6522,N_6487,N_6476);
nor U6523 (N_6523,N_6444,N_6387);
and U6524 (N_6524,N_6449,N_6391);
xnor U6525 (N_6525,N_6480,N_6405);
nand U6526 (N_6526,N_6400,N_6473);
and U6527 (N_6527,N_6457,N_6437);
or U6528 (N_6528,N_6389,N_6479);
and U6529 (N_6529,N_6451,N_6421);
nand U6530 (N_6530,N_6458,N_6398);
or U6531 (N_6531,N_6410,N_6411);
nor U6532 (N_6532,N_6384,N_6452);
and U6533 (N_6533,N_6485,N_6419);
xor U6534 (N_6534,N_6402,N_6490);
nand U6535 (N_6535,N_6495,N_6443);
nor U6536 (N_6536,N_6446,N_6409);
and U6537 (N_6537,N_6436,N_6472);
xor U6538 (N_6538,N_6403,N_6433);
and U6539 (N_6539,N_6441,N_6375);
xor U6540 (N_6540,N_6382,N_6491);
xnor U6541 (N_6541,N_6494,N_6408);
xnor U6542 (N_6542,N_6394,N_6447);
and U6543 (N_6543,N_6484,N_6454);
xor U6544 (N_6544,N_6496,N_6456);
nor U6545 (N_6545,N_6463,N_6483);
xor U6546 (N_6546,N_6376,N_6440);
xor U6547 (N_6547,N_6478,N_6397);
xnor U6548 (N_6548,N_6386,N_6417);
and U6549 (N_6549,N_6425,N_6445);
xor U6550 (N_6550,N_6468,N_6420);
or U6551 (N_6551,N_6477,N_6379);
xor U6552 (N_6552,N_6493,N_6489);
xor U6553 (N_6553,N_6416,N_6428);
or U6554 (N_6554,N_6430,N_6464);
nand U6555 (N_6555,N_6413,N_6395);
and U6556 (N_6556,N_6499,N_6432);
xnor U6557 (N_6557,N_6381,N_6422);
xnor U6558 (N_6558,N_6438,N_6462);
or U6559 (N_6559,N_6423,N_6431);
xnor U6560 (N_6560,N_6442,N_6390);
nor U6561 (N_6561,N_6415,N_6407);
or U6562 (N_6562,N_6429,N_6384);
or U6563 (N_6563,N_6431,N_6460);
nor U6564 (N_6564,N_6434,N_6426);
and U6565 (N_6565,N_6499,N_6476);
nand U6566 (N_6566,N_6418,N_6499);
xnor U6567 (N_6567,N_6441,N_6455);
nor U6568 (N_6568,N_6440,N_6460);
and U6569 (N_6569,N_6430,N_6419);
nor U6570 (N_6570,N_6454,N_6394);
or U6571 (N_6571,N_6440,N_6422);
nand U6572 (N_6572,N_6452,N_6499);
xnor U6573 (N_6573,N_6473,N_6478);
nand U6574 (N_6574,N_6455,N_6424);
nor U6575 (N_6575,N_6452,N_6450);
xnor U6576 (N_6576,N_6494,N_6393);
and U6577 (N_6577,N_6470,N_6390);
or U6578 (N_6578,N_6492,N_6392);
or U6579 (N_6579,N_6390,N_6438);
xor U6580 (N_6580,N_6391,N_6412);
and U6581 (N_6581,N_6421,N_6380);
nor U6582 (N_6582,N_6497,N_6427);
or U6583 (N_6583,N_6425,N_6388);
or U6584 (N_6584,N_6440,N_6382);
nor U6585 (N_6585,N_6419,N_6458);
xnor U6586 (N_6586,N_6492,N_6402);
nand U6587 (N_6587,N_6430,N_6488);
and U6588 (N_6588,N_6459,N_6394);
nand U6589 (N_6589,N_6402,N_6436);
xnor U6590 (N_6590,N_6479,N_6422);
or U6591 (N_6591,N_6410,N_6383);
nand U6592 (N_6592,N_6491,N_6470);
and U6593 (N_6593,N_6492,N_6484);
or U6594 (N_6594,N_6396,N_6488);
xnor U6595 (N_6595,N_6424,N_6423);
xor U6596 (N_6596,N_6426,N_6489);
and U6597 (N_6597,N_6399,N_6489);
and U6598 (N_6598,N_6390,N_6403);
or U6599 (N_6599,N_6428,N_6446);
nor U6600 (N_6600,N_6451,N_6423);
xor U6601 (N_6601,N_6389,N_6456);
xor U6602 (N_6602,N_6491,N_6418);
xor U6603 (N_6603,N_6434,N_6498);
or U6604 (N_6604,N_6379,N_6426);
xor U6605 (N_6605,N_6412,N_6496);
xor U6606 (N_6606,N_6464,N_6399);
nand U6607 (N_6607,N_6408,N_6452);
nor U6608 (N_6608,N_6465,N_6424);
nor U6609 (N_6609,N_6422,N_6472);
and U6610 (N_6610,N_6427,N_6435);
nor U6611 (N_6611,N_6432,N_6475);
and U6612 (N_6612,N_6490,N_6405);
nor U6613 (N_6613,N_6432,N_6453);
xor U6614 (N_6614,N_6403,N_6395);
nand U6615 (N_6615,N_6475,N_6451);
nor U6616 (N_6616,N_6481,N_6420);
xor U6617 (N_6617,N_6443,N_6401);
and U6618 (N_6618,N_6416,N_6384);
or U6619 (N_6619,N_6421,N_6492);
nand U6620 (N_6620,N_6477,N_6417);
nand U6621 (N_6621,N_6446,N_6385);
and U6622 (N_6622,N_6408,N_6446);
nand U6623 (N_6623,N_6464,N_6400);
nor U6624 (N_6624,N_6438,N_6378);
nand U6625 (N_6625,N_6601,N_6597);
and U6626 (N_6626,N_6529,N_6610);
nand U6627 (N_6627,N_6516,N_6503);
or U6628 (N_6628,N_6619,N_6595);
nand U6629 (N_6629,N_6510,N_6535);
and U6630 (N_6630,N_6572,N_6614);
xnor U6631 (N_6631,N_6616,N_6522);
xnor U6632 (N_6632,N_6570,N_6531);
or U6633 (N_6633,N_6590,N_6551);
nand U6634 (N_6634,N_6536,N_6555);
nand U6635 (N_6635,N_6602,N_6620);
and U6636 (N_6636,N_6589,N_6532);
nor U6637 (N_6637,N_6560,N_6534);
xnor U6638 (N_6638,N_6568,N_6507);
or U6639 (N_6639,N_6524,N_6611);
xor U6640 (N_6640,N_6506,N_6544);
nand U6641 (N_6641,N_6617,N_6598);
nand U6642 (N_6642,N_6517,N_6554);
xnor U6643 (N_6643,N_6530,N_6593);
nor U6644 (N_6644,N_6514,N_6591);
and U6645 (N_6645,N_6623,N_6586);
xor U6646 (N_6646,N_6608,N_6582);
xor U6647 (N_6647,N_6546,N_6594);
nor U6648 (N_6648,N_6548,N_6559);
nand U6649 (N_6649,N_6573,N_6520);
xnor U6650 (N_6650,N_6552,N_6508);
or U6651 (N_6651,N_6533,N_6553);
nor U6652 (N_6652,N_6605,N_6621);
nand U6653 (N_6653,N_6521,N_6624);
nand U6654 (N_6654,N_6606,N_6513);
nor U6655 (N_6655,N_6599,N_6509);
or U6656 (N_6656,N_6541,N_6504);
nor U6657 (N_6657,N_6566,N_6575);
nor U6658 (N_6658,N_6558,N_6549);
nand U6659 (N_6659,N_6528,N_6542);
or U6660 (N_6660,N_6584,N_6547);
xor U6661 (N_6661,N_6588,N_6592);
and U6662 (N_6662,N_6604,N_6525);
xor U6663 (N_6663,N_6526,N_6583);
and U6664 (N_6664,N_6515,N_6563);
or U6665 (N_6665,N_6569,N_6519);
or U6666 (N_6666,N_6613,N_6539);
and U6667 (N_6667,N_6587,N_6527);
xnor U6668 (N_6668,N_6543,N_6577);
xnor U6669 (N_6669,N_6580,N_6537);
nor U6670 (N_6670,N_6562,N_6561);
nand U6671 (N_6671,N_6603,N_6550);
nor U6672 (N_6672,N_6556,N_6567);
xor U6673 (N_6673,N_6615,N_6585);
nor U6674 (N_6674,N_6500,N_6596);
and U6675 (N_6675,N_6565,N_6612);
or U6676 (N_6676,N_6578,N_6523);
or U6677 (N_6677,N_6574,N_6518);
nor U6678 (N_6678,N_6607,N_6622);
xnor U6679 (N_6679,N_6511,N_6618);
xnor U6680 (N_6680,N_6579,N_6609);
or U6681 (N_6681,N_6545,N_6505);
xnor U6682 (N_6682,N_6501,N_6540);
or U6683 (N_6683,N_6576,N_6557);
xnor U6684 (N_6684,N_6564,N_6502);
or U6685 (N_6685,N_6538,N_6512);
nor U6686 (N_6686,N_6571,N_6581);
nor U6687 (N_6687,N_6600,N_6544);
or U6688 (N_6688,N_6594,N_6607);
and U6689 (N_6689,N_6550,N_6577);
or U6690 (N_6690,N_6519,N_6590);
and U6691 (N_6691,N_6611,N_6532);
nor U6692 (N_6692,N_6588,N_6507);
xor U6693 (N_6693,N_6607,N_6549);
and U6694 (N_6694,N_6526,N_6524);
nor U6695 (N_6695,N_6595,N_6568);
or U6696 (N_6696,N_6617,N_6520);
nand U6697 (N_6697,N_6505,N_6543);
and U6698 (N_6698,N_6507,N_6532);
or U6699 (N_6699,N_6610,N_6511);
nand U6700 (N_6700,N_6567,N_6590);
nor U6701 (N_6701,N_6513,N_6569);
nand U6702 (N_6702,N_6559,N_6545);
nand U6703 (N_6703,N_6578,N_6561);
and U6704 (N_6704,N_6605,N_6537);
or U6705 (N_6705,N_6519,N_6623);
nor U6706 (N_6706,N_6530,N_6501);
or U6707 (N_6707,N_6598,N_6507);
or U6708 (N_6708,N_6582,N_6546);
and U6709 (N_6709,N_6529,N_6561);
and U6710 (N_6710,N_6585,N_6557);
xor U6711 (N_6711,N_6569,N_6532);
nor U6712 (N_6712,N_6537,N_6574);
nor U6713 (N_6713,N_6547,N_6560);
xnor U6714 (N_6714,N_6529,N_6555);
and U6715 (N_6715,N_6624,N_6561);
and U6716 (N_6716,N_6548,N_6547);
and U6717 (N_6717,N_6553,N_6505);
or U6718 (N_6718,N_6574,N_6597);
and U6719 (N_6719,N_6555,N_6518);
nor U6720 (N_6720,N_6588,N_6598);
nor U6721 (N_6721,N_6594,N_6577);
or U6722 (N_6722,N_6599,N_6508);
xor U6723 (N_6723,N_6519,N_6602);
or U6724 (N_6724,N_6545,N_6526);
or U6725 (N_6725,N_6500,N_6566);
or U6726 (N_6726,N_6512,N_6554);
and U6727 (N_6727,N_6601,N_6578);
nor U6728 (N_6728,N_6527,N_6597);
nor U6729 (N_6729,N_6568,N_6549);
nor U6730 (N_6730,N_6528,N_6518);
nor U6731 (N_6731,N_6600,N_6608);
and U6732 (N_6732,N_6550,N_6534);
xnor U6733 (N_6733,N_6612,N_6567);
xnor U6734 (N_6734,N_6608,N_6577);
nor U6735 (N_6735,N_6586,N_6571);
or U6736 (N_6736,N_6566,N_6550);
or U6737 (N_6737,N_6552,N_6527);
or U6738 (N_6738,N_6614,N_6620);
or U6739 (N_6739,N_6597,N_6506);
xnor U6740 (N_6740,N_6519,N_6560);
and U6741 (N_6741,N_6519,N_6518);
xor U6742 (N_6742,N_6585,N_6522);
xnor U6743 (N_6743,N_6600,N_6547);
or U6744 (N_6744,N_6577,N_6616);
and U6745 (N_6745,N_6587,N_6542);
nor U6746 (N_6746,N_6548,N_6551);
xor U6747 (N_6747,N_6561,N_6505);
xnor U6748 (N_6748,N_6624,N_6546);
xor U6749 (N_6749,N_6530,N_6598);
xor U6750 (N_6750,N_6628,N_6705);
nor U6751 (N_6751,N_6675,N_6749);
nor U6752 (N_6752,N_6687,N_6661);
nor U6753 (N_6753,N_6657,N_6711);
and U6754 (N_6754,N_6654,N_6713);
nand U6755 (N_6755,N_6692,N_6639);
or U6756 (N_6756,N_6652,N_6698);
nand U6757 (N_6757,N_6627,N_6674);
and U6758 (N_6758,N_6699,N_6631);
nor U6759 (N_6759,N_6633,N_6647);
nand U6760 (N_6760,N_6671,N_6640);
and U6761 (N_6761,N_6703,N_6745);
xnor U6762 (N_6762,N_6634,N_6715);
xor U6763 (N_6763,N_6681,N_6744);
and U6764 (N_6764,N_6740,N_6697);
nor U6765 (N_6765,N_6696,N_6719);
or U6766 (N_6766,N_6650,N_6704);
nor U6767 (N_6767,N_6742,N_6673);
xnor U6768 (N_6768,N_6638,N_6667);
or U6769 (N_6769,N_6669,N_6739);
nand U6770 (N_6770,N_6701,N_6645);
nor U6771 (N_6771,N_6642,N_6717);
or U6772 (N_6772,N_6730,N_6664);
nand U6773 (N_6773,N_6649,N_6714);
nor U6774 (N_6774,N_6716,N_6648);
and U6775 (N_6775,N_6731,N_6709);
nor U6776 (N_6776,N_6643,N_6695);
nor U6777 (N_6777,N_6626,N_6637);
xnor U6778 (N_6778,N_6666,N_6712);
nand U6779 (N_6779,N_6720,N_6660);
nand U6780 (N_6780,N_6693,N_6736);
nand U6781 (N_6781,N_6726,N_6632);
xor U6782 (N_6782,N_6700,N_6656);
or U6783 (N_6783,N_6646,N_6672);
and U6784 (N_6784,N_6702,N_6694);
and U6785 (N_6785,N_6734,N_6741);
nor U6786 (N_6786,N_6680,N_6733);
and U6787 (N_6787,N_6724,N_6729);
xor U6788 (N_6788,N_6651,N_6722);
or U6789 (N_6789,N_6653,N_6636);
nor U6790 (N_6790,N_6641,N_6629);
and U6791 (N_6791,N_6748,N_6728);
xor U6792 (N_6792,N_6735,N_6689);
or U6793 (N_6793,N_6679,N_6644);
and U6794 (N_6794,N_6686,N_6706);
xor U6795 (N_6795,N_6710,N_6708);
nor U6796 (N_6796,N_6663,N_6658);
nand U6797 (N_6797,N_6746,N_6668);
nand U6798 (N_6798,N_6630,N_6662);
or U6799 (N_6799,N_6718,N_6691);
or U6800 (N_6800,N_6625,N_6665);
nor U6801 (N_6801,N_6688,N_6683);
xor U6802 (N_6802,N_6721,N_6747);
or U6803 (N_6803,N_6743,N_6737);
xnor U6804 (N_6804,N_6684,N_6678);
or U6805 (N_6805,N_6670,N_6682);
nand U6806 (N_6806,N_6727,N_6723);
xor U6807 (N_6807,N_6685,N_6738);
xor U6808 (N_6808,N_6690,N_6732);
nor U6809 (N_6809,N_6635,N_6676);
and U6810 (N_6810,N_6677,N_6655);
nand U6811 (N_6811,N_6707,N_6659);
xnor U6812 (N_6812,N_6725,N_6669);
or U6813 (N_6813,N_6650,N_6695);
nor U6814 (N_6814,N_6637,N_6650);
xnor U6815 (N_6815,N_6702,N_6689);
nor U6816 (N_6816,N_6638,N_6700);
nor U6817 (N_6817,N_6694,N_6677);
or U6818 (N_6818,N_6668,N_6749);
xnor U6819 (N_6819,N_6634,N_6708);
nor U6820 (N_6820,N_6679,N_6641);
and U6821 (N_6821,N_6656,N_6644);
and U6822 (N_6822,N_6748,N_6670);
xor U6823 (N_6823,N_6649,N_6636);
xnor U6824 (N_6824,N_6663,N_6743);
and U6825 (N_6825,N_6676,N_6641);
nand U6826 (N_6826,N_6629,N_6706);
xnor U6827 (N_6827,N_6657,N_6649);
nand U6828 (N_6828,N_6730,N_6628);
nand U6829 (N_6829,N_6700,N_6632);
nor U6830 (N_6830,N_6697,N_6748);
and U6831 (N_6831,N_6636,N_6657);
nor U6832 (N_6832,N_6647,N_6686);
and U6833 (N_6833,N_6653,N_6722);
nor U6834 (N_6834,N_6725,N_6628);
xnor U6835 (N_6835,N_6705,N_6633);
and U6836 (N_6836,N_6701,N_6665);
or U6837 (N_6837,N_6680,N_6667);
xor U6838 (N_6838,N_6679,N_6658);
and U6839 (N_6839,N_6629,N_6727);
or U6840 (N_6840,N_6648,N_6704);
or U6841 (N_6841,N_6746,N_6685);
and U6842 (N_6842,N_6677,N_6702);
xnor U6843 (N_6843,N_6640,N_6704);
nand U6844 (N_6844,N_6738,N_6676);
nor U6845 (N_6845,N_6668,N_6640);
and U6846 (N_6846,N_6664,N_6628);
nand U6847 (N_6847,N_6681,N_6661);
or U6848 (N_6848,N_6734,N_6728);
and U6849 (N_6849,N_6659,N_6716);
or U6850 (N_6850,N_6628,N_6704);
xnor U6851 (N_6851,N_6644,N_6706);
nor U6852 (N_6852,N_6658,N_6629);
or U6853 (N_6853,N_6695,N_6699);
nor U6854 (N_6854,N_6727,N_6704);
nand U6855 (N_6855,N_6732,N_6678);
nor U6856 (N_6856,N_6650,N_6719);
or U6857 (N_6857,N_6707,N_6739);
and U6858 (N_6858,N_6744,N_6704);
and U6859 (N_6859,N_6718,N_6675);
and U6860 (N_6860,N_6698,N_6744);
and U6861 (N_6861,N_6626,N_6740);
or U6862 (N_6862,N_6665,N_6747);
xor U6863 (N_6863,N_6660,N_6632);
nor U6864 (N_6864,N_6656,N_6675);
xor U6865 (N_6865,N_6654,N_6663);
or U6866 (N_6866,N_6729,N_6653);
or U6867 (N_6867,N_6749,N_6729);
nand U6868 (N_6868,N_6749,N_6644);
or U6869 (N_6869,N_6677,N_6745);
and U6870 (N_6870,N_6665,N_6734);
xnor U6871 (N_6871,N_6659,N_6698);
and U6872 (N_6872,N_6727,N_6666);
nand U6873 (N_6873,N_6735,N_6734);
nor U6874 (N_6874,N_6695,N_6739);
xor U6875 (N_6875,N_6861,N_6782);
or U6876 (N_6876,N_6847,N_6836);
xnor U6877 (N_6877,N_6820,N_6829);
xor U6878 (N_6878,N_6853,N_6802);
nor U6879 (N_6879,N_6821,N_6810);
and U6880 (N_6880,N_6839,N_6794);
or U6881 (N_6881,N_6795,N_6805);
nor U6882 (N_6882,N_6769,N_6848);
or U6883 (N_6883,N_6758,N_6830);
nor U6884 (N_6884,N_6763,N_6822);
or U6885 (N_6885,N_6768,N_6801);
nand U6886 (N_6886,N_6854,N_6779);
and U6887 (N_6887,N_6811,N_6774);
or U6888 (N_6888,N_6814,N_6766);
and U6889 (N_6889,N_6786,N_6813);
nand U6890 (N_6890,N_6784,N_6852);
nor U6891 (N_6891,N_6833,N_6873);
nand U6892 (N_6892,N_6872,N_6751);
xor U6893 (N_6893,N_6849,N_6825);
nor U6894 (N_6894,N_6765,N_6870);
and U6895 (N_6895,N_6753,N_6796);
xor U6896 (N_6896,N_6824,N_6770);
xnor U6897 (N_6897,N_6783,N_6775);
xor U6898 (N_6898,N_6868,N_6874);
xnor U6899 (N_6899,N_6818,N_6855);
nor U6900 (N_6900,N_6759,N_6806);
nor U6901 (N_6901,N_6760,N_6817);
nand U6902 (N_6902,N_6871,N_6793);
or U6903 (N_6903,N_6755,N_6797);
or U6904 (N_6904,N_6842,N_6819);
nor U6905 (N_6905,N_6752,N_6764);
nand U6906 (N_6906,N_6859,N_6767);
xnor U6907 (N_6907,N_6780,N_6851);
or U6908 (N_6908,N_6867,N_6777);
and U6909 (N_6909,N_6808,N_6812);
or U6910 (N_6910,N_6807,N_6773);
xor U6911 (N_6911,N_6831,N_6815);
xor U6912 (N_6912,N_6772,N_6864);
nor U6913 (N_6913,N_6860,N_6840);
or U6914 (N_6914,N_6866,N_6800);
xnor U6915 (N_6915,N_6844,N_6809);
xnor U6916 (N_6916,N_6863,N_6750);
and U6917 (N_6917,N_6835,N_6827);
nor U6918 (N_6918,N_6798,N_6865);
xnor U6919 (N_6919,N_6771,N_6841);
nand U6920 (N_6920,N_6778,N_6799);
xnor U6921 (N_6921,N_6856,N_6869);
xnor U6922 (N_6922,N_6845,N_6787);
and U6923 (N_6923,N_6857,N_6843);
xnor U6924 (N_6924,N_6781,N_6754);
nand U6925 (N_6925,N_6789,N_6823);
nand U6926 (N_6926,N_6785,N_6862);
nor U6927 (N_6927,N_6762,N_6828);
nand U6928 (N_6928,N_6834,N_6846);
and U6929 (N_6929,N_6837,N_6832);
nand U6930 (N_6930,N_6792,N_6790);
nor U6931 (N_6931,N_6756,N_6761);
nor U6932 (N_6932,N_6791,N_6803);
xnor U6933 (N_6933,N_6776,N_6826);
or U6934 (N_6934,N_6804,N_6838);
and U6935 (N_6935,N_6816,N_6788);
and U6936 (N_6936,N_6757,N_6850);
xor U6937 (N_6937,N_6858,N_6830);
nand U6938 (N_6938,N_6851,N_6788);
and U6939 (N_6939,N_6853,N_6869);
nor U6940 (N_6940,N_6756,N_6769);
and U6941 (N_6941,N_6783,N_6863);
and U6942 (N_6942,N_6803,N_6808);
xnor U6943 (N_6943,N_6766,N_6794);
nor U6944 (N_6944,N_6753,N_6850);
xor U6945 (N_6945,N_6864,N_6776);
and U6946 (N_6946,N_6818,N_6831);
nand U6947 (N_6947,N_6790,N_6781);
or U6948 (N_6948,N_6819,N_6853);
or U6949 (N_6949,N_6817,N_6770);
xor U6950 (N_6950,N_6783,N_6802);
and U6951 (N_6951,N_6770,N_6790);
nand U6952 (N_6952,N_6852,N_6796);
or U6953 (N_6953,N_6775,N_6800);
nor U6954 (N_6954,N_6777,N_6828);
and U6955 (N_6955,N_6838,N_6824);
nor U6956 (N_6956,N_6778,N_6769);
xnor U6957 (N_6957,N_6787,N_6782);
nand U6958 (N_6958,N_6867,N_6828);
nor U6959 (N_6959,N_6829,N_6852);
nor U6960 (N_6960,N_6790,N_6783);
or U6961 (N_6961,N_6816,N_6825);
or U6962 (N_6962,N_6853,N_6805);
or U6963 (N_6963,N_6851,N_6772);
nor U6964 (N_6964,N_6820,N_6791);
xor U6965 (N_6965,N_6782,N_6756);
nand U6966 (N_6966,N_6808,N_6864);
nand U6967 (N_6967,N_6813,N_6784);
xnor U6968 (N_6968,N_6847,N_6799);
nor U6969 (N_6969,N_6817,N_6835);
xnor U6970 (N_6970,N_6838,N_6816);
nand U6971 (N_6971,N_6834,N_6814);
xor U6972 (N_6972,N_6843,N_6864);
nand U6973 (N_6973,N_6770,N_6808);
or U6974 (N_6974,N_6774,N_6818);
and U6975 (N_6975,N_6821,N_6792);
and U6976 (N_6976,N_6772,N_6797);
nor U6977 (N_6977,N_6802,N_6836);
or U6978 (N_6978,N_6794,N_6859);
nand U6979 (N_6979,N_6770,N_6869);
and U6980 (N_6980,N_6750,N_6843);
nor U6981 (N_6981,N_6755,N_6836);
xnor U6982 (N_6982,N_6832,N_6836);
xnor U6983 (N_6983,N_6848,N_6856);
and U6984 (N_6984,N_6772,N_6823);
or U6985 (N_6985,N_6855,N_6766);
xor U6986 (N_6986,N_6835,N_6841);
and U6987 (N_6987,N_6785,N_6754);
nand U6988 (N_6988,N_6856,N_6873);
nor U6989 (N_6989,N_6848,N_6786);
nor U6990 (N_6990,N_6762,N_6811);
xnor U6991 (N_6991,N_6810,N_6758);
and U6992 (N_6992,N_6825,N_6845);
xor U6993 (N_6993,N_6777,N_6761);
or U6994 (N_6994,N_6769,N_6761);
xor U6995 (N_6995,N_6780,N_6790);
xor U6996 (N_6996,N_6757,N_6871);
or U6997 (N_6997,N_6854,N_6755);
nor U6998 (N_6998,N_6809,N_6860);
and U6999 (N_6999,N_6820,N_6789);
or U7000 (N_7000,N_6923,N_6921);
nand U7001 (N_7001,N_6978,N_6958);
nand U7002 (N_7002,N_6961,N_6919);
xnor U7003 (N_7003,N_6889,N_6971);
or U7004 (N_7004,N_6894,N_6875);
or U7005 (N_7005,N_6907,N_6989);
xor U7006 (N_7006,N_6892,N_6903);
or U7007 (N_7007,N_6987,N_6933);
nor U7008 (N_7008,N_6905,N_6985);
xnor U7009 (N_7009,N_6886,N_6993);
nand U7010 (N_7010,N_6947,N_6898);
nor U7011 (N_7011,N_6897,N_6916);
xnor U7012 (N_7012,N_6945,N_6992);
nand U7013 (N_7013,N_6977,N_6942);
or U7014 (N_7014,N_6944,N_6909);
nand U7015 (N_7015,N_6952,N_6928);
xor U7016 (N_7016,N_6918,N_6984);
xor U7017 (N_7017,N_6880,N_6973);
nor U7018 (N_7018,N_6899,N_6920);
and U7019 (N_7019,N_6887,N_6934);
nor U7020 (N_7020,N_6990,N_6962);
nand U7021 (N_7021,N_6998,N_6983);
and U7022 (N_7022,N_6884,N_6954);
nand U7023 (N_7023,N_6883,N_6948);
nand U7024 (N_7024,N_6912,N_6915);
nor U7025 (N_7025,N_6931,N_6996);
nand U7026 (N_7026,N_6994,N_6917);
and U7027 (N_7027,N_6890,N_6893);
xnor U7028 (N_7028,N_6911,N_6943);
nand U7029 (N_7029,N_6995,N_6901);
nor U7030 (N_7030,N_6937,N_6949);
nand U7031 (N_7031,N_6950,N_6902);
nand U7032 (N_7032,N_6910,N_6965);
and U7033 (N_7033,N_6975,N_6972);
and U7034 (N_7034,N_6888,N_6939);
xor U7035 (N_7035,N_6963,N_6967);
nand U7036 (N_7036,N_6927,N_6960);
nand U7037 (N_7037,N_6906,N_6951);
or U7038 (N_7038,N_6974,N_6986);
and U7039 (N_7039,N_6957,N_6908);
nor U7040 (N_7040,N_6926,N_6879);
nor U7041 (N_7041,N_6913,N_6964);
xor U7042 (N_7042,N_6999,N_6885);
xnor U7043 (N_7043,N_6922,N_6980);
xor U7044 (N_7044,N_6955,N_6997);
and U7045 (N_7045,N_6925,N_6932);
and U7046 (N_7046,N_6976,N_6991);
and U7047 (N_7047,N_6935,N_6970);
nand U7048 (N_7048,N_6876,N_6968);
nand U7049 (N_7049,N_6966,N_6941);
nor U7050 (N_7050,N_6882,N_6959);
xnor U7051 (N_7051,N_6895,N_6982);
xnor U7052 (N_7052,N_6969,N_6878);
nand U7053 (N_7053,N_6881,N_6896);
or U7054 (N_7054,N_6953,N_6930);
xnor U7055 (N_7055,N_6981,N_6877);
xnor U7056 (N_7056,N_6938,N_6988);
and U7057 (N_7057,N_6979,N_6929);
nor U7058 (N_7058,N_6891,N_6956);
or U7059 (N_7059,N_6936,N_6924);
nand U7060 (N_7060,N_6914,N_6904);
xor U7061 (N_7061,N_6946,N_6900);
nand U7062 (N_7062,N_6940,N_6895);
nor U7063 (N_7063,N_6979,N_6878);
xor U7064 (N_7064,N_6924,N_6927);
or U7065 (N_7065,N_6892,N_6981);
or U7066 (N_7066,N_6991,N_6883);
and U7067 (N_7067,N_6926,N_6941);
nor U7068 (N_7068,N_6890,N_6930);
xnor U7069 (N_7069,N_6907,N_6885);
and U7070 (N_7070,N_6955,N_6946);
and U7071 (N_7071,N_6976,N_6986);
nand U7072 (N_7072,N_6975,N_6916);
nand U7073 (N_7073,N_6927,N_6941);
xnor U7074 (N_7074,N_6923,N_6886);
nor U7075 (N_7075,N_6953,N_6934);
xor U7076 (N_7076,N_6881,N_6995);
nor U7077 (N_7077,N_6986,N_6957);
xnor U7078 (N_7078,N_6960,N_6943);
and U7079 (N_7079,N_6954,N_6887);
and U7080 (N_7080,N_6956,N_6994);
and U7081 (N_7081,N_6926,N_6944);
or U7082 (N_7082,N_6884,N_6892);
or U7083 (N_7083,N_6997,N_6886);
nor U7084 (N_7084,N_6897,N_6954);
or U7085 (N_7085,N_6974,N_6928);
xnor U7086 (N_7086,N_6918,N_6881);
or U7087 (N_7087,N_6928,N_6955);
or U7088 (N_7088,N_6989,N_6913);
nand U7089 (N_7089,N_6992,N_6905);
xnor U7090 (N_7090,N_6904,N_6889);
and U7091 (N_7091,N_6920,N_6980);
or U7092 (N_7092,N_6951,N_6937);
xor U7093 (N_7093,N_6983,N_6886);
nand U7094 (N_7094,N_6899,N_6974);
nor U7095 (N_7095,N_6952,N_6968);
nand U7096 (N_7096,N_6955,N_6977);
xnor U7097 (N_7097,N_6937,N_6975);
nand U7098 (N_7098,N_6907,N_6912);
nor U7099 (N_7099,N_6917,N_6948);
nor U7100 (N_7100,N_6985,N_6887);
nor U7101 (N_7101,N_6933,N_6962);
xor U7102 (N_7102,N_6929,N_6884);
and U7103 (N_7103,N_6909,N_6910);
and U7104 (N_7104,N_6961,N_6964);
xor U7105 (N_7105,N_6897,N_6939);
nand U7106 (N_7106,N_6973,N_6985);
nand U7107 (N_7107,N_6908,N_6982);
nand U7108 (N_7108,N_6903,N_6914);
and U7109 (N_7109,N_6968,N_6888);
xnor U7110 (N_7110,N_6958,N_6892);
nand U7111 (N_7111,N_6890,N_6981);
nand U7112 (N_7112,N_6959,N_6913);
and U7113 (N_7113,N_6889,N_6893);
nor U7114 (N_7114,N_6951,N_6958);
or U7115 (N_7115,N_6910,N_6877);
and U7116 (N_7116,N_6964,N_6901);
xnor U7117 (N_7117,N_6975,N_6899);
nand U7118 (N_7118,N_6975,N_6958);
nand U7119 (N_7119,N_6909,N_6978);
xor U7120 (N_7120,N_6941,N_6939);
nor U7121 (N_7121,N_6924,N_6985);
nand U7122 (N_7122,N_6888,N_6934);
xnor U7123 (N_7123,N_6939,N_6896);
xor U7124 (N_7124,N_6971,N_6982);
nand U7125 (N_7125,N_7038,N_7037);
xnor U7126 (N_7126,N_7010,N_7060);
nand U7127 (N_7127,N_7016,N_7057);
nand U7128 (N_7128,N_7068,N_7006);
xor U7129 (N_7129,N_7073,N_7031);
and U7130 (N_7130,N_7112,N_7113);
and U7131 (N_7131,N_7081,N_7050);
nor U7132 (N_7132,N_7084,N_7028);
nor U7133 (N_7133,N_7047,N_7056);
and U7134 (N_7134,N_7085,N_7062);
and U7135 (N_7135,N_7042,N_7004);
nor U7136 (N_7136,N_7086,N_7049);
xor U7137 (N_7137,N_7080,N_7072);
or U7138 (N_7138,N_7021,N_7012);
nand U7139 (N_7139,N_7015,N_7108);
xnor U7140 (N_7140,N_7058,N_7033);
or U7141 (N_7141,N_7024,N_7071);
and U7142 (N_7142,N_7091,N_7089);
xnor U7143 (N_7143,N_7022,N_7019);
nand U7144 (N_7144,N_7097,N_7110);
nand U7145 (N_7145,N_7053,N_7116);
and U7146 (N_7146,N_7044,N_7120);
nand U7147 (N_7147,N_7040,N_7069);
or U7148 (N_7148,N_7011,N_7105);
nor U7149 (N_7149,N_7079,N_7075);
xor U7150 (N_7150,N_7003,N_7107);
and U7151 (N_7151,N_7046,N_7045);
and U7152 (N_7152,N_7013,N_7017);
xor U7153 (N_7153,N_7009,N_7102);
xor U7154 (N_7154,N_7088,N_7036);
and U7155 (N_7155,N_7121,N_7078);
xor U7156 (N_7156,N_7106,N_7065);
nor U7157 (N_7157,N_7109,N_7008);
xnor U7158 (N_7158,N_7117,N_7066);
nor U7159 (N_7159,N_7101,N_7077);
or U7160 (N_7160,N_7029,N_7026);
nor U7161 (N_7161,N_7055,N_7025);
nand U7162 (N_7162,N_7001,N_7054);
and U7163 (N_7163,N_7114,N_7104);
xor U7164 (N_7164,N_7076,N_7030);
nor U7165 (N_7165,N_7035,N_7043);
and U7166 (N_7166,N_7027,N_7041);
and U7167 (N_7167,N_7103,N_7018);
nand U7168 (N_7168,N_7119,N_7096);
xnor U7169 (N_7169,N_7020,N_7093);
or U7170 (N_7170,N_7034,N_7039);
and U7171 (N_7171,N_7002,N_7122);
xor U7172 (N_7172,N_7082,N_7074);
nand U7173 (N_7173,N_7095,N_7059);
xnor U7174 (N_7174,N_7111,N_7051);
xor U7175 (N_7175,N_7032,N_7052);
or U7176 (N_7176,N_7023,N_7123);
and U7177 (N_7177,N_7118,N_7090);
and U7178 (N_7178,N_7087,N_7063);
xor U7179 (N_7179,N_7098,N_7064);
nand U7180 (N_7180,N_7070,N_7061);
and U7181 (N_7181,N_7083,N_7005);
nand U7182 (N_7182,N_7124,N_7094);
nand U7183 (N_7183,N_7014,N_7067);
or U7184 (N_7184,N_7048,N_7115);
nand U7185 (N_7185,N_7007,N_7100);
and U7186 (N_7186,N_7092,N_7000);
xor U7187 (N_7187,N_7099,N_7032);
xnor U7188 (N_7188,N_7091,N_7057);
or U7189 (N_7189,N_7113,N_7117);
xnor U7190 (N_7190,N_7035,N_7070);
nand U7191 (N_7191,N_7017,N_7018);
or U7192 (N_7192,N_7087,N_7013);
and U7193 (N_7193,N_7048,N_7110);
and U7194 (N_7194,N_7021,N_7052);
or U7195 (N_7195,N_7119,N_7001);
or U7196 (N_7196,N_7010,N_7110);
xor U7197 (N_7197,N_7082,N_7031);
nor U7198 (N_7198,N_7047,N_7081);
nor U7199 (N_7199,N_7045,N_7080);
and U7200 (N_7200,N_7103,N_7043);
nor U7201 (N_7201,N_7113,N_7049);
xnor U7202 (N_7202,N_7117,N_7102);
nor U7203 (N_7203,N_7087,N_7096);
nand U7204 (N_7204,N_7075,N_7000);
or U7205 (N_7205,N_7109,N_7002);
or U7206 (N_7206,N_7024,N_7044);
xor U7207 (N_7207,N_7087,N_7061);
nand U7208 (N_7208,N_7121,N_7076);
or U7209 (N_7209,N_7092,N_7112);
nand U7210 (N_7210,N_7123,N_7017);
xnor U7211 (N_7211,N_7048,N_7020);
nand U7212 (N_7212,N_7007,N_7060);
nor U7213 (N_7213,N_7098,N_7074);
nand U7214 (N_7214,N_7042,N_7089);
or U7215 (N_7215,N_7018,N_7080);
or U7216 (N_7216,N_7099,N_7085);
or U7217 (N_7217,N_7019,N_7103);
or U7218 (N_7218,N_7110,N_7004);
and U7219 (N_7219,N_7117,N_7046);
xnor U7220 (N_7220,N_7034,N_7076);
and U7221 (N_7221,N_7041,N_7065);
xor U7222 (N_7222,N_7104,N_7043);
and U7223 (N_7223,N_7063,N_7096);
nor U7224 (N_7224,N_7073,N_7053);
xnor U7225 (N_7225,N_7021,N_7029);
nor U7226 (N_7226,N_7030,N_7052);
nand U7227 (N_7227,N_7064,N_7013);
or U7228 (N_7228,N_7111,N_7080);
or U7229 (N_7229,N_7106,N_7052);
xnor U7230 (N_7230,N_7075,N_7023);
or U7231 (N_7231,N_7004,N_7122);
nor U7232 (N_7232,N_7106,N_7016);
or U7233 (N_7233,N_7040,N_7063);
nor U7234 (N_7234,N_7001,N_7102);
or U7235 (N_7235,N_7117,N_7019);
xnor U7236 (N_7236,N_7018,N_7086);
nand U7237 (N_7237,N_7015,N_7010);
nand U7238 (N_7238,N_7005,N_7019);
nor U7239 (N_7239,N_7021,N_7058);
xor U7240 (N_7240,N_7047,N_7039);
and U7241 (N_7241,N_7050,N_7012);
and U7242 (N_7242,N_7017,N_7107);
and U7243 (N_7243,N_7084,N_7019);
or U7244 (N_7244,N_7118,N_7018);
or U7245 (N_7245,N_7025,N_7042);
xor U7246 (N_7246,N_7123,N_7046);
xor U7247 (N_7247,N_7115,N_7088);
or U7248 (N_7248,N_7113,N_7057);
xor U7249 (N_7249,N_7019,N_7029);
xnor U7250 (N_7250,N_7141,N_7204);
xor U7251 (N_7251,N_7228,N_7176);
nor U7252 (N_7252,N_7181,N_7174);
xor U7253 (N_7253,N_7206,N_7240);
xnor U7254 (N_7254,N_7218,N_7152);
nand U7255 (N_7255,N_7194,N_7248);
nor U7256 (N_7256,N_7199,N_7170);
nor U7257 (N_7257,N_7167,N_7197);
or U7258 (N_7258,N_7178,N_7144);
and U7259 (N_7259,N_7134,N_7183);
nand U7260 (N_7260,N_7177,N_7130);
and U7261 (N_7261,N_7207,N_7161);
nor U7262 (N_7262,N_7193,N_7237);
and U7263 (N_7263,N_7223,N_7227);
or U7264 (N_7264,N_7157,N_7160);
nor U7265 (N_7265,N_7241,N_7219);
or U7266 (N_7266,N_7151,N_7131);
or U7267 (N_7267,N_7192,N_7224);
nor U7268 (N_7268,N_7213,N_7215);
or U7269 (N_7269,N_7232,N_7225);
nor U7270 (N_7270,N_7165,N_7217);
xnor U7271 (N_7271,N_7236,N_7212);
xnor U7272 (N_7272,N_7139,N_7196);
xor U7273 (N_7273,N_7154,N_7186);
and U7274 (N_7274,N_7247,N_7226);
xor U7275 (N_7275,N_7138,N_7203);
nand U7276 (N_7276,N_7249,N_7171);
and U7277 (N_7277,N_7143,N_7132);
or U7278 (N_7278,N_7244,N_7235);
or U7279 (N_7279,N_7169,N_7209);
xnor U7280 (N_7280,N_7145,N_7173);
and U7281 (N_7281,N_7162,N_7128);
nand U7282 (N_7282,N_7190,N_7175);
or U7283 (N_7283,N_7188,N_7220);
nor U7284 (N_7284,N_7153,N_7168);
and U7285 (N_7285,N_7164,N_7148);
nor U7286 (N_7286,N_7172,N_7125);
and U7287 (N_7287,N_7191,N_7142);
nand U7288 (N_7288,N_7245,N_7229);
nor U7289 (N_7289,N_7208,N_7246);
nand U7290 (N_7290,N_7216,N_7201);
and U7291 (N_7291,N_7233,N_7195);
or U7292 (N_7292,N_7184,N_7211);
nor U7293 (N_7293,N_7182,N_7180);
or U7294 (N_7294,N_7185,N_7230);
or U7295 (N_7295,N_7214,N_7234);
and U7296 (N_7296,N_7243,N_7239);
and U7297 (N_7297,N_7156,N_7150);
and U7298 (N_7298,N_7189,N_7147);
and U7299 (N_7299,N_7136,N_7202);
nor U7300 (N_7300,N_7126,N_7198);
nor U7301 (N_7301,N_7166,N_7137);
nand U7302 (N_7302,N_7158,N_7155);
nand U7303 (N_7303,N_7242,N_7210);
nand U7304 (N_7304,N_7238,N_7231);
xnor U7305 (N_7305,N_7163,N_7127);
xor U7306 (N_7306,N_7179,N_7200);
or U7307 (N_7307,N_7140,N_7205);
and U7308 (N_7308,N_7221,N_7222);
or U7309 (N_7309,N_7149,N_7146);
nand U7310 (N_7310,N_7159,N_7187);
xnor U7311 (N_7311,N_7133,N_7129);
nand U7312 (N_7312,N_7135,N_7246);
or U7313 (N_7313,N_7230,N_7237);
xor U7314 (N_7314,N_7223,N_7142);
nor U7315 (N_7315,N_7242,N_7197);
and U7316 (N_7316,N_7233,N_7140);
and U7317 (N_7317,N_7141,N_7129);
or U7318 (N_7318,N_7152,N_7235);
xnor U7319 (N_7319,N_7205,N_7235);
or U7320 (N_7320,N_7144,N_7162);
xor U7321 (N_7321,N_7129,N_7215);
or U7322 (N_7322,N_7137,N_7225);
nand U7323 (N_7323,N_7216,N_7247);
xor U7324 (N_7324,N_7195,N_7177);
and U7325 (N_7325,N_7232,N_7134);
xnor U7326 (N_7326,N_7217,N_7223);
xnor U7327 (N_7327,N_7183,N_7153);
nand U7328 (N_7328,N_7215,N_7212);
or U7329 (N_7329,N_7223,N_7211);
and U7330 (N_7330,N_7145,N_7166);
nor U7331 (N_7331,N_7238,N_7130);
nand U7332 (N_7332,N_7162,N_7218);
nand U7333 (N_7333,N_7201,N_7191);
xnor U7334 (N_7334,N_7166,N_7146);
xnor U7335 (N_7335,N_7198,N_7245);
xnor U7336 (N_7336,N_7155,N_7219);
nor U7337 (N_7337,N_7195,N_7157);
xnor U7338 (N_7338,N_7224,N_7174);
xnor U7339 (N_7339,N_7156,N_7212);
nand U7340 (N_7340,N_7205,N_7139);
or U7341 (N_7341,N_7214,N_7216);
or U7342 (N_7342,N_7136,N_7201);
or U7343 (N_7343,N_7157,N_7205);
nor U7344 (N_7344,N_7244,N_7223);
or U7345 (N_7345,N_7190,N_7230);
or U7346 (N_7346,N_7249,N_7130);
nand U7347 (N_7347,N_7242,N_7125);
nand U7348 (N_7348,N_7192,N_7235);
xnor U7349 (N_7349,N_7166,N_7159);
nand U7350 (N_7350,N_7245,N_7222);
or U7351 (N_7351,N_7233,N_7231);
xnor U7352 (N_7352,N_7130,N_7141);
nor U7353 (N_7353,N_7236,N_7165);
or U7354 (N_7354,N_7226,N_7154);
nor U7355 (N_7355,N_7194,N_7148);
and U7356 (N_7356,N_7207,N_7249);
or U7357 (N_7357,N_7155,N_7237);
nor U7358 (N_7358,N_7137,N_7249);
and U7359 (N_7359,N_7239,N_7248);
nor U7360 (N_7360,N_7239,N_7207);
xnor U7361 (N_7361,N_7151,N_7210);
xor U7362 (N_7362,N_7147,N_7149);
nor U7363 (N_7363,N_7127,N_7156);
nand U7364 (N_7364,N_7248,N_7131);
and U7365 (N_7365,N_7243,N_7186);
xor U7366 (N_7366,N_7138,N_7201);
nor U7367 (N_7367,N_7126,N_7167);
or U7368 (N_7368,N_7208,N_7145);
nand U7369 (N_7369,N_7128,N_7163);
and U7370 (N_7370,N_7196,N_7193);
or U7371 (N_7371,N_7229,N_7143);
nand U7372 (N_7372,N_7187,N_7173);
nor U7373 (N_7373,N_7249,N_7146);
nand U7374 (N_7374,N_7235,N_7177);
xor U7375 (N_7375,N_7356,N_7360);
nand U7376 (N_7376,N_7336,N_7273);
or U7377 (N_7377,N_7309,N_7329);
or U7378 (N_7378,N_7283,N_7328);
or U7379 (N_7379,N_7359,N_7349);
xor U7380 (N_7380,N_7268,N_7345);
and U7381 (N_7381,N_7352,N_7295);
or U7382 (N_7382,N_7290,N_7306);
and U7383 (N_7383,N_7331,N_7260);
xnor U7384 (N_7384,N_7281,N_7319);
xor U7385 (N_7385,N_7250,N_7298);
nand U7386 (N_7386,N_7316,N_7327);
nand U7387 (N_7387,N_7252,N_7311);
and U7388 (N_7388,N_7255,N_7366);
nor U7389 (N_7389,N_7263,N_7261);
xnor U7390 (N_7390,N_7272,N_7288);
or U7391 (N_7391,N_7346,N_7320);
nor U7392 (N_7392,N_7322,N_7372);
nand U7393 (N_7393,N_7278,N_7284);
nor U7394 (N_7394,N_7315,N_7370);
and U7395 (N_7395,N_7299,N_7353);
and U7396 (N_7396,N_7307,N_7304);
or U7397 (N_7397,N_7364,N_7369);
nand U7398 (N_7398,N_7340,N_7318);
nor U7399 (N_7399,N_7254,N_7310);
xor U7400 (N_7400,N_7287,N_7348);
or U7401 (N_7401,N_7279,N_7267);
xnor U7402 (N_7402,N_7317,N_7374);
nor U7403 (N_7403,N_7256,N_7285);
and U7404 (N_7404,N_7341,N_7308);
nor U7405 (N_7405,N_7297,N_7368);
nand U7406 (N_7406,N_7286,N_7305);
nand U7407 (N_7407,N_7266,N_7262);
or U7408 (N_7408,N_7354,N_7313);
and U7409 (N_7409,N_7338,N_7342);
xor U7410 (N_7410,N_7253,N_7296);
or U7411 (N_7411,N_7339,N_7258);
and U7412 (N_7412,N_7357,N_7294);
nor U7413 (N_7413,N_7257,N_7332);
or U7414 (N_7414,N_7355,N_7303);
nor U7415 (N_7415,N_7302,N_7276);
nor U7416 (N_7416,N_7314,N_7365);
and U7417 (N_7417,N_7343,N_7274);
xnor U7418 (N_7418,N_7337,N_7367);
or U7419 (N_7419,N_7259,N_7289);
or U7420 (N_7420,N_7269,N_7334);
or U7421 (N_7421,N_7280,N_7330);
nor U7422 (N_7422,N_7251,N_7333);
xor U7423 (N_7423,N_7265,N_7291);
and U7424 (N_7424,N_7293,N_7358);
or U7425 (N_7425,N_7350,N_7321);
nor U7426 (N_7426,N_7264,N_7312);
or U7427 (N_7427,N_7271,N_7275);
nand U7428 (N_7428,N_7371,N_7300);
xor U7429 (N_7429,N_7344,N_7301);
nor U7430 (N_7430,N_7347,N_7270);
and U7431 (N_7431,N_7361,N_7363);
and U7432 (N_7432,N_7362,N_7282);
or U7433 (N_7433,N_7324,N_7292);
or U7434 (N_7434,N_7373,N_7351);
xor U7435 (N_7435,N_7326,N_7323);
nand U7436 (N_7436,N_7277,N_7335);
xor U7437 (N_7437,N_7325,N_7307);
and U7438 (N_7438,N_7308,N_7364);
or U7439 (N_7439,N_7272,N_7261);
and U7440 (N_7440,N_7320,N_7344);
or U7441 (N_7441,N_7263,N_7278);
nand U7442 (N_7442,N_7310,N_7261);
xnor U7443 (N_7443,N_7292,N_7326);
nand U7444 (N_7444,N_7318,N_7277);
or U7445 (N_7445,N_7364,N_7261);
xor U7446 (N_7446,N_7274,N_7299);
nor U7447 (N_7447,N_7267,N_7343);
and U7448 (N_7448,N_7257,N_7303);
nand U7449 (N_7449,N_7362,N_7300);
and U7450 (N_7450,N_7373,N_7288);
or U7451 (N_7451,N_7274,N_7268);
or U7452 (N_7452,N_7275,N_7278);
nand U7453 (N_7453,N_7278,N_7252);
nand U7454 (N_7454,N_7272,N_7279);
xnor U7455 (N_7455,N_7329,N_7367);
or U7456 (N_7456,N_7251,N_7301);
nand U7457 (N_7457,N_7367,N_7291);
nor U7458 (N_7458,N_7340,N_7281);
or U7459 (N_7459,N_7254,N_7359);
nor U7460 (N_7460,N_7288,N_7339);
or U7461 (N_7461,N_7298,N_7357);
xnor U7462 (N_7462,N_7308,N_7374);
xor U7463 (N_7463,N_7358,N_7320);
nand U7464 (N_7464,N_7290,N_7348);
or U7465 (N_7465,N_7268,N_7326);
xor U7466 (N_7466,N_7314,N_7319);
xor U7467 (N_7467,N_7279,N_7297);
xnor U7468 (N_7468,N_7310,N_7292);
nor U7469 (N_7469,N_7353,N_7251);
xor U7470 (N_7470,N_7363,N_7321);
and U7471 (N_7471,N_7256,N_7260);
xor U7472 (N_7472,N_7317,N_7262);
xnor U7473 (N_7473,N_7282,N_7332);
and U7474 (N_7474,N_7339,N_7264);
nor U7475 (N_7475,N_7268,N_7329);
and U7476 (N_7476,N_7322,N_7269);
nor U7477 (N_7477,N_7255,N_7353);
nor U7478 (N_7478,N_7317,N_7266);
nor U7479 (N_7479,N_7314,N_7262);
or U7480 (N_7480,N_7285,N_7353);
or U7481 (N_7481,N_7250,N_7299);
xor U7482 (N_7482,N_7355,N_7268);
xor U7483 (N_7483,N_7336,N_7339);
nor U7484 (N_7484,N_7283,N_7251);
nor U7485 (N_7485,N_7256,N_7371);
xnor U7486 (N_7486,N_7268,N_7347);
and U7487 (N_7487,N_7270,N_7294);
and U7488 (N_7488,N_7359,N_7256);
nor U7489 (N_7489,N_7260,N_7354);
nor U7490 (N_7490,N_7301,N_7259);
nand U7491 (N_7491,N_7263,N_7273);
or U7492 (N_7492,N_7316,N_7265);
nor U7493 (N_7493,N_7346,N_7286);
xnor U7494 (N_7494,N_7374,N_7292);
xor U7495 (N_7495,N_7289,N_7342);
and U7496 (N_7496,N_7363,N_7314);
nor U7497 (N_7497,N_7373,N_7279);
or U7498 (N_7498,N_7264,N_7292);
nand U7499 (N_7499,N_7331,N_7277);
or U7500 (N_7500,N_7482,N_7481);
and U7501 (N_7501,N_7497,N_7394);
or U7502 (N_7502,N_7456,N_7432);
xor U7503 (N_7503,N_7443,N_7467);
and U7504 (N_7504,N_7423,N_7480);
nor U7505 (N_7505,N_7403,N_7389);
or U7506 (N_7506,N_7445,N_7421);
or U7507 (N_7507,N_7473,N_7395);
or U7508 (N_7508,N_7495,N_7387);
nand U7509 (N_7509,N_7486,N_7458);
nor U7510 (N_7510,N_7477,N_7379);
xnor U7511 (N_7511,N_7378,N_7487);
nand U7512 (N_7512,N_7459,N_7439);
or U7513 (N_7513,N_7424,N_7400);
xor U7514 (N_7514,N_7382,N_7411);
xor U7515 (N_7515,N_7413,N_7406);
nor U7516 (N_7516,N_7402,N_7409);
nand U7517 (N_7517,N_7476,N_7404);
xnor U7518 (N_7518,N_7390,N_7418);
nand U7519 (N_7519,N_7429,N_7401);
and U7520 (N_7520,N_7433,N_7491);
xnor U7521 (N_7521,N_7492,N_7484);
and U7522 (N_7522,N_7427,N_7489);
nand U7523 (N_7523,N_7410,N_7447);
and U7524 (N_7524,N_7399,N_7455);
or U7525 (N_7525,N_7498,N_7430);
nor U7526 (N_7526,N_7470,N_7425);
and U7527 (N_7527,N_7460,N_7438);
nand U7528 (N_7528,N_7380,N_7466);
xnor U7529 (N_7529,N_7483,N_7414);
nand U7530 (N_7530,N_7468,N_7471);
nand U7531 (N_7531,N_7457,N_7416);
xnor U7532 (N_7532,N_7478,N_7397);
and U7533 (N_7533,N_7435,N_7449);
or U7534 (N_7534,N_7442,N_7388);
or U7535 (N_7535,N_7448,N_7381);
and U7536 (N_7536,N_7415,N_7431);
and U7537 (N_7537,N_7384,N_7446);
or U7538 (N_7538,N_7426,N_7499);
nand U7539 (N_7539,N_7496,N_7469);
nand U7540 (N_7540,N_7419,N_7392);
and U7541 (N_7541,N_7391,N_7398);
nor U7542 (N_7542,N_7422,N_7420);
nand U7543 (N_7543,N_7494,N_7472);
and U7544 (N_7544,N_7461,N_7463);
xor U7545 (N_7545,N_7464,N_7462);
nand U7546 (N_7546,N_7451,N_7490);
nand U7547 (N_7547,N_7493,N_7393);
xnor U7548 (N_7548,N_7396,N_7386);
nand U7549 (N_7549,N_7377,N_7385);
nor U7550 (N_7550,N_7383,N_7485);
nor U7551 (N_7551,N_7454,N_7375);
nand U7552 (N_7552,N_7428,N_7405);
and U7553 (N_7553,N_7407,N_7452);
and U7554 (N_7554,N_7436,N_7441);
or U7555 (N_7555,N_7474,N_7475);
nor U7556 (N_7556,N_7450,N_7465);
nor U7557 (N_7557,N_7376,N_7434);
nor U7558 (N_7558,N_7488,N_7412);
nor U7559 (N_7559,N_7417,N_7440);
nand U7560 (N_7560,N_7408,N_7479);
nor U7561 (N_7561,N_7444,N_7453);
or U7562 (N_7562,N_7437,N_7443);
and U7563 (N_7563,N_7396,N_7449);
nor U7564 (N_7564,N_7450,N_7402);
nand U7565 (N_7565,N_7382,N_7424);
or U7566 (N_7566,N_7453,N_7452);
and U7567 (N_7567,N_7433,N_7376);
xnor U7568 (N_7568,N_7448,N_7414);
nor U7569 (N_7569,N_7455,N_7415);
and U7570 (N_7570,N_7394,N_7413);
or U7571 (N_7571,N_7417,N_7495);
and U7572 (N_7572,N_7440,N_7375);
or U7573 (N_7573,N_7410,N_7450);
and U7574 (N_7574,N_7458,N_7427);
or U7575 (N_7575,N_7417,N_7479);
nand U7576 (N_7576,N_7451,N_7432);
nand U7577 (N_7577,N_7380,N_7472);
nand U7578 (N_7578,N_7440,N_7458);
and U7579 (N_7579,N_7450,N_7429);
and U7580 (N_7580,N_7472,N_7434);
or U7581 (N_7581,N_7450,N_7400);
and U7582 (N_7582,N_7479,N_7468);
or U7583 (N_7583,N_7441,N_7437);
nand U7584 (N_7584,N_7459,N_7478);
and U7585 (N_7585,N_7459,N_7421);
xor U7586 (N_7586,N_7474,N_7450);
xor U7587 (N_7587,N_7463,N_7466);
nor U7588 (N_7588,N_7408,N_7433);
nor U7589 (N_7589,N_7471,N_7480);
and U7590 (N_7590,N_7497,N_7485);
nor U7591 (N_7591,N_7431,N_7429);
or U7592 (N_7592,N_7484,N_7468);
xnor U7593 (N_7593,N_7452,N_7462);
xnor U7594 (N_7594,N_7476,N_7481);
nor U7595 (N_7595,N_7421,N_7384);
nor U7596 (N_7596,N_7466,N_7375);
and U7597 (N_7597,N_7450,N_7395);
and U7598 (N_7598,N_7395,N_7482);
or U7599 (N_7599,N_7456,N_7487);
and U7600 (N_7600,N_7384,N_7423);
nor U7601 (N_7601,N_7432,N_7497);
nor U7602 (N_7602,N_7473,N_7499);
and U7603 (N_7603,N_7399,N_7432);
nor U7604 (N_7604,N_7411,N_7467);
and U7605 (N_7605,N_7451,N_7475);
or U7606 (N_7606,N_7409,N_7398);
xnor U7607 (N_7607,N_7471,N_7383);
or U7608 (N_7608,N_7492,N_7430);
and U7609 (N_7609,N_7400,N_7379);
nand U7610 (N_7610,N_7476,N_7375);
nand U7611 (N_7611,N_7475,N_7400);
xnor U7612 (N_7612,N_7451,N_7422);
nand U7613 (N_7613,N_7424,N_7478);
and U7614 (N_7614,N_7447,N_7405);
nand U7615 (N_7615,N_7407,N_7465);
xnor U7616 (N_7616,N_7419,N_7389);
nor U7617 (N_7617,N_7386,N_7414);
or U7618 (N_7618,N_7406,N_7382);
and U7619 (N_7619,N_7398,N_7458);
nand U7620 (N_7620,N_7432,N_7480);
nor U7621 (N_7621,N_7475,N_7407);
or U7622 (N_7622,N_7433,N_7481);
or U7623 (N_7623,N_7407,N_7466);
or U7624 (N_7624,N_7415,N_7418);
nor U7625 (N_7625,N_7583,N_7517);
nand U7626 (N_7626,N_7600,N_7504);
nor U7627 (N_7627,N_7606,N_7524);
nor U7628 (N_7628,N_7577,N_7533);
and U7629 (N_7629,N_7623,N_7554);
or U7630 (N_7630,N_7591,N_7539);
xor U7631 (N_7631,N_7500,N_7519);
nor U7632 (N_7632,N_7563,N_7514);
nor U7633 (N_7633,N_7515,N_7509);
nor U7634 (N_7634,N_7586,N_7607);
nor U7635 (N_7635,N_7560,N_7604);
and U7636 (N_7636,N_7528,N_7530);
nand U7637 (N_7637,N_7540,N_7572);
or U7638 (N_7638,N_7603,N_7574);
xnor U7639 (N_7639,N_7547,N_7502);
and U7640 (N_7640,N_7520,N_7552);
nor U7641 (N_7641,N_7585,N_7587);
nand U7642 (N_7642,N_7521,N_7523);
nand U7643 (N_7643,N_7513,N_7570);
nor U7644 (N_7644,N_7595,N_7543);
nor U7645 (N_7645,N_7546,N_7569);
xnor U7646 (N_7646,N_7526,N_7592);
nand U7647 (N_7647,N_7567,N_7617);
nand U7648 (N_7648,N_7542,N_7541);
or U7649 (N_7649,N_7624,N_7532);
and U7650 (N_7650,N_7580,N_7564);
and U7651 (N_7651,N_7609,N_7549);
or U7652 (N_7652,N_7551,N_7538);
xor U7653 (N_7653,N_7518,N_7615);
nand U7654 (N_7654,N_7568,N_7608);
and U7655 (N_7655,N_7503,N_7616);
nor U7656 (N_7656,N_7566,N_7550);
nor U7657 (N_7657,N_7605,N_7620);
xor U7658 (N_7658,N_7511,N_7584);
nor U7659 (N_7659,N_7597,N_7562);
and U7660 (N_7660,N_7601,N_7555);
xor U7661 (N_7661,N_7536,N_7505);
xor U7662 (N_7662,N_7622,N_7588);
nor U7663 (N_7663,N_7565,N_7548);
xor U7664 (N_7664,N_7578,N_7561);
xnor U7665 (N_7665,N_7612,N_7618);
nand U7666 (N_7666,N_7573,N_7596);
xor U7667 (N_7667,N_7557,N_7507);
xor U7668 (N_7668,N_7534,N_7556);
nand U7669 (N_7669,N_7611,N_7510);
nor U7670 (N_7670,N_7582,N_7613);
xor U7671 (N_7671,N_7619,N_7590);
nand U7672 (N_7672,N_7558,N_7501);
nand U7673 (N_7673,N_7522,N_7599);
nand U7674 (N_7674,N_7544,N_7506);
nand U7675 (N_7675,N_7598,N_7594);
and U7676 (N_7676,N_7575,N_7525);
or U7677 (N_7677,N_7512,N_7602);
or U7678 (N_7678,N_7571,N_7610);
or U7679 (N_7679,N_7527,N_7508);
nor U7680 (N_7680,N_7516,N_7576);
nor U7681 (N_7681,N_7621,N_7553);
and U7682 (N_7682,N_7535,N_7531);
or U7683 (N_7683,N_7559,N_7614);
nor U7684 (N_7684,N_7579,N_7545);
nand U7685 (N_7685,N_7529,N_7593);
and U7686 (N_7686,N_7581,N_7537);
nor U7687 (N_7687,N_7589,N_7599);
and U7688 (N_7688,N_7503,N_7589);
nand U7689 (N_7689,N_7551,N_7557);
xor U7690 (N_7690,N_7578,N_7595);
nand U7691 (N_7691,N_7608,N_7523);
or U7692 (N_7692,N_7509,N_7593);
nor U7693 (N_7693,N_7620,N_7621);
nand U7694 (N_7694,N_7586,N_7513);
nand U7695 (N_7695,N_7603,N_7596);
and U7696 (N_7696,N_7553,N_7525);
or U7697 (N_7697,N_7505,N_7551);
nor U7698 (N_7698,N_7508,N_7554);
and U7699 (N_7699,N_7515,N_7556);
nand U7700 (N_7700,N_7617,N_7616);
xor U7701 (N_7701,N_7536,N_7568);
nand U7702 (N_7702,N_7516,N_7529);
xor U7703 (N_7703,N_7507,N_7508);
nor U7704 (N_7704,N_7539,N_7513);
and U7705 (N_7705,N_7618,N_7611);
nor U7706 (N_7706,N_7606,N_7564);
nor U7707 (N_7707,N_7616,N_7571);
and U7708 (N_7708,N_7579,N_7622);
and U7709 (N_7709,N_7571,N_7536);
or U7710 (N_7710,N_7517,N_7540);
nor U7711 (N_7711,N_7596,N_7598);
nor U7712 (N_7712,N_7565,N_7528);
nor U7713 (N_7713,N_7540,N_7604);
xor U7714 (N_7714,N_7622,N_7586);
nand U7715 (N_7715,N_7580,N_7539);
and U7716 (N_7716,N_7569,N_7509);
nand U7717 (N_7717,N_7556,N_7604);
nor U7718 (N_7718,N_7528,N_7600);
xnor U7719 (N_7719,N_7560,N_7566);
and U7720 (N_7720,N_7566,N_7503);
xnor U7721 (N_7721,N_7509,N_7506);
nor U7722 (N_7722,N_7582,N_7522);
or U7723 (N_7723,N_7589,N_7583);
or U7724 (N_7724,N_7566,N_7534);
and U7725 (N_7725,N_7576,N_7504);
nor U7726 (N_7726,N_7567,N_7574);
and U7727 (N_7727,N_7564,N_7618);
nor U7728 (N_7728,N_7532,N_7520);
and U7729 (N_7729,N_7550,N_7549);
xor U7730 (N_7730,N_7546,N_7578);
or U7731 (N_7731,N_7619,N_7617);
nor U7732 (N_7732,N_7560,N_7556);
nor U7733 (N_7733,N_7517,N_7619);
nand U7734 (N_7734,N_7551,N_7515);
xor U7735 (N_7735,N_7528,N_7620);
and U7736 (N_7736,N_7540,N_7533);
or U7737 (N_7737,N_7554,N_7615);
and U7738 (N_7738,N_7520,N_7554);
or U7739 (N_7739,N_7515,N_7609);
xnor U7740 (N_7740,N_7587,N_7568);
xnor U7741 (N_7741,N_7546,N_7577);
nand U7742 (N_7742,N_7566,N_7616);
nand U7743 (N_7743,N_7557,N_7541);
and U7744 (N_7744,N_7615,N_7571);
xnor U7745 (N_7745,N_7538,N_7565);
xnor U7746 (N_7746,N_7503,N_7567);
or U7747 (N_7747,N_7589,N_7615);
nand U7748 (N_7748,N_7582,N_7501);
or U7749 (N_7749,N_7513,N_7507);
nor U7750 (N_7750,N_7640,N_7726);
nand U7751 (N_7751,N_7628,N_7699);
nand U7752 (N_7752,N_7703,N_7720);
and U7753 (N_7753,N_7716,N_7649);
nand U7754 (N_7754,N_7634,N_7718);
nor U7755 (N_7755,N_7639,N_7712);
nor U7756 (N_7756,N_7719,N_7741);
nand U7757 (N_7757,N_7705,N_7733);
nor U7758 (N_7758,N_7644,N_7710);
nor U7759 (N_7759,N_7652,N_7681);
xor U7760 (N_7760,N_7687,N_7698);
nand U7761 (N_7761,N_7743,N_7650);
or U7762 (N_7762,N_7737,N_7749);
nand U7763 (N_7763,N_7675,N_7663);
xor U7764 (N_7764,N_7701,N_7682);
nand U7765 (N_7765,N_7633,N_7664);
and U7766 (N_7766,N_7666,N_7691);
nand U7767 (N_7767,N_7642,N_7748);
and U7768 (N_7768,N_7693,N_7714);
nand U7769 (N_7769,N_7648,N_7683);
xnor U7770 (N_7770,N_7643,N_7665);
and U7771 (N_7771,N_7724,N_7653);
nand U7772 (N_7772,N_7686,N_7632);
or U7773 (N_7773,N_7713,N_7630);
nor U7774 (N_7774,N_7722,N_7636);
nand U7775 (N_7775,N_7685,N_7669);
nor U7776 (N_7776,N_7629,N_7674);
xnor U7777 (N_7777,N_7702,N_7739);
or U7778 (N_7778,N_7747,N_7684);
xnor U7779 (N_7779,N_7677,N_7635);
nand U7780 (N_7780,N_7709,N_7732);
xor U7781 (N_7781,N_7658,N_7730);
xnor U7782 (N_7782,N_7727,N_7697);
nand U7783 (N_7783,N_7692,N_7647);
nand U7784 (N_7784,N_7657,N_7641);
or U7785 (N_7785,N_7723,N_7667);
or U7786 (N_7786,N_7696,N_7626);
or U7787 (N_7787,N_7725,N_7660);
xor U7788 (N_7788,N_7740,N_7731);
nand U7789 (N_7789,N_7625,N_7707);
nand U7790 (N_7790,N_7738,N_7715);
nand U7791 (N_7791,N_7728,N_7711);
xor U7792 (N_7792,N_7678,N_7736);
nor U7793 (N_7793,N_7637,N_7679);
nand U7794 (N_7794,N_7729,N_7721);
and U7795 (N_7795,N_7704,N_7655);
and U7796 (N_7796,N_7646,N_7638);
nand U7797 (N_7797,N_7744,N_7746);
or U7798 (N_7798,N_7695,N_7645);
or U7799 (N_7799,N_7706,N_7688);
nor U7800 (N_7800,N_7654,N_7670);
xnor U7801 (N_7801,N_7689,N_7694);
and U7802 (N_7802,N_7700,N_7656);
nand U7803 (N_7803,N_7631,N_7734);
nor U7804 (N_7804,N_7690,N_7672);
and U7805 (N_7805,N_7708,N_7745);
nand U7806 (N_7806,N_7742,N_7668);
nor U7807 (N_7807,N_7676,N_7662);
or U7808 (N_7808,N_7680,N_7735);
nor U7809 (N_7809,N_7627,N_7651);
xnor U7810 (N_7810,N_7673,N_7659);
and U7811 (N_7811,N_7661,N_7671);
xnor U7812 (N_7812,N_7717,N_7729);
and U7813 (N_7813,N_7716,N_7675);
nand U7814 (N_7814,N_7633,N_7745);
nand U7815 (N_7815,N_7700,N_7738);
and U7816 (N_7816,N_7728,N_7681);
and U7817 (N_7817,N_7679,N_7693);
and U7818 (N_7818,N_7635,N_7643);
xnor U7819 (N_7819,N_7627,N_7634);
nand U7820 (N_7820,N_7675,N_7729);
xor U7821 (N_7821,N_7726,N_7672);
nor U7822 (N_7822,N_7647,N_7739);
nor U7823 (N_7823,N_7659,N_7690);
nor U7824 (N_7824,N_7714,N_7712);
and U7825 (N_7825,N_7627,N_7643);
xnor U7826 (N_7826,N_7650,N_7693);
xor U7827 (N_7827,N_7635,N_7658);
xnor U7828 (N_7828,N_7674,N_7669);
and U7829 (N_7829,N_7678,N_7648);
nor U7830 (N_7830,N_7646,N_7744);
xor U7831 (N_7831,N_7741,N_7657);
xnor U7832 (N_7832,N_7686,N_7672);
nand U7833 (N_7833,N_7701,N_7726);
and U7834 (N_7834,N_7676,N_7731);
nor U7835 (N_7835,N_7714,N_7690);
and U7836 (N_7836,N_7705,N_7642);
and U7837 (N_7837,N_7709,N_7660);
nor U7838 (N_7838,N_7697,N_7746);
xnor U7839 (N_7839,N_7639,N_7685);
and U7840 (N_7840,N_7653,N_7634);
nand U7841 (N_7841,N_7746,N_7674);
or U7842 (N_7842,N_7686,N_7699);
nand U7843 (N_7843,N_7662,N_7670);
or U7844 (N_7844,N_7647,N_7720);
nand U7845 (N_7845,N_7699,N_7748);
nand U7846 (N_7846,N_7690,N_7745);
xnor U7847 (N_7847,N_7648,N_7731);
nand U7848 (N_7848,N_7627,N_7745);
and U7849 (N_7849,N_7627,N_7654);
nor U7850 (N_7850,N_7735,N_7631);
or U7851 (N_7851,N_7684,N_7680);
or U7852 (N_7852,N_7708,N_7684);
nor U7853 (N_7853,N_7705,N_7696);
or U7854 (N_7854,N_7713,N_7652);
nor U7855 (N_7855,N_7739,N_7707);
xor U7856 (N_7856,N_7669,N_7706);
nand U7857 (N_7857,N_7706,N_7649);
nand U7858 (N_7858,N_7669,N_7724);
nand U7859 (N_7859,N_7674,N_7722);
and U7860 (N_7860,N_7695,N_7703);
nand U7861 (N_7861,N_7632,N_7626);
xor U7862 (N_7862,N_7749,N_7673);
nand U7863 (N_7863,N_7708,N_7669);
nand U7864 (N_7864,N_7634,N_7658);
or U7865 (N_7865,N_7653,N_7704);
xnor U7866 (N_7866,N_7676,N_7637);
and U7867 (N_7867,N_7746,N_7722);
nand U7868 (N_7868,N_7744,N_7695);
xor U7869 (N_7869,N_7644,N_7719);
nor U7870 (N_7870,N_7670,N_7682);
nor U7871 (N_7871,N_7717,N_7689);
or U7872 (N_7872,N_7669,N_7705);
or U7873 (N_7873,N_7674,N_7648);
and U7874 (N_7874,N_7709,N_7740);
and U7875 (N_7875,N_7831,N_7849);
and U7876 (N_7876,N_7838,N_7834);
nand U7877 (N_7877,N_7858,N_7765);
nor U7878 (N_7878,N_7756,N_7859);
or U7879 (N_7879,N_7827,N_7782);
or U7880 (N_7880,N_7791,N_7781);
xor U7881 (N_7881,N_7794,N_7857);
or U7882 (N_7882,N_7853,N_7776);
and U7883 (N_7883,N_7800,N_7790);
nand U7884 (N_7884,N_7759,N_7854);
nor U7885 (N_7885,N_7763,N_7753);
nor U7886 (N_7886,N_7837,N_7848);
or U7887 (N_7887,N_7841,N_7811);
and U7888 (N_7888,N_7844,N_7860);
and U7889 (N_7889,N_7816,N_7750);
nand U7890 (N_7890,N_7795,N_7845);
nor U7891 (N_7891,N_7784,N_7803);
xor U7892 (N_7892,N_7863,N_7812);
xor U7893 (N_7893,N_7761,N_7852);
nor U7894 (N_7894,N_7783,N_7815);
xor U7895 (N_7895,N_7768,N_7775);
and U7896 (N_7896,N_7767,N_7817);
nor U7897 (N_7897,N_7808,N_7819);
nand U7898 (N_7898,N_7823,N_7826);
nand U7899 (N_7899,N_7786,N_7758);
or U7900 (N_7900,N_7787,N_7867);
and U7901 (N_7901,N_7870,N_7829);
nand U7902 (N_7902,N_7799,N_7805);
or U7903 (N_7903,N_7825,N_7842);
nor U7904 (N_7904,N_7861,N_7828);
nor U7905 (N_7905,N_7809,N_7872);
xor U7906 (N_7906,N_7788,N_7874);
xor U7907 (N_7907,N_7824,N_7843);
nor U7908 (N_7908,N_7754,N_7850);
and U7909 (N_7909,N_7865,N_7773);
nand U7910 (N_7910,N_7832,N_7777);
or U7911 (N_7911,N_7810,N_7833);
or U7912 (N_7912,N_7801,N_7769);
and U7913 (N_7913,N_7873,N_7752);
nor U7914 (N_7914,N_7855,N_7846);
xnor U7915 (N_7915,N_7864,N_7770);
nand U7916 (N_7916,N_7806,N_7796);
nand U7917 (N_7917,N_7851,N_7751);
or U7918 (N_7918,N_7868,N_7820);
nor U7919 (N_7919,N_7762,N_7755);
and U7920 (N_7920,N_7785,N_7798);
xor U7921 (N_7921,N_7771,N_7847);
nor U7922 (N_7922,N_7866,N_7839);
or U7923 (N_7923,N_7778,N_7789);
nand U7924 (N_7924,N_7779,N_7807);
xor U7925 (N_7925,N_7797,N_7764);
nand U7926 (N_7926,N_7835,N_7836);
or U7927 (N_7927,N_7766,N_7774);
and U7928 (N_7928,N_7757,N_7821);
or U7929 (N_7929,N_7856,N_7780);
and U7930 (N_7930,N_7760,N_7830);
or U7931 (N_7931,N_7862,N_7814);
nand U7932 (N_7932,N_7840,N_7804);
or U7933 (N_7933,N_7772,N_7813);
nor U7934 (N_7934,N_7802,N_7869);
nor U7935 (N_7935,N_7871,N_7818);
nand U7936 (N_7936,N_7822,N_7792);
xor U7937 (N_7937,N_7793,N_7786);
nor U7938 (N_7938,N_7814,N_7807);
xnor U7939 (N_7939,N_7789,N_7867);
and U7940 (N_7940,N_7755,N_7754);
and U7941 (N_7941,N_7811,N_7868);
nand U7942 (N_7942,N_7840,N_7761);
and U7943 (N_7943,N_7870,N_7783);
nor U7944 (N_7944,N_7761,N_7789);
xor U7945 (N_7945,N_7842,N_7793);
or U7946 (N_7946,N_7815,N_7854);
xnor U7947 (N_7947,N_7870,N_7859);
nand U7948 (N_7948,N_7811,N_7784);
or U7949 (N_7949,N_7781,N_7768);
and U7950 (N_7950,N_7865,N_7756);
nor U7951 (N_7951,N_7781,N_7844);
nor U7952 (N_7952,N_7792,N_7805);
xnor U7953 (N_7953,N_7847,N_7798);
or U7954 (N_7954,N_7862,N_7770);
nor U7955 (N_7955,N_7811,N_7805);
or U7956 (N_7956,N_7871,N_7840);
nor U7957 (N_7957,N_7795,N_7777);
or U7958 (N_7958,N_7777,N_7818);
nor U7959 (N_7959,N_7872,N_7794);
and U7960 (N_7960,N_7785,N_7799);
and U7961 (N_7961,N_7773,N_7757);
xor U7962 (N_7962,N_7815,N_7850);
nand U7963 (N_7963,N_7869,N_7782);
xor U7964 (N_7964,N_7858,N_7855);
or U7965 (N_7965,N_7805,N_7796);
or U7966 (N_7966,N_7866,N_7859);
and U7967 (N_7967,N_7874,N_7873);
nand U7968 (N_7968,N_7816,N_7866);
and U7969 (N_7969,N_7775,N_7751);
or U7970 (N_7970,N_7780,N_7796);
and U7971 (N_7971,N_7818,N_7857);
nand U7972 (N_7972,N_7750,N_7779);
xnor U7973 (N_7973,N_7838,N_7776);
nand U7974 (N_7974,N_7773,N_7766);
nand U7975 (N_7975,N_7862,N_7782);
nor U7976 (N_7976,N_7750,N_7753);
and U7977 (N_7977,N_7866,N_7765);
or U7978 (N_7978,N_7775,N_7787);
nand U7979 (N_7979,N_7844,N_7842);
xor U7980 (N_7980,N_7778,N_7764);
nand U7981 (N_7981,N_7850,N_7812);
or U7982 (N_7982,N_7835,N_7763);
nor U7983 (N_7983,N_7790,N_7811);
nor U7984 (N_7984,N_7756,N_7781);
nor U7985 (N_7985,N_7779,N_7768);
and U7986 (N_7986,N_7835,N_7793);
or U7987 (N_7987,N_7795,N_7823);
nor U7988 (N_7988,N_7858,N_7751);
nand U7989 (N_7989,N_7766,N_7831);
or U7990 (N_7990,N_7757,N_7874);
nand U7991 (N_7991,N_7814,N_7793);
xor U7992 (N_7992,N_7786,N_7809);
nand U7993 (N_7993,N_7782,N_7854);
or U7994 (N_7994,N_7817,N_7791);
xnor U7995 (N_7995,N_7864,N_7874);
xnor U7996 (N_7996,N_7837,N_7839);
or U7997 (N_7997,N_7763,N_7874);
and U7998 (N_7998,N_7784,N_7845);
and U7999 (N_7999,N_7822,N_7784);
xnor U8000 (N_8000,N_7980,N_7987);
or U8001 (N_8001,N_7997,N_7999);
xor U8002 (N_8002,N_7978,N_7890);
xor U8003 (N_8003,N_7928,N_7889);
nand U8004 (N_8004,N_7900,N_7960);
nand U8005 (N_8005,N_7952,N_7881);
nand U8006 (N_8006,N_7909,N_7969);
nand U8007 (N_8007,N_7977,N_7917);
nor U8008 (N_8008,N_7914,N_7954);
or U8009 (N_8009,N_7883,N_7902);
and U8010 (N_8010,N_7919,N_7947);
and U8011 (N_8011,N_7945,N_7970);
or U8012 (N_8012,N_7916,N_7894);
nor U8013 (N_8013,N_7913,N_7942);
and U8014 (N_8014,N_7925,N_7955);
xnor U8015 (N_8015,N_7912,N_7944);
and U8016 (N_8016,N_7891,N_7921);
or U8017 (N_8017,N_7972,N_7906);
nor U8018 (N_8018,N_7946,N_7983);
xnor U8019 (N_8019,N_7910,N_7967);
nor U8020 (N_8020,N_7887,N_7896);
nand U8021 (N_8021,N_7905,N_7958);
or U8022 (N_8022,N_7982,N_7880);
nand U8023 (N_8023,N_7961,N_7878);
nand U8024 (N_8024,N_7911,N_7901);
nor U8025 (N_8025,N_7938,N_7975);
nand U8026 (N_8026,N_7991,N_7971);
xnor U8027 (N_8027,N_7993,N_7959);
and U8028 (N_8028,N_7932,N_7988);
nand U8029 (N_8029,N_7918,N_7903);
nor U8030 (N_8030,N_7979,N_7985);
xor U8031 (N_8031,N_7892,N_7957);
xnor U8032 (N_8032,N_7943,N_7968);
nand U8033 (N_8033,N_7966,N_7882);
nor U8034 (N_8034,N_7930,N_7907);
xnor U8035 (N_8035,N_7904,N_7996);
nor U8036 (N_8036,N_7965,N_7875);
and U8037 (N_8037,N_7923,N_7939);
and U8038 (N_8038,N_7927,N_7950);
nor U8039 (N_8039,N_7922,N_7924);
and U8040 (N_8040,N_7908,N_7876);
nor U8041 (N_8041,N_7886,N_7964);
nor U8042 (N_8042,N_7899,N_7879);
xor U8043 (N_8043,N_7933,N_7929);
nand U8044 (N_8044,N_7974,N_7888);
nand U8045 (N_8045,N_7998,N_7984);
xor U8046 (N_8046,N_7934,N_7953);
and U8047 (N_8047,N_7962,N_7948);
or U8048 (N_8048,N_7877,N_7981);
and U8049 (N_8049,N_7893,N_7986);
xor U8050 (N_8050,N_7951,N_7898);
nand U8051 (N_8051,N_7884,N_7995);
nand U8052 (N_8052,N_7937,N_7956);
nor U8053 (N_8053,N_7990,N_7941);
nor U8054 (N_8054,N_7949,N_7931);
and U8055 (N_8055,N_7920,N_7940);
and U8056 (N_8056,N_7926,N_7992);
nand U8057 (N_8057,N_7994,N_7885);
or U8058 (N_8058,N_7897,N_7915);
and U8059 (N_8059,N_7936,N_7989);
nand U8060 (N_8060,N_7935,N_7976);
nand U8061 (N_8061,N_7963,N_7973);
and U8062 (N_8062,N_7895,N_7940);
xnor U8063 (N_8063,N_7890,N_7940);
nand U8064 (N_8064,N_7912,N_7951);
and U8065 (N_8065,N_7921,N_7948);
or U8066 (N_8066,N_7943,N_7972);
and U8067 (N_8067,N_7949,N_7903);
nor U8068 (N_8068,N_7929,N_7887);
xnor U8069 (N_8069,N_7973,N_7905);
xnor U8070 (N_8070,N_7982,N_7978);
xnor U8071 (N_8071,N_7963,N_7935);
or U8072 (N_8072,N_7898,N_7904);
nand U8073 (N_8073,N_7906,N_7956);
nor U8074 (N_8074,N_7895,N_7896);
or U8075 (N_8075,N_7919,N_7903);
nor U8076 (N_8076,N_7885,N_7983);
or U8077 (N_8077,N_7910,N_7975);
xor U8078 (N_8078,N_7890,N_7939);
or U8079 (N_8079,N_7896,N_7954);
and U8080 (N_8080,N_7946,N_7915);
nor U8081 (N_8081,N_7996,N_7999);
xnor U8082 (N_8082,N_7900,N_7977);
or U8083 (N_8083,N_7878,N_7934);
and U8084 (N_8084,N_7996,N_7979);
xor U8085 (N_8085,N_7979,N_7878);
xnor U8086 (N_8086,N_7946,N_7891);
xnor U8087 (N_8087,N_7987,N_7941);
nor U8088 (N_8088,N_7953,N_7907);
or U8089 (N_8089,N_7990,N_7983);
xor U8090 (N_8090,N_7893,N_7990);
or U8091 (N_8091,N_7899,N_7980);
nand U8092 (N_8092,N_7966,N_7916);
or U8093 (N_8093,N_7997,N_7960);
nand U8094 (N_8094,N_7908,N_7959);
or U8095 (N_8095,N_7944,N_7911);
or U8096 (N_8096,N_7880,N_7904);
and U8097 (N_8097,N_7925,N_7941);
nand U8098 (N_8098,N_7929,N_7914);
nand U8099 (N_8099,N_7909,N_7910);
and U8100 (N_8100,N_7941,N_7911);
and U8101 (N_8101,N_7951,N_7897);
nand U8102 (N_8102,N_7958,N_7981);
or U8103 (N_8103,N_7905,N_7893);
and U8104 (N_8104,N_7898,N_7957);
and U8105 (N_8105,N_7951,N_7886);
nand U8106 (N_8106,N_7921,N_7942);
nand U8107 (N_8107,N_7980,N_7887);
xnor U8108 (N_8108,N_7971,N_7899);
and U8109 (N_8109,N_7989,N_7995);
and U8110 (N_8110,N_7880,N_7964);
xnor U8111 (N_8111,N_7891,N_7926);
and U8112 (N_8112,N_7992,N_7881);
nor U8113 (N_8113,N_7998,N_7917);
xnor U8114 (N_8114,N_7999,N_7982);
nor U8115 (N_8115,N_7903,N_7889);
nor U8116 (N_8116,N_7974,N_7993);
xor U8117 (N_8117,N_7878,N_7987);
or U8118 (N_8118,N_7920,N_7875);
nand U8119 (N_8119,N_7964,N_7966);
xor U8120 (N_8120,N_7907,N_7878);
and U8121 (N_8121,N_7976,N_7908);
or U8122 (N_8122,N_7934,N_7975);
and U8123 (N_8123,N_7998,N_7897);
or U8124 (N_8124,N_7882,N_7939);
nand U8125 (N_8125,N_8031,N_8117);
and U8126 (N_8126,N_8058,N_8107);
or U8127 (N_8127,N_8060,N_8067);
and U8128 (N_8128,N_8003,N_8001);
nand U8129 (N_8129,N_8114,N_8044);
or U8130 (N_8130,N_8071,N_8122);
or U8131 (N_8131,N_8028,N_8080);
xor U8132 (N_8132,N_8024,N_8059);
nand U8133 (N_8133,N_8035,N_8082);
nand U8134 (N_8134,N_8045,N_8015);
nor U8135 (N_8135,N_8120,N_8008);
or U8136 (N_8136,N_8066,N_8036);
and U8137 (N_8137,N_8017,N_8108);
nor U8138 (N_8138,N_8097,N_8110);
and U8139 (N_8139,N_8075,N_8009);
or U8140 (N_8140,N_8043,N_8014);
xor U8141 (N_8141,N_8033,N_8104);
nand U8142 (N_8142,N_8023,N_8083);
and U8143 (N_8143,N_8091,N_8070);
or U8144 (N_8144,N_8079,N_8111);
nor U8145 (N_8145,N_8016,N_8027);
xor U8146 (N_8146,N_8012,N_8004);
or U8147 (N_8147,N_8092,N_8102);
nand U8148 (N_8148,N_8022,N_8088);
nor U8149 (N_8149,N_8065,N_8018);
nand U8150 (N_8150,N_8096,N_8051);
nor U8151 (N_8151,N_8098,N_8005);
nor U8152 (N_8152,N_8124,N_8034);
and U8153 (N_8153,N_8119,N_8038);
and U8154 (N_8154,N_8068,N_8085);
xnor U8155 (N_8155,N_8006,N_8076);
xnor U8156 (N_8156,N_8052,N_8103);
xor U8157 (N_8157,N_8081,N_8086);
nand U8158 (N_8158,N_8121,N_8020);
xor U8159 (N_8159,N_8115,N_8109);
nor U8160 (N_8160,N_8049,N_8072);
nor U8161 (N_8161,N_8095,N_8074);
nand U8162 (N_8162,N_8078,N_8010);
and U8163 (N_8163,N_8084,N_8040);
nor U8164 (N_8164,N_8077,N_8046);
nor U8165 (N_8165,N_8118,N_8032);
or U8166 (N_8166,N_8047,N_8000);
or U8167 (N_8167,N_8064,N_8093);
nor U8168 (N_8168,N_8073,N_8056);
xor U8169 (N_8169,N_8041,N_8123);
nand U8170 (N_8170,N_8039,N_8021);
nand U8171 (N_8171,N_8048,N_8087);
nor U8172 (N_8172,N_8007,N_8025);
or U8173 (N_8173,N_8029,N_8116);
xnor U8174 (N_8174,N_8026,N_8053);
nor U8175 (N_8175,N_8055,N_8106);
nor U8176 (N_8176,N_8030,N_8019);
and U8177 (N_8177,N_8105,N_8089);
xnor U8178 (N_8178,N_8013,N_8037);
or U8179 (N_8179,N_8063,N_8050);
xnor U8180 (N_8180,N_8061,N_8057);
xnor U8181 (N_8181,N_8054,N_8002);
and U8182 (N_8182,N_8112,N_8042);
xnor U8183 (N_8183,N_8100,N_8113);
nand U8184 (N_8184,N_8090,N_8099);
and U8185 (N_8185,N_8101,N_8062);
nor U8186 (N_8186,N_8094,N_8011);
xor U8187 (N_8187,N_8069,N_8115);
nand U8188 (N_8188,N_8010,N_8019);
or U8189 (N_8189,N_8124,N_8045);
and U8190 (N_8190,N_8008,N_8038);
nor U8191 (N_8191,N_8096,N_8088);
nand U8192 (N_8192,N_8103,N_8077);
xnor U8193 (N_8193,N_8004,N_8014);
xor U8194 (N_8194,N_8049,N_8024);
nor U8195 (N_8195,N_8007,N_8028);
or U8196 (N_8196,N_8009,N_8102);
or U8197 (N_8197,N_8052,N_8016);
or U8198 (N_8198,N_8087,N_8039);
xnor U8199 (N_8199,N_8060,N_8108);
nor U8200 (N_8200,N_8112,N_8002);
xnor U8201 (N_8201,N_8074,N_8117);
nand U8202 (N_8202,N_8046,N_8051);
and U8203 (N_8203,N_8062,N_8043);
or U8204 (N_8204,N_8027,N_8087);
nor U8205 (N_8205,N_8042,N_8113);
xor U8206 (N_8206,N_8056,N_8106);
nand U8207 (N_8207,N_8112,N_8043);
and U8208 (N_8208,N_8004,N_8119);
xor U8209 (N_8209,N_8102,N_8087);
xnor U8210 (N_8210,N_8101,N_8119);
and U8211 (N_8211,N_8074,N_8079);
and U8212 (N_8212,N_8115,N_8027);
or U8213 (N_8213,N_8017,N_8057);
nor U8214 (N_8214,N_8090,N_8110);
nand U8215 (N_8215,N_8099,N_8022);
xnor U8216 (N_8216,N_8055,N_8102);
nor U8217 (N_8217,N_8006,N_8045);
and U8218 (N_8218,N_8015,N_8078);
xnor U8219 (N_8219,N_8029,N_8024);
or U8220 (N_8220,N_8038,N_8114);
xnor U8221 (N_8221,N_8094,N_8032);
xor U8222 (N_8222,N_8057,N_8104);
nand U8223 (N_8223,N_8049,N_8041);
or U8224 (N_8224,N_8067,N_8090);
and U8225 (N_8225,N_8008,N_8002);
or U8226 (N_8226,N_8048,N_8118);
and U8227 (N_8227,N_8095,N_8054);
nand U8228 (N_8228,N_8082,N_8018);
nor U8229 (N_8229,N_8004,N_8038);
and U8230 (N_8230,N_8114,N_8050);
or U8231 (N_8231,N_8099,N_8050);
and U8232 (N_8232,N_8009,N_8116);
xor U8233 (N_8233,N_8037,N_8109);
and U8234 (N_8234,N_8113,N_8034);
xor U8235 (N_8235,N_8011,N_8077);
or U8236 (N_8236,N_8001,N_8059);
and U8237 (N_8237,N_8090,N_8019);
nand U8238 (N_8238,N_8112,N_8108);
nor U8239 (N_8239,N_8088,N_8019);
nand U8240 (N_8240,N_8038,N_8060);
xnor U8241 (N_8241,N_8065,N_8070);
and U8242 (N_8242,N_8042,N_8082);
or U8243 (N_8243,N_8039,N_8056);
and U8244 (N_8244,N_8076,N_8080);
and U8245 (N_8245,N_8072,N_8019);
xnor U8246 (N_8246,N_8018,N_8038);
nor U8247 (N_8247,N_8003,N_8038);
nand U8248 (N_8248,N_8072,N_8108);
nand U8249 (N_8249,N_8057,N_8005);
nor U8250 (N_8250,N_8232,N_8140);
and U8251 (N_8251,N_8137,N_8169);
nor U8252 (N_8252,N_8186,N_8148);
nand U8253 (N_8253,N_8153,N_8167);
nand U8254 (N_8254,N_8180,N_8247);
nand U8255 (N_8255,N_8245,N_8141);
nand U8256 (N_8256,N_8128,N_8156);
nand U8257 (N_8257,N_8204,N_8130);
and U8258 (N_8258,N_8208,N_8143);
nor U8259 (N_8259,N_8243,N_8157);
or U8260 (N_8260,N_8179,N_8209);
nor U8261 (N_8261,N_8249,N_8218);
nand U8262 (N_8262,N_8211,N_8215);
nand U8263 (N_8263,N_8125,N_8166);
xor U8264 (N_8264,N_8146,N_8216);
xnor U8265 (N_8265,N_8160,N_8225);
or U8266 (N_8266,N_8220,N_8237);
xor U8267 (N_8267,N_8154,N_8203);
nor U8268 (N_8268,N_8223,N_8201);
nor U8269 (N_8269,N_8175,N_8142);
nand U8270 (N_8270,N_8162,N_8219);
nand U8271 (N_8271,N_8199,N_8192);
or U8272 (N_8272,N_8177,N_8246);
and U8273 (N_8273,N_8212,N_8244);
nand U8274 (N_8274,N_8144,N_8139);
and U8275 (N_8275,N_8165,N_8164);
and U8276 (N_8276,N_8231,N_8239);
and U8277 (N_8277,N_8221,N_8240);
nor U8278 (N_8278,N_8197,N_8184);
or U8279 (N_8279,N_8126,N_8133);
xnor U8280 (N_8280,N_8233,N_8127);
nand U8281 (N_8281,N_8202,N_8222);
nand U8282 (N_8282,N_8190,N_8168);
nor U8283 (N_8283,N_8174,N_8196);
nor U8284 (N_8284,N_8213,N_8161);
nor U8285 (N_8285,N_8173,N_8207);
nand U8286 (N_8286,N_8129,N_8226);
nor U8287 (N_8287,N_8236,N_8230);
or U8288 (N_8288,N_8151,N_8241);
nand U8289 (N_8289,N_8135,N_8234);
nor U8290 (N_8290,N_8182,N_8136);
nand U8291 (N_8291,N_8229,N_8238);
nand U8292 (N_8292,N_8198,N_8147);
and U8293 (N_8293,N_8228,N_8210);
nand U8294 (N_8294,N_8242,N_8155);
xnor U8295 (N_8295,N_8152,N_8248);
nor U8296 (N_8296,N_8170,N_8178);
or U8297 (N_8297,N_8159,N_8235);
xor U8298 (N_8298,N_8138,N_8134);
nor U8299 (N_8299,N_8181,N_8171);
or U8300 (N_8300,N_8183,N_8163);
or U8301 (N_8301,N_8150,N_8132);
or U8302 (N_8302,N_8206,N_8200);
xor U8303 (N_8303,N_8131,N_8191);
xnor U8304 (N_8304,N_8224,N_8187);
or U8305 (N_8305,N_8217,N_8194);
and U8306 (N_8306,N_8172,N_8188);
nor U8307 (N_8307,N_8149,N_8193);
xor U8308 (N_8308,N_8176,N_8214);
xor U8309 (N_8309,N_8158,N_8145);
xor U8310 (N_8310,N_8205,N_8189);
nand U8311 (N_8311,N_8227,N_8195);
nand U8312 (N_8312,N_8185,N_8148);
or U8313 (N_8313,N_8168,N_8248);
xnor U8314 (N_8314,N_8163,N_8231);
nor U8315 (N_8315,N_8169,N_8232);
nor U8316 (N_8316,N_8161,N_8157);
or U8317 (N_8317,N_8234,N_8142);
nor U8318 (N_8318,N_8155,N_8172);
xnor U8319 (N_8319,N_8176,N_8200);
xnor U8320 (N_8320,N_8132,N_8148);
or U8321 (N_8321,N_8133,N_8172);
xnor U8322 (N_8322,N_8244,N_8218);
xnor U8323 (N_8323,N_8228,N_8128);
or U8324 (N_8324,N_8181,N_8135);
and U8325 (N_8325,N_8189,N_8206);
or U8326 (N_8326,N_8238,N_8202);
or U8327 (N_8327,N_8232,N_8203);
xnor U8328 (N_8328,N_8177,N_8233);
nor U8329 (N_8329,N_8204,N_8188);
xnor U8330 (N_8330,N_8236,N_8201);
nor U8331 (N_8331,N_8228,N_8187);
nand U8332 (N_8332,N_8218,N_8149);
xnor U8333 (N_8333,N_8153,N_8197);
and U8334 (N_8334,N_8170,N_8195);
or U8335 (N_8335,N_8125,N_8236);
nand U8336 (N_8336,N_8195,N_8237);
nor U8337 (N_8337,N_8193,N_8235);
or U8338 (N_8338,N_8177,N_8160);
and U8339 (N_8339,N_8162,N_8144);
or U8340 (N_8340,N_8188,N_8212);
nand U8341 (N_8341,N_8232,N_8220);
nand U8342 (N_8342,N_8143,N_8236);
or U8343 (N_8343,N_8160,N_8192);
xor U8344 (N_8344,N_8248,N_8228);
xor U8345 (N_8345,N_8204,N_8231);
xor U8346 (N_8346,N_8230,N_8182);
nor U8347 (N_8347,N_8210,N_8165);
nor U8348 (N_8348,N_8172,N_8135);
nor U8349 (N_8349,N_8239,N_8158);
nor U8350 (N_8350,N_8249,N_8199);
nor U8351 (N_8351,N_8216,N_8227);
and U8352 (N_8352,N_8176,N_8148);
xnor U8353 (N_8353,N_8234,N_8180);
or U8354 (N_8354,N_8225,N_8143);
nor U8355 (N_8355,N_8184,N_8237);
nand U8356 (N_8356,N_8241,N_8186);
xor U8357 (N_8357,N_8201,N_8192);
nand U8358 (N_8358,N_8158,N_8141);
or U8359 (N_8359,N_8177,N_8144);
nand U8360 (N_8360,N_8246,N_8179);
or U8361 (N_8361,N_8234,N_8181);
and U8362 (N_8362,N_8187,N_8155);
nor U8363 (N_8363,N_8141,N_8167);
or U8364 (N_8364,N_8210,N_8230);
nor U8365 (N_8365,N_8244,N_8243);
and U8366 (N_8366,N_8216,N_8192);
nor U8367 (N_8367,N_8176,N_8219);
or U8368 (N_8368,N_8151,N_8218);
or U8369 (N_8369,N_8168,N_8240);
nor U8370 (N_8370,N_8145,N_8214);
nand U8371 (N_8371,N_8138,N_8150);
or U8372 (N_8372,N_8147,N_8244);
nand U8373 (N_8373,N_8185,N_8189);
or U8374 (N_8374,N_8220,N_8207);
and U8375 (N_8375,N_8368,N_8259);
nor U8376 (N_8376,N_8338,N_8342);
and U8377 (N_8377,N_8344,N_8372);
nand U8378 (N_8378,N_8332,N_8334);
nand U8379 (N_8379,N_8266,N_8349);
nor U8380 (N_8380,N_8252,N_8320);
nor U8381 (N_8381,N_8297,N_8279);
nor U8382 (N_8382,N_8300,N_8305);
and U8383 (N_8383,N_8251,N_8316);
nor U8384 (N_8384,N_8335,N_8365);
and U8385 (N_8385,N_8264,N_8270);
xnor U8386 (N_8386,N_8275,N_8337);
nor U8387 (N_8387,N_8350,N_8281);
nand U8388 (N_8388,N_8352,N_8361);
and U8389 (N_8389,N_8357,N_8295);
nor U8390 (N_8390,N_8364,N_8291);
nand U8391 (N_8391,N_8345,N_8348);
xnor U8392 (N_8392,N_8339,N_8346);
xor U8393 (N_8393,N_8256,N_8315);
xnor U8394 (N_8394,N_8282,N_8347);
nand U8395 (N_8395,N_8258,N_8362);
nand U8396 (N_8396,N_8318,N_8278);
nor U8397 (N_8397,N_8304,N_8296);
or U8398 (N_8398,N_8373,N_8288);
and U8399 (N_8399,N_8292,N_8301);
xor U8400 (N_8400,N_8269,N_8268);
and U8401 (N_8401,N_8330,N_8336);
nor U8402 (N_8402,N_8359,N_8314);
or U8403 (N_8403,N_8333,N_8354);
or U8404 (N_8404,N_8250,N_8293);
and U8405 (N_8405,N_8323,N_8254);
nand U8406 (N_8406,N_8262,N_8286);
nor U8407 (N_8407,N_8331,N_8255);
xor U8408 (N_8408,N_8307,N_8351);
nand U8409 (N_8409,N_8303,N_8273);
or U8410 (N_8410,N_8366,N_8355);
nor U8411 (N_8411,N_8325,N_8272);
or U8412 (N_8412,N_8322,N_8287);
nor U8413 (N_8413,N_8327,N_8371);
nand U8414 (N_8414,N_8261,N_8358);
nand U8415 (N_8415,N_8298,N_8277);
or U8416 (N_8416,N_8290,N_8367);
xor U8417 (N_8417,N_8353,N_8308);
xnor U8418 (N_8418,N_8294,N_8369);
xnor U8419 (N_8419,N_8319,N_8274);
and U8420 (N_8420,N_8329,N_8276);
or U8421 (N_8421,N_8321,N_8328);
or U8422 (N_8422,N_8302,N_8309);
xor U8423 (N_8423,N_8326,N_8299);
or U8424 (N_8424,N_8310,N_8284);
and U8425 (N_8425,N_8265,N_8285);
and U8426 (N_8426,N_8260,N_8283);
or U8427 (N_8427,N_8306,N_8289);
xor U8428 (N_8428,N_8324,N_8370);
and U8429 (N_8429,N_8356,N_8280);
and U8430 (N_8430,N_8312,N_8313);
and U8431 (N_8431,N_8341,N_8363);
nand U8432 (N_8432,N_8317,N_8340);
and U8433 (N_8433,N_8257,N_8360);
nand U8434 (N_8434,N_8253,N_8374);
and U8435 (N_8435,N_8271,N_8267);
and U8436 (N_8436,N_8263,N_8343);
or U8437 (N_8437,N_8311,N_8302);
and U8438 (N_8438,N_8279,N_8303);
or U8439 (N_8439,N_8282,N_8276);
and U8440 (N_8440,N_8266,N_8319);
nor U8441 (N_8441,N_8265,N_8371);
nand U8442 (N_8442,N_8284,N_8293);
nand U8443 (N_8443,N_8296,N_8271);
nor U8444 (N_8444,N_8259,N_8256);
nand U8445 (N_8445,N_8304,N_8358);
nor U8446 (N_8446,N_8313,N_8286);
nand U8447 (N_8447,N_8314,N_8373);
nand U8448 (N_8448,N_8252,N_8347);
nor U8449 (N_8449,N_8326,N_8335);
and U8450 (N_8450,N_8306,N_8363);
nand U8451 (N_8451,N_8265,N_8365);
nand U8452 (N_8452,N_8292,N_8264);
xnor U8453 (N_8453,N_8333,N_8271);
nor U8454 (N_8454,N_8319,N_8288);
nand U8455 (N_8455,N_8311,N_8266);
nand U8456 (N_8456,N_8267,N_8347);
and U8457 (N_8457,N_8346,N_8371);
and U8458 (N_8458,N_8370,N_8282);
xor U8459 (N_8459,N_8319,N_8283);
nor U8460 (N_8460,N_8322,N_8290);
nor U8461 (N_8461,N_8258,N_8342);
or U8462 (N_8462,N_8318,N_8333);
nor U8463 (N_8463,N_8255,N_8284);
nand U8464 (N_8464,N_8339,N_8264);
and U8465 (N_8465,N_8367,N_8259);
or U8466 (N_8466,N_8293,N_8356);
and U8467 (N_8467,N_8297,N_8286);
nor U8468 (N_8468,N_8324,N_8361);
nor U8469 (N_8469,N_8351,N_8342);
nand U8470 (N_8470,N_8270,N_8351);
xor U8471 (N_8471,N_8308,N_8310);
nor U8472 (N_8472,N_8255,N_8272);
or U8473 (N_8473,N_8357,N_8310);
and U8474 (N_8474,N_8272,N_8341);
or U8475 (N_8475,N_8299,N_8346);
nor U8476 (N_8476,N_8314,N_8251);
xnor U8477 (N_8477,N_8254,N_8288);
xor U8478 (N_8478,N_8268,N_8300);
and U8479 (N_8479,N_8357,N_8308);
and U8480 (N_8480,N_8293,N_8352);
or U8481 (N_8481,N_8370,N_8327);
xor U8482 (N_8482,N_8350,N_8334);
and U8483 (N_8483,N_8363,N_8301);
and U8484 (N_8484,N_8356,N_8265);
and U8485 (N_8485,N_8281,N_8258);
xor U8486 (N_8486,N_8339,N_8321);
nor U8487 (N_8487,N_8319,N_8271);
nand U8488 (N_8488,N_8260,N_8309);
nor U8489 (N_8489,N_8344,N_8304);
xnor U8490 (N_8490,N_8332,N_8264);
nor U8491 (N_8491,N_8260,N_8266);
and U8492 (N_8492,N_8268,N_8260);
or U8493 (N_8493,N_8340,N_8358);
or U8494 (N_8494,N_8272,N_8276);
xnor U8495 (N_8495,N_8280,N_8287);
nand U8496 (N_8496,N_8337,N_8289);
nand U8497 (N_8497,N_8328,N_8360);
nand U8498 (N_8498,N_8266,N_8250);
or U8499 (N_8499,N_8357,N_8331);
xnor U8500 (N_8500,N_8425,N_8436);
nand U8501 (N_8501,N_8486,N_8445);
nor U8502 (N_8502,N_8409,N_8424);
xor U8503 (N_8503,N_8498,N_8396);
or U8504 (N_8504,N_8381,N_8423);
or U8505 (N_8505,N_8400,N_8431);
or U8506 (N_8506,N_8482,N_8438);
xnor U8507 (N_8507,N_8399,N_8418);
nor U8508 (N_8508,N_8469,N_8471);
nand U8509 (N_8509,N_8488,N_8407);
and U8510 (N_8510,N_8384,N_8405);
and U8511 (N_8511,N_8394,N_8446);
xor U8512 (N_8512,N_8476,N_8390);
or U8513 (N_8513,N_8376,N_8475);
nor U8514 (N_8514,N_8404,N_8380);
nand U8515 (N_8515,N_8439,N_8412);
or U8516 (N_8516,N_8429,N_8477);
and U8517 (N_8517,N_8467,N_8426);
and U8518 (N_8518,N_8496,N_8462);
and U8519 (N_8519,N_8422,N_8497);
nand U8520 (N_8520,N_8397,N_8444);
xor U8521 (N_8521,N_8440,N_8421);
nor U8522 (N_8522,N_8434,N_8492);
xor U8523 (N_8523,N_8391,N_8389);
nand U8524 (N_8524,N_8479,N_8478);
xor U8525 (N_8525,N_8393,N_8442);
nand U8526 (N_8526,N_8395,N_8448);
or U8527 (N_8527,N_8435,N_8447);
and U8528 (N_8528,N_8408,N_8377);
or U8529 (N_8529,N_8413,N_8464);
nor U8530 (N_8530,N_8490,N_8388);
and U8531 (N_8531,N_8465,N_8455);
xor U8532 (N_8532,N_8375,N_8449);
nand U8533 (N_8533,N_8378,N_8441);
or U8534 (N_8534,N_8417,N_8483);
and U8535 (N_8535,N_8385,N_8398);
or U8536 (N_8536,N_8415,N_8392);
and U8537 (N_8537,N_8432,N_8484);
and U8538 (N_8538,N_8386,N_8493);
or U8539 (N_8539,N_8379,N_8499);
and U8540 (N_8540,N_8420,N_8419);
xor U8541 (N_8541,N_8402,N_8470);
and U8542 (N_8542,N_8458,N_8454);
xor U8543 (N_8543,N_8457,N_8387);
nor U8544 (N_8544,N_8406,N_8494);
or U8545 (N_8545,N_8473,N_8403);
xor U8546 (N_8546,N_8383,N_8414);
nor U8547 (N_8547,N_8463,N_8428);
xnor U8548 (N_8548,N_8411,N_8382);
and U8549 (N_8549,N_8481,N_8453);
nand U8550 (N_8550,N_8437,N_8451);
nor U8551 (N_8551,N_8495,N_8466);
nor U8552 (N_8552,N_8461,N_8487);
nor U8553 (N_8553,N_8491,N_8427);
nand U8554 (N_8554,N_8459,N_8416);
nand U8555 (N_8555,N_8485,N_8456);
nand U8556 (N_8556,N_8474,N_8430);
nor U8557 (N_8557,N_8410,N_8480);
and U8558 (N_8558,N_8401,N_8472);
nor U8559 (N_8559,N_8460,N_8489);
nand U8560 (N_8560,N_8450,N_8433);
and U8561 (N_8561,N_8468,N_8443);
nor U8562 (N_8562,N_8452,N_8499);
and U8563 (N_8563,N_8444,N_8476);
or U8564 (N_8564,N_8451,N_8456);
nand U8565 (N_8565,N_8396,N_8377);
or U8566 (N_8566,N_8490,N_8496);
nand U8567 (N_8567,N_8418,N_8440);
nor U8568 (N_8568,N_8388,N_8491);
or U8569 (N_8569,N_8488,N_8470);
xnor U8570 (N_8570,N_8466,N_8400);
nor U8571 (N_8571,N_8404,N_8470);
and U8572 (N_8572,N_8479,N_8432);
and U8573 (N_8573,N_8448,N_8426);
xnor U8574 (N_8574,N_8481,N_8413);
nor U8575 (N_8575,N_8412,N_8400);
nor U8576 (N_8576,N_8464,N_8492);
xor U8577 (N_8577,N_8408,N_8475);
xnor U8578 (N_8578,N_8444,N_8388);
nor U8579 (N_8579,N_8381,N_8471);
and U8580 (N_8580,N_8481,N_8448);
and U8581 (N_8581,N_8430,N_8444);
xor U8582 (N_8582,N_8376,N_8381);
nand U8583 (N_8583,N_8462,N_8391);
and U8584 (N_8584,N_8480,N_8469);
or U8585 (N_8585,N_8434,N_8464);
and U8586 (N_8586,N_8381,N_8416);
xor U8587 (N_8587,N_8407,N_8379);
and U8588 (N_8588,N_8431,N_8494);
and U8589 (N_8589,N_8450,N_8460);
nand U8590 (N_8590,N_8449,N_8388);
and U8591 (N_8591,N_8384,N_8381);
nand U8592 (N_8592,N_8477,N_8380);
and U8593 (N_8593,N_8462,N_8411);
xor U8594 (N_8594,N_8384,N_8394);
nand U8595 (N_8595,N_8474,N_8421);
xor U8596 (N_8596,N_8448,N_8411);
nand U8597 (N_8597,N_8480,N_8474);
or U8598 (N_8598,N_8484,N_8399);
nand U8599 (N_8599,N_8399,N_8488);
xor U8600 (N_8600,N_8414,N_8425);
and U8601 (N_8601,N_8377,N_8454);
nor U8602 (N_8602,N_8461,N_8430);
xnor U8603 (N_8603,N_8432,N_8471);
and U8604 (N_8604,N_8455,N_8496);
or U8605 (N_8605,N_8426,N_8481);
xnor U8606 (N_8606,N_8432,N_8463);
nor U8607 (N_8607,N_8459,N_8458);
nor U8608 (N_8608,N_8489,N_8378);
and U8609 (N_8609,N_8462,N_8393);
and U8610 (N_8610,N_8491,N_8450);
xor U8611 (N_8611,N_8434,N_8391);
and U8612 (N_8612,N_8466,N_8499);
xnor U8613 (N_8613,N_8386,N_8447);
xnor U8614 (N_8614,N_8498,N_8411);
and U8615 (N_8615,N_8432,N_8487);
or U8616 (N_8616,N_8429,N_8455);
nor U8617 (N_8617,N_8481,N_8411);
or U8618 (N_8618,N_8430,N_8483);
or U8619 (N_8619,N_8475,N_8417);
or U8620 (N_8620,N_8495,N_8398);
and U8621 (N_8621,N_8420,N_8412);
nand U8622 (N_8622,N_8466,N_8484);
xor U8623 (N_8623,N_8382,N_8432);
xor U8624 (N_8624,N_8485,N_8416);
xor U8625 (N_8625,N_8592,N_8621);
nand U8626 (N_8626,N_8515,N_8553);
nand U8627 (N_8627,N_8543,N_8503);
nor U8628 (N_8628,N_8579,N_8505);
nor U8629 (N_8629,N_8518,N_8568);
xor U8630 (N_8630,N_8549,N_8544);
nor U8631 (N_8631,N_8589,N_8508);
nor U8632 (N_8632,N_8601,N_8525);
and U8633 (N_8633,N_8595,N_8623);
xnor U8634 (N_8634,N_8577,N_8521);
and U8635 (N_8635,N_8562,N_8501);
or U8636 (N_8636,N_8593,N_8547);
and U8637 (N_8637,N_8522,N_8587);
and U8638 (N_8638,N_8514,N_8619);
and U8639 (N_8639,N_8517,N_8563);
or U8640 (N_8640,N_8581,N_8590);
and U8641 (N_8641,N_8616,N_8504);
nor U8642 (N_8642,N_8575,N_8560);
and U8643 (N_8643,N_8507,N_8591);
and U8644 (N_8644,N_8510,N_8598);
nor U8645 (N_8645,N_8573,N_8605);
or U8646 (N_8646,N_8618,N_8578);
or U8647 (N_8647,N_8550,N_8541);
or U8648 (N_8648,N_8609,N_8567);
and U8649 (N_8649,N_8536,N_8556);
nand U8650 (N_8650,N_8596,N_8539);
xor U8651 (N_8651,N_8576,N_8540);
and U8652 (N_8652,N_8574,N_8530);
nand U8653 (N_8653,N_8529,N_8570);
xor U8654 (N_8654,N_8512,N_8502);
or U8655 (N_8655,N_8565,N_8607);
or U8656 (N_8656,N_8602,N_8545);
or U8657 (N_8657,N_8594,N_8558);
xnor U8658 (N_8658,N_8604,N_8555);
and U8659 (N_8659,N_8599,N_8569);
xor U8660 (N_8660,N_8585,N_8511);
and U8661 (N_8661,N_8580,N_8561);
xor U8662 (N_8662,N_8532,N_8551);
and U8663 (N_8663,N_8523,N_8614);
and U8664 (N_8664,N_8584,N_8622);
or U8665 (N_8665,N_8611,N_8613);
or U8666 (N_8666,N_8535,N_8608);
and U8667 (N_8667,N_8500,N_8519);
or U8668 (N_8668,N_8528,N_8548);
and U8669 (N_8669,N_8542,N_8624);
nand U8670 (N_8670,N_8583,N_8617);
and U8671 (N_8671,N_8537,N_8524);
xnor U8672 (N_8672,N_8571,N_8620);
nand U8673 (N_8673,N_8506,N_8600);
nand U8674 (N_8674,N_8513,N_8534);
xor U8675 (N_8675,N_8606,N_8586);
and U8676 (N_8676,N_8610,N_8554);
or U8677 (N_8677,N_8588,N_8582);
and U8678 (N_8678,N_8552,N_8603);
and U8679 (N_8679,N_8572,N_8566);
xor U8680 (N_8680,N_8597,N_8557);
and U8681 (N_8681,N_8615,N_8533);
and U8682 (N_8682,N_8612,N_8526);
or U8683 (N_8683,N_8520,N_8516);
nand U8684 (N_8684,N_8509,N_8564);
nand U8685 (N_8685,N_8559,N_8531);
nor U8686 (N_8686,N_8538,N_8527);
nor U8687 (N_8687,N_8546,N_8507);
or U8688 (N_8688,N_8536,N_8520);
nand U8689 (N_8689,N_8558,N_8530);
nand U8690 (N_8690,N_8541,N_8501);
nand U8691 (N_8691,N_8589,N_8518);
or U8692 (N_8692,N_8535,N_8513);
nand U8693 (N_8693,N_8509,N_8563);
nor U8694 (N_8694,N_8610,N_8555);
and U8695 (N_8695,N_8501,N_8623);
nand U8696 (N_8696,N_8582,N_8614);
or U8697 (N_8697,N_8610,N_8596);
xor U8698 (N_8698,N_8582,N_8538);
xor U8699 (N_8699,N_8614,N_8506);
and U8700 (N_8700,N_8555,N_8503);
xor U8701 (N_8701,N_8593,N_8595);
and U8702 (N_8702,N_8580,N_8573);
nand U8703 (N_8703,N_8510,N_8556);
or U8704 (N_8704,N_8604,N_8522);
or U8705 (N_8705,N_8585,N_8530);
nor U8706 (N_8706,N_8595,N_8579);
or U8707 (N_8707,N_8601,N_8587);
xor U8708 (N_8708,N_8603,N_8596);
or U8709 (N_8709,N_8577,N_8576);
and U8710 (N_8710,N_8551,N_8512);
nor U8711 (N_8711,N_8615,N_8599);
xnor U8712 (N_8712,N_8517,N_8616);
nor U8713 (N_8713,N_8519,N_8571);
nand U8714 (N_8714,N_8528,N_8525);
and U8715 (N_8715,N_8579,N_8566);
or U8716 (N_8716,N_8577,N_8545);
nor U8717 (N_8717,N_8621,N_8532);
and U8718 (N_8718,N_8570,N_8517);
and U8719 (N_8719,N_8565,N_8515);
nand U8720 (N_8720,N_8565,N_8604);
or U8721 (N_8721,N_8586,N_8612);
xor U8722 (N_8722,N_8512,N_8573);
nor U8723 (N_8723,N_8502,N_8501);
nand U8724 (N_8724,N_8582,N_8529);
nor U8725 (N_8725,N_8616,N_8601);
and U8726 (N_8726,N_8592,N_8612);
and U8727 (N_8727,N_8532,N_8578);
xor U8728 (N_8728,N_8624,N_8551);
and U8729 (N_8729,N_8528,N_8591);
or U8730 (N_8730,N_8549,N_8502);
nand U8731 (N_8731,N_8555,N_8622);
nor U8732 (N_8732,N_8548,N_8582);
and U8733 (N_8733,N_8536,N_8528);
nor U8734 (N_8734,N_8541,N_8575);
and U8735 (N_8735,N_8526,N_8556);
or U8736 (N_8736,N_8510,N_8562);
and U8737 (N_8737,N_8590,N_8517);
xnor U8738 (N_8738,N_8521,N_8532);
nand U8739 (N_8739,N_8598,N_8558);
nand U8740 (N_8740,N_8514,N_8532);
or U8741 (N_8741,N_8605,N_8591);
and U8742 (N_8742,N_8613,N_8592);
xnor U8743 (N_8743,N_8549,N_8580);
nor U8744 (N_8744,N_8529,N_8504);
or U8745 (N_8745,N_8553,N_8581);
nand U8746 (N_8746,N_8543,N_8585);
or U8747 (N_8747,N_8608,N_8611);
and U8748 (N_8748,N_8572,N_8514);
nor U8749 (N_8749,N_8621,N_8602);
or U8750 (N_8750,N_8668,N_8744);
nand U8751 (N_8751,N_8667,N_8718);
and U8752 (N_8752,N_8637,N_8682);
nor U8753 (N_8753,N_8742,N_8672);
nor U8754 (N_8754,N_8656,N_8648);
xnor U8755 (N_8755,N_8629,N_8707);
nand U8756 (N_8756,N_8642,N_8699);
and U8757 (N_8757,N_8715,N_8678);
xor U8758 (N_8758,N_8709,N_8655);
and U8759 (N_8759,N_8694,N_8743);
or U8760 (N_8760,N_8640,N_8739);
nand U8761 (N_8761,N_8703,N_8677);
or U8762 (N_8762,N_8671,N_8644);
nor U8763 (N_8763,N_8670,N_8734);
xor U8764 (N_8764,N_8690,N_8695);
and U8765 (N_8765,N_8631,N_8686);
xnor U8766 (N_8766,N_8630,N_8635);
and U8767 (N_8767,N_8700,N_8738);
xnor U8768 (N_8768,N_8691,N_8645);
nor U8769 (N_8769,N_8727,N_8654);
xor U8770 (N_8770,N_8701,N_8675);
nor U8771 (N_8771,N_8661,N_8726);
nand U8772 (N_8772,N_8748,N_8721);
or U8773 (N_8773,N_8712,N_8710);
or U8774 (N_8774,N_8662,N_8728);
or U8775 (N_8775,N_8692,N_8716);
and U8776 (N_8776,N_8723,N_8657);
and U8777 (N_8777,N_8674,N_8650);
or U8778 (N_8778,N_8636,N_8646);
nand U8779 (N_8779,N_8653,N_8731);
nor U8780 (N_8780,N_8740,N_8664);
nand U8781 (N_8781,N_8706,N_8689);
nor U8782 (N_8782,N_8651,N_8719);
and U8783 (N_8783,N_8698,N_8736);
and U8784 (N_8784,N_8633,N_8717);
nand U8785 (N_8785,N_8649,N_8685);
or U8786 (N_8786,N_8625,N_8666);
or U8787 (N_8787,N_8659,N_8696);
xor U8788 (N_8788,N_8708,N_8679);
or U8789 (N_8789,N_8724,N_8729);
or U8790 (N_8790,N_8632,N_8628);
nor U8791 (N_8791,N_8722,N_8658);
xnor U8792 (N_8792,N_8673,N_8697);
nor U8793 (N_8793,N_8720,N_8688);
nand U8794 (N_8794,N_8693,N_8730);
nand U8795 (N_8795,N_8735,N_8733);
xor U8796 (N_8796,N_8749,N_8627);
xnor U8797 (N_8797,N_8652,N_8714);
or U8798 (N_8798,N_8745,N_8663);
nand U8799 (N_8799,N_8626,N_8704);
xor U8800 (N_8800,N_8676,N_8669);
xor U8801 (N_8801,N_8741,N_8687);
nor U8802 (N_8802,N_8639,N_8705);
or U8803 (N_8803,N_8747,N_8711);
xor U8804 (N_8804,N_8680,N_8643);
and U8805 (N_8805,N_8732,N_8638);
nand U8806 (N_8806,N_8746,N_8725);
nor U8807 (N_8807,N_8681,N_8737);
nand U8808 (N_8808,N_8684,N_8647);
nor U8809 (N_8809,N_8683,N_8713);
and U8810 (N_8810,N_8660,N_8665);
nand U8811 (N_8811,N_8702,N_8634);
or U8812 (N_8812,N_8641,N_8674);
or U8813 (N_8813,N_8697,N_8643);
and U8814 (N_8814,N_8738,N_8636);
or U8815 (N_8815,N_8713,N_8647);
nor U8816 (N_8816,N_8660,N_8632);
xnor U8817 (N_8817,N_8658,N_8729);
nor U8818 (N_8818,N_8744,N_8699);
and U8819 (N_8819,N_8655,N_8701);
or U8820 (N_8820,N_8732,N_8657);
nand U8821 (N_8821,N_8662,N_8651);
nand U8822 (N_8822,N_8672,N_8749);
nor U8823 (N_8823,N_8691,N_8663);
nand U8824 (N_8824,N_8648,N_8654);
nand U8825 (N_8825,N_8714,N_8646);
or U8826 (N_8826,N_8710,N_8634);
or U8827 (N_8827,N_8658,N_8709);
nor U8828 (N_8828,N_8712,N_8697);
and U8829 (N_8829,N_8743,N_8672);
or U8830 (N_8830,N_8684,N_8701);
nor U8831 (N_8831,N_8720,N_8631);
and U8832 (N_8832,N_8668,N_8639);
and U8833 (N_8833,N_8696,N_8711);
xor U8834 (N_8834,N_8722,N_8640);
nand U8835 (N_8835,N_8675,N_8707);
nand U8836 (N_8836,N_8660,N_8657);
nand U8837 (N_8837,N_8723,N_8647);
and U8838 (N_8838,N_8701,N_8744);
and U8839 (N_8839,N_8643,N_8641);
xor U8840 (N_8840,N_8728,N_8651);
xnor U8841 (N_8841,N_8655,N_8641);
nor U8842 (N_8842,N_8749,N_8659);
nor U8843 (N_8843,N_8713,N_8648);
or U8844 (N_8844,N_8653,N_8663);
xor U8845 (N_8845,N_8648,N_8647);
nand U8846 (N_8846,N_8637,N_8723);
or U8847 (N_8847,N_8680,N_8678);
and U8848 (N_8848,N_8685,N_8645);
nor U8849 (N_8849,N_8741,N_8749);
xor U8850 (N_8850,N_8644,N_8731);
and U8851 (N_8851,N_8749,N_8647);
nor U8852 (N_8852,N_8718,N_8710);
nor U8853 (N_8853,N_8643,N_8705);
or U8854 (N_8854,N_8748,N_8650);
or U8855 (N_8855,N_8692,N_8657);
or U8856 (N_8856,N_8675,N_8700);
or U8857 (N_8857,N_8647,N_8639);
nor U8858 (N_8858,N_8673,N_8666);
and U8859 (N_8859,N_8662,N_8635);
or U8860 (N_8860,N_8645,N_8726);
xnor U8861 (N_8861,N_8729,N_8640);
and U8862 (N_8862,N_8671,N_8631);
nor U8863 (N_8863,N_8700,N_8655);
nor U8864 (N_8864,N_8666,N_8654);
or U8865 (N_8865,N_8730,N_8661);
nor U8866 (N_8866,N_8680,N_8722);
or U8867 (N_8867,N_8695,N_8700);
nand U8868 (N_8868,N_8692,N_8653);
or U8869 (N_8869,N_8668,N_8693);
nor U8870 (N_8870,N_8692,N_8665);
and U8871 (N_8871,N_8730,N_8708);
xor U8872 (N_8872,N_8669,N_8634);
or U8873 (N_8873,N_8643,N_8642);
or U8874 (N_8874,N_8690,N_8703);
nand U8875 (N_8875,N_8796,N_8872);
xnor U8876 (N_8876,N_8808,N_8787);
nor U8877 (N_8877,N_8803,N_8871);
nand U8878 (N_8878,N_8860,N_8790);
nor U8879 (N_8879,N_8859,N_8816);
or U8880 (N_8880,N_8777,N_8858);
xnor U8881 (N_8881,N_8812,N_8759);
or U8882 (N_8882,N_8765,N_8755);
nor U8883 (N_8883,N_8842,N_8753);
nor U8884 (N_8884,N_8768,N_8811);
nor U8885 (N_8885,N_8763,N_8820);
or U8886 (N_8886,N_8774,N_8800);
and U8887 (N_8887,N_8764,N_8813);
xor U8888 (N_8888,N_8769,N_8868);
and U8889 (N_8889,N_8761,N_8821);
xnor U8890 (N_8890,N_8855,N_8861);
and U8891 (N_8891,N_8865,N_8810);
and U8892 (N_8892,N_8791,N_8853);
xnor U8893 (N_8893,N_8815,N_8788);
or U8894 (N_8894,N_8854,N_8819);
and U8895 (N_8895,N_8784,N_8778);
and U8896 (N_8896,N_8832,N_8822);
nand U8897 (N_8897,N_8802,N_8841);
or U8898 (N_8898,N_8845,N_8801);
and U8899 (N_8899,N_8852,N_8838);
or U8900 (N_8900,N_8762,N_8776);
nand U8901 (N_8901,N_8773,N_8869);
xnor U8902 (N_8902,N_8857,N_8798);
and U8903 (N_8903,N_8847,N_8760);
or U8904 (N_8904,N_8794,N_8785);
and U8905 (N_8905,N_8766,N_8837);
nor U8906 (N_8906,N_8767,N_8867);
nor U8907 (N_8907,N_8831,N_8835);
and U8908 (N_8908,N_8848,N_8809);
nor U8909 (N_8909,N_8843,N_8770);
nand U8910 (N_8910,N_8756,N_8817);
or U8911 (N_8911,N_8789,N_8874);
nor U8912 (N_8912,N_8786,N_8829);
xor U8913 (N_8913,N_8870,N_8839);
xnor U8914 (N_8914,N_8846,N_8863);
and U8915 (N_8915,N_8752,N_8873);
or U8916 (N_8916,N_8836,N_8771);
and U8917 (N_8917,N_8782,N_8824);
nor U8918 (N_8918,N_8757,N_8779);
nand U8919 (N_8919,N_8797,N_8783);
nor U8920 (N_8920,N_8856,N_8825);
or U8921 (N_8921,N_8830,N_8754);
and U8922 (N_8922,N_8805,N_8807);
and U8923 (N_8923,N_8781,N_8758);
nor U8924 (N_8924,N_8775,N_8792);
or U8925 (N_8925,N_8862,N_8814);
and U8926 (N_8926,N_8751,N_8780);
and U8927 (N_8927,N_8840,N_8804);
and U8928 (N_8928,N_8799,N_8826);
and U8929 (N_8929,N_8864,N_8806);
or U8930 (N_8930,N_8795,N_8793);
nor U8931 (N_8931,N_8833,N_8823);
or U8932 (N_8932,N_8834,N_8827);
or U8933 (N_8933,N_8828,N_8850);
or U8934 (N_8934,N_8851,N_8750);
and U8935 (N_8935,N_8772,N_8818);
nor U8936 (N_8936,N_8849,N_8866);
or U8937 (N_8937,N_8844,N_8804);
and U8938 (N_8938,N_8863,N_8767);
and U8939 (N_8939,N_8862,N_8769);
xnor U8940 (N_8940,N_8797,N_8765);
nand U8941 (N_8941,N_8780,N_8782);
nand U8942 (N_8942,N_8824,N_8759);
nand U8943 (N_8943,N_8825,N_8860);
xnor U8944 (N_8944,N_8863,N_8788);
xnor U8945 (N_8945,N_8751,N_8804);
or U8946 (N_8946,N_8800,N_8831);
and U8947 (N_8947,N_8872,N_8844);
and U8948 (N_8948,N_8829,N_8864);
nor U8949 (N_8949,N_8772,N_8784);
nor U8950 (N_8950,N_8793,N_8824);
nand U8951 (N_8951,N_8777,N_8841);
or U8952 (N_8952,N_8856,N_8831);
nand U8953 (N_8953,N_8831,N_8793);
and U8954 (N_8954,N_8826,N_8778);
nand U8955 (N_8955,N_8815,N_8843);
nor U8956 (N_8956,N_8757,N_8767);
nor U8957 (N_8957,N_8816,N_8768);
and U8958 (N_8958,N_8794,N_8808);
and U8959 (N_8959,N_8761,N_8846);
or U8960 (N_8960,N_8772,N_8797);
xor U8961 (N_8961,N_8844,N_8823);
xnor U8962 (N_8962,N_8814,N_8797);
xnor U8963 (N_8963,N_8764,N_8799);
and U8964 (N_8964,N_8782,N_8781);
nor U8965 (N_8965,N_8844,N_8765);
nand U8966 (N_8966,N_8758,N_8866);
or U8967 (N_8967,N_8811,N_8830);
nand U8968 (N_8968,N_8832,N_8766);
nor U8969 (N_8969,N_8841,N_8812);
nand U8970 (N_8970,N_8816,N_8775);
and U8971 (N_8971,N_8763,N_8761);
xor U8972 (N_8972,N_8809,N_8783);
or U8973 (N_8973,N_8773,N_8759);
and U8974 (N_8974,N_8761,N_8852);
or U8975 (N_8975,N_8783,N_8769);
xor U8976 (N_8976,N_8756,N_8789);
xnor U8977 (N_8977,N_8829,N_8787);
nor U8978 (N_8978,N_8832,N_8846);
nor U8979 (N_8979,N_8805,N_8779);
or U8980 (N_8980,N_8857,N_8790);
and U8981 (N_8981,N_8776,N_8871);
nor U8982 (N_8982,N_8799,N_8812);
xor U8983 (N_8983,N_8824,N_8830);
nor U8984 (N_8984,N_8818,N_8817);
or U8985 (N_8985,N_8765,N_8823);
nand U8986 (N_8986,N_8799,N_8863);
or U8987 (N_8987,N_8839,N_8841);
xnor U8988 (N_8988,N_8788,N_8829);
or U8989 (N_8989,N_8801,N_8798);
and U8990 (N_8990,N_8814,N_8868);
or U8991 (N_8991,N_8844,N_8856);
xor U8992 (N_8992,N_8762,N_8855);
nand U8993 (N_8993,N_8819,N_8863);
xor U8994 (N_8994,N_8810,N_8789);
nand U8995 (N_8995,N_8872,N_8763);
and U8996 (N_8996,N_8753,N_8762);
or U8997 (N_8997,N_8793,N_8844);
nor U8998 (N_8998,N_8752,N_8841);
or U8999 (N_8999,N_8871,N_8784);
xnor U9000 (N_9000,N_8917,N_8983);
nor U9001 (N_9001,N_8893,N_8885);
nor U9002 (N_9002,N_8891,N_8950);
xor U9003 (N_9003,N_8899,N_8909);
xor U9004 (N_9004,N_8911,N_8970);
and U9005 (N_9005,N_8992,N_8961);
xor U9006 (N_9006,N_8962,N_8916);
xor U9007 (N_9007,N_8995,N_8948);
nand U9008 (N_9008,N_8875,N_8957);
xor U9009 (N_9009,N_8912,N_8902);
nand U9010 (N_9010,N_8939,N_8947);
xnor U9011 (N_9011,N_8982,N_8977);
and U9012 (N_9012,N_8969,N_8920);
nand U9013 (N_9013,N_8965,N_8928);
xor U9014 (N_9014,N_8910,N_8941);
nor U9015 (N_9015,N_8903,N_8888);
or U9016 (N_9016,N_8897,N_8921);
and U9017 (N_9017,N_8998,N_8956);
or U9018 (N_9018,N_8945,N_8879);
or U9019 (N_9019,N_8878,N_8913);
nand U9020 (N_9020,N_8975,N_8937);
and U9021 (N_9021,N_8930,N_8883);
nor U9022 (N_9022,N_8907,N_8966);
or U9023 (N_9023,N_8933,N_8960);
nand U9024 (N_9024,N_8968,N_8896);
xnor U9025 (N_9025,N_8991,N_8889);
xor U9026 (N_9026,N_8989,N_8959);
nand U9027 (N_9027,N_8924,N_8895);
or U9028 (N_9028,N_8876,N_8953);
nand U9029 (N_9029,N_8993,N_8927);
or U9030 (N_9030,N_8944,N_8890);
nand U9031 (N_9031,N_8881,N_8978);
nor U9032 (N_9032,N_8923,N_8931);
nor U9033 (N_9033,N_8922,N_8994);
nand U9034 (N_9034,N_8943,N_8954);
nand U9035 (N_9035,N_8996,N_8882);
or U9036 (N_9036,N_8949,N_8986);
and U9037 (N_9037,N_8951,N_8946);
xor U9038 (N_9038,N_8926,N_8940);
nor U9039 (N_9039,N_8999,N_8990);
xnor U9040 (N_9040,N_8971,N_8886);
nor U9041 (N_9041,N_8898,N_8936);
and U9042 (N_9042,N_8919,N_8938);
xnor U9043 (N_9043,N_8918,N_8894);
and U9044 (N_9044,N_8987,N_8973);
xor U9045 (N_9045,N_8981,N_8932);
nand U9046 (N_9046,N_8901,N_8905);
xnor U9047 (N_9047,N_8972,N_8877);
or U9048 (N_9048,N_8985,N_8892);
or U9049 (N_9049,N_8914,N_8934);
xnor U9050 (N_9050,N_8955,N_8988);
nand U9051 (N_9051,N_8958,N_8979);
xnor U9052 (N_9052,N_8964,N_8963);
nand U9053 (N_9053,N_8929,N_8967);
or U9054 (N_9054,N_8984,N_8906);
nor U9055 (N_9055,N_8880,N_8976);
nand U9056 (N_9056,N_8904,N_8952);
xor U9057 (N_9057,N_8900,N_8908);
or U9058 (N_9058,N_8884,N_8925);
nor U9059 (N_9059,N_8974,N_8942);
or U9060 (N_9060,N_8997,N_8980);
or U9061 (N_9061,N_8915,N_8887);
xor U9062 (N_9062,N_8935,N_8894);
xor U9063 (N_9063,N_8905,N_8921);
and U9064 (N_9064,N_8973,N_8938);
and U9065 (N_9065,N_8938,N_8887);
nor U9066 (N_9066,N_8959,N_8950);
nor U9067 (N_9067,N_8986,N_8959);
nand U9068 (N_9068,N_8896,N_8939);
and U9069 (N_9069,N_8967,N_8882);
xor U9070 (N_9070,N_8981,N_8977);
nor U9071 (N_9071,N_8980,N_8877);
xor U9072 (N_9072,N_8897,N_8968);
xor U9073 (N_9073,N_8935,N_8937);
xnor U9074 (N_9074,N_8997,N_8927);
nand U9075 (N_9075,N_8962,N_8972);
nor U9076 (N_9076,N_8999,N_8886);
nor U9077 (N_9077,N_8943,N_8970);
nand U9078 (N_9078,N_8991,N_8910);
and U9079 (N_9079,N_8964,N_8958);
xor U9080 (N_9080,N_8955,N_8906);
or U9081 (N_9081,N_8968,N_8904);
nand U9082 (N_9082,N_8953,N_8963);
or U9083 (N_9083,N_8985,N_8909);
nand U9084 (N_9084,N_8935,N_8903);
or U9085 (N_9085,N_8985,N_8908);
xnor U9086 (N_9086,N_8904,N_8986);
nand U9087 (N_9087,N_8962,N_8930);
xnor U9088 (N_9088,N_8980,N_8921);
nor U9089 (N_9089,N_8956,N_8935);
xnor U9090 (N_9090,N_8884,N_8997);
xor U9091 (N_9091,N_8998,N_8878);
or U9092 (N_9092,N_8960,N_8973);
nor U9093 (N_9093,N_8890,N_8900);
xnor U9094 (N_9094,N_8956,N_8875);
xnor U9095 (N_9095,N_8904,N_8875);
xnor U9096 (N_9096,N_8907,N_8957);
nand U9097 (N_9097,N_8937,N_8996);
nand U9098 (N_9098,N_8939,N_8940);
nor U9099 (N_9099,N_8917,N_8973);
and U9100 (N_9100,N_8876,N_8928);
nor U9101 (N_9101,N_8992,N_8981);
nand U9102 (N_9102,N_8954,N_8936);
nand U9103 (N_9103,N_8924,N_8923);
or U9104 (N_9104,N_8997,N_8991);
nor U9105 (N_9105,N_8939,N_8899);
nand U9106 (N_9106,N_8995,N_8879);
nand U9107 (N_9107,N_8928,N_8954);
nor U9108 (N_9108,N_8900,N_8931);
nand U9109 (N_9109,N_8886,N_8892);
xor U9110 (N_9110,N_8899,N_8992);
and U9111 (N_9111,N_8929,N_8993);
nor U9112 (N_9112,N_8928,N_8903);
nand U9113 (N_9113,N_8927,N_8885);
xor U9114 (N_9114,N_8946,N_8885);
nor U9115 (N_9115,N_8948,N_8875);
and U9116 (N_9116,N_8970,N_8882);
and U9117 (N_9117,N_8920,N_8946);
and U9118 (N_9118,N_8936,N_8926);
xor U9119 (N_9119,N_8876,N_8924);
and U9120 (N_9120,N_8882,N_8877);
xor U9121 (N_9121,N_8903,N_8944);
xor U9122 (N_9122,N_8944,N_8931);
xnor U9123 (N_9123,N_8990,N_8934);
and U9124 (N_9124,N_8959,N_8951);
or U9125 (N_9125,N_9006,N_9063);
and U9126 (N_9126,N_9044,N_9010);
xnor U9127 (N_9127,N_9085,N_9122);
nand U9128 (N_9128,N_9081,N_9090);
or U9129 (N_9129,N_9113,N_9020);
or U9130 (N_9130,N_9075,N_9109);
or U9131 (N_9131,N_9032,N_9108);
nor U9132 (N_9132,N_9016,N_9118);
xnor U9133 (N_9133,N_9022,N_9028);
and U9134 (N_9134,N_9121,N_9065);
xnor U9135 (N_9135,N_9027,N_9002);
and U9136 (N_9136,N_9106,N_9092);
nand U9137 (N_9137,N_9064,N_9023);
nand U9138 (N_9138,N_9042,N_9116);
nand U9139 (N_9139,N_9001,N_9107);
xor U9140 (N_9140,N_9112,N_9052);
nand U9141 (N_9141,N_9101,N_9005);
xor U9142 (N_9142,N_9040,N_9083);
or U9143 (N_9143,N_9119,N_9031);
and U9144 (N_9144,N_9036,N_9060);
and U9145 (N_9145,N_9067,N_9084);
and U9146 (N_9146,N_9077,N_9007);
nor U9147 (N_9147,N_9009,N_9008);
xor U9148 (N_9148,N_9111,N_9004);
nand U9149 (N_9149,N_9057,N_9114);
nor U9150 (N_9150,N_9079,N_9026);
and U9151 (N_9151,N_9034,N_9073);
nand U9152 (N_9152,N_9033,N_9029);
or U9153 (N_9153,N_9049,N_9050);
nand U9154 (N_9154,N_9070,N_9015);
xor U9155 (N_9155,N_9030,N_9066);
nand U9156 (N_9156,N_9089,N_9071);
and U9157 (N_9157,N_9093,N_9046);
nor U9158 (N_9158,N_9061,N_9014);
xnor U9159 (N_9159,N_9074,N_9000);
nand U9160 (N_9160,N_9123,N_9087);
nor U9161 (N_9161,N_9102,N_9012);
and U9162 (N_9162,N_9105,N_9120);
and U9163 (N_9163,N_9035,N_9094);
nor U9164 (N_9164,N_9037,N_9098);
nor U9165 (N_9165,N_9110,N_9096);
nand U9166 (N_9166,N_9018,N_9099);
nor U9167 (N_9167,N_9059,N_9100);
or U9168 (N_9168,N_9097,N_9080);
nand U9169 (N_9169,N_9086,N_9104);
nor U9170 (N_9170,N_9051,N_9039);
nand U9171 (N_9171,N_9103,N_9024);
nor U9172 (N_9172,N_9047,N_9025);
xnor U9173 (N_9173,N_9056,N_9055);
or U9174 (N_9174,N_9017,N_9043);
or U9175 (N_9175,N_9062,N_9058);
or U9176 (N_9176,N_9021,N_9045);
and U9177 (N_9177,N_9117,N_9078);
xor U9178 (N_9178,N_9013,N_9072);
nor U9179 (N_9179,N_9054,N_9003);
and U9180 (N_9180,N_9011,N_9048);
and U9181 (N_9181,N_9091,N_9069);
or U9182 (N_9182,N_9053,N_9124);
nor U9183 (N_9183,N_9082,N_9041);
xor U9184 (N_9184,N_9019,N_9068);
nand U9185 (N_9185,N_9088,N_9038);
xnor U9186 (N_9186,N_9115,N_9076);
or U9187 (N_9187,N_9095,N_9091);
xnor U9188 (N_9188,N_9041,N_9078);
xor U9189 (N_9189,N_9101,N_9059);
or U9190 (N_9190,N_9060,N_9001);
nor U9191 (N_9191,N_9054,N_9082);
nor U9192 (N_9192,N_9037,N_9026);
nand U9193 (N_9193,N_9006,N_9060);
xnor U9194 (N_9194,N_9120,N_9027);
xor U9195 (N_9195,N_9017,N_9068);
or U9196 (N_9196,N_9004,N_9003);
and U9197 (N_9197,N_9053,N_9008);
or U9198 (N_9198,N_9011,N_9019);
nor U9199 (N_9199,N_9086,N_9097);
nor U9200 (N_9200,N_9065,N_9064);
or U9201 (N_9201,N_9062,N_9039);
or U9202 (N_9202,N_9036,N_9087);
nand U9203 (N_9203,N_9106,N_9033);
nor U9204 (N_9204,N_9024,N_9100);
or U9205 (N_9205,N_9007,N_9076);
or U9206 (N_9206,N_9062,N_9064);
xnor U9207 (N_9207,N_9040,N_9084);
nand U9208 (N_9208,N_9019,N_9099);
and U9209 (N_9209,N_9109,N_9054);
xnor U9210 (N_9210,N_9105,N_9025);
and U9211 (N_9211,N_9122,N_9091);
nand U9212 (N_9212,N_9067,N_9017);
nor U9213 (N_9213,N_9019,N_9037);
and U9214 (N_9214,N_9075,N_9014);
nor U9215 (N_9215,N_9102,N_9005);
nand U9216 (N_9216,N_9038,N_9014);
or U9217 (N_9217,N_9005,N_9021);
nand U9218 (N_9218,N_9027,N_9101);
or U9219 (N_9219,N_9079,N_9064);
nor U9220 (N_9220,N_9110,N_9083);
nor U9221 (N_9221,N_9051,N_9091);
and U9222 (N_9222,N_9084,N_9000);
and U9223 (N_9223,N_9098,N_9114);
nand U9224 (N_9224,N_9109,N_9118);
and U9225 (N_9225,N_9056,N_9042);
nand U9226 (N_9226,N_9031,N_9124);
xor U9227 (N_9227,N_9008,N_9112);
nor U9228 (N_9228,N_9107,N_9015);
xnor U9229 (N_9229,N_9084,N_9081);
or U9230 (N_9230,N_9010,N_9049);
nor U9231 (N_9231,N_9046,N_9028);
or U9232 (N_9232,N_9026,N_9008);
nor U9233 (N_9233,N_9035,N_9038);
nand U9234 (N_9234,N_9077,N_9014);
or U9235 (N_9235,N_9028,N_9035);
and U9236 (N_9236,N_9018,N_9037);
nor U9237 (N_9237,N_9028,N_9062);
nor U9238 (N_9238,N_9105,N_9115);
and U9239 (N_9239,N_9093,N_9054);
nand U9240 (N_9240,N_9004,N_9104);
nand U9241 (N_9241,N_9017,N_9063);
nor U9242 (N_9242,N_9041,N_9006);
and U9243 (N_9243,N_9062,N_9075);
xnor U9244 (N_9244,N_9096,N_9050);
nand U9245 (N_9245,N_9054,N_9030);
nand U9246 (N_9246,N_9089,N_9063);
xnor U9247 (N_9247,N_9107,N_9095);
nor U9248 (N_9248,N_9090,N_9095);
nor U9249 (N_9249,N_9019,N_9001);
or U9250 (N_9250,N_9183,N_9209);
nand U9251 (N_9251,N_9171,N_9249);
xor U9252 (N_9252,N_9133,N_9141);
xor U9253 (N_9253,N_9158,N_9213);
nand U9254 (N_9254,N_9174,N_9159);
and U9255 (N_9255,N_9223,N_9188);
nand U9256 (N_9256,N_9182,N_9177);
and U9257 (N_9257,N_9246,N_9164);
xnor U9258 (N_9258,N_9211,N_9229);
nor U9259 (N_9259,N_9169,N_9204);
nand U9260 (N_9260,N_9201,N_9151);
or U9261 (N_9261,N_9184,N_9138);
nor U9262 (N_9262,N_9137,N_9206);
nand U9263 (N_9263,N_9156,N_9129);
and U9264 (N_9264,N_9203,N_9217);
xnor U9265 (N_9265,N_9163,N_9227);
nand U9266 (N_9266,N_9221,N_9170);
and U9267 (N_9267,N_9236,N_9168);
nand U9268 (N_9268,N_9199,N_9161);
nand U9269 (N_9269,N_9153,N_9136);
xnor U9270 (N_9270,N_9134,N_9140);
or U9271 (N_9271,N_9145,N_9131);
nand U9272 (N_9272,N_9200,N_9150);
and U9273 (N_9273,N_9216,N_9218);
nand U9274 (N_9274,N_9132,N_9152);
and U9275 (N_9275,N_9226,N_9241);
nand U9276 (N_9276,N_9235,N_9245);
nor U9277 (N_9277,N_9202,N_9233);
or U9278 (N_9278,N_9197,N_9157);
nand U9279 (N_9279,N_9191,N_9192);
and U9280 (N_9280,N_9176,N_9194);
and U9281 (N_9281,N_9180,N_9208);
and U9282 (N_9282,N_9173,N_9220);
nor U9283 (N_9283,N_9127,N_9237);
and U9284 (N_9284,N_9231,N_9243);
or U9285 (N_9285,N_9146,N_9219);
or U9286 (N_9286,N_9149,N_9139);
nand U9287 (N_9287,N_9207,N_9125);
and U9288 (N_9288,N_9166,N_9214);
xor U9289 (N_9289,N_9198,N_9155);
xor U9290 (N_9290,N_9135,N_9195);
and U9291 (N_9291,N_9178,N_9228);
xor U9292 (N_9292,N_9160,N_9230);
nor U9293 (N_9293,N_9225,N_9148);
and U9294 (N_9294,N_9143,N_9224);
and U9295 (N_9295,N_9205,N_9185);
xnor U9296 (N_9296,N_9179,N_9187);
nand U9297 (N_9297,N_9128,N_9215);
or U9298 (N_9298,N_9247,N_9189);
nor U9299 (N_9299,N_9144,N_9142);
nand U9300 (N_9300,N_9193,N_9212);
nor U9301 (N_9301,N_9154,N_9172);
nand U9302 (N_9302,N_9162,N_9165);
and U9303 (N_9303,N_9186,N_9210);
or U9304 (N_9304,N_9126,N_9242);
nor U9305 (N_9305,N_9175,N_9240);
or U9306 (N_9306,N_9190,N_9232);
and U9307 (N_9307,N_9244,N_9167);
and U9308 (N_9308,N_9248,N_9234);
xor U9309 (N_9309,N_9196,N_9130);
or U9310 (N_9310,N_9239,N_9147);
nand U9311 (N_9311,N_9222,N_9181);
or U9312 (N_9312,N_9238,N_9246);
xnor U9313 (N_9313,N_9203,N_9142);
nand U9314 (N_9314,N_9165,N_9227);
or U9315 (N_9315,N_9201,N_9226);
or U9316 (N_9316,N_9151,N_9198);
nand U9317 (N_9317,N_9182,N_9170);
nand U9318 (N_9318,N_9217,N_9172);
nor U9319 (N_9319,N_9199,N_9150);
nand U9320 (N_9320,N_9167,N_9191);
and U9321 (N_9321,N_9129,N_9240);
xor U9322 (N_9322,N_9164,N_9134);
or U9323 (N_9323,N_9220,N_9176);
xnor U9324 (N_9324,N_9127,N_9172);
and U9325 (N_9325,N_9152,N_9201);
and U9326 (N_9326,N_9203,N_9198);
xnor U9327 (N_9327,N_9136,N_9211);
nor U9328 (N_9328,N_9177,N_9219);
or U9329 (N_9329,N_9244,N_9218);
nor U9330 (N_9330,N_9211,N_9244);
or U9331 (N_9331,N_9187,N_9166);
nand U9332 (N_9332,N_9171,N_9218);
nand U9333 (N_9333,N_9219,N_9245);
nand U9334 (N_9334,N_9159,N_9169);
nand U9335 (N_9335,N_9205,N_9224);
xor U9336 (N_9336,N_9236,N_9227);
and U9337 (N_9337,N_9179,N_9140);
xnor U9338 (N_9338,N_9156,N_9147);
or U9339 (N_9339,N_9167,N_9208);
xnor U9340 (N_9340,N_9236,N_9161);
nor U9341 (N_9341,N_9230,N_9231);
nor U9342 (N_9342,N_9199,N_9196);
and U9343 (N_9343,N_9182,N_9201);
and U9344 (N_9344,N_9221,N_9176);
and U9345 (N_9345,N_9176,N_9184);
nor U9346 (N_9346,N_9128,N_9135);
xor U9347 (N_9347,N_9225,N_9243);
or U9348 (N_9348,N_9188,N_9140);
nor U9349 (N_9349,N_9197,N_9205);
and U9350 (N_9350,N_9147,N_9187);
nand U9351 (N_9351,N_9223,N_9144);
nand U9352 (N_9352,N_9206,N_9173);
nand U9353 (N_9353,N_9195,N_9139);
nor U9354 (N_9354,N_9165,N_9243);
nand U9355 (N_9355,N_9137,N_9176);
nor U9356 (N_9356,N_9162,N_9191);
nand U9357 (N_9357,N_9176,N_9192);
or U9358 (N_9358,N_9167,N_9234);
nand U9359 (N_9359,N_9128,N_9248);
xnor U9360 (N_9360,N_9183,N_9165);
nor U9361 (N_9361,N_9173,N_9169);
xor U9362 (N_9362,N_9162,N_9177);
and U9363 (N_9363,N_9143,N_9248);
and U9364 (N_9364,N_9214,N_9241);
and U9365 (N_9365,N_9249,N_9244);
xor U9366 (N_9366,N_9191,N_9161);
xnor U9367 (N_9367,N_9176,N_9150);
nor U9368 (N_9368,N_9136,N_9223);
nor U9369 (N_9369,N_9168,N_9183);
nand U9370 (N_9370,N_9127,N_9213);
nor U9371 (N_9371,N_9167,N_9142);
and U9372 (N_9372,N_9178,N_9155);
and U9373 (N_9373,N_9139,N_9188);
nand U9374 (N_9374,N_9231,N_9188);
nor U9375 (N_9375,N_9323,N_9335);
xnor U9376 (N_9376,N_9266,N_9307);
or U9377 (N_9377,N_9352,N_9334);
and U9378 (N_9378,N_9324,N_9288);
nand U9379 (N_9379,N_9330,N_9259);
nor U9380 (N_9380,N_9341,N_9267);
and U9381 (N_9381,N_9325,N_9332);
or U9382 (N_9382,N_9304,N_9361);
and U9383 (N_9383,N_9253,N_9310);
or U9384 (N_9384,N_9260,N_9254);
nand U9385 (N_9385,N_9311,N_9263);
nor U9386 (N_9386,N_9280,N_9312);
and U9387 (N_9387,N_9316,N_9251);
xnor U9388 (N_9388,N_9358,N_9274);
and U9389 (N_9389,N_9337,N_9363);
and U9390 (N_9390,N_9327,N_9355);
or U9391 (N_9391,N_9372,N_9296);
nand U9392 (N_9392,N_9279,N_9318);
or U9393 (N_9393,N_9293,N_9356);
or U9394 (N_9394,N_9328,N_9272);
nand U9395 (N_9395,N_9373,N_9309);
and U9396 (N_9396,N_9333,N_9290);
nor U9397 (N_9397,N_9344,N_9357);
xor U9398 (N_9398,N_9322,N_9367);
nor U9399 (N_9399,N_9340,N_9273);
and U9400 (N_9400,N_9353,N_9368);
nand U9401 (N_9401,N_9350,N_9300);
xor U9402 (N_9402,N_9314,N_9317);
nand U9403 (N_9403,N_9285,N_9366);
nor U9404 (N_9404,N_9264,N_9281);
xnor U9405 (N_9405,N_9354,N_9329);
xor U9406 (N_9406,N_9269,N_9345);
nand U9407 (N_9407,N_9287,N_9255);
nor U9408 (N_9408,N_9326,N_9284);
nor U9409 (N_9409,N_9364,N_9261);
and U9410 (N_9410,N_9374,N_9362);
and U9411 (N_9411,N_9338,N_9351);
and U9412 (N_9412,N_9292,N_9250);
and U9413 (N_9413,N_9301,N_9305);
nor U9414 (N_9414,N_9265,N_9278);
xor U9415 (N_9415,N_9365,N_9319);
xor U9416 (N_9416,N_9331,N_9313);
xor U9417 (N_9417,N_9321,N_9282);
xor U9418 (N_9418,N_9298,N_9262);
nor U9419 (N_9419,N_9342,N_9346);
nor U9420 (N_9420,N_9315,N_9303);
nand U9421 (N_9421,N_9252,N_9348);
nor U9422 (N_9422,N_9320,N_9297);
or U9423 (N_9423,N_9359,N_9294);
or U9424 (N_9424,N_9295,N_9257);
nor U9425 (N_9425,N_9339,N_9349);
nand U9426 (N_9426,N_9291,N_9271);
nand U9427 (N_9427,N_9270,N_9286);
nor U9428 (N_9428,N_9289,N_9371);
xnor U9429 (N_9429,N_9299,N_9283);
or U9430 (N_9430,N_9369,N_9360);
xor U9431 (N_9431,N_9268,N_9277);
or U9432 (N_9432,N_9308,N_9343);
or U9433 (N_9433,N_9347,N_9370);
and U9434 (N_9434,N_9256,N_9306);
and U9435 (N_9435,N_9275,N_9302);
xnor U9436 (N_9436,N_9336,N_9258);
nand U9437 (N_9437,N_9276,N_9322);
nor U9438 (N_9438,N_9283,N_9351);
and U9439 (N_9439,N_9263,N_9327);
and U9440 (N_9440,N_9327,N_9305);
xnor U9441 (N_9441,N_9310,N_9305);
and U9442 (N_9442,N_9345,N_9295);
xor U9443 (N_9443,N_9306,N_9254);
or U9444 (N_9444,N_9268,N_9348);
xnor U9445 (N_9445,N_9254,N_9316);
nor U9446 (N_9446,N_9352,N_9366);
nor U9447 (N_9447,N_9317,N_9253);
xnor U9448 (N_9448,N_9322,N_9252);
xnor U9449 (N_9449,N_9346,N_9313);
or U9450 (N_9450,N_9254,N_9265);
xnor U9451 (N_9451,N_9302,N_9254);
nand U9452 (N_9452,N_9305,N_9341);
nor U9453 (N_9453,N_9322,N_9259);
or U9454 (N_9454,N_9300,N_9361);
and U9455 (N_9455,N_9316,N_9260);
xnor U9456 (N_9456,N_9296,N_9282);
xor U9457 (N_9457,N_9308,N_9332);
or U9458 (N_9458,N_9322,N_9258);
xnor U9459 (N_9459,N_9267,N_9365);
and U9460 (N_9460,N_9329,N_9326);
xnor U9461 (N_9461,N_9349,N_9326);
xnor U9462 (N_9462,N_9292,N_9270);
or U9463 (N_9463,N_9358,N_9365);
and U9464 (N_9464,N_9292,N_9307);
xor U9465 (N_9465,N_9301,N_9316);
xnor U9466 (N_9466,N_9275,N_9344);
nor U9467 (N_9467,N_9329,N_9318);
or U9468 (N_9468,N_9372,N_9257);
nand U9469 (N_9469,N_9337,N_9292);
nor U9470 (N_9470,N_9303,N_9352);
or U9471 (N_9471,N_9359,N_9271);
nor U9472 (N_9472,N_9279,N_9257);
nand U9473 (N_9473,N_9265,N_9292);
and U9474 (N_9474,N_9314,N_9343);
nand U9475 (N_9475,N_9331,N_9337);
xor U9476 (N_9476,N_9282,N_9257);
and U9477 (N_9477,N_9306,N_9274);
xnor U9478 (N_9478,N_9311,N_9257);
and U9479 (N_9479,N_9284,N_9270);
xnor U9480 (N_9480,N_9309,N_9278);
nor U9481 (N_9481,N_9363,N_9345);
and U9482 (N_9482,N_9293,N_9255);
xnor U9483 (N_9483,N_9308,N_9323);
nor U9484 (N_9484,N_9287,N_9365);
nor U9485 (N_9485,N_9373,N_9270);
xor U9486 (N_9486,N_9258,N_9271);
xor U9487 (N_9487,N_9324,N_9333);
xor U9488 (N_9488,N_9374,N_9292);
and U9489 (N_9489,N_9353,N_9322);
or U9490 (N_9490,N_9291,N_9361);
or U9491 (N_9491,N_9302,N_9323);
or U9492 (N_9492,N_9310,N_9250);
and U9493 (N_9493,N_9361,N_9255);
nor U9494 (N_9494,N_9278,N_9345);
xor U9495 (N_9495,N_9255,N_9312);
and U9496 (N_9496,N_9361,N_9349);
nand U9497 (N_9497,N_9359,N_9285);
nand U9498 (N_9498,N_9373,N_9342);
and U9499 (N_9499,N_9280,N_9273);
xor U9500 (N_9500,N_9423,N_9444);
and U9501 (N_9501,N_9436,N_9419);
xnor U9502 (N_9502,N_9461,N_9386);
or U9503 (N_9503,N_9403,N_9466);
or U9504 (N_9504,N_9431,N_9383);
xor U9505 (N_9505,N_9389,N_9434);
nand U9506 (N_9506,N_9428,N_9472);
xnor U9507 (N_9507,N_9498,N_9381);
xor U9508 (N_9508,N_9410,N_9464);
or U9509 (N_9509,N_9407,N_9479);
xor U9510 (N_9510,N_9457,N_9379);
nand U9511 (N_9511,N_9455,N_9451);
nand U9512 (N_9512,N_9405,N_9391);
or U9513 (N_9513,N_9433,N_9401);
nand U9514 (N_9514,N_9487,N_9453);
nand U9515 (N_9515,N_9430,N_9474);
xnor U9516 (N_9516,N_9409,N_9490);
nor U9517 (N_9517,N_9499,N_9488);
and U9518 (N_9518,N_9469,N_9412);
and U9519 (N_9519,N_9489,N_9415);
or U9520 (N_9520,N_9395,N_9492);
nor U9521 (N_9521,N_9429,N_9473);
nor U9522 (N_9522,N_9413,N_9422);
and U9523 (N_9523,N_9446,N_9493);
or U9524 (N_9524,N_9426,N_9445);
or U9525 (N_9525,N_9432,N_9380);
nor U9526 (N_9526,N_9404,N_9462);
or U9527 (N_9527,N_9396,N_9458);
nand U9528 (N_9528,N_9399,N_9424);
or U9529 (N_9529,N_9437,N_9478);
or U9530 (N_9530,N_9497,N_9463);
nor U9531 (N_9531,N_9385,N_9483);
or U9532 (N_9532,N_9420,N_9481);
nor U9533 (N_9533,N_9495,N_9452);
and U9534 (N_9534,N_9475,N_9476);
xnor U9535 (N_9535,N_9416,N_9454);
xnor U9536 (N_9536,N_9491,N_9480);
nand U9537 (N_9537,N_9467,N_9450);
or U9538 (N_9538,N_9397,N_9414);
and U9539 (N_9539,N_9384,N_9443);
nor U9540 (N_9540,N_9494,N_9402);
or U9541 (N_9541,N_9418,N_9390);
and U9542 (N_9542,N_9400,N_9435);
or U9543 (N_9543,N_9411,N_9387);
and U9544 (N_9544,N_9459,N_9392);
xnor U9545 (N_9545,N_9496,N_9447);
nor U9546 (N_9546,N_9442,N_9408);
nand U9547 (N_9547,N_9421,N_9375);
or U9548 (N_9548,N_9449,N_9427);
or U9549 (N_9549,N_9440,N_9382);
and U9550 (N_9550,N_9394,N_9468);
or U9551 (N_9551,N_9377,N_9441);
nand U9552 (N_9552,N_9485,N_9388);
and U9553 (N_9553,N_9484,N_9471);
nand U9554 (N_9554,N_9439,N_9456);
nand U9555 (N_9555,N_9438,N_9406);
nand U9556 (N_9556,N_9482,N_9376);
or U9557 (N_9557,N_9477,N_9398);
and U9558 (N_9558,N_9417,N_9465);
nor U9559 (N_9559,N_9378,N_9448);
nand U9560 (N_9560,N_9393,N_9460);
and U9561 (N_9561,N_9486,N_9470);
xor U9562 (N_9562,N_9425,N_9480);
or U9563 (N_9563,N_9439,N_9482);
and U9564 (N_9564,N_9394,N_9474);
nand U9565 (N_9565,N_9440,N_9456);
and U9566 (N_9566,N_9449,N_9472);
nand U9567 (N_9567,N_9435,N_9378);
or U9568 (N_9568,N_9469,N_9456);
xnor U9569 (N_9569,N_9439,N_9498);
nor U9570 (N_9570,N_9492,N_9481);
nand U9571 (N_9571,N_9407,N_9452);
xnor U9572 (N_9572,N_9405,N_9432);
xnor U9573 (N_9573,N_9490,N_9381);
nor U9574 (N_9574,N_9446,N_9442);
xnor U9575 (N_9575,N_9461,N_9403);
or U9576 (N_9576,N_9440,N_9393);
and U9577 (N_9577,N_9381,N_9429);
or U9578 (N_9578,N_9390,N_9492);
nor U9579 (N_9579,N_9441,N_9482);
or U9580 (N_9580,N_9410,N_9379);
xnor U9581 (N_9581,N_9422,N_9433);
nand U9582 (N_9582,N_9397,N_9419);
xor U9583 (N_9583,N_9471,N_9478);
nor U9584 (N_9584,N_9450,N_9443);
and U9585 (N_9585,N_9458,N_9376);
or U9586 (N_9586,N_9490,N_9398);
or U9587 (N_9587,N_9414,N_9375);
xor U9588 (N_9588,N_9440,N_9471);
or U9589 (N_9589,N_9454,N_9463);
or U9590 (N_9590,N_9497,N_9432);
and U9591 (N_9591,N_9458,N_9489);
nor U9592 (N_9592,N_9472,N_9441);
xor U9593 (N_9593,N_9381,N_9400);
or U9594 (N_9594,N_9446,N_9400);
nand U9595 (N_9595,N_9397,N_9398);
nor U9596 (N_9596,N_9377,N_9434);
nand U9597 (N_9597,N_9386,N_9464);
or U9598 (N_9598,N_9383,N_9385);
or U9599 (N_9599,N_9480,N_9431);
xnor U9600 (N_9600,N_9482,N_9397);
or U9601 (N_9601,N_9478,N_9392);
nand U9602 (N_9602,N_9424,N_9434);
nor U9603 (N_9603,N_9476,N_9458);
or U9604 (N_9604,N_9463,N_9428);
nor U9605 (N_9605,N_9455,N_9379);
nor U9606 (N_9606,N_9469,N_9391);
or U9607 (N_9607,N_9442,N_9452);
or U9608 (N_9608,N_9403,N_9415);
xor U9609 (N_9609,N_9443,N_9389);
nor U9610 (N_9610,N_9467,N_9384);
nor U9611 (N_9611,N_9496,N_9470);
nor U9612 (N_9612,N_9420,N_9498);
or U9613 (N_9613,N_9478,N_9428);
nor U9614 (N_9614,N_9473,N_9407);
xnor U9615 (N_9615,N_9394,N_9441);
nor U9616 (N_9616,N_9422,N_9401);
and U9617 (N_9617,N_9450,N_9463);
nor U9618 (N_9618,N_9384,N_9482);
nor U9619 (N_9619,N_9392,N_9476);
xor U9620 (N_9620,N_9453,N_9431);
nor U9621 (N_9621,N_9472,N_9491);
and U9622 (N_9622,N_9414,N_9411);
nor U9623 (N_9623,N_9378,N_9496);
nand U9624 (N_9624,N_9377,N_9451);
or U9625 (N_9625,N_9532,N_9504);
nand U9626 (N_9626,N_9554,N_9593);
or U9627 (N_9627,N_9542,N_9530);
xor U9628 (N_9628,N_9565,N_9506);
xnor U9629 (N_9629,N_9575,N_9527);
nor U9630 (N_9630,N_9524,N_9590);
xor U9631 (N_9631,N_9514,N_9573);
and U9632 (N_9632,N_9520,N_9548);
nand U9633 (N_9633,N_9586,N_9539);
and U9634 (N_9634,N_9518,N_9513);
xor U9635 (N_9635,N_9580,N_9563);
xor U9636 (N_9636,N_9555,N_9510);
nand U9637 (N_9637,N_9531,N_9574);
or U9638 (N_9638,N_9536,N_9569);
or U9639 (N_9639,N_9547,N_9596);
or U9640 (N_9640,N_9624,N_9576);
and U9641 (N_9641,N_9585,N_9578);
nor U9642 (N_9642,N_9552,N_9617);
and U9643 (N_9643,N_9606,N_9529);
or U9644 (N_9644,N_9605,N_9560);
or U9645 (N_9645,N_9526,N_9544);
or U9646 (N_9646,N_9561,N_9602);
or U9647 (N_9647,N_9621,N_9600);
nor U9648 (N_9648,N_9533,N_9604);
and U9649 (N_9649,N_9577,N_9540);
nor U9650 (N_9650,N_9595,N_9522);
xor U9651 (N_9651,N_9584,N_9556);
and U9652 (N_9652,N_9538,N_9587);
xor U9653 (N_9653,N_9505,N_9521);
xnor U9654 (N_9654,N_9559,N_9568);
nor U9655 (N_9655,N_9551,N_9610);
or U9656 (N_9656,N_9594,N_9616);
nor U9657 (N_9657,N_9528,N_9541);
and U9658 (N_9658,N_9589,N_9515);
and U9659 (N_9659,N_9588,N_9564);
xor U9660 (N_9660,N_9558,N_9549);
nand U9661 (N_9661,N_9612,N_9566);
nand U9662 (N_9662,N_9598,N_9597);
nand U9663 (N_9663,N_9562,N_9572);
and U9664 (N_9664,N_9511,N_9546);
xnor U9665 (N_9665,N_9517,N_9500);
and U9666 (N_9666,N_9516,N_9623);
and U9667 (N_9667,N_9557,N_9545);
or U9668 (N_9668,N_9618,N_9535);
xnor U9669 (N_9669,N_9608,N_9534);
nor U9670 (N_9670,N_9512,N_9603);
xor U9671 (N_9671,N_9503,N_9609);
and U9672 (N_9672,N_9611,N_9622);
and U9673 (N_9673,N_9592,N_9550);
nor U9674 (N_9674,N_9583,N_9508);
xor U9675 (N_9675,N_9525,N_9537);
nor U9676 (N_9676,N_9571,N_9570);
nor U9677 (N_9677,N_9553,N_9509);
xnor U9678 (N_9678,N_9615,N_9599);
nand U9679 (N_9679,N_9581,N_9543);
nand U9680 (N_9680,N_9567,N_9607);
nand U9681 (N_9681,N_9620,N_9523);
nand U9682 (N_9682,N_9501,N_9613);
nor U9683 (N_9683,N_9579,N_9619);
and U9684 (N_9684,N_9519,N_9614);
nand U9685 (N_9685,N_9601,N_9582);
and U9686 (N_9686,N_9507,N_9502);
nand U9687 (N_9687,N_9591,N_9553);
nor U9688 (N_9688,N_9518,N_9550);
nand U9689 (N_9689,N_9524,N_9556);
nor U9690 (N_9690,N_9504,N_9522);
or U9691 (N_9691,N_9533,N_9583);
nor U9692 (N_9692,N_9595,N_9509);
nand U9693 (N_9693,N_9622,N_9522);
nand U9694 (N_9694,N_9590,N_9609);
nand U9695 (N_9695,N_9549,N_9520);
nor U9696 (N_9696,N_9607,N_9577);
and U9697 (N_9697,N_9547,N_9582);
nor U9698 (N_9698,N_9575,N_9577);
nand U9699 (N_9699,N_9544,N_9527);
or U9700 (N_9700,N_9551,N_9546);
or U9701 (N_9701,N_9587,N_9582);
nand U9702 (N_9702,N_9576,N_9597);
and U9703 (N_9703,N_9549,N_9592);
nor U9704 (N_9704,N_9540,N_9617);
nand U9705 (N_9705,N_9581,N_9523);
and U9706 (N_9706,N_9574,N_9507);
and U9707 (N_9707,N_9561,N_9624);
xnor U9708 (N_9708,N_9560,N_9607);
xnor U9709 (N_9709,N_9523,N_9529);
and U9710 (N_9710,N_9549,N_9550);
or U9711 (N_9711,N_9576,N_9583);
nand U9712 (N_9712,N_9564,N_9526);
or U9713 (N_9713,N_9504,N_9569);
and U9714 (N_9714,N_9592,N_9598);
nor U9715 (N_9715,N_9605,N_9556);
and U9716 (N_9716,N_9557,N_9515);
nand U9717 (N_9717,N_9514,N_9606);
xor U9718 (N_9718,N_9512,N_9518);
or U9719 (N_9719,N_9545,N_9576);
xor U9720 (N_9720,N_9569,N_9558);
nor U9721 (N_9721,N_9622,N_9569);
and U9722 (N_9722,N_9535,N_9602);
nand U9723 (N_9723,N_9519,N_9588);
and U9724 (N_9724,N_9614,N_9557);
nand U9725 (N_9725,N_9561,N_9570);
nand U9726 (N_9726,N_9545,N_9570);
or U9727 (N_9727,N_9520,N_9624);
xnor U9728 (N_9728,N_9567,N_9622);
and U9729 (N_9729,N_9506,N_9522);
nand U9730 (N_9730,N_9569,N_9554);
xor U9731 (N_9731,N_9565,N_9536);
or U9732 (N_9732,N_9549,N_9532);
nor U9733 (N_9733,N_9536,N_9563);
or U9734 (N_9734,N_9554,N_9564);
or U9735 (N_9735,N_9611,N_9521);
nor U9736 (N_9736,N_9507,N_9515);
nand U9737 (N_9737,N_9569,N_9561);
and U9738 (N_9738,N_9529,N_9518);
or U9739 (N_9739,N_9576,N_9603);
and U9740 (N_9740,N_9503,N_9573);
xnor U9741 (N_9741,N_9570,N_9513);
nor U9742 (N_9742,N_9525,N_9548);
nor U9743 (N_9743,N_9604,N_9565);
or U9744 (N_9744,N_9509,N_9590);
or U9745 (N_9745,N_9613,N_9614);
nand U9746 (N_9746,N_9508,N_9589);
nand U9747 (N_9747,N_9596,N_9541);
or U9748 (N_9748,N_9539,N_9590);
nor U9749 (N_9749,N_9603,N_9594);
xor U9750 (N_9750,N_9732,N_9674);
or U9751 (N_9751,N_9632,N_9630);
nand U9752 (N_9752,N_9639,N_9681);
xnor U9753 (N_9753,N_9678,N_9635);
or U9754 (N_9754,N_9692,N_9683);
xor U9755 (N_9755,N_9707,N_9708);
nor U9756 (N_9756,N_9636,N_9633);
nor U9757 (N_9757,N_9721,N_9628);
nor U9758 (N_9758,N_9655,N_9689);
nor U9759 (N_9759,N_9699,N_9704);
or U9760 (N_9760,N_9631,N_9737);
nor U9761 (N_9761,N_9680,N_9711);
or U9762 (N_9762,N_9706,N_9685);
nand U9763 (N_9763,N_9728,N_9688);
xnor U9764 (N_9764,N_9626,N_9644);
nor U9765 (N_9765,N_9718,N_9649);
nand U9766 (N_9766,N_9642,N_9673);
or U9767 (N_9767,N_9693,N_9726);
and U9768 (N_9768,N_9686,N_9672);
nand U9769 (N_9769,N_9653,N_9691);
nor U9770 (N_9770,N_9666,N_9733);
and U9771 (N_9771,N_9738,N_9729);
and U9772 (N_9772,N_9629,N_9625);
xnor U9773 (N_9773,N_9677,N_9687);
nand U9774 (N_9774,N_9641,N_9743);
and U9775 (N_9775,N_9651,N_9684);
nand U9776 (N_9776,N_9703,N_9722);
xor U9777 (N_9777,N_9665,N_9660);
nor U9778 (N_9778,N_9645,N_9676);
nor U9779 (N_9779,N_9663,N_9745);
nor U9780 (N_9780,N_9670,N_9662);
and U9781 (N_9781,N_9650,N_9696);
nand U9782 (N_9782,N_9739,N_9705);
nor U9783 (N_9783,N_9658,N_9741);
xor U9784 (N_9784,N_9627,N_9664);
and U9785 (N_9785,N_9640,N_9661);
nor U9786 (N_9786,N_9698,N_9734);
or U9787 (N_9787,N_9715,N_9719);
xnor U9788 (N_9788,N_9714,N_9736);
xnor U9789 (N_9789,N_9643,N_9749);
and U9790 (N_9790,N_9700,N_9695);
nand U9791 (N_9791,N_9652,N_9690);
and U9792 (N_9792,N_9735,N_9679);
xor U9793 (N_9793,N_9747,N_9730);
and U9794 (N_9794,N_9748,N_9646);
nand U9795 (N_9795,N_9668,N_9702);
or U9796 (N_9796,N_9710,N_9723);
nand U9797 (N_9797,N_9724,N_9656);
nand U9798 (N_9798,N_9746,N_9694);
nand U9799 (N_9799,N_9654,N_9697);
xor U9800 (N_9800,N_9712,N_9713);
and U9801 (N_9801,N_9727,N_9637);
or U9802 (N_9802,N_9667,N_9648);
nand U9803 (N_9803,N_9709,N_9634);
nor U9804 (N_9804,N_9657,N_9675);
and U9805 (N_9805,N_9638,N_9717);
xor U9806 (N_9806,N_9647,N_9669);
nand U9807 (N_9807,N_9716,N_9742);
nor U9808 (N_9808,N_9740,N_9731);
and U9809 (N_9809,N_9744,N_9720);
xnor U9810 (N_9810,N_9671,N_9682);
nor U9811 (N_9811,N_9725,N_9659);
nand U9812 (N_9812,N_9701,N_9632);
and U9813 (N_9813,N_9720,N_9697);
nor U9814 (N_9814,N_9714,N_9709);
or U9815 (N_9815,N_9737,N_9719);
or U9816 (N_9816,N_9694,N_9731);
and U9817 (N_9817,N_9690,N_9736);
nand U9818 (N_9818,N_9697,N_9684);
or U9819 (N_9819,N_9670,N_9739);
nand U9820 (N_9820,N_9668,N_9709);
xnor U9821 (N_9821,N_9690,N_9724);
and U9822 (N_9822,N_9648,N_9633);
xnor U9823 (N_9823,N_9735,N_9692);
nor U9824 (N_9824,N_9656,N_9723);
and U9825 (N_9825,N_9690,N_9731);
and U9826 (N_9826,N_9690,N_9716);
nand U9827 (N_9827,N_9674,N_9688);
nand U9828 (N_9828,N_9663,N_9671);
nor U9829 (N_9829,N_9704,N_9670);
nand U9830 (N_9830,N_9634,N_9683);
nor U9831 (N_9831,N_9645,N_9716);
and U9832 (N_9832,N_9745,N_9692);
or U9833 (N_9833,N_9652,N_9713);
nor U9834 (N_9834,N_9739,N_9710);
or U9835 (N_9835,N_9632,N_9683);
xor U9836 (N_9836,N_9625,N_9702);
nor U9837 (N_9837,N_9634,N_9640);
nor U9838 (N_9838,N_9745,N_9705);
and U9839 (N_9839,N_9663,N_9682);
nor U9840 (N_9840,N_9703,N_9667);
and U9841 (N_9841,N_9698,N_9697);
or U9842 (N_9842,N_9733,N_9740);
nor U9843 (N_9843,N_9710,N_9667);
xor U9844 (N_9844,N_9721,N_9719);
nor U9845 (N_9845,N_9709,N_9644);
nor U9846 (N_9846,N_9722,N_9641);
nand U9847 (N_9847,N_9711,N_9735);
nand U9848 (N_9848,N_9657,N_9685);
xnor U9849 (N_9849,N_9649,N_9735);
xor U9850 (N_9850,N_9664,N_9659);
and U9851 (N_9851,N_9675,N_9717);
xnor U9852 (N_9852,N_9717,N_9727);
xnor U9853 (N_9853,N_9708,N_9725);
nor U9854 (N_9854,N_9679,N_9626);
nand U9855 (N_9855,N_9666,N_9676);
and U9856 (N_9856,N_9735,N_9654);
nand U9857 (N_9857,N_9669,N_9706);
xor U9858 (N_9858,N_9732,N_9730);
nor U9859 (N_9859,N_9662,N_9720);
or U9860 (N_9860,N_9738,N_9670);
or U9861 (N_9861,N_9630,N_9725);
nor U9862 (N_9862,N_9677,N_9696);
or U9863 (N_9863,N_9660,N_9700);
xnor U9864 (N_9864,N_9725,N_9696);
nand U9865 (N_9865,N_9726,N_9646);
nand U9866 (N_9866,N_9651,N_9668);
xnor U9867 (N_9867,N_9678,N_9660);
xnor U9868 (N_9868,N_9635,N_9703);
nor U9869 (N_9869,N_9718,N_9693);
nor U9870 (N_9870,N_9743,N_9722);
and U9871 (N_9871,N_9742,N_9749);
xor U9872 (N_9872,N_9714,N_9644);
nor U9873 (N_9873,N_9679,N_9682);
nand U9874 (N_9874,N_9703,N_9660);
and U9875 (N_9875,N_9764,N_9815);
nand U9876 (N_9876,N_9759,N_9843);
xor U9877 (N_9877,N_9827,N_9781);
xnor U9878 (N_9878,N_9808,N_9840);
nand U9879 (N_9879,N_9785,N_9850);
nor U9880 (N_9880,N_9812,N_9857);
nand U9881 (N_9881,N_9866,N_9765);
xnor U9882 (N_9882,N_9761,N_9828);
nor U9883 (N_9883,N_9796,N_9845);
xor U9884 (N_9884,N_9835,N_9768);
nand U9885 (N_9885,N_9816,N_9820);
nor U9886 (N_9886,N_9770,N_9822);
nand U9887 (N_9887,N_9831,N_9751);
or U9888 (N_9888,N_9800,N_9826);
nand U9889 (N_9889,N_9758,N_9795);
nor U9890 (N_9890,N_9868,N_9825);
xnor U9891 (N_9891,N_9794,N_9821);
or U9892 (N_9892,N_9771,N_9851);
nor U9893 (N_9893,N_9792,N_9824);
and U9894 (N_9894,N_9756,N_9823);
xor U9895 (N_9895,N_9814,N_9829);
xor U9896 (N_9896,N_9860,N_9766);
or U9897 (N_9897,N_9760,N_9856);
and U9898 (N_9898,N_9769,N_9779);
nor U9899 (N_9899,N_9784,N_9849);
nand U9900 (N_9900,N_9790,N_9807);
nor U9901 (N_9901,N_9797,N_9842);
xor U9902 (N_9902,N_9855,N_9752);
nand U9903 (N_9903,N_9811,N_9788);
and U9904 (N_9904,N_9861,N_9874);
or U9905 (N_9905,N_9848,N_9854);
nand U9906 (N_9906,N_9783,N_9818);
and U9907 (N_9907,N_9750,N_9799);
nor U9908 (N_9908,N_9806,N_9755);
or U9909 (N_9909,N_9753,N_9846);
or U9910 (N_9910,N_9805,N_9803);
and U9911 (N_9911,N_9780,N_9830);
or U9912 (N_9912,N_9804,N_9793);
or U9913 (N_9913,N_9867,N_9869);
xor U9914 (N_9914,N_9772,N_9798);
nor U9915 (N_9915,N_9774,N_9837);
nand U9916 (N_9916,N_9833,N_9844);
or U9917 (N_9917,N_9834,N_9786);
xor U9918 (N_9918,N_9865,N_9832);
or U9919 (N_9919,N_9767,N_9873);
or U9920 (N_9920,N_9757,N_9776);
nor U9921 (N_9921,N_9853,N_9862);
xnor U9922 (N_9922,N_9852,N_9841);
xnor U9923 (N_9923,N_9777,N_9817);
nor U9924 (N_9924,N_9864,N_9819);
or U9925 (N_9925,N_9773,N_9802);
xor U9926 (N_9926,N_9763,N_9789);
xor U9927 (N_9927,N_9838,N_9775);
and U9928 (N_9928,N_9809,N_9871);
and U9929 (N_9929,N_9836,N_9754);
and U9930 (N_9930,N_9858,N_9782);
nand U9931 (N_9931,N_9778,N_9859);
nand U9932 (N_9932,N_9762,N_9810);
xnor U9933 (N_9933,N_9801,N_9872);
and U9934 (N_9934,N_9787,N_9813);
nor U9935 (N_9935,N_9847,N_9870);
nor U9936 (N_9936,N_9791,N_9863);
nand U9937 (N_9937,N_9839,N_9780);
nor U9938 (N_9938,N_9760,N_9843);
and U9939 (N_9939,N_9778,N_9842);
xnor U9940 (N_9940,N_9831,N_9864);
nand U9941 (N_9941,N_9823,N_9866);
and U9942 (N_9942,N_9796,N_9753);
xnor U9943 (N_9943,N_9789,N_9761);
xnor U9944 (N_9944,N_9752,N_9767);
or U9945 (N_9945,N_9858,N_9797);
and U9946 (N_9946,N_9833,N_9766);
nor U9947 (N_9947,N_9841,N_9785);
nand U9948 (N_9948,N_9785,N_9778);
xor U9949 (N_9949,N_9843,N_9854);
nor U9950 (N_9950,N_9774,N_9825);
and U9951 (N_9951,N_9818,N_9803);
and U9952 (N_9952,N_9842,N_9802);
or U9953 (N_9953,N_9850,N_9796);
xnor U9954 (N_9954,N_9751,N_9841);
and U9955 (N_9955,N_9829,N_9802);
xor U9956 (N_9956,N_9759,N_9790);
or U9957 (N_9957,N_9856,N_9781);
xnor U9958 (N_9958,N_9801,N_9842);
or U9959 (N_9959,N_9811,N_9808);
nand U9960 (N_9960,N_9773,N_9818);
or U9961 (N_9961,N_9807,N_9778);
and U9962 (N_9962,N_9863,N_9847);
or U9963 (N_9963,N_9772,N_9822);
nor U9964 (N_9964,N_9832,N_9873);
nand U9965 (N_9965,N_9840,N_9796);
and U9966 (N_9966,N_9761,N_9826);
xor U9967 (N_9967,N_9759,N_9802);
nand U9968 (N_9968,N_9800,N_9806);
or U9969 (N_9969,N_9809,N_9814);
and U9970 (N_9970,N_9773,N_9850);
and U9971 (N_9971,N_9863,N_9796);
or U9972 (N_9972,N_9782,N_9785);
and U9973 (N_9973,N_9857,N_9865);
and U9974 (N_9974,N_9817,N_9844);
and U9975 (N_9975,N_9825,N_9787);
or U9976 (N_9976,N_9791,N_9838);
or U9977 (N_9977,N_9874,N_9838);
xor U9978 (N_9978,N_9808,N_9825);
xor U9979 (N_9979,N_9865,N_9826);
and U9980 (N_9980,N_9826,N_9828);
nor U9981 (N_9981,N_9810,N_9757);
and U9982 (N_9982,N_9827,N_9856);
xnor U9983 (N_9983,N_9839,N_9762);
nor U9984 (N_9984,N_9785,N_9801);
or U9985 (N_9985,N_9811,N_9784);
xnor U9986 (N_9986,N_9803,N_9864);
or U9987 (N_9987,N_9834,N_9803);
xor U9988 (N_9988,N_9764,N_9874);
nor U9989 (N_9989,N_9807,N_9751);
xnor U9990 (N_9990,N_9810,N_9839);
or U9991 (N_9991,N_9824,N_9810);
nor U9992 (N_9992,N_9850,N_9782);
nor U9993 (N_9993,N_9822,N_9774);
nand U9994 (N_9994,N_9831,N_9856);
and U9995 (N_9995,N_9826,N_9789);
nand U9996 (N_9996,N_9785,N_9802);
or U9997 (N_9997,N_9874,N_9871);
nand U9998 (N_9998,N_9795,N_9828);
nor U9999 (N_9999,N_9787,N_9768);
nand U10000 (N_10000,N_9972,N_9968);
xnor U10001 (N_10001,N_9938,N_9886);
and U10002 (N_10002,N_9911,N_9945);
nor U10003 (N_10003,N_9957,N_9932);
xnor U10004 (N_10004,N_9964,N_9979);
xor U10005 (N_10005,N_9902,N_9885);
nor U10006 (N_10006,N_9915,N_9966);
nand U10007 (N_10007,N_9930,N_9990);
xnor U10008 (N_10008,N_9933,N_9934);
and U10009 (N_10009,N_9876,N_9931);
nor U10010 (N_10010,N_9887,N_9892);
nor U10011 (N_10011,N_9884,N_9924);
or U10012 (N_10012,N_9927,N_9914);
or U10013 (N_10013,N_9950,N_9993);
nor U10014 (N_10014,N_9916,N_9881);
or U10015 (N_10015,N_9973,N_9896);
and U10016 (N_10016,N_9978,N_9910);
nor U10017 (N_10017,N_9956,N_9918);
nand U10018 (N_10018,N_9937,N_9878);
and U10019 (N_10019,N_9941,N_9909);
or U10020 (N_10020,N_9974,N_9913);
xnor U10021 (N_10021,N_9948,N_9997);
nor U10022 (N_10022,N_9904,N_9893);
or U10023 (N_10023,N_9894,N_9880);
and U10024 (N_10024,N_9875,N_9944);
xnor U10025 (N_10025,N_9994,N_9983);
and U10026 (N_10026,N_9883,N_9991);
xnor U10027 (N_10027,N_9903,N_9960);
nor U10028 (N_10028,N_9925,N_9981);
and U10029 (N_10029,N_9985,N_9949);
nor U10030 (N_10030,N_9926,N_9908);
xor U10031 (N_10031,N_9940,N_9921);
nand U10032 (N_10032,N_9900,N_9998);
nand U10033 (N_10033,N_9970,N_9889);
nor U10034 (N_10034,N_9890,N_9917);
nor U10035 (N_10035,N_9897,N_9953);
and U10036 (N_10036,N_9967,N_9954);
or U10037 (N_10037,N_9986,N_9906);
and U10038 (N_10038,N_9971,N_9992);
nor U10039 (N_10039,N_9959,N_9958);
nor U10040 (N_10040,N_9895,N_9987);
nand U10041 (N_10041,N_9984,N_9962);
or U10042 (N_10042,N_9996,N_9882);
or U10043 (N_10043,N_9888,N_9988);
nand U10044 (N_10044,N_9901,N_9939);
xor U10045 (N_10045,N_9989,N_9923);
nand U10046 (N_10046,N_9995,N_9929);
or U10047 (N_10047,N_9922,N_9963);
nor U10048 (N_10048,N_9877,N_9977);
nand U10049 (N_10049,N_9946,N_9912);
nand U10050 (N_10050,N_9980,N_9936);
or U10051 (N_10051,N_9920,N_9975);
nor U10052 (N_10052,N_9976,N_9943);
or U10053 (N_10053,N_9919,N_9947);
xnor U10054 (N_10054,N_9935,N_9965);
and U10055 (N_10055,N_9999,N_9982);
nand U10056 (N_10056,N_9907,N_9879);
or U10057 (N_10057,N_9899,N_9955);
or U10058 (N_10058,N_9942,N_9905);
nor U10059 (N_10059,N_9891,N_9928);
xnor U10060 (N_10060,N_9898,N_9952);
nand U10061 (N_10061,N_9969,N_9951);
or U10062 (N_10062,N_9961,N_9908);
xor U10063 (N_10063,N_9920,N_9999);
or U10064 (N_10064,N_9995,N_9958);
xor U10065 (N_10065,N_9967,N_9918);
nand U10066 (N_10066,N_9940,N_9961);
xor U10067 (N_10067,N_9931,N_9963);
or U10068 (N_10068,N_9965,N_9885);
and U10069 (N_10069,N_9912,N_9949);
nor U10070 (N_10070,N_9943,N_9964);
nor U10071 (N_10071,N_9899,N_9997);
or U10072 (N_10072,N_9946,N_9952);
nand U10073 (N_10073,N_9887,N_9878);
nand U10074 (N_10074,N_9974,N_9956);
xor U10075 (N_10075,N_9920,N_9892);
and U10076 (N_10076,N_9898,N_9939);
nand U10077 (N_10077,N_9961,N_9914);
or U10078 (N_10078,N_9994,N_9884);
and U10079 (N_10079,N_9921,N_9902);
and U10080 (N_10080,N_9990,N_9986);
and U10081 (N_10081,N_9882,N_9876);
nor U10082 (N_10082,N_9947,N_9909);
nor U10083 (N_10083,N_9979,N_9928);
and U10084 (N_10084,N_9965,N_9943);
nor U10085 (N_10085,N_9917,N_9883);
nor U10086 (N_10086,N_9982,N_9941);
or U10087 (N_10087,N_9987,N_9920);
nor U10088 (N_10088,N_9988,N_9926);
and U10089 (N_10089,N_9985,N_9945);
xnor U10090 (N_10090,N_9879,N_9987);
nor U10091 (N_10091,N_9990,N_9981);
xor U10092 (N_10092,N_9897,N_9949);
and U10093 (N_10093,N_9912,N_9950);
and U10094 (N_10094,N_9944,N_9983);
or U10095 (N_10095,N_9968,N_9992);
or U10096 (N_10096,N_9969,N_9954);
and U10097 (N_10097,N_9967,N_9924);
or U10098 (N_10098,N_9977,N_9966);
and U10099 (N_10099,N_9981,N_9985);
nand U10100 (N_10100,N_9906,N_9879);
nor U10101 (N_10101,N_9962,N_9990);
nor U10102 (N_10102,N_9939,N_9962);
or U10103 (N_10103,N_9903,N_9882);
or U10104 (N_10104,N_9923,N_9927);
nor U10105 (N_10105,N_9995,N_9997);
or U10106 (N_10106,N_9936,N_9934);
nand U10107 (N_10107,N_9943,N_9957);
nor U10108 (N_10108,N_9963,N_9993);
and U10109 (N_10109,N_9912,N_9906);
or U10110 (N_10110,N_9948,N_9920);
or U10111 (N_10111,N_9915,N_9918);
and U10112 (N_10112,N_9949,N_9997);
and U10113 (N_10113,N_9887,N_9953);
nand U10114 (N_10114,N_9909,N_9893);
and U10115 (N_10115,N_9932,N_9921);
and U10116 (N_10116,N_9882,N_9922);
or U10117 (N_10117,N_9955,N_9916);
nor U10118 (N_10118,N_9886,N_9931);
nor U10119 (N_10119,N_9919,N_9896);
xnor U10120 (N_10120,N_9907,N_9986);
xor U10121 (N_10121,N_9960,N_9952);
nand U10122 (N_10122,N_9982,N_9890);
nor U10123 (N_10123,N_9943,N_9961);
nand U10124 (N_10124,N_9881,N_9968);
nor U10125 (N_10125,N_10113,N_10011);
xor U10126 (N_10126,N_10103,N_10039);
nand U10127 (N_10127,N_10042,N_10120);
or U10128 (N_10128,N_10025,N_10014);
nor U10129 (N_10129,N_10062,N_10087);
nor U10130 (N_10130,N_10076,N_10102);
and U10131 (N_10131,N_10070,N_10089);
xor U10132 (N_10132,N_10015,N_10035);
and U10133 (N_10133,N_10110,N_10114);
xor U10134 (N_10134,N_10020,N_10098);
xor U10135 (N_10135,N_10115,N_10073);
xor U10136 (N_10136,N_10041,N_10032);
nor U10137 (N_10137,N_10107,N_10085);
and U10138 (N_10138,N_10104,N_10082);
and U10139 (N_10139,N_10094,N_10066);
nand U10140 (N_10140,N_10021,N_10119);
or U10141 (N_10141,N_10096,N_10034);
nand U10142 (N_10142,N_10024,N_10095);
xor U10143 (N_10143,N_10101,N_10077);
or U10144 (N_10144,N_10050,N_10083);
nor U10145 (N_10145,N_10013,N_10045);
nor U10146 (N_10146,N_10047,N_10078);
and U10147 (N_10147,N_10057,N_10022);
nand U10148 (N_10148,N_10090,N_10012);
xor U10149 (N_10149,N_10002,N_10112);
and U10150 (N_10150,N_10040,N_10067);
or U10151 (N_10151,N_10008,N_10064);
and U10152 (N_10152,N_10023,N_10004);
nor U10153 (N_10153,N_10111,N_10093);
and U10154 (N_10154,N_10063,N_10086);
nand U10155 (N_10155,N_10124,N_10118);
nand U10156 (N_10156,N_10030,N_10006);
and U10157 (N_10157,N_10065,N_10044);
xor U10158 (N_10158,N_10049,N_10007);
or U10159 (N_10159,N_10097,N_10088);
or U10160 (N_10160,N_10068,N_10009);
xnor U10161 (N_10161,N_10003,N_10038);
and U10162 (N_10162,N_10080,N_10059);
xor U10163 (N_10163,N_10033,N_10046);
or U10164 (N_10164,N_10075,N_10109);
nand U10165 (N_10165,N_10051,N_10048);
or U10166 (N_10166,N_10117,N_10121);
xnor U10167 (N_10167,N_10026,N_10036);
nand U10168 (N_10168,N_10079,N_10005);
nand U10169 (N_10169,N_10074,N_10056);
and U10170 (N_10170,N_10123,N_10092);
or U10171 (N_10171,N_10071,N_10099);
nor U10172 (N_10172,N_10105,N_10060);
or U10173 (N_10173,N_10018,N_10031);
nand U10174 (N_10174,N_10072,N_10027);
nor U10175 (N_10175,N_10016,N_10084);
nand U10176 (N_10176,N_10058,N_10061);
xor U10177 (N_10177,N_10069,N_10106);
nand U10178 (N_10178,N_10122,N_10001);
or U10179 (N_10179,N_10000,N_10010);
or U10180 (N_10180,N_10028,N_10054);
nand U10181 (N_10181,N_10100,N_10017);
xnor U10182 (N_10182,N_10091,N_10052);
or U10183 (N_10183,N_10029,N_10019);
and U10184 (N_10184,N_10055,N_10108);
or U10185 (N_10185,N_10053,N_10116);
nand U10186 (N_10186,N_10037,N_10081);
xnor U10187 (N_10187,N_10043,N_10017);
nor U10188 (N_10188,N_10062,N_10033);
or U10189 (N_10189,N_10063,N_10118);
nand U10190 (N_10190,N_10017,N_10093);
and U10191 (N_10191,N_10066,N_10036);
xnor U10192 (N_10192,N_10026,N_10114);
or U10193 (N_10193,N_10119,N_10074);
and U10194 (N_10194,N_10124,N_10032);
nor U10195 (N_10195,N_10092,N_10073);
and U10196 (N_10196,N_10011,N_10087);
xor U10197 (N_10197,N_10040,N_10088);
xor U10198 (N_10198,N_10055,N_10008);
xor U10199 (N_10199,N_10089,N_10097);
nand U10200 (N_10200,N_10033,N_10115);
nand U10201 (N_10201,N_10012,N_10119);
xnor U10202 (N_10202,N_10086,N_10041);
xor U10203 (N_10203,N_10004,N_10040);
nand U10204 (N_10204,N_10095,N_10109);
nand U10205 (N_10205,N_10116,N_10079);
nor U10206 (N_10206,N_10019,N_10097);
xor U10207 (N_10207,N_10049,N_10026);
nand U10208 (N_10208,N_10007,N_10011);
nor U10209 (N_10209,N_10019,N_10049);
or U10210 (N_10210,N_10066,N_10097);
nand U10211 (N_10211,N_10086,N_10045);
nor U10212 (N_10212,N_10048,N_10096);
xnor U10213 (N_10213,N_10041,N_10011);
and U10214 (N_10214,N_10042,N_10004);
xnor U10215 (N_10215,N_10119,N_10013);
nor U10216 (N_10216,N_10018,N_10075);
xnor U10217 (N_10217,N_10117,N_10068);
nor U10218 (N_10218,N_10095,N_10011);
xor U10219 (N_10219,N_10076,N_10056);
nor U10220 (N_10220,N_10020,N_10003);
nand U10221 (N_10221,N_10109,N_10030);
nand U10222 (N_10222,N_10016,N_10003);
xnor U10223 (N_10223,N_10021,N_10005);
xor U10224 (N_10224,N_10030,N_10027);
or U10225 (N_10225,N_10104,N_10046);
or U10226 (N_10226,N_10053,N_10042);
and U10227 (N_10227,N_10024,N_10058);
nor U10228 (N_10228,N_10079,N_10121);
nor U10229 (N_10229,N_10103,N_10054);
nor U10230 (N_10230,N_10024,N_10009);
nand U10231 (N_10231,N_10095,N_10123);
and U10232 (N_10232,N_10078,N_10000);
nor U10233 (N_10233,N_10022,N_10089);
nand U10234 (N_10234,N_10012,N_10109);
or U10235 (N_10235,N_10074,N_10028);
nand U10236 (N_10236,N_10057,N_10064);
or U10237 (N_10237,N_10030,N_10000);
and U10238 (N_10238,N_10046,N_10089);
xor U10239 (N_10239,N_10066,N_10012);
or U10240 (N_10240,N_10084,N_10038);
xnor U10241 (N_10241,N_10083,N_10070);
nor U10242 (N_10242,N_10027,N_10074);
xor U10243 (N_10243,N_10025,N_10113);
and U10244 (N_10244,N_10014,N_10038);
nor U10245 (N_10245,N_10095,N_10067);
xnor U10246 (N_10246,N_10121,N_10083);
nor U10247 (N_10247,N_10015,N_10115);
or U10248 (N_10248,N_10019,N_10005);
and U10249 (N_10249,N_10105,N_10079);
xor U10250 (N_10250,N_10232,N_10171);
and U10251 (N_10251,N_10181,N_10214);
nand U10252 (N_10252,N_10185,N_10230);
nand U10253 (N_10253,N_10217,N_10157);
or U10254 (N_10254,N_10163,N_10241);
nand U10255 (N_10255,N_10125,N_10245);
nand U10256 (N_10256,N_10201,N_10182);
or U10257 (N_10257,N_10248,N_10135);
xnor U10258 (N_10258,N_10138,N_10186);
or U10259 (N_10259,N_10192,N_10155);
xnor U10260 (N_10260,N_10190,N_10223);
xnor U10261 (N_10261,N_10169,N_10152);
and U10262 (N_10262,N_10200,N_10141);
nor U10263 (N_10263,N_10151,N_10146);
or U10264 (N_10264,N_10193,N_10249);
nor U10265 (N_10265,N_10161,N_10239);
xor U10266 (N_10266,N_10206,N_10129);
nor U10267 (N_10267,N_10228,N_10132);
nor U10268 (N_10268,N_10220,N_10227);
xnor U10269 (N_10269,N_10172,N_10153);
xor U10270 (N_10270,N_10194,N_10231);
and U10271 (N_10271,N_10224,N_10150);
and U10272 (N_10272,N_10187,N_10188);
and U10273 (N_10273,N_10213,N_10204);
xor U10274 (N_10274,N_10133,N_10134);
nand U10275 (N_10275,N_10203,N_10226);
nor U10276 (N_10276,N_10229,N_10127);
or U10277 (N_10277,N_10158,N_10137);
xor U10278 (N_10278,N_10131,N_10128);
nand U10279 (N_10279,N_10173,N_10196);
xor U10280 (N_10280,N_10234,N_10164);
nor U10281 (N_10281,N_10160,N_10130);
nor U10282 (N_10282,N_10235,N_10195);
nor U10283 (N_10283,N_10143,N_10174);
xnor U10284 (N_10284,N_10215,N_10233);
or U10285 (N_10285,N_10210,N_10209);
nor U10286 (N_10286,N_10205,N_10178);
nor U10287 (N_10287,N_10238,N_10149);
nor U10288 (N_10288,N_10176,N_10179);
nor U10289 (N_10289,N_10198,N_10243);
and U10290 (N_10290,N_10183,N_10170);
nand U10291 (N_10291,N_10236,N_10218);
or U10292 (N_10292,N_10162,N_10154);
and U10293 (N_10293,N_10189,N_10221);
nor U10294 (N_10294,N_10247,N_10126);
xnor U10295 (N_10295,N_10184,N_10147);
and U10296 (N_10296,N_10207,N_10142);
or U10297 (N_10297,N_10202,N_10148);
nand U10298 (N_10298,N_10165,N_10240);
nand U10299 (N_10299,N_10168,N_10212);
or U10300 (N_10300,N_10145,N_10216);
or U10301 (N_10301,N_10219,N_10136);
and U10302 (N_10302,N_10159,N_10225);
nor U10303 (N_10303,N_10191,N_10244);
or U10304 (N_10304,N_10139,N_10167);
or U10305 (N_10305,N_10177,N_10246);
nand U10306 (N_10306,N_10166,N_10237);
xor U10307 (N_10307,N_10180,N_10175);
xor U10308 (N_10308,N_10140,N_10211);
nor U10309 (N_10309,N_10199,N_10197);
or U10310 (N_10310,N_10242,N_10156);
xnor U10311 (N_10311,N_10222,N_10144);
nor U10312 (N_10312,N_10208,N_10196);
xnor U10313 (N_10313,N_10150,N_10135);
and U10314 (N_10314,N_10209,N_10240);
nor U10315 (N_10315,N_10125,N_10213);
and U10316 (N_10316,N_10237,N_10189);
and U10317 (N_10317,N_10229,N_10249);
and U10318 (N_10318,N_10236,N_10129);
nand U10319 (N_10319,N_10244,N_10198);
xor U10320 (N_10320,N_10153,N_10139);
nand U10321 (N_10321,N_10127,N_10206);
nand U10322 (N_10322,N_10221,N_10239);
nand U10323 (N_10323,N_10139,N_10154);
nor U10324 (N_10324,N_10127,N_10143);
xor U10325 (N_10325,N_10234,N_10225);
xnor U10326 (N_10326,N_10183,N_10129);
nor U10327 (N_10327,N_10231,N_10244);
nor U10328 (N_10328,N_10222,N_10200);
and U10329 (N_10329,N_10165,N_10175);
nand U10330 (N_10330,N_10144,N_10151);
nand U10331 (N_10331,N_10246,N_10155);
nor U10332 (N_10332,N_10221,N_10229);
xnor U10333 (N_10333,N_10215,N_10128);
nor U10334 (N_10334,N_10181,N_10227);
nand U10335 (N_10335,N_10132,N_10245);
or U10336 (N_10336,N_10206,N_10131);
or U10337 (N_10337,N_10180,N_10155);
nor U10338 (N_10338,N_10210,N_10246);
nor U10339 (N_10339,N_10244,N_10176);
nor U10340 (N_10340,N_10220,N_10128);
or U10341 (N_10341,N_10213,N_10135);
and U10342 (N_10342,N_10169,N_10143);
nand U10343 (N_10343,N_10210,N_10136);
nor U10344 (N_10344,N_10164,N_10238);
or U10345 (N_10345,N_10159,N_10167);
nand U10346 (N_10346,N_10145,N_10202);
or U10347 (N_10347,N_10236,N_10127);
and U10348 (N_10348,N_10159,N_10162);
or U10349 (N_10349,N_10248,N_10145);
xor U10350 (N_10350,N_10132,N_10234);
xnor U10351 (N_10351,N_10187,N_10237);
nand U10352 (N_10352,N_10190,N_10147);
and U10353 (N_10353,N_10184,N_10212);
or U10354 (N_10354,N_10168,N_10196);
nand U10355 (N_10355,N_10241,N_10225);
or U10356 (N_10356,N_10155,N_10179);
nand U10357 (N_10357,N_10241,N_10168);
nor U10358 (N_10358,N_10174,N_10219);
and U10359 (N_10359,N_10191,N_10209);
xnor U10360 (N_10360,N_10129,N_10164);
or U10361 (N_10361,N_10243,N_10182);
nor U10362 (N_10362,N_10180,N_10213);
nand U10363 (N_10363,N_10174,N_10162);
nand U10364 (N_10364,N_10160,N_10150);
xor U10365 (N_10365,N_10169,N_10196);
nand U10366 (N_10366,N_10222,N_10132);
nand U10367 (N_10367,N_10176,N_10249);
and U10368 (N_10368,N_10186,N_10213);
and U10369 (N_10369,N_10159,N_10228);
xnor U10370 (N_10370,N_10219,N_10238);
xor U10371 (N_10371,N_10143,N_10211);
or U10372 (N_10372,N_10138,N_10193);
xor U10373 (N_10373,N_10236,N_10191);
and U10374 (N_10374,N_10202,N_10201);
and U10375 (N_10375,N_10322,N_10365);
nand U10376 (N_10376,N_10367,N_10331);
nor U10377 (N_10377,N_10257,N_10259);
nor U10378 (N_10378,N_10319,N_10358);
nor U10379 (N_10379,N_10370,N_10303);
nand U10380 (N_10380,N_10260,N_10346);
or U10381 (N_10381,N_10366,N_10361);
nand U10382 (N_10382,N_10280,N_10353);
or U10383 (N_10383,N_10294,N_10283);
nand U10384 (N_10384,N_10332,N_10251);
xor U10385 (N_10385,N_10270,N_10253);
xor U10386 (N_10386,N_10267,N_10325);
nand U10387 (N_10387,N_10344,N_10306);
and U10388 (N_10388,N_10286,N_10314);
and U10389 (N_10389,N_10363,N_10268);
or U10390 (N_10390,N_10310,N_10349);
and U10391 (N_10391,N_10288,N_10289);
and U10392 (N_10392,N_10273,N_10368);
xor U10393 (N_10393,N_10300,N_10277);
xnor U10394 (N_10394,N_10320,N_10296);
nor U10395 (N_10395,N_10278,N_10263);
xor U10396 (N_10396,N_10287,N_10364);
nand U10397 (N_10397,N_10250,N_10282);
xnor U10398 (N_10398,N_10323,N_10359);
xor U10399 (N_10399,N_10254,N_10348);
nand U10400 (N_10400,N_10336,N_10269);
or U10401 (N_10401,N_10338,N_10329);
nand U10402 (N_10402,N_10312,N_10261);
nor U10403 (N_10403,N_10318,N_10255);
and U10404 (N_10404,N_10276,N_10274);
and U10405 (N_10405,N_10295,N_10351);
nor U10406 (N_10406,N_10284,N_10307);
or U10407 (N_10407,N_10374,N_10317);
xnor U10408 (N_10408,N_10357,N_10271);
xor U10409 (N_10409,N_10302,N_10256);
nand U10410 (N_10410,N_10292,N_10293);
nand U10411 (N_10411,N_10321,N_10308);
nand U10412 (N_10412,N_10311,N_10266);
and U10413 (N_10413,N_10356,N_10275);
nand U10414 (N_10414,N_10354,N_10298);
and U10415 (N_10415,N_10315,N_10285);
xnor U10416 (N_10416,N_10258,N_10355);
or U10417 (N_10417,N_10372,N_10337);
or U10418 (N_10418,N_10279,N_10343);
nand U10419 (N_10419,N_10340,N_10262);
xnor U10420 (N_10420,N_10371,N_10335);
and U10421 (N_10421,N_10301,N_10324);
nand U10422 (N_10422,N_10334,N_10339);
nand U10423 (N_10423,N_10330,N_10264);
or U10424 (N_10424,N_10309,N_10347);
nor U10425 (N_10425,N_10345,N_10305);
or U10426 (N_10426,N_10290,N_10326);
nor U10427 (N_10427,N_10297,N_10342);
xor U10428 (N_10428,N_10341,N_10369);
xnor U10429 (N_10429,N_10313,N_10327);
xor U10430 (N_10430,N_10272,N_10328);
and U10431 (N_10431,N_10360,N_10350);
xor U10432 (N_10432,N_10281,N_10291);
or U10433 (N_10433,N_10304,N_10316);
nand U10434 (N_10434,N_10252,N_10299);
xor U10435 (N_10435,N_10373,N_10333);
nand U10436 (N_10436,N_10265,N_10352);
xnor U10437 (N_10437,N_10362,N_10292);
or U10438 (N_10438,N_10305,N_10292);
nand U10439 (N_10439,N_10278,N_10296);
and U10440 (N_10440,N_10300,N_10270);
and U10441 (N_10441,N_10370,N_10271);
nor U10442 (N_10442,N_10337,N_10300);
nand U10443 (N_10443,N_10340,N_10294);
nand U10444 (N_10444,N_10255,N_10360);
or U10445 (N_10445,N_10307,N_10365);
nor U10446 (N_10446,N_10345,N_10284);
nand U10447 (N_10447,N_10290,N_10259);
and U10448 (N_10448,N_10259,N_10354);
and U10449 (N_10449,N_10328,N_10270);
or U10450 (N_10450,N_10327,N_10343);
and U10451 (N_10451,N_10275,N_10359);
and U10452 (N_10452,N_10295,N_10322);
nor U10453 (N_10453,N_10267,N_10254);
nor U10454 (N_10454,N_10335,N_10365);
and U10455 (N_10455,N_10372,N_10265);
xor U10456 (N_10456,N_10282,N_10315);
or U10457 (N_10457,N_10352,N_10256);
and U10458 (N_10458,N_10265,N_10266);
xor U10459 (N_10459,N_10337,N_10306);
and U10460 (N_10460,N_10365,N_10374);
nand U10461 (N_10461,N_10316,N_10298);
xor U10462 (N_10462,N_10354,N_10289);
xor U10463 (N_10463,N_10352,N_10333);
and U10464 (N_10464,N_10293,N_10346);
or U10465 (N_10465,N_10320,N_10335);
nand U10466 (N_10466,N_10259,N_10281);
nor U10467 (N_10467,N_10307,N_10362);
nand U10468 (N_10468,N_10373,N_10318);
and U10469 (N_10469,N_10279,N_10310);
nor U10470 (N_10470,N_10308,N_10324);
nor U10471 (N_10471,N_10334,N_10324);
xnor U10472 (N_10472,N_10274,N_10312);
and U10473 (N_10473,N_10347,N_10336);
nand U10474 (N_10474,N_10369,N_10256);
and U10475 (N_10475,N_10315,N_10259);
nand U10476 (N_10476,N_10363,N_10319);
or U10477 (N_10477,N_10250,N_10363);
nand U10478 (N_10478,N_10348,N_10296);
nand U10479 (N_10479,N_10256,N_10328);
xor U10480 (N_10480,N_10326,N_10366);
nor U10481 (N_10481,N_10302,N_10329);
or U10482 (N_10482,N_10339,N_10252);
xor U10483 (N_10483,N_10270,N_10349);
nand U10484 (N_10484,N_10340,N_10258);
xnor U10485 (N_10485,N_10268,N_10304);
xor U10486 (N_10486,N_10305,N_10294);
and U10487 (N_10487,N_10285,N_10310);
nor U10488 (N_10488,N_10265,N_10261);
nand U10489 (N_10489,N_10310,N_10347);
and U10490 (N_10490,N_10278,N_10307);
or U10491 (N_10491,N_10341,N_10357);
and U10492 (N_10492,N_10368,N_10342);
nand U10493 (N_10493,N_10309,N_10285);
or U10494 (N_10494,N_10321,N_10286);
or U10495 (N_10495,N_10293,N_10356);
or U10496 (N_10496,N_10367,N_10313);
nor U10497 (N_10497,N_10322,N_10287);
xnor U10498 (N_10498,N_10304,N_10277);
nand U10499 (N_10499,N_10261,N_10320);
nand U10500 (N_10500,N_10400,N_10421);
xor U10501 (N_10501,N_10479,N_10438);
nand U10502 (N_10502,N_10485,N_10408);
nand U10503 (N_10503,N_10390,N_10443);
xor U10504 (N_10504,N_10412,N_10460);
or U10505 (N_10505,N_10489,N_10379);
or U10506 (N_10506,N_10447,N_10477);
nand U10507 (N_10507,N_10461,N_10487);
xnor U10508 (N_10508,N_10466,N_10395);
nor U10509 (N_10509,N_10453,N_10486);
xnor U10510 (N_10510,N_10482,N_10493);
nor U10511 (N_10511,N_10449,N_10397);
nor U10512 (N_10512,N_10498,N_10403);
nand U10513 (N_10513,N_10456,N_10441);
and U10514 (N_10514,N_10430,N_10423);
nand U10515 (N_10515,N_10478,N_10474);
and U10516 (N_10516,N_10442,N_10406);
or U10517 (N_10517,N_10391,N_10469);
nand U10518 (N_10518,N_10427,N_10416);
nor U10519 (N_10519,N_10417,N_10378);
and U10520 (N_10520,N_10381,N_10472);
or U10521 (N_10521,N_10413,N_10396);
nor U10522 (N_10522,N_10420,N_10376);
or U10523 (N_10523,N_10422,N_10483);
xnor U10524 (N_10524,N_10384,N_10428);
or U10525 (N_10525,N_10475,N_10492);
or U10526 (N_10526,N_10429,N_10459);
nor U10527 (N_10527,N_10468,N_10457);
and U10528 (N_10528,N_10452,N_10484);
nand U10529 (N_10529,N_10434,N_10424);
or U10530 (N_10530,N_10439,N_10497);
nor U10531 (N_10531,N_10464,N_10377);
nor U10532 (N_10532,N_10436,N_10389);
nand U10533 (N_10533,N_10448,N_10414);
and U10534 (N_10534,N_10445,N_10385);
or U10535 (N_10535,N_10432,N_10399);
and U10536 (N_10536,N_10393,N_10394);
nand U10537 (N_10537,N_10415,N_10481);
nor U10538 (N_10538,N_10496,N_10407);
xor U10539 (N_10539,N_10405,N_10433);
or U10540 (N_10540,N_10435,N_10499);
xnor U10541 (N_10541,N_10387,N_10454);
xnor U10542 (N_10542,N_10470,N_10490);
xor U10543 (N_10543,N_10462,N_10382);
or U10544 (N_10544,N_10473,N_10426);
or U10545 (N_10545,N_10440,N_10404);
or U10546 (N_10546,N_10398,N_10495);
xor U10547 (N_10547,N_10491,N_10431);
or U10548 (N_10548,N_10388,N_10375);
nor U10549 (N_10549,N_10410,N_10463);
or U10550 (N_10550,N_10465,N_10451);
xor U10551 (N_10551,N_10419,N_10446);
or U10552 (N_10552,N_10392,N_10437);
or U10553 (N_10553,N_10476,N_10411);
nand U10554 (N_10554,N_10386,N_10401);
nor U10555 (N_10555,N_10471,N_10380);
nand U10556 (N_10556,N_10480,N_10402);
xor U10557 (N_10557,N_10488,N_10383);
and U10558 (N_10558,N_10425,N_10450);
xnor U10559 (N_10559,N_10455,N_10494);
nand U10560 (N_10560,N_10444,N_10467);
nor U10561 (N_10561,N_10418,N_10458);
xor U10562 (N_10562,N_10409,N_10407);
nand U10563 (N_10563,N_10417,N_10484);
or U10564 (N_10564,N_10394,N_10487);
nand U10565 (N_10565,N_10403,N_10389);
or U10566 (N_10566,N_10452,N_10456);
or U10567 (N_10567,N_10450,N_10493);
and U10568 (N_10568,N_10397,N_10496);
nand U10569 (N_10569,N_10475,N_10488);
nor U10570 (N_10570,N_10384,N_10394);
or U10571 (N_10571,N_10482,N_10453);
and U10572 (N_10572,N_10419,N_10436);
and U10573 (N_10573,N_10392,N_10398);
xnor U10574 (N_10574,N_10472,N_10379);
nand U10575 (N_10575,N_10385,N_10411);
nor U10576 (N_10576,N_10431,N_10487);
nand U10577 (N_10577,N_10454,N_10411);
xnor U10578 (N_10578,N_10424,N_10425);
or U10579 (N_10579,N_10481,N_10454);
xnor U10580 (N_10580,N_10402,N_10378);
and U10581 (N_10581,N_10466,N_10474);
or U10582 (N_10582,N_10409,N_10486);
and U10583 (N_10583,N_10483,N_10417);
nor U10584 (N_10584,N_10410,N_10413);
or U10585 (N_10585,N_10477,N_10446);
or U10586 (N_10586,N_10473,N_10404);
xnor U10587 (N_10587,N_10450,N_10409);
xnor U10588 (N_10588,N_10452,N_10426);
and U10589 (N_10589,N_10438,N_10483);
or U10590 (N_10590,N_10485,N_10419);
xor U10591 (N_10591,N_10380,N_10453);
nor U10592 (N_10592,N_10455,N_10420);
or U10593 (N_10593,N_10385,N_10388);
nand U10594 (N_10594,N_10454,N_10473);
and U10595 (N_10595,N_10476,N_10414);
xor U10596 (N_10596,N_10472,N_10398);
and U10597 (N_10597,N_10486,N_10497);
xnor U10598 (N_10598,N_10406,N_10424);
xor U10599 (N_10599,N_10391,N_10465);
xor U10600 (N_10600,N_10451,N_10402);
or U10601 (N_10601,N_10492,N_10479);
nand U10602 (N_10602,N_10429,N_10454);
or U10603 (N_10603,N_10475,N_10478);
xor U10604 (N_10604,N_10496,N_10443);
and U10605 (N_10605,N_10471,N_10400);
or U10606 (N_10606,N_10377,N_10378);
nor U10607 (N_10607,N_10467,N_10495);
or U10608 (N_10608,N_10453,N_10436);
nor U10609 (N_10609,N_10417,N_10455);
nand U10610 (N_10610,N_10430,N_10448);
nor U10611 (N_10611,N_10486,N_10438);
and U10612 (N_10612,N_10449,N_10461);
and U10613 (N_10613,N_10430,N_10497);
nand U10614 (N_10614,N_10455,N_10402);
nand U10615 (N_10615,N_10387,N_10401);
nand U10616 (N_10616,N_10422,N_10388);
and U10617 (N_10617,N_10493,N_10460);
xor U10618 (N_10618,N_10387,N_10499);
and U10619 (N_10619,N_10484,N_10411);
nand U10620 (N_10620,N_10417,N_10440);
or U10621 (N_10621,N_10490,N_10497);
xor U10622 (N_10622,N_10401,N_10407);
nor U10623 (N_10623,N_10454,N_10397);
nor U10624 (N_10624,N_10468,N_10437);
nor U10625 (N_10625,N_10545,N_10593);
xor U10626 (N_10626,N_10548,N_10518);
nor U10627 (N_10627,N_10575,N_10582);
nor U10628 (N_10628,N_10539,N_10604);
nor U10629 (N_10629,N_10570,N_10577);
nand U10630 (N_10630,N_10574,N_10532);
xor U10631 (N_10631,N_10590,N_10534);
nand U10632 (N_10632,N_10504,N_10503);
or U10633 (N_10633,N_10515,N_10541);
nor U10634 (N_10634,N_10585,N_10528);
and U10635 (N_10635,N_10602,N_10588);
nor U10636 (N_10636,N_10526,N_10546);
nor U10637 (N_10637,N_10563,N_10573);
xnor U10638 (N_10638,N_10513,N_10620);
or U10639 (N_10639,N_10537,N_10603);
nand U10640 (N_10640,N_10512,N_10540);
and U10641 (N_10641,N_10524,N_10578);
or U10642 (N_10642,N_10616,N_10514);
xor U10643 (N_10643,N_10619,N_10567);
xor U10644 (N_10644,N_10591,N_10556);
and U10645 (N_10645,N_10510,N_10558);
nand U10646 (N_10646,N_10505,N_10581);
nand U10647 (N_10647,N_10576,N_10561);
nor U10648 (N_10648,N_10517,N_10615);
nand U10649 (N_10649,N_10564,N_10525);
xnor U10650 (N_10650,N_10552,N_10624);
xor U10651 (N_10651,N_10580,N_10569);
or U10652 (N_10652,N_10613,N_10572);
xor U10653 (N_10653,N_10598,N_10523);
and U10654 (N_10654,N_10543,N_10506);
nand U10655 (N_10655,N_10622,N_10522);
nand U10656 (N_10656,N_10554,N_10511);
xor U10657 (N_10657,N_10562,N_10589);
or U10658 (N_10658,N_10507,N_10536);
or U10659 (N_10659,N_10535,N_10623);
nand U10660 (N_10660,N_10586,N_10520);
xnor U10661 (N_10661,N_10551,N_10607);
xor U10662 (N_10662,N_10583,N_10547);
and U10663 (N_10663,N_10599,N_10521);
nor U10664 (N_10664,N_10542,N_10538);
xor U10665 (N_10665,N_10618,N_10502);
nand U10666 (N_10666,N_10550,N_10519);
and U10667 (N_10667,N_10544,N_10555);
or U10668 (N_10668,N_10533,N_10608);
nor U10669 (N_10669,N_10594,N_10549);
nand U10670 (N_10670,N_10584,N_10531);
xnor U10671 (N_10671,N_10612,N_10508);
xnor U10672 (N_10672,N_10596,N_10529);
xnor U10673 (N_10673,N_10587,N_10571);
or U10674 (N_10674,N_10559,N_10606);
xnor U10675 (N_10675,N_10610,N_10557);
nand U10676 (N_10676,N_10565,N_10566);
and U10677 (N_10677,N_10597,N_10501);
and U10678 (N_10678,N_10617,N_10509);
nor U10679 (N_10679,N_10611,N_10579);
or U10680 (N_10680,N_10516,N_10560);
nor U10681 (N_10681,N_10568,N_10527);
xnor U10682 (N_10682,N_10595,N_10600);
xor U10683 (N_10683,N_10614,N_10621);
and U10684 (N_10684,N_10601,N_10592);
nor U10685 (N_10685,N_10530,N_10500);
or U10686 (N_10686,N_10553,N_10609);
nor U10687 (N_10687,N_10605,N_10542);
nor U10688 (N_10688,N_10524,N_10503);
nand U10689 (N_10689,N_10551,N_10552);
nand U10690 (N_10690,N_10604,N_10607);
nor U10691 (N_10691,N_10599,N_10587);
nor U10692 (N_10692,N_10598,N_10569);
or U10693 (N_10693,N_10544,N_10511);
xnor U10694 (N_10694,N_10576,N_10518);
or U10695 (N_10695,N_10550,N_10617);
nand U10696 (N_10696,N_10577,N_10502);
nand U10697 (N_10697,N_10571,N_10617);
and U10698 (N_10698,N_10578,N_10624);
xor U10699 (N_10699,N_10560,N_10540);
xor U10700 (N_10700,N_10534,N_10550);
and U10701 (N_10701,N_10518,N_10566);
and U10702 (N_10702,N_10503,N_10549);
xnor U10703 (N_10703,N_10504,N_10584);
nand U10704 (N_10704,N_10566,N_10551);
and U10705 (N_10705,N_10588,N_10509);
nand U10706 (N_10706,N_10563,N_10553);
and U10707 (N_10707,N_10598,N_10613);
nor U10708 (N_10708,N_10511,N_10562);
and U10709 (N_10709,N_10540,N_10545);
or U10710 (N_10710,N_10559,N_10597);
and U10711 (N_10711,N_10547,N_10563);
nor U10712 (N_10712,N_10551,N_10622);
xor U10713 (N_10713,N_10524,N_10606);
xnor U10714 (N_10714,N_10621,N_10605);
nand U10715 (N_10715,N_10504,N_10617);
and U10716 (N_10716,N_10541,N_10521);
and U10717 (N_10717,N_10506,N_10525);
nor U10718 (N_10718,N_10586,N_10551);
nor U10719 (N_10719,N_10508,N_10586);
xor U10720 (N_10720,N_10599,N_10557);
and U10721 (N_10721,N_10519,N_10615);
nor U10722 (N_10722,N_10536,N_10612);
xnor U10723 (N_10723,N_10596,N_10554);
or U10724 (N_10724,N_10504,N_10611);
and U10725 (N_10725,N_10597,N_10604);
or U10726 (N_10726,N_10558,N_10531);
xnor U10727 (N_10727,N_10558,N_10544);
nor U10728 (N_10728,N_10553,N_10572);
nand U10729 (N_10729,N_10566,N_10538);
or U10730 (N_10730,N_10532,N_10552);
nand U10731 (N_10731,N_10541,N_10532);
or U10732 (N_10732,N_10592,N_10572);
or U10733 (N_10733,N_10604,N_10510);
or U10734 (N_10734,N_10519,N_10607);
nor U10735 (N_10735,N_10521,N_10558);
or U10736 (N_10736,N_10613,N_10559);
nor U10737 (N_10737,N_10535,N_10531);
nor U10738 (N_10738,N_10511,N_10521);
xnor U10739 (N_10739,N_10522,N_10594);
or U10740 (N_10740,N_10562,N_10538);
nor U10741 (N_10741,N_10603,N_10545);
nand U10742 (N_10742,N_10576,N_10525);
or U10743 (N_10743,N_10572,N_10520);
xnor U10744 (N_10744,N_10598,N_10507);
and U10745 (N_10745,N_10547,N_10544);
xor U10746 (N_10746,N_10572,N_10545);
nor U10747 (N_10747,N_10520,N_10566);
and U10748 (N_10748,N_10552,N_10503);
or U10749 (N_10749,N_10556,N_10570);
nand U10750 (N_10750,N_10649,N_10733);
or U10751 (N_10751,N_10667,N_10743);
nand U10752 (N_10752,N_10734,N_10653);
and U10753 (N_10753,N_10683,N_10626);
nor U10754 (N_10754,N_10638,N_10723);
nor U10755 (N_10755,N_10701,N_10720);
nand U10756 (N_10756,N_10648,N_10738);
or U10757 (N_10757,N_10729,N_10652);
or U10758 (N_10758,N_10680,N_10741);
nor U10759 (N_10759,N_10654,N_10708);
nand U10760 (N_10760,N_10689,N_10742);
and U10761 (N_10761,N_10642,N_10631);
and U10762 (N_10762,N_10677,N_10632);
or U10763 (N_10763,N_10712,N_10727);
xor U10764 (N_10764,N_10684,N_10744);
and U10765 (N_10765,N_10697,N_10656);
nand U10766 (N_10766,N_10692,N_10726);
or U10767 (N_10767,N_10637,N_10629);
nand U10768 (N_10768,N_10661,N_10650);
nor U10769 (N_10769,N_10737,N_10735);
nand U10770 (N_10770,N_10658,N_10685);
xnor U10771 (N_10771,N_10736,N_10625);
or U10772 (N_10772,N_10676,N_10688);
nand U10773 (N_10773,N_10659,N_10678);
nand U10774 (N_10774,N_10731,N_10657);
nor U10775 (N_10775,N_10673,N_10746);
and U10776 (N_10776,N_10663,N_10717);
xor U10777 (N_10777,N_10635,N_10671);
nor U10778 (N_10778,N_10640,N_10698);
nand U10779 (N_10779,N_10662,N_10706);
xor U10780 (N_10780,N_10628,N_10660);
and U10781 (N_10781,N_10721,N_10704);
nand U10782 (N_10782,N_10641,N_10724);
nand U10783 (N_10783,N_10730,N_10747);
and U10784 (N_10784,N_10695,N_10651);
nor U10785 (N_10785,N_10693,N_10655);
nor U10786 (N_10786,N_10687,N_10716);
xor U10787 (N_10787,N_10645,N_10740);
or U10788 (N_10788,N_10728,N_10690);
nand U10789 (N_10789,N_10634,N_10674);
and U10790 (N_10790,N_10679,N_10718);
xnor U10791 (N_10791,N_10696,N_10636);
nand U10792 (N_10792,N_10719,N_10694);
and U10793 (N_10793,N_10745,N_10664);
or U10794 (N_10794,N_10639,N_10666);
or U10795 (N_10795,N_10711,N_10700);
xor U10796 (N_10796,N_10669,N_10691);
nor U10797 (N_10797,N_10665,N_10670);
and U10798 (N_10798,N_10709,N_10748);
and U10799 (N_10799,N_10705,N_10725);
and U10800 (N_10800,N_10722,N_10668);
xnor U10801 (N_10801,N_10710,N_10633);
nand U10802 (N_10802,N_10713,N_10714);
xnor U10803 (N_10803,N_10647,N_10702);
and U10804 (N_10804,N_10732,N_10739);
xnor U10805 (N_10805,N_10630,N_10675);
and U10806 (N_10806,N_10715,N_10707);
xor U10807 (N_10807,N_10699,N_10627);
nor U10808 (N_10808,N_10646,N_10682);
or U10809 (N_10809,N_10686,N_10749);
or U10810 (N_10810,N_10643,N_10703);
or U10811 (N_10811,N_10672,N_10644);
and U10812 (N_10812,N_10681,N_10644);
or U10813 (N_10813,N_10735,N_10641);
or U10814 (N_10814,N_10672,N_10709);
nand U10815 (N_10815,N_10732,N_10662);
nand U10816 (N_10816,N_10660,N_10749);
or U10817 (N_10817,N_10629,N_10723);
and U10818 (N_10818,N_10661,N_10689);
nand U10819 (N_10819,N_10692,N_10638);
nand U10820 (N_10820,N_10749,N_10631);
nand U10821 (N_10821,N_10638,N_10629);
nor U10822 (N_10822,N_10682,N_10654);
or U10823 (N_10823,N_10707,N_10747);
xor U10824 (N_10824,N_10721,N_10646);
xnor U10825 (N_10825,N_10645,N_10739);
xor U10826 (N_10826,N_10697,N_10703);
nand U10827 (N_10827,N_10710,N_10640);
nor U10828 (N_10828,N_10746,N_10638);
or U10829 (N_10829,N_10652,N_10630);
xor U10830 (N_10830,N_10705,N_10711);
nand U10831 (N_10831,N_10707,N_10685);
or U10832 (N_10832,N_10662,N_10631);
nand U10833 (N_10833,N_10656,N_10691);
or U10834 (N_10834,N_10665,N_10642);
nor U10835 (N_10835,N_10666,N_10738);
and U10836 (N_10836,N_10675,N_10626);
nand U10837 (N_10837,N_10631,N_10742);
nand U10838 (N_10838,N_10705,N_10684);
nand U10839 (N_10839,N_10724,N_10656);
or U10840 (N_10840,N_10627,N_10676);
xor U10841 (N_10841,N_10723,N_10709);
or U10842 (N_10842,N_10660,N_10744);
xor U10843 (N_10843,N_10625,N_10707);
nor U10844 (N_10844,N_10721,N_10647);
and U10845 (N_10845,N_10722,N_10744);
or U10846 (N_10846,N_10655,N_10733);
and U10847 (N_10847,N_10705,N_10745);
nand U10848 (N_10848,N_10706,N_10697);
nand U10849 (N_10849,N_10718,N_10658);
and U10850 (N_10850,N_10643,N_10625);
nand U10851 (N_10851,N_10630,N_10744);
nand U10852 (N_10852,N_10747,N_10710);
nor U10853 (N_10853,N_10716,N_10642);
xor U10854 (N_10854,N_10739,N_10725);
and U10855 (N_10855,N_10632,N_10666);
nand U10856 (N_10856,N_10653,N_10709);
nand U10857 (N_10857,N_10733,N_10747);
nor U10858 (N_10858,N_10672,N_10712);
or U10859 (N_10859,N_10717,N_10678);
and U10860 (N_10860,N_10643,N_10636);
nor U10861 (N_10861,N_10697,N_10659);
nor U10862 (N_10862,N_10690,N_10625);
or U10863 (N_10863,N_10738,N_10637);
or U10864 (N_10864,N_10699,N_10721);
or U10865 (N_10865,N_10696,N_10675);
nand U10866 (N_10866,N_10730,N_10679);
and U10867 (N_10867,N_10731,N_10631);
or U10868 (N_10868,N_10739,N_10676);
nand U10869 (N_10869,N_10662,N_10649);
nand U10870 (N_10870,N_10681,N_10746);
xor U10871 (N_10871,N_10641,N_10708);
and U10872 (N_10872,N_10639,N_10654);
xnor U10873 (N_10873,N_10712,N_10633);
and U10874 (N_10874,N_10646,N_10626);
nor U10875 (N_10875,N_10776,N_10795);
xor U10876 (N_10876,N_10778,N_10822);
and U10877 (N_10877,N_10785,N_10773);
xor U10878 (N_10878,N_10844,N_10803);
or U10879 (N_10879,N_10834,N_10760);
and U10880 (N_10880,N_10801,N_10867);
xor U10881 (N_10881,N_10861,N_10824);
nor U10882 (N_10882,N_10807,N_10793);
nand U10883 (N_10883,N_10837,N_10752);
or U10884 (N_10884,N_10839,N_10765);
nand U10885 (N_10885,N_10852,N_10851);
nand U10886 (N_10886,N_10836,N_10854);
nor U10887 (N_10887,N_10857,N_10812);
or U10888 (N_10888,N_10826,N_10869);
xnor U10889 (N_10889,N_10868,N_10823);
nor U10890 (N_10890,N_10790,N_10835);
or U10891 (N_10891,N_10847,N_10753);
nor U10892 (N_10892,N_10865,N_10759);
and U10893 (N_10893,N_10814,N_10859);
and U10894 (N_10894,N_10789,N_10779);
nor U10895 (N_10895,N_10816,N_10802);
nand U10896 (N_10896,N_10827,N_10770);
xor U10897 (N_10897,N_10784,N_10758);
nor U10898 (N_10898,N_10856,N_10870);
or U10899 (N_10899,N_10848,N_10831);
nand U10900 (N_10900,N_10781,N_10833);
and U10901 (N_10901,N_10855,N_10756);
xor U10902 (N_10902,N_10806,N_10841);
and U10903 (N_10903,N_10866,N_10840);
or U10904 (N_10904,N_10761,N_10863);
nand U10905 (N_10905,N_10764,N_10767);
nand U10906 (N_10906,N_10813,N_10750);
and U10907 (N_10907,N_10874,N_10843);
nor U10908 (N_10908,N_10792,N_10860);
and U10909 (N_10909,N_10825,N_10762);
or U10910 (N_10910,N_10809,N_10853);
or U10911 (N_10911,N_10787,N_10820);
or U10912 (N_10912,N_10810,N_10817);
nand U10913 (N_10913,N_10872,N_10766);
xor U10914 (N_10914,N_10811,N_10754);
or U10915 (N_10915,N_10838,N_10828);
nand U10916 (N_10916,N_10786,N_10815);
nor U10917 (N_10917,N_10780,N_10796);
and U10918 (N_10918,N_10804,N_10768);
and U10919 (N_10919,N_10849,N_10800);
nor U10920 (N_10920,N_10783,N_10821);
nand U10921 (N_10921,N_10805,N_10858);
xor U10922 (N_10922,N_10871,N_10799);
and U10923 (N_10923,N_10769,N_10782);
nor U10924 (N_10924,N_10797,N_10788);
xnor U10925 (N_10925,N_10763,N_10846);
xor U10926 (N_10926,N_10772,N_10873);
and U10927 (N_10927,N_10794,N_10755);
nor U10928 (N_10928,N_10830,N_10845);
xnor U10929 (N_10929,N_10757,N_10818);
nand U10930 (N_10930,N_10862,N_10832);
xor U10931 (N_10931,N_10819,N_10771);
nand U10932 (N_10932,N_10774,N_10864);
nand U10933 (N_10933,N_10775,N_10791);
or U10934 (N_10934,N_10808,N_10777);
or U10935 (N_10935,N_10798,N_10850);
and U10936 (N_10936,N_10829,N_10751);
xnor U10937 (N_10937,N_10842,N_10751);
nor U10938 (N_10938,N_10857,N_10865);
nor U10939 (N_10939,N_10842,N_10763);
nand U10940 (N_10940,N_10769,N_10832);
xnor U10941 (N_10941,N_10767,N_10795);
and U10942 (N_10942,N_10796,N_10832);
and U10943 (N_10943,N_10768,N_10758);
and U10944 (N_10944,N_10811,N_10797);
or U10945 (N_10945,N_10757,N_10862);
nor U10946 (N_10946,N_10855,N_10781);
or U10947 (N_10947,N_10844,N_10865);
nor U10948 (N_10948,N_10765,N_10853);
xor U10949 (N_10949,N_10787,N_10844);
or U10950 (N_10950,N_10838,N_10790);
or U10951 (N_10951,N_10815,N_10752);
xor U10952 (N_10952,N_10792,N_10812);
or U10953 (N_10953,N_10805,N_10788);
xnor U10954 (N_10954,N_10764,N_10784);
or U10955 (N_10955,N_10753,N_10795);
and U10956 (N_10956,N_10830,N_10807);
xor U10957 (N_10957,N_10770,N_10767);
xor U10958 (N_10958,N_10855,N_10801);
nand U10959 (N_10959,N_10827,N_10822);
xor U10960 (N_10960,N_10860,N_10845);
or U10961 (N_10961,N_10865,N_10815);
nor U10962 (N_10962,N_10869,N_10778);
nand U10963 (N_10963,N_10800,N_10869);
xor U10964 (N_10964,N_10796,N_10837);
nand U10965 (N_10965,N_10760,N_10871);
or U10966 (N_10966,N_10827,N_10818);
xnor U10967 (N_10967,N_10811,N_10771);
and U10968 (N_10968,N_10773,N_10834);
or U10969 (N_10969,N_10867,N_10823);
or U10970 (N_10970,N_10804,N_10854);
nand U10971 (N_10971,N_10836,N_10870);
nor U10972 (N_10972,N_10821,N_10792);
xor U10973 (N_10973,N_10859,N_10813);
nor U10974 (N_10974,N_10751,N_10849);
xor U10975 (N_10975,N_10814,N_10758);
xor U10976 (N_10976,N_10825,N_10856);
xor U10977 (N_10977,N_10831,N_10796);
or U10978 (N_10978,N_10835,N_10872);
and U10979 (N_10979,N_10869,N_10846);
nor U10980 (N_10980,N_10850,N_10774);
or U10981 (N_10981,N_10855,N_10836);
nor U10982 (N_10982,N_10848,N_10861);
nand U10983 (N_10983,N_10817,N_10853);
xnor U10984 (N_10984,N_10847,N_10791);
xnor U10985 (N_10985,N_10801,N_10839);
nor U10986 (N_10986,N_10856,N_10809);
or U10987 (N_10987,N_10827,N_10826);
and U10988 (N_10988,N_10752,N_10800);
nor U10989 (N_10989,N_10838,N_10762);
xnor U10990 (N_10990,N_10864,N_10791);
or U10991 (N_10991,N_10859,N_10756);
nor U10992 (N_10992,N_10831,N_10800);
or U10993 (N_10993,N_10820,N_10811);
nand U10994 (N_10994,N_10824,N_10797);
nor U10995 (N_10995,N_10855,N_10869);
or U10996 (N_10996,N_10798,N_10797);
nand U10997 (N_10997,N_10809,N_10810);
nand U10998 (N_10998,N_10819,N_10780);
or U10999 (N_10999,N_10858,N_10860);
nand U11000 (N_11000,N_10876,N_10879);
nor U11001 (N_11001,N_10890,N_10967);
nor U11002 (N_11002,N_10958,N_10990);
or U11003 (N_11003,N_10977,N_10918);
and U11004 (N_11004,N_10933,N_10941);
nor U11005 (N_11005,N_10943,N_10966);
nand U11006 (N_11006,N_10982,N_10908);
or U11007 (N_11007,N_10914,N_10999);
and U11008 (N_11008,N_10994,N_10916);
or U11009 (N_11009,N_10940,N_10934);
xor U11010 (N_11010,N_10885,N_10892);
or U11011 (N_11011,N_10944,N_10878);
xor U11012 (N_11012,N_10884,N_10900);
nand U11013 (N_11013,N_10959,N_10950);
nor U11014 (N_11014,N_10995,N_10954);
or U11015 (N_11015,N_10920,N_10919);
nor U11016 (N_11016,N_10921,N_10927);
and U11017 (N_11017,N_10924,N_10964);
nor U11018 (N_11018,N_10997,N_10989);
nor U11019 (N_11019,N_10893,N_10962);
nor U11020 (N_11020,N_10985,N_10925);
xnor U11021 (N_11021,N_10975,N_10883);
or U11022 (N_11022,N_10948,N_10942);
nand U11023 (N_11023,N_10993,N_10928);
xnor U11024 (N_11024,N_10889,N_10988);
and U11025 (N_11025,N_10930,N_10904);
and U11026 (N_11026,N_10937,N_10931);
nand U11027 (N_11027,N_10875,N_10996);
or U11028 (N_11028,N_10979,N_10935);
or U11029 (N_11029,N_10926,N_10902);
nand U11030 (N_11030,N_10923,N_10907);
nor U11031 (N_11031,N_10909,N_10957);
nor U11032 (N_11032,N_10955,N_10968);
and U11033 (N_11033,N_10915,N_10986);
or U11034 (N_11034,N_10932,N_10929);
nor U11035 (N_11035,N_10898,N_10961);
nor U11036 (N_11036,N_10887,N_10947);
xnor U11037 (N_11037,N_10877,N_10973);
xor U11038 (N_11038,N_10992,N_10984);
nand U11039 (N_11039,N_10891,N_10910);
nand U11040 (N_11040,N_10980,N_10946);
nor U11041 (N_11041,N_10991,N_10906);
xor U11042 (N_11042,N_10911,N_10983);
and U11043 (N_11043,N_10951,N_10903);
nor U11044 (N_11044,N_10978,N_10888);
nand U11045 (N_11045,N_10972,N_10939);
nand U11046 (N_11046,N_10945,N_10901);
xnor U11047 (N_11047,N_10952,N_10969);
nand U11048 (N_11048,N_10905,N_10949);
nor U11049 (N_11049,N_10917,N_10882);
nor U11050 (N_11050,N_10897,N_10953);
nand U11051 (N_11051,N_10894,N_10998);
nand U11052 (N_11052,N_10886,N_10987);
xnor U11053 (N_11053,N_10912,N_10963);
nand U11054 (N_11054,N_10970,N_10896);
nor U11055 (N_11055,N_10974,N_10881);
nand U11056 (N_11056,N_10899,N_10965);
nand U11057 (N_11057,N_10922,N_10895);
and U11058 (N_11058,N_10880,N_10938);
nor U11059 (N_11059,N_10913,N_10960);
and U11060 (N_11060,N_10936,N_10971);
and U11061 (N_11061,N_10976,N_10981);
nor U11062 (N_11062,N_10956,N_10991);
nor U11063 (N_11063,N_10923,N_10912);
nor U11064 (N_11064,N_10894,N_10911);
or U11065 (N_11065,N_10895,N_10878);
xnor U11066 (N_11066,N_10999,N_10888);
or U11067 (N_11067,N_10938,N_10999);
nor U11068 (N_11068,N_10916,N_10969);
xor U11069 (N_11069,N_10878,N_10949);
nor U11070 (N_11070,N_10937,N_10910);
or U11071 (N_11071,N_10968,N_10910);
or U11072 (N_11072,N_10911,N_10939);
or U11073 (N_11073,N_10913,N_10963);
nand U11074 (N_11074,N_10932,N_10965);
nor U11075 (N_11075,N_10887,N_10932);
xor U11076 (N_11076,N_10972,N_10907);
or U11077 (N_11077,N_10950,N_10886);
or U11078 (N_11078,N_10876,N_10966);
xor U11079 (N_11079,N_10974,N_10933);
nor U11080 (N_11080,N_10968,N_10936);
xnor U11081 (N_11081,N_10880,N_10893);
and U11082 (N_11082,N_10970,N_10931);
nand U11083 (N_11083,N_10946,N_10885);
nand U11084 (N_11084,N_10947,N_10925);
nor U11085 (N_11085,N_10930,N_10978);
xnor U11086 (N_11086,N_10971,N_10919);
nand U11087 (N_11087,N_10932,N_10991);
xor U11088 (N_11088,N_10994,N_10963);
nor U11089 (N_11089,N_10897,N_10956);
nand U11090 (N_11090,N_10994,N_10923);
or U11091 (N_11091,N_10994,N_10952);
nand U11092 (N_11092,N_10948,N_10933);
and U11093 (N_11093,N_10901,N_10938);
nand U11094 (N_11094,N_10999,N_10985);
nand U11095 (N_11095,N_10888,N_10916);
nor U11096 (N_11096,N_10977,N_10877);
nand U11097 (N_11097,N_10937,N_10896);
xor U11098 (N_11098,N_10932,N_10995);
and U11099 (N_11099,N_10892,N_10876);
nand U11100 (N_11100,N_10969,N_10991);
or U11101 (N_11101,N_10915,N_10972);
and U11102 (N_11102,N_10922,N_10960);
nor U11103 (N_11103,N_10961,N_10933);
xor U11104 (N_11104,N_10959,N_10977);
nand U11105 (N_11105,N_10955,N_10877);
nor U11106 (N_11106,N_10994,N_10986);
xnor U11107 (N_11107,N_10896,N_10980);
nor U11108 (N_11108,N_10904,N_10990);
xnor U11109 (N_11109,N_10998,N_10991);
xnor U11110 (N_11110,N_10879,N_10949);
nor U11111 (N_11111,N_10999,N_10984);
nor U11112 (N_11112,N_10974,N_10942);
xor U11113 (N_11113,N_10958,N_10991);
nor U11114 (N_11114,N_10955,N_10882);
and U11115 (N_11115,N_10980,N_10909);
xnor U11116 (N_11116,N_10878,N_10877);
and U11117 (N_11117,N_10996,N_10923);
or U11118 (N_11118,N_10994,N_10992);
nand U11119 (N_11119,N_10955,N_10994);
nand U11120 (N_11120,N_10999,N_10923);
xnor U11121 (N_11121,N_10927,N_10952);
xor U11122 (N_11122,N_10893,N_10900);
or U11123 (N_11123,N_10950,N_10992);
or U11124 (N_11124,N_10899,N_10883);
nor U11125 (N_11125,N_11106,N_11103);
or U11126 (N_11126,N_11097,N_11049);
and U11127 (N_11127,N_11005,N_11083);
nand U11128 (N_11128,N_11002,N_11111);
nand U11129 (N_11129,N_11012,N_11124);
xor U11130 (N_11130,N_11088,N_11112);
nand U11131 (N_11131,N_11039,N_11122);
and U11132 (N_11132,N_11040,N_11009);
nor U11133 (N_11133,N_11030,N_11027);
nor U11134 (N_11134,N_11090,N_11067);
xor U11135 (N_11135,N_11000,N_11015);
xor U11136 (N_11136,N_11048,N_11072);
nand U11137 (N_11137,N_11007,N_11028);
xor U11138 (N_11138,N_11034,N_11063);
nand U11139 (N_11139,N_11047,N_11074);
and U11140 (N_11140,N_11080,N_11035);
nand U11141 (N_11141,N_11004,N_11084);
xor U11142 (N_11142,N_11033,N_11079);
and U11143 (N_11143,N_11056,N_11024);
or U11144 (N_11144,N_11026,N_11093);
nand U11145 (N_11145,N_11031,N_11116);
and U11146 (N_11146,N_11094,N_11019);
or U11147 (N_11147,N_11029,N_11041);
and U11148 (N_11148,N_11021,N_11082);
and U11149 (N_11149,N_11114,N_11022);
nor U11150 (N_11150,N_11046,N_11062);
nor U11151 (N_11151,N_11104,N_11081);
nor U11152 (N_11152,N_11098,N_11060);
xnor U11153 (N_11153,N_11011,N_11014);
nand U11154 (N_11154,N_11050,N_11107);
xnor U11155 (N_11155,N_11037,N_11078);
xnor U11156 (N_11156,N_11055,N_11010);
and U11157 (N_11157,N_11036,N_11095);
and U11158 (N_11158,N_11110,N_11073);
or U11159 (N_11159,N_11096,N_11101);
nor U11160 (N_11160,N_11059,N_11053);
xor U11161 (N_11161,N_11086,N_11087);
nor U11162 (N_11162,N_11085,N_11061);
or U11163 (N_11163,N_11077,N_11069);
xor U11164 (N_11164,N_11065,N_11051);
or U11165 (N_11165,N_11075,N_11091);
and U11166 (N_11166,N_11064,N_11044);
xnor U11167 (N_11167,N_11058,N_11017);
xnor U11168 (N_11168,N_11025,N_11117);
or U11169 (N_11169,N_11071,N_11045);
and U11170 (N_11170,N_11115,N_11052);
or U11171 (N_11171,N_11057,N_11054);
nand U11172 (N_11172,N_11032,N_11001);
and U11173 (N_11173,N_11038,N_11100);
and U11174 (N_11174,N_11121,N_11016);
nand U11175 (N_11175,N_11003,N_11076);
nand U11176 (N_11176,N_11008,N_11113);
xnor U11177 (N_11177,N_11118,N_11018);
nor U11178 (N_11178,N_11109,N_11006);
nand U11179 (N_11179,N_11023,N_11123);
and U11180 (N_11180,N_11099,N_11119);
and U11181 (N_11181,N_11013,N_11070);
nor U11182 (N_11182,N_11120,N_11020);
xnor U11183 (N_11183,N_11043,N_11092);
xor U11184 (N_11184,N_11108,N_11042);
nand U11185 (N_11185,N_11068,N_11066);
or U11186 (N_11186,N_11102,N_11089);
xor U11187 (N_11187,N_11105,N_11095);
xor U11188 (N_11188,N_11037,N_11094);
nand U11189 (N_11189,N_11053,N_11123);
or U11190 (N_11190,N_11068,N_11017);
nand U11191 (N_11191,N_11055,N_11080);
xnor U11192 (N_11192,N_11092,N_11018);
or U11193 (N_11193,N_11095,N_11026);
nand U11194 (N_11194,N_11090,N_11012);
xnor U11195 (N_11195,N_11117,N_11084);
or U11196 (N_11196,N_11086,N_11103);
xor U11197 (N_11197,N_11076,N_11101);
xor U11198 (N_11198,N_11002,N_11062);
nor U11199 (N_11199,N_11093,N_11040);
nand U11200 (N_11200,N_11082,N_11002);
or U11201 (N_11201,N_11025,N_11066);
and U11202 (N_11202,N_11035,N_11045);
xor U11203 (N_11203,N_11024,N_11095);
and U11204 (N_11204,N_11089,N_11082);
xnor U11205 (N_11205,N_11009,N_11073);
or U11206 (N_11206,N_11089,N_11050);
and U11207 (N_11207,N_11042,N_11053);
nand U11208 (N_11208,N_11001,N_11040);
nor U11209 (N_11209,N_11041,N_11108);
nor U11210 (N_11210,N_11012,N_11039);
xnor U11211 (N_11211,N_11049,N_11103);
xnor U11212 (N_11212,N_11059,N_11020);
nor U11213 (N_11213,N_11051,N_11000);
xor U11214 (N_11214,N_11083,N_11120);
nor U11215 (N_11215,N_11107,N_11057);
or U11216 (N_11216,N_11034,N_11044);
xor U11217 (N_11217,N_11107,N_11124);
nand U11218 (N_11218,N_11116,N_11105);
nand U11219 (N_11219,N_11106,N_11062);
or U11220 (N_11220,N_11023,N_11040);
nor U11221 (N_11221,N_11029,N_11052);
nand U11222 (N_11222,N_11043,N_11102);
and U11223 (N_11223,N_11066,N_11123);
xnor U11224 (N_11224,N_11065,N_11084);
xnor U11225 (N_11225,N_11021,N_11104);
or U11226 (N_11226,N_11057,N_11009);
and U11227 (N_11227,N_11079,N_11094);
nand U11228 (N_11228,N_11123,N_11082);
nand U11229 (N_11229,N_11119,N_11098);
and U11230 (N_11230,N_11048,N_11085);
and U11231 (N_11231,N_11058,N_11022);
and U11232 (N_11232,N_11079,N_11044);
and U11233 (N_11233,N_11017,N_11019);
nand U11234 (N_11234,N_11092,N_11119);
nor U11235 (N_11235,N_11072,N_11018);
and U11236 (N_11236,N_11101,N_11104);
xor U11237 (N_11237,N_11123,N_11017);
and U11238 (N_11238,N_11076,N_11111);
nor U11239 (N_11239,N_11068,N_11078);
nor U11240 (N_11240,N_11102,N_11123);
and U11241 (N_11241,N_11042,N_11002);
nand U11242 (N_11242,N_11034,N_11108);
nor U11243 (N_11243,N_11017,N_11114);
or U11244 (N_11244,N_11024,N_11090);
nand U11245 (N_11245,N_11047,N_11051);
xnor U11246 (N_11246,N_11028,N_11044);
xor U11247 (N_11247,N_11098,N_11004);
nand U11248 (N_11248,N_11002,N_11070);
or U11249 (N_11249,N_11076,N_11098);
nand U11250 (N_11250,N_11224,N_11206);
nand U11251 (N_11251,N_11241,N_11213);
xor U11252 (N_11252,N_11226,N_11199);
or U11253 (N_11253,N_11178,N_11209);
xnor U11254 (N_11254,N_11216,N_11182);
and U11255 (N_11255,N_11139,N_11181);
nor U11256 (N_11256,N_11239,N_11125);
xor U11257 (N_11257,N_11200,N_11208);
nor U11258 (N_11258,N_11203,N_11212);
or U11259 (N_11259,N_11165,N_11246);
nor U11260 (N_11260,N_11193,N_11196);
xor U11261 (N_11261,N_11233,N_11162);
nor U11262 (N_11262,N_11211,N_11231);
nand U11263 (N_11263,N_11167,N_11133);
or U11264 (N_11264,N_11190,N_11232);
and U11265 (N_11265,N_11187,N_11177);
xor U11266 (N_11266,N_11204,N_11126);
xor U11267 (N_11267,N_11130,N_11179);
or U11268 (N_11268,N_11159,N_11142);
nor U11269 (N_11269,N_11153,N_11192);
or U11270 (N_11270,N_11236,N_11152);
nor U11271 (N_11271,N_11248,N_11234);
nor U11272 (N_11272,N_11219,N_11147);
nand U11273 (N_11273,N_11180,N_11151);
or U11274 (N_11274,N_11128,N_11244);
nand U11275 (N_11275,N_11191,N_11225);
xor U11276 (N_11276,N_11235,N_11161);
nor U11277 (N_11277,N_11156,N_11205);
nand U11278 (N_11278,N_11145,N_11132);
or U11279 (N_11279,N_11210,N_11188);
or U11280 (N_11280,N_11154,N_11229);
and U11281 (N_11281,N_11172,N_11218);
nand U11282 (N_11282,N_11127,N_11217);
or U11283 (N_11283,N_11136,N_11131);
or U11284 (N_11284,N_11155,N_11148);
nor U11285 (N_11285,N_11168,N_11230);
nor U11286 (N_11286,N_11138,N_11242);
nand U11287 (N_11287,N_11198,N_11245);
and U11288 (N_11288,N_11158,N_11222);
nor U11289 (N_11289,N_11185,N_11174);
xnor U11290 (N_11290,N_11141,N_11135);
nand U11291 (N_11291,N_11137,N_11171);
nand U11292 (N_11292,N_11207,N_11183);
nor U11293 (N_11293,N_11129,N_11163);
and U11294 (N_11294,N_11164,N_11160);
nand U11295 (N_11295,N_11227,N_11146);
nor U11296 (N_11296,N_11134,N_11176);
xnor U11297 (N_11297,N_11157,N_11150);
nand U11298 (N_11298,N_11143,N_11240);
nand U11299 (N_11299,N_11223,N_11169);
nand U11300 (N_11300,N_11184,N_11215);
xnor U11301 (N_11301,N_11189,N_11140);
nor U11302 (N_11302,N_11144,N_11197);
and U11303 (N_11303,N_11149,N_11186);
and U11304 (N_11304,N_11228,N_11170);
nor U11305 (N_11305,N_11249,N_11220);
or U11306 (N_11306,N_11175,N_11166);
and U11307 (N_11307,N_11173,N_11194);
nand U11308 (N_11308,N_11195,N_11243);
or U11309 (N_11309,N_11237,N_11238);
nand U11310 (N_11310,N_11214,N_11221);
xor U11311 (N_11311,N_11202,N_11201);
nand U11312 (N_11312,N_11247,N_11182);
nor U11313 (N_11313,N_11139,N_11239);
xor U11314 (N_11314,N_11163,N_11156);
nor U11315 (N_11315,N_11181,N_11165);
nand U11316 (N_11316,N_11148,N_11242);
nor U11317 (N_11317,N_11213,N_11154);
nand U11318 (N_11318,N_11131,N_11145);
and U11319 (N_11319,N_11195,N_11143);
and U11320 (N_11320,N_11153,N_11189);
nor U11321 (N_11321,N_11249,N_11152);
nand U11322 (N_11322,N_11149,N_11137);
and U11323 (N_11323,N_11146,N_11204);
xnor U11324 (N_11324,N_11248,N_11233);
or U11325 (N_11325,N_11158,N_11175);
and U11326 (N_11326,N_11229,N_11188);
nand U11327 (N_11327,N_11209,N_11140);
xor U11328 (N_11328,N_11131,N_11162);
or U11329 (N_11329,N_11213,N_11162);
or U11330 (N_11330,N_11166,N_11156);
nand U11331 (N_11331,N_11191,N_11227);
or U11332 (N_11332,N_11130,N_11205);
or U11333 (N_11333,N_11206,N_11139);
or U11334 (N_11334,N_11209,N_11185);
xnor U11335 (N_11335,N_11140,N_11149);
nand U11336 (N_11336,N_11128,N_11207);
or U11337 (N_11337,N_11204,N_11131);
nand U11338 (N_11338,N_11191,N_11201);
xnor U11339 (N_11339,N_11243,N_11226);
xnor U11340 (N_11340,N_11167,N_11183);
xor U11341 (N_11341,N_11232,N_11220);
and U11342 (N_11342,N_11130,N_11220);
xnor U11343 (N_11343,N_11148,N_11210);
nor U11344 (N_11344,N_11245,N_11151);
nand U11345 (N_11345,N_11159,N_11214);
and U11346 (N_11346,N_11174,N_11198);
xnor U11347 (N_11347,N_11144,N_11139);
nand U11348 (N_11348,N_11149,N_11243);
nor U11349 (N_11349,N_11208,N_11202);
xor U11350 (N_11350,N_11241,N_11197);
xnor U11351 (N_11351,N_11207,N_11233);
and U11352 (N_11352,N_11182,N_11209);
nor U11353 (N_11353,N_11186,N_11226);
nor U11354 (N_11354,N_11232,N_11249);
or U11355 (N_11355,N_11225,N_11214);
and U11356 (N_11356,N_11236,N_11211);
or U11357 (N_11357,N_11224,N_11126);
nor U11358 (N_11358,N_11210,N_11238);
xnor U11359 (N_11359,N_11202,N_11158);
nor U11360 (N_11360,N_11142,N_11180);
and U11361 (N_11361,N_11227,N_11240);
nor U11362 (N_11362,N_11247,N_11206);
xor U11363 (N_11363,N_11174,N_11183);
nand U11364 (N_11364,N_11202,N_11144);
or U11365 (N_11365,N_11168,N_11191);
nor U11366 (N_11366,N_11200,N_11190);
nor U11367 (N_11367,N_11149,N_11181);
xor U11368 (N_11368,N_11180,N_11128);
and U11369 (N_11369,N_11141,N_11231);
or U11370 (N_11370,N_11242,N_11171);
nor U11371 (N_11371,N_11126,N_11207);
nor U11372 (N_11372,N_11212,N_11126);
xnor U11373 (N_11373,N_11229,N_11139);
nand U11374 (N_11374,N_11172,N_11153);
and U11375 (N_11375,N_11336,N_11350);
or U11376 (N_11376,N_11252,N_11274);
xnor U11377 (N_11377,N_11257,N_11288);
and U11378 (N_11378,N_11295,N_11308);
or U11379 (N_11379,N_11273,N_11359);
nor U11380 (N_11380,N_11309,N_11369);
or U11381 (N_11381,N_11267,N_11300);
xnor U11382 (N_11382,N_11301,N_11285);
nor U11383 (N_11383,N_11293,N_11271);
nand U11384 (N_11384,N_11298,N_11343);
nor U11385 (N_11385,N_11263,N_11357);
nand U11386 (N_11386,N_11280,N_11256);
nor U11387 (N_11387,N_11352,N_11290);
or U11388 (N_11388,N_11270,N_11344);
nand U11389 (N_11389,N_11327,N_11259);
nor U11390 (N_11390,N_11321,N_11340);
or U11391 (N_11391,N_11262,N_11348);
or U11392 (N_11392,N_11330,N_11260);
nor U11393 (N_11393,N_11349,N_11353);
and U11394 (N_11394,N_11341,N_11306);
nand U11395 (N_11395,N_11269,N_11304);
nor U11396 (N_11396,N_11307,N_11338);
or U11397 (N_11397,N_11335,N_11294);
xnor U11398 (N_11398,N_11323,N_11361);
nor U11399 (N_11399,N_11356,N_11342);
and U11400 (N_11400,N_11325,N_11326);
nor U11401 (N_11401,N_11358,N_11318);
nand U11402 (N_11402,N_11368,N_11302);
nand U11403 (N_11403,N_11251,N_11364);
nor U11404 (N_11404,N_11333,N_11360);
nor U11405 (N_11405,N_11347,N_11367);
nand U11406 (N_11406,N_11287,N_11265);
nor U11407 (N_11407,N_11272,N_11284);
xor U11408 (N_11408,N_11264,N_11310);
xor U11409 (N_11409,N_11339,N_11283);
nand U11410 (N_11410,N_11313,N_11355);
or U11411 (N_11411,N_11305,N_11261);
and U11412 (N_11412,N_11374,N_11250);
xor U11413 (N_11413,N_11282,N_11299);
or U11414 (N_11414,N_11315,N_11297);
or U11415 (N_11415,N_11289,N_11322);
and U11416 (N_11416,N_11320,N_11303);
or U11417 (N_11417,N_11253,N_11372);
xnor U11418 (N_11418,N_11316,N_11281);
and U11419 (N_11419,N_11268,N_11337);
or U11420 (N_11420,N_11311,N_11351);
nand U11421 (N_11421,N_11332,N_11334);
and U11422 (N_11422,N_11319,N_11275);
or U11423 (N_11423,N_11366,N_11317);
and U11424 (N_11424,N_11296,N_11278);
nand U11425 (N_11425,N_11354,N_11277);
nand U11426 (N_11426,N_11276,N_11373);
or U11427 (N_11427,N_11286,N_11255);
or U11428 (N_11428,N_11363,N_11329);
nor U11429 (N_11429,N_11312,N_11331);
xnor U11430 (N_11430,N_11370,N_11324);
nand U11431 (N_11431,N_11258,N_11292);
nand U11432 (N_11432,N_11314,N_11362);
or U11433 (N_11433,N_11346,N_11345);
nor U11434 (N_11434,N_11291,N_11371);
nand U11435 (N_11435,N_11266,N_11279);
and U11436 (N_11436,N_11365,N_11328);
and U11437 (N_11437,N_11254,N_11333);
xor U11438 (N_11438,N_11261,N_11332);
and U11439 (N_11439,N_11271,N_11279);
xnor U11440 (N_11440,N_11314,N_11334);
nand U11441 (N_11441,N_11258,N_11302);
nand U11442 (N_11442,N_11316,N_11340);
xor U11443 (N_11443,N_11267,N_11367);
or U11444 (N_11444,N_11292,N_11287);
xor U11445 (N_11445,N_11315,N_11371);
nand U11446 (N_11446,N_11312,N_11296);
nand U11447 (N_11447,N_11266,N_11303);
or U11448 (N_11448,N_11339,N_11329);
nand U11449 (N_11449,N_11305,N_11335);
nor U11450 (N_11450,N_11265,N_11266);
nand U11451 (N_11451,N_11374,N_11286);
and U11452 (N_11452,N_11275,N_11355);
nor U11453 (N_11453,N_11333,N_11281);
nand U11454 (N_11454,N_11275,N_11341);
and U11455 (N_11455,N_11256,N_11302);
xnor U11456 (N_11456,N_11292,N_11368);
nand U11457 (N_11457,N_11313,N_11327);
and U11458 (N_11458,N_11293,N_11326);
and U11459 (N_11459,N_11263,N_11352);
xor U11460 (N_11460,N_11311,N_11372);
or U11461 (N_11461,N_11302,N_11301);
nor U11462 (N_11462,N_11340,N_11330);
nand U11463 (N_11463,N_11317,N_11347);
xor U11464 (N_11464,N_11325,N_11271);
nor U11465 (N_11465,N_11316,N_11326);
and U11466 (N_11466,N_11268,N_11346);
or U11467 (N_11467,N_11297,N_11316);
nand U11468 (N_11468,N_11262,N_11275);
nor U11469 (N_11469,N_11354,N_11349);
nor U11470 (N_11470,N_11271,N_11258);
nand U11471 (N_11471,N_11295,N_11301);
and U11472 (N_11472,N_11360,N_11295);
or U11473 (N_11473,N_11259,N_11306);
and U11474 (N_11474,N_11329,N_11298);
nor U11475 (N_11475,N_11263,N_11369);
and U11476 (N_11476,N_11279,N_11265);
xor U11477 (N_11477,N_11298,N_11302);
nand U11478 (N_11478,N_11360,N_11297);
or U11479 (N_11479,N_11269,N_11325);
nand U11480 (N_11480,N_11324,N_11296);
xnor U11481 (N_11481,N_11358,N_11344);
xnor U11482 (N_11482,N_11253,N_11297);
nor U11483 (N_11483,N_11347,N_11293);
xor U11484 (N_11484,N_11343,N_11334);
nor U11485 (N_11485,N_11340,N_11261);
nand U11486 (N_11486,N_11250,N_11331);
and U11487 (N_11487,N_11300,N_11301);
xor U11488 (N_11488,N_11269,N_11347);
xnor U11489 (N_11489,N_11356,N_11368);
or U11490 (N_11490,N_11289,N_11255);
xor U11491 (N_11491,N_11354,N_11288);
or U11492 (N_11492,N_11372,N_11315);
xor U11493 (N_11493,N_11320,N_11262);
and U11494 (N_11494,N_11345,N_11299);
or U11495 (N_11495,N_11351,N_11335);
or U11496 (N_11496,N_11301,N_11308);
and U11497 (N_11497,N_11374,N_11364);
and U11498 (N_11498,N_11298,N_11348);
and U11499 (N_11499,N_11292,N_11267);
or U11500 (N_11500,N_11438,N_11478);
and U11501 (N_11501,N_11405,N_11460);
nand U11502 (N_11502,N_11434,N_11482);
and U11503 (N_11503,N_11446,N_11413);
or U11504 (N_11504,N_11393,N_11427);
xor U11505 (N_11505,N_11467,N_11382);
xor U11506 (N_11506,N_11429,N_11403);
xor U11507 (N_11507,N_11406,N_11465);
or U11508 (N_11508,N_11471,N_11395);
nand U11509 (N_11509,N_11417,N_11424);
nand U11510 (N_11510,N_11383,N_11481);
and U11511 (N_11511,N_11414,N_11411);
nor U11512 (N_11512,N_11420,N_11499);
xnor U11513 (N_11513,N_11404,N_11483);
xnor U11514 (N_11514,N_11387,N_11394);
nand U11515 (N_11515,N_11407,N_11380);
nand U11516 (N_11516,N_11397,N_11496);
or U11517 (N_11517,N_11445,N_11491);
nand U11518 (N_11518,N_11477,N_11443);
or U11519 (N_11519,N_11488,N_11435);
or U11520 (N_11520,N_11418,N_11449);
and U11521 (N_11521,N_11480,N_11390);
nand U11522 (N_11522,N_11389,N_11400);
nand U11523 (N_11523,N_11379,N_11437);
nand U11524 (N_11524,N_11410,N_11448);
nand U11525 (N_11525,N_11422,N_11470);
nor U11526 (N_11526,N_11396,N_11384);
xor U11527 (N_11527,N_11442,N_11469);
nor U11528 (N_11528,N_11428,N_11416);
nor U11529 (N_11529,N_11388,N_11475);
xnor U11530 (N_11530,N_11433,N_11408);
nand U11531 (N_11531,N_11494,N_11402);
and U11532 (N_11532,N_11462,N_11450);
nor U11533 (N_11533,N_11484,N_11493);
or U11534 (N_11534,N_11485,N_11455);
nor U11535 (N_11535,N_11412,N_11440);
xnor U11536 (N_11536,N_11430,N_11498);
nand U11537 (N_11537,N_11425,N_11386);
nand U11538 (N_11538,N_11376,N_11495);
xor U11539 (N_11539,N_11399,N_11375);
and U11540 (N_11540,N_11401,N_11432);
xor U11541 (N_11541,N_11468,N_11447);
or U11542 (N_11542,N_11453,N_11439);
xnor U11543 (N_11543,N_11444,N_11385);
or U11544 (N_11544,N_11466,N_11441);
or U11545 (N_11545,N_11489,N_11474);
nor U11546 (N_11546,N_11486,N_11454);
nor U11547 (N_11547,N_11426,N_11391);
nand U11548 (N_11548,N_11459,N_11473);
nor U11549 (N_11549,N_11431,N_11492);
and U11550 (N_11550,N_11381,N_11451);
nand U11551 (N_11551,N_11419,N_11479);
or U11552 (N_11552,N_11415,N_11487);
or U11553 (N_11553,N_11458,N_11490);
nand U11554 (N_11554,N_11456,N_11378);
or U11555 (N_11555,N_11464,N_11409);
xor U11556 (N_11556,N_11421,N_11457);
xor U11557 (N_11557,N_11398,N_11392);
nor U11558 (N_11558,N_11472,N_11436);
xor U11559 (N_11559,N_11463,N_11476);
and U11560 (N_11560,N_11377,N_11497);
or U11561 (N_11561,N_11452,N_11461);
and U11562 (N_11562,N_11423,N_11387);
and U11563 (N_11563,N_11459,N_11464);
nand U11564 (N_11564,N_11484,N_11384);
nand U11565 (N_11565,N_11465,N_11440);
or U11566 (N_11566,N_11491,N_11424);
nor U11567 (N_11567,N_11499,N_11454);
nand U11568 (N_11568,N_11462,N_11391);
and U11569 (N_11569,N_11474,N_11430);
xnor U11570 (N_11570,N_11378,N_11382);
or U11571 (N_11571,N_11420,N_11390);
and U11572 (N_11572,N_11383,N_11457);
nor U11573 (N_11573,N_11377,N_11420);
nand U11574 (N_11574,N_11497,N_11430);
and U11575 (N_11575,N_11495,N_11473);
nor U11576 (N_11576,N_11472,N_11480);
nand U11577 (N_11577,N_11468,N_11395);
xor U11578 (N_11578,N_11411,N_11375);
nor U11579 (N_11579,N_11393,N_11418);
xnor U11580 (N_11580,N_11418,N_11479);
nor U11581 (N_11581,N_11478,N_11468);
nor U11582 (N_11582,N_11487,N_11435);
and U11583 (N_11583,N_11438,N_11376);
or U11584 (N_11584,N_11456,N_11414);
nand U11585 (N_11585,N_11429,N_11488);
or U11586 (N_11586,N_11424,N_11489);
nor U11587 (N_11587,N_11379,N_11446);
and U11588 (N_11588,N_11436,N_11498);
or U11589 (N_11589,N_11453,N_11419);
or U11590 (N_11590,N_11434,N_11413);
nor U11591 (N_11591,N_11497,N_11493);
and U11592 (N_11592,N_11433,N_11476);
or U11593 (N_11593,N_11474,N_11440);
xnor U11594 (N_11594,N_11397,N_11385);
and U11595 (N_11595,N_11458,N_11464);
or U11596 (N_11596,N_11462,N_11479);
nand U11597 (N_11597,N_11476,N_11483);
or U11598 (N_11598,N_11492,N_11478);
and U11599 (N_11599,N_11498,N_11445);
nor U11600 (N_11600,N_11393,N_11459);
or U11601 (N_11601,N_11476,N_11408);
or U11602 (N_11602,N_11469,N_11459);
nand U11603 (N_11603,N_11468,N_11412);
or U11604 (N_11604,N_11414,N_11481);
nand U11605 (N_11605,N_11458,N_11414);
xor U11606 (N_11606,N_11378,N_11444);
and U11607 (N_11607,N_11479,N_11474);
and U11608 (N_11608,N_11444,N_11397);
nand U11609 (N_11609,N_11482,N_11389);
nand U11610 (N_11610,N_11387,N_11432);
nand U11611 (N_11611,N_11498,N_11471);
or U11612 (N_11612,N_11479,N_11395);
xnor U11613 (N_11613,N_11388,N_11480);
nor U11614 (N_11614,N_11480,N_11450);
and U11615 (N_11615,N_11483,N_11387);
or U11616 (N_11616,N_11396,N_11379);
nand U11617 (N_11617,N_11447,N_11481);
nand U11618 (N_11618,N_11394,N_11460);
or U11619 (N_11619,N_11379,N_11451);
nor U11620 (N_11620,N_11425,N_11471);
and U11621 (N_11621,N_11455,N_11388);
xnor U11622 (N_11622,N_11462,N_11423);
and U11623 (N_11623,N_11484,N_11417);
nor U11624 (N_11624,N_11380,N_11386);
nand U11625 (N_11625,N_11578,N_11624);
xor U11626 (N_11626,N_11620,N_11576);
nor U11627 (N_11627,N_11536,N_11512);
xnor U11628 (N_11628,N_11586,N_11545);
nand U11629 (N_11629,N_11503,N_11525);
nor U11630 (N_11630,N_11584,N_11605);
nor U11631 (N_11631,N_11534,N_11521);
nand U11632 (N_11632,N_11526,N_11532);
xor U11633 (N_11633,N_11509,N_11592);
and U11634 (N_11634,N_11587,N_11535);
or U11635 (N_11635,N_11611,N_11504);
xor U11636 (N_11636,N_11610,N_11612);
and U11637 (N_11637,N_11569,N_11539);
xnor U11638 (N_11638,N_11585,N_11523);
or U11639 (N_11639,N_11538,N_11554);
xnor U11640 (N_11640,N_11608,N_11597);
or U11641 (N_11641,N_11547,N_11562);
xnor U11642 (N_11642,N_11552,N_11515);
and U11643 (N_11643,N_11550,N_11507);
xor U11644 (N_11644,N_11517,N_11575);
nor U11645 (N_11645,N_11528,N_11533);
xor U11646 (N_11646,N_11500,N_11513);
nand U11647 (N_11647,N_11582,N_11524);
and U11648 (N_11648,N_11542,N_11516);
nor U11649 (N_11649,N_11558,N_11591);
and U11650 (N_11650,N_11589,N_11604);
nor U11651 (N_11651,N_11501,N_11601);
or U11652 (N_11652,N_11595,N_11622);
or U11653 (N_11653,N_11564,N_11508);
xor U11654 (N_11654,N_11561,N_11556);
or U11655 (N_11655,N_11615,N_11510);
nor U11656 (N_11656,N_11520,N_11583);
nor U11657 (N_11657,N_11544,N_11621);
and U11658 (N_11658,N_11567,N_11598);
xnor U11659 (N_11659,N_11505,N_11566);
and U11660 (N_11660,N_11572,N_11593);
nor U11661 (N_11661,N_11580,N_11609);
nand U11662 (N_11662,N_11581,N_11537);
nor U11663 (N_11663,N_11519,N_11599);
xor U11664 (N_11664,N_11514,N_11596);
nor U11665 (N_11665,N_11518,N_11590);
and U11666 (N_11666,N_11588,N_11619);
nand U11667 (N_11667,N_11541,N_11614);
nand U11668 (N_11668,N_11502,N_11570);
and U11669 (N_11669,N_11565,N_11553);
or U11670 (N_11670,N_11549,N_11522);
and U11671 (N_11671,N_11574,N_11616);
and U11672 (N_11672,N_11527,N_11579);
xnor U11673 (N_11673,N_11613,N_11623);
xnor U11674 (N_11674,N_11594,N_11577);
and U11675 (N_11675,N_11560,N_11573);
xor U11676 (N_11676,N_11563,N_11531);
or U11677 (N_11677,N_11602,N_11543);
or U11678 (N_11678,N_11548,N_11571);
and U11679 (N_11679,N_11557,N_11607);
xor U11680 (N_11680,N_11618,N_11606);
nor U11681 (N_11681,N_11530,N_11511);
and U11682 (N_11682,N_11603,N_11540);
and U11683 (N_11683,N_11551,N_11617);
nand U11684 (N_11684,N_11568,N_11555);
and U11685 (N_11685,N_11600,N_11559);
xnor U11686 (N_11686,N_11546,N_11506);
or U11687 (N_11687,N_11529,N_11613);
or U11688 (N_11688,N_11511,N_11615);
nor U11689 (N_11689,N_11610,N_11623);
and U11690 (N_11690,N_11567,N_11515);
or U11691 (N_11691,N_11578,N_11509);
nor U11692 (N_11692,N_11565,N_11618);
nand U11693 (N_11693,N_11537,N_11576);
xor U11694 (N_11694,N_11553,N_11576);
xor U11695 (N_11695,N_11620,N_11551);
or U11696 (N_11696,N_11544,N_11527);
nor U11697 (N_11697,N_11607,N_11582);
or U11698 (N_11698,N_11527,N_11574);
or U11699 (N_11699,N_11502,N_11501);
or U11700 (N_11700,N_11523,N_11564);
or U11701 (N_11701,N_11606,N_11505);
nand U11702 (N_11702,N_11597,N_11623);
nor U11703 (N_11703,N_11574,N_11518);
or U11704 (N_11704,N_11556,N_11584);
and U11705 (N_11705,N_11553,N_11546);
or U11706 (N_11706,N_11533,N_11511);
and U11707 (N_11707,N_11551,N_11587);
xor U11708 (N_11708,N_11538,N_11562);
and U11709 (N_11709,N_11534,N_11602);
and U11710 (N_11710,N_11576,N_11503);
xnor U11711 (N_11711,N_11546,N_11531);
nand U11712 (N_11712,N_11547,N_11514);
nand U11713 (N_11713,N_11555,N_11593);
xor U11714 (N_11714,N_11529,N_11578);
nand U11715 (N_11715,N_11579,N_11567);
nand U11716 (N_11716,N_11612,N_11568);
or U11717 (N_11717,N_11608,N_11535);
nor U11718 (N_11718,N_11509,N_11600);
xor U11719 (N_11719,N_11500,N_11544);
nand U11720 (N_11720,N_11605,N_11587);
nor U11721 (N_11721,N_11528,N_11504);
or U11722 (N_11722,N_11545,N_11503);
or U11723 (N_11723,N_11564,N_11519);
nor U11724 (N_11724,N_11562,N_11566);
nor U11725 (N_11725,N_11567,N_11501);
or U11726 (N_11726,N_11598,N_11600);
or U11727 (N_11727,N_11525,N_11519);
or U11728 (N_11728,N_11521,N_11542);
or U11729 (N_11729,N_11505,N_11605);
nand U11730 (N_11730,N_11548,N_11514);
or U11731 (N_11731,N_11608,N_11574);
nand U11732 (N_11732,N_11543,N_11533);
nor U11733 (N_11733,N_11624,N_11552);
nor U11734 (N_11734,N_11579,N_11542);
nor U11735 (N_11735,N_11506,N_11597);
or U11736 (N_11736,N_11562,N_11611);
xnor U11737 (N_11737,N_11583,N_11555);
and U11738 (N_11738,N_11511,N_11518);
xor U11739 (N_11739,N_11615,N_11590);
nor U11740 (N_11740,N_11563,N_11605);
xnor U11741 (N_11741,N_11515,N_11557);
nor U11742 (N_11742,N_11608,N_11553);
xnor U11743 (N_11743,N_11607,N_11511);
nor U11744 (N_11744,N_11592,N_11528);
nor U11745 (N_11745,N_11514,N_11508);
or U11746 (N_11746,N_11572,N_11587);
xor U11747 (N_11747,N_11550,N_11508);
nand U11748 (N_11748,N_11532,N_11560);
and U11749 (N_11749,N_11540,N_11601);
xor U11750 (N_11750,N_11712,N_11747);
xor U11751 (N_11751,N_11729,N_11745);
nor U11752 (N_11752,N_11727,N_11661);
nand U11753 (N_11753,N_11679,N_11673);
nand U11754 (N_11754,N_11692,N_11701);
nand U11755 (N_11755,N_11658,N_11640);
nor U11756 (N_11756,N_11654,N_11741);
or U11757 (N_11757,N_11703,N_11651);
xnor U11758 (N_11758,N_11686,N_11704);
xnor U11759 (N_11759,N_11698,N_11631);
and U11760 (N_11760,N_11726,N_11664);
or U11761 (N_11761,N_11714,N_11718);
xor U11762 (N_11762,N_11665,N_11713);
xor U11763 (N_11763,N_11700,N_11743);
and U11764 (N_11764,N_11715,N_11632);
nor U11765 (N_11765,N_11737,N_11643);
xor U11766 (N_11766,N_11724,N_11742);
nor U11767 (N_11767,N_11630,N_11675);
or U11768 (N_11768,N_11716,N_11668);
nor U11769 (N_11769,N_11634,N_11659);
nand U11770 (N_11770,N_11705,N_11663);
nor U11771 (N_11771,N_11655,N_11689);
nand U11772 (N_11772,N_11674,N_11633);
nand U11773 (N_11773,N_11721,N_11735);
xor U11774 (N_11774,N_11738,N_11736);
xnor U11775 (N_11775,N_11676,N_11670);
nor U11776 (N_11776,N_11642,N_11707);
or U11777 (N_11777,N_11723,N_11626);
or U11778 (N_11778,N_11667,N_11652);
and U11779 (N_11779,N_11711,N_11706);
or U11780 (N_11780,N_11656,N_11641);
nor U11781 (N_11781,N_11681,N_11746);
or U11782 (N_11782,N_11683,N_11671);
xnor U11783 (N_11783,N_11709,N_11625);
nor U11784 (N_11784,N_11722,N_11694);
nor U11785 (N_11785,N_11720,N_11734);
or U11786 (N_11786,N_11628,N_11696);
or U11787 (N_11787,N_11740,N_11647);
and U11788 (N_11788,N_11744,N_11639);
and U11789 (N_11789,N_11645,N_11646);
and U11790 (N_11790,N_11672,N_11725);
and U11791 (N_11791,N_11660,N_11748);
xor U11792 (N_11792,N_11731,N_11691);
nand U11793 (N_11793,N_11739,N_11695);
or U11794 (N_11794,N_11680,N_11693);
nand U11795 (N_11795,N_11650,N_11719);
or U11796 (N_11796,N_11697,N_11636);
xor U11797 (N_11797,N_11708,N_11684);
or U11798 (N_11798,N_11728,N_11688);
nand U11799 (N_11799,N_11648,N_11687);
and U11800 (N_11800,N_11657,N_11678);
nand U11801 (N_11801,N_11717,N_11749);
or U11802 (N_11802,N_11710,N_11635);
and U11803 (N_11803,N_11644,N_11637);
nor U11804 (N_11804,N_11732,N_11649);
nor U11805 (N_11805,N_11699,N_11682);
xnor U11806 (N_11806,N_11638,N_11627);
nand U11807 (N_11807,N_11653,N_11629);
nand U11808 (N_11808,N_11690,N_11730);
xnor U11809 (N_11809,N_11702,N_11666);
xor U11810 (N_11810,N_11685,N_11662);
or U11811 (N_11811,N_11669,N_11733);
or U11812 (N_11812,N_11677,N_11638);
xnor U11813 (N_11813,N_11705,N_11686);
and U11814 (N_11814,N_11679,N_11677);
and U11815 (N_11815,N_11664,N_11657);
nand U11816 (N_11816,N_11639,N_11719);
nand U11817 (N_11817,N_11626,N_11649);
or U11818 (N_11818,N_11667,N_11681);
nand U11819 (N_11819,N_11727,N_11682);
nand U11820 (N_11820,N_11659,N_11651);
and U11821 (N_11821,N_11743,N_11703);
and U11822 (N_11822,N_11634,N_11653);
or U11823 (N_11823,N_11647,N_11733);
or U11824 (N_11824,N_11699,N_11693);
nor U11825 (N_11825,N_11671,N_11637);
or U11826 (N_11826,N_11707,N_11634);
or U11827 (N_11827,N_11657,N_11659);
nand U11828 (N_11828,N_11672,N_11659);
nor U11829 (N_11829,N_11694,N_11709);
xnor U11830 (N_11830,N_11662,N_11646);
nand U11831 (N_11831,N_11744,N_11659);
xor U11832 (N_11832,N_11638,N_11685);
xnor U11833 (N_11833,N_11686,N_11732);
and U11834 (N_11834,N_11744,N_11745);
or U11835 (N_11835,N_11693,N_11746);
or U11836 (N_11836,N_11703,N_11748);
and U11837 (N_11837,N_11681,N_11698);
nand U11838 (N_11838,N_11635,N_11669);
and U11839 (N_11839,N_11732,N_11725);
xor U11840 (N_11840,N_11708,N_11692);
xnor U11841 (N_11841,N_11644,N_11640);
nor U11842 (N_11842,N_11700,N_11722);
nor U11843 (N_11843,N_11742,N_11748);
nor U11844 (N_11844,N_11744,N_11702);
nand U11845 (N_11845,N_11659,N_11707);
xnor U11846 (N_11846,N_11643,N_11688);
nand U11847 (N_11847,N_11732,N_11704);
or U11848 (N_11848,N_11675,N_11730);
or U11849 (N_11849,N_11654,N_11669);
nor U11850 (N_11850,N_11664,N_11633);
and U11851 (N_11851,N_11656,N_11678);
and U11852 (N_11852,N_11678,N_11723);
and U11853 (N_11853,N_11716,N_11733);
xor U11854 (N_11854,N_11695,N_11649);
xnor U11855 (N_11855,N_11721,N_11748);
xnor U11856 (N_11856,N_11669,N_11651);
nand U11857 (N_11857,N_11663,N_11667);
and U11858 (N_11858,N_11743,N_11689);
or U11859 (N_11859,N_11631,N_11666);
xnor U11860 (N_11860,N_11701,N_11642);
xnor U11861 (N_11861,N_11736,N_11655);
or U11862 (N_11862,N_11685,N_11697);
and U11863 (N_11863,N_11637,N_11730);
nor U11864 (N_11864,N_11643,N_11631);
nor U11865 (N_11865,N_11646,N_11713);
nand U11866 (N_11866,N_11716,N_11707);
nor U11867 (N_11867,N_11710,N_11741);
nand U11868 (N_11868,N_11733,N_11748);
and U11869 (N_11869,N_11639,N_11642);
nand U11870 (N_11870,N_11742,N_11729);
xor U11871 (N_11871,N_11629,N_11690);
nor U11872 (N_11872,N_11712,N_11647);
and U11873 (N_11873,N_11639,N_11688);
or U11874 (N_11874,N_11653,N_11689);
and U11875 (N_11875,N_11826,N_11781);
nor U11876 (N_11876,N_11842,N_11863);
xor U11877 (N_11877,N_11773,N_11866);
nand U11878 (N_11878,N_11852,N_11869);
nor U11879 (N_11879,N_11823,N_11831);
xor U11880 (N_11880,N_11828,N_11797);
or U11881 (N_11881,N_11815,N_11820);
or U11882 (N_11882,N_11832,N_11859);
nor U11883 (N_11883,N_11854,N_11760);
nor U11884 (N_11884,N_11814,N_11864);
xor U11885 (N_11885,N_11771,N_11766);
nand U11886 (N_11886,N_11867,N_11801);
nor U11887 (N_11887,N_11779,N_11834);
nor U11888 (N_11888,N_11767,N_11861);
or U11889 (N_11889,N_11868,N_11860);
nor U11890 (N_11890,N_11757,N_11786);
or U11891 (N_11891,N_11802,N_11870);
xnor U11892 (N_11892,N_11783,N_11873);
or U11893 (N_11893,N_11787,N_11849);
or U11894 (N_11894,N_11857,N_11793);
xnor U11895 (N_11895,N_11764,N_11838);
and U11896 (N_11896,N_11821,N_11794);
or U11897 (N_11897,N_11853,N_11872);
xor U11898 (N_11898,N_11813,N_11829);
xor U11899 (N_11899,N_11795,N_11843);
nand U11900 (N_11900,N_11776,N_11761);
and U11901 (N_11901,N_11777,N_11855);
and U11902 (N_11902,N_11789,N_11839);
nor U11903 (N_11903,N_11811,N_11835);
nor U11904 (N_11904,N_11871,N_11753);
nor U11905 (N_11905,N_11807,N_11769);
nor U11906 (N_11906,N_11763,N_11837);
or U11907 (N_11907,N_11816,N_11822);
nor U11908 (N_11908,N_11836,N_11780);
nor U11909 (N_11909,N_11841,N_11812);
nor U11910 (N_11910,N_11790,N_11840);
xor U11911 (N_11911,N_11818,N_11848);
nor U11912 (N_11912,N_11874,N_11799);
nand U11913 (N_11913,N_11845,N_11800);
xor U11914 (N_11914,N_11778,N_11782);
nand U11915 (N_11915,N_11770,N_11851);
and U11916 (N_11916,N_11756,N_11844);
nand U11917 (N_11917,N_11850,N_11755);
xor U11918 (N_11918,N_11752,N_11754);
or U11919 (N_11919,N_11751,N_11804);
and U11920 (N_11920,N_11824,N_11827);
nand U11921 (N_11921,N_11862,N_11808);
and U11922 (N_11922,N_11774,N_11784);
xor U11923 (N_11923,N_11825,N_11759);
or U11924 (N_11924,N_11847,N_11846);
or U11925 (N_11925,N_11762,N_11803);
nand U11926 (N_11926,N_11791,N_11768);
xnor U11927 (N_11927,N_11788,N_11830);
and U11928 (N_11928,N_11792,N_11858);
xor U11929 (N_11929,N_11796,N_11772);
xnor U11930 (N_11930,N_11785,N_11765);
xor U11931 (N_11931,N_11750,N_11833);
and U11932 (N_11932,N_11806,N_11758);
nand U11933 (N_11933,N_11810,N_11775);
or U11934 (N_11934,N_11819,N_11798);
or U11935 (N_11935,N_11805,N_11817);
nor U11936 (N_11936,N_11856,N_11865);
and U11937 (N_11937,N_11809,N_11757);
and U11938 (N_11938,N_11821,N_11772);
or U11939 (N_11939,N_11784,N_11838);
and U11940 (N_11940,N_11773,N_11783);
and U11941 (N_11941,N_11812,N_11800);
nor U11942 (N_11942,N_11841,N_11752);
xor U11943 (N_11943,N_11776,N_11762);
or U11944 (N_11944,N_11759,N_11817);
and U11945 (N_11945,N_11798,N_11815);
xor U11946 (N_11946,N_11816,N_11844);
nand U11947 (N_11947,N_11777,N_11829);
xnor U11948 (N_11948,N_11828,N_11776);
nor U11949 (N_11949,N_11785,N_11759);
xor U11950 (N_11950,N_11821,N_11764);
or U11951 (N_11951,N_11844,N_11788);
nor U11952 (N_11952,N_11834,N_11755);
and U11953 (N_11953,N_11753,N_11799);
nand U11954 (N_11954,N_11859,N_11853);
nor U11955 (N_11955,N_11792,N_11794);
and U11956 (N_11956,N_11807,N_11852);
nand U11957 (N_11957,N_11788,N_11786);
or U11958 (N_11958,N_11804,N_11773);
or U11959 (N_11959,N_11856,N_11759);
nor U11960 (N_11960,N_11811,N_11867);
nand U11961 (N_11961,N_11844,N_11801);
and U11962 (N_11962,N_11773,N_11757);
xnor U11963 (N_11963,N_11759,N_11846);
nor U11964 (N_11964,N_11859,N_11780);
and U11965 (N_11965,N_11811,N_11866);
or U11966 (N_11966,N_11812,N_11815);
xor U11967 (N_11967,N_11854,N_11809);
or U11968 (N_11968,N_11851,N_11804);
xor U11969 (N_11969,N_11785,N_11789);
nor U11970 (N_11970,N_11753,N_11794);
nor U11971 (N_11971,N_11843,N_11847);
xnor U11972 (N_11972,N_11872,N_11816);
xnor U11973 (N_11973,N_11828,N_11813);
nor U11974 (N_11974,N_11789,N_11768);
nor U11975 (N_11975,N_11793,N_11814);
nand U11976 (N_11976,N_11872,N_11848);
and U11977 (N_11977,N_11782,N_11859);
xnor U11978 (N_11978,N_11777,N_11771);
nand U11979 (N_11979,N_11815,N_11785);
xnor U11980 (N_11980,N_11796,N_11866);
xnor U11981 (N_11981,N_11764,N_11844);
nor U11982 (N_11982,N_11781,N_11870);
nand U11983 (N_11983,N_11841,N_11865);
nor U11984 (N_11984,N_11853,N_11854);
or U11985 (N_11985,N_11849,N_11843);
nor U11986 (N_11986,N_11759,N_11847);
xnor U11987 (N_11987,N_11862,N_11856);
and U11988 (N_11988,N_11750,N_11791);
and U11989 (N_11989,N_11854,N_11812);
and U11990 (N_11990,N_11856,N_11786);
and U11991 (N_11991,N_11800,N_11853);
and U11992 (N_11992,N_11863,N_11818);
or U11993 (N_11993,N_11819,N_11830);
xnor U11994 (N_11994,N_11791,N_11760);
nor U11995 (N_11995,N_11795,N_11790);
or U11996 (N_11996,N_11777,N_11845);
xnor U11997 (N_11997,N_11753,N_11771);
and U11998 (N_11998,N_11850,N_11823);
or U11999 (N_11999,N_11824,N_11834);
nand U12000 (N_12000,N_11967,N_11990);
or U12001 (N_12001,N_11942,N_11908);
or U12002 (N_12002,N_11906,N_11935);
and U12003 (N_12003,N_11950,N_11954);
and U12004 (N_12004,N_11897,N_11986);
and U12005 (N_12005,N_11925,N_11888);
or U12006 (N_12006,N_11907,N_11877);
and U12007 (N_12007,N_11900,N_11885);
and U12008 (N_12008,N_11914,N_11997);
nand U12009 (N_12009,N_11875,N_11913);
nor U12010 (N_12010,N_11893,N_11890);
nand U12011 (N_12011,N_11947,N_11994);
and U12012 (N_12012,N_11878,N_11936);
and U12013 (N_12013,N_11971,N_11983);
nand U12014 (N_12014,N_11923,N_11985);
nor U12015 (N_12015,N_11970,N_11987);
or U12016 (N_12016,N_11937,N_11951);
nor U12017 (N_12017,N_11980,N_11892);
and U12018 (N_12018,N_11920,N_11880);
nor U12019 (N_12019,N_11895,N_11918);
or U12020 (N_12020,N_11969,N_11992);
xnor U12021 (N_12021,N_11904,N_11917);
and U12022 (N_12022,N_11924,N_11929);
xor U12023 (N_12023,N_11887,N_11926);
nor U12024 (N_12024,N_11968,N_11958);
xor U12025 (N_12025,N_11910,N_11953);
nand U12026 (N_12026,N_11981,N_11955);
and U12027 (N_12027,N_11965,N_11934);
or U12028 (N_12028,N_11945,N_11933);
or U12029 (N_12029,N_11995,N_11889);
nand U12030 (N_12030,N_11876,N_11886);
and U12031 (N_12031,N_11999,N_11972);
nand U12032 (N_12032,N_11941,N_11949);
and U12033 (N_12033,N_11978,N_11946);
nor U12034 (N_12034,N_11989,N_11976);
and U12035 (N_12035,N_11993,N_11905);
or U12036 (N_12036,N_11931,N_11884);
nand U12037 (N_12037,N_11939,N_11960);
xnor U12038 (N_12038,N_11991,N_11883);
and U12039 (N_12039,N_11961,N_11881);
nand U12040 (N_12040,N_11956,N_11952);
and U12041 (N_12041,N_11975,N_11921);
nand U12042 (N_12042,N_11916,N_11938);
nor U12043 (N_12043,N_11996,N_11898);
xnor U12044 (N_12044,N_11928,N_11932);
nor U12045 (N_12045,N_11964,N_11977);
nand U12046 (N_12046,N_11943,N_11982);
or U12047 (N_12047,N_11922,N_11963);
nand U12048 (N_12048,N_11948,N_11915);
nand U12049 (N_12049,N_11940,N_11901);
xnor U12050 (N_12050,N_11894,N_11909);
nor U12051 (N_12051,N_11988,N_11930);
or U12052 (N_12052,N_11962,N_11902);
or U12053 (N_12053,N_11903,N_11912);
nand U12054 (N_12054,N_11998,N_11896);
nor U12055 (N_12055,N_11984,N_11919);
xor U12056 (N_12056,N_11974,N_11973);
or U12057 (N_12057,N_11899,N_11959);
nor U12058 (N_12058,N_11979,N_11882);
or U12059 (N_12059,N_11891,N_11944);
or U12060 (N_12060,N_11911,N_11879);
nand U12061 (N_12061,N_11927,N_11957);
or U12062 (N_12062,N_11966,N_11956);
xnor U12063 (N_12063,N_11876,N_11937);
xnor U12064 (N_12064,N_11934,N_11994);
xor U12065 (N_12065,N_11907,N_11893);
nand U12066 (N_12066,N_11974,N_11899);
or U12067 (N_12067,N_11919,N_11927);
nor U12068 (N_12068,N_11910,N_11902);
nor U12069 (N_12069,N_11953,N_11917);
xnor U12070 (N_12070,N_11929,N_11902);
or U12071 (N_12071,N_11898,N_11914);
and U12072 (N_12072,N_11944,N_11931);
xnor U12073 (N_12073,N_11938,N_11941);
and U12074 (N_12074,N_11921,N_11908);
or U12075 (N_12075,N_11938,N_11989);
nand U12076 (N_12076,N_11958,N_11877);
nor U12077 (N_12077,N_11941,N_11960);
nor U12078 (N_12078,N_11875,N_11963);
xor U12079 (N_12079,N_11996,N_11915);
and U12080 (N_12080,N_11894,N_11937);
and U12081 (N_12081,N_11991,N_11890);
or U12082 (N_12082,N_11972,N_11951);
nand U12083 (N_12083,N_11909,N_11971);
nand U12084 (N_12084,N_11954,N_11988);
or U12085 (N_12085,N_11994,N_11886);
xnor U12086 (N_12086,N_11917,N_11966);
nand U12087 (N_12087,N_11912,N_11956);
nor U12088 (N_12088,N_11887,N_11994);
and U12089 (N_12089,N_11931,N_11994);
nand U12090 (N_12090,N_11908,N_11938);
nand U12091 (N_12091,N_11904,N_11978);
xor U12092 (N_12092,N_11964,N_11941);
xnor U12093 (N_12093,N_11985,N_11966);
nor U12094 (N_12094,N_11939,N_11979);
nor U12095 (N_12095,N_11923,N_11885);
or U12096 (N_12096,N_11943,N_11892);
xnor U12097 (N_12097,N_11898,N_11876);
or U12098 (N_12098,N_11884,N_11969);
and U12099 (N_12099,N_11997,N_11974);
nand U12100 (N_12100,N_11948,N_11953);
or U12101 (N_12101,N_11876,N_11953);
and U12102 (N_12102,N_11976,N_11889);
nor U12103 (N_12103,N_11931,N_11950);
and U12104 (N_12104,N_11894,N_11897);
or U12105 (N_12105,N_11963,N_11895);
xnor U12106 (N_12106,N_11926,N_11944);
xnor U12107 (N_12107,N_11878,N_11979);
nand U12108 (N_12108,N_11882,N_11968);
and U12109 (N_12109,N_11886,N_11929);
or U12110 (N_12110,N_11903,N_11991);
or U12111 (N_12111,N_11915,N_11944);
or U12112 (N_12112,N_11998,N_11987);
or U12113 (N_12113,N_11955,N_11947);
xor U12114 (N_12114,N_11933,N_11915);
or U12115 (N_12115,N_11995,N_11993);
xor U12116 (N_12116,N_11920,N_11967);
and U12117 (N_12117,N_11921,N_11951);
nand U12118 (N_12118,N_11896,N_11986);
xnor U12119 (N_12119,N_11900,N_11902);
nand U12120 (N_12120,N_11991,N_11953);
or U12121 (N_12121,N_11924,N_11980);
and U12122 (N_12122,N_11977,N_11916);
xor U12123 (N_12123,N_11957,N_11878);
xor U12124 (N_12124,N_11916,N_11904);
or U12125 (N_12125,N_12118,N_12110);
or U12126 (N_12126,N_12019,N_12072);
xnor U12127 (N_12127,N_12045,N_12076);
and U12128 (N_12128,N_12078,N_12006);
nand U12129 (N_12129,N_12040,N_12060);
nand U12130 (N_12130,N_12075,N_12105);
xor U12131 (N_12131,N_12086,N_12096);
xnor U12132 (N_12132,N_12095,N_12124);
or U12133 (N_12133,N_12066,N_12107);
and U12134 (N_12134,N_12013,N_12106);
nand U12135 (N_12135,N_12100,N_12021);
or U12136 (N_12136,N_12082,N_12032);
xnor U12137 (N_12137,N_12069,N_12053);
nand U12138 (N_12138,N_12074,N_12079);
nor U12139 (N_12139,N_12000,N_12098);
and U12140 (N_12140,N_12055,N_12004);
and U12141 (N_12141,N_12023,N_12009);
and U12142 (N_12142,N_12065,N_12102);
or U12143 (N_12143,N_12025,N_12062);
xnor U12144 (N_12144,N_12026,N_12061);
nor U12145 (N_12145,N_12070,N_12093);
nor U12146 (N_12146,N_12015,N_12018);
nand U12147 (N_12147,N_12014,N_12020);
xnor U12148 (N_12148,N_12092,N_12029);
or U12149 (N_12149,N_12104,N_12089);
xnor U12150 (N_12150,N_12041,N_12056);
nor U12151 (N_12151,N_12058,N_12064);
xor U12152 (N_12152,N_12037,N_12054);
and U12153 (N_12153,N_12017,N_12005);
nor U12154 (N_12154,N_12010,N_12071);
or U12155 (N_12155,N_12115,N_12049);
nor U12156 (N_12156,N_12113,N_12034);
and U12157 (N_12157,N_12044,N_12039);
and U12158 (N_12158,N_12068,N_12038);
xnor U12159 (N_12159,N_12036,N_12031);
xnor U12160 (N_12160,N_12114,N_12063);
nand U12161 (N_12161,N_12099,N_12073);
nand U12162 (N_12162,N_12024,N_12002);
xor U12163 (N_12163,N_12122,N_12111);
xnor U12164 (N_12164,N_12047,N_12091);
and U12165 (N_12165,N_12090,N_12052);
and U12166 (N_12166,N_12085,N_12094);
nor U12167 (N_12167,N_12077,N_12048);
xor U12168 (N_12168,N_12042,N_12116);
xnor U12169 (N_12169,N_12088,N_12081);
or U12170 (N_12170,N_12033,N_12112);
or U12171 (N_12171,N_12050,N_12008);
and U12172 (N_12172,N_12057,N_12028);
or U12173 (N_12173,N_12087,N_12012);
nor U12174 (N_12174,N_12035,N_12119);
xnor U12175 (N_12175,N_12101,N_12117);
and U12176 (N_12176,N_12011,N_12097);
nand U12177 (N_12177,N_12003,N_12007);
and U12178 (N_12178,N_12022,N_12120);
xnor U12179 (N_12179,N_12051,N_12001);
xor U12180 (N_12180,N_12109,N_12083);
nor U12181 (N_12181,N_12059,N_12084);
nand U12182 (N_12182,N_12121,N_12027);
nand U12183 (N_12183,N_12043,N_12123);
xor U12184 (N_12184,N_12030,N_12103);
nor U12185 (N_12185,N_12016,N_12108);
nand U12186 (N_12186,N_12067,N_12080);
and U12187 (N_12187,N_12046,N_12072);
xor U12188 (N_12188,N_12030,N_12003);
and U12189 (N_12189,N_12016,N_12101);
or U12190 (N_12190,N_12089,N_12122);
nand U12191 (N_12191,N_12094,N_12010);
nand U12192 (N_12192,N_12115,N_12096);
nand U12193 (N_12193,N_12025,N_12049);
or U12194 (N_12194,N_12060,N_12116);
and U12195 (N_12195,N_12041,N_12025);
or U12196 (N_12196,N_12025,N_12024);
and U12197 (N_12197,N_12097,N_12076);
nand U12198 (N_12198,N_12043,N_12107);
or U12199 (N_12199,N_12107,N_12064);
or U12200 (N_12200,N_12004,N_12044);
nand U12201 (N_12201,N_12113,N_12056);
or U12202 (N_12202,N_12004,N_12101);
or U12203 (N_12203,N_12079,N_12000);
xor U12204 (N_12204,N_12025,N_12089);
and U12205 (N_12205,N_12074,N_12052);
nand U12206 (N_12206,N_12083,N_12035);
nand U12207 (N_12207,N_12088,N_12105);
nand U12208 (N_12208,N_12084,N_12032);
or U12209 (N_12209,N_12027,N_12065);
nand U12210 (N_12210,N_12065,N_12044);
and U12211 (N_12211,N_12092,N_12008);
xor U12212 (N_12212,N_12056,N_12103);
nand U12213 (N_12213,N_12012,N_12050);
xnor U12214 (N_12214,N_12008,N_12100);
and U12215 (N_12215,N_12096,N_12028);
or U12216 (N_12216,N_12029,N_12120);
nand U12217 (N_12217,N_12118,N_12102);
nand U12218 (N_12218,N_12036,N_12065);
nor U12219 (N_12219,N_12043,N_12029);
nand U12220 (N_12220,N_12111,N_12027);
nand U12221 (N_12221,N_12004,N_12094);
or U12222 (N_12222,N_12071,N_12039);
nor U12223 (N_12223,N_12020,N_12077);
and U12224 (N_12224,N_12072,N_12038);
or U12225 (N_12225,N_12056,N_12082);
nor U12226 (N_12226,N_12108,N_12026);
xnor U12227 (N_12227,N_12058,N_12121);
nor U12228 (N_12228,N_12022,N_12029);
nand U12229 (N_12229,N_12051,N_12063);
xnor U12230 (N_12230,N_12097,N_12022);
nor U12231 (N_12231,N_12040,N_12071);
and U12232 (N_12232,N_12028,N_12011);
nor U12233 (N_12233,N_12048,N_12033);
and U12234 (N_12234,N_12089,N_12096);
nand U12235 (N_12235,N_12106,N_12022);
nor U12236 (N_12236,N_12011,N_12074);
nand U12237 (N_12237,N_12079,N_12019);
and U12238 (N_12238,N_12054,N_12048);
nand U12239 (N_12239,N_12018,N_12013);
nand U12240 (N_12240,N_12010,N_12009);
nand U12241 (N_12241,N_12041,N_12072);
nand U12242 (N_12242,N_12123,N_12074);
or U12243 (N_12243,N_12059,N_12009);
nor U12244 (N_12244,N_12020,N_12023);
nand U12245 (N_12245,N_12015,N_12027);
xnor U12246 (N_12246,N_12020,N_12045);
nand U12247 (N_12247,N_12037,N_12031);
xor U12248 (N_12248,N_12093,N_12107);
nand U12249 (N_12249,N_12004,N_12099);
nand U12250 (N_12250,N_12186,N_12145);
or U12251 (N_12251,N_12164,N_12235);
or U12252 (N_12252,N_12191,N_12185);
nor U12253 (N_12253,N_12147,N_12197);
or U12254 (N_12254,N_12130,N_12211);
xor U12255 (N_12255,N_12146,N_12196);
nor U12256 (N_12256,N_12214,N_12229);
and U12257 (N_12257,N_12226,N_12232);
or U12258 (N_12258,N_12135,N_12246);
xnor U12259 (N_12259,N_12248,N_12141);
nand U12260 (N_12260,N_12139,N_12176);
and U12261 (N_12261,N_12210,N_12206);
nand U12262 (N_12262,N_12160,N_12205);
or U12263 (N_12263,N_12129,N_12181);
and U12264 (N_12264,N_12138,N_12223);
xnor U12265 (N_12265,N_12167,N_12231);
xor U12266 (N_12266,N_12132,N_12208);
or U12267 (N_12267,N_12236,N_12249);
nand U12268 (N_12268,N_12207,N_12243);
or U12269 (N_12269,N_12137,N_12184);
nand U12270 (N_12270,N_12165,N_12194);
and U12271 (N_12271,N_12242,N_12199);
nor U12272 (N_12272,N_12162,N_12180);
xor U12273 (N_12273,N_12217,N_12134);
nor U12274 (N_12274,N_12193,N_12169);
xnor U12275 (N_12275,N_12155,N_12200);
and U12276 (N_12276,N_12238,N_12245);
nor U12277 (N_12277,N_12140,N_12189);
or U12278 (N_12278,N_12183,N_12168);
and U12279 (N_12279,N_12133,N_12212);
xnor U12280 (N_12280,N_12178,N_12225);
xor U12281 (N_12281,N_12126,N_12218);
nand U12282 (N_12282,N_12241,N_12131);
and U12283 (N_12283,N_12239,N_12209);
and U12284 (N_12284,N_12159,N_12203);
nor U12285 (N_12285,N_12222,N_12244);
xor U12286 (N_12286,N_12173,N_12128);
nand U12287 (N_12287,N_12221,N_12237);
and U12288 (N_12288,N_12188,N_12195);
nor U12289 (N_12289,N_12192,N_12153);
nor U12290 (N_12290,N_12148,N_12198);
xor U12291 (N_12291,N_12172,N_12202);
or U12292 (N_12292,N_12174,N_12143);
nor U12293 (N_12293,N_12127,N_12158);
nand U12294 (N_12294,N_12233,N_12136);
nand U12295 (N_12295,N_12201,N_12170);
nor U12296 (N_12296,N_12216,N_12163);
nand U12297 (N_12297,N_12166,N_12213);
nor U12298 (N_12298,N_12224,N_12179);
and U12299 (N_12299,N_12150,N_12157);
and U12300 (N_12300,N_12230,N_12152);
nor U12301 (N_12301,N_12125,N_12151);
xnor U12302 (N_12302,N_12154,N_12247);
nor U12303 (N_12303,N_12228,N_12240);
nor U12304 (N_12304,N_12187,N_12161);
xor U12305 (N_12305,N_12177,N_12142);
nor U12306 (N_12306,N_12219,N_12171);
nand U12307 (N_12307,N_12204,N_12182);
nand U12308 (N_12308,N_12215,N_12220);
and U12309 (N_12309,N_12227,N_12149);
xor U12310 (N_12310,N_12175,N_12190);
nand U12311 (N_12311,N_12144,N_12234);
nand U12312 (N_12312,N_12156,N_12188);
and U12313 (N_12313,N_12162,N_12248);
and U12314 (N_12314,N_12194,N_12192);
or U12315 (N_12315,N_12133,N_12175);
and U12316 (N_12316,N_12154,N_12158);
and U12317 (N_12317,N_12183,N_12198);
and U12318 (N_12318,N_12235,N_12145);
xor U12319 (N_12319,N_12145,N_12249);
nand U12320 (N_12320,N_12185,N_12196);
xor U12321 (N_12321,N_12139,N_12217);
and U12322 (N_12322,N_12188,N_12189);
or U12323 (N_12323,N_12220,N_12130);
nand U12324 (N_12324,N_12135,N_12143);
and U12325 (N_12325,N_12187,N_12178);
nor U12326 (N_12326,N_12178,N_12173);
and U12327 (N_12327,N_12212,N_12208);
nand U12328 (N_12328,N_12225,N_12230);
nor U12329 (N_12329,N_12188,N_12224);
nand U12330 (N_12330,N_12159,N_12145);
nor U12331 (N_12331,N_12171,N_12221);
and U12332 (N_12332,N_12190,N_12219);
nand U12333 (N_12333,N_12246,N_12176);
nor U12334 (N_12334,N_12218,N_12144);
xnor U12335 (N_12335,N_12212,N_12150);
nand U12336 (N_12336,N_12159,N_12243);
or U12337 (N_12337,N_12199,N_12184);
nor U12338 (N_12338,N_12241,N_12249);
xor U12339 (N_12339,N_12198,N_12249);
nand U12340 (N_12340,N_12134,N_12179);
nand U12341 (N_12341,N_12197,N_12245);
or U12342 (N_12342,N_12207,N_12141);
or U12343 (N_12343,N_12191,N_12242);
or U12344 (N_12344,N_12133,N_12197);
nand U12345 (N_12345,N_12213,N_12178);
and U12346 (N_12346,N_12221,N_12174);
nand U12347 (N_12347,N_12133,N_12230);
xor U12348 (N_12348,N_12177,N_12149);
or U12349 (N_12349,N_12127,N_12192);
and U12350 (N_12350,N_12247,N_12128);
xor U12351 (N_12351,N_12226,N_12244);
nor U12352 (N_12352,N_12170,N_12192);
or U12353 (N_12353,N_12248,N_12207);
nand U12354 (N_12354,N_12181,N_12174);
and U12355 (N_12355,N_12208,N_12228);
nor U12356 (N_12356,N_12168,N_12132);
and U12357 (N_12357,N_12128,N_12160);
xnor U12358 (N_12358,N_12190,N_12242);
xnor U12359 (N_12359,N_12197,N_12186);
xor U12360 (N_12360,N_12207,N_12153);
or U12361 (N_12361,N_12165,N_12230);
and U12362 (N_12362,N_12198,N_12244);
and U12363 (N_12363,N_12161,N_12205);
and U12364 (N_12364,N_12217,N_12130);
xor U12365 (N_12365,N_12155,N_12206);
and U12366 (N_12366,N_12234,N_12198);
or U12367 (N_12367,N_12140,N_12234);
or U12368 (N_12368,N_12231,N_12171);
and U12369 (N_12369,N_12202,N_12171);
nand U12370 (N_12370,N_12217,N_12135);
or U12371 (N_12371,N_12214,N_12183);
xor U12372 (N_12372,N_12244,N_12151);
and U12373 (N_12373,N_12141,N_12129);
xor U12374 (N_12374,N_12156,N_12220);
nor U12375 (N_12375,N_12301,N_12332);
and U12376 (N_12376,N_12279,N_12310);
nand U12377 (N_12377,N_12293,N_12267);
nand U12378 (N_12378,N_12352,N_12339);
xnor U12379 (N_12379,N_12254,N_12300);
nor U12380 (N_12380,N_12365,N_12262);
and U12381 (N_12381,N_12329,N_12304);
xor U12382 (N_12382,N_12324,N_12303);
xnor U12383 (N_12383,N_12348,N_12311);
nor U12384 (N_12384,N_12359,N_12306);
and U12385 (N_12385,N_12255,N_12354);
and U12386 (N_12386,N_12307,N_12314);
and U12387 (N_12387,N_12288,N_12369);
nor U12388 (N_12388,N_12295,N_12276);
and U12389 (N_12389,N_12264,N_12260);
and U12390 (N_12390,N_12292,N_12312);
nand U12391 (N_12391,N_12258,N_12290);
nand U12392 (N_12392,N_12252,N_12286);
xnor U12393 (N_12393,N_12297,N_12257);
or U12394 (N_12394,N_12305,N_12294);
nor U12395 (N_12395,N_12298,N_12280);
xnor U12396 (N_12396,N_12334,N_12350);
or U12397 (N_12397,N_12275,N_12336);
nand U12398 (N_12398,N_12368,N_12321);
nor U12399 (N_12399,N_12362,N_12357);
xor U12400 (N_12400,N_12281,N_12341);
and U12401 (N_12401,N_12272,N_12331);
nor U12402 (N_12402,N_12338,N_12256);
nor U12403 (N_12403,N_12284,N_12340);
or U12404 (N_12404,N_12363,N_12253);
and U12405 (N_12405,N_12372,N_12318);
xor U12406 (N_12406,N_12335,N_12351);
xnor U12407 (N_12407,N_12342,N_12358);
or U12408 (N_12408,N_12323,N_12355);
or U12409 (N_12409,N_12271,N_12366);
or U12410 (N_12410,N_12309,N_12337);
nand U12411 (N_12411,N_12317,N_12364);
or U12412 (N_12412,N_12373,N_12270);
and U12413 (N_12413,N_12299,N_12282);
or U12414 (N_12414,N_12269,N_12333);
nand U12415 (N_12415,N_12349,N_12259);
or U12416 (N_12416,N_12325,N_12313);
and U12417 (N_12417,N_12273,N_12308);
xnor U12418 (N_12418,N_12371,N_12367);
or U12419 (N_12419,N_12326,N_12347);
nand U12420 (N_12420,N_12328,N_12361);
nor U12421 (N_12421,N_12296,N_12291);
or U12422 (N_12422,N_12343,N_12250);
nor U12423 (N_12423,N_12370,N_12268);
nand U12424 (N_12424,N_12353,N_12346);
nor U12425 (N_12425,N_12330,N_12263);
or U12426 (N_12426,N_12261,N_12278);
nand U12427 (N_12427,N_12265,N_12289);
or U12428 (N_12428,N_12285,N_12251);
xnor U12429 (N_12429,N_12316,N_12322);
and U12430 (N_12430,N_12277,N_12327);
and U12431 (N_12431,N_12287,N_12274);
or U12432 (N_12432,N_12320,N_12302);
nand U12433 (N_12433,N_12345,N_12356);
or U12434 (N_12434,N_12266,N_12344);
and U12435 (N_12435,N_12319,N_12374);
nand U12436 (N_12436,N_12315,N_12360);
or U12437 (N_12437,N_12283,N_12269);
and U12438 (N_12438,N_12275,N_12357);
nor U12439 (N_12439,N_12290,N_12372);
and U12440 (N_12440,N_12374,N_12339);
or U12441 (N_12441,N_12309,N_12255);
nand U12442 (N_12442,N_12285,N_12316);
nor U12443 (N_12443,N_12263,N_12270);
xor U12444 (N_12444,N_12270,N_12316);
and U12445 (N_12445,N_12320,N_12339);
or U12446 (N_12446,N_12348,N_12354);
or U12447 (N_12447,N_12262,N_12357);
nor U12448 (N_12448,N_12341,N_12352);
and U12449 (N_12449,N_12354,N_12323);
or U12450 (N_12450,N_12293,N_12282);
and U12451 (N_12451,N_12340,N_12293);
xor U12452 (N_12452,N_12273,N_12364);
nand U12453 (N_12453,N_12318,N_12312);
nor U12454 (N_12454,N_12370,N_12346);
nand U12455 (N_12455,N_12280,N_12323);
or U12456 (N_12456,N_12311,N_12371);
nor U12457 (N_12457,N_12339,N_12350);
or U12458 (N_12458,N_12338,N_12366);
or U12459 (N_12459,N_12313,N_12283);
xnor U12460 (N_12460,N_12274,N_12330);
and U12461 (N_12461,N_12363,N_12336);
and U12462 (N_12462,N_12330,N_12283);
and U12463 (N_12463,N_12281,N_12320);
nor U12464 (N_12464,N_12370,N_12292);
xor U12465 (N_12465,N_12252,N_12337);
or U12466 (N_12466,N_12329,N_12367);
xnor U12467 (N_12467,N_12260,N_12348);
xnor U12468 (N_12468,N_12340,N_12302);
and U12469 (N_12469,N_12339,N_12319);
and U12470 (N_12470,N_12351,N_12337);
xor U12471 (N_12471,N_12352,N_12270);
nand U12472 (N_12472,N_12315,N_12304);
nand U12473 (N_12473,N_12358,N_12315);
xnor U12474 (N_12474,N_12273,N_12353);
xnor U12475 (N_12475,N_12261,N_12305);
nand U12476 (N_12476,N_12319,N_12354);
xnor U12477 (N_12477,N_12289,N_12364);
nor U12478 (N_12478,N_12326,N_12253);
xor U12479 (N_12479,N_12258,N_12367);
and U12480 (N_12480,N_12271,N_12348);
and U12481 (N_12481,N_12366,N_12273);
nor U12482 (N_12482,N_12263,N_12342);
nor U12483 (N_12483,N_12309,N_12347);
nor U12484 (N_12484,N_12258,N_12273);
or U12485 (N_12485,N_12289,N_12257);
xnor U12486 (N_12486,N_12372,N_12264);
nor U12487 (N_12487,N_12318,N_12257);
nand U12488 (N_12488,N_12317,N_12348);
nor U12489 (N_12489,N_12337,N_12370);
and U12490 (N_12490,N_12352,N_12366);
and U12491 (N_12491,N_12264,N_12257);
xnor U12492 (N_12492,N_12348,N_12319);
or U12493 (N_12493,N_12293,N_12254);
xnor U12494 (N_12494,N_12346,N_12279);
or U12495 (N_12495,N_12320,N_12285);
nand U12496 (N_12496,N_12368,N_12300);
xor U12497 (N_12497,N_12276,N_12255);
xnor U12498 (N_12498,N_12257,N_12258);
nand U12499 (N_12499,N_12261,N_12272);
and U12500 (N_12500,N_12389,N_12432);
xor U12501 (N_12501,N_12461,N_12387);
and U12502 (N_12502,N_12433,N_12472);
or U12503 (N_12503,N_12490,N_12487);
nor U12504 (N_12504,N_12396,N_12406);
and U12505 (N_12505,N_12405,N_12457);
nor U12506 (N_12506,N_12446,N_12424);
xnor U12507 (N_12507,N_12449,N_12417);
nor U12508 (N_12508,N_12496,N_12482);
or U12509 (N_12509,N_12467,N_12408);
xor U12510 (N_12510,N_12392,N_12412);
nor U12511 (N_12511,N_12464,N_12498);
or U12512 (N_12512,N_12455,N_12398);
and U12513 (N_12513,N_12441,N_12439);
and U12514 (N_12514,N_12428,N_12375);
nor U12515 (N_12515,N_12429,N_12471);
and U12516 (N_12516,N_12415,N_12409);
or U12517 (N_12517,N_12474,N_12488);
and U12518 (N_12518,N_12481,N_12463);
nand U12519 (N_12519,N_12478,N_12475);
nor U12520 (N_12520,N_12466,N_12425);
nor U12521 (N_12521,N_12489,N_12494);
and U12522 (N_12522,N_12447,N_12442);
and U12523 (N_12523,N_12423,N_12401);
or U12524 (N_12524,N_12460,N_12410);
xnor U12525 (N_12525,N_12480,N_12391);
nand U12526 (N_12526,N_12380,N_12384);
xnor U12527 (N_12527,N_12402,N_12453);
and U12528 (N_12528,N_12434,N_12451);
and U12529 (N_12529,N_12414,N_12397);
xor U12530 (N_12530,N_12435,N_12470);
or U12531 (N_12531,N_12438,N_12493);
xnor U12532 (N_12532,N_12473,N_12459);
nand U12533 (N_12533,N_12476,N_12400);
and U12534 (N_12534,N_12426,N_12382);
or U12535 (N_12535,N_12492,N_12421);
nor U12536 (N_12536,N_12445,N_12416);
xnor U12537 (N_12537,N_12378,N_12484);
and U12538 (N_12538,N_12443,N_12468);
nand U12539 (N_12539,N_12379,N_12394);
nor U12540 (N_12540,N_12427,N_12404);
and U12541 (N_12541,N_12413,N_12462);
nor U12542 (N_12542,N_12407,N_12390);
and U12543 (N_12543,N_12381,N_12483);
and U12544 (N_12544,N_12377,N_12479);
xor U12545 (N_12545,N_12436,N_12419);
xor U12546 (N_12546,N_12450,N_12403);
nor U12547 (N_12547,N_12491,N_12422);
or U12548 (N_12548,N_12437,N_12440);
nor U12549 (N_12549,N_12495,N_12458);
xor U12550 (N_12550,N_12485,N_12395);
xor U12551 (N_12551,N_12465,N_12420);
xor U12552 (N_12552,N_12376,N_12411);
nor U12553 (N_12553,N_12383,N_12452);
nor U12554 (N_12554,N_12393,N_12385);
and U12555 (N_12555,N_12499,N_12477);
xor U12556 (N_12556,N_12456,N_12486);
nor U12557 (N_12557,N_12454,N_12386);
xnor U12558 (N_12558,N_12469,N_12448);
xor U12559 (N_12559,N_12388,N_12431);
nand U12560 (N_12560,N_12430,N_12444);
and U12561 (N_12561,N_12497,N_12399);
and U12562 (N_12562,N_12418,N_12490);
nand U12563 (N_12563,N_12419,N_12429);
nor U12564 (N_12564,N_12391,N_12390);
xor U12565 (N_12565,N_12406,N_12445);
or U12566 (N_12566,N_12483,N_12403);
or U12567 (N_12567,N_12434,N_12445);
or U12568 (N_12568,N_12407,N_12483);
xnor U12569 (N_12569,N_12381,N_12464);
and U12570 (N_12570,N_12491,N_12493);
nor U12571 (N_12571,N_12386,N_12458);
nand U12572 (N_12572,N_12402,N_12484);
nor U12573 (N_12573,N_12432,N_12482);
nor U12574 (N_12574,N_12445,N_12447);
and U12575 (N_12575,N_12383,N_12467);
or U12576 (N_12576,N_12386,N_12375);
nor U12577 (N_12577,N_12413,N_12456);
nor U12578 (N_12578,N_12404,N_12394);
nand U12579 (N_12579,N_12440,N_12455);
nand U12580 (N_12580,N_12448,N_12437);
and U12581 (N_12581,N_12440,N_12377);
xnor U12582 (N_12582,N_12432,N_12475);
nand U12583 (N_12583,N_12390,N_12441);
nand U12584 (N_12584,N_12449,N_12379);
nand U12585 (N_12585,N_12415,N_12392);
or U12586 (N_12586,N_12499,N_12396);
nand U12587 (N_12587,N_12431,N_12423);
nor U12588 (N_12588,N_12445,N_12421);
or U12589 (N_12589,N_12441,N_12397);
nand U12590 (N_12590,N_12376,N_12409);
or U12591 (N_12591,N_12408,N_12395);
nand U12592 (N_12592,N_12436,N_12390);
nand U12593 (N_12593,N_12497,N_12474);
nand U12594 (N_12594,N_12445,N_12432);
xor U12595 (N_12595,N_12398,N_12478);
xor U12596 (N_12596,N_12423,N_12454);
nand U12597 (N_12597,N_12479,N_12496);
and U12598 (N_12598,N_12379,N_12462);
or U12599 (N_12599,N_12461,N_12497);
and U12600 (N_12600,N_12420,N_12476);
nor U12601 (N_12601,N_12420,N_12425);
xnor U12602 (N_12602,N_12474,N_12470);
nand U12603 (N_12603,N_12435,N_12452);
nand U12604 (N_12604,N_12493,N_12382);
nand U12605 (N_12605,N_12408,N_12421);
or U12606 (N_12606,N_12476,N_12384);
and U12607 (N_12607,N_12380,N_12376);
nand U12608 (N_12608,N_12411,N_12396);
or U12609 (N_12609,N_12434,N_12381);
and U12610 (N_12610,N_12446,N_12441);
nor U12611 (N_12611,N_12469,N_12408);
or U12612 (N_12612,N_12432,N_12466);
and U12613 (N_12613,N_12452,N_12463);
and U12614 (N_12614,N_12413,N_12429);
and U12615 (N_12615,N_12434,N_12497);
and U12616 (N_12616,N_12445,N_12462);
xnor U12617 (N_12617,N_12389,N_12427);
xnor U12618 (N_12618,N_12376,N_12421);
nor U12619 (N_12619,N_12479,N_12434);
nor U12620 (N_12620,N_12425,N_12481);
nand U12621 (N_12621,N_12383,N_12470);
and U12622 (N_12622,N_12415,N_12478);
or U12623 (N_12623,N_12491,N_12381);
xnor U12624 (N_12624,N_12420,N_12403);
nand U12625 (N_12625,N_12605,N_12608);
and U12626 (N_12626,N_12571,N_12532);
and U12627 (N_12627,N_12594,N_12592);
or U12628 (N_12628,N_12504,N_12609);
nand U12629 (N_12629,N_12517,N_12610);
nor U12630 (N_12630,N_12513,N_12531);
and U12631 (N_12631,N_12558,N_12549);
xnor U12632 (N_12632,N_12550,N_12535);
xor U12633 (N_12633,N_12599,N_12556);
nand U12634 (N_12634,N_12507,N_12617);
xnor U12635 (N_12635,N_12520,N_12501);
xnor U12636 (N_12636,N_12590,N_12611);
xor U12637 (N_12637,N_12509,N_12525);
xor U12638 (N_12638,N_12578,N_12546);
or U12639 (N_12639,N_12575,N_12506);
and U12640 (N_12640,N_12576,N_12552);
nor U12641 (N_12641,N_12559,N_12580);
xnor U12642 (N_12642,N_12540,N_12574);
and U12643 (N_12643,N_12566,N_12616);
nand U12644 (N_12644,N_12544,N_12555);
nor U12645 (N_12645,N_12533,N_12606);
or U12646 (N_12646,N_12557,N_12584);
or U12647 (N_12647,N_12621,N_12563);
and U12648 (N_12648,N_12624,N_12591);
nand U12649 (N_12649,N_12593,N_12514);
nor U12650 (N_12650,N_12620,N_12613);
nor U12651 (N_12651,N_12551,N_12553);
or U12652 (N_12652,N_12602,N_12595);
nor U12653 (N_12653,N_12545,N_12615);
and U12654 (N_12654,N_12526,N_12561);
nand U12655 (N_12655,N_12565,N_12618);
xnor U12656 (N_12656,N_12541,N_12585);
nor U12657 (N_12657,N_12607,N_12573);
or U12658 (N_12658,N_12523,N_12587);
xor U12659 (N_12659,N_12581,N_12515);
xor U12660 (N_12660,N_12572,N_12589);
nor U12661 (N_12661,N_12582,N_12601);
or U12662 (N_12662,N_12564,N_12530);
nand U12663 (N_12663,N_12534,N_12598);
or U12664 (N_12664,N_12612,N_12569);
xnor U12665 (N_12665,N_12500,N_12511);
nand U12666 (N_12666,N_12579,N_12529);
nor U12667 (N_12667,N_12512,N_12568);
nor U12668 (N_12668,N_12597,N_12596);
nor U12669 (N_12669,N_12503,N_12508);
nor U12670 (N_12670,N_12600,N_12586);
xor U12671 (N_12671,N_12537,N_12567);
and U12672 (N_12672,N_12619,N_12539);
and U12673 (N_12673,N_12604,N_12547);
and U12674 (N_12674,N_12622,N_12570);
and U12675 (N_12675,N_12623,N_12548);
xor U12676 (N_12676,N_12614,N_12502);
and U12677 (N_12677,N_12518,N_12543);
or U12678 (N_12678,N_12528,N_12577);
nor U12679 (N_12679,N_12510,N_12538);
xor U12680 (N_12680,N_12516,N_12527);
and U12681 (N_12681,N_12603,N_12505);
nor U12682 (N_12682,N_12522,N_12560);
and U12683 (N_12683,N_12562,N_12521);
xor U12684 (N_12684,N_12583,N_12519);
nor U12685 (N_12685,N_12588,N_12554);
xnor U12686 (N_12686,N_12536,N_12524);
xor U12687 (N_12687,N_12542,N_12583);
or U12688 (N_12688,N_12539,N_12523);
and U12689 (N_12689,N_12613,N_12565);
nor U12690 (N_12690,N_12522,N_12624);
and U12691 (N_12691,N_12577,N_12520);
xnor U12692 (N_12692,N_12583,N_12599);
xnor U12693 (N_12693,N_12595,N_12566);
xnor U12694 (N_12694,N_12590,N_12584);
xor U12695 (N_12695,N_12537,N_12513);
nand U12696 (N_12696,N_12623,N_12624);
and U12697 (N_12697,N_12592,N_12591);
nor U12698 (N_12698,N_12579,N_12568);
xor U12699 (N_12699,N_12502,N_12518);
xnor U12700 (N_12700,N_12519,N_12553);
xor U12701 (N_12701,N_12562,N_12583);
nor U12702 (N_12702,N_12616,N_12598);
xor U12703 (N_12703,N_12599,N_12572);
or U12704 (N_12704,N_12526,N_12504);
or U12705 (N_12705,N_12594,N_12550);
or U12706 (N_12706,N_12573,N_12523);
nor U12707 (N_12707,N_12563,N_12512);
nor U12708 (N_12708,N_12617,N_12599);
nor U12709 (N_12709,N_12508,N_12614);
or U12710 (N_12710,N_12588,N_12612);
or U12711 (N_12711,N_12603,N_12594);
and U12712 (N_12712,N_12578,N_12597);
nand U12713 (N_12713,N_12617,N_12564);
or U12714 (N_12714,N_12600,N_12531);
or U12715 (N_12715,N_12611,N_12580);
xor U12716 (N_12716,N_12582,N_12605);
nand U12717 (N_12717,N_12544,N_12546);
nor U12718 (N_12718,N_12500,N_12605);
nand U12719 (N_12719,N_12596,N_12524);
and U12720 (N_12720,N_12532,N_12608);
nor U12721 (N_12721,N_12531,N_12532);
or U12722 (N_12722,N_12509,N_12560);
and U12723 (N_12723,N_12600,N_12545);
nand U12724 (N_12724,N_12525,N_12516);
nor U12725 (N_12725,N_12530,N_12560);
and U12726 (N_12726,N_12546,N_12553);
nor U12727 (N_12727,N_12513,N_12538);
or U12728 (N_12728,N_12593,N_12541);
or U12729 (N_12729,N_12591,N_12539);
xor U12730 (N_12730,N_12598,N_12589);
and U12731 (N_12731,N_12610,N_12576);
nand U12732 (N_12732,N_12558,N_12568);
or U12733 (N_12733,N_12531,N_12569);
nor U12734 (N_12734,N_12623,N_12608);
nand U12735 (N_12735,N_12570,N_12509);
nor U12736 (N_12736,N_12536,N_12551);
xnor U12737 (N_12737,N_12505,N_12527);
xnor U12738 (N_12738,N_12540,N_12573);
nor U12739 (N_12739,N_12597,N_12544);
xor U12740 (N_12740,N_12524,N_12609);
nor U12741 (N_12741,N_12563,N_12525);
or U12742 (N_12742,N_12614,N_12603);
nor U12743 (N_12743,N_12563,N_12618);
xor U12744 (N_12744,N_12615,N_12590);
or U12745 (N_12745,N_12596,N_12605);
nor U12746 (N_12746,N_12501,N_12582);
xor U12747 (N_12747,N_12521,N_12590);
xnor U12748 (N_12748,N_12532,N_12612);
or U12749 (N_12749,N_12593,N_12587);
nand U12750 (N_12750,N_12723,N_12735);
xor U12751 (N_12751,N_12661,N_12724);
nand U12752 (N_12752,N_12733,N_12708);
or U12753 (N_12753,N_12682,N_12725);
nor U12754 (N_12754,N_12703,N_12651);
nor U12755 (N_12755,N_12629,N_12743);
xnor U12756 (N_12756,N_12746,N_12670);
nand U12757 (N_12757,N_12689,N_12704);
nor U12758 (N_12758,N_12730,N_12666);
and U12759 (N_12759,N_12678,N_12654);
and U12760 (N_12760,N_12676,N_12736);
and U12761 (N_12761,N_12732,N_12718);
nor U12762 (N_12762,N_12700,N_12660);
nand U12763 (N_12763,N_12693,N_12745);
or U12764 (N_12764,N_12740,N_12681);
and U12765 (N_12765,N_12635,N_12728);
and U12766 (N_12766,N_12719,N_12630);
xor U12767 (N_12767,N_12639,N_12652);
or U12768 (N_12768,N_12748,N_12679);
xnor U12769 (N_12769,N_12687,N_12749);
xor U12770 (N_12770,N_12707,N_12712);
or U12771 (N_12771,N_12628,N_12706);
and U12772 (N_12772,N_12716,N_12636);
xor U12773 (N_12773,N_12662,N_12633);
and U12774 (N_12774,N_12717,N_12640);
or U12775 (N_12775,N_12720,N_12638);
nand U12776 (N_12776,N_12664,N_12697);
xor U12777 (N_12777,N_12727,N_12741);
nand U12778 (N_12778,N_12675,N_12691);
nor U12779 (N_12779,N_12684,N_12726);
nor U12780 (N_12780,N_12713,N_12737);
or U12781 (N_12781,N_12715,N_12722);
and U12782 (N_12782,N_12702,N_12686);
nor U12783 (N_12783,N_12710,N_12705);
nand U12784 (N_12784,N_12690,N_12742);
nor U12785 (N_12785,N_12729,N_12644);
nand U12786 (N_12786,N_12626,N_12731);
or U12787 (N_12787,N_12663,N_12685);
and U12788 (N_12788,N_12721,N_12739);
nor U12789 (N_12789,N_12650,N_12655);
and U12790 (N_12790,N_12641,N_12637);
nor U12791 (N_12791,N_12659,N_12714);
nor U12792 (N_12792,N_12744,N_12631);
nor U12793 (N_12793,N_12649,N_12657);
or U12794 (N_12794,N_12692,N_12688);
or U12795 (N_12795,N_12647,N_12673);
or U12796 (N_12796,N_12671,N_12658);
and U12797 (N_12797,N_12642,N_12656);
and U12798 (N_12798,N_12627,N_12668);
and U12799 (N_12799,N_12672,N_12698);
nand U12800 (N_12800,N_12680,N_12634);
and U12801 (N_12801,N_12674,N_12645);
xnor U12802 (N_12802,N_12667,N_12709);
or U12803 (N_12803,N_12747,N_12677);
nand U12804 (N_12804,N_12699,N_12734);
and U12805 (N_12805,N_12665,N_12696);
xnor U12806 (N_12806,N_12643,N_12695);
nor U12807 (N_12807,N_12669,N_12653);
or U12808 (N_12808,N_12632,N_12711);
nor U12809 (N_12809,N_12701,N_12648);
xnor U12810 (N_12810,N_12694,N_12683);
or U12811 (N_12811,N_12646,N_12625);
nor U12812 (N_12812,N_12738,N_12648);
nor U12813 (N_12813,N_12648,N_12672);
or U12814 (N_12814,N_12628,N_12640);
nor U12815 (N_12815,N_12730,N_12682);
or U12816 (N_12816,N_12693,N_12678);
or U12817 (N_12817,N_12720,N_12656);
and U12818 (N_12818,N_12695,N_12671);
nor U12819 (N_12819,N_12657,N_12741);
or U12820 (N_12820,N_12667,N_12642);
nand U12821 (N_12821,N_12749,N_12695);
nor U12822 (N_12822,N_12714,N_12727);
xnor U12823 (N_12823,N_12687,N_12705);
nor U12824 (N_12824,N_12662,N_12729);
nor U12825 (N_12825,N_12682,N_12640);
nand U12826 (N_12826,N_12674,N_12636);
nor U12827 (N_12827,N_12697,N_12727);
xnor U12828 (N_12828,N_12727,N_12662);
nor U12829 (N_12829,N_12734,N_12693);
or U12830 (N_12830,N_12691,N_12708);
xnor U12831 (N_12831,N_12710,N_12656);
nand U12832 (N_12832,N_12689,N_12748);
xor U12833 (N_12833,N_12668,N_12710);
nand U12834 (N_12834,N_12656,N_12682);
and U12835 (N_12835,N_12734,N_12670);
nor U12836 (N_12836,N_12695,N_12669);
and U12837 (N_12837,N_12647,N_12658);
xor U12838 (N_12838,N_12704,N_12709);
or U12839 (N_12839,N_12706,N_12642);
and U12840 (N_12840,N_12693,N_12701);
or U12841 (N_12841,N_12746,N_12647);
nor U12842 (N_12842,N_12657,N_12692);
nor U12843 (N_12843,N_12650,N_12714);
nand U12844 (N_12844,N_12655,N_12631);
nand U12845 (N_12845,N_12653,N_12656);
nand U12846 (N_12846,N_12641,N_12653);
nand U12847 (N_12847,N_12716,N_12669);
xor U12848 (N_12848,N_12693,N_12655);
and U12849 (N_12849,N_12630,N_12659);
and U12850 (N_12850,N_12626,N_12676);
nand U12851 (N_12851,N_12713,N_12724);
xnor U12852 (N_12852,N_12650,N_12687);
nand U12853 (N_12853,N_12660,N_12687);
xor U12854 (N_12854,N_12741,N_12662);
xnor U12855 (N_12855,N_12721,N_12664);
nor U12856 (N_12856,N_12701,N_12736);
nand U12857 (N_12857,N_12696,N_12739);
xnor U12858 (N_12858,N_12636,N_12698);
nand U12859 (N_12859,N_12661,N_12725);
nor U12860 (N_12860,N_12709,N_12743);
or U12861 (N_12861,N_12689,N_12658);
xor U12862 (N_12862,N_12744,N_12743);
and U12863 (N_12863,N_12712,N_12715);
and U12864 (N_12864,N_12632,N_12643);
and U12865 (N_12865,N_12637,N_12728);
nor U12866 (N_12866,N_12677,N_12660);
nand U12867 (N_12867,N_12672,N_12649);
or U12868 (N_12868,N_12705,N_12667);
nand U12869 (N_12869,N_12693,N_12676);
nor U12870 (N_12870,N_12692,N_12690);
nand U12871 (N_12871,N_12637,N_12629);
nor U12872 (N_12872,N_12628,N_12667);
and U12873 (N_12873,N_12693,N_12660);
or U12874 (N_12874,N_12721,N_12643);
xnor U12875 (N_12875,N_12832,N_12791);
or U12876 (N_12876,N_12846,N_12854);
or U12877 (N_12877,N_12760,N_12822);
nor U12878 (N_12878,N_12858,N_12873);
nor U12879 (N_12879,N_12838,N_12774);
nand U12880 (N_12880,N_12757,N_12755);
xnor U12881 (N_12881,N_12835,N_12866);
nand U12882 (N_12882,N_12786,N_12834);
xor U12883 (N_12883,N_12762,N_12753);
or U12884 (N_12884,N_12847,N_12754);
xnor U12885 (N_12885,N_12848,N_12856);
and U12886 (N_12886,N_12767,N_12845);
nand U12887 (N_12887,N_12789,N_12833);
nand U12888 (N_12888,N_12826,N_12808);
nor U12889 (N_12889,N_12758,N_12855);
xnor U12890 (N_12890,N_12868,N_12788);
nand U12891 (N_12891,N_12836,N_12853);
xnor U12892 (N_12892,N_12844,N_12790);
or U12893 (N_12893,N_12830,N_12859);
nand U12894 (N_12894,N_12817,N_12870);
nor U12895 (N_12895,N_12860,N_12752);
nor U12896 (N_12896,N_12764,N_12829);
nor U12897 (N_12897,N_12796,N_12781);
xnor U12898 (N_12898,N_12850,N_12863);
or U12899 (N_12899,N_12807,N_12841);
nand U12900 (N_12900,N_12825,N_12823);
and U12901 (N_12901,N_12864,N_12811);
nand U12902 (N_12902,N_12843,N_12827);
nand U12903 (N_12903,N_12805,N_12766);
xnor U12904 (N_12904,N_12750,N_12759);
xnor U12905 (N_12905,N_12865,N_12824);
nor U12906 (N_12906,N_12828,N_12837);
nor U12907 (N_12907,N_12782,N_12794);
xor U12908 (N_12908,N_12756,N_12775);
or U12909 (N_12909,N_12798,N_12819);
nor U12910 (N_12910,N_12783,N_12812);
nor U12911 (N_12911,N_12771,N_12768);
nand U12912 (N_12912,N_12872,N_12773);
nand U12913 (N_12913,N_12869,N_12867);
nor U12914 (N_12914,N_12797,N_12862);
xor U12915 (N_12915,N_12799,N_12849);
and U12916 (N_12916,N_12802,N_12772);
nand U12917 (N_12917,N_12821,N_12861);
nor U12918 (N_12918,N_12816,N_12803);
and U12919 (N_12919,N_12777,N_12785);
xor U12920 (N_12920,N_12787,N_12831);
nand U12921 (N_12921,N_12793,N_12776);
nand U12922 (N_12922,N_12871,N_12769);
xnor U12923 (N_12923,N_12779,N_12801);
nor U12924 (N_12924,N_12815,N_12806);
xor U12925 (N_12925,N_12780,N_12842);
nand U12926 (N_12926,N_12839,N_12804);
nor U12927 (N_12927,N_12852,N_12763);
and U12928 (N_12928,N_12840,N_12751);
and U12929 (N_12929,N_12814,N_12851);
nor U12930 (N_12930,N_12820,N_12770);
nor U12931 (N_12931,N_12800,N_12813);
and U12932 (N_12932,N_12765,N_12857);
or U12933 (N_12933,N_12874,N_12792);
nor U12934 (N_12934,N_12795,N_12809);
or U12935 (N_12935,N_12778,N_12761);
nor U12936 (N_12936,N_12810,N_12818);
or U12937 (N_12937,N_12784,N_12804);
or U12938 (N_12938,N_12762,N_12801);
or U12939 (N_12939,N_12865,N_12768);
and U12940 (N_12940,N_12829,N_12857);
xnor U12941 (N_12941,N_12754,N_12765);
nand U12942 (N_12942,N_12796,N_12767);
nor U12943 (N_12943,N_12806,N_12837);
xor U12944 (N_12944,N_12820,N_12774);
xnor U12945 (N_12945,N_12834,N_12833);
xor U12946 (N_12946,N_12869,N_12874);
xor U12947 (N_12947,N_12787,N_12801);
xnor U12948 (N_12948,N_12765,N_12828);
nand U12949 (N_12949,N_12808,N_12844);
or U12950 (N_12950,N_12797,N_12792);
nand U12951 (N_12951,N_12753,N_12863);
and U12952 (N_12952,N_12817,N_12871);
or U12953 (N_12953,N_12776,N_12814);
xnor U12954 (N_12954,N_12842,N_12764);
or U12955 (N_12955,N_12847,N_12869);
xnor U12956 (N_12956,N_12836,N_12764);
nand U12957 (N_12957,N_12795,N_12874);
nand U12958 (N_12958,N_12806,N_12811);
nand U12959 (N_12959,N_12857,N_12816);
and U12960 (N_12960,N_12807,N_12760);
nand U12961 (N_12961,N_12759,N_12773);
nand U12962 (N_12962,N_12776,N_12797);
and U12963 (N_12963,N_12873,N_12826);
xnor U12964 (N_12964,N_12764,N_12808);
or U12965 (N_12965,N_12794,N_12868);
and U12966 (N_12966,N_12853,N_12865);
or U12967 (N_12967,N_12766,N_12798);
nor U12968 (N_12968,N_12758,N_12817);
nor U12969 (N_12969,N_12794,N_12789);
nor U12970 (N_12970,N_12818,N_12796);
or U12971 (N_12971,N_12818,N_12820);
nand U12972 (N_12972,N_12856,N_12766);
nand U12973 (N_12973,N_12871,N_12818);
nand U12974 (N_12974,N_12759,N_12783);
or U12975 (N_12975,N_12829,N_12839);
nand U12976 (N_12976,N_12845,N_12840);
nand U12977 (N_12977,N_12807,N_12872);
nand U12978 (N_12978,N_12829,N_12791);
xnor U12979 (N_12979,N_12780,N_12855);
xor U12980 (N_12980,N_12815,N_12797);
and U12981 (N_12981,N_12867,N_12801);
nand U12982 (N_12982,N_12862,N_12772);
and U12983 (N_12983,N_12865,N_12806);
or U12984 (N_12984,N_12782,N_12773);
or U12985 (N_12985,N_12828,N_12779);
nor U12986 (N_12986,N_12854,N_12776);
nand U12987 (N_12987,N_12835,N_12830);
and U12988 (N_12988,N_12752,N_12756);
xor U12989 (N_12989,N_12827,N_12766);
xor U12990 (N_12990,N_12870,N_12796);
nand U12991 (N_12991,N_12860,N_12798);
nand U12992 (N_12992,N_12831,N_12873);
xor U12993 (N_12993,N_12763,N_12787);
or U12994 (N_12994,N_12806,N_12761);
and U12995 (N_12995,N_12849,N_12813);
nor U12996 (N_12996,N_12821,N_12828);
and U12997 (N_12997,N_12775,N_12815);
and U12998 (N_12998,N_12810,N_12870);
nor U12999 (N_12999,N_12807,N_12781);
nand U13000 (N_13000,N_12935,N_12932);
nand U13001 (N_13001,N_12978,N_12894);
xnor U13002 (N_13002,N_12891,N_12889);
and U13003 (N_13003,N_12923,N_12887);
nand U13004 (N_13004,N_12877,N_12985);
or U13005 (N_13005,N_12921,N_12886);
or U13006 (N_13006,N_12961,N_12981);
nand U13007 (N_13007,N_12915,N_12954);
xor U13008 (N_13008,N_12948,N_12922);
nand U13009 (N_13009,N_12912,N_12958);
nor U13010 (N_13010,N_12969,N_12914);
xor U13011 (N_13011,N_12946,N_12930);
xnor U13012 (N_13012,N_12918,N_12890);
xor U13013 (N_13013,N_12907,N_12945);
or U13014 (N_13014,N_12972,N_12933);
xor U13015 (N_13015,N_12967,N_12908);
and U13016 (N_13016,N_12942,N_12899);
xnor U13017 (N_13017,N_12976,N_12993);
nand U13018 (N_13018,N_12951,N_12916);
or U13019 (N_13019,N_12936,N_12911);
and U13020 (N_13020,N_12938,N_12926);
or U13021 (N_13021,N_12953,N_12917);
nor U13022 (N_13022,N_12971,N_12984);
or U13023 (N_13023,N_12919,N_12939);
nor U13024 (N_13024,N_12964,N_12878);
nand U13025 (N_13025,N_12924,N_12988);
or U13026 (N_13026,N_12898,N_12997);
nor U13027 (N_13027,N_12944,N_12965);
or U13028 (N_13028,N_12928,N_12943);
xnor U13029 (N_13029,N_12909,N_12910);
xor U13030 (N_13030,N_12986,N_12995);
xor U13031 (N_13031,N_12884,N_12987);
and U13032 (N_13032,N_12994,N_12885);
or U13033 (N_13033,N_12966,N_12880);
nand U13034 (N_13034,N_12881,N_12974);
xor U13035 (N_13035,N_12888,N_12925);
nor U13036 (N_13036,N_12934,N_12906);
or U13037 (N_13037,N_12876,N_12940);
nor U13038 (N_13038,N_12893,N_12920);
or U13039 (N_13039,N_12962,N_12960);
and U13040 (N_13040,N_12902,N_12975);
or U13041 (N_13041,N_12979,N_12977);
xor U13042 (N_13042,N_12913,N_12882);
nand U13043 (N_13043,N_12999,N_12955);
xor U13044 (N_13044,N_12903,N_12875);
nor U13045 (N_13045,N_12901,N_12973);
nor U13046 (N_13046,N_12929,N_12947);
xnor U13047 (N_13047,N_12879,N_12895);
nor U13048 (N_13048,N_12996,N_12998);
nand U13049 (N_13049,N_12950,N_12892);
nand U13050 (N_13050,N_12989,N_12970);
or U13051 (N_13051,N_12980,N_12927);
and U13052 (N_13052,N_12931,N_12896);
nand U13053 (N_13053,N_12904,N_12897);
nand U13054 (N_13054,N_12941,N_12959);
nor U13055 (N_13055,N_12883,N_12957);
nand U13056 (N_13056,N_12983,N_12963);
xor U13057 (N_13057,N_12952,N_12968);
or U13058 (N_13058,N_12982,N_12900);
or U13059 (N_13059,N_12937,N_12905);
nand U13060 (N_13060,N_12992,N_12991);
and U13061 (N_13061,N_12949,N_12956);
nand U13062 (N_13062,N_12990,N_12957);
xnor U13063 (N_13063,N_12971,N_12956);
and U13064 (N_13064,N_12979,N_12944);
xor U13065 (N_13065,N_12929,N_12935);
nand U13066 (N_13066,N_12888,N_12909);
or U13067 (N_13067,N_12969,N_12907);
and U13068 (N_13068,N_12970,N_12987);
nor U13069 (N_13069,N_12931,N_12986);
nand U13070 (N_13070,N_12991,N_12925);
or U13071 (N_13071,N_12888,N_12979);
and U13072 (N_13072,N_12979,N_12984);
nor U13073 (N_13073,N_12909,N_12962);
and U13074 (N_13074,N_12985,N_12945);
nand U13075 (N_13075,N_12908,N_12963);
and U13076 (N_13076,N_12952,N_12924);
and U13077 (N_13077,N_12893,N_12974);
or U13078 (N_13078,N_12930,N_12952);
nor U13079 (N_13079,N_12932,N_12982);
and U13080 (N_13080,N_12963,N_12961);
nand U13081 (N_13081,N_12931,N_12886);
xnor U13082 (N_13082,N_12984,N_12908);
nand U13083 (N_13083,N_12900,N_12907);
and U13084 (N_13084,N_12907,N_12997);
and U13085 (N_13085,N_12986,N_12948);
nand U13086 (N_13086,N_12923,N_12973);
nor U13087 (N_13087,N_12951,N_12887);
nand U13088 (N_13088,N_12938,N_12928);
nor U13089 (N_13089,N_12956,N_12959);
xor U13090 (N_13090,N_12908,N_12968);
or U13091 (N_13091,N_12914,N_12890);
or U13092 (N_13092,N_12928,N_12886);
nand U13093 (N_13093,N_12942,N_12977);
nand U13094 (N_13094,N_12989,N_12919);
or U13095 (N_13095,N_12965,N_12877);
and U13096 (N_13096,N_12898,N_12987);
xor U13097 (N_13097,N_12875,N_12982);
nand U13098 (N_13098,N_12969,N_12983);
xor U13099 (N_13099,N_12916,N_12997);
nand U13100 (N_13100,N_12998,N_12976);
and U13101 (N_13101,N_12907,N_12948);
or U13102 (N_13102,N_12997,N_12938);
xor U13103 (N_13103,N_12881,N_12982);
or U13104 (N_13104,N_12921,N_12994);
xnor U13105 (N_13105,N_12903,N_12948);
or U13106 (N_13106,N_12926,N_12939);
nand U13107 (N_13107,N_12905,N_12982);
and U13108 (N_13108,N_12981,N_12933);
nor U13109 (N_13109,N_12998,N_12883);
nor U13110 (N_13110,N_12912,N_12968);
xor U13111 (N_13111,N_12986,N_12894);
or U13112 (N_13112,N_12913,N_12982);
and U13113 (N_13113,N_12978,N_12961);
or U13114 (N_13114,N_12926,N_12935);
nor U13115 (N_13115,N_12912,N_12908);
nand U13116 (N_13116,N_12949,N_12924);
nor U13117 (N_13117,N_12942,N_12937);
xor U13118 (N_13118,N_12978,N_12896);
and U13119 (N_13119,N_12993,N_12914);
nand U13120 (N_13120,N_12986,N_12952);
or U13121 (N_13121,N_12989,N_12914);
nand U13122 (N_13122,N_12974,N_12946);
or U13123 (N_13123,N_12977,N_12904);
and U13124 (N_13124,N_12906,N_12982);
nand U13125 (N_13125,N_13099,N_13003);
nand U13126 (N_13126,N_13107,N_13088);
xor U13127 (N_13127,N_13106,N_13046);
nor U13128 (N_13128,N_13056,N_13032);
nor U13129 (N_13129,N_13113,N_13121);
and U13130 (N_13130,N_13023,N_13093);
and U13131 (N_13131,N_13105,N_13020);
nor U13132 (N_13132,N_13074,N_13005);
nor U13133 (N_13133,N_13052,N_13114);
nor U13134 (N_13134,N_13024,N_13049);
nand U13135 (N_13135,N_13048,N_13089);
xor U13136 (N_13136,N_13076,N_13071);
nor U13137 (N_13137,N_13043,N_13039);
and U13138 (N_13138,N_13102,N_13031);
nand U13139 (N_13139,N_13066,N_13119);
nand U13140 (N_13140,N_13051,N_13103);
nand U13141 (N_13141,N_13041,N_13094);
nor U13142 (N_13142,N_13063,N_13018);
or U13143 (N_13143,N_13029,N_13069);
nand U13144 (N_13144,N_13015,N_13042);
nor U13145 (N_13145,N_13091,N_13004);
or U13146 (N_13146,N_13006,N_13096);
or U13147 (N_13147,N_13082,N_13011);
nor U13148 (N_13148,N_13059,N_13012);
xor U13149 (N_13149,N_13057,N_13028);
and U13150 (N_13150,N_13061,N_13021);
nor U13151 (N_13151,N_13067,N_13007);
and U13152 (N_13152,N_13002,N_13072);
nor U13153 (N_13153,N_13079,N_13097);
xor U13154 (N_13154,N_13084,N_13075);
nand U13155 (N_13155,N_13080,N_13077);
xnor U13156 (N_13156,N_13060,N_13090);
nand U13157 (N_13157,N_13095,N_13036);
nor U13158 (N_13158,N_13124,N_13053);
nor U13159 (N_13159,N_13000,N_13073);
or U13160 (N_13160,N_13026,N_13111);
nand U13161 (N_13161,N_13008,N_13001);
or U13162 (N_13162,N_13118,N_13017);
or U13163 (N_13163,N_13085,N_13025);
xnor U13164 (N_13164,N_13013,N_13050);
xor U13165 (N_13165,N_13064,N_13100);
or U13166 (N_13166,N_13092,N_13045);
or U13167 (N_13167,N_13033,N_13083);
nor U13168 (N_13168,N_13108,N_13009);
nor U13169 (N_13169,N_13037,N_13117);
or U13170 (N_13170,N_13040,N_13035);
xnor U13171 (N_13171,N_13078,N_13054);
nor U13172 (N_13172,N_13122,N_13038);
or U13173 (N_13173,N_13019,N_13055);
nor U13174 (N_13174,N_13027,N_13110);
xnor U13175 (N_13175,N_13115,N_13070);
nand U13176 (N_13176,N_13065,N_13109);
xnor U13177 (N_13177,N_13104,N_13044);
or U13178 (N_13178,N_13087,N_13034);
nor U13179 (N_13179,N_13030,N_13098);
nor U13180 (N_13180,N_13101,N_13112);
xor U13181 (N_13181,N_13010,N_13116);
xor U13182 (N_13182,N_13062,N_13120);
nor U13183 (N_13183,N_13068,N_13058);
or U13184 (N_13184,N_13123,N_13014);
and U13185 (N_13185,N_13022,N_13081);
xor U13186 (N_13186,N_13016,N_13047);
nor U13187 (N_13187,N_13086,N_13016);
nand U13188 (N_13188,N_13052,N_13105);
or U13189 (N_13189,N_13029,N_13008);
and U13190 (N_13190,N_13084,N_13077);
nand U13191 (N_13191,N_13032,N_13093);
and U13192 (N_13192,N_13009,N_13033);
and U13193 (N_13193,N_13103,N_13006);
nand U13194 (N_13194,N_13123,N_13065);
and U13195 (N_13195,N_13046,N_13079);
nor U13196 (N_13196,N_13025,N_13116);
xor U13197 (N_13197,N_13072,N_13052);
and U13198 (N_13198,N_13106,N_13050);
nand U13199 (N_13199,N_13065,N_13052);
xor U13200 (N_13200,N_13027,N_13099);
or U13201 (N_13201,N_13047,N_13025);
xnor U13202 (N_13202,N_13124,N_13114);
and U13203 (N_13203,N_13053,N_13012);
and U13204 (N_13204,N_13040,N_13034);
or U13205 (N_13205,N_13091,N_13025);
nand U13206 (N_13206,N_13014,N_13015);
nand U13207 (N_13207,N_13043,N_13003);
nor U13208 (N_13208,N_13028,N_13120);
xor U13209 (N_13209,N_13018,N_13113);
nor U13210 (N_13210,N_13010,N_13102);
nor U13211 (N_13211,N_13048,N_13056);
and U13212 (N_13212,N_13034,N_13039);
nand U13213 (N_13213,N_13006,N_13116);
nand U13214 (N_13214,N_13099,N_13039);
and U13215 (N_13215,N_13108,N_13018);
nand U13216 (N_13216,N_13108,N_13011);
nor U13217 (N_13217,N_13058,N_13006);
nor U13218 (N_13218,N_13089,N_13116);
xor U13219 (N_13219,N_13113,N_13118);
nor U13220 (N_13220,N_13053,N_13087);
nand U13221 (N_13221,N_13073,N_13037);
nand U13222 (N_13222,N_13003,N_13017);
xor U13223 (N_13223,N_13004,N_13090);
and U13224 (N_13224,N_13000,N_13066);
xor U13225 (N_13225,N_13002,N_13105);
or U13226 (N_13226,N_13079,N_13068);
nor U13227 (N_13227,N_13023,N_13020);
xor U13228 (N_13228,N_13052,N_13111);
and U13229 (N_13229,N_13020,N_13002);
and U13230 (N_13230,N_13034,N_13089);
xor U13231 (N_13231,N_13064,N_13008);
xor U13232 (N_13232,N_13071,N_13107);
or U13233 (N_13233,N_13122,N_13091);
nor U13234 (N_13234,N_13070,N_13096);
xor U13235 (N_13235,N_13098,N_13066);
and U13236 (N_13236,N_13080,N_13059);
or U13237 (N_13237,N_13115,N_13053);
or U13238 (N_13238,N_13100,N_13051);
xor U13239 (N_13239,N_13021,N_13028);
nand U13240 (N_13240,N_13051,N_13121);
nand U13241 (N_13241,N_13015,N_13114);
nand U13242 (N_13242,N_13113,N_13081);
and U13243 (N_13243,N_13094,N_13011);
nor U13244 (N_13244,N_13110,N_13007);
nand U13245 (N_13245,N_13078,N_13030);
or U13246 (N_13246,N_13115,N_13110);
or U13247 (N_13247,N_13103,N_13040);
and U13248 (N_13248,N_13070,N_13109);
xnor U13249 (N_13249,N_13083,N_13071);
or U13250 (N_13250,N_13129,N_13239);
and U13251 (N_13251,N_13224,N_13248);
or U13252 (N_13252,N_13146,N_13221);
and U13253 (N_13253,N_13215,N_13246);
nand U13254 (N_13254,N_13192,N_13143);
nor U13255 (N_13255,N_13194,N_13195);
nand U13256 (N_13256,N_13241,N_13132);
xnor U13257 (N_13257,N_13147,N_13141);
nand U13258 (N_13258,N_13164,N_13227);
nor U13259 (N_13259,N_13242,N_13174);
nand U13260 (N_13260,N_13139,N_13200);
and U13261 (N_13261,N_13183,N_13196);
and U13262 (N_13262,N_13236,N_13175);
or U13263 (N_13263,N_13230,N_13220);
nor U13264 (N_13264,N_13185,N_13206);
nand U13265 (N_13265,N_13222,N_13157);
and U13266 (N_13266,N_13162,N_13219);
xnor U13267 (N_13267,N_13186,N_13148);
xnor U13268 (N_13268,N_13182,N_13159);
nor U13269 (N_13269,N_13201,N_13173);
nand U13270 (N_13270,N_13178,N_13212);
nand U13271 (N_13271,N_13187,N_13211);
and U13272 (N_13272,N_13213,N_13126);
xor U13273 (N_13273,N_13223,N_13163);
and U13274 (N_13274,N_13172,N_13135);
and U13275 (N_13275,N_13134,N_13180);
or U13276 (N_13276,N_13152,N_13137);
or U13277 (N_13277,N_13234,N_13168);
or U13278 (N_13278,N_13210,N_13214);
nor U13279 (N_13279,N_13161,N_13233);
nor U13280 (N_13280,N_13188,N_13176);
or U13281 (N_13281,N_13156,N_13136);
xnor U13282 (N_13282,N_13240,N_13127);
or U13283 (N_13283,N_13225,N_13167);
xor U13284 (N_13284,N_13149,N_13198);
xor U13285 (N_13285,N_13142,N_13209);
nand U13286 (N_13286,N_13217,N_13190);
xnor U13287 (N_13287,N_13243,N_13131);
and U13288 (N_13288,N_13249,N_13169);
nor U13289 (N_13289,N_13229,N_13155);
and U13290 (N_13290,N_13171,N_13238);
nand U13291 (N_13291,N_13128,N_13140);
xnor U13292 (N_13292,N_13170,N_13144);
and U13293 (N_13293,N_13247,N_13166);
or U13294 (N_13294,N_13216,N_13202);
xor U13295 (N_13295,N_13181,N_13125);
nand U13296 (N_13296,N_13177,N_13199);
nor U13297 (N_13297,N_13237,N_13160);
xnor U13298 (N_13298,N_13205,N_13154);
or U13299 (N_13299,N_13153,N_13138);
xnor U13300 (N_13300,N_13130,N_13218);
or U13301 (N_13301,N_13208,N_13179);
and U13302 (N_13302,N_13232,N_13207);
and U13303 (N_13303,N_13228,N_13158);
nand U13304 (N_13304,N_13245,N_13204);
nand U13305 (N_13305,N_13226,N_13203);
and U13306 (N_13306,N_13197,N_13150);
nand U13307 (N_13307,N_13193,N_13151);
or U13308 (N_13308,N_13191,N_13133);
nor U13309 (N_13309,N_13244,N_13145);
or U13310 (N_13310,N_13184,N_13231);
xor U13311 (N_13311,N_13235,N_13189);
xnor U13312 (N_13312,N_13165,N_13232);
or U13313 (N_13313,N_13225,N_13235);
or U13314 (N_13314,N_13232,N_13240);
and U13315 (N_13315,N_13195,N_13170);
or U13316 (N_13316,N_13231,N_13239);
xnor U13317 (N_13317,N_13233,N_13157);
nor U13318 (N_13318,N_13186,N_13190);
and U13319 (N_13319,N_13209,N_13227);
xor U13320 (N_13320,N_13151,N_13205);
or U13321 (N_13321,N_13225,N_13203);
nand U13322 (N_13322,N_13237,N_13244);
and U13323 (N_13323,N_13154,N_13150);
or U13324 (N_13324,N_13142,N_13198);
or U13325 (N_13325,N_13149,N_13193);
and U13326 (N_13326,N_13183,N_13176);
xor U13327 (N_13327,N_13165,N_13151);
and U13328 (N_13328,N_13192,N_13186);
or U13329 (N_13329,N_13187,N_13185);
nor U13330 (N_13330,N_13226,N_13200);
and U13331 (N_13331,N_13222,N_13217);
xor U13332 (N_13332,N_13215,N_13221);
xnor U13333 (N_13333,N_13226,N_13179);
and U13334 (N_13334,N_13177,N_13175);
nor U13335 (N_13335,N_13215,N_13241);
nor U13336 (N_13336,N_13162,N_13223);
xor U13337 (N_13337,N_13163,N_13171);
and U13338 (N_13338,N_13181,N_13224);
and U13339 (N_13339,N_13160,N_13171);
nand U13340 (N_13340,N_13129,N_13126);
nand U13341 (N_13341,N_13190,N_13224);
and U13342 (N_13342,N_13234,N_13183);
and U13343 (N_13343,N_13131,N_13228);
nand U13344 (N_13344,N_13183,N_13190);
nand U13345 (N_13345,N_13197,N_13137);
and U13346 (N_13346,N_13208,N_13231);
or U13347 (N_13347,N_13161,N_13153);
nor U13348 (N_13348,N_13130,N_13244);
nor U13349 (N_13349,N_13246,N_13165);
xnor U13350 (N_13350,N_13162,N_13144);
xor U13351 (N_13351,N_13150,N_13163);
or U13352 (N_13352,N_13194,N_13203);
nand U13353 (N_13353,N_13236,N_13206);
or U13354 (N_13354,N_13182,N_13157);
and U13355 (N_13355,N_13127,N_13192);
or U13356 (N_13356,N_13242,N_13159);
xor U13357 (N_13357,N_13166,N_13184);
or U13358 (N_13358,N_13206,N_13180);
nand U13359 (N_13359,N_13228,N_13215);
xnor U13360 (N_13360,N_13232,N_13226);
xnor U13361 (N_13361,N_13164,N_13206);
nand U13362 (N_13362,N_13171,N_13152);
and U13363 (N_13363,N_13238,N_13155);
and U13364 (N_13364,N_13130,N_13239);
nor U13365 (N_13365,N_13153,N_13235);
nand U13366 (N_13366,N_13153,N_13149);
and U13367 (N_13367,N_13194,N_13177);
and U13368 (N_13368,N_13196,N_13194);
and U13369 (N_13369,N_13132,N_13235);
nand U13370 (N_13370,N_13220,N_13176);
nor U13371 (N_13371,N_13133,N_13130);
or U13372 (N_13372,N_13155,N_13164);
and U13373 (N_13373,N_13221,N_13202);
and U13374 (N_13374,N_13240,N_13212);
nand U13375 (N_13375,N_13269,N_13362);
and U13376 (N_13376,N_13356,N_13343);
nand U13377 (N_13377,N_13331,N_13255);
xnor U13378 (N_13378,N_13347,N_13370);
nand U13379 (N_13379,N_13346,N_13271);
or U13380 (N_13380,N_13282,N_13254);
and U13381 (N_13381,N_13264,N_13294);
nor U13382 (N_13382,N_13299,N_13320);
nor U13383 (N_13383,N_13277,N_13258);
nor U13384 (N_13384,N_13300,N_13361);
and U13385 (N_13385,N_13263,N_13252);
and U13386 (N_13386,N_13368,N_13292);
nand U13387 (N_13387,N_13297,N_13287);
or U13388 (N_13388,N_13309,N_13359);
and U13389 (N_13389,N_13253,N_13304);
or U13390 (N_13390,N_13279,N_13327);
xnor U13391 (N_13391,N_13291,N_13322);
nor U13392 (N_13392,N_13372,N_13310);
xor U13393 (N_13393,N_13260,N_13314);
xor U13394 (N_13394,N_13349,N_13358);
nor U13395 (N_13395,N_13357,N_13261);
nor U13396 (N_13396,N_13371,N_13326);
or U13397 (N_13397,N_13289,N_13280);
or U13398 (N_13398,N_13259,N_13367);
xor U13399 (N_13399,N_13328,N_13315);
and U13400 (N_13400,N_13284,N_13313);
xor U13401 (N_13401,N_13273,N_13266);
and U13402 (N_13402,N_13302,N_13306);
xnor U13403 (N_13403,N_13268,N_13251);
xor U13404 (N_13404,N_13272,N_13323);
nor U13405 (N_13405,N_13335,N_13286);
and U13406 (N_13406,N_13338,N_13329);
nor U13407 (N_13407,N_13369,N_13307);
or U13408 (N_13408,N_13250,N_13342);
nand U13409 (N_13409,N_13353,N_13324);
or U13410 (N_13410,N_13325,N_13374);
and U13411 (N_13411,N_13312,N_13311);
nand U13412 (N_13412,N_13290,N_13305);
and U13413 (N_13413,N_13373,N_13283);
or U13414 (N_13414,N_13256,N_13276);
nor U13415 (N_13415,N_13334,N_13363);
nor U13416 (N_13416,N_13317,N_13319);
and U13417 (N_13417,N_13257,N_13270);
xor U13418 (N_13418,N_13339,N_13332);
or U13419 (N_13419,N_13274,N_13285);
and U13420 (N_13420,N_13296,N_13355);
or U13421 (N_13421,N_13344,N_13267);
or U13422 (N_13422,N_13308,N_13281);
nand U13423 (N_13423,N_13336,N_13301);
or U13424 (N_13424,N_13364,N_13265);
nand U13425 (N_13425,N_13298,N_13341);
and U13426 (N_13426,N_13366,N_13340);
or U13427 (N_13427,N_13333,N_13365);
or U13428 (N_13428,N_13321,N_13288);
nor U13429 (N_13429,N_13262,N_13278);
or U13430 (N_13430,N_13295,N_13318);
or U13431 (N_13431,N_13352,N_13337);
and U13432 (N_13432,N_13354,N_13360);
nand U13433 (N_13433,N_13350,N_13316);
xor U13434 (N_13434,N_13293,N_13348);
nand U13435 (N_13435,N_13330,N_13351);
or U13436 (N_13436,N_13345,N_13275);
xor U13437 (N_13437,N_13303,N_13257);
and U13438 (N_13438,N_13367,N_13360);
nand U13439 (N_13439,N_13315,N_13364);
nor U13440 (N_13440,N_13256,N_13352);
and U13441 (N_13441,N_13267,N_13327);
nand U13442 (N_13442,N_13362,N_13275);
xnor U13443 (N_13443,N_13374,N_13251);
xor U13444 (N_13444,N_13260,N_13347);
or U13445 (N_13445,N_13371,N_13281);
nand U13446 (N_13446,N_13365,N_13339);
or U13447 (N_13447,N_13253,N_13309);
and U13448 (N_13448,N_13288,N_13251);
nand U13449 (N_13449,N_13349,N_13332);
xor U13450 (N_13450,N_13272,N_13338);
and U13451 (N_13451,N_13261,N_13369);
and U13452 (N_13452,N_13335,N_13274);
and U13453 (N_13453,N_13271,N_13344);
and U13454 (N_13454,N_13361,N_13355);
or U13455 (N_13455,N_13255,N_13315);
xnor U13456 (N_13456,N_13358,N_13324);
and U13457 (N_13457,N_13281,N_13324);
or U13458 (N_13458,N_13362,N_13266);
nor U13459 (N_13459,N_13280,N_13302);
nor U13460 (N_13460,N_13334,N_13311);
nand U13461 (N_13461,N_13368,N_13366);
or U13462 (N_13462,N_13257,N_13299);
nor U13463 (N_13463,N_13304,N_13366);
xor U13464 (N_13464,N_13335,N_13333);
xor U13465 (N_13465,N_13333,N_13321);
xnor U13466 (N_13466,N_13314,N_13350);
or U13467 (N_13467,N_13327,N_13284);
and U13468 (N_13468,N_13281,N_13286);
xnor U13469 (N_13469,N_13250,N_13255);
or U13470 (N_13470,N_13363,N_13271);
or U13471 (N_13471,N_13329,N_13363);
nor U13472 (N_13472,N_13369,N_13321);
nand U13473 (N_13473,N_13364,N_13289);
or U13474 (N_13474,N_13288,N_13285);
nand U13475 (N_13475,N_13353,N_13342);
or U13476 (N_13476,N_13296,N_13261);
nand U13477 (N_13477,N_13279,N_13364);
or U13478 (N_13478,N_13263,N_13329);
or U13479 (N_13479,N_13362,N_13363);
nor U13480 (N_13480,N_13310,N_13323);
nand U13481 (N_13481,N_13303,N_13363);
xnor U13482 (N_13482,N_13317,N_13310);
or U13483 (N_13483,N_13334,N_13318);
or U13484 (N_13484,N_13293,N_13313);
or U13485 (N_13485,N_13359,N_13368);
nor U13486 (N_13486,N_13255,N_13345);
nand U13487 (N_13487,N_13260,N_13254);
and U13488 (N_13488,N_13255,N_13291);
nor U13489 (N_13489,N_13322,N_13293);
nand U13490 (N_13490,N_13254,N_13296);
nor U13491 (N_13491,N_13283,N_13372);
nor U13492 (N_13492,N_13317,N_13262);
nor U13493 (N_13493,N_13338,N_13275);
nor U13494 (N_13494,N_13278,N_13319);
nand U13495 (N_13495,N_13275,N_13259);
or U13496 (N_13496,N_13277,N_13281);
and U13497 (N_13497,N_13294,N_13282);
nand U13498 (N_13498,N_13360,N_13357);
xnor U13499 (N_13499,N_13329,N_13281);
xnor U13500 (N_13500,N_13489,N_13391);
nor U13501 (N_13501,N_13410,N_13379);
and U13502 (N_13502,N_13496,N_13459);
and U13503 (N_13503,N_13386,N_13390);
xnor U13504 (N_13504,N_13424,N_13464);
xnor U13505 (N_13505,N_13411,N_13385);
xor U13506 (N_13506,N_13414,N_13431);
or U13507 (N_13507,N_13405,N_13393);
or U13508 (N_13508,N_13481,N_13449);
nand U13509 (N_13509,N_13387,N_13401);
nor U13510 (N_13510,N_13480,N_13428);
nor U13511 (N_13511,N_13397,N_13445);
nor U13512 (N_13512,N_13409,N_13479);
nor U13513 (N_13513,N_13378,N_13487);
nor U13514 (N_13514,N_13392,N_13376);
and U13515 (N_13515,N_13488,N_13412);
nand U13516 (N_13516,N_13476,N_13415);
nor U13517 (N_13517,N_13485,N_13426);
nand U13518 (N_13518,N_13438,N_13429);
and U13519 (N_13519,N_13472,N_13450);
or U13520 (N_13520,N_13474,N_13477);
and U13521 (N_13521,N_13465,N_13478);
nand U13522 (N_13522,N_13475,N_13382);
nand U13523 (N_13523,N_13470,N_13420);
nand U13524 (N_13524,N_13381,N_13448);
nor U13525 (N_13525,N_13463,N_13404);
nand U13526 (N_13526,N_13469,N_13398);
nand U13527 (N_13527,N_13399,N_13402);
nor U13528 (N_13528,N_13403,N_13407);
and U13529 (N_13529,N_13486,N_13444);
xnor U13530 (N_13530,N_13451,N_13384);
and U13531 (N_13531,N_13394,N_13377);
or U13532 (N_13532,N_13439,N_13455);
xnor U13533 (N_13533,N_13396,N_13471);
nand U13534 (N_13534,N_13497,N_13380);
nand U13535 (N_13535,N_13413,N_13383);
nand U13536 (N_13536,N_13454,N_13388);
nor U13537 (N_13537,N_13389,N_13435);
nor U13538 (N_13538,N_13462,N_13427);
or U13539 (N_13539,N_13400,N_13416);
or U13540 (N_13540,N_13491,N_13473);
xor U13541 (N_13541,N_13437,N_13408);
and U13542 (N_13542,N_13484,N_13433);
or U13543 (N_13543,N_13458,N_13425);
nand U13544 (N_13544,N_13467,N_13432);
or U13545 (N_13545,N_13453,N_13493);
or U13546 (N_13546,N_13456,N_13441);
xnor U13547 (N_13547,N_13466,N_13461);
nor U13548 (N_13548,N_13421,N_13442);
or U13549 (N_13549,N_13419,N_13468);
nand U13550 (N_13550,N_13452,N_13482);
nand U13551 (N_13551,N_13499,N_13498);
and U13552 (N_13552,N_13422,N_13492);
and U13553 (N_13553,N_13436,N_13495);
xnor U13554 (N_13554,N_13395,N_13423);
nor U13555 (N_13555,N_13434,N_13457);
xnor U13556 (N_13556,N_13417,N_13446);
and U13557 (N_13557,N_13460,N_13406);
and U13558 (N_13558,N_13443,N_13418);
and U13559 (N_13559,N_13483,N_13440);
xnor U13560 (N_13560,N_13447,N_13430);
nand U13561 (N_13561,N_13494,N_13375);
or U13562 (N_13562,N_13490,N_13469);
nand U13563 (N_13563,N_13442,N_13445);
xor U13564 (N_13564,N_13377,N_13472);
and U13565 (N_13565,N_13461,N_13431);
nor U13566 (N_13566,N_13405,N_13398);
nor U13567 (N_13567,N_13399,N_13432);
nand U13568 (N_13568,N_13435,N_13430);
or U13569 (N_13569,N_13445,N_13423);
nand U13570 (N_13570,N_13422,N_13427);
or U13571 (N_13571,N_13448,N_13440);
xnor U13572 (N_13572,N_13461,N_13468);
and U13573 (N_13573,N_13436,N_13483);
or U13574 (N_13574,N_13384,N_13481);
xnor U13575 (N_13575,N_13389,N_13491);
nor U13576 (N_13576,N_13378,N_13493);
nor U13577 (N_13577,N_13406,N_13451);
xor U13578 (N_13578,N_13456,N_13401);
nand U13579 (N_13579,N_13444,N_13423);
and U13580 (N_13580,N_13381,N_13475);
xor U13581 (N_13581,N_13488,N_13477);
nor U13582 (N_13582,N_13396,N_13467);
and U13583 (N_13583,N_13394,N_13479);
xor U13584 (N_13584,N_13449,N_13487);
and U13585 (N_13585,N_13414,N_13417);
and U13586 (N_13586,N_13436,N_13379);
nand U13587 (N_13587,N_13382,N_13463);
nor U13588 (N_13588,N_13447,N_13419);
xor U13589 (N_13589,N_13490,N_13405);
xor U13590 (N_13590,N_13424,N_13488);
xor U13591 (N_13591,N_13425,N_13473);
nand U13592 (N_13592,N_13418,N_13477);
and U13593 (N_13593,N_13385,N_13480);
or U13594 (N_13594,N_13398,N_13442);
and U13595 (N_13595,N_13477,N_13427);
and U13596 (N_13596,N_13412,N_13393);
nand U13597 (N_13597,N_13420,N_13476);
and U13598 (N_13598,N_13481,N_13490);
or U13599 (N_13599,N_13494,N_13386);
xor U13600 (N_13600,N_13436,N_13393);
nand U13601 (N_13601,N_13497,N_13438);
nor U13602 (N_13602,N_13413,N_13493);
or U13603 (N_13603,N_13472,N_13438);
nor U13604 (N_13604,N_13451,N_13381);
nand U13605 (N_13605,N_13428,N_13409);
xnor U13606 (N_13606,N_13469,N_13467);
xnor U13607 (N_13607,N_13428,N_13493);
nand U13608 (N_13608,N_13434,N_13441);
or U13609 (N_13609,N_13435,N_13394);
nor U13610 (N_13610,N_13492,N_13409);
or U13611 (N_13611,N_13455,N_13420);
xor U13612 (N_13612,N_13467,N_13417);
nand U13613 (N_13613,N_13471,N_13440);
nor U13614 (N_13614,N_13476,N_13438);
nor U13615 (N_13615,N_13461,N_13420);
nand U13616 (N_13616,N_13496,N_13465);
xor U13617 (N_13617,N_13398,N_13409);
nand U13618 (N_13618,N_13427,N_13491);
nand U13619 (N_13619,N_13380,N_13456);
nand U13620 (N_13620,N_13467,N_13498);
nand U13621 (N_13621,N_13377,N_13433);
nand U13622 (N_13622,N_13487,N_13455);
or U13623 (N_13623,N_13392,N_13464);
and U13624 (N_13624,N_13484,N_13436);
nand U13625 (N_13625,N_13564,N_13540);
nor U13626 (N_13626,N_13521,N_13551);
nand U13627 (N_13627,N_13529,N_13615);
nand U13628 (N_13628,N_13552,N_13570);
xor U13629 (N_13629,N_13608,N_13567);
and U13630 (N_13630,N_13612,N_13623);
or U13631 (N_13631,N_13512,N_13587);
and U13632 (N_13632,N_13539,N_13621);
and U13633 (N_13633,N_13532,N_13501);
nor U13634 (N_13634,N_13610,N_13533);
and U13635 (N_13635,N_13580,N_13578);
nor U13636 (N_13636,N_13550,N_13522);
xnor U13637 (N_13637,N_13618,N_13536);
nand U13638 (N_13638,N_13613,N_13557);
nor U13639 (N_13639,N_13617,N_13606);
xor U13640 (N_13640,N_13599,N_13517);
nor U13641 (N_13641,N_13559,N_13537);
and U13642 (N_13642,N_13500,N_13585);
nand U13643 (N_13643,N_13514,N_13598);
or U13644 (N_13644,N_13568,N_13505);
nor U13645 (N_13645,N_13614,N_13561);
nor U13646 (N_13646,N_13591,N_13502);
and U13647 (N_13647,N_13601,N_13574);
nand U13648 (N_13648,N_13544,N_13510);
or U13649 (N_13649,N_13604,N_13503);
nand U13650 (N_13650,N_13520,N_13575);
and U13651 (N_13651,N_13518,N_13507);
nand U13652 (N_13652,N_13595,N_13609);
and U13653 (N_13653,N_13605,N_13603);
nand U13654 (N_13654,N_13593,N_13583);
nor U13655 (N_13655,N_13597,N_13586);
nor U13656 (N_13656,N_13513,N_13619);
nor U13657 (N_13657,N_13543,N_13506);
or U13658 (N_13658,N_13547,N_13535);
and U13659 (N_13659,N_13624,N_13516);
and U13660 (N_13660,N_13620,N_13554);
nand U13661 (N_13661,N_13553,N_13527);
xor U13662 (N_13662,N_13545,N_13602);
nor U13663 (N_13663,N_13579,N_13515);
and U13664 (N_13664,N_13596,N_13590);
and U13665 (N_13665,N_13538,N_13508);
and U13666 (N_13666,N_13531,N_13611);
nor U13667 (N_13667,N_13524,N_13576);
and U13668 (N_13668,N_13556,N_13541);
xnor U13669 (N_13669,N_13594,N_13511);
or U13670 (N_13670,N_13588,N_13530);
and U13671 (N_13671,N_13528,N_13525);
and U13672 (N_13672,N_13509,N_13573);
xor U13673 (N_13673,N_13565,N_13558);
or U13674 (N_13674,N_13504,N_13542);
nand U13675 (N_13675,N_13616,N_13600);
nor U13676 (N_13676,N_13546,N_13572);
nand U13677 (N_13677,N_13581,N_13569);
nand U13678 (N_13678,N_13548,N_13584);
xor U13679 (N_13679,N_13607,N_13562);
xnor U13680 (N_13680,N_13534,N_13523);
xor U13681 (N_13681,N_13519,N_13549);
and U13682 (N_13682,N_13526,N_13571);
and U13683 (N_13683,N_13592,N_13566);
or U13684 (N_13684,N_13589,N_13555);
nand U13685 (N_13685,N_13563,N_13560);
or U13686 (N_13686,N_13582,N_13577);
nor U13687 (N_13687,N_13622,N_13516);
nor U13688 (N_13688,N_13523,N_13591);
nand U13689 (N_13689,N_13552,N_13584);
and U13690 (N_13690,N_13510,N_13613);
and U13691 (N_13691,N_13535,N_13523);
nand U13692 (N_13692,N_13603,N_13537);
nor U13693 (N_13693,N_13589,N_13570);
or U13694 (N_13694,N_13543,N_13557);
nand U13695 (N_13695,N_13574,N_13528);
nand U13696 (N_13696,N_13560,N_13593);
nor U13697 (N_13697,N_13516,N_13500);
and U13698 (N_13698,N_13619,N_13516);
nand U13699 (N_13699,N_13520,N_13582);
or U13700 (N_13700,N_13551,N_13593);
nand U13701 (N_13701,N_13526,N_13566);
and U13702 (N_13702,N_13536,N_13608);
and U13703 (N_13703,N_13540,N_13560);
xnor U13704 (N_13704,N_13541,N_13620);
or U13705 (N_13705,N_13522,N_13500);
or U13706 (N_13706,N_13503,N_13586);
or U13707 (N_13707,N_13528,N_13521);
nor U13708 (N_13708,N_13614,N_13513);
and U13709 (N_13709,N_13546,N_13545);
nand U13710 (N_13710,N_13617,N_13552);
xnor U13711 (N_13711,N_13587,N_13601);
or U13712 (N_13712,N_13520,N_13523);
nor U13713 (N_13713,N_13588,N_13624);
and U13714 (N_13714,N_13589,N_13520);
nand U13715 (N_13715,N_13538,N_13544);
nor U13716 (N_13716,N_13603,N_13516);
nand U13717 (N_13717,N_13543,N_13606);
nor U13718 (N_13718,N_13530,N_13571);
and U13719 (N_13719,N_13584,N_13583);
xnor U13720 (N_13720,N_13619,N_13562);
nand U13721 (N_13721,N_13574,N_13557);
and U13722 (N_13722,N_13583,N_13595);
xnor U13723 (N_13723,N_13507,N_13554);
or U13724 (N_13724,N_13618,N_13507);
nor U13725 (N_13725,N_13578,N_13617);
nand U13726 (N_13726,N_13513,N_13507);
and U13727 (N_13727,N_13615,N_13607);
xnor U13728 (N_13728,N_13541,N_13606);
nor U13729 (N_13729,N_13595,N_13528);
and U13730 (N_13730,N_13602,N_13583);
xnor U13731 (N_13731,N_13560,N_13537);
and U13732 (N_13732,N_13518,N_13541);
and U13733 (N_13733,N_13509,N_13613);
nand U13734 (N_13734,N_13580,N_13531);
or U13735 (N_13735,N_13561,N_13516);
and U13736 (N_13736,N_13585,N_13555);
nor U13737 (N_13737,N_13571,N_13592);
xor U13738 (N_13738,N_13603,N_13600);
xor U13739 (N_13739,N_13540,N_13507);
xor U13740 (N_13740,N_13527,N_13510);
xor U13741 (N_13741,N_13508,N_13523);
and U13742 (N_13742,N_13564,N_13515);
and U13743 (N_13743,N_13574,N_13570);
or U13744 (N_13744,N_13543,N_13615);
xor U13745 (N_13745,N_13584,N_13517);
nand U13746 (N_13746,N_13582,N_13619);
or U13747 (N_13747,N_13610,N_13506);
or U13748 (N_13748,N_13550,N_13578);
xor U13749 (N_13749,N_13538,N_13547);
nor U13750 (N_13750,N_13691,N_13746);
or U13751 (N_13751,N_13715,N_13641);
nand U13752 (N_13752,N_13717,N_13693);
xnor U13753 (N_13753,N_13663,N_13630);
nor U13754 (N_13754,N_13634,N_13666);
nand U13755 (N_13755,N_13657,N_13731);
and U13756 (N_13756,N_13643,N_13709);
or U13757 (N_13757,N_13724,N_13696);
or U13758 (N_13758,N_13627,N_13711);
nand U13759 (N_13759,N_13727,N_13682);
nand U13760 (N_13760,N_13637,N_13674);
nand U13761 (N_13761,N_13739,N_13676);
nand U13762 (N_13762,N_13699,N_13667);
and U13763 (N_13763,N_13644,N_13672);
xor U13764 (N_13764,N_13688,N_13648);
and U13765 (N_13765,N_13629,N_13707);
or U13766 (N_13766,N_13675,N_13636);
xnor U13767 (N_13767,N_13661,N_13652);
and U13768 (N_13768,N_13744,N_13705);
and U13769 (N_13769,N_13633,N_13635);
nand U13770 (N_13770,N_13710,N_13665);
or U13771 (N_13771,N_13712,N_13720);
and U13772 (N_13772,N_13730,N_13698);
nand U13773 (N_13773,N_13726,N_13631);
or U13774 (N_13774,N_13694,N_13639);
nor U13775 (N_13775,N_13654,N_13677);
nand U13776 (N_13776,N_13695,N_13625);
nor U13777 (N_13777,N_13734,N_13683);
or U13778 (N_13778,N_13626,N_13743);
and U13779 (N_13779,N_13745,N_13701);
and U13780 (N_13780,N_13653,N_13718);
xor U13781 (N_13781,N_13700,N_13687);
xor U13782 (N_13782,N_13640,N_13685);
nand U13783 (N_13783,N_13690,N_13662);
nand U13784 (N_13784,N_13741,N_13702);
xnor U13785 (N_13785,N_13673,N_13689);
nand U13786 (N_13786,N_13722,N_13658);
or U13787 (N_13787,N_13728,N_13738);
nor U13788 (N_13788,N_13681,N_13628);
nor U13789 (N_13789,N_13729,N_13748);
nand U13790 (N_13790,N_13642,N_13638);
nor U13791 (N_13791,N_13692,N_13723);
nand U13792 (N_13792,N_13679,N_13732);
and U13793 (N_13793,N_13740,N_13706);
or U13794 (N_13794,N_13659,N_13664);
nand U13795 (N_13795,N_13651,N_13735);
nand U13796 (N_13796,N_13697,N_13713);
or U13797 (N_13797,N_13646,N_13655);
nand U13798 (N_13798,N_13737,N_13736);
and U13799 (N_13799,N_13725,N_13714);
nor U13800 (N_13800,N_13650,N_13632);
nand U13801 (N_13801,N_13719,N_13716);
xor U13802 (N_13802,N_13656,N_13649);
and U13803 (N_13803,N_13742,N_13721);
xor U13804 (N_13804,N_13703,N_13670);
nand U13805 (N_13805,N_13647,N_13749);
or U13806 (N_13806,N_13747,N_13684);
nor U13807 (N_13807,N_13708,N_13678);
xor U13808 (N_13808,N_13669,N_13668);
nor U13809 (N_13809,N_13686,N_13704);
nor U13810 (N_13810,N_13645,N_13733);
nand U13811 (N_13811,N_13671,N_13660);
nand U13812 (N_13812,N_13680,N_13729);
or U13813 (N_13813,N_13659,N_13663);
xor U13814 (N_13814,N_13698,N_13715);
or U13815 (N_13815,N_13695,N_13629);
xnor U13816 (N_13816,N_13694,N_13721);
xnor U13817 (N_13817,N_13650,N_13640);
or U13818 (N_13818,N_13737,N_13693);
nor U13819 (N_13819,N_13714,N_13734);
nand U13820 (N_13820,N_13632,N_13674);
and U13821 (N_13821,N_13670,N_13674);
xor U13822 (N_13822,N_13637,N_13682);
xor U13823 (N_13823,N_13690,N_13710);
and U13824 (N_13824,N_13647,N_13748);
or U13825 (N_13825,N_13689,N_13633);
nor U13826 (N_13826,N_13645,N_13730);
or U13827 (N_13827,N_13729,N_13635);
or U13828 (N_13828,N_13681,N_13640);
or U13829 (N_13829,N_13715,N_13701);
nor U13830 (N_13830,N_13666,N_13722);
nand U13831 (N_13831,N_13736,N_13658);
or U13832 (N_13832,N_13722,N_13656);
nor U13833 (N_13833,N_13684,N_13625);
nand U13834 (N_13834,N_13734,N_13695);
xnor U13835 (N_13835,N_13730,N_13664);
and U13836 (N_13836,N_13685,N_13728);
or U13837 (N_13837,N_13638,N_13695);
nor U13838 (N_13838,N_13680,N_13712);
nor U13839 (N_13839,N_13713,N_13630);
and U13840 (N_13840,N_13681,N_13705);
nand U13841 (N_13841,N_13660,N_13673);
nor U13842 (N_13842,N_13646,N_13727);
nand U13843 (N_13843,N_13687,N_13740);
and U13844 (N_13844,N_13710,N_13737);
nor U13845 (N_13845,N_13711,N_13632);
nand U13846 (N_13846,N_13746,N_13673);
or U13847 (N_13847,N_13645,N_13719);
xnor U13848 (N_13848,N_13713,N_13749);
or U13849 (N_13849,N_13695,N_13641);
nor U13850 (N_13850,N_13691,N_13741);
or U13851 (N_13851,N_13649,N_13658);
or U13852 (N_13852,N_13684,N_13726);
nor U13853 (N_13853,N_13638,N_13669);
nand U13854 (N_13854,N_13653,N_13701);
xnor U13855 (N_13855,N_13694,N_13719);
or U13856 (N_13856,N_13731,N_13710);
or U13857 (N_13857,N_13741,N_13729);
nor U13858 (N_13858,N_13681,N_13738);
or U13859 (N_13859,N_13636,N_13711);
nand U13860 (N_13860,N_13651,N_13742);
or U13861 (N_13861,N_13663,N_13735);
or U13862 (N_13862,N_13674,N_13748);
and U13863 (N_13863,N_13734,N_13661);
xnor U13864 (N_13864,N_13699,N_13627);
or U13865 (N_13865,N_13629,N_13733);
nor U13866 (N_13866,N_13694,N_13744);
or U13867 (N_13867,N_13686,N_13703);
or U13868 (N_13868,N_13716,N_13744);
nand U13869 (N_13869,N_13659,N_13730);
xnor U13870 (N_13870,N_13741,N_13680);
and U13871 (N_13871,N_13652,N_13714);
and U13872 (N_13872,N_13731,N_13629);
nor U13873 (N_13873,N_13713,N_13693);
nor U13874 (N_13874,N_13668,N_13638);
nor U13875 (N_13875,N_13775,N_13790);
or U13876 (N_13876,N_13769,N_13805);
or U13877 (N_13877,N_13752,N_13755);
nand U13878 (N_13878,N_13801,N_13840);
nor U13879 (N_13879,N_13868,N_13847);
and U13880 (N_13880,N_13866,N_13807);
or U13881 (N_13881,N_13750,N_13844);
or U13882 (N_13882,N_13864,N_13767);
and U13883 (N_13883,N_13802,N_13781);
and U13884 (N_13884,N_13776,N_13788);
nor U13885 (N_13885,N_13861,N_13819);
nand U13886 (N_13886,N_13772,N_13867);
nor U13887 (N_13887,N_13850,N_13773);
and U13888 (N_13888,N_13761,N_13827);
and U13889 (N_13889,N_13838,N_13785);
or U13890 (N_13890,N_13835,N_13809);
nand U13891 (N_13891,N_13799,N_13758);
nand U13892 (N_13892,N_13810,N_13791);
xor U13893 (N_13893,N_13831,N_13806);
nand U13894 (N_13894,N_13762,N_13869);
nand U13895 (N_13895,N_13856,N_13778);
and U13896 (N_13896,N_13820,N_13872);
or U13897 (N_13897,N_13789,N_13765);
xnor U13898 (N_13898,N_13766,N_13759);
or U13899 (N_13899,N_13754,N_13782);
xor U13900 (N_13900,N_13841,N_13796);
nand U13901 (N_13901,N_13860,N_13795);
and U13902 (N_13902,N_13792,N_13859);
nor U13903 (N_13903,N_13824,N_13794);
nand U13904 (N_13904,N_13821,N_13822);
nand U13905 (N_13905,N_13839,N_13828);
nand U13906 (N_13906,N_13798,N_13811);
nand U13907 (N_13907,N_13849,N_13757);
and U13908 (N_13908,N_13783,N_13817);
and U13909 (N_13909,N_13818,N_13857);
or U13910 (N_13910,N_13768,N_13763);
and U13911 (N_13911,N_13756,N_13764);
nor U13912 (N_13912,N_13854,N_13846);
nand U13913 (N_13913,N_13804,N_13753);
nand U13914 (N_13914,N_13863,N_13833);
nand U13915 (N_13915,N_13855,N_13770);
nand U13916 (N_13916,N_13845,N_13843);
nor U13917 (N_13917,N_13813,N_13834);
and U13918 (N_13918,N_13816,N_13842);
nor U13919 (N_13919,N_13829,N_13865);
nand U13920 (N_13920,N_13797,N_13832);
nor U13921 (N_13921,N_13786,N_13830);
or U13922 (N_13922,N_13852,N_13851);
xnor U13923 (N_13923,N_13771,N_13793);
xnor U13924 (N_13924,N_13848,N_13774);
or U13925 (N_13925,N_13784,N_13836);
nor U13926 (N_13926,N_13825,N_13837);
and U13927 (N_13927,N_13826,N_13871);
and U13928 (N_13928,N_13873,N_13803);
nor U13929 (N_13929,N_13787,N_13751);
nand U13930 (N_13930,N_13853,N_13812);
nor U13931 (N_13931,N_13777,N_13800);
and U13932 (N_13932,N_13760,N_13823);
xor U13933 (N_13933,N_13858,N_13780);
and U13934 (N_13934,N_13874,N_13814);
and U13935 (N_13935,N_13808,N_13870);
and U13936 (N_13936,N_13815,N_13862);
xor U13937 (N_13937,N_13779,N_13838);
or U13938 (N_13938,N_13782,N_13799);
xor U13939 (N_13939,N_13797,N_13815);
nor U13940 (N_13940,N_13822,N_13865);
and U13941 (N_13941,N_13821,N_13788);
nand U13942 (N_13942,N_13783,N_13864);
xor U13943 (N_13943,N_13756,N_13871);
and U13944 (N_13944,N_13801,N_13761);
nand U13945 (N_13945,N_13869,N_13759);
or U13946 (N_13946,N_13859,N_13816);
or U13947 (N_13947,N_13807,N_13763);
nand U13948 (N_13948,N_13771,N_13800);
xor U13949 (N_13949,N_13850,N_13776);
and U13950 (N_13950,N_13776,N_13834);
nor U13951 (N_13951,N_13791,N_13814);
and U13952 (N_13952,N_13784,N_13778);
or U13953 (N_13953,N_13842,N_13834);
or U13954 (N_13954,N_13762,N_13840);
or U13955 (N_13955,N_13785,N_13824);
xor U13956 (N_13956,N_13806,N_13867);
nand U13957 (N_13957,N_13782,N_13785);
or U13958 (N_13958,N_13774,N_13866);
xor U13959 (N_13959,N_13825,N_13751);
nand U13960 (N_13960,N_13773,N_13757);
xnor U13961 (N_13961,N_13799,N_13873);
nor U13962 (N_13962,N_13828,N_13806);
and U13963 (N_13963,N_13816,N_13786);
or U13964 (N_13964,N_13808,N_13788);
xor U13965 (N_13965,N_13767,N_13802);
or U13966 (N_13966,N_13812,N_13835);
nand U13967 (N_13967,N_13868,N_13840);
xor U13968 (N_13968,N_13808,N_13795);
and U13969 (N_13969,N_13843,N_13846);
or U13970 (N_13970,N_13793,N_13818);
xor U13971 (N_13971,N_13830,N_13796);
or U13972 (N_13972,N_13783,N_13862);
and U13973 (N_13973,N_13872,N_13815);
xnor U13974 (N_13974,N_13847,N_13778);
and U13975 (N_13975,N_13870,N_13765);
and U13976 (N_13976,N_13768,N_13842);
xor U13977 (N_13977,N_13822,N_13797);
xnor U13978 (N_13978,N_13806,N_13819);
and U13979 (N_13979,N_13762,N_13852);
and U13980 (N_13980,N_13848,N_13810);
nand U13981 (N_13981,N_13772,N_13750);
nor U13982 (N_13982,N_13852,N_13812);
nor U13983 (N_13983,N_13788,N_13874);
nor U13984 (N_13984,N_13845,N_13750);
or U13985 (N_13985,N_13765,N_13869);
nand U13986 (N_13986,N_13819,N_13868);
nor U13987 (N_13987,N_13801,N_13757);
or U13988 (N_13988,N_13859,N_13791);
nand U13989 (N_13989,N_13855,N_13814);
or U13990 (N_13990,N_13849,N_13833);
and U13991 (N_13991,N_13758,N_13772);
and U13992 (N_13992,N_13839,N_13835);
nor U13993 (N_13993,N_13770,N_13872);
and U13994 (N_13994,N_13822,N_13804);
xnor U13995 (N_13995,N_13766,N_13820);
xor U13996 (N_13996,N_13774,N_13789);
or U13997 (N_13997,N_13829,N_13854);
or U13998 (N_13998,N_13760,N_13820);
nor U13999 (N_13999,N_13827,N_13838);
xnor U14000 (N_14000,N_13907,N_13946);
xor U14001 (N_14001,N_13915,N_13959);
nor U14002 (N_14002,N_13958,N_13994);
xnor U14003 (N_14003,N_13929,N_13914);
xor U14004 (N_14004,N_13970,N_13876);
nand U14005 (N_14005,N_13913,N_13947);
or U14006 (N_14006,N_13996,N_13896);
nor U14007 (N_14007,N_13980,N_13988);
nor U14008 (N_14008,N_13995,N_13962);
nor U14009 (N_14009,N_13880,N_13993);
xnor U14010 (N_14010,N_13930,N_13983);
nor U14011 (N_14011,N_13977,N_13926);
xor U14012 (N_14012,N_13903,N_13881);
nand U14013 (N_14013,N_13890,N_13968);
nand U14014 (N_14014,N_13900,N_13951);
nor U14015 (N_14015,N_13992,N_13948);
and U14016 (N_14016,N_13935,N_13888);
nor U14017 (N_14017,N_13942,N_13990);
nor U14018 (N_14018,N_13899,N_13918);
xor U14019 (N_14019,N_13895,N_13953);
nand U14020 (N_14020,N_13908,N_13911);
nand U14021 (N_14021,N_13875,N_13941);
or U14022 (N_14022,N_13904,N_13998);
and U14023 (N_14023,N_13957,N_13940);
nand U14024 (N_14024,N_13969,N_13887);
nand U14025 (N_14025,N_13949,N_13933);
xnor U14026 (N_14026,N_13905,N_13960);
nor U14027 (N_14027,N_13938,N_13989);
or U14028 (N_14028,N_13923,N_13909);
and U14029 (N_14029,N_13902,N_13950);
nand U14030 (N_14030,N_13936,N_13885);
and U14031 (N_14031,N_13964,N_13879);
xnor U14032 (N_14032,N_13987,N_13906);
nor U14033 (N_14033,N_13932,N_13943);
and U14034 (N_14034,N_13955,N_13891);
nor U14035 (N_14035,N_13975,N_13889);
xor U14036 (N_14036,N_13910,N_13997);
nor U14037 (N_14037,N_13893,N_13877);
xnor U14038 (N_14038,N_13898,N_13920);
xnor U14039 (N_14039,N_13919,N_13928);
nor U14040 (N_14040,N_13965,N_13901);
nand U14041 (N_14041,N_13967,N_13884);
xnor U14042 (N_14042,N_13917,N_13937);
nor U14043 (N_14043,N_13921,N_13974);
and U14044 (N_14044,N_13883,N_13981);
nand U14045 (N_14045,N_13963,N_13924);
xor U14046 (N_14046,N_13945,N_13897);
xnor U14047 (N_14047,N_13886,N_13939);
or U14048 (N_14048,N_13952,N_13916);
nand U14049 (N_14049,N_13954,N_13956);
xnor U14050 (N_14050,N_13931,N_13966);
and U14051 (N_14051,N_13971,N_13972);
nor U14052 (N_14052,N_13991,N_13878);
nand U14053 (N_14053,N_13934,N_13976);
xnor U14054 (N_14054,N_13961,N_13979);
and U14055 (N_14055,N_13925,N_13892);
nand U14056 (N_14056,N_13922,N_13973);
or U14057 (N_14057,N_13985,N_13944);
xnor U14058 (N_14058,N_13912,N_13999);
or U14059 (N_14059,N_13986,N_13894);
xor U14060 (N_14060,N_13984,N_13978);
and U14061 (N_14061,N_13927,N_13982);
or U14062 (N_14062,N_13882,N_13997);
and U14063 (N_14063,N_13978,N_13988);
or U14064 (N_14064,N_13959,N_13991);
nor U14065 (N_14065,N_13971,N_13904);
xor U14066 (N_14066,N_13961,N_13950);
or U14067 (N_14067,N_13956,N_13910);
nor U14068 (N_14068,N_13914,N_13972);
nand U14069 (N_14069,N_13995,N_13917);
and U14070 (N_14070,N_13878,N_13888);
nand U14071 (N_14071,N_13944,N_13951);
or U14072 (N_14072,N_13925,N_13961);
xor U14073 (N_14073,N_13985,N_13973);
nor U14074 (N_14074,N_13962,N_13882);
xnor U14075 (N_14075,N_13952,N_13892);
and U14076 (N_14076,N_13990,N_13915);
xor U14077 (N_14077,N_13913,N_13879);
nor U14078 (N_14078,N_13990,N_13888);
or U14079 (N_14079,N_13881,N_13885);
and U14080 (N_14080,N_13991,N_13890);
or U14081 (N_14081,N_13983,N_13896);
nand U14082 (N_14082,N_13948,N_13981);
or U14083 (N_14083,N_13968,N_13963);
nand U14084 (N_14084,N_13988,N_13918);
nor U14085 (N_14085,N_13886,N_13976);
nand U14086 (N_14086,N_13900,N_13998);
xnor U14087 (N_14087,N_13898,N_13959);
xor U14088 (N_14088,N_13896,N_13916);
nor U14089 (N_14089,N_13952,N_13932);
nand U14090 (N_14090,N_13984,N_13947);
xnor U14091 (N_14091,N_13887,N_13992);
or U14092 (N_14092,N_13905,N_13878);
or U14093 (N_14093,N_13891,N_13972);
or U14094 (N_14094,N_13902,N_13982);
nand U14095 (N_14095,N_13943,N_13941);
or U14096 (N_14096,N_13881,N_13970);
xor U14097 (N_14097,N_13904,N_13994);
nor U14098 (N_14098,N_13974,N_13951);
or U14099 (N_14099,N_13971,N_13897);
nor U14100 (N_14100,N_13924,N_13907);
nor U14101 (N_14101,N_13912,N_13896);
nor U14102 (N_14102,N_13910,N_13898);
nor U14103 (N_14103,N_13914,N_13979);
xor U14104 (N_14104,N_13934,N_13940);
nand U14105 (N_14105,N_13908,N_13900);
or U14106 (N_14106,N_13988,N_13899);
and U14107 (N_14107,N_13986,N_13995);
xnor U14108 (N_14108,N_13927,N_13890);
xor U14109 (N_14109,N_13976,N_13883);
nand U14110 (N_14110,N_13971,N_13990);
nor U14111 (N_14111,N_13972,N_13966);
or U14112 (N_14112,N_13915,N_13884);
xnor U14113 (N_14113,N_13956,N_13876);
or U14114 (N_14114,N_13891,N_13910);
nor U14115 (N_14115,N_13957,N_13975);
xor U14116 (N_14116,N_13946,N_13949);
or U14117 (N_14117,N_13984,N_13960);
and U14118 (N_14118,N_13955,N_13898);
or U14119 (N_14119,N_13940,N_13969);
nand U14120 (N_14120,N_13884,N_13957);
xnor U14121 (N_14121,N_13983,N_13919);
or U14122 (N_14122,N_13889,N_13937);
or U14123 (N_14123,N_13922,N_13992);
xnor U14124 (N_14124,N_13954,N_13920);
nand U14125 (N_14125,N_14124,N_14036);
nand U14126 (N_14126,N_14025,N_14033);
and U14127 (N_14127,N_14063,N_14110);
and U14128 (N_14128,N_14048,N_14089);
nand U14129 (N_14129,N_14093,N_14106);
or U14130 (N_14130,N_14068,N_14045);
nand U14131 (N_14131,N_14051,N_14069);
and U14132 (N_14132,N_14088,N_14043);
or U14133 (N_14133,N_14072,N_14001);
xnor U14134 (N_14134,N_14018,N_14096);
and U14135 (N_14135,N_14003,N_14105);
and U14136 (N_14136,N_14019,N_14080);
nand U14137 (N_14137,N_14037,N_14079);
or U14138 (N_14138,N_14076,N_14087);
and U14139 (N_14139,N_14057,N_14059);
xnor U14140 (N_14140,N_14021,N_14086);
or U14141 (N_14141,N_14008,N_14010);
nand U14142 (N_14142,N_14119,N_14074);
or U14143 (N_14143,N_14012,N_14009);
nor U14144 (N_14144,N_14042,N_14077);
xor U14145 (N_14145,N_14100,N_14041);
xor U14146 (N_14146,N_14030,N_14116);
xnor U14147 (N_14147,N_14084,N_14066);
or U14148 (N_14148,N_14052,N_14095);
xnor U14149 (N_14149,N_14017,N_14058);
nand U14150 (N_14150,N_14115,N_14090);
and U14151 (N_14151,N_14028,N_14082);
or U14152 (N_14152,N_14007,N_14044);
and U14153 (N_14153,N_14014,N_14020);
xor U14154 (N_14154,N_14081,N_14002);
and U14155 (N_14155,N_14098,N_14073);
nor U14156 (N_14156,N_14099,N_14047);
nor U14157 (N_14157,N_14092,N_14065);
or U14158 (N_14158,N_14109,N_14085);
nand U14159 (N_14159,N_14078,N_14102);
or U14160 (N_14160,N_14123,N_14050);
or U14161 (N_14161,N_14111,N_14006);
nor U14162 (N_14162,N_14013,N_14094);
nand U14163 (N_14163,N_14062,N_14061);
nand U14164 (N_14164,N_14070,N_14113);
or U14165 (N_14165,N_14083,N_14122);
nand U14166 (N_14166,N_14114,N_14053);
or U14167 (N_14167,N_14040,N_14027);
nor U14168 (N_14168,N_14004,N_14024);
nor U14169 (N_14169,N_14049,N_14064);
and U14170 (N_14170,N_14075,N_14032);
and U14171 (N_14171,N_14016,N_14035);
and U14172 (N_14172,N_14026,N_14091);
or U14173 (N_14173,N_14067,N_14117);
nor U14174 (N_14174,N_14034,N_14118);
nand U14175 (N_14175,N_14038,N_14101);
nor U14176 (N_14176,N_14005,N_14011);
and U14177 (N_14177,N_14056,N_14121);
and U14178 (N_14178,N_14029,N_14031);
xor U14179 (N_14179,N_14108,N_14054);
nand U14180 (N_14180,N_14097,N_14104);
nor U14181 (N_14181,N_14055,N_14120);
nor U14182 (N_14182,N_14022,N_14071);
nand U14183 (N_14183,N_14112,N_14103);
or U14184 (N_14184,N_14046,N_14015);
nand U14185 (N_14185,N_14000,N_14060);
nand U14186 (N_14186,N_14039,N_14023);
and U14187 (N_14187,N_14107,N_14065);
nor U14188 (N_14188,N_14110,N_14016);
and U14189 (N_14189,N_14025,N_14117);
nand U14190 (N_14190,N_14071,N_14081);
or U14191 (N_14191,N_14087,N_14089);
nand U14192 (N_14192,N_14112,N_14075);
and U14193 (N_14193,N_14105,N_14007);
nor U14194 (N_14194,N_14122,N_14113);
or U14195 (N_14195,N_14033,N_14023);
and U14196 (N_14196,N_14093,N_14116);
nand U14197 (N_14197,N_14032,N_14006);
or U14198 (N_14198,N_14092,N_14037);
or U14199 (N_14199,N_14123,N_14117);
and U14200 (N_14200,N_14026,N_14085);
xor U14201 (N_14201,N_14047,N_14055);
nor U14202 (N_14202,N_14108,N_14026);
xor U14203 (N_14203,N_14045,N_14075);
nand U14204 (N_14204,N_14060,N_14080);
or U14205 (N_14205,N_14056,N_14030);
or U14206 (N_14206,N_14061,N_14058);
nor U14207 (N_14207,N_14005,N_14004);
xor U14208 (N_14208,N_14009,N_14088);
and U14209 (N_14209,N_14116,N_14115);
and U14210 (N_14210,N_14112,N_14061);
or U14211 (N_14211,N_14007,N_14056);
xnor U14212 (N_14212,N_14101,N_14004);
or U14213 (N_14213,N_14110,N_14031);
nor U14214 (N_14214,N_14124,N_14061);
nor U14215 (N_14215,N_14069,N_14111);
and U14216 (N_14216,N_14001,N_14087);
or U14217 (N_14217,N_14073,N_14046);
nor U14218 (N_14218,N_14093,N_14050);
nand U14219 (N_14219,N_14081,N_14107);
nor U14220 (N_14220,N_14062,N_14098);
nand U14221 (N_14221,N_14090,N_14065);
or U14222 (N_14222,N_14087,N_14121);
xnor U14223 (N_14223,N_14104,N_14091);
or U14224 (N_14224,N_14014,N_14019);
xnor U14225 (N_14225,N_14036,N_14118);
nand U14226 (N_14226,N_14105,N_14062);
or U14227 (N_14227,N_14007,N_14010);
nor U14228 (N_14228,N_14002,N_14054);
nand U14229 (N_14229,N_14022,N_14012);
xnor U14230 (N_14230,N_14038,N_14097);
xnor U14231 (N_14231,N_14103,N_14106);
nand U14232 (N_14232,N_14080,N_14044);
or U14233 (N_14233,N_14090,N_14109);
and U14234 (N_14234,N_14020,N_14078);
xnor U14235 (N_14235,N_14072,N_14005);
and U14236 (N_14236,N_14086,N_14103);
nand U14237 (N_14237,N_14071,N_14034);
or U14238 (N_14238,N_14097,N_14080);
or U14239 (N_14239,N_14082,N_14102);
nor U14240 (N_14240,N_14074,N_14002);
nand U14241 (N_14241,N_14041,N_14000);
and U14242 (N_14242,N_14078,N_14077);
nand U14243 (N_14243,N_14061,N_14045);
xor U14244 (N_14244,N_14118,N_14029);
nor U14245 (N_14245,N_14014,N_14023);
xnor U14246 (N_14246,N_14045,N_14065);
xnor U14247 (N_14247,N_14090,N_14103);
nor U14248 (N_14248,N_14031,N_14034);
or U14249 (N_14249,N_14080,N_14090);
and U14250 (N_14250,N_14138,N_14125);
and U14251 (N_14251,N_14141,N_14220);
nor U14252 (N_14252,N_14156,N_14207);
or U14253 (N_14253,N_14153,N_14175);
nor U14254 (N_14254,N_14139,N_14247);
xnor U14255 (N_14255,N_14239,N_14228);
and U14256 (N_14256,N_14197,N_14238);
xnor U14257 (N_14257,N_14164,N_14200);
and U14258 (N_14258,N_14204,N_14174);
nor U14259 (N_14259,N_14243,N_14151);
or U14260 (N_14260,N_14245,N_14193);
xor U14261 (N_14261,N_14183,N_14190);
and U14262 (N_14262,N_14231,N_14201);
xnor U14263 (N_14263,N_14154,N_14214);
nand U14264 (N_14264,N_14180,N_14194);
nor U14265 (N_14265,N_14127,N_14130);
nor U14266 (N_14266,N_14129,N_14215);
xor U14267 (N_14267,N_14167,N_14165);
and U14268 (N_14268,N_14218,N_14172);
nand U14269 (N_14269,N_14150,N_14142);
xnor U14270 (N_14270,N_14176,N_14186);
or U14271 (N_14271,N_14248,N_14226);
and U14272 (N_14272,N_14152,N_14162);
and U14273 (N_14273,N_14241,N_14136);
xnor U14274 (N_14274,N_14206,N_14184);
or U14275 (N_14275,N_14211,N_14224);
or U14276 (N_14276,N_14232,N_14143);
nand U14277 (N_14277,N_14229,N_14182);
and U14278 (N_14278,N_14179,N_14168);
or U14279 (N_14279,N_14192,N_14210);
xnor U14280 (N_14280,N_14219,N_14170);
nand U14281 (N_14281,N_14134,N_14177);
and U14282 (N_14282,N_14155,N_14133);
nand U14283 (N_14283,N_14242,N_14209);
nand U14284 (N_14284,N_14149,N_14185);
and U14285 (N_14285,N_14159,N_14249);
and U14286 (N_14286,N_14246,N_14233);
or U14287 (N_14287,N_14208,N_14198);
and U14288 (N_14288,N_14145,N_14160);
nor U14289 (N_14289,N_14158,N_14216);
nand U14290 (N_14290,N_14166,N_14181);
xnor U14291 (N_14291,N_14178,N_14234);
nor U14292 (N_14292,N_14157,N_14230);
nor U14293 (N_14293,N_14128,N_14169);
or U14294 (N_14294,N_14240,N_14222);
and U14295 (N_14295,N_14188,N_14135);
nand U14296 (N_14296,N_14173,N_14202);
and U14297 (N_14297,N_14213,N_14131);
xnor U14298 (N_14298,N_14195,N_14140);
or U14299 (N_14299,N_14161,N_14146);
xnor U14300 (N_14300,N_14163,N_14199);
nor U14301 (N_14301,N_14187,N_14144);
and U14302 (N_14302,N_14205,N_14212);
and U14303 (N_14303,N_14196,N_14148);
and U14304 (N_14304,N_14244,N_14137);
xor U14305 (N_14305,N_14225,N_14235);
nor U14306 (N_14306,N_14237,N_14227);
or U14307 (N_14307,N_14203,N_14189);
or U14308 (N_14308,N_14236,N_14191);
or U14309 (N_14309,N_14223,N_14171);
or U14310 (N_14310,N_14132,N_14217);
xor U14311 (N_14311,N_14126,N_14147);
nand U14312 (N_14312,N_14221,N_14219);
nor U14313 (N_14313,N_14164,N_14173);
nor U14314 (N_14314,N_14246,N_14158);
and U14315 (N_14315,N_14232,N_14144);
nand U14316 (N_14316,N_14134,N_14200);
or U14317 (N_14317,N_14189,N_14158);
xor U14318 (N_14318,N_14180,N_14178);
nor U14319 (N_14319,N_14126,N_14244);
and U14320 (N_14320,N_14151,N_14132);
nand U14321 (N_14321,N_14128,N_14202);
xor U14322 (N_14322,N_14217,N_14198);
and U14323 (N_14323,N_14142,N_14238);
xor U14324 (N_14324,N_14135,N_14152);
nand U14325 (N_14325,N_14142,N_14141);
nor U14326 (N_14326,N_14158,N_14209);
nand U14327 (N_14327,N_14196,N_14190);
xnor U14328 (N_14328,N_14125,N_14227);
nor U14329 (N_14329,N_14214,N_14150);
nand U14330 (N_14330,N_14230,N_14191);
nand U14331 (N_14331,N_14195,N_14156);
or U14332 (N_14332,N_14248,N_14179);
or U14333 (N_14333,N_14188,N_14196);
and U14334 (N_14334,N_14223,N_14231);
xnor U14335 (N_14335,N_14133,N_14195);
xor U14336 (N_14336,N_14140,N_14213);
or U14337 (N_14337,N_14206,N_14191);
nand U14338 (N_14338,N_14129,N_14217);
and U14339 (N_14339,N_14193,N_14246);
nand U14340 (N_14340,N_14192,N_14183);
and U14341 (N_14341,N_14200,N_14199);
or U14342 (N_14342,N_14126,N_14176);
and U14343 (N_14343,N_14149,N_14240);
or U14344 (N_14344,N_14245,N_14232);
xor U14345 (N_14345,N_14133,N_14148);
xnor U14346 (N_14346,N_14192,N_14204);
or U14347 (N_14347,N_14224,N_14158);
xor U14348 (N_14348,N_14228,N_14245);
and U14349 (N_14349,N_14139,N_14164);
or U14350 (N_14350,N_14244,N_14206);
xnor U14351 (N_14351,N_14175,N_14146);
and U14352 (N_14352,N_14135,N_14141);
and U14353 (N_14353,N_14154,N_14208);
nor U14354 (N_14354,N_14246,N_14128);
nand U14355 (N_14355,N_14212,N_14193);
xor U14356 (N_14356,N_14187,N_14203);
and U14357 (N_14357,N_14246,N_14221);
xor U14358 (N_14358,N_14245,N_14236);
or U14359 (N_14359,N_14183,N_14240);
nor U14360 (N_14360,N_14236,N_14220);
or U14361 (N_14361,N_14195,N_14229);
nor U14362 (N_14362,N_14196,N_14242);
nand U14363 (N_14363,N_14190,N_14143);
xor U14364 (N_14364,N_14163,N_14157);
or U14365 (N_14365,N_14164,N_14225);
xor U14366 (N_14366,N_14206,N_14173);
xor U14367 (N_14367,N_14171,N_14142);
xor U14368 (N_14368,N_14179,N_14241);
xor U14369 (N_14369,N_14238,N_14236);
xnor U14370 (N_14370,N_14128,N_14147);
nand U14371 (N_14371,N_14247,N_14235);
or U14372 (N_14372,N_14173,N_14184);
and U14373 (N_14373,N_14243,N_14170);
or U14374 (N_14374,N_14133,N_14181);
nor U14375 (N_14375,N_14276,N_14286);
or U14376 (N_14376,N_14265,N_14255);
xnor U14377 (N_14377,N_14284,N_14343);
or U14378 (N_14378,N_14351,N_14317);
and U14379 (N_14379,N_14269,N_14352);
or U14380 (N_14380,N_14369,N_14282);
and U14381 (N_14381,N_14370,N_14260);
and U14382 (N_14382,N_14258,N_14318);
or U14383 (N_14383,N_14266,N_14353);
or U14384 (N_14384,N_14251,N_14270);
nand U14385 (N_14385,N_14336,N_14302);
or U14386 (N_14386,N_14280,N_14347);
and U14387 (N_14387,N_14346,N_14323);
nand U14388 (N_14388,N_14335,N_14363);
xor U14389 (N_14389,N_14366,N_14309);
or U14390 (N_14390,N_14296,N_14281);
nor U14391 (N_14391,N_14263,N_14274);
nand U14392 (N_14392,N_14345,N_14254);
nor U14393 (N_14393,N_14287,N_14359);
and U14394 (N_14394,N_14354,N_14292);
or U14395 (N_14395,N_14277,N_14315);
and U14396 (N_14396,N_14331,N_14340);
nand U14397 (N_14397,N_14332,N_14334);
nand U14398 (N_14398,N_14365,N_14278);
nand U14399 (N_14399,N_14283,N_14356);
xor U14400 (N_14400,N_14301,N_14322);
nor U14401 (N_14401,N_14294,N_14355);
and U14402 (N_14402,N_14314,N_14350);
and U14403 (N_14403,N_14261,N_14305);
and U14404 (N_14404,N_14275,N_14295);
nand U14405 (N_14405,N_14297,N_14316);
or U14406 (N_14406,N_14325,N_14358);
nand U14407 (N_14407,N_14298,N_14371);
nor U14408 (N_14408,N_14306,N_14267);
nor U14409 (N_14409,N_14373,N_14273);
or U14410 (N_14410,N_14364,N_14360);
or U14411 (N_14411,N_14310,N_14327);
or U14412 (N_14412,N_14328,N_14253);
and U14413 (N_14413,N_14341,N_14338);
nor U14414 (N_14414,N_14256,N_14361);
or U14415 (N_14415,N_14257,N_14362);
xnor U14416 (N_14416,N_14290,N_14324);
nor U14417 (N_14417,N_14259,N_14329);
xnor U14418 (N_14418,N_14285,N_14303);
xnor U14419 (N_14419,N_14372,N_14319);
xnor U14420 (N_14420,N_14252,N_14279);
and U14421 (N_14421,N_14271,N_14288);
xor U14422 (N_14422,N_14357,N_14313);
or U14423 (N_14423,N_14374,N_14333);
nand U14424 (N_14424,N_14368,N_14342);
nand U14425 (N_14425,N_14272,N_14262);
xor U14426 (N_14426,N_14307,N_14344);
or U14427 (N_14427,N_14299,N_14339);
and U14428 (N_14428,N_14300,N_14304);
xnor U14429 (N_14429,N_14337,N_14367);
nand U14430 (N_14430,N_14320,N_14326);
xor U14431 (N_14431,N_14311,N_14250);
or U14432 (N_14432,N_14291,N_14349);
nand U14433 (N_14433,N_14312,N_14264);
xnor U14434 (N_14434,N_14321,N_14289);
nand U14435 (N_14435,N_14293,N_14348);
xor U14436 (N_14436,N_14330,N_14308);
or U14437 (N_14437,N_14268,N_14329);
or U14438 (N_14438,N_14327,N_14292);
xor U14439 (N_14439,N_14369,N_14258);
nand U14440 (N_14440,N_14279,N_14308);
and U14441 (N_14441,N_14369,N_14279);
and U14442 (N_14442,N_14365,N_14326);
or U14443 (N_14443,N_14367,N_14267);
nor U14444 (N_14444,N_14358,N_14351);
or U14445 (N_14445,N_14279,N_14322);
nand U14446 (N_14446,N_14361,N_14319);
xnor U14447 (N_14447,N_14361,N_14314);
nand U14448 (N_14448,N_14251,N_14333);
xor U14449 (N_14449,N_14345,N_14291);
nand U14450 (N_14450,N_14275,N_14369);
and U14451 (N_14451,N_14304,N_14269);
or U14452 (N_14452,N_14274,N_14363);
xnor U14453 (N_14453,N_14358,N_14355);
or U14454 (N_14454,N_14330,N_14276);
and U14455 (N_14455,N_14263,N_14348);
and U14456 (N_14456,N_14290,N_14362);
nor U14457 (N_14457,N_14345,N_14371);
and U14458 (N_14458,N_14365,N_14349);
xnor U14459 (N_14459,N_14251,N_14358);
xor U14460 (N_14460,N_14277,N_14302);
nand U14461 (N_14461,N_14325,N_14341);
nor U14462 (N_14462,N_14287,N_14250);
xor U14463 (N_14463,N_14269,N_14355);
or U14464 (N_14464,N_14297,N_14274);
nand U14465 (N_14465,N_14309,N_14357);
or U14466 (N_14466,N_14278,N_14311);
and U14467 (N_14467,N_14287,N_14293);
nand U14468 (N_14468,N_14339,N_14357);
or U14469 (N_14469,N_14319,N_14362);
nor U14470 (N_14470,N_14340,N_14304);
xor U14471 (N_14471,N_14260,N_14335);
or U14472 (N_14472,N_14253,N_14339);
or U14473 (N_14473,N_14333,N_14295);
xor U14474 (N_14474,N_14337,N_14284);
xnor U14475 (N_14475,N_14359,N_14342);
xnor U14476 (N_14476,N_14304,N_14323);
or U14477 (N_14477,N_14275,N_14298);
nand U14478 (N_14478,N_14371,N_14297);
xnor U14479 (N_14479,N_14350,N_14261);
and U14480 (N_14480,N_14369,N_14370);
or U14481 (N_14481,N_14304,N_14369);
or U14482 (N_14482,N_14300,N_14331);
nand U14483 (N_14483,N_14330,N_14351);
nand U14484 (N_14484,N_14312,N_14355);
xnor U14485 (N_14485,N_14315,N_14346);
nand U14486 (N_14486,N_14355,N_14321);
and U14487 (N_14487,N_14267,N_14294);
nand U14488 (N_14488,N_14274,N_14275);
and U14489 (N_14489,N_14350,N_14366);
nor U14490 (N_14490,N_14305,N_14306);
nand U14491 (N_14491,N_14291,N_14256);
or U14492 (N_14492,N_14305,N_14370);
and U14493 (N_14493,N_14324,N_14352);
xor U14494 (N_14494,N_14312,N_14353);
or U14495 (N_14495,N_14360,N_14374);
or U14496 (N_14496,N_14271,N_14354);
nand U14497 (N_14497,N_14316,N_14329);
nor U14498 (N_14498,N_14355,N_14328);
or U14499 (N_14499,N_14293,N_14262);
and U14500 (N_14500,N_14460,N_14413);
and U14501 (N_14501,N_14399,N_14391);
or U14502 (N_14502,N_14436,N_14467);
nand U14503 (N_14503,N_14459,N_14455);
and U14504 (N_14504,N_14468,N_14435);
nand U14505 (N_14505,N_14397,N_14481);
xnor U14506 (N_14506,N_14480,N_14404);
nand U14507 (N_14507,N_14419,N_14433);
and U14508 (N_14508,N_14462,N_14389);
nor U14509 (N_14509,N_14422,N_14424);
and U14510 (N_14510,N_14484,N_14445);
nor U14511 (N_14511,N_14466,N_14492);
nand U14512 (N_14512,N_14438,N_14425);
nand U14513 (N_14513,N_14418,N_14412);
and U14514 (N_14514,N_14448,N_14390);
or U14515 (N_14515,N_14449,N_14488);
or U14516 (N_14516,N_14495,N_14405);
and U14517 (N_14517,N_14382,N_14375);
or U14518 (N_14518,N_14417,N_14434);
xnor U14519 (N_14519,N_14421,N_14446);
nand U14520 (N_14520,N_14470,N_14420);
xnor U14521 (N_14521,N_14496,N_14443);
or U14522 (N_14522,N_14478,N_14393);
and U14523 (N_14523,N_14472,N_14416);
or U14524 (N_14524,N_14498,N_14442);
nor U14525 (N_14525,N_14441,N_14396);
xor U14526 (N_14526,N_14447,N_14483);
xnor U14527 (N_14527,N_14471,N_14402);
and U14528 (N_14528,N_14497,N_14401);
and U14529 (N_14529,N_14426,N_14380);
or U14530 (N_14530,N_14384,N_14487);
and U14531 (N_14531,N_14394,N_14407);
and U14532 (N_14532,N_14437,N_14415);
nor U14533 (N_14533,N_14388,N_14482);
xnor U14534 (N_14534,N_14423,N_14489);
nand U14535 (N_14535,N_14414,N_14486);
nand U14536 (N_14536,N_14385,N_14476);
nor U14537 (N_14537,N_14464,N_14469);
xor U14538 (N_14538,N_14477,N_14461);
xor U14539 (N_14539,N_14458,N_14465);
or U14540 (N_14540,N_14453,N_14395);
nor U14541 (N_14541,N_14444,N_14411);
nand U14542 (N_14542,N_14432,N_14406);
and U14543 (N_14543,N_14451,N_14427);
nand U14544 (N_14544,N_14439,N_14463);
or U14545 (N_14545,N_14403,N_14378);
nor U14546 (N_14546,N_14392,N_14376);
or U14547 (N_14547,N_14377,N_14499);
nand U14548 (N_14548,N_14383,N_14440);
and U14549 (N_14549,N_14409,N_14457);
or U14550 (N_14550,N_14479,N_14473);
nand U14551 (N_14551,N_14410,N_14381);
nand U14552 (N_14552,N_14379,N_14386);
xor U14553 (N_14553,N_14456,N_14454);
and U14554 (N_14554,N_14490,N_14387);
or U14555 (N_14555,N_14475,N_14430);
or U14556 (N_14556,N_14474,N_14400);
xnor U14557 (N_14557,N_14431,N_14494);
or U14558 (N_14558,N_14452,N_14428);
nand U14559 (N_14559,N_14429,N_14398);
and U14560 (N_14560,N_14491,N_14450);
nor U14561 (N_14561,N_14485,N_14493);
or U14562 (N_14562,N_14408,N_14418);
or U14563 (N_14563,N_14468,N_14453);
or U14564 (N_14564,N_14443,N_14499);
nand U14565 (N_14565,N_14429,N_14422);
nor U14566 (N_14566,N_14441,N_14477);
and U14567 (N_14567,N_14462,N_14413);
nand U14568 (N_14568,N_14470,N_14404);
or U14569 (N_14569,N_14468,N_14482);
nand U14570 (N_14570,N_14413,N_14383);
xnor U14571 (N_14571,N_14488,N_14406);
or U14572 (N_14572,N_14438,N_14408);
nand U14573 (N_14573,N_14492,N_14499);
and U14574 (N_14574,N_14412,N_14465);
nand U14575 (N_14575,N_14489,N_14389);
or U14576 (N_14576,N_14400,N_14435);
nand U14577 (N_14577,N_14377,N_14458);
xor U14578 (N_14578,N_14459,N_14428);
and U14579 (N_14579,N_14397,N_14406);
nand U14580 (N_14580,N_14432,N_14437);
nand U14581 (N_14581,N_14445,N_14389);
nor U14582 (N_14582,N_14377,N_14375);
nor U14583 (N_14583,N_14379,N_14402);
nor U14584 (N_14584,N_14426,N_14457);
nand U14585 (N_14585,N_14461,N_14395);
or U14586 (N_14586,N_14376,N_14481);
nand U14587 (N_14587,N_14434,N_14377);
or U14588 (N_14588,N_14375,N_14434);
nor U14589 (N_14589,N_14449,N_14477);
and U14590 (N_14590,N_14490,N_14400);
and U14591 (N_14591,N_14413,N_14455);
or U14592 (N_14592,N_14421,N_14427);
and U14593 (N_14593,N_14461,N_14496);
and U14594 (N_14594,N_14428,N_14407);
nand U14595 (N_14595,N_14433,N_14386);
xnor U14596 (N_14596,N_14499,N_14410);
nor U14597 (N_14597,N_14379,N_14466);
xnor U14598 (N_14598,N_14385,N_14393);
nand U14599 (N_14599,N_14479,N_14418);
and U14600 (N_14600,N_14431,N_14490);
nand U14601 (N_14601,N_14468,N_14459);
or U14602 (N_14602,N_14375,N_14453);
nor U14603 (N_14603,N_14427,N_14411);
nand U14604 (N_14604,N_14466,N_14388);
nor U14605 (N_14605,N_14431,N_14378);
nand U14606 (N_14606,N_14450,N_14461);
or U14607 (N_14607,N_14404,N_14460);
nand U14608 (N_14608,N_14468,N_14478);
nor U14609 (N_14609,N_14466,N_14432);
and U14610 (N_14610,N_14436,N_14400);
nand U14611 (N_14611,N_14441,N_14390);
and U14612 (N_14612,N_14486,N_14467);
xnor U14613 (N_14613,N_14475,N_14401);
xnor U14614 (N_14614,N_14468,N_14432);
or U14615 (N_14615,N_14395,N_14423);
xor U14616 (N_14616,N_14460,N_14431);
nand U14617 (N_14617,N_14480,N_14398);
or U14618 (N_14618,N_14462,N_14477);
or U14619 (N_14619,N_14429,N_14431);
and U14620 (N_14620,N_14402,N_14414);
and U14621 (N_14621,N_14470,N_14432);
nand U14622 (N_14622,N_14396,N_14394);
and U14623 (N_14623,N_14410,N_14480);
nor U14624 (N_14624,N_14493,N_14437);
or U14625 (N_14625,N_14519,N_14583);
or U14626 (N_14626,N_14586,N_14502);
or U14627 (N_14627,N_14546,N_14600);
xnor U14628 (N_14628,N_14537,N_14524);
and U14629 (N_14629,N_14580,N_14515);
or U14630 (N_14630,N_14509,N_14530);
xnor U14631 (N_14631,N_14598,N_14545);
and U14632 (N_14632,N_14501,N_14541);
xnor U14633 (N_14633,N_14592,N_14581);
or U14634 (N_14634,N_14578,N_14516);
or U14635 (N_14635,N_14603,N_14565);
xnor U14636 (N_14636,N_14500,N_14594);
or U14637 (N_14637,N_14513,N_14508);
nand U14638 (N_14638,N_14596,N_14538);
xor U14639 (N_14639,N_14582,N_14607);
nor U14640 (N_14640,N_14557,N_14620);
nor U14641 (N_14641,N_14611,N_14564);
xor U14642 (N_14642,N_14561,N_14510);
nor U14643 (N_14643,N_14505,N_14601);
or U14644 (N_14644,N_14528,N_14593);
nor U14645 (N_14645,N_14577,N_14506);
and U14646 (N_14646,N_14597,N_14514);
xnor U14647 (N_14647,N_14532,N_14571);
nand U14648 (N_14648,N_14552,N_14518);
xnor U14649 (N_14649,N_14614,N_14605);
xor U14650 (N_14650,N_14588,N_14563);
nor U14651 (N_14651,N_14566,N_14599);
xor U14652 (N_14652,N_14619,N_14584);
and U14653 (N_14653,N_14573,N_14572);
nand U14654 (N_14654,N_14555,N_14504);
nor U14655 (N_14655,N_14560,N_14520);
xor U14656 (N_14656,N_14534,N_14525);
and U14657 (N_14657,N_14527,N_14604);
nand U14658 (N_14658,N_14547,N_14535);
and U14659 (N_14659,N_14543,N_14544);
or U14660 (N_14660,N_14602,N_14550);
or U14661 (N_14661,N_14562,N_14569);
nand U14662 (N_14662,N_14589,N_14531);
and U14663 (N_14663,N_14591,N_14533);
xor U14664 (N_14664,N_14553,N_14606);
or U14665 (N_14665,N_14612,N_14609);
or U14666 (N_14666,N_14556,N_14568);
nor U14667 (N_14667,N_14559,N_14529);
or U14668 (N_14668,N_14521,N_14549);
and U14669 (N_14669,N_14539,N_14503);
xor U14670 (N_14670,N_14507,N_14617);
xor U14671 (N_14671,N_14570,N_14608);
nand U14672 (N_14672,N_14623,N_14574);
nor U14673 (N_14673,N_14616,N_14613);
nand U14674 (N_14674,N_14558,N_14615);
and U14675 (N_14675,N_14575,N_14579);
nand U14676 (N_14676,N_14622,N_14554);
nor U14677 (N_14677,N_14523,N_14595);
and U14678 (N_14678,N_14548,N_14536);
and U14679 (N_14679,N_14587,N_14621);
or U14680 (N_14680,N_14522,N_14540);
nand U14681 (N_14681,N_14610,N_14551);
or U14682 (N_14682,N_14567,N_14512);
nor U14683 (N_14683,N_14576,N_14511);
nand U14684 (N_14684,N_14517,N_14542);
and U14685 (N_14685,N_14618,N_14624);
nand U14686 (N_14686,N_14526,N_14590);
or U14687 (N_14687,N_14585,N_14539);
or U14688 (N_14688,N_14581,N_14614);
nand U14689 (N_14689,N_14545,N_14601);
nand U14690 (N_14690,N_14521,N_14509);
nand U14691 (N_14691,N_14535,N_14609);
xnor U14692 (N_14692,N_14525,N_14594);
nor U14693 (N_14693,N_14598,N_14524);
xnor U14694 (N_14694,N_14580,N_14507);
xor U14695 (N_14695,N_14549,N_14562);
xor U14696 (N_14696,N_14614,N_14521);
xnor U14697 (N_14697,N_14617,N_14576);
nand U14698 (N_14698,N_14526,N_14605);
and U14699 (N_14699,N_14543,N_14553);
nor U14700 (N_14700,N_14534,N_14593);
nor U14701 (N_14701,N_14517,N_14569);
and U14702 (N_14702,N_14607,N_14509);
nor U14703 (N_14703,N_14540,N_14512);
nand U14704 (N_14704,N_14520,N_14543);
and U14705 (N_14705,N_14506,N_14547);
and U14706 (N_14706,N_14616,N_14500);
and U14707 (N_14707,N_14599,N_14535);
or U14708 (N_14708,N_14558,N_14623);
or U14709 (N_14709,N_14589,N_14547);
nor U14710 (N_14710,N_14570,N_14520);
nor U14711 (N_14711,N_14598,N_14530);
and U14712 (N_14712,N_14605,N_14510);
nand U14713 (N_14713,N_14582,N_14544);
and U14714 (N_14714,N_14612,N_14533);
or U14715 (N_14715,N_14607,N_14574);
xor U14716 (N_14716,N_14613,N_14590);
nor U14717 (N_14717,N_14501,N_14551);
nand U14718 (N_14718,N_14550,N_14593);
nor U14719 (N_14719,N_14585,N_14580);
and U14720 (N_14720,N_14618,N_14602);
xnor U14721 (N_14721,N_14595,N_14582);
nand U14722 (N_14722,N_14607,N_14624);
xor U14723 (N_14723,N_14537,N_14510);
or U14724 (N_14724,N_14558,N_14530);
nand U14725 (N_14725,N_14595,N_14610);
xor U14726 (N_14726,N_14555,N_14503);
nor U14727 (N_14727,N_14598,N_14513);
or U14728 (N_14728,N_14608,N_14574);
or U14729 (N_14729,N_14520,N_14541);
nand U14730 (N_14730,N_14620,N_14542);
nand U14731 (N_14731,N_14562,N_14583);
nor U14732 (N_14732,N_14505,N_14621);
xor U14733 (N_14733,N_14546,N_14581);
nand U14734 (N_14734,N_14612,N_14521);
and U14735 (N_14735,N_14604,N_14602);
xnor U14736 (N_14736,N_14608,N_14543);
nor U14737 (N_14737,N_14539,N_14544);
nor U14738 (N_14738,N_14595,N_14563);
or U14739 (N_14739,N_14608,N_14620);
nor U14740 (N_14740,N_14578,N_14520);
nand U14741 (N_14741,N_14581,N_14531);
xnor U14742 (N_14742,N_14591,N_14608);
nor U14743 (N_14743,N_14536,N_14535);
nor U14744 (N_14744,N_14612,N_14582);
nor U14745 (N_14745,N_14550,N_14546);
nor U14746 (N_14746,N_14565,N_14592);
nand U14747 (N_14747,N_14621,N_14618);
nand U14748 (N_14748,N_14534,N_14528);
and U14749 (N_14749,N_14533,N_14613);
xor U14750 (N_14750,N_14720,N_14683);
nand U14751 (N_14751,N_14687,N_14678);
nand U14752 (N_14752,N_14668,N_14728);
xnor U14753 (N_14753,N_14741,N_14730);
nor U14754 (N_14754,N_14738,N_14709);
nand U14755 (N_14755,N_14724,N_14639);
or U14756 (N_14756,N_14640,N_14712);
and U14757 (N_14757,N_14707,N_14731);
and U14758 (N_14758,N_14722,N_14705);
and U14759 (N_14759,N_14627,N_14658);
xor U14760 (N_14760,N_14636,N_14637);
xor U14761 (N_14761,N_14727,N_14682);
or U14762 (N_14762,N_14650,N_14746);
nand U14763 (N_14763,N_14744,N_14739);
xor U14764 (N_14764,N_14663,N_14659);
and U14765 (N_14765,N_14716,N_14725);
or U14766 (N_14766,N_14625,N_14657);
xor U14767 (N_14767,N_14713,N_14695);
xnor U14768 (N_14768,N_14647,N_14743);
nor U14769 (N_14769,N_14673,N_14643);
xor U14770 (N_14770,N_14737,N_14654);
or U14771 (N_14771,N_14645,N_14630);
nand U14772 (N_14772,N_14642,N_14680);
nand U14773 (N_14773,N_14688,N_14626);
and U14774 (N_14774,N_14653,N_14651);
and U14775 (N_14775,N_14661,N_14646);
nand U14776 (N_14776,N_14676,N_14635);
or U14777 (N_14777,N_14671,N_14702);
nand U14778 (N_14778,N_14748,N_14628);
nor U14779 (N_14779,N_14719,N_14641);
and U14780 (N_14780,N_14706,N_14694);
xnor U14781 (N_14781,N_14669,N_14740);
and U14782 (N_14782,N_14670,N_14633);
nand U14783 (N_14783,N_14699,N_14689);
or U14784 (N_14784,N_14736,N_14649);
or U14785 (N_14785,N_14708,N_14697);
nand U14786 (N_14786,N_14747,N_14717);
nor U14787 (N_14787,N_14703,N_14652);
or U14788 (N_14788,N_14693,N_14692);
nand U14789 (N_14789,N_14674,N_14648);
and U14790 (N_14790,N_14742,N_14729);
nand U14791 (N_14791,N_14685,N_14691);
or U14792 (N_14792,N_14665,N_14632);
nor U14793 (N_14793,N_14672,N_14660);
or U14794 (N_14794,N_14745,N_14700);
xnor U14795 (N_14795,N_14634,N_14734);
xnor U14796 (N_14796,N_14644,N_14662);
or U14797 (N_14797,N_14733,N_14629);
and U14798 (N_14798,N_14690,N_14749);
xnor U14799 (N_14799,N_14698,N_14655);
nand U14800 (N_14800,N_14667,N_14677);
nand U14801 (N_14801,N_14711,N_14735);
xnor U14802 (N_14802,N_14723,N_14681);
nor U14803 (N_14803,N_14679,N_14638);
and U14804 (N_14804,N_14675,N_14656);
and U14805 (N_14805,N_14721,N_14696);
nor U14806 (N_14806,N_14686,N_14710);
or U14807 (N_14807,N_14732,N_14701);
xnor U14808 (N_14808,N_14714,N_14726);
nor U14809 (N_14809,N_14631,N_14664);
and U14810 (N_14810,N_14666,N_14704);
xnor U14811 (N_14811,N_14718,N_14715);
nor U14812 (N_14812,N_14684,N_14655);
and U14813 (N_14813,N_14681,N_14722);
and U14814 (N_14814,N_14715,N_14675);
nand U14815 (N_14815,N_14637,N_14668);
and U14816 (N_14816,N_14682,N_14722);
nand U14817 (N_14817,N_14627,N_14747);
and U14818 (N_14818,N_14723,N_14729);
nor U14819 (N_14819,N_14666,N_14691);
xnor U14820 (N_14820,N_14740,N_14639);
or U14821 (N_14821,N_14682,N_14638);
xor U14822 (N_14822,N_14699,N_14647);
xnor U14823 (N_14823,N_14721,N_14724);
nor U14824 (N_14824,N_14662,N_14697);
xnor U14825 (N_14825,N_14685,N_14719);
and U14826 (N_14826,N_14747,N_14700);
nor U14827 (N_14827,N_14733,N_14680);
or U14828 (N_14828,N_14671,N_14734);
or U14829 (N_14829,N_14681,N_14633);
or U14830 (N_14830,N_14627,N_14694);
nor U14831 (N_14831,N_14632,N_14741);
or U14832 (N_14832,N_14744,N_14663);
nor U14833 (N_14833,N_14693,N_14626);
nor U14834 (N_14834,N_14682,N_14695);
nor U14835 (N_14835,N_14706,N_14683);
nor U14836 (N_14836,N_14694,N_14747);
nand U14837 (N_14837,N_14737,N_14648);
nor U14838 (N_14838,N_14631,N_14713);
xor U14839 (N_14839,N_14645,N_14672);
and U14840 (N_14840,N_14693,N_14644);
and U14841 (N_14841,N_14630,N_14705);
or U14842 (N_14842,N_14667,N_14681);
or U14843 (N_14843,N_14654,N_14694);
and U14844 (N_14844,N_14675,N_14699);
and U14845 (N_14845,N_14678,N_14671);
and U14846 (N_14846,N_14648,N_14706);
xor U14847 (N_14847,N_14713,N_14643);
or U14848 (N_14848,N_14637,N_14681);
xnor U14849 (N_14849,N_14636,N_14704);
nor U14850 (N_14850,N_14634,N_14720);
nor U14851 (N_14851,N_14737,N_14630);
and U14852 (N_14852,N_14626,N_14674);
nand U14853 (N_14853,N_14730,N_14714);
xor U14854 (N_14854,N_14700,N_14634);
and U14855 (N_14855,N_14730,N_14691);
or U14856 (N_14856,N_14722,N_14664);
nand U14857 (N_14857,N_14633,N_14647);
nor U14858 (N_14858,N_14709,N_14686);
nor U14859 (N_14859,N_14698,N_14654);
and U14860 (N_14860,N_14636,N_14709);
or U14861 (N_14861,N_14726,N_14736);
or U14862 (N_14862,N_14644,N_14684);
nand U14863 (N_14863,N_14648,N_14693);
or U14864 (N_14864,N_14699,N_14731);
or U14865 (N_14865,N_14668,N_14686);
xnor U14866 (N_14866,N_14683,N_14679);
or U14867 (N_14867,N_14716,N_14649);
and U14868 (N_14868,N_14712,N_14708);
and U14869 (N_14869,N_14725,N_14703);
or U14870 (N_14870,N_14654,N_14682);
nand U14871 (N_14871,N_14704,N_14685);
nand U14872 (N_14872,N_14743,N_14711);
xor U14873 (N_14873,N_14676,N_14694);
xor U14874 (N_14874,N_14625,N_14659);
xnor U14875 (N_14875,N_14753,N_14785);
nor U14876 (N_14876,N_14850,N_14774);
or U14877 (N_14877,N_14846,N_14752);
nand U14878 (N_14878,N_14855,N_14760);
nor U14879 (N_14879,N_14809,N_14873);
or U14880 (N_14880,N_14867,N_14853);
nand U14881 (N_14881,N_14811,N_14847);
nor U14882 (N_14882,N_14839,N_14860);
and U14883 (N_14883,N_14821,N_14815);
nand U14884 (N_14884,N_14824,N_14805);
and U14885 (N_14885,N_14865,N_14828);
xnor U14886 (N_14886,N_14807,N_14827);
nand U14887 (N_14887,N_14831,N_14848);
or U14888 (N_14888,N_14755,N_14808);
and U14889 (N_14889,N_14854,N_14750);
and U14890 (N_14890,N_14864,N_14758);
nor U14891 (N_14891,N_14757,N_14789);
nor U14892 (N_14892,N_14803,N_14840);
xnor U14893 (N_14893,N_14790,N_14842);
or U14894 (N_14894,N_14862,N_14826);
nand U14895 (N_14895,N_14813,N_14830);
or U14896 (N_14896,N_14858,N_14779);
and U14897 (N_14897,N_14765,N_14849);
or U14898 (N_14898,N_14817,N_14861);
nor U14899 (N_14899,N_14791,N_14777);
or U14900 (N_14900,N_14795,N_14764);
or U14901 (N_14901,N_14823,N_14773);
or U14902 (N_14902,N_14759,N_14783);
nand U14903 (N_14903,N_14812,N_14868);
nand U14904 (N_14904,N_14851,N_14814);
xnor U14905 (N_14905,N_14781,N_14838);
nor U14906 (N_14906,N_14775,N_14804);
xnor U14907 (N_14907,N_14754,N_14784);
or U14908 (N_14908,N_14786,N_14810);
xnor U14909 (N_14909,N_14798,N_14834);
and U14910 (N_14910,N_14778,N_14761);
nor U14911 (N_14911,N_14822,N_14780);
xnor U14912 (N_14912,N_14806,N_14866);
nand U14913 (N_14913,N_14871,N_14872);
nand U14914 (N_14914,N_14802,N_14857);
and U14915 (N_14915,N_14816,N_14841);
nand U14916 (N_14916,N_14776,N_14819);
xor U14917 (N_14917,N_14829,N_14856);
nor U14918 (N_14918,N_14762,N_14756);
and U14919 (N_14919,N_14852,N_14782);
xor U14920 (N_14920,N_14766,N_14833);
or U14921 (N_14921,N_14836,N_14793);
and U14922 (N_14922,N_14859,N_14800);
xor U14923 (N_14923,N_14787,N_14771);
xor U14924 (N_14924,N_14751,N_14788);
xnor U14925 (N_14925,N_14845,N_14843);
xor U14926 (N_14926,N_14844,N_14763);
and U14927 (N_14927,N_14797,N_14870);
or U14928 (N_14928,N_14799,N_14818);
xor U14929 (N_14929,N_14767,N_14869);
and U14930 (N_14930,N_14874,N_14792);
and U14931 (N_14931,N_14863,N_14796);
or U14932 (N_14932,N_14794,N_14772);
or U14933 (N_14933,N_14835,N_14832);
nand U14934 (N_14934,N_14769,N_14801);
nor U14935 (N_14935,N_14820,N_14837);
or U14936 (N_14936,N_14825,N_14768);
or U14937 (N_14937,N_14770,N_14812);
or U14938 (N_14938,N_14816,N_14796);
nand U14939 (N_14939,N_14756,N_14840);
nor U14940 (N_14940,N_14783,N_14869);
and U14941 (N_14941,N_14800,N_14860);
and U14942 (N_14942,N_14864,N_14819);
nor U14943 (N_14943,N_14825,N_14797);
nand U14944 (N_14944,N_14752,N_14851);
and U14945 (N_14945,N_14855,N_14823);
xnor U14946 (N_14946,N_14825,N_14764);
nand U14947 (N_14947,N_14792,N_14775);
nor U14948 (N_14948,N_14781,N_14862);
or U14949 (N_14949,N_14752,N_14870);
xnor U14950 (N_14950,N_14801,N_14833);
xor U14951 (N_14951,N_14864,N_14855);
and U14952 (N_14952,N_14852,N_14830);
nand U14953 (N_14953,N_14797,N_14769);
xor U14954 (N_14954,N_14779,N_14834);
and U14955 (N_14955,N_14863,N_14788);
nand U14956 (N_14956,N_14794,N_14797);
xor U14957 (N_14957,N_14792,N_14837);
nand U14958 (N_14958,N_14826,N_14800);
and U14959 (N_14959,N_14859,N_14865);
and U14960 (N_14960,N_14870,N_14750);
or U14961 (N_14961,N_14787,N_14858);
nor U14962 (N_14962,N_14759,N_14859);
and U14963 (N_14963,N_14857,N_14791);
nand U14964 (N_14964,N_14828,N_14786);
xnor U14965 (N_14965,N_14779,N_14773);
nand U14966 (N_14966,N_14852,N_14828);
and U14967 (N_14967,N_14834,N_14750);
xor U14968 (N_14968,N_14838,N_14866);
xor U14969 (N_14969,N_14847,N_14763);
nor U14970 (N_14970,N_14790,N_14776);
nand U14971 (N_14971,N_14853,N_14787);
nor U14972 (N_14972,N_14860,N_14759);
nor U14973 (N_14973,N_14788,N_14804);
xnor U14974 (N_14974,N_14801,N_14830);
or U14975 (N_14975,N_14759,N_14784);
xnor U14976 (N_14976,N_14812,N_14864);
nand U14977 (N_14977,N_14820,N_14846);
xor U14978 (N_14978,N_14800,N_14816);
and U14979 (N_14979,N_14865,N_14852);
or U14980 (N_14980,N_14817,N_14862);
xnor U14981 (N_14981,N_14758,N_14815);
nand U14982 (N_14982,N_14866,N_14750);
nor U14983 (N_14983,N_14859,N_14760);
and U14984 (N_14984,N_14859,N_14822);
and U14985 (N_14985,N_14818,N_14785);
xnor U14986 (N_14986,N_14821,N_14824);
nand U14987 (N_14987,N_14859,N_14798);
nand U14988 (N_14988,N_14771,N_14758);
nand U14989 (N_14989,N_14750,N_14846);
nor U14990 (N_14990,N_14824,N_14791);
and U14991 (N_14991,N_14874,N_14768);
or U14992 (N_14992,N_14841,N_14829);
nand U14993 (N_14993,N_14789,N_14867);
xnor U14994 (N_14994,N_14791,N_14870);
xor U14995 (N_14995,N_14828,N_14757);
and U14996 (N_14996,N_14853,N_14862);
nor U14997 (N_14997,N_14792,N_14867);
nor U14998 (N_14998,N_14757,N_14770);
nand U14999 (N_14999,N_14845,N_14823);
nor UO_0 (O_0,N_14896,N_14986);
nand UO_1 (O_1,N_14977,N_14897);
nor UO_2 (O_2,N_14902,N_14997);
nand UO_3 (O_3,N_14990,N_14877);
nand UO_4 (O_4,N_14968,N_14899);
nor UO_5 (O_5,N_14921,N_14912);
nor UO_6 (O_6,N_14885,N_14953);
xnor UO_7 (O_7,N_14945,N_14911);
nor UO_8 (O_8,N_14969,N_14925);
and UO_9 (O_9,N_14995,N_14973);
nand UO_10 (O_10,N_14949,N_14930);
nor UO_11 (O_11,N_14891,N_14958);
or UO_12 (O_12,N_14914,N_14935);
nor UO_13 (O_13,N_14999,N_14898);
nor UO_14 (O_14,N_14884,N_14892);
and UO_15 (O_15,N_14940,N_14964);
and UO_16 (O_16,N_14882,N_14886);
or UO_17 (O_17,N_14889,N_14883);
nand UO_18 (O_18,N_14970,N_14926);
and UO_19 (O_19,N_14957,N_14992);
xnor UO_20 (O_20,N_14907,N_14916);
xor UO_21 (O_21,N_14934,N_14900);
nor UO_22 (O_22,N_14947,N_14939);
nand UO_23 (O_23,N_14888,N_14895);
nand UO_24 (O_24,N_14981,N_14928);
and UO_25 (O_25,N_14963,N_14943);
xnor UO_26 (O_26,N_14965,N_14946);
nand UO_27 (O_27,N_14959,N_14980);
and UO_28 (O_28,N_14944,N_14987);
and UO_29 (O_29,N_14910,N_14982);
xor UO_30 (O_30,N_14908,N_14954);
or UO_31 (O_31,N_14893,N_14971);
nor UO_32 (O_32,N_14881,N_14972);
xor UO_33 (O_33,N_14978,N_14966);
nand UO_34 (O_34,N_14938,N_14894);
xor UO_35 (O_35,N_14936,N_14956);
nand UO_36 (O_36,N_14950,N_14979);
and UO_37 (O_37,N_14876,N_14920);
xor UO_38 (O_38,N_14922,N_14983);
xnor UO_39 (O_39,N_14994,N_14890);
nor UO_40 (O_40,N_14932,N_14941);
and UO_41 (O_41,N_14975,N_14923);
nor UO_42 (O_42,N_14924,N_14976);
and UO_43 (O_43,N_14974,N_14905);
nand UO_44 (O_44,N_14903,N_14984);
nand UO_45 (O_45,N_14960,N_14880);
and UO_46 (O_46,N_14933,N_14967);
nand UO_47 (O_47,N_14988,N_14875);
or UO_48 (O_48,N_14909,N_14961);
or UO_49 (O_49,N_14942,N_14879);
xnor UO_50 (O_50,N_14985,N_14998);
and UO_51 (O_51,N_14931,N_14906);
xor UO_52 (O_52,N_14927,N_14993);
and UO_53 (O_53,N_14929,N_14989);
or UO_54 (O_54,N_14878,N_14991);
xnor UO_55 (O_55,N_14913,N_14948);
or UO_56 (O_56,N_14901,N_14951);
and UO_57 (O_57,N_14962,N_14937);
xnor UO_58 (O_58,N_14915,N_14952);
nand UO_59 (O_59,N_14904,N_14919);
nand UO_60 (O_60,N_14955,N_14996);
xnor UO_61 (O_61,N_14917,N_14887);
nand UO_62 (O_62,N_14918,N_14965);
xnor UO_63 (O_63,N_14896,N_14949);
nand UO_64 (O_64,N_14898,N_14915);
nor UO_65 (O_65,N_14913,N_14950);
or UO_66 (O_66,N_14991,N_14905);
nand UO_67 (O_67,N_14956,N_14896);
and UO_68 (O_68,N_14923,N_14911);
and UO_69 (O_69,N_14970,N_14937);
and UO_70 (O_70,N_14971,N_14980);
and UO_71 (O_71,N_14989,N_14878);
xnor UO_72 (O_72,N_14911,N_14982);
nor UO_73 (O_73,N_14926,N_14907);
and UO_74 (O_74,N_14909,N_14905);
or UO_75 (O_75,N_14991,N_14990);
nand UO_76 (O_76,N_14946,N_14974);
xnor UO_77 (O_77,N_14993,N_14942);
xnor UO_78 (O_78,N_14941,N_14973);
nor UO_79 (O_79,N_14993,N_14970);
nor UO_80 (O_80,N_14894,N_14945);
xor UO_81 (O_81,N_14964,N_14895);
xor UO_82 (O_82,N_14889,N_14938);
nand UO_83 (O_83,N_14877,N_14952);
nand UO_84 (O_84,N_14949,N_14941);
and UO_85 (O_85,N_14934,N_14954);
and UO_86 (O_86,N_14932,N_14933);
and UO_87 (O_87,N_14899,N_14988);
or UO_88 (O_88,N_14991,N_14969);
nand UO_89 (O_89,N_14880,N_14950);
nor UO_90 (O_90,N_14981,N_14945);
or UO_91 (O_91,N_14955,N_14900);
or UO_92 (O_92,N_14964,N_14928);
nand UO_93 (O_93,N_14978,N_14947);
or UO_94 (O_94,N_14951,N_14998);
or UO_95 (O_95,N_14960,N_14908);
xor UO_96 (O_96,N_14997,N_14986);
xnor UO_97 (O_97,N_14974,N_14880);
and UO_98 (O_98,N_14891,N_14981);
nor UO_99 (O_99,N_14887,N_14894);
nand UO_100 (O_100,N_14895,N_14940);
xor UO_101 (O_101,N_14988,N_14922);
nor UO_102 (O_102,N_14951,N_14914);
or UO_103 (O_103,N_14999,N_14994);
or UO_104 (O_104,N_14978,N_14934);
nor UO_105 (O_105,N_14916,N_14933);
and UO_106 (O_106,N_14975,N_14967);
or UO_107 (O_107,N_14913,N_14979);
nor UO_108 (O_108,N_14904,N_14982);
xnor UO_109 (O_109,N_14944,N_14977);
nand UO_110 (O_110,N_14963,N_14884);
and UO_111 (O_111,N_14883,N_14936);
xnor UO_112 (O_112,N_14980,N_14923);
nor UO_113 (O_113,N_14988,N_14960);
or UO_114 (O_114,N_14944,N_14971);
nand UO_115 (O_115,N_14876,N_14944);
xor UO_116 (O_116,N_14989,N_14882);
xnor UO_117 (O_117,N_14914,N_14969);
and UO_118 (O_118,N_14969,N_14999);
and UO_119 (O_119,N_14899,N_14911);
or UO_120 (O_120,N_14920,N_14917);
nand UO_121 (O_121,N_14980,N_14990);
nand UO_122 (O_122,N_14936,N_14968);
nand UO_123 (O_123,N_14879,N_14882);
nor UO_124 (O_124,N_14977,N_14965);
or UO_125 (O_125,N_14907,N_14921);
nand UO_126 (O_126,N_14893,N_14900);
nand UO_127 (O_127,N_14921,N_14995);
nand UO_128 (O_128,N_14891,N_14920);
xnor UO_129 (O_129,N_14933,N_14936);
xor UO_130 (O_130,N_14905,N_14878);
and UO_131 (O_131,N_14878,N_14914);
or UO_132 (O_132,N_14986,N_14974);
and UO_133 (O_133,N_14954,N_14893);
or UO_134 (O_134,N_14973,N_14885);
or UO_135 (O_135,N_14940,N_14957);
or UO_136 (O_136,N_14918,N_14943);
and UO_137 (O_137,N_14954,N_14922);
nand UO_138 (O_138,N_14998,N_14989);
nand UO_139 (O_139,N_14941,N_14915);
and UO_140 (O_140,N_14934,N_14979);
nor UO_141 (O_141,N_14982,N_14966);
nor UO_142 (O_142,N_14912,N_14881);
or UO_143 (O_143,N_14941,N_14892);
nor UO_144 (O_144,N_14983,N_14935);
xnor UO_145 (O_145,N_14963,N_14888);
nor UO_146 (O_146,N_14900,N_14892);
and UO_147 (O_147,N_14902,N_14964);
nand UO_148 (O_148,N_14878,N_14923);
nor UO_149 (O_149,N_14927,N_14945);
and UO_150 (O_150,N_14897,N_14972);
nor UO_151 (O_151,N_14908,N_14922);
and UO_152 (O_152,N_14946,N_14970);
nor UO_153 (O_153,N_14898,N_14951);
or UO_154 (O_154,N_14896,N_14944);
or UO_155 (O_155,N_14876,N_14881);
or UO_156 (O_156,N_14980,N_14927);
and UO_157 (O_157,N_14948,N_14927);
nor UO_158 (O_158,N_14977,N_14884);
nand UO_159 (O_159,N_14903,N_14978);
nand UO_160 (O_160,N_14909,N_14906);
nor UO_161 (O_161,N_14998,N_14886);
and UO_162 (O_162,N_14890,N_14912);
nand UO_163 (O_163,N_14959,N_14903);
nor UO_164 (O_164,N_14898,N_14997);
nor UO_165 (O_165,N_14890,N_14949);
and UO_166 (O_166,N_14939,N_14934);
or UO_167 (O_167,N_14910,N_14939);
nor UO_168 (O_168,N_14978,N_14884);
xnor UO_169 (O_169,N_14896,N_14965);
nor UO_170 (O_170,N_14957,N_14984);
nor UO_171 (O_171,N_14877,N_14907);
and UO_172 (O_172,N_14920,N_14956);
nand UO_173 (O_173,N_14944,N_14892);
nand UO_174 (O_174,N_14986,N_14969);
nor UO_175 (O_175,N_14986,N_14982);
nor UO_176 (O_176,N_14919,N_14931);
nand UO_177 (O_177,N_14948,N_14963);
nor UO_178 (O_178,N_14882,N_14898);
and UO_179 (O_179,N_14909,N_14967);
xnor UO_180 (O_180,N_14987,N_14952);
nand UO_181 (O_181,N_14900,N_14901);
nand UO_182 (O_182,N_14982,N_14993);
and UO_183 (O_183,N_14930,N_14978);
xor UO_184 (O_184,N_14923,N_14984);
or UO_185 (O_185,N_14876,N_14979);
and UO_186 (O_186,N_14922,N_14978);
nand UO_187 (O_187,N_14929,N_14912);
xor UO_188 (O_188,N_14973,N_14897);
nor UO_189 (O_189,N_14959,N_14875);
and UO_190 (O_190,N_14921,N_14887);
or UO_191 (O_191,N_14982,N_14937);
and UO_192 (O_192,N_14990,N_14982);
nand UO_193 (O_193,N_14961,N_14884);
and UO_194 (O_194,N_14993,N_14886);
or UO_195 (O_195,N_14906,N_14998);
or UO_196 (O_196,N_14957,N_14935);
nor UO_197 (O_197,N_14982,N_14932);
nor UO_198 (O_198,N_14886,N_14999);
or UO_199 (O_199,N_14976,N_14932);
xor UO_200 (O_200,N_14913,N_14995);
or UO_201 (O_201,N_14949,N_14968);
and UO_202 (O_202,N_14930,N_14907);
or UO_203 (O_203,N_14922,N_14898);
nand UO_204 (O_204,N_14998,N_14897);
or UO_205 (O_205,N_14980,N_14943);
or UO_206 (O_206,N_14920,N_14888);
nand UO_207 (O_207,N_14908,N_14958);
xor UO_208 (O_208,N_14946,N_14880);
xor UO_209 (O_209,N_14902,N_14993);
or UO_210 (O_210,N_14884,N_14986);
nor UO_211 (O_211,N_14994,N_14949);
nand UO_212 (O_212,N_14977,N_14983);
or UO_213 (O_213,N_14995,N_14992);
nor UO_214 (O_214,N_14921,N_14914);
xnor UO_215 (O_215,N_14899,N_14980);
nor UO_216 (O_216,N_14978,N_14977);
and UO_217 (O_217,N_14908,N_14929);
and UO_218 (O_218,N_14991,N_14983);
nand UO_219 (O_219,N_14995,N_14966);
or UO_220 (O_220,N_14949,N_14931);
nand UO_221 (O_221,N_14942,N_14933);
and UO_222 (O_222,N_14943,N_14986);
xnor UO_223 (O_223,N_14958,N_14942);
and UO_224 (O_224,N_14893,N_14943);
and UO_225 (O_225,N_14915,N_14935);
or UO_226 (O_226,N_14999,N_14992);
and UO_227 (O_227,N_14966,N_14967);
nor UO_228 (O_228,N_14921,N_14952);
nor UO_229 (O_229,N_14913,N_14882);
and UO_230 (O_230,N_14897,N_14904);
nand UO_231 (O_231,N_14883,N_14941);
xnor UO_232 (O_232,N_14995,N_14901);
nor UO_233 (O_233,N_14987,N_14983);
xor UO_234 (O_234,N_14927,N_14917);
nor UO_235 (O_235,N_14971,N_14890);
and UO_236 (O_236,N_14892,N_14982);
nor UO_237 (O_237,N_14954,N_14942);
nand UO_238 (O_238,N_14984,N_14941);
or UO_239 (O_239,N_14931,N_14916);
nand UO_240 (O_240,N_14906,N_14963);
nor UO_241 (O_241,N_14953,N_14908);
nor UO_242 (O_242,N_14942,N_14880);
nand UO_243 (O_243,N_14875,N_14891);
or UO_244 (O_244,N_14945,N_14999);
xor UO_245 (O_245,N_14992,N_14967);
and UO_246 (O_246,N_14897,N_14935);
nand UO_247 (O_247,N_14938,N_14901);
nor UO_248 (O_248,N_14917,N_14895);
nand UO_249 (O_249,N_14917,N_14969);
nand UO_250 (O_250,N_14990,N_14938);
nand UO_251 (O_251,N_14893,N_14914);
and UO_252 (O_252,N_14961,N_14916);
xor UO_253 (O_253,N_14924,N_14902);
and UO_254 (O_254,N_14933,N_14941);
xnor UO_255 (O_255,N_14904,N_14902);
nor UO_256 (O_256,N_14956,N_14915);
nand UO_257 (O_257,N_14905,N_14990);
and UO_258 (O_258,N_14940,N_14970);
nand UO_259 (O_259,N_14982,N_14967);
or UO_260 (O_260,N_14981,N_14967);
xnor UO_261 (O_261,N_14942,N_14940);
and UO_262 (O_262,N_14973,N_14937);
and UO_263 (O_263,N_14931,N_14988);
or UO_264 (O_264,N_14905,N_14917);
and UO_265 (O_265,N_14955,N_14991);
nand UO_266 (O_266,N_14977,N_14971);
and UO_267 (O_267,N_14904,N_14907);
xor UO_268 (O_268,N_14944,N_14980);
and UO_269 (O_269,N_14975,N_14958);
nand UO_270 (O_270,N_14967,N_14884);
nand UO_271 (O_271,N_14995,N_14969);
nand UO_272 (O_272,N_14898,N_14878);
nand UO_273 (O_273,N_14968,N_14886);
nor UO_274 (O_274,N_14892,N_14936);
or UO_275 (O_275,N_14935,N_14958);
xor UO_276 (O_276,N_14940,N_14982);
xnor UO_277 (O_277,N_14949,N_14976);
and UO_278 (O_278,N_14939,N_14952);
nor UO_279 (O_279,N_14880,N_14917);
xnor UO_280 (O_280,N_14962,N_14986);
or UO_281 (O_281,N_14896,N_14991);
and UO_282 (O_282,N_14948,N_14943);
xnor UO_283 (O_283,N_14911,N_14974);
xnor UO_284 (O_284,N_14902,N_14990);
nor UO_285 (O_285,N_14915,N_14978);
nand UO_286 (O_286,N_14876,N_14898);
or UO_287 (O_287,N_14989,N_14894);
xnor UO_288 (O_288,N_14890,N_14916);
or UO_289 (O_289,N_14944,N_14959);
nor UO_290 (O_290,N_14996,N_14875);
xnor UO_291 (O_291,N_14978,N_14982);
xor UO_292 (O_292,N_14928,N_14963);
xor UO_293 (O_293,N_14916,N_14894);
and UO_294 (O_294,N_14936,N_14993);
nand UO_295 (O_295,N_14908,N_14977);
nand UO_296 (O_296,N_14922,N_14963);
and UO_297 (O_297,N_14937,N_14898);
nand UO_298 (O_298,N_14915,N_14965);
xor UO_299 (O_299,N_14986,N_14893);
and UO_300 (O_300,N_14975,N_14902);
and UO_301 (O_301,N_14940,N_14892);
or UO_302 (O_302,N_14883,N_14960);
nand UO_303 (O_303,N_14986,N_14882);
and UO_304 (O_304,N_14885,N_14962);
or UO_305 (O_305,N_14897,N_14932);
and UO_306 (O_306,N_14962,N_14966);
nor UO_307 (O_307,N_14986,N_14990);
xor UO_308 (O_308,N_14976,N_14894);
nand UO_309 (O_309,N_14991,N_14916);
nor UO_310 (O_310,N_14924,N_14943);
and UO_311 (O_311,N_14934,N_14881);
nor UO_312 (O_312,N_14925,N_14946);
nand UO_313 (O_313,N_14976,N_14887);
or UO_314 (O_314,N_14935,N_14996);
or UO_315 (O_315,N_14888,N_14944);
xnor UO_316 (O_316,N_14972,N_14956);
or UO_317 (O_317,N_14992,N_14942);
nor UO_318 (O_318,N_14993,N_14968);
xnor UO_319 (O_319,N_14884,N_14911);
nor UO_320 (O_320,N_14888,N_14896);
or UO_321 (O_321,N_14990,N_14939);
xnor UO_322 (O_322,N_14979,N_14900);
nand UO_323 (O_323,N_14990,N_14951);
or UO_324 (O_324,N_14875,N_14909);
or UO_325 (O_325,N_14968,N_14894);
or UO_326 (O_326,N_14911,N_14877);
nor UO_327 (O_327,N_14932,N_14895);
or UO_328 (O_328,N_14995,N_14965);
and UO_329 (O_329,N_14967,N_14923);
nor UO_330 (O_330,N_14892,N_14999);
or UO_331 (O_331,N_14989,N_14906);
or UO_332 (O_332,N_14893,N_14918);
nor UO_333 (O_333,N_14909,N_14921);
nor UO_334 (O_334,N_14917,N_14942);
nor UO_335 (O_335,N_14915,N_14928);
nor UO_336 (O_336,N_14987,N_14949);
or UO_337 (O_337,N_14967,N_14892);
nand UO_338 (O_338,N_14893,N_14926);
or UO_339 (O_339,N_14930,N_14996);
nor UO_340 (O_340,N_14922,N_14936);
xor UO_341 (O_341,N_14961,N_14997);
and UO_342 (O_342,N_14995,N_14960);
xor UO_343 (O_343,N_14910,N_14965);
and UO_344 (O_344,N_14906,N_14929);
nand UO_345 (O_345,N_14891,N_14971);
nand UO_346 (O_346,N_14949,N_14993);
nor UO_347 (O_347,N_14890,N_14926);
or UO_348 (O_348,N_14879,N_14941);
xor UO_349 (O_349,N_14921,N_14881);
and UO_350 (O_350,N_14935,N_14948);
and UO_351 (O_351,N_14928,N_14906);
nand UO_352 (O_352,N_14977,N_14998);
xor UO_353 (O_353,N_14932,N_14965);
and UO_354 (O_354,N_14911,N_14952);
or UO_355 (O_355,N_14879,N_14897);
nand UO_356 (O_356,N_14877,N_14942);
nor UO_357 (O_357,N_14893,N_14888);
and UO_358 (O_358,N_14875,N_14961);
xnor UO_359 (O_359,N_14878,N_14907);
xnor UO_360 (O_360,N_14902,N_14889);
nor UO_361 (O_361,N_14937,N_14916);
nor UO_362 (O_362,N_14975,N_14899);
nor UO_363 (O_363,N_14960,N_14985);
xnor UO_364 (O_364,N_14879,N_14990);
or UO_365 (O_365,N_14938,N_14977);
or UO_366 (O_366,N_14996,N_14897);
and UO_367 (O_367,N_14900,N_14913);
and UO_368 (O_368,N_14877,N_14972);
xnor UO_369 (O_369,N_14937,N_14977);
nor UO_370 (O_370,N_14896,N_14904);
xor UO_371 (O_371,N_14916,N_14984);
and UO_372 (O_372,N_14957,N_14989);
nor UO_373 (O_373,N_14945,N_14920);
and UO_374 (O_374,N_14978,N_14909);
nor UO_375 (O_375,N_14986,N_14930);
nand UO_376 (O_376,N_14894,N_14913);
xor UO_377 (O_377,N_14914,N_14994);
or UO_378 (O_378,N_14882,N_14877);
or UO_379 (O_379,N_14924,N_14950);
xor UO_380 (O_380,N_14923,N_14882);
and UO_381 (O_381,N_14901,N_14981);
xor UO_382 (O_382,N_14927,N_14918);
and UO_383 (O_383,N_14974,N_14998);
nand UO_384 (O_384,N_14879,N_14936);
or UO_385 (O_385,N_14944,N_14941);
nand UO_386 (O_386,N_14960,N_14936);
and UO_387 (O_387,N_14891,N_14888);
nand UO_388 (O_388,N_14953,N_14879);
xor UO_389 (O_389,N_14909,N_14997);
nor UO_390 (O_390,N_14988,N_14896);
and UO_391 (O_391,N_14960,N_14932);
and UO_392 (O_392,N_14964,N_14957);
and UO_393 (O_393,N_14924,N_14954);
or UO_394 (O_394,N_14904,N_14885);
nor UO_395 (O_395,N_14910,N_14962);
nor UO_396 (O_396,N_14946,N_14895);
xnor UO_397 (O_397,N_14937,N_14950);
nand UO_398 (O_398,N_14941,N_14963);
nand UO_399 (O_399,N_14927,N_14891);
and UO_400 (O_400,N_14988,N_14921);
and UO_401 (O_401,N_14958,N_14894);
nand UO_402 (O_402,N_14962,N_14945);
nor UO_403 (O_403,N_14913,N_14981);
nor UO_404 (O_404,N_14895,N_14914);
xor UO_405 (O_405,N_14919,N_14927);
nand UO_406 (O_406,N_14958,N_14932);
nor UO_407 (O_407,N_14962,N_14950);
xnor UO_408 (O_408,N_14913,N_14898);
and UO_409 (O_409,N_14912,N_14995);
nand UO_410 (O_410,N_14900,N_14916);
or UO_411 (O_411,N_14992,N_14902);
nor UO_412 (O_412,N_14948,N_14996);
or UO_413 (O_413,N_14911,N_14941);
and UO_414 (O_414,N_14901,N_14883);
and UO_415 (O_415,N_14965,N_14889);
nor UO_416 (O_416,N_14913,N_14938);
and UO_417 (O_417,N_14877,N_14883);
nand UO_418 (O_418,N_14959,N_14885);
xnor UO_419 (O_419,N_14891,N_14998);
or UO_420 (O_420,N_14893,N_14920);
xor UO_421 (O_421,N_14899,N_14992);
and UO_422 (O_422,N_14875,N_14892);
or UO_423 (O_423,N_14948,N_14959);
and UO_424 (O_424,N_14914,N_14948);
or UO_425 (O_425,N_14962,N_14949);
and UO_426 (O_426,N_14967,N_14907);
or UO_427 (O_427,N_14983,N_14889);
or UO_428 (O_428,N_14996,N_14990);
and UO_429 (O_429,N_14883,N_14982);
xor UO_430 (O_430,N_14970,N_14954);
nor UO_431 (O_431,N_14933,N_14979);
and UO_432 (O_432,N_14921,N_14990);
nand UO_433 (O_433,N_14909,N_14896);
nor UO_434 (O_434,N_14906,N_14899);
or UO_435 (O_435,N_14967,N_14988);
xnor UO_436 (O_436,N_14896,N_14947);
nor UO_437 (O_437,N_14910,N_14980);
and UO_438 (O_438,N_14957,N_14980);
or UO_439 (O_439,N_14971,N_14910);
or UO_440 (O_440,N_14913,N_14983);
or UO_441 (O_441,N_14934,N_14896);
xnor UO_442 (O_442,N_14967,N_14964);
nand UO_443 (O_443,N_14908,N_14890);
and UO_444 (O_444,N_14956,N_14950);
and UO_445 (O_445,N_14880,N_14956);
xnor UO_446 (O_446,N_14903,N_14910);
nand UO_447 (O_447,N_14882,N_14983);
nand UO_448 (O_448,N_14940,N_14888);
xnor UO_449 (O_449,N_14928,N_14984);
nand UO_450 (O_450,N_14875,N_14925);
or UO_451 (O_451,N_14888,N_14950);
xnor UO_452 (O_452,N_14966,N_14954);
nand UO_453 (O_453,N_14885,N_14908);
nand UO_454 (O_454,N_14999,N_14934);
xor UO_455 (O_455,N_14970,N_14925);
and UO_456 (O_456,N_14903,N_14951);
nand UO_457 (O_457,N_14895,N_14911);
or UO_458 (O_458,N_14903,N_14975);
xor UO_459 (O_459,N_14953,N_14999);
and UO_460 (O_460,N_14925,N_14895);
and UO_461 (O_461,N_14955,N_14966);
nand UO_462 (O_462,N_14943,N_14905);
or UO_463 (O_463,N_14983,N_14948);
and UO_464 (O_464,N_14928,N_14903);
and UO_465 (O_465,N_14934,N_14982);
xnor UO_466 (O_466,N_14924,N_14988);
or UO_467 (O_467,N_14970,N_14903);
nand UO_468 (O_468,N_14997,N_14977);
xor UO_469 (O_469,N_14972,N_14883);
and UO_470 (O_470,N_14989,N_14927);
or UO_471 (O_471,N_14900,N_14885);
and UO_472 (O_472,N_14972,N_14986);
and UO_473 (O_473,N_14927,N_14879);
or UO_474 (O_474,N_14928,N_14989);
or UO_475 (O_475,N_14995,N_14974);
and UO_476 (O_476,N_14940,N_14878);
and UO_477 (O_477,N_14916,N_14939);
xnor UO_478 (O_478,N_14876,N_14927);
nor UO_479 (O_479,N_14976,N_14957);
nand UO_480 (O_480,N_14969,N_14971);
nor UO_481 (O_481,N_14914,N_14876);
and UO_482 (O_482,N_14898,N_14934);
nand UO_483 (O_483,N_14916,N_14992);
xor UO_484 (O_484,N_14932,N_14974);
xor UO_485 (O_485,N_14899,N_14951);
and UO_486 (O_486,N_14958,N_14890);
nand UO_487 (O_487,N_14994,N_14905);
nand UO_488 (O_488,N_14896,N_14979);
nand UO_489 (O_489,N_14963,N_14894);
nor UO_490 (O_490,N_14891,N_14907);
nand UO_491 (O_491,N_14959,N_14899);
nand UO_492 (O_492,N_14995,N_14962);
and UO_493 (O_493,N_14914,N_14980);
nand UO_494 (O_494,N_14930,N_14929);
nor UO_495 (O_495,N_14947,N_14909);
nor UO_496 (O_496,N_14911,N_14883);
nand UO_497 (O_497,N_14897,N_14944);
and UO_498 (O_498,N_14926,N_14963);
or UO_499 (O_499,N_14899,N_14881);
nor UO_500 (O_500,N_14949,N_14995);
or UO_501 (O_501,N_14901,N_14956);
xnor UO_502 (O_502,N_14943,N_14931);
nor UO_503 (O_503,N_14951,N_14969);
or UO_504 (O_504,N_14881,N_14895);
nor UO_505 (O_505,N_14923,N_14941);
xnor UO_506 (O_506,N_14928,N_14994);
and UO_507 (O_507,N_14917,N_14954);
nand UO_508 (O_508,N_14931,N_14879);
nand UO_509 (O_509,N_14949,N_14989);
nand UO_510 (O_510,N_14924,N_14878);
nand UO_511 (O_511,N_14966,N_14933);
nor UO_512 (O_512,N_14894,N_14947);
or UO_513 (O_513,N_14982,N_14931);
and UO_514 (O_514,N_14969,N_14920);
or UO_515 (O_515,N_14987,N_14919);
xor UO_516 (O_516,N_14991,N_14912);
nand UO_517 (O_517,N_14967,N_14998);
nor UO_518 (O_518,N_14998,N_14959);
nor UO_519 (O_519,N_14988,N_14893);
or UO_520 (O_520,N_14935,N_14919);
xnor UO_521 (O_521,N_14935,N_14962);
xor UO_522 (O_522,N_14890,N_14879);
nor UO_523 (O_523,N_14911,N_14875);
and UO_524 (O_524,N_14959,N_14890);
or UO_525 (O_525,N_14884,N_14989);
and UO_526 (O_526,N_14894,N_14898);
xnor UO_527 (O_527,N_14937,N_14876);
xor UO_528 (O_528,N_14880,N_14967);
xor UO_529 (O_529,N_14930,N_14968);
or UO_530 (O_530,N_14946,N_14945);
nor UO_531 (O_531,N_14956,N_14983);
xnor UO_532 (O_532,N_14972,N_14980);
or UO_533 (O_533,N_14946,N_14989);
xor UO_534 (O_534,N_14953,N_14962);
nand UO_535 (O_535,N_14974,N_14994);
nand UO_536 (O_536,N_14987,N_14923);
nor UO_537 (O_537,N_14898,N_14929);
nand UO_538 (O_538,N_14933,N_14999);
xor UO_539 (O_539,N_14964,N_14907);
and UO_540 (O_540,N_14983,N_14892);
nand UO_541 (O_541,N_14877,N_14967);
or UO_542 (O_542,N_14937,N_14975);
xnor UO_543 (O_543,N_14956,N_14908);
xor UO_544 (O_544,N_14989,N_14910);
nand UO_545 (O_545,N_14967,N_14978);
nor UO_546 (O_546,N_14972,N_14981);
nor UO_547 (O_547,N_14953,N_14897);
nor UO_548 (O_548,N_14969,N_14979);
nand UO_549 (O_549,N_14884,N_14948);
xnor UO_550 (O_550,N_14955,N_14976);
or UO_551 (O_551,N_14992,N_14895);
or UO_552 (O_552,N_14924,N_14983);
and UO_553 (O_553,N_14977,N_14961);
and UO_554 (O_554,N_14947,N_14995);
nand UO_555 (O_555,N_14930,N_14976);
or UO_556 (O_556,N_14967,N_14949);
xnor UO_557 (O_557,N_14897,N_14954);
xor UO_558 (O_558,N_14969,N_14881);
xor UO_559 (O_559,N_14939,N_14909);
nor UO_560 (O_560,N_14886,N_14960);
nand UO_561 (O_561,N_14968,N_14876);
nor UO_562 (O_562,N_14990,N_14945);
nor UO_563 (O_563,N_14966,N_14987);
or UO_564 (O_564,N_14924,N_14938);
xor UO_565 (O_565,N_14913,N_14875);
nor UO_566 (O_566,N_14993,N_14991);
or UO_567 (O_567,N_14924,N_14992);
nor UO_568 (O_568,N_14945,N_14929);
xor UO_569 (O_569,N_14891,N_14943);
nor UO_570 (O_570,N_14916,N_14889);
or UO_571 (O_571,N_14969,N_14875);
nor UO_572 (O_572,N_14959,N_14981);
and UO_573 (O_573,N_14963,N_14917);
xor UO_574 (O_574,N_14937,N_14926);
nand UO_575 (O_575,N_14901,N_14990);
nand UO_576 (O_576,N_14917,N_14884);
nand UO_577 (O_577,N_14881,N_14957);
nand UO_578 (O_578,N_14974,N_14983);
nor UO_579 (O_579,N_14927,N_14880);
or UO_580 (O_580,N_14904,N_14913);
nor UO_581 (O_581,N_14952,N_14998);
nor UO_582 (O_582,N_14919,N_14944);
nand UO_583 (O_583,N_14893,N_14913);
or UO_584 (O_584,N_14903,N_14884);
and UO_585 (O_585,N_14938,N_14975);
nand UO_586 (O_586,N_14895,N_14878);
xor UO_587 (O_587,N_14878,N_14922);
nor UO_588 (O_588,N_14910,N_14881);
and UO_589 (O_589,N_14907,N_14989);
xnor UO_590 (O_590,N_14882,N_14984);
xor UO_591 (O_591,N_14984,N_14972);
or UO_592 (O_592,N_14955,N_14887);
or UO_593 (O_593,N_14891,N_14917);
and UO_594 (O_594,N_14911,N_14932);
or UO_595 (O_595,N_14981,N_14910);
or UO_596 (O_596,N_14954,N_14881);
xor UO_597 (O_597,N_14944,N_14920);
and UO_598 (O_598,N_14894,N_14969);
nor UO_599 (O_599,N_14941,N_14875);
xnor UO_600 (O_600,N_14955,N_14892);
and UO_601 (O_601,N_14965,N_14948);
and UO_602 (O_602,N_14898,N_14989);
and UO_603 (O_603,N_14979,N_14882);
nand UO_604 (O_604,N_14900,N_14887);
nand UO_605 (O_605,N_14880,N_14962);
and UO_606 (O_606,N_14990,N_14878);
and UO_607 (O_607,N_14927,N_14899);
nor UO_608 (O_608,N_14909,N_14974);
xor UO_609 (O_609,N_14915,N_14991);
xnor UO_610 (O_610,N_14880,N_14929);
nand UO_611 (O_611,N_14944,N_14894);
xor UO_612 (O_612,N_14904,N_14942);
and UO_613 (O_613,N_14998,N_14887);
nor UO_614 (O_614,N_14925,N_14932);
nand UO_615 (O_615,N_14961,N_14914);
xor UO_616 (O_616,N_14955,N_14928);
or UO_617 (O_617,N_14970,N_14962);
nor UO_618 (O_618,N_14972,N_14966);
nand UO_619 (O_619,N_14963,N_14947);
and UO_620 (O_620,N_14912,N_14946);
and UO_621 (O_621,N_14974,N_14915);
nand UO_622 (O_622,N_14944,N_14986);
nand UO_623 (O_623,N_14957,N_14971);
or UO_624 (O_624,N_14988,N_14956);
and UO_625 (O_625,N_14882,N_14997);
xor UO_626 (O_626,N_14927,N_14929);
or UO_627 (O_627,N_14940,N_14945);
nor UO_628 (O_628,N_14875,N_14895);
and UO_629 (O_629,N_14904,N_14999);
and UO_630 (O_630,N_14936,N_14998);
nor UO_631 (O_631,N_14970,N_14924);
nor UO_632 (O_632,N_14975,N_14892);
nor UO_633 (O_633,N_14987,N_14899);
nand UO_634 (O_634,N_14905,N_14910);
nand UO_635 (O_635,N_14949,N_14961);
xor UO_636 (O_636,N_14933,N_14943);
and UO_637 (O_637,N_14884,N_14912);
nand UO_638 (O_638,N_14996,N_14954);
and UO_639 (O_639,N_14910,N_14990);
or UO_640 (O_640,N_14887,N_14977);
nor UO_641 (O_641,N_14886,N_14899);
nor UO_642 (O_642,N_14975,N_14962);
nand UO_643 (O_643,N_14943,N_14976);
nor UO_644 (O_644,N_14922,N_14981);
or UO_645 (O_645,N_14938,N_14877);
nand UO_646 (O_646,N_14901,N_14882);
nor UO_647 (O_647,N_14922,N_14976);
or UO_648 (O_648,N_14915,N_14999);
xnor UO_649 (O_649,N_14933,N_14894);
xnor UO_650 (O_650,N_14943,N_14960);
nand UO_651 (O_651,N_14928,N_14970);
xor UO_652 (O_652,N_14995,N_14976);
nor UO_653 (O_653,N_14970,N_14904);
nand UO_654 (O_654,N_14919,N_14929);
and UO_655 (O_655,N_14996,N_14963);
xor UO_656 (O_656,N_14957,N_14924);
nor UO_657 (O_657,N_14904,N_14953);
nor UO_658 (O_658,N_14959,N_14973);
xor UO_659 (O_659,N_14921,N_14983);
xnor UO_660 (O_660,N_14998,N_14880);
or UO_661 (O_661,N_14885,N_14976);
and UO_662 (O_662,N_14901,N_14942);
nand UO_663 (O_663,N_14916,N_14976);
nand UO_664 (O_664,N_14958,N_14889);
nor UO_665 (O_665,N_14961,N_14952);
or UO_666 (O_666,N_14912,N_14894);
nor UO_667 (O_667,N_14913,N_14941);
and UO_668 (O_668,N_14903,N_14893);
and UO_669 (O_669,N_14904,N_14929);
and UO_670 (O_670,N_14979,N_14943);
nand UO_671 (O_671,N_14911,N_14929);
nor UO_672 (O_672,N_14984,N_14953);
nand UO_673 (O_673,N_14883,N_14891);
and UO_674 (O_674,N_14977,N_14879);
and UO_675 (O_675,N_14926,N_14909);
or UO_676 (O_676,N_14948,N_14917);
xor UO_677 (O_677,N_14903,N_14920);
nor UO_678 (O_678,N_14921,N_14947);
and UO_679 (O_679,N_14967,N_14922);
nor UO_680 (O_680,N_14984,N_14885);
nor UO_681 (O_681,N_14998,N_14892);
nand UO_682 (O_682,N_14951,N_14979);
nand UO_683 (O_683,N_14926,N_14900);
nor UO_684 (O_684,N_14990,N_14946);
xnor UO_685 (O_685,N_14956,N_14890);
nor UO_686 (O_686,N_14982,N_14943);
nand UO_687 (O_687,N_14918,N_14944);
nor UO_688 (O_688,N_14884,N_14984);
or UO_689 (O_689,N_14904,N_14898);
nor UO_690 (O_690,N_14972,N_14906);
nor UO_691 (O_691,N_14920,N_14923);
nor UO_692 (O_692,N_14999,N_14944);
or UO_693 (O_693,N_14916,N_14904);
and UO_694 (O_694,N_14953,N_14892);
xnor UO_695 (O_695,N_14907,N_14922);
xor UO_696 (O_696,N_14980,N_14960);
nand UO_697 (O_697,N_14885,N_14918);
nor UO_698 (O_698,N_14883,N_14890);
nor UO_699 (O_699,N_14917,N_14932);
or UO_700 (O_700,N_14883,N_14954);
and UO_701 (O_701,N_14925,N_14881);
nor UO_702 (O_702,N_14939,N_14975);
and UO_703 (O_703,N_14935,N_14952);
nor UO_704 (O_704,N_14908,N_14991);
nor UO_705 (O_705,N_14897,N_14988);
and UO_706 (O_706,N_14972,N_14995);
and UO_707 (O_707,N_14929,N_14939);
nand UO_708 (O_708,N_14926,N_14896);
and UO_709 (O_709,N_14970,N_14981);
nor UO_710 (O_710,N_14935,N_14975);
nor UO_711 (O_711,N_14929,N_14965);
or UO_712 (O_712,N_14876,N_14949);
and UO_713 (O_713,N_14971,N_14935);
or UO_714 (O_714,N_14926,N_14978);
nand UO_715 (O_715,N_14894,N_14905);
xnor UO_716 (O_716,N_14962,N_14968);
and UO_717 (O_717,N_14950,N_14931);
nand UO_718 (O_718,N_14929,N_14926);
xnor UO_719 (O_719,N_14883,N_14971);
xor UO_720 (O_720,N_14967,N_14906);
or UO_721 (O_721,N_14981,N_14985);
nor UO_722 (O_722,N_14908,N_14999);
xor UO_723 (O_723,N_14976,N_14977);
nand UO_724 (O_724,N_14939,N_14928);
and UO_725 (O_725,N_14889,N_14962);
and UO_726 (O_726,N_14949,N_14973);
nand UO_727 (O_727,N_14918,N_14985);
and UO_728 (O_728,N_14983,N_14969);
xnor UO_729 (O_729,N_14953,N_14975);
nand UO_730 (O_730,N_14890,N_14895);
and UO_731 (O_731,N_14999,N_14987);
xor UO_732 (O_732,N_14937,N_14889);
nor UO_733 (O_733,N_14966,N_14901);
nand UO_734 (O_734,N_14917,N_14913);
nand UO_735 (O_735,N_14925,N_14928);
nor UO_736 (O_736,N_14875,N_14894);
nand UO_737 (O_737,N_14931,N_14918);
or UO_738 (O_738,N_14930,N_14962);
or UO_739 (O_739,N_14887,N_14980);
nor UO_740 (O_740,N_14989,N_14903);
xnor UO_741 (O_741,N_14969,N_14915);
nand UO_742 (O_742,N_14971,N_14958);
nor UO_743 (O_743,N_14986,N_14906);
and UO_744 (O_744,N_14957,N_14905);
xor UO_745 (O_745,N_14914,N_14979);
nor UO_746 (O_746,N_14993,N_14944);
nor UO_747 (O_747,N_14985,N_14980);
or UO_748 (O_748,N_14960,N_14999);
nand UO_749 (O_749,N_14946,N_14897);
or UO_750 (O_750,N_14968,N_14985);
xnor UO_751 (O_751,N_14944,N_14964);
and UO_752 (O_752,N_14905,N_14913);
xnor UO_753 (O_753,N_14905,N_14964);
and UO_754 (O_754,N_14877,N_14984);
nor UO_755 (O_755,N_14989,N_14876);
or UO_756 (O_756,N_14959,N_14918);
or UO_757 (O_757,N_14977,N_14970);
or UO_758 (O_758,N_14981,N_14933);
nand UO_759 (O_759,N_14969,N_14958);
nand UO_760 (O_760,N_14968,N_14934);
nor UO_761 (O_761,N_14990,N_14983);
nor UO_762 (O_762,N_14920,N_14929);
and UO_763 (O_763,N_14900,N_14930);
nand UO_764 (O_764,N_14945,N_14974);
and UO_765 (O_765,N_14900,N_14938);
or UO_766 (O_766,N_14956,N_14984);
xnor UO_767 (O_767,N_14993,N_14996);
nor UO_768 (O_768,N_14899,N_14989);
nor UO_769 (O_769,N_14975,N_14944);
xor UO_770 (O_770,N_14903,N_14925);
nor UO_771 (O_771,N_14890,N_14891);
or UO_772 (O_772,N_14904,N_14962);
nand UO_773 (O_773,N_14930,N_14972);
xnor UO_774 (O_774,N_14937,N_14985);
or UO_775 (O_775,N_14939,N_14883);
and UO_776 (O_776,N_14985,N_14943);
or UO_777 (O_777,N_14995,N_14948);
nor UO_778 (O_778,N_14904,N_14901);
or UO_779 (O_779,N_14927,N_14968);
and UO_780 (O_780,N_14970,N_14930);
and UO_781 (O_781,N_14933,N_14957);
nor UO_782 (O_782,N_14898,N_14964);
nand UO_783 (O_783,N_14933,N_14921);
and UO_784 (O_784,N_14908,N_14986);
nand UO_785 (O_785,N_14908,N_14906);
or UO_786 (O_786,N_14939,N_14992);
or UO_787 (O_787,N_14927,N_14990);
xor UO_788 (O_788,N_14935,N_14974);
xor UO_789 (O_789,N_14982,N_14929);
nand UO_790 (O_790,N_14996,N_14977);
nor UO_791 (O_791,N_14965,N_14891);
xnor UO_792 (O_792,N_14975,N_14996);
nand UO_793 (O_793,N_14991,N_14920);
nor UO_794 (O_794,N_14968,N_14997);
nor UO_795 (O_795,N_14983,N_14893);
nor UO_796 (O_796,N_14882,N_14959);
or UO_797 (O_797,N_14894,N_14970);
or UO_798 (O_798,N_14910,N_14951);
or UO_799 (O_799,N_14915,N_14900);
xnor UO_800 (O_800,N_14989,N_14991);
and UO_801 (O_801,N_14910,N_14887);
or UO_802 (O_802,N_14901,N_14947);
nor UO_803 (O_803,N_14981,N_14951);
nand UO_804 (O_804,N_14895,N_14891);
nand UO_805 (O_805,N_14974,N_14969);
or UO_806 (O_806,N_14889,N_14888);
nand UO_807 (O_807,N_14943,N_14940);
nor UO_808 (O_808,N_14969,N_14963);
xnor UO_809 (O_809,N_14890,N_14975);
or UO_810 (O_810,N_14933,N_14935);
and UO_811 (O_811,N_14998,N_14965);
and UO_812 (O_812,N_14977,N_14911);
and UO_813 (O_813,N_14969,N_14893);
or UO_814 (O_814,N_14933,N_14893);
xnor UO_815 (O_815,N_14876,N_14971);
xnor UO_816 (O_816,N_14883,N_14974);
or UO_817 (O_817,N_14879,N_14972);
nor UO_818 (O_818,N_14968,N_14889);
xor UO_819 (O_819,N_14981,N_14957);
nor UO_820 (O_820,N_14971,N_14990);
or UO_821 (O_821,N_14956,N_14904);
or UO_822 (O_822,N_14952,N_14985);
nor UO_823 (O_823,N_14989,N_14920);
xor UO_824 (O_824,N_14941,N_14956);
or UO_825 (O_825,N_14952,N_14940);
nand UO_826 (O_826,N_14932,N_14961);
and UO_827 (O_827,N_14894,N_14904);
nand UO_828 (O_828,N_14959,N_14967);
xor UO_829 (O_829,N_14932,N_14994);
and UO_830 (O_830,N_14974,N_14951);
or UO_831 (O_831,N_14957,N_14936);
and UO_832 (O_832,N_14962,N_14892);
or UO_833 (O_833,N_14911,N_14991);
nand UO_834 (O_834,N_14921,N_14931);
nor UO_835 (O_835,N_14940,N_14994);
nor UO_836 (O_836,N_14941,N_14987);
nor UO_837 (O_837,N_14923,N_14957);
xnor UO_838 (O_838,N_14919,N_14879);
and UO_839 (O_839,N_14921,N_14985);
nor UO_840 (O_840,N_14937,N_14964);
nand UO_841 (O_841,N_14995,N_14986);
xnor UO_842 (O_842,N_14878,N_14973);
nor UO_843 (O_843,N_14993,N_14891);
or UO_844 (O_844,N_14993,N_14971);
and UO_845 (O_845,N_14897,N_14901);
nor UO_846 (O_846,N_14891,N_14990);
xor UO_847 (O_847,N_14879,N_14951);
nand UO_848 (O_848,N_14879,N_14946);
and UO_849 (O_849,N_14979,N_14938);
nand UO_850 (O_850,N_14964,N_14900);
xor UO_851 (O_851,N_14946,N_14892);
nor UO_852 (O_852,N_14919,N_14952);
xor UO_853 (O_853,N_14937,N_14980);
nor UO_854 (O_854,N_14926,N_14985);
or UO_855 (O_855,N_14960,N_14913);
xnor UO_856 (O_856,N_14963,N_14932);
nand UO_857 (O_857,N_14902,N_14972);
nand UO_858 (O_858,N_14973,N_14926);
nand UO_859 (O_859,N_14885,N_14909);
or UO_860 (O_860,N_14942,N_14973);
or UO_861 (O_861,N_14880,N_14923);
or UO_862 (O_862,N_14932,N_14985);
and UO_863 (O_863,N_14925,N_14945);
or UO_864 (O_864,N_14877,N_14951);
or UO_865 (O_865,N_14998,N_14984);
and UO_866 (O_866,N_14896,N_14929);
xor UO_867 (O_867,N_14942,N_14885);
xor UO_868 (O_868,N_14911,N_14995);
or UO_869 (O_869,N_14949,N_14914);
and UO_870 (O_870,N_14951,N_14949);
or UO_871 (O_871,N_14973,N_14891);
nor UO_872 (O_872,N_14939,N_14998);
and UO_873 (O_873,N_14877,N_14974);
nand UO_874 (O_874,N_14951,N_14922);
nand UO_875 (O_875,N_14928,N_14960);
nor UO_876 (O_876,N_14930,N_14984);
xnor UO_877 (O_877,N_14981,N_14889);
and UO_878 (O_878,N_14988,N_14918);
and UO_879 (O_879,N_14976,N_14876);
xnor UO_880 (O_880,N_14906,N_14952);
nor UO_881 (O_881,N_14902,N_14948);
and UO_882 (O_882,N_14935,N_14930);
and UO_883 (O_883,N_14973,N_14923);
nand UO_884 (O_884,N_14967,N_14939);
xor UO_885 (O_885,N_14881,N_14983);
nand UO_886 (O_886,N_14969,N_14892);
nand UO_887 (O_887,N_14949,N_14956);
or UO_888 (O_888,N_14986,N_14904);
or UO_889 (O_889,N_14901,N_14960);
nor UO_890 (O_890,N_14942,N_14875);
xor UO_891 (O_891,N_14922,N_14910);
and UO_892 (O_892,N_14879,N_14945);
nand UO_893 (O_893,N_14925,N_14880);
xor UO_894 (O_894,N_14965,N_14983);
or UO_895 (O_895,N_14988,N_14948);
nand UO_896 (O_896,N_14927,N_14940);
or UO_897 (O_897,N_14970,N_14911);
nor UO_898 (O_898,N_14877,N_14912);
xor UO_899 (O_899,N_14901,N_14974);
nand UO_900 (O_900,N_14953,N_14998);
and UO_901 (O_901,N_14996,N_14902);
nand UO_902 (O_902,N_14995,N_14953);
xor UO_903 (O_903,N_14937,N_14979);
nor UO_904 (O_904,N_14922,N_14943);
nand UO_905 (O_905,N_14962,N_14906);
nand UO_906 (O_906,N_14902,N_14994);
xor UO_907 (O_907,N_14977,N_14958);
xnor UO_908 (O_908,N_14953,N_14933);
xor UO_909 (O_909,N_14985,N_14915);
or UO_910 (O_910,N_14919,N_14942);
nand UO_911 (O_911,N_14935,N_14943);
xor UO_912 (O_912,N_14982,N_14885);
and UO_913 (O_913,N_14970,N_14921);
nand UO_914 (O_914,N_14913,N_14881);
xnor UO_915 (O_915,N_14974,N_14916);
nand UO_916 (O_916,N_14885,N_14951);
nand UO_917 (O_917,N_14949,N_14918);
nand UO_918 (O_918,N_14917,N_14878);
and UO_919 (O_919,N_14959,N_14876);
or UO_920 (O_920,N_14894,N_14948);
and UO_921 (O_921,N_14952,N_14990);
nand UO_922 (O_922,N_14909,N_14901);
and UO_923 (O_923,N_14879,N_14893);
nand UO_924 (O_924,N_14879,N_14991);
and UO_925 (O_925,N_14880,N_14963);
or UO_926 (O_926,N_14938,N_14981);
and UO_927 (O_927,N_14932,N_14876);
nand UO_928 (O_928,N_14883,N_14946);
or UO_929 (O_929,N_14932,N_14942);
xor UO_930 (O_930,N_14976,N_14918);
and UO_931 (O_931,N_14888,N_14973);
nor UO_932 (O_932,N_14976,N_14925);
nor UO_933 (O_933,N_14912,N_14940);
nor UO_934 (O_934,N_14956,N_14995);
nand UO_935 (O_935,N_14900,N_14912);
and UO_936 (O_936,N_14906,N_14918);
and UO_937 (O_937,N_14994,N_14903);
or UO_938 (O_938,N_14906,N_14914);
nand UO_939 (O_939,N_14995,N_14978);
nand UO_940 (O_940,N_14991,N_14971);
nand UO_941 (O_941,N_14884,N_14973);
nor UO_942 (O_942,N_14906,N_14884);
or UO_943 (O_943,N_14937,N_14952);
xor UO_944 (O_944,N_14923,N_14909);
xor UO_945 (O_945,N_14926,N_14990);
nor UO_946 (O_946,N_14989,N_14881);
xnor UO_947 (O_947,N_14887,N_14988);
and UO_948 (O_948,N_14992,N_14994);
or UO_949 (O_949,N_14938,N_14911);
and UO_950 (O_950,N_14908,N_14881);
and UO_951 (O_951,N_14930,N_14974);
xnor UO_952 (O_952,N_14950,N_14890);
nand UO_953 (O_953,N_14877,N_14937);
nor UO_954 (O_954,N_14880,N_14876);
nand UO_955 (O_955,N_14996,N_14890);
or UO_956 (O_956,N_14881,N_14884);
nor UO_957 (O_957,N_14927,N_14942);
and UO_958 (O_958,N_14905,N_14877);
or UO_959 (O_959,N_14879,N_14937);
nor UO_960 (O_960,N_14937,N_14943);
nand UO_961 (O_961,N_14876,N_14975);
xor UO_962 (O_962,N_14973,N_14875);
and UO_963 (O_963,N_14920,N_14892);
nor UO_964 (O_964,N_14879,N_14952);
nor UO_965 (O_965,N_14964,N_14981);
and UO_966 (O_966,N_14917,N_14951);
or UO_967 (O_967,N_14952,N_14964);
xor UO_968 (O_968,N_14920,N_14982);
and UO_969 (O_969,N_14877,N_14903);
xnor UO_970 (O_970,N_14958,N_14909);
xnor UO_971 (O_971,N_14970,N_14956);
nand UO_972 (O_972,N_14975,N_14950);
nor UO_973 (O_973,N_14886,N_14934);
nor UO_974 (O_974,N_14881,N_14951);
xnor UO_975 (O_975,N_14917,N_14961);
xnor UO_976 (O_976,N_14954,N_14952);
nor UO_977 (O_977,N_14973,N_14997);
and UO_978 (O_978,N_14929,N_14990);
xnor UO_979 (O_979,N_14890,N_14948);
xor UO_980 (O_980,N_14994,N_14959);
nor UO_981 (O_981,N_14919,N_14995);
and UO_982 (O_982,N_14903,N_14934);
and UO_983 (O_983,N_14896,N_14894);
nand UO_984 (O_984,N_14942,N_14929);
or UO_985 (O_985,N_14910,N_14929);
nor UO_986 (O_986,N_14918,N_14876);
xnor UO_987 (O_987,N_14956,N_14884);
nand UO_988 (O_988,N_14937,N_14918);
nor UO_989 (O_989,N_14916,N_14888);
nand UO_990 (O_990,N_14929,N_14962);
nor UO_991 (O_991,N_14904,N_14879);
nor UO_992 (O_992,N_14939,N_14970);
or UO_993 (O_993,N_14916,N_14942);
or UO_994 (O_994,N_14905,N_14915);
and UO_995 (O_995,N_14879,N_14922);
nand UO_996 (O_996,N_14920,N_14896);
or UO_997 (O_997,N_14907,N_14952);
or UO_998 (O_998,N_14980,N_14895);
xnor UO_999 (O_999,N_14886,N_14938);
and UO_1000 (O_1000,N_14990,N_14882);
or UO_1001 (O_1001,N_14950,N_14894);
or UO_1002 (O_1002,N_14895,N_14931);
nand UO_1003 (O_1003,N_14936,N_14906);
xnor UO_1004 (O_1004,N_14987,N_14988);
nor UO_1005 (O_1005,N_14887,N_14985);
nand UO_1006 (O_1006,N_14992,N_14901);
or UO_1007 (O_1007,N_14905,N_14886);
xnor UO_1008 (O_1008,N_14883,N_14885);
xnor UO_1009 (O_1009,N_14948,N_14971);
nand UO_1010 (O_1010,N_14941,N_14954);
and UO_1011 (O_1011,N_14943,N_14957);
xnor UO_1012 (O_1012,N_14956,N_14902);
nor UO_1013 (O_1013,N_14887,N_14906);
or UO_1014 (O_1014,N_14889,N_14920);
or UO_1015 (O_1015,N_14974,N_14990);
xnor UO_1016 (O_1016,N_14920,N_14885);
xnor UO_1017 (O_1017,N_14912,N_14947);
nor UO_1018 (O_1018,N_14999,N_14885);
or UO_1019 (O_1019,N_14958,N_14986);
nor UO_1020 (O_1020,N_14919,N_14877);
xor UO_1021 (O_1021,N_14972,N_14977);
nor UO_1022 (O_1022,N_14984,N_14921);
nand UO_1023 (O_1023,N_14982,N_14981);
nand UO_1024 (O_1024,N_14934,N_14892);
nor UO_1025 (O_1025,N_14940,N_14896);
nand UO_1026 (O_1026,N_14890,N_14937);
xor UO_1027 (O_1027,N_14912,N_14917);
nand UO_1028 (O_1028,N_14878,N_14899);
or UO_1029 (O_1029,N_14977,N_14943);
xnor UO_1030 (O_1030,N_14988,N_14975);
or UO_1031 (O_1031,N_14956,N_14912);
and UO_1032 (O_1032,N_14969,N_14942);
and UO_1033 (O_1033,N_14921,N_14924);
and UO_1034 (O_1034,N_14920,N_14933);
or UO_1035 (O_1035,N_14964,N_14887);
xnor UO_1036 (O_1036,N_14950,N_14974);
xnor UO_1037 (O_1037,N_14991,N_14951);
and UO_1038 (O_1038,N_14929,N_14983);
xor UO_1039 (O_1039,N_14985,N_14963);
and UO_1040 (O_1040,N_14953,N_14880);
and UO_1041 (O_1041,N_14985,N_14882);
nand UO_1042 (O_1042,N_14911,N_14984);
nor UO_1043 (O_1043,N_14905,N_14951);
nand UO_1044 (O_1044,N_14984,N_14985);
and UO_1045 (O_1045,N_14896,N_14884);
or UO_1046 (O_1046,N_14955,N_14993);
or UO_1047 (O_1047,N_14935,N_14963);
nor UO_1048 (O_1048,N_14876,N_14946);
and UO_1049 (O_1049,N_14893,N_14942);
xnor UO_1050 (O_1050,N_14948,N_14969);
xnor UO_1051 (O_1051,N_14912,N_14930);
nor UO_1052 (O_1052,N_14889,N_14892);
or UO_1053 (O_1053,N_14955,N_14899);
xor UO_1054 (O_1054,N_14903,N_14886);
xor UO_1055 (O_1055,N_14985,N_14991);
nor UO_1056 (O_1056,N_14887,N_14958);
nand UO_1057 (O_1057,N_14963,N_14954);
nand UO_1058 (O_1058,N_14978,N_14880);
nor UO_1059 (O_1059,N_14976,N_14967);
or UO_1060 (O_1060,N_14901,N_14916);
or UO_1061 (O_1061,N_14887,N_14936);
or UO_1062 (O_1062,N_14969,N_14985);
and UO_1063 (O_1063,N_14932,N_14916);
xnor UO_1064 (O_1064,N_14994,N_14897);
or UO_1065 (O_1065,N_14897,N_14967);
xnor UO_1066 (O_1066,N_14984,N_14992);
xnor UO_1067 (O_1067,N_14992,N_14896);
nand UO_1068 (O_1068,N_14942,N_14977);
nor UO_1069 (O_1069,N_14907,N_14943);
and UO_1070 (O_1070,N_14916,N_14981);
nor UO_1071 (O_1071,N_14919,N_14979);
nor UO_1072 (O_1072,N_14935,N_14940);
and UO_1073 (O_1073,N_14968,N_14900);
and UO_1074 (O_1074,N_14939,N_14937);
and UO_1075 (O_1075,N_14879,N_14944);
and UO_1076 (O_1076,N_14987,N_14935);
xor UO_1077 (O_1077,N_14916,N_14941);
nand UO_1078 (O_1078,N_14925,N_14920);
nand UO_1079 (O_1079,N_14984,N_14970);
xnor UO_1080 (O_1080,N_14988,N_14938);
nand UO_1081 (O_1081,N_14878,N_14928);
and UO_1082 (O_1082,N_14895,N_14916);
and UO_1083 (O_1083,N_14953,N_14926);
xor UO_1084 (O_1084,N_14990,N_14976);
nor UO_1085 (O_1085,N_14931,N_14894);
nand UO_1086 (O_1086,N_14905,N_14947);
xnor UO_1087 (O_1087,N_14982,N_14952);
or UO_1088 (O_1088,N_14893,N_14978);
and UO_1089 (O_1089,N_14918,N_14925);
nand UO_1090 (O_1090,N_14880,N_14926);
and UO_1091 (O_1091,N_14889,N_14913);
nand UO_1092 (O_1092,N_14908,N_14901);
xnor UO_1093 (O_1093,N_14946,N_14991);
nand UO_1094 (O_1094,N_14957,N_14948);
nor UO_1095 (O_1095,N_14992,N_14904);
nor UO_1096 (O_1096,N_14951,N_14984);
or UO_1097 (O_1097,N_14938,N_14932);
xor UO_1098 (O_1098,N_14944,N_14985);
nand UO_1099 (O_1099,N_14908,N_14883);
nand UO_1100 (O_1100,N_14924,N_14964);
nand UO_1101 (O_1101,N_14912,N_14908);
and UO_1102 (O_1102,N_14925,N_14886);
xor UO_1103 (O_1103,N_14981,N_14912);
and UO_1104 (O_1104,N_14988,N_14923);
and UO_1105 (O_1105,N_14885,N_14932);
xnor UO_1106 (O_1106,N_14918,N_14884);
nor UO_1107 (O_1107,N_14894,N_14901);
and UO_1108 (O_1108,N_14982,N_14963);
xnor UO_1109 (O_1109,N_14916,N_14938);
and UO_1110 (O_1110,N_14912,N_14952);
nor UO_1111 (O_1111,N_14897,N_14921);
nor UO_1112 (O_1112,N_14876,N_14992);
xor UO_1113 (O_1113,N_14883,N_14957);
xor UO_1114 (O_1114,N_14923,N_14991);
or UO_1115 (O_1115,N_14946,N_14916);
xnor UO_1116 (O_1116,N_14939,N_14987);
xnor UO_1117 (O_1117,N_14987,N_14888);
and UO_1118 (O_1118,N_14998,N_14882);
xor UO_1119 (O_1119,N_14930,N_14999);
xnor UO_1120 (O_1120,N_14912,N_14899);
and UO_1121 (O_1121,N_14976,N_14901);
nor UO_1122 (O_1122,N_14937,N_14891);
and UO_1123 (O_1123,N_14987,N_14900);
xnor UO_1124 (O_1124,N_14961,N_14927);
and UO_1125 (O_1125,N_14883,N_14956);
and UO_1126 (O_1126,N_14908,N_14888);
nand UO_1127 (O_1127,N_14934,N_14915);
nor UO_1128 (O_1128,N_14997,N_14922);
nor UO_1129 (O_1129,N_14971,N_14914);
and UO_1130 (O_1130,N_14914,N_14973);
or UO_1131 (O_1131,N_14991,N_14957);
xor UO_1132 (O_1132,N_14907,N_14931);
nand UO_1133 (O_1133,N_14959,N_14906);
nand UO_1134 (O_1134,N_14999,N_14957);
nor UO_1135 (O_1135,N_14999,N_14997);
and UO_1136 (O_1136,N_14921,N_14888);
nand UO_1137 (O_1137,N_14893,N_14881);
xor UO_1138 (O_1138,N_14967,N_14984);
nor UO_1139 (O_1139,N_14997,N_14940);
xnor UO_1140 (O_1140,N_14964,N_14976);
nor UO_1141 (O_1141,N_14997,N_14949);
or UO_1142 (O_1142,N_14989,N_14960);
or UO_1143 (O_1143,N_14961,N_14957);
xnor UO_1144 (O_1144,N_14960,N_14898);
nand UO_1145 (O_1145,N_14949,N_14965);
and UO_1146 (O_1146,N_14977,N_14924);
or UO_1147 (O_1147,N_14979,N_14917);
nand UO_1148 (O_1148,N_14890,N_14995);
nand UO_1149 (O_1149,N_14911,N_14966);
and UO_1150 (O_1150,N_14996,N_14912);
or UO_1151 (O_1151,N_14927,N_14907);
nand UO_1152 (O_1152,N_14918,N_14991);
nand UO_1153 (O_1153,N_14955,N_14954);
nor UO_1154 (O_1154,N_14889,N_14914);
xnor UO_1155 (O_1155,N_14951,N_14955);
xor UO_1156 (O_1156,N_14932,N_14922);
and UO_1157 (O_1157,N_14925,N_14987);
nor UO_1158 (O_1158,N_14880,N_14995);
nand UO_1159 (O_1159,N_14951,N_14997);
xnor UO_1160 (O_1160,N_14931,N_14888);
xnor UO_1161 (O_1161,N_14976,N_14965);
nand UO_1162 (O_1162,N_14932,N_14884);
xor UO_1163 (O_1163,N_14943,N_14954);
xor UO_1164 (O_1164,N_14897,N_14969);
nor UO_1165 (O_1165,N_14912,N_14931);
or UO_1166 (O_1166,N_14936,N_14902);
nand UO_1167 (O_1167,N_14950,N_14934);
xnor UO_1168 (O_1168,N_14960,N_14947);
and UO_1169 (O_1169,N_14896,N_14983);
nand UO_1170 (O_1170,N_14917,N_14983);
xnor UO_1171 (O_1171,N_14951,N_14986);
and UO_1172 (O_1172,N_14955,N_14911);
nor UO_1173 (O_1173,N_14989,N_14938);
or UO_1174 (O_1174,N_14898,N_14959);
or UO_1175 (O_1175,N_14901,N_14903);
or UO_1176 (O_1176,N_14898,N_14881);
and UO_1177 (O_1177,N_14926,N_14915);
xor UO_1178 (O_1178,N_14958,N_14923);
nand UO_1179 (O_1179,N_14882,N_14950);
nor UO_1180 (O_1180,N_14987,N_14998);
or UO_1181 (O_1181,N_14951,N_14960);
nor UO_1182 (O_1182,N_14897,N_14936);
or UO_1183 (O_1183,N_14905,N_14898);
xor UO_1184 (O_1184,N_14963,N_14995);
nor UO_1185 (O_1185,N_14962,N_14875);
or UO_1186 (O_1186,N_14991,N_14927);
xor UO_1187 (O_1187,N_14906,N_14943);
nor UO_1188 (O_1188,N_14900,N_14922);
and UO_1189 (O_1189,N_14974,N_14936);
and UO_1190 (O_1190,N_14946,N_14913);
nand UO_1191 (O_1191,N_14931,N_14897);
xnor UO_1192 (O_1192,N_14885,N_14888);
and UO_1193 (O_1193,N_14894,N_14964);
xnor UO_1194 (O_1194,N_14925,N_14890);
nand UO_1195 (O_1195,N_14934,N_14925);
xor UO_1196 (O_1196,N_14989,N_14993);
nor UO_1197 (O_1197,N_14973,N_14972);
nand UO_1198 (O_1198,N_14929,N_14994);
or UO_1199 (O_1199,N_14989,N_14973);
and UO_1200 (O_1200,N_14902,N_14913);
or UO_1201 (O_1201,N_14964,N_14893);
nor UO_1202 (O_1202,N_14917,N_14881);
and UO_1203 (O_1203,N_14876,N_14963);
and UO_1204 (O_1204,N_14949,N_14898);
nand UO_1205 (O_1205,N_14994,N_14981);
and UO_1206 (O_1206,N_14977,N_14928);
or UO_1207 (O_1207,N_14893,N_14923);
xor UO_1208 (O_1208,N_14978,N_14952);
nor UO_1209 (O_1209,N_14974,N_14944);
xor UO_1210 (O_1210,N_14885,N_14992);
nand UO_1211 (O_1211,N_14926,N_14898);
nand UO_1212 (O_1212,N_14966,N_14980);
and UO_1213 (O_1213,N_14965,N_14980);
nand UO_1214 (O_1214,N_14902,N_14944);
nor UO_1215 (O_1215,N_14891,N_14999);
xor UO_1216 (O_1216,N_14902,N_14912);
or UO_1217 (O_1217,N_14971,N_14950);
or UO_1218 (O_1218,N_14908,N_14898);
nand UO_1219 (O_1219,N_14977,N_14994);
nand UO_1220 (O_1220,N_14945,N_14924);
or UO_1221 (O_1221,N_14885,N_14928);
and UO_1222 (O_1222,N_14906,N_14941);
nor UO_1223 (O_1223,N_14965,N_14999);
nand UO_1224 (O_1224,N_14941,N_14947);
nor UO_1225 (O_1225,N_14884,N_14920);
xor UO_1226 (O_1226,N_14953,N_14987);
nand UO_1227 (O_1227,N_14951,N_14989);
or UO_1228 (O_1228,N_14963,N_14895);
or UO_1229 (O_1229,N_14943,N_14928);
xnor UO_1230 (O_1230,N_14982,N_14909);
nand UO_1231 (O_1231,N_14935,N_14946);
and UO_1232 (O_1232,N_14937,N_14894);
nor UO_1233 (O_1233,N_14960,N_14957);
xnor UO_1234 (O_1234,N_14980,N_14973);
nand UO_1235 (O_1235,N_14945,N_14902);
xor UO_1236 (O_1236,N_14966,N_14936);
and UO_1237 (O_1237,N_14894,N_14934);
or UO_1238 (O_1238,N_14925,N_14914);
nand UO_1239 (O_1239,N_14979,N_14993);
or UO_1240 (O_1240,N_14879,N_14935);
and UO_1241 (O_1241,N_14982,N_14889);
and UO_1242 (O_1242,N_14988,N_14913);
or UO_1243 (O_1243,N_14962,N_14912);
nand UO_1244 (O_1244,N_14948,N_14921);
or UO_1245 (O_1245,N_14933,N_14897);
or UO_1246 (O_1246,N_14893,N_14958);
xor UO_1247 (O_1247,N_14960,N_14912);
nor UO_1248 (O_1248,N_14913,N_14980);
nand UO_1249 (O_1249,N_14975,N_14912);
and UO_1250 (O_1250,N_14907,N_14883);
and UO_1251 (O_1251,N_14972,N_14978);
nand UO_1252 (O_1252,N_14956,N_14930);
xnor UO_1253 (O_1253,N_14994,N_14990);
xor UO_1254 (O_1254,N_14941,N_14976);
or UO_1255 (O_1255,N_14903,N_14960);
nor UO_1256 (O_1256,N_14886,N_14955);
and UO_1257 (O_1257,N_14929,N_14900);
and UO_1258 (O_1258,N_14928,N_14979);
or UO_1259 (O_1259,N_14959,N_14974);
or UO_1260 (O_1260,N_14992,N_14893);
nand UO_1261 (O_1261,N_14919,N_14998);
or UO_1262 (O_1262,N_14923,N_14889);
or UO_1263 (O_1263,N_14945,N_14992);
xnor UO_1264 (O_1264,N_14936,N_14949);
and UO_1265 (O_1265,N_14988,N_14941);
or UO_1266 (O_1266,N_14946,N_14981);
and UO_1267 (O_1267,N_14989,N_14945);
or UO_1268 (O_1268,N_14945,N_14971);
or UO_1269 (O_1269,N_14921,N_14959);
xor UO_1270 (O_1270,N_14888,N_14965);
and UO_1271 (O_1271,N_14881,N_14998);
and UO_1272 (O_1272,N_14946,N_14927);
or UO_1273 (O_1273,N_14933,N_14899);
xnor UO_1274 (O_1274,N_14977,N_14913);
or UO_1275 (O_1275,N_14896,N_14955);
xnor UO_1276 (O_1276,N_14902,N_14881);
or UO_1277 (O_1277,N_14884,N_14891);
and UO_1278 (O_1278,N_14980,N_14882);
and UO_1279 (O_1279,N_14897,N_14943);
xor UO_1280 (O_1280,N_14903,N_14954);
or UO_1281 (O_1281,N_14985,N_14889);
xor UO_1282 (O_1282,N_14896,N_14963);
or UO_1283 (O_1283,N_14907,N_14901);
nand UO_1284 (O_1284,N_14981,N_14877);
nand UO_1285 (O_1285,N_14991,N_14952);
nor UO_1286 (O_1286,N_14948,N_14968);
and UO_1287 (O_1287,N_14952,N_14895);
nand UO_1288 (O_1288,N_14929,N_14948);
nor UO_1289 (O_1289,N_14999,N_14926);
or UO_1290 (O_1290,N_14924,N_14942);
nor UO_1291 (O_1291,N_14944,N_14958);
nand UO_1292 (O_1292,N_14974,N_14926);
xnor UO_1293 (O_1293,N_14978,N_14953);
xor UO_1294 (O_1294,N_14933,N_14878);
nand UO_1295 (O_1295,N_14967,N_14942);
xnor UO_1296 (O_1296,N_14991,N_14919);
or UO_1297 (O_1297,N_14908,N_14963);
and UO_1298 (O_1298,N_14978,N_14985);
xnor UO_1299 (O_1299,N_14968,N_14920);
and UO_1300 (O_1300,N_14918,N_14963);
xnor UO_1301 (O_1301,N_14977,N_14888);
or UO_1302 (O_1302,N_14946,N_14889);
nand UO_1303 (O_1303,N_14927,N_14937);
nor UO_1304 (O_1304,N_14878,N_14903);
nor UO_1305 (O_1305,N_14945,N_14878);
nor UO_1306 (O_1306,N_14966,N_14924);
nor UO_1307 (O_1307,N_14949,N_14924);
nor UO_1308 (O_1308,N_14931,N_14954);
xor UO_1309 (O_1309,N_14896,N_14984);
nor UO_1310 (O_1310,N_14982,N_14984);
or UO_1311 (O_1311,N_14958,N_14925);
nor UO_1312 (O_1312,N_14889,N_14924);
xor UO_1313 (O_1313,N_14924,N_14961);
xnor UO_1314 (O_1314,N_14905,N_14952);
xnor UO_1315 (O_1315,N_14929,N_14986);
nand UO_1316 (O_1316,N_14912,N_14926);
or UO_1317 (O_1317,N_14953,N_14982);
or UO_1318 (O_1318,N_14936,N_14881);
and UO_1319 (O_1319,N_14922,N_14883);
nand UO_1320 (O_1320,N_14942,N_14925);
nor UO_1321 (O_1321,N_14949,N_14938);
or UO_1322 (O_1322,N_14936,N_14928);
and UO_1323 (O_1323,N_14904,N_14954);
and UO_1324 (O_1324,N_14995,N_14957);
xnor UO_1325 (O_1325,N_14952,N_14892);
nor UO_1326 (O_1326,N_14882,N_14900);
or UO_1327 (O_1327,N_14986,N_14909);
xor UO_1328 (O_1328,N_14976,N_14921);
nand UO_1329 (O_1329,N_14961,N_14963);
or UO_1330 (O_1330,N_14973,N_14911);
xnor UO_1331 (O_1331,N_14941,N_14893);
xor UO_1332 (O_1332,N_14941,N_14908);
nand UO_1333 (O_1333,N_14935,N_14899);
or UO_1334 (O_1334,N_14917,N_14875);
or UO_1335 (O_1335,N_14975,N_14955);
xor UO_1336 (O_1336,N_14881,N_14901);
or UO_1337 (O_1337,N_14886,N_14990);
nor UO_1338 (O_1338,N_14986,N_14947);
and UO_1339 (O_1339,N_14898,N_14883);
xnor UO_1340 (O_1340,N_14921,N_14986);
nand UO_1341 (O_1341,N_14932,N_14987);
or UO_1342 (O_1342,N_14935,N_14986);
nand UO_1343 (O_1343,N_14988,N_14957);
or UO_1344 (O_1344,N_14934,N_14918);
xor UO_1345 (O_1345,N_14902,N_14935);
and UO_1346 (O_1346,N_14984,N_14948);
or UO_1347 (O_1347,N_14926,N_14886);
nand UO_1348 (O_1348,N_14875,N_14914);
or UO_1349 (O_1349,N_14943,N_14970);
and UO_1350 (O_1350,N_14952,N_14994);
nor UO_1351 (O_1351,N_14986,N_14932);
or UO_1352 (O_1352,N_14892,N_14986);
nand UO_1353 (O_1353,N_14903,N_14942);
nand UO_1354 (O_1354,N_14879,N_14903);
nor UO_1355 (O_1355,N_14879,N_14924);
or UO_1356 (O_1356,N_14944,N_14931);
or UO_1357 (O_1357,N_14905,N_14995);
xnor UO_1358 (O_1358,N_14919,N_14909);
xor UO_1359 (O_1359,N_14927,N_14883);
and UO_1360 (O_1360,N_14976,N_14956);
xnor UO_1361 (O_1361,N_14990,N_14957);
or UO_1362 (O_1362,N_14983,N_14930);
nor UO_1363 (O_1363,N_14981,N_14934);
nor UO_1364 (O_1364,N_14884,N_14879);
or UO_1365 (O_1365,N_14977,N_14950);
xnor UO_1366 (O_1366,N_14906,N_14886);
nor UO_1367 (O_1367,N_14987,N_14884);
and UO_1368 (O_1368,N_14988,N_14990);
or UO_1369 (O_1369,N_14948,N_14924);
xnor UO_1370 (O_1370,N_14992,N_14933);
xor UO_1371 (O_1371,N_14967,N_14937);
nand UO_1372 (O_1372,N_14985,N_14974);
or UO_1373 (O_1373,N_14970,N_14881);
or UO_1374 (O_1374,N_14962,N_14905);
or UO_1375 (O_1375,N_14930,N_14989);
nor UO_1376 (O_1376,N_14938,N_14925);
nor UO_1377 (O_1377,N_14976,N_14881);
nand UO_1378 (O_1378,N_14986,N_14888);
nor UO_1379 (O_1379,N_14999,N_14980);
nor UO_1380 (O_1380,N_14997,N_14928);
nand UO_1381 (O_1381,N_14890,N_14965);
xor UO_1382 (O_1382,N_14919,N_14918);
nand UO_1383 (O_1383,N_14953,N_14947);
nor UO_1384 (O_1384,N_14956,N_14927);
nand UO_1385 (O_1385,N_14974,N_14958);
xnor UO_1386 (O_1386,N_14968,N_14909);
and UO_1387 (O_1387,N_14929,N_14992);
xnor UO_1388 (O_1388,N_14965,N_14884);
and UO_1389 (O_1389,N_14884,N_14945);
nor UO_1390 (O_1390,N_14878,N_14953);
nand UO_1391 (O_1391,N_14889,N_14970);
and UO_1392 (O_1392,N_14983,N_14944);
xnor UO_1393 (O_1393,N_14976,N_14898);
nand UO_1394 (O_1394,N_14933,N_14926);
or UO_1395 (O_1395,N_14990,N_14987);
nor UO_1396 (O_1396,N_14999,N_14921);
and UO_1397 (O_1397,N_14936,N_14983);
xnor UO_1398 (O_1398,N_14891,N_14910);
nor UO_1399 (O_1399,N_14875,N_14889);
or UO_1400 (O_1400,N_14875,N_14932);
xnor UO_1401 (O_1401,N_14967,N_14924);
nand UO_1402 (O_1402,N_14966,N_14992);
and UO_1403 (O_1403,N_14936,N_14890);
xnor UO_1404 (O_1404,N_14884,N_14923);
and UO_1405 (O_1405,N_14949,N_14878);
nand UO_1406 (O_1406,N_14966,N_14974);
nand UO_1407 (O_1407,N_14957,N_14910);
and UO_1408 (O_1408,N_14973,N_14917);
nand UO_1409 (O_1409,N_14949,N_14943);
or UO_1410 (O_1410,N_14992,N_14996);
nand UO_1411 (O_1411,N_14999,N_14912);
nand UO_1412 (O_1412,N_14883,N_14965);
and UO_1413 (O_1413,N_14947,N_14875);
xnor UO_1414 (O_1414,N_14988,N_14965);
and UO_1415 (O_1415,N_14979,N_14973);
or UO_1416 (O_1416,N_14930,N_14879);
xor UO_1417 (O_1417,N_14930,N_14977);
nand UO_1418 (O_1418,N_14983,N_14971);
xnor UO_1419 (O_1419,N_14898,N_14953);
xor UO_1420 (O_1420,N_14953,N_14983);
and UO_1421 (O_1421,N_14964,N_14968);
nand UO_1422 (O_1422,N_14930,N_14991);
or UO_1423 (O_1423,N_14882,N_14938);
or UO_1424 (O_1424,N_14882,N_14949);
xnor UO_1425 (O_1425,N_14898,N_14965);
nor UO_1426 (O_1426,N_14978,N_14898);
xor UO_1427 (O_1427,N_14949,N_14908);
xnor UO_1428 (O_1428,N_14879,N_14973);
and UO_1429 (O_1429,N_14937,N_14907);
or UO_1430 (O_1430,N_14922,N_14996);
and UO_1431 (O_1431,N_14962,N_14964);
nand UO_1432 (O_1432,N_14984,N_14946);
nand UO_1433 (O_1433,N_14997,N_14919);
nand UO_1434 (O_1434,N_14940,N_14890);
or UO_1435 (O_1435,N_14976,N_14951);
nor UO_1436 (O_1436,N_14899,N_14891);
nor UO_1437 (O_1437,N_14983,N_14937);
or UO_1438 (O_1438,N_14975,N_14997);
nor UO_1439 (O_1439,N_14908,N_14935);
nand UO_1440 (O_1440,N_14987,N_14967);
and UO_1441 (O_1441,N_14989,N_14921);
and UO_1442 (O_1442,N_14995,N_14938);
nand UO_1443 (O_1443,N_14918,N_14994);
or UO_1444 (O_1444,N_14887,N_14877);
xnor UO_1445 (O_1445,N_14883,N_14992);
or UO_1446 (O_1446,N_14966,N_14960);
nor UO_1447 (O_1447,N_14979,N_14999);
and UO_1448 (O_1448,N_14911,N_14933);
nand UO_1449 (O_1449,N_14892,N_14931);
nand UO_1450 (O_1450,N_14994,N_14912);
and UO_1451 (O_1451,N_14916,N_14994);
xor UO_1452 (O_1452,N_14889,N_14969);
or UO_1453 (O_1453,N_14916,N_14977);
xor UO_1454 (O_1454,N_14877,N_14915);
nand UO_1455 (O_1455,N_14959,N_14992);
xor UO_1456 (O_1456,N_14979,N_14912);
or UO_1457 (O_1457,N_14945,N_14897);
or UO_1458 (O_1458,N_14890,N_14979);
or UO_1459 (O_1459,N_14978,N_14937);
nor UO_1460 (O_1460,N_14887,N_14961);
and UO_1461 (O_1461,N_14879,N_14883);
nor UO_1462 (O_1462,N_14918,N_14905);
xnor UO_1463 (O_1463,N_14917,N_14999);
and UO_1464 (O_1464,N_14925,N_14994);
and UO_1465 (O_1465,N_14995,N_14884);
and UO_1466 (O_1466,N_14952,N_14969);
and UO_1467 (O_1467,N_14972,N_14960);
nand UO_1468 (O_1468,N_14931,N_14966);
xor UO_1469 (O_1469,N_14900,N_14996);
nor UO_1470 (O_1470,N_14916,N_14896);
and UO_1471 (O_1471,N_14932,N_14950);
xor UO_1472 (O_1472,N_14939,N_14999);
or UO_1473 (O_1473,N_14997,N_14969);
nor UO_1474 (O_1474,N_14942,N_14878);
or UO_1475 (O_1475,N_14953,N_14955);
nor UO_1476 (O_1476,N_14991,N_14897);
and UO_1477 (O_1477,N_14962,N_14895);
and UO_1478 (O_1478,N_14994,N_14956);
nand UO_1479 (O_1479,N_14970,N_14923);
and UO_1480 (O_1480,N_14967,N_14997);
nor UO_1481 (O_1481,N_14970,N_14953);
and UO_1482 (O_1482,N_14904,N_14968);
or UO_1483 (O_1483,N_14960,N_14978);
or UO_1484 (O_1484,N_14934,N_14909);
and UO_1485 (O_1485,N_14977,N_14883);
xor UO_1486 (O_1486,N_14952,N_14936);
and UO_1487 (O_1487,N_14895,N_14966);
xnor UO_1488 (O_1488,N_14905,N_14927);
or UO_1489 (O_1489,N_14998,N_14997);
or UO_1490 (O_1490,N_14947,N_14937);
or UO_1491 (O_1491,N_14958,N_14983);
or UO_1492 (O_1492,N_14988,N_14949);
nor UO_1493 (O_1493,N_14892,N_14994);
nor UO_1494 (O_1494,N_14910,N_14969);
xor UO_1495 (O_1495,N_14953,N_14965);
and UO_1496 (O_1496,N_14990,N_14981);
nand UO_1497 (O_1497,N_14971,N_14934);
or UO_1498 (O_1498,N_14951,N_14894);
or UO_1499 (O_1499,N_14990,N_14947);
xnor UO_1500 (O_1500,N_14919,N_14960);
xnor UO_1501 (O_1501,N_14982,N_14917);
nand UO_1502 (O_1502,N_14999,N_14998);
xor UO_1503 (O_1503,N_14895,N_14905);
nor UO_1504 (O_1504,N_14877,N_14947);
xnor UO_1505 (O_1505,N_14900,N_14945);
nor UO_1506 (O_1506,N_14934,N_14921);
nor UO_1507 (O_1507,N_14881,N_14919);
and UO_1508 (O_1508,N_14908,N_14936);
nand UO_1509 (O_1509,N_14905,N_14885);
or UO_1510 (O_1510,N_14887,N_14956);
nor UO_1511 (O_1511,N_14918,N_14913);
and UO_1512 (O_1512,N_14961,N_14904);
xor UO_1513 (O_1513,N_14962,N_14974);
xnor UO_1514 (O_1514,N_14974,N_14913);
or UO_1515 (O_1515,N_14950,N_14896);
or UO_1516 (O_1516,N_14890,N_14957);
xor UO_1517 (O_1517,N_14988,N_14917);
nor UO_1518 (O_1518,N_14969,N_14953);
or UO_1519 (O_1519,N_14954,N_14936);
nand UO_1520 (O_1520,N_14947,N_14993);
nand UO_1521 (O_1521,N_14935,N_14978);
xnor UO_1522 (O_1522,N_14984,N_14881);
nor UO_1523 (O_1523,N_14972,N_14875);
nor UO_1524 (O_1524,N_14982,N_14875);
and UO_1525 (O_1525,N_14923,N_14943);
or UO_1526 (O_1526,N_14882,N_14943);
or UO_1527 (O_1527,N_14993,N_14961);
nor UO_1528 (O_1528,N_14903,N_14918);
xor UO_1529 (O_1529,N_14999,N_14928);
or UO_1530 (O_1530,N_14878,N_14971);
xor UO_1531 (O_1531,N_14918,N_14930);
nor UO_1532 (O_1532,N_14988,N_14905);
xor UO_1533 (O_1533,N_14920,N_14898);
nand UO_1534 (O_1534,N_14990,N_14893);
and UO_1535 (O_1535,N_14978,N_14881);
or UO_1536 (O_1536,N_14999,N_14967);
nand UO_1537 (O_1537,N_14880,N_14932);
and UO_1538 (O_1538,N_14979,N_14936);
or UO_1539 (O_1539,N_14971,N_14997);
or UO_1540 (O_1540,N_14940,N_14951);
nand UO_1541 (O_1541,N_14903,N_14947);
and UO_1542 (O_1542,N_14992,N_14951);
and UO_1543 (O_1543,N_14876,N_14887);
or UO_1544 (O_1544,N_14963,N_14953);
or UO_1545 (O_1545,N_14953,N_14883);
nand UO_1546 (O_1546,N_14936,N_14940);
nor UO_1547 (O_1547,N_14942,N_14978);
nand UO_1548 (O_1548,N_14960,N_14884);
and UO_1549 (O_1549,N_14952,N_14983);
nor UO_1550 (O_1550,N_14955,N_14943);
and UO_1551 (O_1551,N_14901,N_14972);
or UO_1552 (O_1552,N_14909,N_14945);
nor UO_1553 (O_1553,N_14956,N_14933);
or UO_1554 (O_1554,N_14954,N_14915);
and UO_1555 (O_1555,N_14946,N_14959);
and UO_1556 (O_1556,N_14967,N_14893);
or UO_1557 (O_1557,N_14932,N_14882);
or UO_1558 (O_1558,N_14973,N_14999);
nor UO_1559 (O_1559,N_14877,N_14929);
xor UO_1560 (O_1560,N_14912,N_14916);
nand UO_1561 (O_1561,N_14954,N_14993);
and UO_1562 (O_1562,N_14968,N_14996);
nor UO_1563 (O_1563,N_14923,N_14927);
nor UO_1564 (O_1564,N_14986,N_14948);
xnor UO_1565 (O_1565,N_14882,N_14903);
or UO_1566 (O_1566,N_14987,N_14969);
nor UO_1567 (O_1567,N_14899,N_14986);
nor UO_1568 (O_1568,N_14899,N_14949);
nand UO_1569 (O_1569,N_14960,N_14953);
nand UO_1570 (O_1570,N_14880,N_14892);
or UO_1571 (O_1571,N_14951,N_14939);
xor UO_1572 (O_1572,N_14925,N_14910);
nand UO_1573 (O_1573,N_14954,N_14990);
or UO_1574 (O_1574,N_14990,N_14935);
nor UO_1575 (O_1575,N_14904,N_14921);
nor UO_1576 (O_1576,N_14931,N_14953);
and UO_1577 (O_1577,N_14916,N_14892);
nand UO_1578 (O_1578,N_14907,N_14956);
or UO_1579 (O_1579,N_14995,N_14909);
xnor UO_1580 (O_1580,N_14982,N_14983);
xor UO_1581 (O_1581,N_14934,N_14929);
nand UO_1582 (O_1582,N_14937,N_14971);
nand UO_1583 (O_1583,N_14982,N_14994);
or UO_1584 (O_1584,N_14980,N_14898);
and UO_1585 (O_1585,N_14875,N_14955);
nor UO_1586 (O_1586,N_14940,N_14926);
and UO_1587 (O_1587,N_14920,N_14918);
nand UO_1588 (O_1588,N_14943,N_14912);
and UO_1589 (O_1589,N_14936,N_14994);
xnor UO_1590 (O_1590,N_14926,N_14980);
nand UO_1591 (O_1591,N_14988,N_14989);
or UO_1592 (O_1592,N_14970,N_14994);
nand UO_1593 (O_1593,N_14931,N_14963);
or UO_1594 (O_1594,N_14931,N_14901);
xor UO_1595 (O_1595,N_14962,N_14967);
and UO_1596 (O_1596,N_14964,N_14916);
nand UO_1597 (O_1597,N_14964,N_14946);
nand UO_1598 (O_1598,N_14991,N_14995);
or UO_1599 (O_1599,N_14989,N_14981);
or UO_1600 (O_1600,N_14949,N_14950);
xnor UO_1601 (O_1601,N_14927,N_14895);
and UO_1602 (O_1602,N_14916,N_14995);
nor UO_1603 (O_1603,N_14904,N_14909);
xnor UO_1604 (O_1604,N_14968,N_14893);
nand UO_1605 (O_1605,N_14880,N_14943);
or UO_1606 (O_1606,N_14960,N_14879);
xnor UO_1607 (O_1607,N_14908,N_14933);
nand UO_1608 (O_1608,N_14970,N_14887);
nand UO_1609 (O_1609,N_14933,N_14958);
xor UO_1610 (O_1610,N_14945,N_14939);
nor UO_1611 (O_1611,N_14986,N_14920);
and UO_1612 (O_1612,N_14900,N_14974);
nand UO_1613 (O_1613,N_14995,N_14955);
xor UO_1614 (O_1614,N_14992,N_14940);
xnor UO_1615 (O_1615,N_14886,N_14943);
nor UO_1616 (O_1616,N_14909,N_14916);
xnor UO_1617 (O_1617,N_14919,N_14910);
nand UO_1618 (O_1618,N_14974,N_14903);
and UO_1619 (O_1619,N_14988,N_14916);
or UO_1620 (O_1620,N_14941,N_14889);
or UO_1621 (O_1621,N_14981,N_14979);
or UO_1622 (O_1622,N_14968,N_14963);
xor UO_1623 (O_1623,N_14907,N_14940);
nor UO_1624 (O_1624,N_14951,N_14956);
or UO_1625 (O_1625,N_14930,N_14975);
or UO_1626 (O_1626,N_14878,N_14927);
nor UO_1627 (O_1627,N_14948,N_14946);
xnor UO_1628 (O_1628,N_14909,N_14898);
xnor UO_1629 (O_1629,N_14978,N_14959);
nand UO_1630 (O_1630,N_14996,N_14896);
nor UO_1631 (O_1631,N_14974,N_14920);
xor UO_1632 (O_1632,N_14993,N_14884);
xor UO_1633 (O_1633,N_14923,N_14953);
or UO_1634 (O_1634,N_14963,N_14962);
nand UO_1635 (O_1635,N_14935,N_14985);
nor UO_1636 (O_1636,N_14887,N_14945);
nor UO_1637 (O_1637,N_14960,N_14892);
and UO_1638 (O_1638,N_14908,N_14894);
xnor UO_1639 (O_1639,N_14983,N_14878);
xor UO_1640 (O_1640,N_14931,N_14979);
and UO_1641 (O_1641,N_14942,N_14949);
and UO_1642 (O_1642,N_14900,N_14906);
and UO_1643 (O_1643,N_14908,N_14913);
nand UO_1644 (O_1644,N_14985,N_14884);
nand UO_1645 (O_1645,N_14991,N_14947);
nor UO_1646 (O_1646,N_14969,N_14965);
nor UO_1647 (O_1647,N_14962,N_14888);
nor UO_1648 (O_1648,N_14961,N_14935);
nand UO_1649 (O_1649,N_14960,N_14984);
and UO_1650 (O_1650,N_14940,N_14948);
and UO_1651 (O_1651,N_14995,N_14942);
or UO_1652 (O_1652,N_14889,N_14966);
and UO_1653 (O_1653,N_14944,N_14965);
nand UO_1654 (O_1654,N_14937,N_14992);
or UO_1655 (O_1655,N_14969,N_14887);
nor UO_1656 (O_1656,N_14913,N_14919);
and UO_1657 (O_1657,N_14930,N_14994);
or UO_1658 (O_1658,N_14956,N_14965);
and UO_1659 (O_1659,N_14881,N_14885);
xnor UO_1660 (O_1660,N_14889,N_14989);
xnor UO_1661 (O_1661,N_14939,N_14908);
and UO_1662 (O_1662,N_14895,N_14941);
xnor UO_1663 (O_1663,N_14912,N_14910);
and UO_1664 (O_1664,N_14924,N_14960);
nand UO_1665 (O_1665,N_14918,N_14912);
xnor UO_1666 (O_1666,N_14881,N_14992);
or UO_1667 (O_1667,N_14904,N_14963);
nand UO_1668 (O_1668,N_14876,N_14897);
nand UO_1669 (O_1669,N_14935,N_14901);
xnor UO_1670 (O_1670,N_14996,N_14974);
xnor UO_1671 (O_1671,N_14919,N_14980);
and UO_1672 (O_1672,N_14888,N_14957);
or UO_1673 (O_1673,N_14995,N_14917);
nand UO_1674 (O_1674,N_14965,N_14982);
nand UO_1675 (O_1675,N_14993,N_14956);
nor UO_1676 (O_1676,N_14881,N_14944);
nand UO_1677 (O_1677,N_14921,N_14939);
nor UO_1678 (O_1678,N_14997,N_14912);
xor UO_1679 (O_1679,N_14989,N_14961);
nand UO_1680 (O_1680,N_14958,N_14964);
and UO_1681 (O_1681,N_14918,N_14982);
xnor UO_1682 (O_1682,N_14894,N_14889);
and UO_1683 (O_1683,N_14984,N_14931);
or UO_1684 (O_1684,N_14972,N_14985);
nor UO_1685 (O_1685,N_14942,N_14918);
nor UO_1686 (O_1686,N_14924,N_14932);
nand UO_1687 (O_1687,N_14957,N_14983);
xnor UO_1688 (O_1688,N_14933,N_14976);
nand UO_1689 (O_1689,N_14945,N_14977);
nor UO_1690 (O_1690,N_14981,N_14894);
nor UO_1691 (O_1691,N_14964,N_14972);
nand UO_1692 (O_1692,N_14993,N_14918);
xnor UO_1693 (O_1693,N_14984,N_14994);
and UO_1694 (O_1694,N_14889,N_14948);
or UO_1695 (O_1695,N_14899,N_14877);
nor UO_1696 (O_1696,N_14997,N_14918);
nand UO_1697 (O_1697,N_14935,N_14955);
xor UO_1698 (O_1698,N_14924,N_14965);
nand UO_1699 (O_1699,N_14876,N_14991);
nand UO_1700 (O_1700,N_14979,N_14905);
or UO_1701 (O_1701,N_14929,N_14972);
xnor UO_1702 (O_1702,N_14998,N_14981);
or UO_1703 (O_1703,N_14940,N_14962);
or UO_1704 (O_1704,N_14929,N_14975);
xor UO_1705 (O_1705,N_14878,N_14910);
nand UO_1706 (O_1706,N_14928,N_14951);
nor UO_1707 (O_1707,N_14907,N_14914);
nor UO_1708 (O_1708,N_14931,N_14993);
xnor UO_1709 (O_1709,N_14962,N_14991);
or UO_1710 (O_1710,N_14993,N_14999);
xor UO_1711 (O_1711,N_14931,N_14964);
xor UO_1712 (O_1712,N_14919,N_14889);
nand UO_1713 (O_1713,N_14980,N_14941);
nor UO_1714 (O_1714,N_14883,N_14918);
xor UO_1715 (O_1715,N_14938,N_14987);
and UO_1716 (O_1716,N_14975,N_14965);
nor UO_1717 (O_1717,N_14981,N_14898);
nand UO_1718 (O_1718,N_14975,N_14971);
xnor UO_1719 (O_1719,N_14953,N_14934);
nor UO_1720 (O_1720,N_14885,N_14884);
and UO_1721 (O_1721,N_14985,N_14988);
xor UO_1722 (O_1722,N_14983,N_14986);
and UO_1723 (O_1723,N_14917,N_14914);
nand UO_1724 (O_1724,N_14992,N_14968);
or UO_1725 (O_1725,N_14880,N_14969);
and UO_1726 (O_1726,N_14931,N_14978);
and UO_1727 (O_1727,N_14899,N_14893);
and UO_1728 (O_1728,N_14920,N_14932);
or UO_1729 (O_1729,N_14913,N_14903);
and UO_1730 (O_1730,N_14988,N_14961);
nand UO_1731 (O_1731,N_14916,N_14877);
xor UO_1732 (O_1732,N_14979,N_14991);
nor UO_1733 (O_1733,N_14956,N_14935);
nand UO_1734 (O_1734,N_14896,N_14879);
and UO_1735 (O_1735,N_14987,N_14947);
or UO_1736 (O_1736,N_14930,N_14928);
or UO_1737 (O_1737,N_14886,N_14995);
or UO_1738 (O_1738,N_14995,N_14985);
nor UO_1739 (O_1739,N_14960,N_14959);
or UO_1740 (O_1740,N_14925,N_14912);
and UO_1741 (O_1741,N_14996,N_14944);
or UO_1742 (O_1742,N_14998,N_14958);
and UO_1743 (O_1743,N_14956,N_14905);
or UO_1744 (O_1744,N_14960,N_14998);
and UO_1745 (O_1745,N_14964,N_14903);
and UO_1746 (O_1746,N_14901,N_14884);
nor UO_1747 (O_1747,N_14933,N_14879);
and UO_1748 (O_1748,N_14974,N_14904);
and UO_1749 (O_1749,N_14910,N_14913);
nor UO_1750 (O_1750,N_14953,N_14888);
nand UO_1751 (O_1751,N_14880,N_14896);
or UO_1752 (O_1752,N_14974,N_14982);
xor UO_1753 (O_1753,N_14943,N_14899);
nor UO_1754 (O_1754,N_14970,N_14890);
nand UO_1755 (O_1755,N_14975,N_14966);
or UO_1756 (O_1756,N_14969,N_14975);
and UO_1757 (O_1757,N_14928,N_14987);
nor UO_1758 (O_1758,N_14995,N_14970);
or UO_1759 (O_1759,N_14933,N_14959);
or UO_1760 (O_1760,N_14880,N_14875);
or UO_1761 (O_1761,N_14926,N_14942);
nor UO_1762 (O_1762,N_14953,N_14877);
and UO_1763 (O_1763,N_14986,N_14881);
or UO_1764 (O_1764,N_14939,N_14896);
xor UO_1765 (O_1765,N_14913,N_14911);
nor UO_1766 (O_1766,N_14901,N_14887);
and UO_1767 (O_1767,N_14929,N_14915);
or UO_1768 (O_1768,N_14952,N_14887);
nor UO_1769 (O_1769,N_14943,N_14901);
or UO_1770 (O_1770,N_14982,N_14957);
nand UO_1771 (O_1771,N_14893,N_14997);
nand UO_1772 (O_1772,N_14881,N_14888);
nor UO_1773 (O_1773,N_14913,N_14930);
nand UO_1774 (O_1774,N_14991,N_14933);
nand UO_1775 (O_1775,N_14879,N_14988);
and UO_1776 (O_1776,N_14936,N_14978);
or UO_1777 (O_1777,N_14939,N_14974);
nand UO_1778 (O_1778,N_14986,N_14879);
nor UO_1779 (O_1779,N_14942,N_14923);
or UO_1780 (O_1780,N_14992,N_14910);
nor UO_1781 (O_1781,N_14922,N_14923);
nand UO_1782 (O_1782,N_14898,N_14939);
nand UO_1783 (O_1783,N_14966,N_14905);
and UO_1784 (O_1784,N_14876,N_14983);
and UO_1785 (O_1785,N_14999,N_14896);
nor UO_1786 (O_1786,N_14881,N_14918);
and UO_1787 (O_1787,N_14998,N_14890);
or UO_1788 (O_1788,N_14938,N_14885);
nor UO_1789 (O_1789,N_14943,N_14888);
xnor UO_1790 (O_1790,N_14938,N_14954);
or UO_1791 (O_1791,N_14927,N_14978);
xor UO_1792 (O_1792,N_14918,N_14962);
and UO_1793 (O_1793,N_14918,N_14983);
nor UO_1794 (O_1794,N_14890,N_14917);
xnor UO_1795 (O_1795,N_14950,N_14897);
nand UO_1796 (O_1796,N_14880,N_14881);
and UO_1797 (O_1797,N_14956,N_14964);
nand UO_1798 (O_1798,N_14989,N_14912);
xor UO_1799 (O_1799,N_14942,N_14962);
nand UO_1800 (O_1800,N_14923,N_14960);
or UO_1801 (O_1801,N_14881,N_14891);
or UO_1802 (O_1802,N_14968,N_14922);
nand UO_1803 (O_1803,N_14983,N_14951);
nor UO_1804 (O_1804,N_14986,N_14890);
nor UO_1805 (O_1805,N_14880,N_14996);
and UO_1806 (O_1806,N_14900,N_14878);
nor UO_1807 (O_1807,N_14987,N_14916);
nor UO_1808 (O_1808,N_14953,N_14889);
nand UO_1809 (O_1809,N_14914,N_14938);
and UO_1810 (O_1810,N_14936,N_14941);
nor UO_1811 (O_1811,N_14921,N_14940);
or UO_1812 (O_1812,N_14929,N_14993);
or UO_1813 (O_1813,N_14950,N_14915);
xnor UO_1814 (O_1814,N_14875,N_14885);
nor UO_1815 (O_1815,N_14996,N_14972);
nand UO_1816 (O_1816,N_14980,N_14969);
and UO_1817 (O_1817,N_14915,N_14961);
xor UO_1818 (O_1818,N_14962,N_14989);
nor UO_1819 (O_1819,N_14980,N_14916);
nand UO_1820 (O_1820,N_14959,N_14922);
nor UO_1821 (O_1821,N_14930,N_14886);
and UO_1822 (O_1822,N_14884,N_14897);
xnor UO_1823 (O_1823,N_14938,N_14902);
xnor UO_1824 (O_1824,N_14951,N_14968);
and UO_1825 (O_1825,N_14977,N_14984);
and UO_1826 (O_1826,N_14984,N_14938);
nand UO_1827 (O_1827,N_14937,N_14999);
nand UO_1828 (O_1828,N_14952,N_14992);
xor UO_1829 (O_1829,N_14970,N_14986);
or UO_1830 (O_1830,N_14925,N_14898);
nand UO_1831 (O_1831,N_14917,N_14889);
xor UO_1832 (O_1832,N_14936,N_14943);
nor UO_1833 (O_1833,N_14927,N_14947);
or UO_1834 (O_1834,N_14968,N_14984);
nor UO_1835 (O_1835,N_14960,N_14981);
and UO_1836 (O_1836,N_14947,N_14952);
or UO_1837 (O_1837,N_14879,N_14895);
and UO_1838 (O_1838,N_14985,N_14896);
or UO_1839 (O_1839,N_14970,N_14989);
nor UO_1840 (O_1840,N_14994,N_14964);
xor UO_1841 (O_1841,N_14932,N_14893);
xnor UO_1842 (O_1842,N_14885,N_14996);
and UO_1843 (O_1843,N_14892,N_14985);
nor UO_1844 (O_1844,N_14988,N_14976);
nand UO_1845 (O_1845,N_14944,N_14880);
nor UO_1846 (O_1846,N_14940,N_14922);
or UO_1847 (O_1847,N_14943,N_14993);
nor UO_1848 (O_1848,N_14878,N_14894);
nor UO_1849 (O_1849,N_14875,N_14983);
nor UO_1850 (O_1850,N_14896,N_14989);
nor UO_1851 (O_1851,N_14914,N_14959);
or UO_1852 (O_1852,N_14891,N_14896);
nand UO_1853 (O_1853,N_14985,N_14994);
or UO_1854 (O_1854,N_14888,N_14917);
nand UO_1855 (O_1855,N_14930,N_14965);
nor UO_1856 (O_1856,N_14880,N_14913);
and UO_1857 (O_1857,N_14994,N_14893);
xnor UO_1858 (O_1858,N_14926,N_14996);
nand UO_1859 (O_1859,N_14944,N_14930);
and UO_1860 (O_1860,N_14975,N_14896);
and UO_1861 (O_1861,N_14892,N_14937);
or UO_1862 (O_1862,N_14954,N_14882);
nor UO_1863 (O_1863,N_14899,N_14875);
xnor UO_1864 (O_1864,N_14927,N_14910);
and UO_1865 (O_1865,N_14936,N_14976);
nand UO_1866 (O_1866,N_14925,N_14915);
nand UO_1867 (O_1867,N_14947,N_14899);
nor UO_1868 (O_1868,N_14988,N_14919);
nand UO_1869 (O_1869,N_14994,N_14946);
or UO_1870 (O_1870,N_14998,N_14969);
xor UO_1871 (O_1871,N_14925,N_14902);
xor UO_1872 (O_1872,N_14950,N_14999);
nor UO_1873 (O_1873,N_14961,N_14891);
and UO_1874 (O_1874,N_14935,N_14876);
nand UO_1875 (O_1875,N_14993,N_14988);
and UO_1876 (O_1876,N_14888,N_14967);
xnor UO_1877 (O_1877,N_14906,N_14876);
xnor UO_1878 (O_1878,N_14926,N_14928);
or UO_1879 (O_1879,N_14973,N_14908);
xnor UO_1880 (O_1880,N_14887,N_14996);
nor UO_1881 (O_1881,N_14884,N_14955);
or UO_1882 (O_1882,N_14895,N_14939);
nor UO_1883 (O_1883,N_14961,N_14877);
xnor UO_1884 (O_1884,N_14899,N_14929);
or UO_1885 (O_1885,N_14921,N_14946);
nor UO_1886 (O_1886,N_14999,N_14951);
or UO_1887 (O_1887,N_14912,N_14983);
or UO_1888 (O_1888,N_14982,N_14977);
or UO_1889 (O_1889,N_14936,N_14939);
nand UO_1890 (O_1890,N_14898,N_14892);
and UO_1891 (O_1891,N_14879,N_14954);
xnor UO_1892 (O_1892,N_14987,N_14904);
xor UO_1893 (O_1893,N_14919,N_14945);
nor UO_1894 (O_1894,N_14985,N_14930);
nand UO_1895 (O_1895,N_14975,N_14904);
nor UO_1896 (O_1896,N_14975,N_14959);
and UO_1897 (O_1897,N_14962,N_14943);
and UO_1898 (O_1898,N_14956,N_14944);
xor UO_1899 (O_1899,N_14897,N_14875);
xnor UO_1900 (O_1900,N_14922,N_14985);
and UO_1901 (O_1901,N_14934,N_14943);
nor UO_1902 (O_1902,N_14904,N_14941);
nor UO_1903 (O_1903,N_14883,N_14975);
xnor UO_1904 (O_1904,N_14948,N_14899);
nor UO_1905 (O_1905,N_14875,N_14971);
nor UO_1906 (O_1906,N_14886,N_14994);
or UO_1907 (O_1907,N_14922,N_14915);
nor UO_1908 (O_1908,N_14875,N_14929);
nand UO_1909 (O_1909,N_14952,N_14966);
nor UO_1910 (O_1910,N_14945,N_14964);
xor UO_1911 (O_1911,N_14979,N_14983);
nand UO_1912 (O_1912,N_14948,N_14985);
and UO_1913 (O_1913,N_14875,N_14993);
xnor UO_1914 (O_1914,N_14894,N_14949);
nor UO_1915 (O_1915,N_14996,N_14951);
nor UO_1916 (O_1916,N_14890,N_14980);
xnor UO_1917 (O_1917,N_14917,N_14904);
or UO_1918 (O_1918,N_14981,N_14952);
nor UO_1919 (O_1919,N_14917,N_14947);
or UO_1920 (O_1920,N_14999,N_14946);
or UO_1921 (O_1921,N_14933,N_14904);
and UO_1922 (O_1922,N_14876,N_14999);
and UO_1923 (O_1923,N_14897,N_14962);
nand UO_1924 (O_1924,N_14900,N_14939);
nand UO_1925 (O_1925,N_14905,N_14924);
and UO_1926 (O_1926,N_14896,N_14925);
nand UO_1927 (O_1927,N_14946,N_14924);
xnor UO_1928 (O_1928,N_14951,N_14888);
xor UO_1929 (O_1929,N_14958,N_14984);
or UO_1930 (O_1930,N_14911,N_14985);
nand UO_1931 (O_1931,N_14900,N_14877);
nand UO_1932 (O_1932,N_14973,N_14967);
nand UO_1933 (O_1933,N_14913,N_14916);
nand UO_1934 (O_1934,N_14935,N_14965);
or UO_1935 (O_1935,N_14908,N_14930);
and UO_1936 (O_1936,N_14949,N_14999);
and UO_1937 (O_1937,N_14961,N_14897);
and UO_1938 (O_1938,N_14880,N_14891);
nand UO_1939 (O_1939,N_14927,N_14926);
and UO_1940 (O_1940,N_14923,N_14885);
nor UO_1941 (O_1941,N_14876,N_14990);
nor UO_1942 (O_1942,N_14902,N_14958);
nand UO_1943 (O_1943,N_14987,N_14963);
and UO_1944 (O_1944,N_14929,N_14887);
or UO_1945 (O_1945,N_14884,N_14919);
or UO_1946 (O_1946,N_14971,N_14992);
or UO_1947 (O_1947,N_14941,N_14940);
nand UO_1948 (O_1948,N_14901,N_14980);
nand UO_1949 (O_1949,N_14895,N_14902);
nor UO_1950 (O_1950,N_14923,N_14951);
nand UO_1951 (O_1951,N_14997,N_14876);
and UO_1952 (O_1952,N_14939,N_14894);
nor UO_1953 (O_1953,N_14926,N_14979);
nor UO_1954 (O_1954,N_14969,N_14946);
and UO_1955 (O_1955,N_14993,N_14960);
and UO_1956 (O_1956,N_14998,N_14903);
nand UO_1957 (O_1957,N_14923,N_14961);
nor UO_1958 (O_1958,N_14922,N_14966);
xnor UO_1959 (O_1959,N_14941,N_14896);
nand UO_1960 (O_1960,N_14956,N_14875);
nor UO_1961 (O_1961,N_14965,N_14950);
xor UO_1962 (O_1962,N_14983,N_14907);
or UO_1963 (O_1963,N_14927,N_14996);
and UO_1964 (O_1964,N_14981,N_14936);
nand UO_1965 (O_1965,N_14922,N_14986);
and UO_1966 (O_1966,N_14908,N_14970);
and UO_1967 (O_1967,N_14998,N_14938);
nor UO_1968 (O_1968,N_14956,N_14878);
or UO_1969 (O_1969,N_14946,N_14929);
nand UO_1970 (O_1970,N_14886,N_14902);
nand UO_1971 (O_1971,N_14887,N_14934);
and UO_1972 (O_1972,N_14906,N_14975);
and UO_1973 (O_1973,N_14997,N_14963);
and UO_1974 (O_1974,N_14972,N_14913);
or UO_1975 (O_1975,N_14991,N_14904);
or UO_1976 (O_1976,N_14894,N_14918);
nand UO_1977 (O_1977,N_14931,N_14960);
and UO_1978 (O_1978,N_14940,N_14930);
or UO_1979 (O_1979,N_14924,N_14968);
nor UO_1980 (O_1980,N_14975,N_14885);
nor UO_1981 (O_1981,N_14920,N_14995);
nand UO_1982 (O_1982,N_14929,N_14960);
and UO_1983 (O_1983,N_14939,N_14989);
nor UO_1984 (O_1984,N_14878,N_14969);
nand UO_1985 (O_1985,N_14900,N_14897);
or UO_1986 (O_1986,N_14976,N_14926);
nor UO_1987 (O_1987,N_14931,N_14973);
nor UO_1988 (O_1988,N_14956,N_14986);
nand UO_1989 (O_1989,N_14949,N_14877);
and UO_1990 (O_1990,N_14961,N_14978);
nor UO_1991 (O_1991,N_14895,N_14896);
xor UO_1992 (O_1992,N_14972,N_14937);
and UO_1993 (O_1993,N_14925,N_14947);
or UO_1994 (O_1994,N_14940,N_14967);
and UO_1995 (O_1995,N_14885,N_14964);
or UO_1996 (O_1996,N_14931,N_14926);
or UO_1997 (O_1997,N_14969,N_14877);
and UO_1998 (O_1998,N_14915,N_14953);
nor UO_1999 (O_1999,N_14920,N_14935);
endmodule