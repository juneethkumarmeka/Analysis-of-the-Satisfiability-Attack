module basic_1000_10000_1500_5_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_253,In_543);
nand U1 (N_1,In_73,In_259);
and U2 (N_2,In_148,In_539);
nand U3 (N_3,In_561,In_646);
and U4 (N_4,In_940,In_87);
nand U5 (N_5,In_487,In_584);
nand U6 (N_6,In_521,In_637);
nor U7 (N_7,In_121,In_753);
nor U8 (N_8,In_633,In_871);
nand U9 (N_9,In_306,In_271);
and U10 (N_10,In_309,In_188);
or U11 (N_11,In_298,In_251);
or U12 (N_12,In_33,In_609);
nor U13 (N_13,In_716,In_709);
nor U14 (N_14,In_685,In_975);
nor U15 (N_15,In_836,In_173);
nor U16 (N_16,In_913,In_14);
or U17 (N_17,In_9,In_725);
and U18 (N_18,In_761,In_311);
nand U19 (N_19,In_332,In_362);
and U20 (N_20,In_981,In_401);
nand U21 (N_21,In_420,In_974);
or U22 (N_22,In_195,In_741);
xor U23 (N_23,In_484,In_961);
or U24 (N_24,In_270,In_428);
and U25 (N_25,In_766,In_81);
nand U26 (N_26,In_804,In_547);
and U27 (N_27,In_27,In_25);
nor U28 (N_28,In_814,In_673);
nor U29 (N_29,In_582,In_792);
or U30 (N_30,In_107,In_509);
nor U31 (N_31,In_468,In_1);
or U32 (N_32,In_357,In_337);
nor U33 (N_33,In_34,In_686);
or U34 (N_34,In_751,In_890);
and U35 (N_35,In_876,In_129);
nand U36 (N_36,In_954,In_841);
and U37 (N_37,In_677,In_506);
and U38 (N_38,In_808,In_229);
or U39 (N_39,In_134,In_736);
and U40 (N_40,In_347,In_647);
nor U41 (N_41,In_3,In_218);
nand U42 (N_42,In_381,In_409);
or U43 (N_43,In_755,In_331);
or U44 (N_44,In_432,In_608);
nor U45 (N_45,In_15,In_921);
nor U46 (N_46,In_439,In_953);
or U47 (N_47,In_930,In_241);
and U48 (N_48,In_386,In_247);
or U49 (N_49,In_597,In_292);
and U50 (N_50,In_127,In_430);
nand U51 (N_51,In_210,In_705);
or U52 (N_52,In_457,In_977);
or U53 (N_53,In_242,In_211);
and U54 (N_54,In_344,In_986);
or U55 (N_55,In_451,In_626);
nor U56 (N_56,In_462,In_289);
and U57 (N_57,In_868,In_290);
or U58 (N_58,In_361,In_589);
nand U59 (N_59,In_693,In_248);
or U60 (N_60,In_689,In_743);
nor U61 (N_61,In_510,In_485);
nor U62 (N_62,In_669,In_861);
nand U63 (N_63,In_398,In_67);
nor U64 (N_64,In_959,In_200);
or U65 (N_65,In_98,In_583);
and U66 (N_66,In_748,In_826);
and U67 (N_67,In_21,In_789);
nor U68 (N_68,In_72,In_448);
nand U69 (N_69,In_447,In_778);
nand U70 (N_70,In_989,In_313);
or U71 (N_71,In_117,In_84);
nor U72 (N_72,In_275,In_927);
or U73 (N_73,In_681,In_197);
and U74 (N_74,In_214,In_215);
or U75 (N_75,In_631,In_412);
nand U76 (N_76,In_665,In_153);
nor U77 (N_77,In_246,In_122);
nor U78 (N_78,In_407,In_380);
and U79 (N_79,In_904,In_972);
and U80 (N_80,In_834,In_529);
nor U81 (N_81,In_45,In_138);
nand U82 (N_82,In_657,In_243);
nand U83 (N_83,In_666,In_415);
and U84 (N_84,In_262,In_221);
nand U85 (N_85,In_823,In_226);
nor U86 (N_86,In_49,In_966);
nor U87 (N_87,In_302,In_334);
nand U88 (N_88,In_548,In_264);
nand U89 (N_89,In_391,In_674);
or U90 (N_90,In_797,In_827);
and U91 (N_91,In_592,In_653);
or U92 (N_92,In_739,In_844);
or U93 (N_93,In_18,In_553);
and U94 (N_94,In_329,In_463);
and U95 (N_95,In_414,In_902);
nand U96 (N_96,In_581,In_704);
nor U97 (N_97,In_518,In_175);
or U98 (N_98,In_212,In_41);
and U99 (N_99,In_923,In_907);
or U100 (N_100,In_857,In_364);
or U101 (N_101,In_874,In_824);
nand U102 (N_102,In_503,In_520);
nand U103 (N_103,In_13,In_256);
and U104 (N_104,In_860,In_898);
nand U105 (N_105,In_452,In_55);
nor U106 (N_106,In_103,In_632);
or U107 (N_107,In_239,In_108);
nand U108 (N_108,In_57,In_760);
or U109 (N_109,In_537,In_99);
or U110 (N_110,In_472,In_842);
and U111 (N_111,In_651,In_796);
nand U112 (N_112,In_636,In_956);
and U113 (N_113,In_356,In_11);
nand U114 (N_114,In_206,In_908);
nand U115 (N_115,In_723,In_943);
and U116 (N_116,In_979,In_312);
nand U117 (N_117,In_319,In_812);
nor U118 (N_118,In_737,In_277);
nor U119 (N_119,In_567,In_119);
nand U120 (N_120,In_38,In_531);
or U121 (N_121,In_629,In_238);
nor U122 (N_122,In_562,In_590);
nand U123 (N_123,In_28,In_746);
nand U124 (N_124,In_763,In_697);
and U125 (N_125,In_997,In_130);
or U126 (N_126,In_110,In_217);
and U127 (N_127,In_0,In_397);
or U128 (N_128,In_799,In_282);
nand U129 (N_129,In_726,In_151);
and U130 (N_130,In_433,In_516);
nor U131 (N_131,In_599,In_640);
and U132 (N_132,In_528,In_578);
nor U133 (N_133,In_170,In_479);
nand U134 (N_134,In_152,In_111);
nor U135 (N_135,In_490,In_780);
or U136 (N_136,In_384,In_639);
or U137 (N_137,In_51,In_32);
nand U138 (N_138,In_141,In_707);
or U139 (N_139,In_189,In_106);
and U140 (N_140,In_931,In_910);
nor U141 (N_141,In_996,In_788);
nor U142 (N_142,In_534,In_877);
and U143 (N_143,In_690,In_892);
nor U144 (N_144,In_621,In_196);
nor U145 (N_145,In_867,In_245);
and U146 (N_146,In_475,In_37);
nor U147 (N_147,In_586,In_885);
and U148 (N_148,In_752,In_419);
and U149 (N_149,In_848,In_889);
or U150 (N_150,In_557,In_157);
nor U151 (N_151,In_533,In_555);
or U152 (N_152,In_502,In_566);
and U153 (N_153,In_610,In_375);
nand U154 (N_154,In_692,In_900);
or U155 (N_155,In_650,In_496);
and U156 (N_156,In_740,In_678);
nor U157 (N_157,In_444,In_434);
nor U158 (N_158,In_64,In_388);
and U159 (N_159,In_299,In_688);
nor U160 (N_160,In_287,In_494);
nor U161 (N_161,In_321,In_711);
nand U162 (N_162,In_389,In_135);
and U163 (N_163,In_802,In_425);
nand U164 (N_164,In_155,In_83);
and U165 (N_165,In_483,In_635);
nand U166 (N_166,In_209,In_658);
or U167 (N_167,In_851,In_4);
nor U168 (N_168,In_782,In_437);
nor U169 (N_169,In_58,In_252);
and U170 (N_170,In_205,In_202);
nand U171 (N_171,In_71,In_887);
nand U172 (N_172,In_875,In_465);
nand U173 (N_173,In_895,In_617);
nor U174 (N_174,In_638,In_995);
and U175 (N_175,In_883,In_42);
and U176 (N_176,In_288,In_661);
nor U177 (N_177,In_317,In_225);
nor U178 (N_178,In_770,In_449);
and U179 (N_179,In_982,In_351);
and U180 (N_180,In_594,In_527);
nand U181 (N_181,In_493,In_233);
nor U182 (N_182,In_691,In_560);
nor U183 (N_183,In_291,In_140);
or U184 (N_184,In_395,In_336);
and U185 (N_185,In_934,In_749);
nor U186 (N_186,In_142,In_227);
or U187 (N_187,In_858,In_694);
and U188 (N_188,In_964,In_787);
nor U189 (N_189,In_345,In_145);
nor U190 (N_190,In_61,In_575);
and U191 (N_191,In_837,In_216);
or U192 (N_192,In_869,In_684);
nor U193 (N_193,In_456,In_91);
nand U194 (N_194,In_474,In_240);
or U195 (N_195,In_777,In_269);
nand U196 (N_196,In_757,In_295);
or U197 (N_197,In_879,In_286);
or U198 (N_198,In_112,In_652);
nand U199 (N_199,In_564,In_458);
nor U200 (N_200,In_68,In_840);
nand U201 (N_201,In_261,In_565);
nor U202 (N_202,In_466,In_664);
or U203 (N_203,In_471,In_146);
nand U204 (N_204,In_497,In_498);
nor U205 (N_205,In_76,In_2);
and U206 (N_206,In_893,In_349);
and U207 (N_207,In_236,In_371);
and U208 (N_208,In_769,In_358);
or U209 (N_209,In_19,In_230);
and U210 (N_210,In_634,In_192);
and U211 (N_211,In_849,In_396);
and U212 (N_212,In_476,In_399);
or U213 (N_213,In_62,In_687);
nand U214 (N_214,In_624,In_160);
and U215 (N_215,In_696,In_801);
or U216 (N_216,In_36,In_459);
nand U217 (N_217,In_998,In_17);
and U218 (N_218,In_266,In_143);
or U219 (N_219,In_411,In_701);
and U220 (N_220,In_779,In_720);
or U221 (N_221,In_668,In_558);
nand U222 (N_222,In_862,In_622);
nand U223 (N_223,In_194,In_949);
nand U224 (N_224,In_759,In_204);
nand U225 (N_225,In_526,In_50);
nor U226 (N_226,In_971,In_601);
nor U227 (N_227,In_273,In_5);
and U228 (N_228,In_393,In_817);
nor U229 (N_229,In_523,In_208);
and U230 (N_230,In_220,In_545);
nand U231 (N_231,In_815,In_552);
and U232 (N_232,In_951,In_181);
or U233 (N_233,In_785,In_939);
nand U234 (N_234,In_481,In_810);
nand U235 (N_235,In_265,In_501);
and U236 (N_236,In_672,In_655);
and U237 (N_237,In_405,In_825);
and U238 (N_238,In_944,In_920);
or U239 (N_239,In_762,In_846);
or U240 (N_240,In_783,In_864);
and U241 (N_241,In_570,In_571);
and U242 (N_242,In_427,In_508);
or U243 (N_243,In_641,In_343);
nor U244 (N_244,In_917,In_147);
nor U245 (N_245,In_764,In_137);
or U246 (N_246,In_89,In_870);
and U247 (N_247,In_69,In_886);
and U248 (N_248,In_219,In_372);
and U249 (N_249,In_104,In_85);
nand U250 (N_250,In_832,In_424);
and U251 (N_251,In_422,In_161);
nand U252 (N_252,In_267,In_207);
or U253 (N_253,In_616,In_314);
and U254 (N_254,In_663,In_65);
nand U255 (N_255,In_660,In_576);
or U256 (N_256,In_588,In_254);
or U257 (N_257,In_721,In_714);
and U258 (N_258,In_52,In_791);
or U259 (N_259,In_550,In_744);
or U260 (N_260,In_307,In_625);
or U261 (N_261,In_324,In_78);
or U262 (N_262,In_232,In_504);
nand U263 (N_263,In_203,In_719);
nand U264 (N_264,In_962,In_790);
nor U265 (N_265,In_198,In_530);
or U266 (N_266,In_854,In_183);
and U267 (N_267,In_618,In_228);
nand U268 (N_268,In_549,In_492);
nor U269 (N_269,In_320,In_56);
or U270 (N_270,In_43,In_585);
nor U271 (N_271,In_572,In_352);
nor U272 (N_272,In_710,In_470);
and U273 (N_273,In_340,In_35);
nand U274 (N_274,In_469,In_237);
and U275 (N_275,In_999,In_990);
or U276 (N_276,In_360,In_738);
nor U277 (N_277,In_105,In_654);
nor U278 (N_278,In_699,In_569);
nand U279 (N_279,In_53,In_850);
or U280 (N_280,In_554,In_477);
or U281 (N_281,In_40,In_540);
nor U282 (N_282,In_855,In_813);
and U283 (N_283,In_775,In_774);
or U284 (N_284,In_191,In_342);
nor U285 (N_285,In_919,In_70);
nand U286 (N_286,In_519,In_906);
nand U287 (N_287,In_922,In_577);
or U288 (N_288,In_281,In_423);
nand U289 (N_289,In_376,In_359);
or U290 (N_290,In_991,In_676);
or U291 (N_291,In_865,In_538);
xnor U292 (N_292,In_274,In_614);
or U293 (N_293,In_95,In_31);
and U294 (N_294,In_436,In_128);
or U295 (N_295,In_830,In_645);
or U296 (N_296,In_662,In_441);
nor U297 (N_297,In_912,In_819);
and U298 (N_298,In_733,In_952);
nand U299 (N_299,In_184,In_888);
and U300 (N_300,In_994,In_149);
nor U301 (N_301,In_522,In_960);
nand U302 (N_302,In_708,In_325);
nor U303 (N_303,In_901,In_10);
and U304 (N_304,In_935,In_715);
and U305 (N_305,In_628,In_820);
or U306 (N_306,In_406,In_48);
or U307 (N_307,In_491,In_185);
or U308 (N_308,In_285,In_426);
nand U309 (N_309,In_899,In_947);
xor U310 (N_310,In_682,In_937);
nand U311 (N_311,In_330,In_294);
nand U312 (N_312,In_698,In_392);
and U313 (N_313,In_440,In_683);
and U314 (N_314,In_310,In_988);
nand U315 (N_315,In_679,In_442);
or U316 (N_316,In_500,In_524);
or U317 (N_317,In_374,In_542);
nor U318 (N_318,In_993,In_59);
and U319 (N_319,In_656,In_158);
nand U320 (N_320,In_431,In_911);
and U321 (N_321,In_171,In_963);
and U322 (N_322,In_421,In_366);
and U323 (N_323,In_495,In_443);
and U324 (N_324,In_353,In_283);
nand U325 (N_325,In_144,In_512);
nor U326 (N_326,In_563,In_354);
nand U327 (N_327,In_47,In_26);
and U328 (N_328,In_505,In_296);
or U329 (N_329,In_118,In_318);
and U330 (N_330,In_732,In_132);
nand U331 (N_331,In_909,In_776);
and U332 (N_332,In_260,In_168);
nor U333 (N_333,In_323,In_24);
nand U334 (N_334,In_297,In_120);
or U335 (N_335,In_446,In_74);
nand U336 (N_336,In_435,In_793);
nor U337 (N_337,In_822,In_809);
or U338 (N_338,In_728,In_880);
nor U339 (N_339,In_124,In_773);
nor U340 (N_340,In_918,In_852);
nand U341 (N_341,In_976,In_544);
and U342 (N_342,In_123,In_182);
and U343 (N_343,In_619,In_671);
nand U344 (N_344,In_758,In_786);
and U345 (N_345,In_600,In_604);
and U346 (N_346,In_373,In_587);
or U347 (N_347,In_328,In_418);
or U348 (N_348,In_897,In_455);
nor U349 (N_349,In_172,In_659);
nand U350 (N_350,In_536,In_190);
nor U351 (N_351,In_978,In_623);
or U352 (N_352,In_100,In_385);
nand U353 (N_353,In_873,In_402);
nand U354 (N_354,In_174,In_845);
and U355 (N_355,In_713,In_514);
and U356 (N_356,In_928,In_747);
nor U357 (N_357,In_593,In_598);
and U358 (N_358,In_79,In_113);
nor U359 (N_359,In_224,In_821);
nand U360 (N_360,In_304,In_131);
nor U361 (N_361,In_387,In_882);
or U362 (N_362,In_416,In_630);
and U363 (N_363,In_163,In_369);
nand U364 (N_364,In_517,In_515);
nor U365 (N_365,In_765,In_80);
nand U366 (N_366,In_66,In_829);
and U367 (N_367,In_811,In_133);
xor U368 (N_368,In_44,In_367);
nand U369 (N_369,In_46,In_63);
and U370 (N_370,In_379,In_363);
nor U371 (N_371,In_109,In_333);
or U372 (N_372,In_675,In_938);
nor U373 (N_373,In_750,In_16);
nand U374 (N_374,In_835,In_370);
or U375 (N_375,In_250,In_278);
and U376 (N_376,In_905,In_644);
nor U377 (N_377,In_284,In_335);
nand U378 (N_378,In_394,In_933);
nand U379 (N_379,In_805,In_97);
nor U380 (N_380,In_159,In_177);
nor U381 (N_381,In_568,In_305);
nor U382 (N_382,In_8,In_950);
nor U383 (N_383,In_754,In_847);
nand U384 (N_384,In_595,In_818);
nor U385 (N_385,In_532,In_383);
nand U386 (N_386,In_965,In_856);
xnor U387 (N_387,In_473,In_772);
nor U388 (N_388,In_438,In_176);
and U389 (N_389,In_169,In_948);
or U390 (N_390,In_178,In_591);
or U391 (N_391,In_390,In_489);
or U392 (N_392,In_162,In_115);
nand U393 (N_393,In_116,In_573);
and U394 (N_394,In_139,In_878);
and U395 (N_395,In_718,In_30);
nand U396 (N_396,In_165,In_445);
and U397 (N_397,In_724,In_125);
or U398 (N_398,In_90,In_894);
and U399 (N_399,In_39,In_382);
and U400 (N_400,In_969,In_803);
and U401 (N_401,In_613,In_955);
or U402 (N_402,In_199,In_186);
or U403 (N_403,In_179,In_92);
nand U404 (N_404,In_244,In_722);
nor U405 (N_405,In_326,In_499);
nor U406 (N_406,In_756,In_695);
nor U407 (N_407,In_461,In_642);
nand U408 (N_408,In_20,In_798);
and U409 (N_409,In_136,In_315);
and U410 (N_410,In_350,In_417);
nand U411 (N_411,In_667,In_800);
nor U412 (N_412,In_745,In_486);
nor U413 (N_413,In_932,In_670);
nand U414 (N_414,In_859,In_513);
or U415 (N_415,In_276,In_453);
nor U416 (N_416,In_559,In_903);
nand U417 (N_417,In_941,In_82);
xor U418 (N_418,In_23,In_413);
and U419 (N_419,In_712,In_828);
or U420 (N_420,In_702,In_967);
nor U421 (N_421,In_863,In_968);
or U422 (N_422,In_156,In_987);
and U423 (N_423,In_88,In_742);
nor U424 (N_424,In_126,In_958);
and U425 (N_425,In_884,In_403);
xor U426 (N_426,In_460,In_93);
or U427 (N_427,In_213,In_408);
and U428 (N_428,In_308,In_322);
nand U429 (N_429,In_794,In_925);
nand U430 (N_430,In_896,In_75);
or U431 (N_431,In_551,In_327);
nor U432 (N_432,In_627,In_546);
nor U433 (N_433,In_257,In_488);
nand U434 (N_434,In_280,In_164);
and U435 (N_435,In_154,In_293);
and U436 (N_436,In_480,In_467);
or U437 (N_437,In_22,In_201);
nor U438 (N_438,In_429,In_535);
nand U439 (N_439,In_450,In_365);
nor U440 (N_440,In_872,In_339);
nor U441 (N_441,In_839,In_580);
and U442 (N_442,In_234,In_101);
and U443 (N_443,In_924,In_942);
and U444 (N_444,In_404,In_180);
or U445 (N_445,In_222,In_649);
nor U446 (N_446,In_464,In_94);
or U447 (N_447,In_936,In_231);
or U448 (N_448,In_378,In_96);
nand U449 (N_449,In_612,In_914);
or U450 (N_450,In_316,In_574);
nand U451 (N_451,In_301,In_258);
or U452 (N_452,In_77,In_482);
and U453 (N_453,In_511,In_970);
and U454 (N_454,In_735,In_167);
nand U455 (N_455,In_926,In_60);
and U456 (N_456,In_929,In_605);
or U457 (N_457,In_806,In_731);
and U458 (N_458,In_303,In_946);
and U459 (N_459,In_957,In_984);
or U460 (N_460,In_166,In_346);
or U461 (N_461,In_992,In_341);
or U462 (N_462,In_150,In_915);
nor U463 (N_463,In_368,In_235);
nor U464 (N_464,In_54,In_717);
or U465 (N_465,In_29,In_795);
or U466 (N_466,In_525,In_843);
or U467 (N_467,In_541,In_703);
nor U468 (N_468,In_891,In_838);
nand U469 (N_469,In_973,In_853);
or U470 (N_470,In_833,In_86);
nand U471 (N_471,In_507,In_377);
and U472 (N_472,In_983,In_729);
nand U473 (N_473,In_980,In_249);
nor U474 (N_474,In_187,In_781);
nand U475 (N_475,In_866,In_596);
or U476 (N_476,In_400,In_771);
and U477 (N_477,In_784,In_615);
or U478 (N_478,In_881,In_102);
or U479 (N_479,In_348,In_602);
nand U480 (N_480,In_700,In_7);
nor U481 (N_481,In_985,In_831);
and U482 (N_482,In_454,In_730);
nor U483 (N_483,In_648,In_611);
or U484 (N_484,In_706,In_255);
nor U485 (N_485,In_6,In_556);
or U486 (N_486,In_807,In_410);
nor U487 (N_487,In_223,In_355);
or U488 (N_488,In_268,In_579);
nor U489 (N_489,In_114,In_767);
nor U490 (N_490,In_916,In_620);
and U491 (N_491,In_193,In_643);
nor U492 (N_492,In_734,In_680);
nand U493 (N_493,In_606,In_272);
nand U494 (N_494,In_945,In_300);
and U495 (N_495,In_603,In_768);
nor U496 (N_496,In_478,In_263);
and U497 (N_497,In_279,In_727);
or U498 (N_498,In_12,In_816);
nand U499 (N_499,In_338,In_607);
nor U500 (N_500,In_459,In_520);
nor U501 (N_501,In_251,In_702);
or U502 (N_502,In_607,In_251);
and U503 (N_503,In_162,In_445);
nor U504 (N_504,In_611,In_345);
or U505 (N_505,In_983,In_406);
nor U506 (N_506,In_162,In_572);
and U507 (N_507,In_19,In_110);
or U508 (N_508,In_929,In_749);
or U509 (N_509,In_937,In_959);
or U510 (N_510,In_239,In_741);
or U511 (N_511,In_536,In_234);
or U512 (N_512,In_247,In_717);
and U513 (N_513,In_286,In_889);
nor U514 (N_514,In_798,In_577);
nor U515 (N_515,In_627,In_46);
and U516 (N_516,In_232,In_702);
or U517 (N_517,In_464,In_929);
nor U518 (N_518,In_729,In_413);
and U519 (N_519,In_830,In_680);
and U520 (N_520,In_550,In_355);
or U521 (N_521,In_945,In_555);
or U522 (N_522,In_227,In_260);
and U523 (N_523,In_340,In_77);
nor U524 (N_524,In_544,In_683);
and U525 (N_525,In_30,In_737);
and U526 (N_526,In_644,In_901);
or U527 (N_527,In_603,In_289);
nand U528 (N_528,In_16,In_273);
nand U529 (N_529,In_478,In_936);
or U530 (N_530,In_765,In_968);
nor U531 (N_531,In_122,In_158);
and U532 (N_532,In_670,In_205);
nor U533 (N_533,In_391,In_817);
nor U534 (N_534,In_320,In_347);
nand U535 (N_535,In_766,In_912);
and U536 (N_536,In_965,In_911);
and U537 (N_537,In_696,In_704);
nand U538 (N_538,In_558,In_410);
or U539 (N_539,In_427,In_748);
or U540 (N_540,In_825,In_74);
xor U541 (N_541,In_496,In_306);
or U542 (N_542,In_529,In_569);
and U543 (N_543,In_87,In_72);
nor U544 (N_544,In_547,In_28);
nor U545 (N_545,In_665,In_159);
or U546 (N_546,In_781,In_659);
or U547 (N_547,In_491,In_12);
and U548 (N_548,In_133,In_599);
and U549 (N_549,In_882,In_29);
or U550 (N_550,In_735,In_609);
or U551 (N_551,In_751,In_395);
and U552 (N_552,In_527,In_294);
or U553 (N_553,In_653,In_42);
nor U554 (N_554,In_204,In_862);
nor U555 (N_555,In_669,In_101);
nor U556 (N_556,In_780,In_655);
and U557 (N_557,In_169,In_328);
nand U558 (N_558,In_426,In_819);
nor U559 (N_559,In_739,In_113);
nand U560 (N_560,In_10,In_214);
or U561 (N_561,In_520,In_731);
nand U562 (N_562,In_879,In_902);
nor U563 (N_563,In_533,In_746);
and U564 (N_564,In_529,In_182);
nor U565 (N_565,In_247,In_553);
and U566 (N_566,In_547,In_723);
nand U567 (N_567,In_961,In_886);
or U568 (N_568,In_416,In_253);
nand U569 (N_569,In_484,In_114);
nor U570 (N_570,In_458,In_596);
nand U571 (N_571,In_492,In_20);
or U572 (N_572,In_957,In_499);
or U573 (N_573,In_242,In_290);
nor U574 (N_574,In_853,In_29);
or U575 (N_575,In_363,In_176);
and U576 (N_576,In_782,In_467);
nand U577 (N_577,In_577,In_113);
or U578 (N_578,In_433,In_200);
nor U579 (N_579,In_294,In_836);
or U580 (N_580,In_83,In_720);
and U581 (N_581,In_233,In_819);
nor U582 (N_582,In_821,In_581);
nor U583 (N_583,In_344,In_912);
nand U584 (N_584,In_589,In_776);
or U585 (N_585,In_419,In_84);
nand U586 (N_586,In_740,In_725);
nand U587 (N_587,In_73,In_301);
and U588 (N_588,In_810,In_764);
or U589 (N_589,In_432,In_453);
or U590 (N_590,In_390,In_554);
nand U591 (N_591,In_447,In_597);
nor U592 (N_592,In_191,In_900);
or U593 (N_593,In_851,In_371);
or U594 (N_594,In_534,In_828);
nor U595 (N_595,In_39,In_673);
nand U596 (N_596,In_829,In_195);
and U597 (N_597,In_230,In_68);
nand U598 (N_598,In_642,In_309);
and U599 (N_599,In_457,In_369);
or U600 (N_600,In_872,In_184);
nand U601 (N_601,In_808,In_299);
and U602 (N_602,In_608,In_531);
nor U603 (N_603,In_315,In_258);
nor U604 (N_604,In_817,In_512);
nand U605 (N_605,In_203,In_535);
nand U606 (N_606,In_654,In_79);
nor U607 (N_607,In_271,In_54);
or U608 (N_608,In_710,In_567);
or U609 (N_609,In_313,In_575);
nand U610 (N_610,In_348,In_372);
or U611 (N_611,In_602,In_998);
or U612 (N_612,In_453,In_614);
and U613 (N_613,In_637,In_233);
or U614 (N_614,In_766,In_955);
or U615 (N_615,In_195,In_132);
nand U616 (N_616,In_177,In_513);
nor U617 (N_617,In_359,In_63);
nor U618 (N_618,In_203,In_692);
nor U619 (N_619,In_942,In_934);
and U620 (N_620,In_544,In_196);
and U621 (N_621,In_798,In_386);
nor U622 (N_622,In_800,In_354);
and U623 (N_623,In_65,In_484);
and U624 (N_624,In_950,In_961);
and U625 (N_625,In_254,In_208);
nand U626 (N_626,In_594,In_76);
and U627 (N_627,In_807,In_558);
nand U628 (N_628,In_686,In_599);
or U629 (N_629,In_208,In_911);
nand U630 (N_630,In_702,In_706);
or U631 (N_631,In_996,In_979);
nor U632 (N_632,In_941,In_587);
nor U633 (N_633,In_304,In_178);
or U634 (N_634,In_307,In_299);
nor U635 (N_635,In_630,In_775);
or U636 (N_636,In_371,In_327);
or U637 (N_637,In_426,In_187);
and U638 (N_638,In_338,In_832);
and U639 (N_639,In_411,In_151);
nor U640 (N_640,In_117,In_816);
nand U641 (N_641,In_368,In_690);
or U642 (N_642,In_496,In_90);
nor U643 (N_643,In_319,In_116);
nor U644 (N_644,In_660,In_264);
or U645 (N_645,In_622,In_929);
nor U646 (N_646,In_660,In_23);
or U647 (N_647,In_146,In_560);
nor U648 (N_648,In_106,In_575);
or U649 (N_649,In_487,In_796);
or U650 (N_650,In_406,In_550);
or U651 (N_651,In_664,In_580);
and U652 (N_652,In_844,In_862);
and U653 (N_653,In_791,In_474);
or U654 (N_654,In_375,In_418);
nor U655 (N_655,In_298,In_518);
or U656 (N_656,In_359,In_33);
and U657 (N_657,In_219,In_825);
or U658 (N_658,In_518,In_160);
nor U659 (N_659,In_57,In_252);
nor U660 (N_660,In_955,In_458);
nand U661 (N_661,In_902,In_225);
and U662 (N_662,In_189,In_958);
nand U663 (N_663,In_42,In_251);
and U664 (N_664,In_990,In_12);
nand U665 (N_665,In_317,In_562);
nor U666 (N_666,In_148,In_365);
nand U667 (N_667,In_331,In_857);
nand U668 (N_668,In_420,In_565);
nor U669 (N_669,In_168,In_240);
and U670 (N_670,In_602,In_242);
or U671 (N_671,In_874,In_747);
and U672 (N_672,In_666,In_468);
and U673 (N_673,In_157,In_969);
nand U674 (N_674,In_185,In_633);
and U675 (N_675,In_719,In_143);
and U676 (N_676,In_307,In_159);
nor U677 (N_677,In_241,In_321);
nand U678 (N_678,In_546,In_36);
nand U679 (N_679,In_795,In_754);
or U680 (N_680,In_636,In_578);
nand U681 (N_681,In_657,In_941);
or U682 (N_682,In_793,In_326);
and U683 (N_683,In_774,In_430);
nor U684 (N_684,In_676,In_765);
nor U685 (N_685,In_486,In_906);
nor U686 (N_686,In_347,In_186);
or U687 (N_687,In_983,In_197);
and U688 (N_688,In_956,In_571);
and U689 (N_689,In_579,In_775);
nand U690 (N_690,In_520,In_651);
or U691 (N_691,In_97,In_444);
nor U692 (N_692,In_279,In_929);
or U693 (N_693,In_956,In_925);
or U694 (N_694,In_14,In_250);
or U695 (N_695,In_406,In_53);
nand U696 (N_696,In_911,In_38);
and U697 (N_697,In_556,In_839);
nand U698 (N_698,In_504,In_675);
nor U699 (N_699,In_910,In_485);
nand U700 (N_700,In_395,In_772);
nand U701 (N_701,In_570,In_647);
nand U702 (N_702,In_973,In_251);
or U703 (N_703,In_305,In_774);
or U704 (N_704,In_25,In_555);
and U705 (N_705,In_186,In_390);
nand U706 (N_706,In_319,In_10);
nand U707 (N_707,In_786,In_950);
nand U708 (N_708,In_223,In_279);
or U709 (N_709,In_624,In_920);
or U710 (N_710,In_384,In_66);
and U711 (N_711,In_559,In_468);
nand U712 (N_712,In_904,In_886);
nand U713 (N_713,In_561,In_892);
nand U714 (N_714,In_492,In_224);
nand U715 (N_715,In_445,In_241);
and U716 (N_716,In_261,In_499);
and U717 (N_717,In_831,In_669);
nor U718 (N_718,In_82,In_787);
nor U719 (N_719,In_83,In_983);
nand U720 (N_720,In_567,In_798);
nand U721 (N_721,In_903,In_329);
nand U722 (N_722,In_839,In_436);
and U723 (N_723,In_234,In_960);
nand U724 (N_724,In_459,In_764);
nand U725 (N_725,In_63,In_409);
nand U726 (N_726,In_892,In_448);
or U727 (N_727,In_414,In_556);
or U728 (N_728,In_868,In_151);
or U729 (N_729,In_351,In_888);
or U730 (N_730,In_323,In_860);
nand U731 (N_731,In_736,In_906);
or U732 (N_732,In_270,In_288);
nor U733 (N_733,In_543,In_69);
or U734 (N_734,In_351,In_320);
or U735 (N_735,In_606,In_787);
or U736 (N_736,In_944,In_33);
or U737 (N_737,In_77,In_278);
nand U738 (N_738,In_708,In_983);
or U739 (N_739,In_922,In_760);
nor U740 (N_740,In_604,In_952);
or U741 (N_741,In_188,In_92);
or U742 (N_742,In_29,In_321);
or U743 (N_743,In_801,In_398);
or U744 (N_744,In_864,In_775);
nand U745 (N_745,In_955,In_284);
and U746 (N_746,In_982,In_462);
nand U747 (N_747,In_536,In_308);
and U748 (N_748,In_34,In_404);
or U749 (N_749,In_347,In_420);
nor U750 (N_750,In_681,In_133);
and U751 (N_751,In_110,In_63);
nand U752 (N_752,In_70,In_324);
and U753 (N_753,In_633,In_290);
nor U754 (N_754,In_36,In_474);
and U755 (N_755,In_546,In_945);
and U756 (N_756,In_829,In_638);
nand U757 (N_757,In_393,In_785);
or U758 (N_758,In_433,In_534);
nand U759 (N_759,In_550,In_76);
or U760 (N_760,In_940,In_78);
nand U761 (N_761,In_548,In_119);
or U762 (N_762,In_43,In_697);
and U763 (N_763,In_807,In_340);
nand U764 (N_764,In_507,In_941);
and U765 (N_765,In_38,In_435);
and U766 (N_766,In_20,In_508);
nand U767 (N_767,In_815,In_479);
and U768 (N_768,In_39,In_93);
nor U769 (N_769,In_652,In_445);
nand U770 (N_770,In_373,In_660);
nand U771 (N_771,In_570,In_838);
nand U772 (N_772,In_705,In_702);
or U773 (N_773,In_534,In_95);
nand U774 (N_774,In_303,In_768);
or U775 (N_775,In_654,In_124);
nand U776 (N_776,In_15,In_31);
nand U777 (N_777,In_183,In_49);
and U778 (N_778,In_626,In_105);
or U779 (N_779,In_578,In_741);
or U780 (N_780,In_71,In_49);
and U781 (N_781,In_727,In_521);
nand U782 (N_782,In_316,In_565);
and U783 (N_783,In_5,In_939);
and U784 (N_784,In_62,In_924);
nor U785 (N_785,In_10,In_995);
nor U786 (N_786,In_344,In_77);
nand U787 (N_787,In_26,In_96);
nor U788 (N_788,In_50,In_670);
nor U789 (N_789,In_428,In_251);
nand U790 (N_790,In_984,In_912);
nand U791 (N_791,In_485,In_225);
nand U792 (N_792,In_591,In_17);
nand U793 (N_793,In_265,In_86);
and U794 (N_794,In_595,In_700);
or U795 (N_795,In_847,In_725);
and U796 (N_796,In_706,In_698);
nor U797 (N_797,In_177,In_25);
nor U798 (N_798,In_1,In_991);
and U799 (N_799,In_390,In_454);
nand U800 (N_800,In_118,In_484);
nor U801 (N_801,In_106,In_80);
or U802 (N_802,In_236,In_447);
or U803 (N_803,In_106,In_415);
nor U804 (N_804,In_540,In_936);
and U805 (N_805,In_852,In_507);
xnor U806 (N_806,In_176,In_28);
nor U807 (N_807,In_950,In_600);
and U808 (N_808,In_275,In_230);
or U809 (N_809,In_486,In_887);
nor U810 (N_810,In_553,In_654);
and U811 (N_811,In_855,In_306);
nand U812 (N_812,In_547,In_380);
nor U813 (N_813,In_491,In_307);
and U814 (N_814,In_196,In_625);
and U815 (N_815,In_151,In_344);
nand U816 (N_816,In_864,In_589);
nor U817 (N_817,In_751,In_290);
or U818 (N_818,In_600,In_14);
and U819 (N_819,In_712,In_160);
nand U820 (N_820,In_889,In_5);
nand U821 (N_821,In_300,In_43);
or U822 (N_822,In_997,In_183);
nor U823 (N_823,In_226,In_706);
nor U824 (N_824,In_433,In_609);
nand U825 (N_825,In_414,In_553);
nor U826 (N_826,In_837,In_892);
nand U827 (N_827,In_182,In_345);
and U828 (N_828,In_131,In_814);
nand U829 (N_829,In_75,In_320);
and U830 (N_830,In_945,In_128);
and U831 (N_831,In_738,In_439);
or U832 (N_832,In_430,In_96);
nor U833 (N_833,In_382,In_844);
nor U834 (N_834,In_841,In_555);
and U835 (N_835,In_275,In_466);
nor U836 (N_836,In_546,In_524);
and U837 (N_837,In_308,In_343);
nand U838 (N_838,In_185,In_539);
nand U839 (N_839,In_787,In_925);
nand U840 (N_840,In_740,In_973);
or U841 (N_841,In_52,In_76);
and U842 (N_842,In_236,In_214);
nor U843 (N_843,In_905,In_555);
nor U844 (N_844,In_734,In_354);
nor U845 (N_845,In_121,In_846);
nand U846 (N_846,In_484,In_924);
nor U847 (N_847,In_192,In_411);
nor U848 (N_848,In_585,In_101);
nor U849 (N_849,In_665,In_406);
and U850 (N_850,In_189,In_100);
nor U851 (N_851,In_434,In_505);
nand U852 (N_852,In_126,In_82);
or U853 (N_853,In_376,In_743);
or U854 (N_854,In_779,In_226);
nand U855 (N_855,In_74,In_337);
or U856 (N_856,In_361,In_742);
nand U857 (N_857,In_261,In_318);
and U858 (N_858,In_819,In_701);
nor U859 (N_859,In_404,In_758);
nor U860 (N_860,In_817,In_516);
and U861 (N_861,In_600,In_731);
or U862 (N_862,In_782,In_580);
and U863 (N_863,In_117,In_869);
nor U864 (N_864,In_157,In_196);
nand U865 (N_865,In_612,In_55);
and U866 (N_866,In_96,In_260);
nand U867 (N_867,In_166,In_894);
and U868 (N_868,In_164,In_657);
and U869 (N_869,In_258,In_495);
and U870 (N_870,In_209,In_773);
nand U871 (N_871,In_91,In_708);
and U872 (N_872,In_769,In_423);
or U873 (N_873,In_635,In_630);
or U874 (N_874,In_701,In_910);
or U875 (N_875,In_186,In_296);
or U876 (N_876,In_810,In_319);
and U877 (N_877,In_912,In_537);
nand U878 (N_878,In_366,In_948);
and U879 (N_879,In_495,In_645);
or U880 (N_880,In_436,In_207);
nor U881 (N_881,In_931,In_60);
and U882 (N_882,In_852,In_996);
nor U883 (N_883,In_754,In_771);
or U884 (N_884,In_354,In_755);
or U885 (N_885,In_219,In_858);
or U886 (N_886,In_462,In_384);
and U887 (N_887,In_199,In_933);
xor U888 (N_888,In_490,In_799);
or U889 (N_889,In_650,In_305);
or U890 (N_890,In_365,In_517);
nand U891 (N_891,In_194,In_362);
nand U892 (N_892,In_571,In_813);
or U893 (N_893,In_721,In_967);
nor U894 (N_894,In_114,In_491);
or U895 (N_895,In_937,In_591);
nand U896 (N_896,In_288,In_733);
and U897 (N_897,In_913,In_401);
and U898 (N_898,In_807,In_504);
nor U899 (N_899,In_731,In_800);
nand U900 (N_900,In_364,In_198);
nor U901 (N_901,In_90,In_786);
and U902 (N_902,In_80,In_640);
nand U903 (N_903,In_168,In_819);
and U904 (N_904,In_267,In_782);
or U905 (N_905,In_79,In_952);
or U906 (N_906,In_680,In_202);
and U907 (N_907,In_908,In_857);
and U908 (N_908,In_776,In_97);
and U909 (N_909,In_418,In_590);
or U910 (N_910,In_336,In_662);
nand U911 (N_911,In_702,In_102);
and U912 (N_912,In_967,In_462);
nor U913 (N_913,In_340,In_283);
or U914 (N_914,In_995,In_801);
nand U915 (N_915,In_645,In_946);
or U916 (N_916,In_894,In_845);
or U917 (N_917,In_708,In_514);
or U918 (N_918,In_919,In_772);
or U919 (N_919,In_43,In_136);
or U920 (N_920,In_687,In_805);
nand U921 (N_921,In_388,In_163);
nor U922 (N_922,In_85,In_183);
nand U923 (N_923,In_924,In_982);
or U924 (N_924,In_945,In_557);
and U925 (N_925,In_960,In_878);
and U926 (N_926,In_380,In_622);
nand U927 (N_927,In_510,In_432);
nor U928 (N_928,In_333,In_548);
nand U929 (N_929,In_651,In_226);
and U930 (N_930,In_85,In_419);
xnor U931 (N_931,In_590,In_627);
nand U932 (N_932,In_47,In_805);
and U933 (N_933,In_639,In_427);
and U934 (N_934,In_178,In_357);
nor U935 (N_935,In_931,In_325);
and U936 (N_936,In_592,In_184);
and U937 (N_937,In_468,In_391);
nor U938 (N_938,In_840,In_304);
nor U939 (N_939,In_51,In_111);
nor U940 (N_940,In_733,In_598);
or U941 (N_941,In_639,In_267);
nor U942 (N_942,In_326,In_212);
and U943 (N_943,In_443,In_652);
nand U944 (N_944,In_877,In_330);
or U945 (N_945,In_959,In_797);
nor U946 (N_946,In_218,In_236);
nand U947 (N_947,In_410,In_917);
nor U948 (N_948,In_916,In_829);
nand U949 (N_949,In_797,In_245);
xnor U950 (N_950,In_668,In_934);
and U951 (N_951,In_842,In_832);
or U952 (N_952,In_256,In_67);
and U953 (N_953,In_844,In_552);
nor U954 (N_954,In_282,In_785);
and U955 (N_955,In_122,In_721);
and U956 (N_956,In_145,In_95);
nor U957 (N_957,In_619,In_894);
nor U958 (N_958,In_947,In_488);
and U959 (N_959,In_7,In_8);
nor U960 (N_960,In_106,In_592);
nand U961 (N_961,In_446,In_287);
or U962 (N_962,In_257,In_505);
nor U963 (N_963,In_738,In_838);
nor U964 (N_964,In_643,In_288);
or U965 (N_965,In_415,In_157);
or U966 (N_966,In_446,In_563);
or U967 (N_967,In_174,In_759);
nor U968 (N_968,In_396,In_851);
or U969 (N_969,In_352,In_68);
and U970 (N_970,In_826,In_368);
nor U971 (N_971,In_286,In_72);
nor U972 (N_972,In_100,In_278);
and U973 (N_973,In_264,In_774);
nor U974 (N_974,In_540,In_674);
nor U975 (N_975,In_435,In_810);
nand U976 (N_976,In_510,In_343);
nor U977 (N_977,In_622,In_181);
nor U978 (N_978,In_103,In_540);
or U979 (N_979,In_249,In_292);
nor U980 (N_980,In_409,In_28);
or U981 (N_981,In_466,In_18);
or U982 (N_982,In_306,In_368);
or U983 (N_983,In_369,In_973);
or U984 (N_984,In_781,In_311);
nand U985 (N_985,In_681,In_86);
and U986 (N_986,In_581,In_488);
and U987 (N_987,In_250,In_666);
nor U988 (N_988,In_752,In_640);
nand U989 (N_989,In_811,In_385);
nor U990 (N_990,In_945,In_75);
nor U991 (N_991,In_90,In_966);
and U992 (N_992,In_530,In_953);
and U993 (N_993,In_223,In_221);
nor U994 (N_994,In_186,In_194);
nor U995 (N_995,In_92,In_762);
or U996 (N_996,In_407,In_142);
or U997 (N_997,In_75,In_734);
nand U998 (N_998,In_96,In_321);
nor U999 (N_999,In_900,In_896);
nor U1000 (N_1000,In_416,In_586);
nor U1001 (N_1001,In_126,In_209);
nor U1002 (N_1002,In_27,In_502);
nand U1003 (N_1003,In_441,In_367);
and U1004 (N_1004,In_138,In_898);
nor U1005 (N_1005,In_940,In_227);
or U1006 (N_1006,In_93,In_961);
nand U1007 (N_1007,In_528,In_743);
and U1008 (N_1008,In_582,In_511);
nand U1009 (N_1009,In_366,In_779);
xnor U1010 (N_1010,In_606,In_172);
or U1011 (N_1011,In_803,In_584);
or U1012 (N_1012,In_395,In_763);
nor U1013 (N_1013,In_433,In_769);
and U1014 (N_1014,In_728,In_298);
nand U1015 (N_1015,In_864,In_432);
nand U1016 (N_1016,In_336,In_949);
nor U1017 (N_1017,In_549,In_192);
nor U1018 (N_1018,In_403,In_421);
nand U1019 (N_1019,In_846,In_680);
nand U1020 (N_1020,In_246,In_721);
or U1021 (N_1021,In_343,In_698);
nand U1022 (N_1022,In_934,In_845);
and U1023 (N_1023,In_826,In_716);
nand U1024 (N_1024,In_47,In_815);
and U1025 (N_1025,In_603,In_410);
nand U1026 (N_1026,In_254,In_945);
or U1027 (N_1027,In_949,In_255);
or U1028 (N_1028,In_833,In_384);
and U1029 (N_1029,In_500,In_41);
nor U1030 (N_1030,In_670,In_399);
nand U1031 (N_1031,In_488,In_849);
nand U1032 (N_1032,In_610,In_767);
nand U1033 (N_1033,In_896,In_691);
or U1034 (N_1034,In_915,In_690);
or U1035 (N_1035,In_238,In_377);
and U1036 (N_1036,In_623,In_636);
and U1037 (N_1037,In_218,In_545);
nand U1038 (N_1038,In_711,In_151);
or U1039 (N_1039,In_536,In_738);
and U1040 (N_1040,In_454,In_768);
or U1041 (N_1041,In_113,In_88);
or U1042 (N_1042,In_431,In_134);
and U1043 (N_1043,In_144,In_556);
xnor U1044 (N_1044,In_598,In_936);
and U1045 (N_1045,In_724,In_704);
and U1046 (N_1046,In_411,In_612);
nor U1047 (N_1047,In_98,In_717);
nor U1048 (N_1048,In_979,In_585);
or U1049 (N_1049,In_837,In_286);
and U1050 (N_1050,In_261,In_54);
nand U1051 (N_1051,In_303,In_440);
nand U1052 (N_1052,In_932,In_560);
and U1053 (N_1053,In_126,In_280);
or U1054 (N_1054,In_795,In_945);
and U1055 (N_1055,In_211,In_735);
or U1056 (N_1056,In_560,In_631);
or U1057 (N_1057,In_523,In_947);
nor U1058 (N_1058,In_177,In_238);
nand U1059 (N_1059,In_513,In_207);
or U1060 (N_1060,In_143,In_653);
and U1061 (N_1061,In_977,In_374);
or U1062 (N_1062,In_602,In_383);
and U1063 (N_1063,In_584,In_999);
and U1064 (N_1064,In_807,In_640);
nor U1065 (N_1065,In_753,In_417);
nand U1066 (N_1066,In_808,In_70);
and U1067 (N_1067,In_405,In_26);
or U1068 (N_1068,In_633,In_162);
and U1069 (N_1069,In_18,In_931);
or U1070 (N_1070,In_388,In_625);
nor U1071 (N_1071,In_677,In_752);
or U1072 (N_1072,In_410,In_490);
nor U1073 (N_1073,In_511,In_376);
and U1074 (N_1074,In_615,In_787);
nand U1075 (N_1075,In_920,In_478);
or U1076 (N_1076,In_854,In_855);
nand U1077 (N_1077,In_42,In_521);
nor U1078 (N_1078,In_219,In_461);
or U1079 (N_1079,In_657,In_636);
nor U1080 (N_1080,In_363,In_872);
nand U1081 (N_1081,In_373,In_254);
nor U1082 (N_1082,In_929,In_959);
or U1083 (N_1083,In_281,In_911);
or U1084 (N_1084,In_834,In_43);
nand U1085 (N_1085,In_655,In_623);
nor U1086 (N_1086,In_156,In_908);
nand U1087 (N_1087,In_64,In_174);
and U1088 (N_1088,In_473,In_967);
and U1089 (N_1089,In_952,In_972);
and U1090 (N_1090,In_433,In_626);
nand U1091 (N_1091,In_884,In_523);
or U1092 (N_1092,In_305,In_625);
nand U1093 (N_1093,In_752,In_669);
nand U1094 (N_1094,In_264,In_700);
or U1095 (N_1095,In_172,In_538);
nand U1096 (N_1096,In_285,In_680);
and U1097 (N_1097,In_359,In_250);
or U1098 (N_1098,In_294,In_491);
nor U1099 (N_1099,In_922,In_859);
nor U1100 (N_1100,In_32,In_798);
or U1101 (N_1101,In_629,In_901);
nand U1102 (N_1102,In_850,In_596);
or U1103 (N_1103,In_148,In_917);
nor U1104 (N_1104,In_764,In_332);
nor U1105 (N_1105,In_71,In_344);
nor U1106 (N_1106,In_345,In_364);
or U1107 (N_1107,In_946,In_992);
nand U1108 (N_1108,In_269,In_373);
nor U1109 (N_1109,In_558,In_26);
nand U1110 (N_1110,In_218,In_984);
nand U1111 (N_1111,In_26,In_389);
nor U1112 (N_1112,In_686,In_443);
and U1113 (N_1113,In_983,In_794);
or U1114 (N_1114,In_450,In_806);
or U1115 (N_1115,In_194,In_298);
and U1116 (N_1116,In_266,In_737);
or U1117 (N_1117,In_675,In_795);
and U1118 (N_1118,In_454,In_594);
xnor U1119 (N_1119,In_714,In_25);
nand U1120 (N_1120,In_807,In_207);
or U1121 (N_1121,In_118,In_127);
or U1122 (N_1122,In_417,In_805);
and U1123 (N_1123,In_131,In_607);
and U1124 (N_1124,In_172,In_724);
or U1125 (N_1125,In_593,In_332);
nor U1126 (N_1126,In_983,In_716);
nand U1127 (N_1127,In_815,In_717);
nor U1128 (N_1128,In_867,In_187);
or U1129 (N_1129,In_463,In_356);
nand U1130 (N_1130,In_390,In_442);
or U1131 (N_1131,In_24,In_465);
and U1132 (N_1132,In_361,In_512);
and U1133 (N_1133,In_204,In_64);
and U1134 (N_1134,In_503,In_87);
and U1135 (N_1135,In_40,In_860);
nand U1136 (N_1136,In_229,In_273);
xor U1137 (N_1137,In_670,In_132);
nand U1138 (N_1138,In_981,In_602);
nor U1139 (N_1139,In_802,In_434);
nand U1140 (N_1140,In_173,In_216);
or U1141 (N_1141,In_240,In_421);
nor U1142 (N_1142,In_321,In_449);
or U1143 (N_1143,In_415,In_909);
xor U1144 (N_1144,In_805,In_182);
and U1145 (N_1145,In_546,In_973);
nor U1146 (N_1146,In_143,In_778);
nand U1147 (N_1147,In_125,In_75);
or U1148 (N_1148,In_989,In_462);
nor U1149 (N_1149,In_523,In_529);
nand U1150 (N_1150,In_453,In_239);
and U1151 (N_1151,In_578,In_325);
and U1152 (N_1152,In_754,In_958);
nor U1153 (N_1153,In_26,In_709);
and U1154 (N_1154,In_612,In_650);
or U1155 (N_1155,In_675,In_34);
and U1156 (N_1156,In_388,In_337);
xnor U1157 (N_1157,In_161,In_319);
or U1158 (N_1158,In_247,In_784);
nor U1159 (N_1159,In_114,In_942);
and U1160 (N_1160,In_19,In_76);
nand U1161 (N_1161,In_99,In_943);
nand U1162 (N_1162,In_509,In_996);
nand U1163 (N_1163,In_303,In_283);
nor U1164 (N_1164,In_126,In_853);
or U1165 (N_1165,In_537,In_427);
nand U1166 (N_1166,In_156,In_644);
nand U1167 (N_1167,In_273,In_296);
nor U1168 (N_1168,In_844,In_418);
nor U1169 (N_1169,In_954,In_629);
and U1170 (N_1170,In_357,In_289);
nand U1171 (N_1171,In_83,In_397);
or U1172 (N_1172,In_274,In_781);
and U1173 (N_1173,In_186,In_703);
and U1174 (N_1174,In_271,In_141);
nor U1175 (N_1175,In_925,In_917);
and U1176 (N_1176,In_446,In_671);
and U1177 (N_1177,In_320,In_477);
or U1178 (N_1178,In_582,In_175);
or U1179 (N_1179,In_106,In_186);
nor U1180 (N_1180,In_519,In_968);
nor U1181 (N_1181,In_648,In_282);
or U1182 (N_1182,In_734,In_660);
nand U1183 (N_1183,In_710,In_355);
nor U1184 (N_1184,In_761,In_16);
or U1185 (N_1185,In_828,In_613);
nor U1186 (N_1186,In_288,In_856);
nor U1187 (N_1187,In_858,In_71);
nor U1188 (N_1188,In_632,In_854);
nand U1189 (N_1189,In_327,In_999);
nand U1190 (N_1190,In_223,In_83);
nand U1191 (N_1191,In_621,In_371);
nor U1192 (N_1192,In_438,In_654);
or U1193 (N_1193,In_308,In_698);
nor U1194 (N_1194,In_711,In_64);
and U1195 (N_1195,In_404,In_278);
nor U1196 (N_1196,In_891,In_382);
and U1197 (N_1197,In_332,In_755);
nand U1198 (N_1198,In_397,In_378);
nor U1199 (N_1199,In_730,In_248);
or U1200 (N_1200,In_743,In_850);
and U1201 (N_1201,In_989,In_357);
nor U1202 (N_1202,In_56,In_851);
nand U1203 (N_1203,In_622,In_35);
or U1204 (N_1204,In_372,In_418);
nor U1205 (N_1205,In_539,In_378);
or U1206 (N_1206,In_619,In_74);
or U1207 (N_1207,In_495,In_1);
nand U1208 (N_1208,In_122,In_841);
and U1209 (N_1209,In_834,In_779);
or U1210 (N_1210,In_403,In_97);
nand U1211 (N_1211,In_817,In_905);
nand U1212 (N_1212,In_744,In_754);
or U1213 (N_1213,In_232,In_906);
nor U1214 (N_1214,In_148,In_305);
or U1215 (N_1215,In_273,In_436);
nand U1216 (N_1216,In_916,In_831);
and U1217 (N_1217,In_43,In_850);
or U1218 (N_1218,In_51,In_800);
nand U1219 (N_1219,In_347,In_292);
or U1220 (N_1220,In_942,In_538);
or U1221 (N_1221,In_990,In_476);
or U1222 (N_1222,In_730,In_59);
and U1223 (N_1223,In_95,In_19);
or U1224 (N_1224,In_284,In_706);
and U1225 (N_1225,In_345,In_764);
and U1226 (N_1226,In_451,In_527);
or U1227 (N_1227,In_674,In_765);
and U1228 (N_1228,In_248,In_789);
nand U1229 (N_1229,In_808,In_767);
nand U1230 (N_1230,In_312,In_463);
or U1231 (N_1231,In_552,In_367);
or U1232 (N_1232,In_565,In_626);
nor U1233 (N_1233,In_157,In_268);
and U1234 (N_1234,In_382,In_654);
and U1235 (N_1235,In_167,In_745);
and U1236 (N_1236,In_791,In_368);
nor U1237 (N_1237,In_325,In_301);
or U1238 (N_1238,In_38,In_530);
and U1239 (N_1239,In_55,In_474);
nor U1240 (N_1240,In_539,In_991);
or U1241 (N_1241,In_153,In_402);
nand U1242 (N_1242,In_381,In_612);
nand U1243 (N_1243,In_480,In_239);
or U1244 (N_1244,In_584,In_301);
and U1245 (N_1245,In_637,In_99);
nor U1246 (N_1246,In_124,In_250);
nand U1247 (N_1247,In_360,In_528);
or U1248 (N_1248,In_365,In_434);
and U1249 (N_1249,In_156,In_767);
nand U1250 (N_1250,In_257,In_432);
xor U1251 (N_1251,In_512,In_830);
and U1252 (N_1252,In_673,In_453);
nand U1253 (N_1253,In_907,In_618);
and U1254 (N_1254,In_260,In_223);
nand U1255 (N_1255,In_243,In_719);
or U1256 (N_1256,In_623,In_595);
and U1257 (N_1257,In_775,In_802);
nor U1258 (N_1258,In_149,In_584);
nand U1259 (N_1259,In_566,In_429);
nand U1260 (N_1260,In_833,In_435);
nor U1261 (N_1261,In_823,In_225);
nand U1262 (N_1262,In_339,In_955);
and U1263 (N_1263,In_539,In_939);
nor U1264 (N_1264,In_469,In_422);
or U1265 (N_1265,In_948,In_466);
and U1266 (N_1266,In_623,In_654);
nand U1267 (N_1267,In_294,In_477);
or U1268 (N_1268,In_709,In_105);
and U1269 (N_1269,In_894,In_861);
and U1270 (N_1270,In_210,In_774);
nand U1271 (N_1271,In_215,In_278);
nor U1272 (N_1272,In_371,In_393);
or U1273 (N_1273,In_327,In_691);
and U1274 (N_1274,In_439,In_611);
nand U1275 (N_1275,In_758,In_686);
nor U1276 (N_1276,In_356,In_992);
nor U1277 (N_1277,In_522,In_7);
nand U1278 (N_1278,In_152,In_675);
nand U1279 (N_1279,In_970,In_257);
or U1280 (N_1280,In_420,In_766);
and U1281 (N_1281,In_524,In_893);
and U1282 (N_1282,In_996,In_525);
nand U1283 (N_1283,In_230,In_573);
and U1284 (N_1284,In_547,In_213);
nor U1285 (N_1285,In_325,In_137);
or U1286 (N_1286,In_855,In_417);
and U1287 (N_1287,In_291,In_892);
and U1288 (N_1288,In_844,In_554);
or U1289 (N_1289,In_533,In_438);
or U1290 (N_1290,In_299,In_702);
and U1291 (N_1291,In_175,In_462);
or U1292 (N_1292,In_222,In_31);
nand U1293 (N_1293,In_558,In_180);
nor U1294 (N_1294,In_546,In_640);
nor U1295 (N_1295,In_568,In_905);
nand U1296 (N_1296,In_767,In_24);
nor U1297 (N_1297,In_511,In_462);
and U1298 (N_1298,In_912,In_29);
nand U1299 (N_1299,In_29,In_145);
or U1300 (N_1300,In_333,In_526);
or U1301 (N_1301,In_446,In_646);
nor U1302 (N_1302,In_316,In_976);
nor U1303 (N_1303,In_427,In_640);
or U1304 (N_1304,In_427,In_657);
nand U1305 (N_1305,In_300,In_128);
and U1306 (N_1306,In_701,In_358);
xnor U1307 (N_1307,In_395,In_482);
nor U1308 (N_1308,In_560,In_251);
or U1309 (N_1309,In_960,In_128);
nand U1310 (N_1310,In_413,In_873);
and U1311 (N_1311,In_496,In_533);
nor U1312 (N_1312,In_514,In_400);
nand U1313 (N_1313,In_182,In_996);
xor U1314 (N_1314,In_308,In_569);
or U1315 (N_1315,In_31,In_895);
nand U1316 (N_1316,In_58,In_162);
or U1317 (N_1317,In_91,In_464);
nand U1318 (N_1318,In_570,In_133);
and U1319 (N_1319,In_64,In_714);
or U1320 (N_1320,In_693,In_237);
or U1321 (N_1321,In_87,In_449);
nand U1322 (N_1322,In_476,In_530);
and U1323 (N_1323,In_291,In_820);
nor U1324 (N_1324,In_302,In_655);
nor U1325 (N_1325,In_13,In_725);
nand U1326 (N_1326,In_823,In_490);
nor U1327 (N_1327,In_583,In_471);
and U1328 (N_1328,In_359,In_860);
nand U1329 (N_1329,In_243,In_128);
and U1330 (N_1330,In_323,In_673);
nand U1331 (N_1331,In_676,In_205);
nand U1332 (N_1332,In_455,In_563);
or U1333 (N_1333,In_601,In_257);
and U1334 (N_1334,In_644,In_442);
and U1335 (N_1335,In_356,In_308);
and U1336 (N_1336,In_889,In_439);
and U1337 (N_1337,In_628,In_988);
nand U1338 (N_1338,In_793,In_154);
nor U1339 (N_1339,In_728,In_185);
or U1340 (N_1340,In_176,In_904);
nor U1341 (N_1341,In_139,In_100);
xor U1342 (N_1342,In_11,In_496);
or U1343 (N_1343,In_413,In_796);
nor U1344 (N_1344,In_611,In_151);
nand U1345 (N_1345,In_409,In_250);
or U1346 (N_1346,In_559,In_792);
nand U1347 (N_1347,In_433,In_51);
or U1348 (N_1348,In_296,In_158);
nor U1349 (N_1349,In_448,In_363);
and U1350 (N_1350,In_387,In_15);
or U1351 (N_1351,In_13,In_955);
nand U1352 (N_1352,In_905,In_632);
or U1353 (N_1353,In_808,In_549);
and U1354 (N_1354,In_453,In_57);
and U1355 (N_1355,In_993,In_966);
nand U1356 (N_1356,In_702,In_932);
nor U1357 (N_1357,In_482,In_474);
xor U1358 (N_1358,In_618,In_719);
or U1359 (N_1359,In_818,In_908);
nor U1360 (N_1360,In_819,In_484);
or U1361 (N_1361,In_106,In_431);
nor U1362 (N_1362,In_851,In_120);
nor U1363 (N_1363,In_474,In_467);
or U1364 (N_1364,In_400,In_232);
or U1365 (N_1365,In_199,In_254);
nand U1366 (N_1366,In_831,In_423);
or U1367 (N_1367,In_438,In_121);
and U1368 (N_1368,In_293,In_155);
nand U1369 (N_1369,In_510,In_459);
and U1370 (N_1370,In_41,In_731);
or U1371 (N_1371,In_948,In_892);
nand U1372 (N_1372,In_322,In_665);
or U1373 (N_1373,In_801,In_581);
or U1374 (N_1374,In_502,In_905);
nor U1375 (N_1375,In_547,In_400);
nor U1376 (N_1376,In_138,In_610);
or U1377 (N_1377,In_610,In_956);
and U1378 (N_1378,In_767,In_961);
nand U1379 (N_1379,In_486,In_184);
nor U1380 (N_1380,In_811,In_230);
and U1381 (N_1381,In_937,In_563);
or U1382 (N_1382,In_275,In_606);
nor U1383 (N_1383,In_96,In_442);
or U1384 (N_1384,In_485,In_655);
nor U1385 (N_1385,In_736,In_415);
and U1386 (N_1386,In_906,In_411);
and U1387 (N_1387,In_483,In_244);
nand U1388 (N_1388,In_904,In_848);
nand U1389 (N_1389,In_615,In_63);
nor U1390 (N_1390,In_220,In_20);
nand U1391 (N_1391,In_515,In_577);
nor U1392 (N_1392,In_438,In_247);
and U1393 (N_1393,In_706,In_17);
nor U1394 (N_1394,In_62,In_682);
nor U1395 (N_1395,In_687,In_623);
or U1396 (N_1396,In_479,In_441);
nand U1397 (N_1397,In_785,In_580);
nand U1398 (N_1398,In_854,In_686);
nand U1399 (N_1399,In_40,In_426);
nor U1400 (N_1400,In_943,In_660);
and U1401 (N_1401,In_222,In_660);
and U1402 (N_1402,In_775,In_931);
and U1403 (N_1403,In_852,In_797);
nand U1404 (N_1404,In_991,In_358);
nand U1405 (N_1405,In_751,In_989);
nand U1406 (N_1406,In_872,In_802);
nand U1407 (N_1407,In_78,In_653);
nor U1408 (N_1408,In_843,In_464);
nor U1409 (N_1409,In_955,In_24);
and U1410 (N_1410,In_206,In_109);
nor U1411 (N_1411,In_744,In_323);
nand U1412 (N_1412,In_471,In_516);
nand U1413 (N_1413,In_8,In_103);
nand U1414 (N_1414,In_515,In_458);
and U1415 (N_1415,In_200,In_383);
nand U1416 (N_1416,In_361,In_530);
and U1417 (N_1417,In_955,In_945);
nor U1418 (N_1418,In_107,In_961);
or U1419 (N_1419,In_769,In_442);
and U1420 (N_1420,In_263,In_346);
or U1421 (N_1421,In_204,In_94);
or U1422 (N_1422,In_844,In_453);
or U1423 (N_1423,In_322,In_951);
nor U1424 (N_1424,In_950,In_565);
or U1425 (N_1425,In_616,In_250);
nor U1426 (N_1426,In_169,In_828);
xor U1427 (N_1427,In_639,In_259);
nor U1428 (N_1428,In_305,In_187);
xor U1429 (N_1429,In_584,In_229);
and U1430 (N_1430,In_354,In_454);
or U1431 (N_1431,In_758,In_691);
and U1432 (N_1432,In_489,In_809);
or U1433 (N_1433,In_737,In_530);
or U1434 (N_1434,In_539,In_276);
nand U1435 (N_1435,In_404,In_399);
and U1436 (N_1436,In_596,In_680);
nor U1437 (N_1437,In_224,In_309);
or U1438 (N_1438,In_409,In_194);
nand U1439 (N_1439,In_626,In_561);
nand U1440 (N_1440,In_863,In_402);
or U1441 (N_1441,In_878,In_403);
or U1442 (N_1442,In_323,In_947);
and U1443 (N_1443,In_227,In_679);
or U1444 (N_1444,In_840,In_969);
nand U1445 (N_1445,In_443,In_169);
or U1446 (N_1446,In_470,In_674);
nor U1447 (N_1447,In_794,In_986);
nand U1448 (N_1448,In_8,In_377);
and U1449 (N_1449,In_535,In_199);
and U1450 (N_1450,In_866,In_477);
nor U1451 (N_1451,In_138,In_381);
or U1452 (N_1452,In_549,In_459);
nor U1453 (N_1453,In_942,In_68);
nor U1454 (N_1454,In_410,In_223);
and U1455 (N_1455,In_267,In_717);
nand U1456 (N_1456,In_308,In_390);
nand U1457 (N_1457,In_952,In_936);
or U1458 (N_1458,In_975,In_699);
nand U1459 (N_1459,In_958,In_665);
or U1460 (N_1460,In_234,In_533);
or U1461 (N_1461,In_681,In_748);
and U1462 (N_1462,In_712,In_594);
or U1463 (N_1463,In_966,In_659);
nand U1464 (N_1464,In_768,In_531);
nand U1465 (N_1465,In_496,In_694);
and U1466 (N_1466,In_889,In_75);
nor U1467 (N_1467,In_500,In_877);
and U1468 (N_1468,In_780,In_468);
nor U1469 (N_1469,In_408,In_722);
or U1470 (N_1470,In_914,In_399);
and U1471 (N_1471,In_818,In_993);
nand U1472 (N_1472,In_71,In_204);
nor U1473 (N_1473,In_593,In_260);
or U1474 (N_1474,In_441,In_740);
nand U1475 (N_1475,In_354,In_29);
and U1476 (N_1476,In_435,In_220);
nor U1477 (N_1477,In_939,In_803);
or U1478 (N_1478,In_910,In_778);
and U1479 (N_1479,In_182,In_135);
and U1480 (N_1480,In_285,In_393);
nor U1481 (N_1481,In_265,In_824);
or U1482 (N_1482,In_915,In_252);
nand U1483 (N_1483,In_302,In_10);
and U1484 (N_1484,In_412,In_238);
nand U1485 (N_1485,In_732,In_541);
nor U1486 (N_1486,In_737,In_227);
and U1487 (N_1487,In_871,In_118);
nor U1488 (N_1488,In_301,In_82);
or U1489 (N_1489,In_873,In_613);
nand U1490 (N_1490,In_576,In_394);
or U1491 (N_1491,In_225,In_708);
nor U1492 (N_1492,In_660,In_390);
nand U1493 (N_1493,In_330,In_933);
nand U1494 (N_1494,In_768,In_723);
nand U1495 (N_1495,In_48,In_142);
nor U1496 (N_1496,In_426,In_92);
or U1497 (N_1497,In_161,In_445);
or U1498 (N_1498,In_86,In_785);
or U1499 (N_1499,In_777,In_82);
and U1500 (N_1500,In_87,In_930);
nor U1501 (N_1501,In_853,In_620);
or U1502 (N_1502,In_93,In_68);
and U1503 (N_1503,In_628,In_802);
and U1504 (N_1504,In_381,In_664);
nor U1505 (N_1505,In_867,In_330);
nand U1506 (N_1506,In_894,In_786);
and U1507 (N_1507,In_298,In_649);
or U1508 (N_1508,In_118,In_82);
nor U1509 (N_1509,In_987,In_340);
and U1510 (N_1510,In_976,In_79);
and U1511 (N_1511,In_778,In_123);
nor U1512 (N_1512,In_496,In_96);
nand U1513 (N_1513,In_759,In_589);
nor U1514 (N_1514,In_482,In_36);
nand U1515 (N_1515,In_516,In_124);
or U1516 (N_1516,In_899,In_751);
nand U1517 (N_1517,In_531,In_6);
nor U1518 (N_1518,In_946,In_628);
nand U1519 (N_1519,In_977,In_665);
and U1520 (N_1520,In_364,In_292);
nand U1521 (N_1521,In_997,In_681);
nand U1522 (N_1522,In_756,In_61);
nand U1523 (N_1523,In_56,In_0);
or U1524 (N_1524,In_990,In_279);
and U1525 (N_1525,In_480,In_732);
xor U1526 (N_1526,In_523,In_679);
or U1527 (N_1527,In_947,In_698);
nand U1528 (N_1528,In_866,In_887);
and U1529 (N_1529,In_771,In_829);
nor U1530 (N_1530,In_150,In_757);
and U1531 (N_1531,In_409,In_11);
nand U1532 (N_1532,In_571,In_3);
and U1533 (N_1533,In_684,In_363);
or U1534 (N_1534,In_156,In_963);
or U1535 (N_1535,In_470,In_864);
or U1536 (N_1536,In_670,In_96);
nand U1537 (N_1537,In_722,In_477);
nor U1538 (N_1538,In_337,In_924);
nand U1539 (N_1539,In_726,In_851);
and U1540 (N_1540,In_511,In_148);
and U1541 (N_1541,In_205,In_403);
nand U1542 (N_1542,In_556,In_380);
nand U1543 (N_1543,In_591,In_149);
nor U1544 (N_1544,In_866,In_638);
nand U1545 (N_1545,In_604,In_855);
and U1546 (N_1546,In_826,In_353);
or U1547 (N_1547,In_598,In_966);
nor U1548 (N_1548,In_925,In_298);
nor U1549 (N_1549,In_46,In_964);
or U1550 (N_1550,In_436,In_252);
and U1551 (N_1551,In_840,In_264);
nand U1552 (N_1552,In_441,In_798);
nor U1553 (N_1553,In_781,In_955);
and U1554 (N_1554,In_827,In_245);
or U1555 (N_1555,In_503,In_875);
nand U1556 (N_1556,In_7,In_593);
or U1557 (N_1557,In_510,In_306);
or U1558 (N_1558,In_510,In_420);
and U1559 (N_1559,In_235,In_453);
nor U1560 (N_1560,In_387,In_628);
nor U1561 (N_1561,In_578,In_44);
nand U1562 (N_1562,In_347,In_948);
nand U1563 (N_1563,In_579,In_315);
nor U1564 (N_1564,In_396,In_982);
nor U1565 (N_1565,In_165,In_728);
nand U1566 (N_1566,In_68,In_217);
nor U1567 (N_1567,In_663,In_804);
nand U1568 (N_1568,In_743,In_600);
or U1569 (N_1569,In_909,In_867);
and U1570 (N_1570,In_195,In_608);
and U1571 (N_1571,In_477,In_173);
nand U1572 (N_1572,In_38,In_701);
or U1573 (N_1573,In_328,In_514);
or U1574 (N_1574,In_454,In_930);
nor U1575 (N_1575,In_912,In_38);
nand U1576 (N_1576,In_135,In_412);
nor U1577 (N_1577,In_103,In_1);
nor U1578 (N_1578,In_433,In_228);
nand U1579 (N_1579,In_985,In_232);
nor U1580 (N_1580,In_5,In_537);
or U1581 (N_1581,In_107,In_609);
and U1582 (N_1582,In_896,In_453);
or U1583 (N_1583,In_991,In_108);
nand U1584 (N_1584,In_407,In_228);
or U1585 (N_1585,In_426,In_118);
nand U1586 (N_1586,In_154,In_905);
nor U1587 (N_1587,In_540,In_121);
nor U1588 (N_1588,In_220,In_766);
and U1589 (N_1589,In_810,In_60);
nand U1590 (N_1590,In_391,In_447);
nand U1591 (N_1591,In_344,In_490);
or U1592 (N_1592,In_607,In_195);
or U1593 (N_1593,In_382,In_148);
or U1594 (N_1594,In_468,In_223);
nand U1595 (N_1595,In_219,In_524);
or U1596 (N_1596,In_388,In_804);
or U1597 (N_1597,In_871,In_656);
nor U1598 (N_1598,In_366,In_333);
or U1599 (N_1599,In_362,In_619);
nor U1600 (N_1600,In_666,In_271);
or U1601 (N_1601,In_951,In_170);
nor U1602 (N_1602,In_263,In_868);
and U1603 (N_1603,In_295,In_553);
and U1604 (N_1604,In_73,In_40);
nor U1605 (N_1605,In_164,In_431);
and U1606 (N_1606,In_333,In_922);
nand U1607 (N_1607,In_678,In_692);
and U1608 (N_1608,In_787,In_486);
nor U1609 (N_1609,In_575,In_647);
nor U1610 (N_1610,In_261,In_956);
nor U1611 (N_1611,In_264,In_702);
or U1612 (N_1612,In_617,In_603);
nor U1613 (N_1613,In_526,In_646);
or U1614 (N_1614,In_172,In_957);
and U1615 (N_1615,In_904,In_737);
and U1616 (N_1616,In_348,In_762);
nand U1617 (N_1617,In_394,In_218);
and U1618 (N_1618,In_833,In_998);
nor U1619 (N_1619,In_908,In_663);
nor U1620 (N_1620,In_477,In_361);
or U1621 (N_1621,In_588,In_599);
nor U1622 (N_1622,In_938,In_479);
nand U1623 (N_1623,In_323,In_328);
nand U1624 (N_1624,In_772,In_699);
and U1625 (N_1625,In_776,In_890);
or U1626 (N_1626,In_311,In_981);
or U1627 (N_1627,In_574,In_403);
and U1628 (N_1628,In_646,In_24);
and U1629 (N_1629,In_555,In_228);
or U1630 (N_1630,In_409,In_299);
and U1631 (N_1631,In_157,In_542);
or U1632 (N_1632,In_738,In_964);
nor U1633 (N_1633,In_685,In_84);
and U1634 (N_1634,In_525,In_731);
nand U1635 (N_1635,In_563,In_818);
nand U1636 (N_1636,In_76,In_637);
and U1637 (N_1637,In_270,In_68);
nand U1638 (N_1638,In_65,In_510);
and U1639 (N_1639,In_92,In_34);
and U1640 (N_1640,In_941,In_819);
and U1641 (N_1641,In_736,In_760);
and U1642 (N_1642,In_34,In_21);
and U1643 (N_1643,In_703,In_217);
and U1644 (N_1644,In_990,In_115);
and U1645 (N_1645,In_511,In_420);
nor U1646 (N_1646,In_481,In_732);
or U1647 (N_1647,In_326,In_413);
nor U1648 (N_1648,In_500,In_726);
nor U1649 (N_1649,In_397,In_362);
xor U1650 (N_1650,In_615,In_721);
nand U1651 (N_1651,In_266,In_643);
or U1652 (N_1652,In_899,In_257);
and U1653 (N_1653,In_938,In_642);
nand U1654 (N_1654,In_650,In_982);
or U1655 (N_1655,In_17,In_450);
nor U1656 (N_1656,In_929,In_923);
or U1657 (N_1657,In_346,In_456);
or U1658 (N_1658,In_760,In_577);
or U1659 (N_1659,In_567,In_131);
and U1660 (N_1660,In_695,In_813);
or U1661 (N_1661,In_321,In_161);
nand U1662 (N_1662,In_961,In_470);
nand U1663 (N_1663,In_416,In_581);
and U1664 (N_1664,In_797,In_685);
xnor U1665 (N_1665,In_293,In_356);
nor U1666 (N_1666,In_498,In_606);
or U1667 (N_1667,In_537,In_2);
nor U1668 (N_1668,In_108,In_501);
and U1669 (N_1669,In_428,In_267);
and U1670 (N_1670,In_654,In_416);
nor U1671 (N_1671,In_224,In_555);
and U1672 (N_1672,In_615,In_280);
and U1673 (N_1673,In_24,In_979);
nor U1674 (N_1674,In_254,In_751);
nor U1675 (N_1675,In_714,In_231);
nor U1676 (N_1676,In_10,In_853);
nand U1677 (N_1677,In_234,In_920);
and U1678 (N_1678,In_525,In_190);
nor U1679 (N_1679,In_6,In_965);
and U1680 (N_1680,In_767,In_989);
nand U1681 (N_1681,In_376,In_405);
nor U1682 (N_1682,In_467,In_149);
and U1683 (N_1683,In_193,In_800);
nor U1684 (N_1684,In_260,In_755);
and U1685 (N_1685,In_387,In_510);
or U1686 (N_1686,In_975,In_96);
and U1687 (N_1687,In_834,In_583);
and U1688 (N_1688,In_390,In_987);
nand U1689 (N_1689,In_403,In_139);
or U1690 (N_1690,In_604,In_311);
nand U1691 (N_1691,In_687,In_123);
or U1692 (N_1692,In_737,In_168);
nor U1693 (N_1693,In_791,In_655);
or U1694 (N_1694,In_523,In_698);
and U1695 (N_1695,In_464,In_37);
and U1696 (N_1696,In_281,In_885);
nand U1697 (N_1697,In_352,In_931);
and U1698 (N_1698,In_761,In_461);
nand U1699 (N_1699,In_120,In_767);
and U1700 (N_1700,In_821,In_158);
nor U1701 (N_1701,In_480,In_824);
or U1702 (N_1702,In_991,In_144);
or U1703 (N_1703,In_73,In_334);
and U1704 (N_1704,In_592,In_502);
or U1705 (N_1705,In_83,In_347);
nand U1706 (N_1706,In_683,In_191);
nand U1707 (N_1707,In_86,In_18);
nor U1708 (N_1708,In_43,In_59);
or U1709 (N_1709,In_56,In_975);
nor U1710 (N_1710,In_782,In_146);
or U1711 (N_1711,In_162,In_107);
or U1712 (N_1712,In_289,In_790);
xor U1713 (N_1713,In_669,In_976);
or U1714 (N_1714,In_235,In_898);
nand U1715 (N_1715,In_483,In_762);
nand U1716 (N_1716,In_628,In_162);
or U1717 (N_1717,In_759,In_555);
nor U1718 (N_1718,In_743,In_891);
and U1719 (N_1719,In_475,In_216);
or U1720 (N_1720,In_918,In_822);
and U1721 (N_1721,In_406,In_960);
or U1722 (N_1722,In_443,In_700);
nor U1723 (N_1723,In_655,In_642);
and U1724 (N_1724,In_367,In_288);
and U1725 (N_1725,In_29,In_894);
and U1726 (N_1726,In_895,In_806);
or U1727 (N_1727,In_152,In_15);
nand U1728 (N_1728,In_713,In_303);
or U1729 (N_1729,In_580,In_175);
nor U1730 (N_1730,In_171,In_215);
or U1731 (N_1731,In_39,In_703);
nor U1732 (N_1732,In_724,In_541);
nand U1733 (N_1733,In_402,In_478);
or U1734 (N_1734,In_427,In_779);
nor U1735 (N_1735,In_179,In_290);
or U1736 (N_1736,In_893,In_804);
or U1737 (N_1737,In_120,In_274);
nor U1738 (N_1738,In_921,In_248);
and U1739 (N_1739,In_648,In_948);
and U1740 (N_1740,In_838,In_413);
and U1741 (N_1741,In_300,In_210);
or U1742 (N_1742,In_727,In_423);
nor U1743 (N_1743,In_272,In_833);
nand U1744 (N_1744,In_775,In_819);
nand U1745 (N_1745,In_643,In_856);
or U1746 (N_1746,In_617,In_427);
and U1747 (N_1747,In_374,In_131);
and U1748 (N_1748,In_658,In_257);
nand U1749 (N_1749,In_472,In_862);
and U1750 (N_1750,In_117,In_83);
xnor U1751 (N_1751,In_872,In_165);
nor U1752 (N_1752,In_454,In_881);
xnor U1753 (N_1753,In_164,In_868);
nand U1754 (N_1754,In_446,In_479);
and U1755 (N_1755,In_627,In_119);
and U1756 (N_1756,In_253,In_86);
nand U1757 (N_1757,In_598,In_796);
nor U1758 (N_1758,In_30,In_141);
nand U1759 (N_1759,In_64,In_502);
xnor U1760 (N_1760,In_603,In_186);
nor U1761 (N_1761,In_19,In_166);
nand U1762 (N_1762,In_271,In_53);
or U1763 (N_1763,In_427,In_918);
nor U1764 (N_1764,In_407,In_616);
or U1765 (N_1765,In_507,In_691);
or U1766 (N_1766,In_447,In_94);
nor U1767 (N_1767,In_116,In_541);
xor U1768 (N_1768,In_521,In_791);
and U1769 (N_1769,In_48,In_81);
and U1770 (N_1770,In_810,In_836);
and U1771 (N_1771,In_938,In_147);
and U1772 (N_1772,In_746,In_52);
or U1773 (N_1773,In_678,In_406);
and U1774 (N_1774,In_306,In_607);
nor U1775 (N_1775,In_939,In_14);
or U1776 (N_1776,In_353,In_571);
and U1777 (N_1777,In_36,In_72);
nor U1778 (N_1778,In_969,In_698);
nand U1779 (N_1779,In_156,In_581);
and U1780 (N_1780,In_20,In_693);
nor U1781 (N_1781,In_729,In_717);
or U1782 (N_1782,In_457,In_973);
nand U1783 (N_1783,In_248,In_238);
nand U1784 (N_1784,In_888,In_274);
and U1785 (N_1785,In_777,In_411);
nand U1786 (N_1786,In_354,In_152);
and U1787 (N_1787,In_763,In_104);
and U1788 (N_1788,In_690,In_392);
or U1789 (N_1789,In_121,In_288);
or U1790 (N_1790,In_462,In_278);
and U1791 (N_1791,In_741,In_191);
and U1792 (N_1792,In_145,In_623);
or U1793 (N_1793,In_763,In_50);
nand U1794 (N_1794,In_997,In_156);
or U1795 (N_1795,In_222,In_740);
or U1796 (N_1796,In_615,In_557);
nand U1797 (N_1797,In_169,In_385);
or U1798 (N_1798,In_548,In_767);
or U1799 (N_1799,In_465,In_240);
or U1800 (N_1800,In_233,In_46);
xor U1801 (N_1801,In_751,In_660);
nor U1802 (N_1802,In_381,In_313);
or U1803 (N_1803,In_290,In_816);
or U1804 (N_1804,In_343,In_186);
nand U1805 (N_1805,In_281,In_217);
and U1806 (N_1806,In_738,In_136);
and U1807 (N_1807,In_419,In_8);
nand U1808 (N_1808,In_254,In_297);
and U1809 (N_1809,In_741,In_854);
or U1810 (N_1810,In_720,In_299);
nor U1811 (N_1811,In_930,In_267);
nor U1812 (N_1812,In_845,In_883);
nand U1813 (N_1813,In_184,In_84);
nor U1814 (N_1814,In_368,In_546);
nand U1815 (N_1815,In_518,In_68);
or U1816 (N_1816,In_177,In_583);
nor U1817 (N_1817,In_112,In_618);
nand U1818 (N_1818,In_33,In_664);
or U1819 (N_1819,In_215,In_95);
nor U1820 (N_1820,In_4,In_500);
and U1821 (N_1821,In_438,In_683);
and U1822 (N_1822,In_32,In_398);
and U1823 (N_1823,In_900,In_542);
nor U1824 (N_1824,In_797,In_342);
nor U1825 (N_1825,In_595,In_577);
and U1826 (N_1826,In_521,In_535);
nand U1827 (N_1827,In_446,In_926);
nand U1828 (N_1828,In_605,In_365);
or U1829 (N_1829,In_779,In_29);
nand U1830 (N_1830,In_571,In_319);
xor U1831 (N_1831,In_892,In_815);
nor U1832 (N_1832,In_178,In_89);
nand U1833 (N_1833,In_5,In_521);
or U1834 (N_1834,In_175,In_760);
and U1835 (N_1835,In_257,In_112);
or U1836 (N_1836,In_864,In_506);
nor U1837 (N_1837,In_137,In_84);
nor U1838 (N_1838,In_955,In_435);
nand U1839 (N_1839,In_814,In_187);
nand U1840 (N_1840,In_1,In_87);
or U1841 (N_1841,In_818,In_397);
or U1842 (N_1842,In_944,In_108);
nor U1843 (N_1843,In_977,In_514);
and U1844 (N_1844,In_222,In_330);
and U1845 (N_1845,In_337,In_372);
and U1846 (N_1846,In_143,In_382);
and U1847 (N_1847,In_529,In_922);
and U1848 (N_1848,In_827,In_446);
nor U1849 (N_1849,In_717,In_260);
and U1850 (N_1850,In_251,In_568);
and U1851 (N_1851,In_964,In_896);
nor U1852 (N_1852,In_2,In_93);
nand U1853 (N_1853,In_539,In_718);
nand U1854 (N_1854,In_918,In_71);
and U1855 (N_1855,In_176,In_996);
nor U1856 (N_1856,In_759,In_347);
or U1857 (N_1857,In_787,In_918);
or U1858 (N_1858,In_387,In_802);
nor U1859 (N_1859,In_809,In_443);
or U1860 (N_1860,In_775,In_730);
nor U1861 (N_1861,In_60,In_368);
or U1862 (N_1862,In_845,In_142);
nor U1863 (N_1863,In_974,In_479);
nand U1864 (N_1864,In_156,In_503);
and U1865 (N_1865,In_775,In_594);
nand U1866 (N_1866,In_874,In_916);
and U1867 (N_1867,In_399,In_794);
nand U1868 (N_1868,In_220,In_453);
nor U1869 (N_1869,In_705,In_245);
nand U1870 (N_1870,In_626,In_666);
and U1871 (N_1871,In_948,In_795);
nor U1872 (N_1872,In_869,In_43);
and U1873 (N_1873,In_868,In_846);
and U1874 (N_1874,In_344,In_589);
nand U1875 (N_1875,In_734,In_693);
nand U1876 (N_1876,In_25,In_577);
nand U1877 (N_1877,In_764,In_839);
nor U1878 (N_1878,In_515,In_595);
or U1879 (N_1879,In_139,In_451);
or U1880 (N_1880,In_385,In_836);
or U1881 (N_1881,In_92,In_926);
or U1882 (N_1882,In_161,In_203);
nand U1883 (N_1883,In_242,In_867);
nor U1884 (N_1884,In_192,In_16);
nand U1885 (N_1885,In_413,In_331);
nor U1886 (N_1886,In_855,In_30);
or U1887 (N_1887,In_29,In_985);
and U1888 (N_1888,In_340,In_890);
or U1889 (N_1889,In_127,In_697);
and U1890 (N_1890,In_273,In_501);
nor U1891 (N_1891,In_846,In_739);
nand U1892 (N_1892,In_500,In_36);
nor U1893 (N_1893,In_743,In_265);
xor U1894 (N_1894,In_763,In_712);
nand U1895 (N_1895,In_435,In_502);
nor U1896 (N_1896,In_589,In_97);
or U1897 (N_1897,In_2,In_998);
nor U1898 (N_1898,In_321,In_591);
nor U1899 (N_1899,In_278,In_913);
and U1900 (N_1900,In_390,In_62);
or U1901 (N_1901,In_673,In_595);
and U1902 (N_1902,In_754,In_56);
nor U1903 (N_1903,In_366,In_162);
or U1904 (N_1904,In_977,In_670);
or U1905 (N_1905,In_115,In_289);
nand U1906 (N_1906,In_407,In_562);
nor U1907 (N_1907,In_458,In_781);
and U1908 (N_1908,In_992,In_296);
or U1909 (N_1909,In_690,In_367);
and U1910 (N_1910,In_711,In_478);
nor U1911 (N_1911,In_437,In_612);
nor U1912 (N_1912,In_361,In_524);
and U1913 (N_1913,In_423,In_584);
nand U1914 (N_1914,In_857,In_465);
nand U1915 (N_1915,In_666,In_622);
nor U1916 (N_1916,In_110,In_26);
nor U1917 (N_1917,In_93,In_992);
nand U1918 (N_1918,In_242,In_713);
nor U1919 (N_1919,In_176,In_797);
and U1920 (N_1920,In_718,In_68);
nor U1921 (N_1921,In_362,In_284);
and U1922 (N_1922,In_548,In_712);
and U1923 (N_1923,In_951,In_597);
nor U1924 (N_1924,In_140,In_68);
nand U1925 (N_1925,In_300,In_36);
nor U1926 (N_1926,In_656,In_425);
nand U1927 (N_1927,In_479,In_547);
or U1928 (N_1928,In_99,In_680);
or U1929 (N_1929,In_142,In_748);
nand U1930 (N_1930,In_807,In_840);
nand U1931 (N_1931,In_164,In_118);
nor U1932 (N_1932,In_130,In_315);
and U1933 (N_1933,In_928,In_443);
or U1934 (N_1934,In_164,In_15);
nor U1935 (N_1935,In_274,In_458);
nand U1936 (N_1936,In_175,In_90);
nand U1937 (N_1937,In_645,In_491);
or U1938 (N_1938,In_966,In_688);
or U1939 (N_1939,In_447,In_788);
or U1940 (N_1940,In_30,In_443);
or U1941 (N_1941,In_424,In_785);
nor U1942 (N_1942,In_287,In_157);
nand U1943 (N_1943,In_689,In_483);
or U1944 (N_1944,In_105,In_534);
nand U1945 (N_1945,In_2,In_528);
nor U1946 (N_1946,In_439,In_553);
nor U1947 (N_1947,In_820,In_809);
nor U1948 (N_1948,In_536,In_473);
nor U1949 (N_1949,In_786,In_907);
or U1950 (N_1950,In_285,In_49);
nand U1951 (N_1951,In_878,In_371);
nor U1952 (N_1952,In_164,In_421);
or U1953 (N_1953,In_144,In_683);
nor U1954 (N_1954,In_8,In_244);
nor U1955 (N_1955,In_887,In_350);
or U1956 (N_1956,In_89,In_678);
and U1957 (N_1957,In_112,In_34);
and U1958 (N_1958,In_574,In_322);
and U1959 (N_1959,In_441,In_800);
or U1960 (N_1960,In_264,In_747);
nor U1961 (N_1961,In_815,In_674);
and U1962 (N_1962,In_973,In_466);
nand U1963 (N_1963,In_939,In_23);
and U1964 (N_1964,In_472,In_236);
nor U1965 (N_1965,In_216,In_343);
nor U1966 (N_1966,In_983,In_741);
nand U1967 (N_1967,In_157,In_889);
and U1968 (N_1968,In_139,In_791);
or U1969 (N_1969,In_504,In_458);
or U1970 (N_1970,In_576,In_539);
and U1971 (N_1971,In_67,In_134);
nor U1972 (N_1972,In_646,In_748);
nand U1973 (N_1973,In_987,In_77);
nor U1974 (N_1974,In_897,In_24);
nand U1975 (N_1975,In_515,In_125);
or U1976 (N_1976,In_396,In_324);
and U1977 (N_1977,In_861,In_653);
and U1978 (N_1978,In_369,In_264);
nor U1979 (N_1979,In_156,In_280);
or U1980 (N_1980,In_227,In_507);
xnor U1981 (N_1981,In_436,In_410);
and U1982 (N_1982,In_812,In_689);
and U1983 (N_1983,In_833,In_440);
and U1984 (N_1984,In_508,In_892);
or U1985 (N_1985,In_671,In_675);
nand U1986 (N_1986,In_482,In_372);
or U1987 (N_1987,In_851,In_890);
nor U1988 (N_1988,In_778,In_919);
or U1989 (N_1989,In_642,In_319);
nor U1990 (N_1990,In_400,In_785);
nor U1991 (N_1991,In_134,In_734);
nand U1992 (N_1992,In_983,In_875);
nand U1993 (N_1993,In_110,In_759);
or U1994 (N_1994,In_589,In_710);
nor U1995 (N_1995,In_470,In_52);
nor U1996 (N_1996,In_809,In_365);
nand U1997 (N_1997,In_408,In_642);
nand U1998 (N_1998,In_91,In_226);
xnor U1999 (N_1999,In_348,In_728);
nand U2000 (N_2000,N_1456,N_1723);
or U2001 (N_2001,N_411,N_402);
nand U2002 (N_2002,N_433,N_23);
nor U2003 (N_2003,N_445,N_1133);
or U2004 (N_2004,N_1236,N_861);
xnor U2005 (N_2005,N_212,N_657);
nand U2006 (N_2006,N_264,N_1654);
or U2007 (N_2007,N_57,N_1614);
and U2008 (N_2008,N_419,N_432);
nand U2009 (N_2009,N_1651,N_1936);
or U2010 (N_2010,N_1288,N_438);
xnor U2011 (N_2011,N_1954,N_590);
and U2012 (N_2012,N_1672,N_564);
nand U2013 (N_2013,N_1246,N_348);
or U2014 (N_2014,N_986,N_8);
nor U2015 (N_2015,N_532,N_1466);
and U2016 (N_2016,N_1960,N_1009);
and U2017 (N_2017,N_450,N_1607);
nor U2018 (N_2018,N_1532,N_759);
nand U2019 (N_2019,N_1568,N_1766);
or U2020 (N_2020,N_1197,N_1241);
nand U2021 (N_2021,N_73,N_887);
nand U2022 (N_2022,N_1116,N_260);
and U2023 (N_2023,N_1036,N_1214);
and U2024 (N_2024,N_1351,N_1294);
or U2025 (N_2025,N_1734,N_1743);
or U2026 (N_2026,N_689,N_32);
or U2027 (N_2027,N_1777,N_454);
and U2028 (N_2028,N_1496,N_701);
nor U2029 (N_2029,N_1562,N_725);
or U2030 (N_2030,N_1567,N_124);
nand U2031 (N_2031,N_386,N_601);
nand U2032 (N_2032,N_1634,N_1015);
and U2033 (N_2033,N_1978,N_525);
or U2034 (N_2034,N_1038,N_1268);
nand U2035 (N_2035,N_1608,N_681);
or U2036 (N_2036,N_1367,N_153);
and U2037 (N_2037,N_1691,N_1625);
or U2038 (N_2038,N_1779,N_847);
or U2039 (N_2039,N_731,N_1179);
or U2040 (N_2040,N_1517,N_279);
and U2041 (N_2041,N_1098,N_739);
or U2042 (N_2042,N_1760,N_1878);
or U2043 (N_2043,N_453,N_206);
or U2044 (N_2044,N_1077,N_1257);
nor U2045 (N_2045,N_1836,N_545);
nor U2046 (N_2046,N_1000,N_1380);
or U2047 (N_2047,N_1492,N_918);
nand U2048 (N_2048,N_1850,N_1443);
nor U2049 (N_2049,N_479,N_1021);
nor U2050 (N_2050,N_1315,N_219);
xor U2051 (N_2051,N_1928,N_553);
or U2052 (N_2052,N_742,N_1353);
or U2053 (N_2053,N_458,N_435);
nor U2054 (N_2054,N_1616,N_1992);
nor U2055 (N_2055,N_1307,N_224);
or U2056 (N_2056,N_1363,N_877);
or U2057 (N_2057,N_334,N_1172);
nor U2058 (N_2058,N_888,N_1627);
nor U2059 (N_2059,N_785,N_2);
nand U2060 (N_2060,N_608,N_188);
or U2061 (N_2061,N_1995,N_1054);
nand U2062 (N_2062,N_1925,N_1695);
nand U2063 (N_2063,N_697,N_1579);
nand U2064 (N_2064,N_145,N_449);
and U2065 (N_2065,N_794,N_710);
nor U2066 (N_2066,N_1907,N_1153);
nor U2067 (N_2067,N_31,N_1684);
nor U2068 (N_2068,N_1096,N_614);
or U2069 (N_2069,N_1027,N_1780);
nand U2070 (N_2070,N_492,N_65);
or U2071 (N_2071,N_651,N_1285);
and U2072 (N_2072,N_1822,N_754);
and U2073 (N_2073,N_974,N_1437);
or U2074 (N_2074,N_586,N_838);
or U2075 (N_2075,N_829,N_753);
nand U2076 (N_2076,N_1430,N_985);
and U2077 (N_2077,N_15,N_71);
and U2078 (N_2078,N_1377,N_159);
nand U2079 (N_2079,N_598,N_1753);
xnor U2080 (N_2080,N_957,N_373);
or U2081 (N_2081,N_14,N_1180);
nor U2082 (N_2082,N_1089,N_142);
nand U2083 (N_2083,N_782,N_854);
nand U2084 (N_2084,N_883,N_497);
nor U2085 (N_2085,N_685,N_610);
nor U2086 (N_2086,N_975,N_592);
or U2087 (N_2087,N_1170,N_1208);
or U2088 (N_2088,N_1427,N_1795);
nand U2089 (N_2089,N_254,N_997);
nand U2090 (N_2090,N_851,N_1313);
xor U2091 (N_2091,N_1452,N_1768);
or U2092 (N_2092,N_104,N_95);
nand U2093 (N_2093,N_240,N_1258);
nand U2094 (N_2094,N_626,N_1201);
or U2095 (N_2095,N_1174,N_1609);
and U2096 (N_2096,N_1410,N_1716);
nor U2097 (N_2097,N_305,N_835);
and U2098 (N_2098,N_1516,N_283);
nor U2099 (N_2099,N_1722,N_1647);
nand U2100 (N_2100,N_319,N_1896);
nand U2101 (N_2101,N_1524,N_1886);
nand U2102 (N_2102,N_815,N_728);
and U2103 (N_2103,N_619,N_434);
or U2104 (N_2104,N_1439,N_1699);
and U2105 (N_2105,N_1053,N_267);
and U2106 (N_2106,N_834,N_331);
nor U2107 (N_2107,N_155,N_1185);
nand U2108 (N_2108,N_1321,N_182);
and U2109 (N_2109,N_79,N_366);
or U2110 (N_2110,N_1937,N_1655);
nor U2111 (N_2111,N_857,N_825);
or U2112 (N_2112,N_1704,N_1838);
or U2113 (N_2113,N_1227,N_370);
nor U2114 (N_2114,N_583,N_580);
or U2115 (N_2115,N_674,N_646);
nand U2116 (N_2116,N_88,N_396);
nor U2117 (N_2117,N_1047,N_459);
xnor U2118 (N_2118,N_1057,N_1113);
nor U2119 (N_2119,N_1088,N_1093);
or U2120 (N_2120,N_1166,N_100);
nor U2121 (N_2121,N_168,N_539);
and U2122 (N_2122,N_1973,N_1981);
nand U2123 (N_2123,N_549,N_1013);
or U2124 (N_2124,N_1479,N_536);
and U2125 (N_2125,N_1656,N_1284);
nand U2126 (N_2126,N_72,N_636);
nand U2127 (N_2127,N_889,N_746);
or U2128 (N_2128,N_924,N_1518);
and U2129 (N_2129,N_1677,N_66);
nor U2130 (N_2130,N_650,N_132);
nand U2131 (N_2131,N_784,N_1248);
nand U2132 (N_2132,N_620,N_734);
or U2133 (N_2133,N_1551,N_578);
and U2134 (N_2134,N_1167,N_1163);
or U2135 (N_2135,N_358,N_919);
or U2136 (N_2136,N_1260,N_1793);
or U2137 (N_2137,N_1191,N_1228);
nor U2138 (N_2138,N_290,N_302);
nor U2139 (N_2139,N_477,N_1323);
and U2140 (N_2140,N_47,N_484);
or U2141 (N_2141,N_1824,N_1661);
nand U2142 (N_2142,N_171,N_486);
nand U2143 (N_2143,N_1948,N_1868);
and U2144 (N_2144,N_75,N_1792);
or U2145 (N_2145,N_1,N_916);
and U2146 (N_2146,N_1557,N_1658);
nand U2147 (N_2147,N_1306,N_467);
or U2148 (N_2148,N_695,N_1339);
nor U2149 (N_2149,N_1788,N_347);
and U2150 (N_2150,N_1223,N_29);
and U2151 (N_2151,N_481,N_1271);
nand U2152 (N_2152,N_1225,N_1342);
nor U2153 (N_2153,N_355,N_1933);
nand U2154 (N_2154,N_1891,N_900);
nand U2155 (N_2155,N_1305,N_647);
nand U2156 (N_2156,N_1388,N_382);
nand U2157 (N_2157,N_1597,N_1066);
or U2158 (N_2158,N_134,N_801);
nor U2159 (N_2159,N_663,N_472);
nor U2160 (N_2160,N_1657,N_711);
and U2161 (N_2161,N_1650,N_1909);
nand U2162 (N_2162,N_664,N_1414);
or U2163 (N_2163,N_365,N_360);
or U2164 (N_2164,N_1890,N_1359);
nand U2165 (N_2165,N_1150,N_228);
or U2166 (N_2166,N_1952,N_716);
nand U2167 (N_2167,N_1611,N_1527);
nor U2168 (N_2168,N_1571,N_1504);
and U2169 (N_2169,N_1846,N_1026);
and U2170 (N_2170,N_1593,N_1690);
or U2171 (N_2171,N_275,N_117);
nand U2172 (N_2172,N_27,N_77);
and U2173 (N_2173,N_504,N_1964);
and U2174 (N_2174,N_771,N_1697);
and U2175 (N_2175,N_138,N_1253);
nand U2176 (N_2176,N_624,N_1441);
nand U2177 (N_2177,N_788,N_426);
nand U2178 (N_2178,N_1635,N_740);
nand U2179 (N_2179,N_1478,N_1999);
and U2180 (N_2180,N_705,N_766);
nor U2181 (N_2181,N_1195,N_1485);
nor U2182 (N_2182,N_589,N_520);
and U2183 (N_2183,N_1162,N_1622);
and U2184 (N_2184,N_1512,N_1087);
nor U2185 (N_2185,N_1598,N_869);
nand U2186 (N_2186,N_495,N_1786);
and U2187 (N_2187,N_1880,N_1408);
or U2188 (N_2188,N_1979,N_1790);
nand U2189 (N_2189,N_519,N_1636);
nor U2190 (N_2190,N_1942,N_522);
nand U2191 (N_2191,N_491,N_1910);
nor U2192 (N_2192,N_896,N_1784);
nand U2193 (N_2193,N_1075,N_1887);
nand U2194 (N_2194,N_1894,N_409);
nand U2195 (N_2195,N_541,N_1375);
nand U2196 (N_2196,N_19,N_1633);
nor U2197 (N_2197,N_747,N_855);
nor U2198 (N_2198,N_1210,N_1052);
or U2199 (N_2199,N_1537,N_461);
nand U2200 (N_2200,N_1619,N_1831);
nor U2201 (N_2201,N_1728,N_908);
nor U2202 (N_2202,N_1433,N_242);
and U2203 (N_2203,N_871,N_1549);
xor U2204 (N_2204,N_346,N_4);
nor U2205 (N_2205,N_556,N_1930);
nand U2206 (N_2206,N_707,N_143);
nor U2207 (N_2207,N_1024,N_1807);
or U2208 (N_2208,N_1381,N_1854);
or U2209 (N_2209,N_1624,N_1333);
nor U2210 (N_2210,N_1461,N_1368);
and U2211 (N_2211,N_1161,N_1319);
nor U2212 (N_2212,N_92,N_1261);
or U2213 (N_2213,N_1142,N_1781);
nor U2214 (N_2214,N_1175,N_289);
or U2215 (N_2215,N_1763,N_1346);
nand U2216 (N_2216,N_200,N_1233);
nand U2217 (N_2217,N_251,N_414);
and U2218 (N_2218,N_727,N_1095);
and U2219 (N_2219,N_687,N_1159);
or U2220 (N_2220,N_616,N_1529);
nand U2221 (N_2221,N_136,N_327);
or U2222 (N_2222,N_1758,N_1639);
and U2223 (N_2223,N_1269,N_87);
nor U2224 (N_2224,N_485,N_356);
or U2225 (N_2225,N_1188,N_907);
nor U2226 (N_2226,N_1975,N_991);
nand U2227 (N_2227,N_44,N_508);
nand U2228 (N_2228,N_1812,N_1299);
nor U2229 (N_2229,N_1630,N_1546);
or U2230 (N_2230,N_34,N_1139);
nand U2231 (N_2231,N_530,N_1957);
nor U2232 (N_2232,N_1971,N_10);
nor U2233 (N_2233,N_934,N_169);
nor U2234 (N_2234,N_107,N_1901);
nor U2235 (N_2235,N_1314,N_1158);
and U2236 (N_2236,N_118,N_1031);
nand U2237 (N_2237,N_1666,N_1502);
nand U2238 (N_2238,N_1757,N_1705);
and U2239 (N_2239,N_1062,N_533);
nand U2240 (N_2240,N_42,N_550);
nand U2241 (N_2241,N_1435,N_587);
nor U2242 (N_2242,N_82,N_554);
nand U2243 (N_2243,N_712,N_170);
and U2244 (N_2244,N_1984,N_312);
and U2245 (N_2245,N_1500,N_670);
nand U2246 (N_2246,N_723,N_548);
or U2247 (N_2247,N_1157,N_1827);
nor U2248 (N_2248,N_1732,N_1085);
and U2249 (N_2249,N_1458,N_1645);
or U2250 (N_2250,N_1640,N_1004);
or U2251 (N_2251,N_89,N_1395);
nand U2252 (N_2252,N_1097,N_904);
or U2253 (N_2253,N_1869,N_154);
nand U2254 (N_2254,N_421,N_547);
nand U2255 (N_2255,N_1164,N_1130);
nor U2256 (N_2256,N_1545,N_1450);
nor U2257 (N_2257,N_194,N_1415);
nand U2258 (N_2258,N_654,N_1371);
nand U2259 (N_2259,N_1023,N_1821);
and U2260 (N_2260,N_1472,N_1224);
or U2261 (N_2261,N_645,N_992);
nand U2262 (N_2262,N_1962,N_1751);
nor U2263 (N_2263,N_330,N_1421);
and U2264 (N_2264,N_769,N_1349);
nand U2265 (N_2265,N_1550,N_535);
nor U2266 (N_2266,N_1686,N_637);
or U2267 (N_2267,N_469,N_1362);
nand U2268 (N_2268,N_85,N_1376);
and U2269 (N_2269,N_1839,N_1570);
nand U2270 (N_2270,N_860,N_959);
or U2271 (N_2271,N_127,N_1037);
nor U2272 (N_2272,N_1345,N_938);
nand U2273 (N_2273,N_81,N_229);
and U2274 (N_2274,N_1426,N_37);
nand U2275 (N_2275,N_1033,N_1365);
nand U2276 (N_2276,N_678,N_777);
or U2277 (N_2277,N_466,N_1470);
nand U2278 (N_2278,N_1542,N_1382);
nor U2279 (N_2279,N_597,N_1219);
or U2280 (N_2280,N_822,N_1772);
and U2281 (N_2281,N_1252,N_76);
or U2282 (N_2282,N_1638,N_1515);
or U2283 (N_2283,N_1112,N_1741);
nor U2284 (N_2284,N_572,N_1072);
or U2285 (N_2285,N_1444,N_756);
nor U2286 (N_2286,N_1950,N_537);
or U2287 (N_2287,N_1276,N_1584);
nand U2288 (N_2288,N_186,N_1914);
nor U2289 (N_2289,N_377,N_571);
and U2290 (N_2290,N_1538,N_634);
or U2291 (N_2291,N_179,N_677);
nand U2292 (N_2292,N_828,N_962);
nand U2293 (N_2293,N_1673,N_557);
and U2294 (N_2294,N_1182,N_1463);
and U2295 (N_2295,N_1264,N_1561);
nor U2296 (N_2296,N_1857,N_1663);
or U2297 (N_2297,N_611,N_146);
and U2298 (N_2298,N_973,N_909);
and U2299 (N_2299,N_802,N_1211);
nor U2300 (N_2300,N_1509,N_1423);
or U2301 (N_2301,N_425,N_1966);
and U2302 (N_2302,N_816,N_1165);
or U2303 (N_2303,N_25,N_679);
nor U2304 (N_2304,N_1863,N_1132);
and U2305 (N_2305,N_1671,N_1249);
and U2306 (N_2306,N_1767,N_1387);
nor U2307 (N_2307,N_1533,N_1856);
or U2308 (N_2308,N_790,N_1669);
or U2309 (N_2309,N_1724,N_1416);
nand U2310 (N_2310,N_9,N_846);
nor U2311 (N_2311,N_721,N_427);
nor U2312 (N_2312,N_776,N_1540);
nor U2313 (N_2313,N_499,N_1316);
nand U2314 (N_2314,N_227,N_1070);
nand U2315 (N_2315,N_666,N_1621);
and U2316 (N_2316,N_948,N_1370);
nand U2317 (N_2317,N_1255,N_1017);
nand U2318 (N_2318,N_686,N_1424);
nand U2319 (N_2319,N_1895,N_706);
nor U2320 (N_2320,N_653,N_609);
or U2321 (N_2321,N_139,N_691);
and U2322 (N_2322,N_1006,N_531);
or U2323 (N_2323,N_1393,N_1587);
nor U2324 (N_2324,N_713,N_1577);
nand U2325 (N_2325,N_898,N_1446);
or U2326 (N_2326,N_1727,N_1733);
and U2327 (N_2327,N_1646,N_294);
nor U2328 (N_2328,N_30,N_884);
nand U2329 (N_2329,N_199,N_881);
or U2330 (N_2330,N_1069,N_1385);
nor U2331 (N_2331,N_595,N_1254);
and U2332 (N_2332,N_1216,N_1325);
or U2333 (N_2333,N_1591,N_446);
nor U2334 (N_2334,N_1202,N_245);
or U2335 (N_2335,N_131,N_755);
and U2336 (N_2336,N_462,N_1875);
nand U2337 (N_2337,N_70,N_394);
and U2338 (N_2338,N_791,N_1858);
or U2339 (N_2339,N_1800,N_464);
nor U2340 (N_2340,N_671,N_367);
and U2341 (N_2341,N_503,N_999);
and U2342 (N_2342,N_428,N_488);
or U2343 (N_2343,N_1056,N_872);
nor U2344 (N_2344,N_936,N_1776);
nand U2345 (N_2345,N_830,N_915);
and U2346 (N_2346,N_1696,N_950);
nand U2347 (N_2347,N_201,N_1469);
nor U2348 (N_2348,N_383,N_501);
nand U2349 (N_2349,N_996,N_960);
or U2350 (N_2350,N_783,N_1744);
nand U2351 (N_2351,N_1837,N_1338);
or U2352 (N_2352,N_287,N_86);
or U2353 (N_2353,N_588,N_1694);
nor U2354 (N_2354,N_1468,N_1337);
or U2355 (N_2355,N_209,N_1553);
or U2356 (N_2356,N_106,N_593);
or U2357 (N_2357,N_1281,N_1231);
and U2358 (N_2358,N_406,N_803);
nand U2359 (N_2359,N_1808,N_927);
nor U2360 (N_2360,N_1402,N_1110);
and U2361 (N_2361,N_1620,N_1399);
nor U2362 (N_2362,N_630,N_5);
nand U2363 (N_2363,N_1143,N_1022);
or U2364 (N_2364,N_1632,N_1422);
nand U2365 (N_2365,N_1756,N_1154);
nand U2366 (N_2366,N_1580,N_84);
nand U2367 (N_2367,N_187,N_208);
or U2368 (N_2368,N_112,N_1046);
nand U2369 (N_2369,N_596,N_281);
nor U2370 (N_2370,N_845,N_844);
nor U2371 (N_2371,N_125,N_1340);
nand U2372 (N_2372,N_54,N_1302);
nor U2373 (N_2373,N_1643,N_998);
nand U2374 (N_2374,N_239,N_848);
and U2375 (N_2375,N_473,N_1924);
or U2376 (N_2376,N_1637,N_489);
nand U2377 (N_2377,N_880,N_780);
nand U2378 (N_2378,N_1711,N_1406);
nor U2379 (N_2379,N_318,N_1523);
nor U2380 (N_2380,N_1592,N_853);
nor U2381 (N_2381,N_910,N_1754);
nor U2382 (N_2382,N_817,N_1477);
nand U2383 (N_2383,N_863,N_352);
nor U2384 (N_2384,N_980,N_1938);
or U2385 (N_2385,N_412,N_1358);
nor U2386 (N_2386,N_1105,N_1566);
or U2387 (N_2387,N_1662,N_758);
nand U2388 (N_2388,N_1117,N_16);
or U2389 (N_2389,N_1169,N_388);
or U2390 (N_2390,N_837,N_510);
nand U2391 (N_2391,N_1953,N_726);
nor U2392 (N_2392,N_652,N_717);
xor U2393 (N_2393,N_41,N_841);
nand U2394 (N_2394,N_1731,N_1932);
and U2395 (N_2395,N_1206,N_1042);
or U2396 (N_2396,N_1149,N_1604);
or U2397 (N_2397,N_988,N_234);
and U2398 (N_2398,N_1121,N_1360);
and U2399 (N_2399,N_603,N_1140);
nor U2400 (N_2400,N_527,N_437);
nor U2401 (N_2401,N_990,N_165);
nand U2402 (N_2402,N_399,N_604);
nand U2403 (N_2403,N_1060,N_1573);
and U2404 (N_2404,N_983,N_1802);
and U2405 (N_2405,N_369,N_1081);
xnor U2406 (N_2406,N_1151,N_658);
nor U2407 (N_2407,N_1606,N_225);
nand U2408 (N_2408,N_1974,N_1934);
nand U2409 (N_2409,N_53,N_271);
and U2410 (N_2410,N_1785,N_1805);
and U2411 (N_2411,N_204,N_172);
and U2412 (N_2412,N_576,N_475);
nand U2413 (N_2413,N_1204,N_995);
nor U2414 (N_2414,N_137,N_339);
or U2415 (N_2415,N_1526,N_1407);
or U2416 (N_2416,N_529,N_672);
or U2417 (N_2417,N_296,N_929);
nor U2418 (N_2418,N_220,N_190);
and U2419 (N_2419,N_476,N_509);
nor U2420 (N_2420,N_833,N_600);
and U2421 (N_2421,N_1670,N_43);
nand U2422 (N_2422,N_751,N_1687);
or U2423 (N_2423,N_966,N_1816);
or U2424 (N_2424,N_625,N_1138);
nor U2425 (N_2425,N_1941,N_615);
and U2426 (N_2426,N_633,N_1915);
or U2427 (N_2427,N_585,N_393);
and U2428 (N_2428,N_1109,N_1397);
nor U2429 (N_2429,N_1676,N_984);
or U2430 (N_2430,N_1002,N_255);
nor U2431 (N_2431,N_1083,N_1730);
and U2432 (N_2432,N_304,N_252);
or U2433 (N_2433,N_1798,N_133);
or U2434 (N_2434,N_818,N_613);
or U2435 (N_2435,N_856,N_268);
nor U2436 (N_2436,N_507,N_1156);
and U2437 (N_2437,N_1243,N_876);
and U2438 (N_2438,N_873,N_1303);
nor U2439 (N_2439,N_431,N_1289);
nor U2440 (N_2440,N_1374,N_1575);
nand U2441 (N_2441,N_1521,N_1475);
and U2442 (N_2442,N_668,N_805);
nor U2443 (N_2443,N_185,N_1882);
or U2444 (N_2444,N_1187,N_1976);
and U2445 (N_2445,N_1679,N_1739);
nand U2446 (N_2446,N_878,N_1605);
and U2447 (N_2447,N_982,N_135);
nor U2448 (N_2448,N_1209,N_1877);
nand U2449 (N_2449,N_528,N_457);
nand U2450 (N_2450,N_1865,N_116);
xor U2451 (N_2451,N_1811,N_1355);
and U2452 (N_2452,N_511,N_521);
nand U2453 (N_2453,N_1725,N_111);
or U2454 (N_2454,N_789,N_364);
nor U2455 (N_2455,N_1438,N_1912);
nor U2456 (N_2456,N_444,N_1683);
nor U2457 (N_2457,N_836,N_178);
and U2458 (N_2458,N_1107,N_1213);
and U2459 (N_2459,N_1205,N_774);
nor U2460 (N_2460,N_892,N_420);
nand U2461 (N_2461,N_1350,N_94);
and U2462 (N_2462,N_291,N_979);
nand U2463 (N_2463,N_1445,N_961);
and U2464 (N_2464,N_90,N_1762);
nor U2465 (N_2465,N_494,N_78);
or U2466 (N_2466,N_1840,N_1124);
nand U2467 (N_2467,N_1775,N_628);
xor U2468 (N_2468,N_7,N_1278);
nor U2469 (N_2469,N_1797,N_429);
or U2470 (N_2470,N_1250,N_384);
nor U2471 (N_2471,N_1996,N_413);
nor U2472 (N_2472,N_1554,N_690);
or U2473 (N_2473,N_1931,N_28);
nand U2474 (N_2474,N_946,N_558);
and U2475 (N_2475,N_1834,N_1789);
nand U2476 (N_2476,N_534,N_269);
and U2477 (N_2477,N_993,N_1883);
nor U2478 (N_2478,N_1530,N_1823);
nand U2479 (N_2479,N_1011,N_1576);
nor U2480 (N_2480,N_1983,N_1746);
and U2481 (N_2481,N_978,N_902);
nor U2482 (N_2482,N_248,N_729);
nor U2483 (N_2483,N_1487,N_1310);
and U2484 (N_2484,N_417,N_708);
and U2485 (N_2485,N_1674,N_971);
or U2486 (N_2486,N_490,N_213);
xnor U2487 (N_2487,N_1127,N_256);
and U2488 (N_2488,N_1879,N_602);
nand U2489 (N_2489,N_932,N_584);
or U2490 (N_2490,N_448,N_972);
nor U2491 (N_2491,N_1552,N_235);
nand U2492 (N_2492,N_923,N_343);
nand U2493 (N_2493,N_123,N_1943);
or U2494 (N_2494,N_1588,N_442);
and U2495 (N_2495,N_441,N_1970);
or U2496 (N_2496,N_233,N_1084);
or U2497 (N_2497,N_885,N_1090);
and U2498 (N_2498,N_1301,N_1274);
nand U2499 (N_2499,N_1238,N_1495);
and U2500 (N_2500,N_1326,N_575);
nand U2501 (N_2501,N_1872,N_309);
nand U2502 (N_2502,N_901,N_1327);
or U2503 (N_2503,N_1612,N_760);
nor U2504 (N_2504,N_1270,N_11);
and U2505 (N_2505,N_195,N_565);
nand U2506 (N_2506,N_763,N_1356);
and U2507 (N_2507,N_618,N_1404);
and U2508 (N_2508,N_1900,N_1290);
or U2509 (N_2509,N_744,N_40);
and U2510 (N_2510,N_1898,N_714);
or U2511 (N_2511,N_792,N_1578);
nor U2512 (N_2512,N_1372,N_102);
or U2513 (N_2513,N_389,N_317);
and U2514 (N_2514,N_308,N_1644);
or U2515 (N_2515,N_45,N_1405);
nor U2516 (N_2516,N_612,N_1688);
or U2517 (N_2517,N_1594,N_390);
or U2518 (N_2518,N_1177,N_1714);
nand U2519 (N_2519,N_1918,N_307);
nor U2520 (N_2520,N_381,N_404);
or U2521 (N_2521,N_1417,N_1300);
or U2522 (N_2522,N_1548,N_175);
nand U2523 (N_2523,N_121,N_483);
nor U2524 (N_2524,N_920,N_1884);
nand U2525 (N_2525,N_1226,N_850);
or U2526 (N_2526,N_1431,N_840);
nand U2527 (N_2527,N_917,N_243);
xor U2528 (N_2528,N_1759,N_814);
nor U2529 (N_2529,N_276,N_768);
and U2530 (N_2530,N_1409,N_544);
nand U2531 (N_2531,N_694,N_1520);
nand U2532 (N_2532,N_1851,N_1222);
or U2533 (N_2533,N_262,N_1825);
and U2534 (N_2534,N_669,N_1968);
or U2535 (N_2535,N_1184,N_894);
and U2536 (N_2536,N_958,N_865);
and U2537 (N_2537,N_1813,N_60);
nor U2538 (N_2538,N_105,N_342);
nand U2539 (N_2539,N_591,N_749);
nor U2540 (N_2540,N_247,N_743);
or U2541 (N_2541,N_1160,N_500);
or U2542 (N_2542,N_1428,N_1379);
or U2543 (N_2543,N_1985,N_63);
nor U2544 (N_2544,N_258,N_64);
nor U2545 (N_2545,N_362,N_1357);
nor U2546 (N_2546,N_831,N_368);
or U2547 (N_2547,N_676,N_987);
or U2548 (N_2548,N_1710,N_1599);
nand U2549 (N_2549,N_724,N_1459);
and U2550 (N_2550,N_222,N_324);
nor U2551 (N_2551,N_1993,N_284);
or U2552 (N_2552,N_156,N_843);
or U2553 (N_2553,N_1929,N_1860);
nand U2554 (N_2554,N_1432,N_1481);
nor U2555 (N_2555,N_196,N_897);
nor U2556 (N_2556,N_354,N_1086);
nand U2557 (N_2557,N_879,N_1425);
or U2558 (N_2558,N_1221,N_1448);
and U2559 (N_2559,N_1008,N_1787);
and U2560 (N_2560,N_20,N_1990);
and U2561 (N_2561,N_1944,N_1806);
nand U2562 (N_2562,N_517,N_1764);
or U2563 (N_2563,N_141,N_767);
nand U2564 (N_2564,N_1920,N_1708);
nor U2565 (N_2565,N_1955,N_266);
nor U2566 (N_2566,N_1641,N_12);
and U2567 (N_2567,N_286,N_523);
nor U2568 (N_2568,N_667,N_1455);
and U2569 (N_2569,N_1675,N_1178);
nand U2570 (N_2570,N_895,N_1510);
nand U2571 (N_2571,N_1297,N_1080);
or U2572 (N_2572,N_1596,N_1659);
nor U2573 (N_2573,N_1859,N_1242);
nand U2574 (N_2574,N_1118,N_292);
nand U2575 (N_2575,N_1967,N_1718);
or U2576 (N_2576,N_736,N_1262);
and U2577 (N_2577,N_218,N_956);
or U2578 (N_2578,N_311,N_632);
nand U2579 (N_2579,N_50,N_478);
or U2580 (N_2580,N_1074,N_1010);
nand U2581 (N_2581,N_1652,N_1040);
or U2582 (N_2582,N_1146,N_1122);
or U2583 (N_2583,N_567,N_568);
nor U2584 (N_2584,N_954,N_1283);
nor U2585 (N_2585,N_1508,N_1335);
nor U2586 (N_2586,N_1012,N_1791);
nor U2587 (N_2587,N_313,N_480);
nor U2588 (N_2588,N_157,N_1199);
and U2589 (N_2589,N_1911,N_273);
and U2590 (N_2590,N_376,N_989);
xnor U2591 (N_2591,N_1702,N_719);
or U2592 (N_2592,N_977,N_439);
and U2593 (N_2593,N_1501,N_1750);
or U2594 (N_2594,N_238,N_1665);
and U2595 (N_2595,N_379,N_1092);
and U2596 (N_2596,N_207,N_1876);
nor U2597 (N_2597,N_1841,N_1873);
and U2598 (N_2598,N_1803,N_1043);
and U2599 (N_2599,N_1847,N_704);
and U2600 (N_2600,N_1005,N_1603);
nor U2601 (N_2601,N_819,N_810);
and U2602 (N_2602,N_397,N_378);
nand U2603 (N_2603,N_150,N_1473);
or U2604 (N_2604,N_1001,N_1332);
and U2605 (N_2605,N_867,N_513);
or U2606 (N_2606,N_1778,N_1623);
nand U2607 (N_2607,N_849,N_91);
nor U2608 (N_2608,N_1531,N_675);
and U2609 (N_2609,N_1480,N_1927);
nor U2610 (N_2610,N_1558,N_173);
and U2611 (N_2611,N_1308,N_471);
nand U2612 (N_2612,N_935,N_1522);
and U2613 (N_2613,N_1678,N_1881);
and U2614 (N_2614,N_665,N_804);
or U2615 (N_2615,N_336,N_424);
nor U2616 (N_2616,N_1352,N_1101);
or U2617 (N_2617,N_1528,N_1343);
and U2618 (N_2618,N_1864,N_1078);
nand U2619 (N_2619,N_52,N_1899);
and U2620 (N_2620,N_1835,N_144);
nor U2621 (N_2621,N_1701,N_1239);
nand U2622 (N_2622,N_944,N_272);
or U2623 (N_2623,N_344,N_74);
or U2624 (N_2624,N_931,N_1273);
nand U2625 (N_2625,N_1212,N_1245);
nor U2626 (N_2626,N_322,N_551);
and U2627 (N_2627,N_1689,N_303);
or U2628 (N_2628,N_1503,N_1462);
and U2629 (N_2629,N_177,N_49);
nand U2630 (N_2630,N_474,N_1190);
nor U2631 (N_2631,N_216,N_237);
nor U2632 (N_2632,N_1513,N_928);
or U2633 (N_2633,N_1293,N_968);
or U2634 (N_2634,N_1324,N_67);
nor U2635 (N_2635,N_13,N_1392);
nor U2636 (N_2636,N_278,N_1749);
nor U2637 (N_2637,N_1770,N_809);
nor U2638 (N_2638,N_436,N_1296);
nor U2639 (N_2639,N_1347,N_372);
nor U2640 (N_2640,N_298,N_1506);
or U2641 (N_2641,N_1988,N_823);
or U2642 (N_2642,N_18,N_524);
nor U2643 (N_2643,N_361,N_1247);
nand U2644 (N_2644,N_732,N_1680);
and U2645 (N_2645,N_905,N_1099);
nor U2646 (N_2646,N_1103,N_1007);
and U2647 (N_2647,N_217,N_1144);
or U2648 (N_2648,N_1707,N_1064);
nand U2649 (N_2649,N_1519,N_1574);
nand U2650 (N_2650,N_59,N_101);
nor U2651 (N_2651,N_1980,N_109);
or U2652 (N_2652,N_1145,N_947);
or U2653 (N_2653,N_577,N_148);
nor U2654 (N_2654,N_48,N_174);
nor U2655 (N_2655,N_796,N_1949);
nand U2656 (N_2656,N_215,N_1765);
and U2657 (N_2657,N_1555,N_1493);
nor U2658 (N_2658,N_1141,N_1600);
or U2659 (N_2659,N_1713,N_1003);
or U2660 (N_2660,N_1498,N_696);
or U2661 (N_2661,N_899,N_1390);
nor U2662 (N_2662,N_93,N_332);
nand U2663 (N_2663,N_97,N_1100);
and U2664 (N_2664,N_265,N_698);
and U2665 (N_2665,N_408,N_1998);
or U2666 (N_2666,N_1067,N_1457);
nor U2667 (N_2667,N_569,N_120);
or U2668 (N_2668,N_1735,N_1063);
and U2669 (N_2669,N_1065,N_1820);
and U2670 (N_2670,N_244,N_1048);
or U2671 (N_2671,N_1071,N_231);
nor U2672 (N_2672,N_230,N_1685);
nor U2673 (N_2673,N_55,N_1035);
and U2674 (N_2674,N_1511,N_737);
nand U2675 (N_2675,N_594,N_733);
and U2676 (N_2676,N_1491,N_320);
nor U2677 (N_2677,N_410,N_648);
nand U2678 (N_2678,N_661,N_570);
or U2679 (N_2679,N_1277,N_1369);
and U2680 (N_2680,N_660,N_191);
nand U2681 (N_2681,N_1842,N_128);
and U2682 (N_2682,N_942,N_1693);
or U2683 (N_2683,N_80,N_1041);
nor U2684 (N_2684,N_913,N_566);
and U2685 (N_2685,N_1922,N_1965);
nor U2686 (N_2686,N_1908,N_1488);
nand U2687 (N_2687,N_1581,N_1698);
nand U2688 (N_2688,N_1050,N_1945);
and U2689 (N_2689,N_1874,N_692);
and U2690 (N_2690,N_852,N_1391);
nor U2691 (N_2691,N_821,N_210);
or U2692 (N_2692,N_149,N_259);
nand U2693 (N_2693,N_46,N_192);
nor U2694 (N_2694,N_543,N_1994);
or U2695 (N_2695,N_1460,N_1344);
and U2696 (N_2696,N_1401,N_1505);
or U2697 (N_2697,N_405,N_874);
and U2698 (N_2698,N_189,N_1830);
nor U2699 (N_2699,N_812,N_1796);
and U2700 (N_2700,N_58,N_316);
and U2701 (N_2701,N_1218,N_1181);
or U2702 (N_2702,N_1986,N_1411);
nor U2703 (N_2703,N_0,N_1715);
and U2704 (N_2704,N_221,N_582);
nor U2705 (N_2705,N_69,N_1709);
nand U2706 (N_2706,N_1987,N_1464);
nand U2707 (N_2707,N_114,N_398);
and U2708 (N_2708,N_1018,N_781);
nand U2709 (N_2709,N_1913,N_1068);
or U2710 (N_2710,N_1499,N_456);
and U2711 (N_2711,N_1155,N_606);
nand U2712 (N_2712,N_526,N_516);
nor U2713 (N_2713,N_353,N_176);
nand U2714 (N_2714,N_644,N_1617);
and U2715 (N_2715,N_338,N_1094);
or U2716 (N_2716,N_1280,N_1186);
nor U2717 (N_2717,N_1189,N_1320);
or U2718 (N_2718,N_181,N_1586);
nor U2719 (N_2719,N_198,N_1171);
and U2720 (N_2720,N_68,N_1809);
nor U2721 (N_2721,N_232,N_193);
and U2722 (N_2722,N_1436,N_1176);
nand U2723 (N_2723,N_463,N_579);
nand U2724 (N_2724,N_939,N_323);
or U2725 (N_2725,N_1721,N_1585);
and U2726 (N_2726,N_720,N_1681);
nor U2727 (N_2727,N_460,N_487);
or U2728 (N_2728,N_371,N_773);
and U2729 (N_2729,N_357,N_953);
and U2730 (N_2730,N_1489,N_807);
nor U2731 (N_2731,N_709,N_1590);
nand U2732 (N_2732,N_310,N_1341);
and U2733 (N_2733,N_1736,N_1547);
and U2734 (N_2734,N_1849,N_321);
xor U2735 (N_2735,N_295,N_778);
nand U2736 (N_2736,N_1569,N_1152);
nand U2737 (N_2737,N_798,N_799);
or U2738 (N_2738,N_1719,N_518);
or U2739 (N_2739,N_455,N_864);
nand U2740 (N_2740,N_797,N_1137);
or U2741 (N_2741,N_482,N_748);
or U2742 (N_2742,N_119,N_787);
and U2743 (N_2743,N_643,N_1853);
and U2744 (N_2744,N_1329,N_1168);
and U2745 (N_2745,N_793,N_515);
nand U2746 (N_2746,N_1761,N_1667);
and U2747 (N_2747,N_282,N_418);
nand U2748 (N_2748,N_1649,N_981);
nand U2749 (N_2749,N_1128,N_1400);
nand U2750 (N_2750,N_1818,N_1304);
and U2751 (N_2751,N_683,N_1742);
or U2752 (N_2752,N_1729,N_1773);
nand U2753 (N_2753,N_1451,N_401);
nor U2754 (N_2754,N_890,N_36);
nor U2755 (N_2755,N_937,N_51);
and U2756 (N_2756,N_1266,N_162);
and U2757 (N_2757,N_1234,N_167);
nor U2758 (N_2758,N_1091,N_680);
nand U2759 (N_2759,N_561,N_1565);
or U2760 (N_2760,N_1025,N_868);
or U2761 (N_2761,N_1419,N_808);
or U2762 (N_2762,N_241,N_1682);
nor U2763 (N_2763,N_546,N_1885);
nor U2764 (N_2764,N_1595,N_1398);
and U2765 (N_2765,N_1251,N_1867);
or U2766 (N_2766,N_1660,N_451);
and U2767 (N_2767,N_1183,N_555);
nor U2768 (N_2768,N_1292,N_1051);
nor U2769 (N_2769,N_1474,N_1921);
or U2770 (N_2770,N_1828,N_573);
and U2771 (N_2771,N_35,N_1720);
nor U2772 (N_2772,N_757,N_375);
nor U2773 (N_2773,N_1514,N_1102);
nand U2774 (N_2774,N_839,N_1192);
nand U2775 (N_2775,N_226,N_314);
nor U2776 (N_2776,N_735,N_1535);
or U2777 (N_2777,N_1737,N_627);
or U2778 (N_2778,N_1601,N_933);
nand U2779 (N_2779,N_552,N_263);
or U2780 (N_2780,N_96,N_1819);
nor U2781 (N_2781,N_659,N_911);
and U2782 (N_2782,N_211,N_1916);
and U2783 (N_2783,N_1465,N_180);
and U2784 (N_2784,N_649,N_779);
nor U2785 (N_2785,N_113,N_1559);
nor U2786 (N_2786,N_440,N_965);
nand U2787 (N_2787,N_1471,N_1563);
nand U2788 (N_2788,N_250,N_1173);
and U2789 (N_2789,N_293,N_98);
nor U2790 (N_2790,N_967,N_300);
or U2791 (N_2791,N_560,N_832);
nor U2792 (N_2792,N_811,N_1897);
and U2793 (N_2793,N_1507,N_1700);
or U2794 (N_2794,N_514,N_1279);
nor U2795 (N_2795,N_824,N_1738);
or U2796 (N_2796,N_351,N_1951);
nor U2797 (N_2797,N_1237,N_1801);
and U2798 (N_2798,N_1311,N_1076);
nor U2799 (N_2799,N_1740,N_641);
or U2800 (N_2800,N_297,N_1692);
or U2801 (N_2801,N_385,N_498);
nand U2802 (N_2802,N_1378,N_1275);
and U2803 (N_2803,N_638,N_1030);
nor U2804 (N_2804,N_1134,N_1020);
and U2805 (N_2805,N_538,N_22);
and U2806 (N_2806,N_1905,N_1194);
nand U2807 (N_2807,N_1230,N_745);
and U2808 (N_2808,N_1969,N_617);
nand U2809 (N_2809,N_1291,N_129);
nor U2810 (N_2810,N_329,N_1354);
nand U2811 (N_2811,N_115,N_416);
nand U2812 (N_2812,N_1120,N_1703);
and U2813 (N_2813,N_1203,N_1044);
and U2814 (N_2814,N_761,N_1866);
nor U2815 (N_2815,N_1845,N_642);
nor U2816 (N_2816,N_1282,N_468);
or U2817 (N_2817,N_1602,N_607);
nor U2818 (N_2818,N_1997,N_859);
nor U2819 (N_2819,N_882,N_1855);
nor U2820 (N_2820,N_1628,N_622);
or U2821 (N_2821,N_1972,N_1833);
nor U2822 (N_2822,N_1108,N_629);
nor U2823 (N_2823,N_415,N_827);
nor U2824 (N_2824,N_1016,N_1539);
and U2825 (N_2825,N_1582,N_328);
and U2826 (N_2826,N_1106,N_1804);
or U2827 (N_2827,N_306,N_866);
or U2828 (N_2828,N_99,N_1129);
and U2829 (N_2829,N_1295,N_770);
nor U2830 (N_2830,N_1484,N_6);
or U2831 (N_2831,N_1958,N_1902);
and U2832 (N_2832,N_1039,N_341);
nor U2833 (N_2833,N_1564,N_1482);
nor U2834 (N_2834,N_1543,N_430);
or U2835 (N_2835,N_943,N_563);
nand U2836 (N_2836,N_108,N_21);
nand U2837 (N_2837,N_1111,N_1019);
xnor U2838 (N_2838,N_1336,N_820);
and U2839 (N_2839,N_1923,N_1244);
and U2840 (N_2840,N_1774,N_1453);
nor U2841 (N_2841,N_684,N_858);
or U2842 (N_2842,N_1131,N_1613);
or U2843 (N_2843,N_1848,N_1028);
or U2844 (N_2844,N_914,N_33);
and U2845 (N_2845,N_465,N_955);
or U2846 (N_2846,N_655,N_1418);
nor U2847 (N_2847,N_1615,N_110);
nand U2848 (N_2848,N_1373,N_340);
and U2849 (N_2849,N_1318,N_1755);
nand U2850 (N_2850,N_447,N_274);
nor U2851 (N_2851,N_61,N_775);
nor U2852 (N_2852,N_1904,N_1259);
or U2853 (N_2853,N_1926,N_1544);
and U2854 (N_2854,N_280,N_3);
and U2855 (N_2855,N_926,N_83);
or U2856 (N_2856,N_921,N_1229);
or U2857 (N_2857,N_1888,N_1783);
nor U2858 (N_2858,N_1748,N_964);
nand U2859 (N_2859,N_1536,N_349);
and U2860 (N_2860,N_1123,N_1940);
nand U2861 (N_2861,N_205,N_1298);
nor U2862 (N_2862,N_994,N_1826);
nand U2863 (N_2863,N_400,N_1442);
or U2864 (N_2864,N_202,N_1844);
nor U2865 (N_2865,N_337,N_502);
nand U2866 (N_2866,N_1668,N_270);
nor U2867 (N_2867,N_1525,N_640);
nor U2868 (N_2868,N_1892,N_1331);
nand U2869 (N_2869,N_891,N_1889);
nor U2870 (N_2870,N_1361,N_1196);
nand U2871 (N_2871,N_38,N_257);
nor U2872 (N_2872,N_1384,N_1317);
nor U2873 (N_2873,N_1045,N_1235);
nand U2874 (N_2874,N_1215,N_688);
and U2875 (N_2875,N_1114,N_103);
or U2876 (N_2876,N_1494,N_941);
or U2877 (N_2877,N_325,N_285);
or U2878 (N_2878,N_197,N_184);
or U2879 (N_2879,N_1348,N_249);
nand U2880 (N_2880,N_496,N_599);
xnor U2881 (N_2881,N_951,N_970);
and U2882 (N_2882,N_605,N_1256);
nor U2883 (N_2883,N_952,N_1815);
and U2884 (N_2884,N_1817,N_1726);
nand U2885 (N_2885,N_505,N_147);
nor U2886 (N_2886,N_772,N_623);
nand U2887 (N_2887,N_277,N_1717);
xor U2888 (N_2888,N_903,N_639);
and U2889 (N_2889,N_765,N_1490);
and U2890 (N_2890,N_1467,N_24);
or U2891 (N_2891,N_1125,N_1956);
and U2892 (N_2892,N_1272,N_682);
or U2893 (N_2893,N_1664,N_1312);
or U2894 (N_2894,N_1642,N_922);
and U2895 (N_2895,N_963,N_1483);
nor U2896 (N_2896,N_1771,N_1752);
nor U2897 (N_2897,N_730,N_1631);
or U2898 (N_2898,N_1287,N_1413);
nand U2899 (N_2899,N_1263,N_1745);
or U2900 (N_2900,N_752,N_718);
and U2901 (N_2901,N_1906,N_1058);
and U2902 (N_2902,N_656,N_1814);
and U2903 (N_2903,N_1403,N_976);
nand U2904 (N_2904,N_1207,N_422);
nor U2905 (N_2905,N_722,N_126);
and U2906 (N_2906,N_1769,N_214);
or U2907 (N_2907,N_715,N_826);
nor U2908 (N_2908,N_1486,N_164);
nand U2909 (N_2909,N_246,N_1947);
and U2910 (N_2910,N_1629,N_1394);
nor U2911 (N_2911,N_183,N_540);
nand U2912 (N_2912,N_17,N_1082);
nor U2913 (N_2913,N_1712,N_1747);
and U2914 (N_2914,N_786,N_1653);
nor U2915 (N_2915,N_1961,N_1989);
or U2916 (N_2916,N_26,N_800);
nor U2917 (N_2917,N_1079,N_631);
nor U2918 (N_2918,N_1917,N_940);
or U2919 (N_2919,N_574,N_806);
or U2920 (N_2920,N_423,N_1440);
and U2921 (N_2921,N_542,N_335);
nor U2922 (N_2922,N_1794,N_912);
or U2923 (N_2923,N_1217,N_969);
or U2924 (N_2924,N_1115,N_1055);
or U2925 (N_2925,N_930,N_1014);
and U2926 (N_2926,N_813,N_326);
nand U2927 (N_2927,N_363,N_1977);
nor U2928 (N_2928,N_392,N_1782);
nor U2929 (N_2929,N_1583,N_161);
and U2930 (N_2930,N_1982,N_1059);
and U2931 (N_2931,N_261,N_130);
and U2932 (N_2932,N_762,N_1198);
and U2933 (N_2933,N_288,N_152);
nand U2934 (N_2934,N_158,N_443);
and U2935 (N_2935,N_1618,N_673);
or U2936 (N_2936,N_374,N_203);
nor U2937 (N_2937,N_1447,N_345);
or U2938 (N_2938,N_1903,N_1136);
and U2939 (N_2939,N_1383,N_299);
or U2940 (N_2940,N_906,N_1648);
and U2941 (N_2941,N_452,N_1220);
or U2942 (N_2942,N_493,N_407);
nand U2943 (N_2943,N_301,N_140);
nor U2944 (N_2944,N_1049,N_1919);
or U2945 (N_2945,N_693,N_395);
nand U2946 (N_2946,N_1389,N_166);
and U2947 (N_2947,N_1556,N_1232);
nor U2948 (N_2948,N_562,N_741);
and U2949 (N_2949,N_359,N_1386);
nand U2950 (N_2950,N_1119,N_380);
nor U2951 (N_2951,N_662,N_1364);
and U2952 (N_2952,N_1893,N_1193);
nor U2953 (N_2953,N_56,N_1935);
nand U2954 (N_2954,N_403,N_1330);
nand U2955 (N_2955,N_1991,N_1240);
or U2956 (N_2956,N_1541,N_1843);
or U2957 (N_2957,N_62,N_1832);
or U2958 (N_2958,N_1126,N_1104);
and U2959 (N_2959,N_949,N_1810);
nor U2960 (N_2960,N_160,N_1706);
nand U2961 (N_2961,N_1829,N_893);
or U2962 (N_2962,N_223,N_1366);
and U2963 (N_2963,N_1572,N_1135);
nor U2964 (N_2964,N_1334,N_163);
nand U2965 (N_2965,N_1939,N_1610);
nor U2966 (N_2966,N_1799,N_151);
or U2967 (N_2967,N_391,N_1589);
nor U2968 (N_2968,N_559,N_795);
and U2969 (N_2969,N_699,N_1870);
nor U2970 (N_2970,N_1073,N_1429);
and U2971 (N_2971,N_1265,N_1148);
nand U2972 (N_2972,N_1029,N_1626);
or U2973 (N_2973,N_1434,N_506);
nand U2974 (N_2974,N_1959,N_1061);
nand U2975 (N_2975,N_875,N_122);
nor U2976 (N_2976,N_700,N_1396);
or U2977 (N_2977,N_703,N_1861);
and U2978 (N_2978,N_581,N_1871);
nor U2979 (N_2979,N_315,N_387);
nand U2980 (N_2980,N_1449,N_738);
or U2981 (N_2981,N_1309,N_1497);
nor U2982 (N_2982,N_621,N_470);
nand U2983 (N_2983,N_1560,N_870);
nand U2984 (N_2984,N_1946,N_253);
nor U2985 (N_2985,N_1963,N_1147);
and U2986 (N_2986,N_1420,N_764);
or U2987 (N_2987,N_1852,N_350);
or U2988 (N_2988,N_1032,N_1328);
or U2989 (N_2989,N_1476,N_1454);
or U2990 (N_2990,N_1267,N_39);
and U2991 (N_2991,N_512,N_635);
nor U2992 (N_2992,N_1534,N_1322);
or U2993 (N_2993,N_1862,N_750);
and U2994 (N_2994,N_236,N_1286);
or U2995 (N_2995,N_1412,N_925);
or U2996 (N_2996,N_945,N_886);
or U2997 (N_2997,N_702,N_1034);
and U2998 (N_2998,N_333,N_1200);
or U2999 (N_2999,N_842,N_862);
nand U3000 (N_3000,N_224,N_54);
nand U3001 (N_3001,N_227,N_1083);
and U3002 (N_3002,N_857,N_183);
and U3003 (N_3003,N_733,N_1802);
nor U3004 (N_3004,N_545,N_1334);
nand U3005 (N_3005,N_41,N_1132);
nand U3006 (N_3006,N_139,N_898);
or U3007 (N_3007,N_458,N_1045);
nor U3008 (N_3008,N_1208,N_1088);
nor U3009 (N_3009,N_318,N_35);
and U3010 (N_3010,N_381,N_69);
nand U3011 (N_3011,N_316,N_1945);
nand U3012 (N_3012,N_349,N_961);
nor U3013 (N_3013,N_1985,N_359);
nor U3014 (N_3014,N_1978,N_212);
and U3015 (N_3015,N_1209,N_1819);
nand U3016 (N_3016,N_1706,N_1174);
or U3017 (N_3017,N_16,N_1505);
and U3018 (N_3018,N_1721,N_1792);
nand U3019 (N_3019,N_1372,N_793);
or U3020 (N_3020,N_1995,N_1765);
or U3021 (N_3021,N_1205,N_1225);
or U3022 (N_3022,N_1096,N_71);
or U3023 (N_3023,N_1072,N_859);
nor U3024 (N_3024,N_769,N_664);
nor U3025 (N_3025,N_1309,N_1583);
and U3026 (N_3026,N_661,N_894);
or U3027 (N_3027,N_1773,N_1919);
or U3028 (N_3028,N_1088,N_301);
or U3029 (N_3029,N_217,N_878);
and U3030 (N_3030,N_1179,N_506);
and U3031 (N_3031,N_1557,N_733);
nor U3032 (N_3032,N_326,N_1218);
and U3033 (N_3033,N_1705,N_395);
nor U3034 (N_3034,N_251,N_1109);
nand U3035 (N_3035,N_117,N_81);
nor U3036 (N_3036,N_1898,N_1210);
nor U3037 (N_3037,N_603,N_192);
nand U3038 (N_3038,N_847,N_1369);
nand U3039 (N_3039,N_1312,N_933);
or U3040 (N_3040,N_368,N_369);
and U3041 (N_3041,N_1639,N_286);
or U3042 (N_3042,N_342,N_351);
and U3043 (N_3043,N_1239,N_1933);
nand U3044 (N_3044,N_280,N_1475);
nand U3045 (N_3045,N_1242,N_1282);
nor U3046 (N_3046,N_1938,N_1203);
nor U3047 (N_3047,N_1103,N_1628);
xnor U3048 (N_3048,N_174,N_1742);
or U3049 (N_3049,N_1573,N_1341);
nor U3050 (N_3050,N_54,N_1161);
nand U3051 (N_3051,N_1599,N_550);
nand U3052 (N_3052,N_954,N_1573);
or U3053 (N_3053,N_597,N_1596);
or U3054 (N_3054,N_458,N_27);
and U3055 (N_3055,N_429,N_1700);
or U3056 (N_3056,N_1233,N_1596);
or U3057 (N_3057,N_1621,N_671);
nor U3058 (N_3058,N_1998,N_821);
nor U3059 (N_3059,N_669,N_68);
nand U3060 (N_3060,N_865,N_1786);
nand U3061 (N_3061,N_1273,N_1909);
and U3062 (N_3062,N_627,N_1484);
nand U3063 (N_3063,N_643,N_1512);
nand U3064 (N_3064,N_341,N_1716);
nor U3065 (N_3065,N_462,N_447);
and U3066 (N_3066,N_1005,N_925);
and U3067 (N_3067,N_459,N_265);
or U3068 (N_3068,N_117,N_1480);
nand U3069 (N_3069,N_39,N_104);
or U3070 (N_3070,N_1628,N_1731);
and U3071 (N_3071,N_1720,N_241);
nand U3072 (N_3072,N_490,N_1592);
nand U3073 (N_3073,N_265,N_1528);
nand U3074 (N_3074,N_1182,N_1857);
or U3075 (N_3075,N_1863,N_1502);
nand U3076 (N_3076,N_550,N_1883);
nand U3077 (N_3077,N_105,N_1810);
nand U3078 (N_3078,N_1481,N_989);
or U3079 (N_3079,N_1135,N_53);
nand U3080 (N_3080,N_1052,N_1712);
nor U3081 (N_3081,N_121,N_981);
nor U3082 (N_3082,N_27,N_946);
nand U3083 (N_3083,N_1978,N_1143);
nand U3084 (N_3084,N_1500,N_1000);
or U3085 (N_3085,N_974,N_502);
nand U3086 (N_3086,N_300,N_1521);
nand U3087 (N_3087,N_181,N_46);
or U3088 (N_3088,N_1275,N_14);
nor U3089 (N_3089,N_474,N_386);
nor U3090 (N_3090,N_207,N_1898);
and U3091 (N_3091,N_1087,N_726);
nor U3092 (N_3092,N_1300,N_850);
or U3093 (N_3093,N_1332,N_1561);
and U3094 (N_3094,N_641,N_375);
nor U3095 (N_3095,N_1441,N_1869);
nor U3096 (N_3096,N_253,N_1715);
or U3097 (N_3097,N_264,N_1276);
or U3098 (N_3098,N_219,N_1678);
nor U3099 (N_3099,N_1756,N_198);
or U3100 (N_3100,N_1240,N_274);
and U3101 (N_3101,N_1013,N_1631);
nor U3102 (N_3102,N_1483,N_470);
or U3103 (N_3103,N_420,N_458);
or U3104 (N_3104,N_140,N_510);
or U3105 (N_3105,N_1215,N_1871);
nor U3106 (N_3106,N_1528,N_24);
and U3107 (N_3107,N_1288,N_1117);
and U3108 (N_3108,N_1621,N_1078);
or U3109 (N_3109,N_555,N_1312);
and U3110 (N_3110,N_1428,N_603);
and U3111 (N_3111,N_1816,N_982);
and U3112 (N_3112,N_796,N_660);
nor U3113 (N_3113,N_239,N_701);
nand U3114 (N_3114,N_486,N_1174);
nand U3115 (N_3115,N_784,N_1301);
or U3116 (N_3116,N_731,N_1884);
nand U3117 (N_3117,N_926,N_1334);
and U3118 (N_3118,N_1010,N_1148);
nor U3119 (N_3119,N_38,N_1111);
nor U3120 (N_3120,N_39,N_1957);
nand U3121 (N_3121,N_1558,N_987);
and U3122 (N_3122,N_26,N_385);
xor U3123 (N_3123,N_352,N_1794);
nand U3124 (N_3124,N_1287,N_29);
or U3125 (N_3125,N_417,N_1197);
or U3126 (N_3126,N_346,N_897);
xnor U3127 (N_3127,N_181,N_1842);
nor U3128 (N_3128,N_1422,N_831);
or U3129 (N_3129,N_1440,N_1588);
nor U3130 (N_3130,N_1230,N_1459);
xor U3131 (N_3131,N_1516,N_1949);
or U3132 (N_3132,N_1738,N_1802);
and U3133 (N_3133,N_1754,N_932);
nand U3134 (N_3134,N_39,N_818);
and U3135 (N_3135,N_1286,N_1786);
nor U3136 (N_3136,N_1864,N_772);
xor U3137 (N_3137,N_1596,N_1692);
or U3138 (N_3138,N_575,N_1919);
and U3139 (N_3139,N_1074,N_458);
or U3140 (N_3140,N_1307,N_1016);
and U3141 (N_3141,N_1178,N_776);
nand U3142 (N_3142,N_1235,N_23);
nor U3143 (N_3143,N_418,N_1044);
nor U3144 (N_3144,N_1708,N_736);
or U3145 (N_3145,N_1617,N_1317);
and U3146 (N_3146,N_1153,N_1166);
and U3147 (N_3147,N_1641,N_1167);
nor U3148 (N_3148,N_1835,N_1778);
or U3149 (N_3149,N_235,N_792);
nor U3150 (N_3150,N_417,N_794);
or U3151 (N_3151,N_1112,N_570);
nand U3152 (N_3152,N_1470,N_586);
nand U3153 (N_3153,N_1513,N_1311);
nor U3154 (N_3154,N_1180,N_1718);
nor U3155 (N_3155,N_221,N_198);
nor U3156 (N_3156,N_1089,N_1802);
and U3157 (N_3157,N_768,N_1118);
nor U3158 (N_3158,N_1472,N_960);
nor U3159 (N_3159,N_495,N_195);
nor U3160 (N_3160,N_1852,N_280);
and U3161 (N_3161,N_1967,N_748);
nand U3162 (N_3162,N_1754,N_1071);
or U3163 (N_3163,N_284,N_1925);
nand U3164 (N_3164,N_310,N_1429);
and U3165 (N_3165,N_1921,N_1129);
nand U3166 (N_3166,N_668,N_1258);
and U3167 (N_3167,N_1286,N_1882);
and U3168 (N_3168,N_1577,N_568);
nand U3169 (N_3169,N_276,N_390);
and U3170 (N_3170,N_1920,N_1555);
or U3171 (N_3171,N_631,N_276);
or U3172 (N_3172,N_1257,N_535);
and U3173 (N_3173,N_893,N_930);
nor U3174 (N_3174,N_1977,N_1181);
xnor U3175 (N_3175,N_1747,N_445);
or U3176 (N_3176,N_321,N_664);
or U3177 (N_3177,N_1652,N_113);
nand U3178 (N_3178,N_1280,N_696);
nand U3179 (N_3179,N_1845,N_997);
nand U3180 (N_3180,N_1907,N_1984);
and U3181 (N_3181,N_936,N_1563);
nor U3182 (N_3182,N_1138,N_1218);
nor U3183 (N_3183,N_663,N_1273);
or U3184 (N_3184,N_1681,N_1146);
or U3185 (N_3185,N_150,N_1651);
and U3186 (N_3186,N_1993,N_1476);
nor U3187 (N_3187,N_1338,N_330);
or U3188 (N_3188,N_778,N_1163);
or U3189 (N_3189,N_1061,N_115);
nor U3190 (N_3190,N_95,N_1158);
and U3191 (N_3191,N_752,N_1276);
and U3192 (N_3192,N_1805,N_636);
nand U3193 (N_3193,N_509,N_524);
nand U3194 (N_3194,N_801,N_770);
nor U3195 (N_3195,N_1165,N_590);
and U3196 (N_3196,N_208,N_1095);
and U3197 (N_3197,N_849,N_1671);
nor U3198 (N_3198,N_424,N_1446);
nand U3199 (N_3199,N_583,N_1227);
nor U3200 (N_3200,N_89,N_1909);
or U3201 (N_3201,N_274,N_1587);
or U3202 (N_3202,N_812,N_1265);
or U3203 (N_3203,N_997,N_1267);
nand U3204 (N_3204,N_1605,N_1789);
or U3205 (N_3205,N_1590,N_552);
and U3206 (N_3206,N_361,N_848);
and U3207 (N_3207,N_1419,N_945);
nand U3208 (N_3208,N_1093,N_1562);
nand U3209 (N_3209,N_1179,N_1476);
nand U3210 (N_3210,N_1994,N_131);
nand U3211 (N_3211,N_258,N_447);
nand U3212 (N_3212,N_535,N_1557);
or U3213 (N_3213,N_1104,N_1999);
and U3214 (N_3214,N_172,N_109);
nand U3215 (N_3215,N_1449,N_1612);
and U3216 (N_3216,N_307,N_1305);
nor U3217 (N_3217,N_1212,N_320);
or U3218 (N_3218,N_55,N_178);
or U3219 (N_3219,N_1191,N_332);
nor U3220 (N_3220,N_293,N_82);
nor U3221 (N_3221,N_1816,N_1056);
nor U3222 (N_3222,N_1063,N_1611);
nor U3223 (N_3223,N_1044,N_755);
nor U3224 (N_3224,N_724,N_1118);
and U3225 (N_3225,N_666,N_1865);
nor U3226 (N_3226,N_1920,N_1214);
or U3227 (N_3227,N_186,N_660);
or U3228 (N_3228,N_250,N_1741);
nor U3229 (N_3229,N_1342,N_296);
and U3230 (N_3230,N_517,N_961);
nor U3231 (N_3231,N_329,N_1686);
and U3232 (N_3232,N_1885,N_1001);
nand U3233 (N_3233,N_337,N_992);
nor U3234 (N_3234,N_1661,N_1530);
and U3235 (N_3235,N_1871,N_595);
and U3236 (N_3236,N_164,N_652);
or U3237 (N_3237,N_1213,N_342);
nor U3238 (N_3238,N_421,N_1280);
nand U3239 (N_3239,N_1566,N_1747);
or U3240 (N_3240,N_1677,N_1482);
and U3241 (N_3241,N_1564,N_1715);
and U3242 (N_3242,N_461,N_91);
or U3243 (N_3243,N_1838,N_1889);
and U3244 (N_3244,N_1998,N_265);
and U3245 (N_3245,N_1750,N_1129);
or U3246 (N_3246,N_1866,N_632);
nand U3247 (N_3247,N_43,N_1415);
nor U3248 (N_3248,N_1229,N_1859);
nor U3249 (N_3249,N_1776,N_1021);
or U3250 (N_3250,N_1650,N_440);
or U3251 (N_3251,N_1388,N_1395);
nand U3252 (N_3252,N_156,N_1827);
and U3253 (N_3253,N_133,N_1127);
nand U3254 (N_3254,N_974,N_920);
and U3255 (N_3255,N_250,N_1169);
and U3256 (N_3256,N_1156,N_848);
nand U3257 (N_3257,N_823,N_1853);
or U3258 (N_3258,N_1730,N_747);
or U3259 (N_3259,N_1357,N_1505);
nand U3260 (N_3260,N_6,N_1571);
and U3261 (N_3261,N_337,N_660);
or U3262 (N_3262,N_1988,N_1537);
or U3263 (N_3263,N_1010,N_842);
or U3264 (N_3264,N_817,N_1859);
or U3265 (N_3265,N_1888,N_229);
and U3266 (N_3266,N_524,N_1212);
and U3267 (N_3267,N_959,N_358);
and U3268 (N_3268,N_20,N_38);
or U3269 (N_3269,N_852,N_267);
and U3270 (N_3270,N_1601,N_325);
and U3271 (N_3271,N_547,N_544);
nand U3272 (N_3272,N_1145,N_1758);
or U3273 (N_3273,N_93,N_847);
and U3274 (N_3274,N_378,N_5);
nor U3275 (N_3275,N_1586,N_1985);
and U3276 (N_3276,N_1411,N_1288);
nor U3277 (N_3277,N_1403,N_958);
or U3278 (N_3278,N_1976,N_645);
xnor U3279 (N_3279,N_846,N_894);
or U3280 (N_3280,N_1950,N_1577);
and U3281 (N_3281,N_251,N_436);
nand U3282 (N_3282,N_881,N_1445);
or U3283 (N_3283,N_170,N_173);
and U3284 (N_3284,N_1158,N_986);
nor U3285 (N_3285,N_108,N_276);
or U3286 (N_3286,N_1066,N_1250);
and U3287 (N_3287,N_725,N_1152);
nand U3288 (N_3288,N_655,N_432);
nor U3289 (N_3289,N_567,N_846);
nand U3290 (N_3290,N_206,N_1215);
or U3291 (N_3291,N_723,N_340);
or U3292 (N_3292,N_1912,N_814);
and U3293 (N_3293,N_1030,N_485);
nor U3294 (N_3294,N_1854,N_547);
nand U3295 (N_3295,N_1158,N_1843);
nor U3296 (N_3296,N_181,N_1943);
nor U3297 (N_3297,N_788,N_1307);
nand U3298 (N_3298,N_1825,N_1631);
and U3299 (N_3299,N_173,N_867);
and U3300 (N_3300,N_655,N_1699);
and U3301 (N_3301,N_722,N_797);
nor U3302 (N_3302,N_1003,N_544);
nor U3303 (N_3303,N_1461,N_137);
and U3304 (N_3304,N_210,N_1702);
nand U3305 (N_3305,N_1086,N_506);
nor U3306 (N_3306,N_1785,N_663);
and U3307 (N_3307,N_1812,N_1166);
nand U3308 (N_3308,N_1548,N_411);
nor U3309 (N_3309,N_281,N_263);
nand U3310 (N_3310,N_1181,N_1919);
or U3311 (N_3311,N_1904,N_970);
nand U3312 (N_3312,N_453,N_203);
nor U3313 (N_3313,N_1569,N_57);
nand U3314 (N_3314,N_1184,N_539);
or U3315 (N_3315,N_1479,N_903);
nor U3316 (N_3316,N_561,N_1464);
nor U3317 (N_3317,N_1515,N_1394);
nor U3318 (N_3318,N_1671,N_911);
nor U3319 (N_3319,N_832,N_1712);
or U3320 (N_3320,N_1036,N_164);
and U3321 (N_3321,N_404,N_405);
or U3322 (N_3322,N_989,N_441);
and U3323 (N_3323,N_467,N_302);
and U3324 (N_3324,N_239,N_1950);
and U3325 (N_3325,N_1495,N_736);
nor U3326 (N_3326,N_1992,N_1561);
nor U3327 (N_3327,N_1848,N_1192);
nand U3328 (N_3328,N_671,N_1524);
nand U3329 (N_3329,N_1840,N_1825);
nor U3330 (N_3330,N_1110,N_1951);
nor U3331 (N_3331,N_1876,N_791);
nand U3332 (N_3332,N_649,N_1081);
or U3333 (N_3333,N_827,N_1311);
nand U3334 (N_3334,N_855,N_645);
nand U3335 (N_3335,N_1465,N_453);
nand U3336 (N_3336,N_792,N_1393);
nand U3337 (N_3337,N_1849,N_1330);
nand U3338 (N_3338,N_1870,N_1260);
nor U3339 (N_3339,N_1543,N_1019);
nand U3340 (N_3340,N_817,N_1887);
xnor U3341 (N_3341,N_1670,N_336);
or U3342 (N_3342,N_1718,N_422);
or U3343 (N_3343,N_368,N_1448);
and U3344 (N_3344,N_1805,N_258);
nand U3345 (N_3345,N_1559,N_1908);
or U3346 (N_3346,N_1139,N_51);
or U3347 (N_3347,N_615,N_185);
or U3348 (N_3348,N_833,N_964);
nor U3349 (N_3349,N_337,N_745);
or U3350 (N_3350,N_321,N_9);
and U3351 (N_3351,N_112,N_525);
nand U3352 (N_3352,N_1812,N_432);
or U3353 (N_3353,N_1459,N_312);
and U3354 (N_3354,N_1734,N_1237);
nand U3355 (N_3355,N_1323,N_462);
nand U3356 (N_3356,N_419,N_501);
or U3357 (N_3357,N_1048,N_452);
or U3358 (N_3358,N_116,N_463);
nor U3359 (N_3359,N_445,N_284);
or U3360 (N_3360,N_138,N_1097);
or U3361 (N_3361,N_534,N_1860);
nor U3362 (N_3362,N_679,N_1870);
or U3363 (N_3363,N_1256,N_590);
and U3364 (N_3364,N_1409,N_1157);
nand U3365 (N_3365,N_1523,N_334);
or U3366 (N_3366,N_1198,N_241);
nand U3367 (N_3367,N_678,N_1146);
or U3368 (N_3368,N_83,N_1079);
nor U3369 (N_3369,N_264,N_1521);
nand U3370 (N_3370,N_153,N_85);
and U3371 (N_3371,N_484,N_960);
nand U3372 (N_3372,N_720,N_1283);
or U3373 (N_3373,N_1815,N_1093);
nand U3374 (N_3374,N_679,N_51);
or U3375 (N_3375,N_1495,N_1015);
and U3376 (N_3376,N_1051,N_1487);
nor U3377 (N_3377,N_1522,N_1437);
nand U3378 (N_3378,N_1762,N_1866);
or U3379 (N_3379,N_1325,N_1695);
nor U3380 (N_3380,N_512,N_1724);
nand U3381 (N_3381,N_1504,N_1644);
and U3382 (N_3382,N_887,N_1112);
or U3383 (N_3383,N_886,N_1294);
nor U3384 (N_3384,N_1120,N_890);
and U3385 (N_3385,N_1346,N_1454);
nor U3386 (N_3386,N_392,N_427);
or U3387 (N_3387,N_1481,N_958);
nor U3388 (N_3388,N_298,N_112);
nand U3389 (N_3389,N_653,N_729);
and U3390 (N_3390,N_910,N_943);
and U3391 (N_3391,N_1721,N_1162);
nor U3392 (N_3392,N_146,N_63);
or U3393 (N_3393,N_1044,N_1042);
nand U3394 (N_3394,N_1680,N_1166);
or U3395 (N_3395,N_1381,N_1270);
nor U3396 (N_3396,N_414,N_182);
nor U3397 (N_3397,N_1394,N_1886);
or U3398 (N_3398,N_418,N_1771);
nor U3399 (N_3399,N_959,N_390);
or U3400 (N_3400,N_1735,N_596);
and U3401 (N_3401,N_554,N_1927);
and U3402 (N_3402,N_149,N_550);
and U3403 (N_3403,N_155,N_1887);
nand U3404 (N_3404,N_1410,N_1267);
or U3405 (N_3405,N_727,N_1538);
nor U3406 (N_3406,N_331,N_1695);
and U3407 (N_3407,N_811,N_334);
or U3408 (N_3408,N_367,N_931);
nand U3409 (N_3409,N_1572,N_27);
nor U3410 (N_3410,N_192,N_581);
nor U3411 (N_3411,N_612,N_1705);
and U3412 (N_3412,N_1125,N_741);
nand U3413 (N_3413,N_1048,N_1835);
and U3414 (N_3414,N_1979,N_1608);
or U3415 (N_3415,N_604,N_949);
nand U3416 (N_3416,N_1784,N_626);
or U3417 (N_3417,N_214,N_1926);
nor U3418 (N_3418,N_871,N_1723);
nand U3419 (N_3419,N_1765,N_117);
nor U3420 (N_3420,N_980,N_889);
nand U3421 (N_3421,N_614,N_33);
and U3422 (N_3422,N_747,N_1957);
nand U3423 (N_3423,N_544,N_273);
nand U3424 (N_3424,N_1141,N_1110);
and U3425 (N_3425,N_162,N_544);
or U3426 (N_3426,N_99,N_1775);
or U3427 (N_3427,N_176,N_1185);
xnor U3428 (N_3428,N_1480,N_1538);
or U3429 (N_3429,N_498,N_1662);
nand U3430 (N_3430,N_678,N_1568);
nor U3431 (N_3431,N_1915,N_1541);
and U3432 (N_3432,N_1415,N_247);
and U3433 (N_3433,N_738,N_1982);
nand U3434 (N_3434,N_514,N_336);
and U3435 (N_3435,N_191,N_313);
and U3436 (N_3436,N_403,N_1132);
or U3437 (N_3437,N_311,N_1714);
nand U3438 (N_3438,N_1923,N_952);
nor U3439 (N_3439,N_1866,N_1514);
or U3440 (N_3440,N_37,N_144);
or U3441 (N_3441,N_1165,N_660);
nand U3442 (N_3442,N_1089,N_218);
nand U3443 (N_3443,N_618,N_1845);
nor U3444 (N_3444,N_1411,N_272);
nand U3445 (N_3445,N_190,N_1225);
and U3446 (N_3446,N_820,N_1534);
or U3447 (N_3447,N_528,N_403);
nand U3448 (N_3448,N_1924,N_1054);
and U3449 (N_3449,N_1874,N_1579);
nand U3450 (N_3450,N_1124,N_1562);
nor U3451 (N_3451,N_1485,N_225);
or U3452 (N_3452,N_1365,N_865);
and U3453 (N_3453,N_616,N_1989);
or U3454 (N_3454,N_1832,N_904);
nor U3455 (N_3455,N_1199,N_116);
nor U3456 (N_3456,N_1970,N_1123);
nand U3457 (N_3457,N_1199,N_902);
or U3458 (N_3458,N_265,N_1669);
nor U3459 (N_3459,N_1266,N_1883);
and U3460 (N_3460,N_1070,N_1008);
or U3461 (N_3461,N_1536,N_1077);
nand U3462 (N_3462,N_407,N_210);
or U3463 (N_3463,N_993,N_61);
nor U3464 (N_3464,N_956,N_1702);
and U3465 (N_3465,N_536,N_29);
nor U3466 (N_3466,N_1729,N_1686);
and U3467 (N_3467,N_656,N_728);
or U3468 (N_3468,N_1444,N_1759);
nand U3469 (N_3469,N_600,N_1298);
and U3470 (N_3470,N_118,N_926);
nor U3471 (N_3471,N_633,N_1873);
or U3472 (N_3472,N_1652,N_136);
nand U3473 (N_3473,N_1181,N_1561);
or U3474 (N_3474,N_1993,N_1905);
nor U3475 (N_3475,N_158,N_1028);
nor U3476 (N_3476,N_1123,N_98);
and U3477 (N_3477,N_236,N_305);
or U3478 (N_3478,N_564,N_1202);
or U3479 (N_3479,N_314,N_555);
or U3480 (N_3480,N_578,N_1996);
and U3481 (N_3481,N_39,N_1597);
nand U3482 (N_3482,N_430,N_1869);
and U3483 (N_3483,N_406,N_1606);
nor U3484 (N_3484,N_1614,N_867);
nor U3485 (N_3485,N_71,N_1361);
nand U3486 (N_3486,N_1245,N_1922);
nand U3487 (N_3487,N_277,N_385);
nand U3488 (N_3488,N_1243,N_1091);
nand U3489 (N_3489,N_382,N_1691);
or U3490 (N_3490,N_1171,N_756);
or U3491 (N_3491,N_709,N_642);
nor U3492 (N_3492,N_169,N_964);
nand U3493 (N_3493,N_302,N_734);
or U3494 (N_3494,N_1905,N_1724);
nor U3495 (N_3495,N_919,N_251);
or U3496 (N_3496,N_1322,N_313);
nor U3497 (N_3497,N_1157,N_662);
and U3498 (N_3498,N_112,N_1126);
and U3499 (N_3499,N_1084,N_461);
and U3500 (N_3500,N_565,N_759);
nor U3501 (N_3501,N_553,N_146);
and U3502 (N_3502,N_1112,N_237);
xor U3503 (N_3503,N_1370,N_561);
and U3504 (N_3504,N_547,N_984);
and U3505 (N_3505,N_816,N_1898);
nor U3506 (N_3506,N_529,N_739);
or U3507 (N_3507,N_1455,N_397);
and U3508 (N_3508,N_954,N_1644);
nand U3509 (N_3509,N_614,N_310);
nor U3510 (N_3510,N_1034,N_364);
or U3511 (N_3511,N_435,N_5);
nor U3512 (N_3512,N_393,N_1726);
nor U3513 (N_3513,N_179,N_840);
and U3514 (N_3514,N_1469,N_520);
or U3515 (N_3515,N_1819,N_312);
nand U3516 (N_3516,N_1216,N_527);
and U3517 (N_3517,N_380,N_1890);
or U3518 (N_3518,N_464,N_328);
or U3519 (N_3519,N_445,N_113);
or U3520 (N_3520,N_264,N_1565);
or U3521 (N_3521,N_1665,N_1499);
nand U3522 (N_3522,N_484,N_208);
and U3523 (N_3523,N_1306,N_1688);
nor U3524 (N_3524,N_785,N_1898);
nor U3525 (N_3525,N_419,N_932);
or U3526 (N_3526,N_1746,N_1349);
or U3527 (N_3527,N_387,N_779);
nand U3528 (N_3528,N_1338,N_662);
or U3529 (N_3529,N_1079,N_1468);
and U3530 (N_3530,N_612,N_292);
or U3531 (N_3531,N_186,N_138);
nor U3532 (N_3532,N_1556,N_767);
nor U3533 (N_3533,N_1773,N_1385);
xor U3534 (N_3534,N_322,N_803);
or U3535 (N_3535,N_1930,N_911);
nand U3536 (N_3536,N_1110,N_358);
nand U3537 (N_3537,N_493,N_247);
or U3538 (N_3538,N_105,N_12);
nor U3539 (N_3539,N_1976,N_530);
nand U3540 (N_3540,N_1523,N_623);
and U3541 (N_3541,N_787,N_488);
nor U3542 (N_3542,N_1260,N_1991);
or U3543 (N_3543,N_465,N_1381);
nor U3544 (N_3544,N_1901,N_42);
nand U3545 (N_3545,N_1427,N_1074);
and U3546 (N_3546,N_554,N_321);
and U3547 (N_3547,N_1812,N_420);
or U3548 (N_3548,N_578,N_963);
or U3549 (N_3549,N_970,N_1591);
nand U3550 (N_3550,N_1727,N_699);
nor U3551 (N_3551,N_685,N_937);
or U3552 (N_3552,N_1991,N_1440);
nand U3553 (N_3553,N_1113,N_1746);
nor U3554 (N_3554,N_1864,N_722);
and U3555 (N_3555,N_1901,N_118);
or U3556 (N_3556,N_1186,N_551);
and U3557 (N_3557,N_1482,N_1633);
or U3558 (N_3558,N_264,N_1266);
and U3559 (N_3559,N_491,N_1365);
or U3560 (N_3560,N_1921,N_1113);
nand U3561 (N_3561,N_826,N_0);
nand U3562 (N_3562,N_1380,N_1502);
nor U3563 (N_3563,N_1321,N_1481);
and U3564 (N_3564,N_632,N_1307);
nor U3565 (N_3565,N_584,N_78);
or U3566 (N_3566,N_1098,N_865);
nor U3567 (N_3567,N_378,N_1056);
or U3568 (N_3568,N_1999,N_1719);
nand U3569 (N_3569,N_1520,N_1237);
and U3570 (N_3570,N_1125,N_1900);
or U3571 (N_3571,N_813,N_1527);
nor U3572 (N_3572,N_1841,N_867);
and U3573 (N_3573,N_954,N_25);
or U3574 (N_3574,N_1623,N_1503);
nand U3575 (N_3575,N_114,N_1160);
or U3576 (N_3576,N_1386,N_12);
or U3577 (N_3577,N_1417,N_405);
nand U3578 (N_3578,N_76,N_1032);
nor U3579 (N_3579,N_33,N_1334);
xor U3580 (N_3580,N_296,N_407);
or U3581 (N_3581,N_1044,N_185);
nand U3582 (N_3582,N_1193,N_608);
and U3583 (N_3583,N_1533,N_72);
nand U3584 (N_3584,N_1872,N_897);
nor U3585 (N_3585,N_1580,N_1803);
nand U3586 (N_3586,N_1800,N_955);
or U3587 (N_3587,N_1362,N_649);
and U3588 (N_3588,N_45,N_321);
and U3589 (N_3589,N_724,N_272);
nor U3590 (N_3590,N_1034,N_1338);
and U3591 (N_3591,N_556,N_1669);
and U3592 (N_3592,N_995,N_176);
nor U3593 (N_3593,N_321,N_1974);
nor U3594 (N_3594,N_229,N_1325);
nor U3595 (N_3595,N_1598,N_1275);
and U3596 (N_3596,N_1270,N_335);
nor U3597 (N_3597,N_1753,N_1238);
xnor U3598 (N_3598,N_1304,N_72);
nand U3599 (N_3599,N_1301,N_203);
nor U3600 (N_3600,N_407,N_1899);
nand U3601 (N_3601,N_267,N_1088);
and U3602 (N_3602,N_1347,N_929);
nor U3603 (N_3603,N_1927,N_207);
or U3604 (N_3604,N_992,N_733);
nor U3605 (N_3605,N_1284,N_82);
and U3606 (N_3606,N_762,N_1189);
nor U3607 (N_3607,N_164,N_1661);
nor U3608 (N_3608,N_260,N_1738);
or U3609 (N_3609,N_30,N_1624);
nor U3610 (N_3610,N_434,N_1238);
nand U3611 (N_3611,N_1067,N_1149);
or U3612 (N_3612,N_579,N_1892);
nand U3613 (N_3613,N_1489,N_1357);
and U3614 (N_3614,N_559,N_1087);
or U3615 (N_3615,N_1482,N_1529);
and U3616 (N_3616,N_1291,N_550);
nor U3617 (N_3617,N_594,N_1144);
nor U3618 (N_3618,N_673,N_823);
nand U3619 (N_3619,N_25,N_1567);
nand U3620 (N_3620,N_1123,N_1944);
or U3621 (N_3621,N_343,N_1718);
and U3622 (N_3622,N_1,N_611);
and U3623 (N_3623,N_602,N_1477);
nor U3624 (N_3624,N_1926,N_754);
and U3625 (N_3625,N_1549,N_294);
nand U3626 (N_3626,N_1457,N_186);
nor U3627 (N_3627,N_1893,N_310);
nand U3628 (N_3628,N_1231,N_147);
and U3629 (N_3629,N_1836,N_1736);
and U3630 (N_3630,N_1672,N_1316);
and U3631 (N_3631,N_1287,N_1439);
nor U3632 (N_3632,N_439,N_940);
and U3633 (N_3633,N_51,N_374);
or U3634 (N_3634,N_160,N_826);
or U3635 (N_3635,N_1126,N_526);
nand U3636 (N_3636,N_845,N_1784);
nor U3637 (N_3637,N_1871,N_1764);
and U3638 (N_3638,N_104,N_732);
or U3639 (N_3639,N_897,N_1744);
nand U3640 (N_3640,N_103,N_1743);
nand U3641 (N_3641,N_907,N_1003);
nand U3642 (N_3642,N_1189,N_1379);
nand U3643 (N_3643,N_1161,N_609);
and U3644 (N_3644,N_1121,N_89);
and U3645 (N_3645,N_318,N_752);
or U3646 (N_3646,N_600,N_1280);
xnor U3647 (N_3647,N_1359,N_1325);
nor U3648 (N_3648,N_521,N_1796);
or U3649 (N_3649,N_158,N_84);
nand U3650 (N_3650,N_256,N_1096);
or U3651 (N_3651,N_711,N_999);
nor U3652 (N_3652,N_1774,N_828);
and U3653 (N_3653,N_209,N_512);
nand U3654 (N_3654,N_1889,N_978);
and U3655 (N_3655,N_360,N_271);
nor U3656 (N_3656,N_695,N_768);
or U3657 (N_3657,N_1786,N_1965);
xor U3658 (N_3658,N_1402,N_109);
nor U3659 (N_3659,N_420,N_953);
and U3660 (N_3660,N_1708,N_1295);
nand U3661 (N_3661,N_1157,N_1914);
nor U3662 (N_3662,N_1974,N_574);
nand U3663 (N_3663,N_416,N_174);
nand U3664 (N_3664,N_1561,N_677);
nand U3665 (N_3665,N_1339,N_1840);
and U3666 (N_3666,N_1315,N_115);
nand U3667 (N_3667,N_985,N_1306);
nand U3668 (N_3668,N_925,N_990);
nor U3669 (N_3669,N_924,N_105);
nor U3670 (N_3670,N_1459,N_234);
and U3671 (N_3671,N_790,N_531);
or U3672 (N_3672,N_417,N_564);
or U3673 (N_3673,N_1211,N_570);
nor U3674 (N_3674,N_1666,N_501);
nor U3675 (N_3675,N_540,N_1004);
nand U3676 (N_3676,N_1110,N_896);
and U3677 (N_3677,N_865,N_1052);
nand U3678 (N_3678,N_1470,N_959);
and U3679 (N_3679,N_178,N_362);
and U3680 (N_3680,N_71,N_468);
nand U3681 (N_3681,N_1034,N_1193);
xnor U3682 (N_3682,N_571,N_435);
nand U3683 (N_3683,N_1068,N_844);
nand U3684 (N_3684,N_1957,N_1808);
or U3685 (N_3685,N_273,N_1941);
nand U3686 (N_3686,N_405,N_345);
nor U3687 (N_3687,N_195,N_460);
and U3688 (N_3688,N_1223,N_659);
nor U3689 (N_3689,N_1197,N_390);
nand U3690 (N_3690,N_158,N_1218);
or U3691 (N_3691,N_1256,N_427);
nand U3692 (N_3692,N_1914,N_821);
nand U3693 (N_3693,N_1907,N_932);
and U3694 (N_3694,N_1543,N_1652);
nand U3695 (N_3695,N_955,N_985);
nand U3696 (N_3696,N_93,N_943);
nor U3697 (N_3697,N_1145,N_1507);
xor U3698 (N_3698,N_1351,N_902);
nor U3699 (N_3699,N_83,N_225);
or U3700 (N_3700,N_931,N_1737);
nand U3701 (N_3701,N_1443,N_1879);
nor U3702 (N_3702,N_406,N_1503);
or U3703 (N_3703,N_1282,N_378);
or U3704 (N_3704,N_1773,N_250);
nand U3705 (N_3705,N_974,N_1893);
or U3706 (N_3706,N_883,N_251);
and U3707 (N_3707,N_694,N_1310);
nor U3708 (N_3708,N_23,N_601);
or U3709 (N_3709,N_1053,N_482);
or U3710 (N_3710,N_10,N_1270);
nand U3711 (N_3711,N_1922,N_226);
nor U3712 (N_3712,N_555,N_838);
nand U3713 (N_3713,N_878,N_380);
nor U3714 (N_3714,N_1935,N_1096);
and U3715 (N_3715,N_380,N_383);
or U3716 (N_3716,N_1123,N_1543);
nand U3717 (N_3717,N_2,N_1508);
nand U3718 (N_3718,N_1075,N_20);
and U3719 (N_3719,N_619,N_410);
nand U3720 (N_3720,N_1228,N_117);
nand U3721 (N_3721,N_1270,N_430);
nand U3722 (N_3722,N_1916,N_1940);
nand U3723 (N_3723,N_1265,N_594);
or U3724 (N_3724,N_979,N_723);
or U3725 (N_3725,N_1020,N_1936);
or U3726 (N_3726,N_504,N_238);
or U3727 (N_3727,N_1389,N_693);
and U3728 (N_3728,N_424,N_67);
or U3729 (N_3729,N_456,N_1449);
nor U3730 (N_3730,N_1466,N_1696);
nor U3731 (N_3731,N_1966,N_1416);
and U3732 (N_3732,N_1971,N_695);
and U3733 (N_3733,N_853,N_1544);
and U3734 (N_3734,N_1743,N_1272);
or U3735 (N_3735,N_1372,N_1865);
or U3736 (N_3736,N_59,N_522);
nand U3737 (N_3737,N_473,N_1400);
nor U3738 (N_3738,N_396,N_643);
and U3739 (N_3739,N_1117,N_508);
and U3740 (N_3740,N_455,N_754);
nor U3741 (N_3741,N_1284,N_457);
xnor U3742 (N_3742,N_1788,N_860);
or U3743 (N_3743,N_92,N_1057);
nand U3744 (N_3744,N_201,N_1535);
and U3745 (N_3745,N_492,N_847);
and U3746 (N_3746,N_1758,N_966);
nand U3747 (N_3747,N_541,N_1757);
nor U3748 (N_3748,N_67,N_324);
or U3749 (N_3749,N_1567,N_1394);
or U3750 (N_3750,N_1395,N_1966);
and U3751 (N_3751,N_1856,N_1799);
and U3752 (N_3752,N_1037,N_1185);
nor U3753 (N_3753,N_689,N_1397);
or U3754 (N_3754,N_479,N_1733);
nand U3755 (N_3755,N_373,N_1811);
or U3756 (N_3756,N_1554,N_756);
nand U3757 (N_3757,N_139,N_295);
or U3758 (N_3758,N_251,N_600);
nand U3759 (N_3759,N_797,N_627);
or U3760 (N_3760,N_1269,N_352);
nand U3761 (N_3761,N_848,N_1742);
nand U3762 (N_3762,N_683,N_620);
and U3763 (N_3763,N_282,N_1623);
and U3764 (N_3764,N_1113,N_1444);
or U3765 (N_3765,N_348,N_675);
nor U3766 (N_3766,N_1332,N_1167);
and U3767 (N_3767,N_1493,N_1540);
nand U3768 (N_3768,N_266,N_1849);
nand U3769 (N_3769,N_1694,N_126);
nor U3770 (N_3770,N_1771,N_1634);
or U3771 (N_3771,N_1782,N_786);
or U3772 (N_3772,N_1281,N_1686);
and U3773 (N_3773,N_1916,N_1401);
or U3774 (N_3774,N_1687,N_1289);
or U3775 (N_3775,N_653,N_1352);
nor U3776 (N_3776,N_761,N_1582);
or U3777 (N_3777,N_1219,N_410);
and U3778 (N_3778,N_569,N_1238);
xor U3779 (N_3779,N_544,N_751);
or U3780 (N_3780,N_308,N_134);
nor U3781 (N_3781,N_1729,N_1263);
nand U3782 (N_3782,N_590,N_1371);
or U3783 (N_3783,N_913,N_1518);
nor U3784 (N_3784,N_1427,N_133);
nand U3785 (N_3785,N_541,N_227);
nand U3786 (N_3786,N_524,N_1566);
and U3787 (N_3787,N_366,N_269);
nand U3788 (N_3788,N_1263,N_1183);
nor U3789 (N_3789,N_732,N_1036);
and U3790 (N_3790,N_386,N_1035);
nand U3791 (N_3791,N_342,N_1412);
nand U3792 (N_3792,N_1375,N_1924);
or U3793 (N_3793,N_1851,N_702);
nor U3794 (N_3794,N_1346,N_181);
or U3795 (N_3795,N_1248,N_1112);
nand U3796 (N_3796,N_1666,N_150);
and U3797 (N_3797,N_528,N_1212);
and U3798 (N_3798,N_741,N_63);
and U3799 (N_3799,N_778,N_851);
or U3800 (N_3800,N_622,N_1132);
and U3801 (N_3801,N_578,N_1485);
or U3802 (N_3802,N_1509,N_1829);
and U3803 (N_3803,N_1909,N_43);
and U3804 (N_3804,N_1518,N_1007);
nand U3805 (N_3805,N_1453,N_790);
and U3806 (N_3806,N_1591,N_1451);
nor U3807 (N_3807,N_880,N_1024);
or U3808 (N_3808,N_1431,N_1834);
nor U3809 (N_3809,N_1528,N_151);
xnor U3810 (N_3810,N_784,N_998);
nor U3811 (N_3811,N_194,N_1461);
and U3812 (N_3812,N_769,N_469);
and U3813 (N_3813,N_782,N_137);
and U3814 (N_3814,N_856,N_1058);
nand U3815 (N_3815,N_355,N_638);
nor U3816 (N_3816,N_1402,N_1487);
nor U3817 (N_3817,N_1651,N_677);
and U3818 (N_3818,N_1949,N_134);
or U3819 (N_3819,N_308,N_1798);
nand U3820 (N_3820,N_532,N_1537);
nor U3821 (N_3821,N_1969,N_1835);
or U3822 (N_3822,N_1370,N_1300);
and U3823 (N_3823,N_313,N_399);
nand U3824 (N_3824,N_852,N_974);
and U3825 (N_3825,N_894,N_1532);
nand U3826 (N_3826,N_1088,N_190);
or U3827 (N_3827,N_1495,N_1654);
or U3828 (N_3828,N_267,N_1079);
or U3829 (N_3829,N_560,N_1420);
and U3830 (N_3830,N_1289,N_1428);
and U3831 (N_3831,N_1392,N_1741);
nor U3832 (N_3832,N_1388,N_257);
nand U3833 (N_3833,N_1005,N_91);
nand U3834 (N_3834,N_1862,N_1484);
nand U3835 (N_3835,N_1767,N_1197);
or U3836 (N_3836,N_1643,N_1159);
or U3837 (N_3837,N_1526,N_214);
nor U3838 (N_3838,N_1410,N_618);
xnor U3839 (N_3839,N_697,N_1146);
nor U3840 (N_3840,N_1117,N_1614);
nor U3841 (N_3841,N_1034,N_1846);
or U3842 (N_3842,N_908,N_1335);
nor U3843 (N_3843,N_724,N_1796);
xor U3844 (N_3844,N_925,N_884);
xor U3845 (N_3845,N_706,N_99);
nand U3846 (N_3846,N_421,N_174);
nor U3847 (N_3847,N_1700,N_298);
or U3848 (N_3848,N_1242,N_1653);
nor U3849 (N_3849,N_1418,N_1033);
or U3850 (N_3850,N_1216,N_1720);
nand U3851 (N_3851,N_1061,N_738);
or U3852 (N_3852,N_1872,N_536);
nand U3853 (N_3853,N_409,N_299);
nor U3854 (N_3854,N_80,N_1957);
nor U3855 (N_3855,N_8,N_217);
and U3856 (N_3856,N_1595,N_673);
or U3857 (N_3857,N_1734,N_343);
nand U3858 (N_3858,N_34,N_1630);
and U3859 (N_3859,N_533,N_134);
nand U3860 (N_3860,N_231,N_1388);
nor U3861 (N_3861,N_819,N_928);
nor U3862 (N_3862,N_187,N_1635);
nand U3863 (N_3863,N_275,N_1169);
nand U3864 (N_3864,N_1497,N_873);
nand U3865 (N_3865,N_940,N_319);
and U3866 (N_3866,N_699,N_297);
nor U3867 (N_3867,N_1714,N_1046);
nand U3868 (N_3868,N_1071,N_1432);
nor U3869 (N_3869,N_894,N_1599);
and U3870 (N_3870,N_197,N_1658);
nor U3871 (N_3871,N_565,N_168);
and U3872 (N_3872,N_1788,N_659);
nand U3873 (N_3873,N_360,N_447);
nor U3874 (N_3874,N_1726,N_159);
nor U3875 (N_3875,N_1904,N_135);
nand U3876 (N_3876,N_863,N_786);
or U3877 (N_3877,N_1409,N_865);
nand U3878 (N_3878,N_375,N_525);
or U3879 (N_3879,N_1157,N_1512);
nor U3880 (N_3880,N_1034,N_732);
nand U3881 (N_3881,N_1328,N_1691);
nand U3882 (N_3882,N_1385,N_772);
or U3883 (N_3883,N_1365,N_862);
and U3884 (N_3884,N_1377,N_248);
or U3885 (N_3885,N_1692,N_1420);
nand U3886 (N_3886,N_986,N_1493);
nand U3887 (N_3887,N_479,N_1521);
nand U3888 (N_3888,N_1132,N_503);
nor U3889 (N_3889,N_815,N_1253);
nor U3890 (N_3890,N_1164,N_1371);
xor U3891 (N_3891,N_18,N_1442);
and U3892 (N_3892,N_219,N_888);
nor U3893 (N_3893,N_1685,N_1301);
or U3894 (N_3894,N_873,N_915);
and U3895 (N_3895,N_573,N_1232);
or U3896 (N_3896,N_893,N_1417);
nor U3897 (N_3897,N_1233,N_792);
or U3898 (N_3898,N_1146,N_1156);
nor U3899 (N_3899,N_583,N_544);
and U3900 (N_3900,N_1382,N_291);
nor U3901 (N_3901,N_461,N_980);
and U3902 (N_3902,N_341,N_1877);
and U3903 (N_3903,N_1832,N_1069);
nand U3904 (N_3904,N_438,N_98);
nand U3905 (N_3905,N_979,N_1054);
nand U3906 (N_3906,N_1286,N_121);
nor U3907 (N_3907,N_295,N_1269);
nand U3908 (N_3908,N_447,N_1812);
or U3909 (N_3909,N_820,N_36);
or U3910 (N_3910,N_1718,N_1222);
nor U3911 (N_3911,N_1192,N_1161);
or U3912 (N_3912,N_260,N_560);
nor U3913 (N_3913,N_547,N_356);
or U3914 (N_3914,N_1151,N_921);
or U3915 (N_3915,N_1759,N_1796);
nor U3916 (N_3916,N_773,N_1101);
nor U3917 (N_3917,N_807,N_802);
and U3918 (N_3918,N_1857,N_503);
or U3919 (N_3919,N_1001,N_963);
nor U3920 (N_3920,N_944,N_1186);
and U3921 (N_3921,N_1908,N_1783);
xnor U3922 (N_3922,N_119,N_128);
nand U3923 (N_3923,N_58,N_615);
and U3924 (N_3924,N_454,N_1033);
and U3925 (N_3925,N_1958,N_258);
and U3926 (N_3926,N_1908,N_1274);
and U3927 (N_3927,N_752,N_207);
and U3928 (N_3928,N_498,N_804);
and U3929 (N_3929,N_1063,N_974);
and U3930 (N_3930,N_1780,N_1667);
and U3931 (N_3931,N_1250,N_936);
or U3932 (N_3932,N_110,N_1804);
nor U3933 (N_3933,N_949,N_396);
nand U3934 (N_3934,N_1432,N_1272);
nand U3935 (N_3935,N_1888,N_1107);
nand U3936 (N_3936,N_632,N_1436);
or U3937 (N_3937,N_1845,N_1802);
or U3938 (N_3938,N_1963,N_305);
or U3939 (N_3939,N_1205,N_222);
and U3940 (N_3940,N_1125,N_1929);
and U3941 (N_3941,N_1601,N_755);
and U3942 (N_3942,N_1563,N_101);
or U3943 (N_3943,N_1188,N_994);
nor U3944 (N_3944,N_1362,N_204);
nand U3945 (N_3945,N_559,N_349);
nor U3946 (N_3946,N_1445,N_518);
nand U3947 (N_3947,N_1496,N_521);
nor U3948 (N_3948,N_1474,N_704);
nand U3949 (N_3949,N_992,N_1754);
or U3950 (N_3950,N_1963,N_711);
nand U3951 (N_3951,N_1999,N_1682);
and U3952 (N_3952,N_347,N_11);
nor U3953 (N_3953,N_1454,N_1568);
or U3954 (N_3954,N_1362,N_129);
or U3955 (N_3955,N_490,N_175);
nand U3956 (N_3956,N_136,N_1788);
nor U3957 (N_3957,N_912,N_242);
or U3958 (N_3958,N_1517,N_576);
and U3959 (N_3959,N_1071,N_1755);
or U3960 (N_3960,N_1857,N_704);
nor U3961 (N_3961,N_171,N_1780);
nor U3962 (N_3962,N_1589,N_1218);
nor U3963 (N_3963,N_147,N_1785);
nand U3964 (N_3964,N_1427,N_69);
nor U3965 (N_3965,N_1306,N_1375);
nand U3966 (N_3966,N_1935,N_277);
and U3967 (N_3967,N_346,N_1448);
nand U3968 (N_3968,N_288,N_136);
or U3969 (N_3969,N_1640,N_64);
nand U3970 (N_3970,N_1589,N_1906);
and U3971 (N_3971,N_857,N_1510);
or U3972 (N_3972,N_369,N_1412);
and U3973 (N_3973,N_106,N_1207);
nor U3974 (N_3974,N_658,N_1917);
or U3975 (N_3975,N_540,N_369);
and U3976 (N_3976,N_1781,N_1191);
nor U3977 (N_3977,N_696,N_646);
and U3978 (N_3978,N_1708,N_1457);
or U3979 (N_3979,N_1835,N_1386);
nand U3980 (N_3980,N_1879,N_1838);
and U3981 (N_3981,N_1240,N_408);
nor U3982 (N_3982,N_968,N_187);
or U3983 (N_3983,N_1699,N_1988);
nand U3984 (N_3984,N_36,N_1579);
nor U3985 (N_3985,N_411,N_888);
nand U3986 (N_3986,N_1401,N_1564);
and U3987 (N_3987,N_1391,N_1935);
nor U3988 (N_3988,N_1075,N_751);
nor U3989 (N_3989,N_575,N_208);
nor U3990 (N_3990,N_1404,N_338);
or U3991 (N_3991,N_1342,N_1459);
nand U3992 (N_3992,N_1820,N_1651);
or U3993 (N_3993,N_1850,N_30);
and U3994 (N_3994,N_1654,N_1693);
nand U3995 (N_3995,N_1783,N_1417);
nor U3996 (N_3996,N_1472,N_1889);
nand U3997 (N_3997,N_1040,N_878);
and U3998 (N_3998,N_233,N_425);
and U3999 (N_3999,N_1972,N_686);
nand U4000 (N_4000,N_3654,N_3319);
or U4001 (N_4001,N_2572,N_2714);
nor U4002 (N_4002,N_3786,N_3927);
nor U4003 (N_4003,N_3692,N_2448);
or U4004 (N_4004,N_2590,N_3346);
and U4005 (N_4005,N_3584,N_3945);
or U4006 (N_4006,N_2452,N_2753);
or U4007 (N_4007,N_3822,N_2420);
nor U4008 (N_4008,N_2567,N_3394);
nand U4009 (N_4009,N_2256,N_3116);
nor U4010 (N_4010,N_3600,N_2973);
or U4011 (N_4011,N_3196,N_2806);
and U4012 (N_4012,N_2575,N_2770);
or U4013 (N_4013,N_3241,N_2199);
nor U4014 (N_4014,N_2493,N_3579);
and U4015 (N_4015,N_2334,N_3976);
and U4016 (N_4016,N_3258,N_3094);
or U4017 (N_4017,N_3146,N_3256);
or U4018 (N_4018,N_3881,N_3973);
and U4019 (N_4019,N_2805,N_3395);
nor U4020 (N_4020,N_2869,N_2369);
and U4021 (N_4021,N_3819,N_3040);
nor U4022 (N_4022,N_2482,N_3556);
nor U4023 (N_4023,N_3087,N_2297);
nand U4024 (N_4024,N_2883,N_2060);
nand U4025 (N_4025,N_2579,N_2386);
or U4026 (N_4026,N_3707,N_2103);
or U4027 (N_4027,N_2155,N_3598);
and U4028 (N_4028,N_3417,N_3679);
and U4029 (N_4029,N_2004,N_3029);
nor U4030 (N_4030,N_2915,N_2043);
or U4031 (N_4031,N_3179,N_2121);
and U4032 (N_4032,N_3864,N_3495);
nand U4033 (N_4033,N_2917,N_3035);
xnor U4034 (N_4034,N_3878,N_2732);
nand U4035 (N_4035,N_2023,N_3203);
and U4036 (N_4036,N_2472,N_3139);
nand U4037 (N_4037,N_2494,N_2135);
nand U4038 (N_4038,N_3624,N_3308);
or U4039 (N_4039,N_2412,N_2694);
nand U4040 (N_4040,N_3709,N_3371);
or U4041 (N_4041,N_3360,N_2514);
or U4042 (N_4042,N_2440,N_3657);
and U4043 (N_4043,N_3675,N_2641);
or U4044 (N_4044,N_2588,N_3633);
nor U4045 (N_4045,N_3861,N_3820);
nor U4046 (N_4046,N_3583,N_3772);
or U4047 (N_4047,N_2849,N_2112);
and U4048 (N_4048,N_2381,N_2008);
nor U4049 (N_4049,N_2231,N_2290);
nand U4050 (N_4050,N_2524,N_2578);
and U4051 (N_4051,N_3586,N_2106);
nor U4052 (N_4052,N_3199,N_2128);
nand U4053 (N_4053,N_3362,N_2619);
nand U4054 (N_4054,N_2266,N_3745);
and U4055 (N_4055,N_2158,N_2115);
nor U4056 (N_4056,N_3970,N_3984);
and U4057 (N_4057,N_3949,N_2082);
xnor U4058 (N_4058,N_3374,N_2267);
nand U4059 (N_4059,N_2337,N_2505);
or U4060 (N_4060,N_3439,N_3158);
and U4061 (N_4061,N_2400,N_2399);
nor U4062 (N_4062,N_3272,N_2916);
nand U4063 (N_4063,N_3212,N_3160);
and U4064 (N_4064,N_2413,N_2767);
nand U4065 (N_4065,N_3658,N_3079);
or U4066 (N_4066,N_2855,N_2913);
nor U4067 (N_4067,N_3390,N_3687);
nand U4068 (N_4068,N_3490,N_3553);
nand U4069 (N_4069,N_2015,N_3218);
or U4070 (N_4070,N_3313,N_2934);
nor U4071 (N_4071,N_2397,N_2327);
or U4072 (N_4072,N_3081,N_2954);
or U4073 (N_4073,N_2117,N_3236);
nor U4074 (N_4074,N_3150,N_2515);
nor U4075 (N_4075,N_3255,N_2224);
nand U4076 (N_4076,N_2678,N_2792);
nor U4077 (N_4077,N_3427,N_2722);
nor U4078 (N_4078,N_3876,N_3612);
or U4079 (N_4079,N_2238,N_3232);
nor U4080 (N_4080,N_2891,N_2316);
nor U4081 (N_4081,N_3590,N_3428);
and U4082 (N_4082,N_2846,N_3110);
nand U4083 (N_4083,N_2387,N_2690);
or U4084 (N_4084,N_2245,N_2374);
or U4085 (N_4085,N_2250,N_3606);
nor U4086 (N_4086,N_2780,N_3036);
nand U4087 (N_4087,N_2312,N_3183);
and U4088 (N_4088,N_2888,N_3863);
nand U4089 (N_4089,N_3172,N_3726);
nand U4090 (N_4090,N_3339,N_3091);
nor U4091 (N_4091,N_3473,N_3266);
and U4092 (N_4092,N_2286,N_2313);
nand U4093 (N_4093,N_2603,N_2003);
nor U4094 (N_4094,N_2717,N_2630);
nor U4095 (N_4095,N_2563,N_3985);
and U4096 (N_4096,N_3460,N_2396);
nor U4097 (N_4097,N_2465,N_3135);
nor U4098 (N_4098,N_3959,N_2914);
nand U4099 (N_4099,N_2812,N_3324);
nor U4100 (N_4100,N_2584,N_2686);
nor U4101 (N_4101,N_3813,N_2942);
and U4102 (N_4102,N_3857,N_2451);
and U4103 (N_4103,N_2086,N_3835);
and U4104 (N_4104,N_3092,N_3049);
nand U4105 (N_4105,N_2002,N_2293);
nand U4106 (N_4106,N_3044,N_2701);
or U4107 (N_4107,N_3787,N_3830);
and U4108 (N_4108,N_3843,N_2994);
or U4109 (N_4109,N_2054,N_2168);
nor U4110 (N_4110,N_3301,N_3210);
or U4111 (N_4111,N_3983,N_2956);
nand U4112 (N_4112,N_3373,N_3570);
or U4113 (N_4113,N_3481,N_2191);
nor U4114 (N_4114,N_2298,N_2443);
and U4115 (N_4115,N_2618,N_3603);
and U4116 (N_4116,N_3856,N_2164);
and U4117 (N_4117,N_2719,N_3560);
or U4118 (N_4118,N_2657,N_3765);
or U4119 (N_4119,N_3462,N_3482);
xnor U4120 (N_4120,N_2670,N_3415);
nor U4121 (N_4121,N_3444,N_2402);
nand U4122 (N_4122,N_2393,N_2063);
or U4123 (N_4123,N_2787,N_3803);
or U4124 (N_4124,N_2559,N_2895);
nand U4125 (N_4125,N_3205,N_2172);
and U4126 (N_4126,N_3350,N_3790);
nor U4127 (N_4127,N_2309,N_3464);
xnor U4128 (N_4128,N_3454,N_2553);
and U4129 (N_4129,N_3562,N_3076);
nor U4130 (N_4130,N_2186,N_3678);
nor U4131 (N_4131,N_2308,N_2639);
nand U4132 (N_4132,N_2148,N_3320);
and U4133 (N_4133,N_3702,N_3154);
nor U4134 (N_4134,N_2940,N_3963);
and U4135 (N_4135,N_2088,N_2808);
nand U4136 (N_4136,N_2113,N_2742);
nand U4137 (N_4137,N_2348,N_2009);
nand U4138 (N_4138,N_3396,N_2543);
nor U4139 (N_4139,N_2344,N_2053);
nand U4140 (N_4140,N_2646,N_2713);
and U4141 (N_4141,N_2281,N_2886);
nand U4142 (N_4142,N_3795,N_3336);
nand U4143 (N_4143,N_2785,N_3997);
and U4144 (N_4144,N_2189,N_3144);
xnor U4145 (N_4145,N_3222,N_2810);
nor U4146 (N_4146,N_3870,N_2061);
nand U4147 (N_4147,N_3892,N_2017);
and U4148 (N_4148,N_3214,N_2119);
and U4149 (N_4149,N_3342,N_2398);
xor U4150 (N_4150,N_3652,N_2633);
nor U4151 (N_4151,N_2236,N_2253);
and U4152 (N_4152,N_2304,N_3451);
or U4153 (N_4153,N_3867,N_2361);
or U4154 (N_4154,N_2907,N_2987);
or U4155 (N_4155,N_2391,N_2547);
nand U4156 (N_4156,N_3541,N_3750);
nor U4157 (N_4157,N_3289,N_2985);
or U4158 (N_4158,N_2969,N_2663);
and U4159 (N_4159,N_2232,N_3178);
nand U4160 (N_4160,N_3185,N_3215);
nor U4161 (N_4161,N_2356,N_2190);
or U4162 (N_4162,N_2279,N_3884);
or U4163 (N_4163,N_3838,N_3351);
nand U4164 (N_4164,N_3851,N_3779);
or U4165 (N_4165,N_2066,N_2209);
and U4166 (N_4166,N_3906,N_3907);
and U4167 (N_4167,N_3776,N_3459);
nor U4168 (N_4168,N_3502,N_3964);
or U4169 (N_4169,N_3340,N_2275);
or U4170 (N_4170,N_2163,N_2542);
nor U4171 (N_4171,N_3596,N_2634);
nor U4172 (N_4172,N_2950,N_3620);
nand U4173 (N_4173,N_2020,N_2496);
nand U4174 (N_4174,N_2703,N_3519);
or U4175 (N_4175,N_2478,N_2471);
or U4176 (N_4176,N_3228,N_3254);
nand U4177 (N_4177,N_3968,N_2607);
nand U4178 (N_4178,N_2372,N_3510);
and U4179 (N_4179,N_2779,N_3500);
nand U4180 (N_4180,N_3085,N_3602);
nor U4181 (N_4181,N_3499,N_3257);
and U4182 (N_4182,N_3170,N_3405);
and U4183 (N_4183,N_3694,N_2574);
nor U4184 (N_4184,N_2140,N_2355);
or U4185 (N_4185,N_2264,N_2754);
nand U4186 (N_4186,N_2062,N_3735);
nand U4187 (N_4187,N_3681,N_3914);
and U4188 (N_4188,N_2414,N_3032);
and U4189 (N_4189,N_3849,N_2893);
nor U4190 (N_4190,N_2375,N_2509);
or U4191 (N_4191,N_2027,N_2594);
and U4192 (N_4192,N_2675,N_2098);
nand U4193 (N_4193,N_2862,N_3465);
or U4194 (N_4194,N_2876,N_2890);
nor U4195 (N_4195,N_2724,N_2145);
or U4196 (N_4196,N_3385,N_2255);
and U4197 (N_4197,N_3453,N_3994);
and U4198 (N_4198,N_3089,N_2160);
or U4199 (N_4199,N_3124,N_3470);
nand U4200 (N_4200,N_2814,N_2022);
or U4201 (N_4201,N_3788,N_3563);
nor U4202 (N_4202,N_3552,N_2909);
and U4203 (N_4203,N_2852,N_2137);
nor U4204 (N_4204,N_3662,N_2360);
nand U4205 (N_4205,N_2674,N_2406);
and U4206 (N_4206,N_3516,N_2366);
nand U4207 (N_4207,N_2211,N_3523);
and U4208 (N_4208,N_2798,N_3548);
and U4209 (N_4209,N_2395,N_2188);
and U4210 (N_4210,N_3733,N_2863);
and U4211 (N_4211,N_2616,N_2651);
and U4212 (N_4212,N_2442,N_2995);
nand U4213 (N_4213,N_3007,N_3068);
and U4214 (N_4214,N_2101,N_3644);
or U4215 (N_4215,N_2492,N_2200);
or U4216 (N_4216,N_3167,N_3078);
and U4217 (N_4217,N_2453,N_2411);
nand U4218 (N_4218,N_2433,N_3278);
and U4219 (N_4219,N_2169,N_3645);
and U4220 (N_4220,N_2303,N_2735);
nand U4221 (N_4221,N_2242,N_3375);
and U4222 (N_4222,N_3794,N_2625);
and U4223 (N_4223,N_3842,N_3151);
nand U4224 (N_4224,N_2367,N_2766);
and U4225 (N_4225,N_2282,N_3656);
nand U4226 (N_4226,N_2394,N_2809);
nand U4227 (N_4227,N_3780,N_3286);
nand U4228 (N_4228,N_2860,N_2599);
or U4229 (N_4229,N_3069,N_2006);
and U4230 (N_4230,N_3555,N_3609);
nor U4231 (N_4231,N_3245,N_3920);
nor U4232 (N_4232,N_2997,N_2796);
nor U4233 (N_4233,N_3659,N_2823);
or U4234 (N_4234,N_2908,N_3941);
or U4235 (N_4235,N_2564,N_3288);
or U4236 (N_4236,N_3230,N_3244);
nor U4237 (N_4237,N_3275,N_2070);
nand U4238 (N_4238,N_3507,N_2447);
or U4239 (N_4239,N_3104,N_2235);
nand U4240 (N_4240,N_2981,N_2929);
or U4241 (N_4241,N_3243,N_3883);
nor U4242 (N_4242,N_3897,N_3568);
and U4243 (N_4243,N_2300,N_3270);
or U4244 (N_4244,N_3446,N_3448);
nor U4245 (N_4245,N_2602,N_3751);
and U4246 (N_4246,N_2432,N_2270);
and U4247 (N_4247,N_3386,N_3996);
nor U4248 (N_4248,N_2058,N_3877);
nor U4249 (N_4249,N_2436,N_2130);
or U4250 (N_4250,N_3269,N_3753);
nor U4251 (N_4251,N_2044,N_3489);
nand U4252 (N_4252,N_3743,N_2228);
nor U4253 (N_4253,N_2382,N_3281);
nand U4254 (N_4254,N_3755,N_2935);
nand U4255 (N_4255,N_2426,N_2109);
nand U4256 (N_4256,N_3058,N_2632);
or U4257 (N_4257,N_2434,N_3117);
and U4258 (N_4258,N_3280,N_2610);
or U4259 (N_4259,N_2655,N_3801);
nand U4260 (N_4260,N_2133,N_3220);
nand U4261 (N_4261,N_3207,N_2029);
and U4262 (N_4262,N_3197,N_2198);
nor U4263 (N_4263,N_2193,N_3237);
nor U4264 (N_4264,N_3233,N_2152);
or U4265 (N_4265,N_2644,N_3194);
nor U4266 (N_4266,N_2497,N_2761);
nor U4267 (N_4267,N_2569,N_3223);
xnor U4268 (N_4268,N_3926,N_2181);
nor U4269 (N_4269,N_2662,N_3474);
nand U4270 (N_4270,N_2437,N_3588);
and U4271 (N_4271,N_3497,N_3629);
and U4272 (N_4272,N_3585,N_3296);
nand U4273 (N_4273,N_3824,N_2455);
xnor U4274 (N_4274,N_2491,N_2676);
or U4275 (N_4275,N_3231,N_2763);
nand U4276 (N_4276,N_2979,N_2800);
nand U4277 (N_4277,N_2949,N_2410);
and U4278 (N_4278,N_2107,N_2952);
and U4279 (N_4279,N_2955,N_2904);
and U4280 (N_4280,N_3971,N_2790);
or U4281 (N_4281,N_3325,N_3565);
or U4282 (N_4282,N_2507,N_3388);
and U4283 (N_4283,N_2582,N_3993);
nor U4284 (N_4284,N_2214,N_2899);
and U4285 (N_4285,N_2483,N_2839);
nand U4286 (N_4286,N_3334,N_2357);
nand U4287 (N_4287,N_3471,N_2331);
nand U4288 (N_4288,N_3761,N_2162);
nand U4289 (N_4289,N_2252,N_3577);
nand U4290 (N_4290,N_2278,N_3639);
nor U4291 (N_4291,N_3689,N_2537);
and U4292 (N_4292,N_2516,N_2990);
nor U4293 (N_4293,N_3125,N_3487);
nor U4294 (N_4294,N_3802,N_3498);
or U4295 (N_4295,N_3812,N_2404);
and U4296 (N_4296,N_3744,N_2457);
nor U4297 (N_4297,N_2338,N_2081);
or U4298 (N_4298,N_3521,N_3153);
or U4299 (N_4299,N_2998,N_3595);
and U4300 (N_4300,N_3770,N_2237);
nor U4301 (N_4301,N_3947,N_2332);
or U4302 (N_4302,N_2512,N_3890);
nor U4303 (N_4303,N_3111,N_3528);
or U4304 (N_4304,N_3328,N_3114);
nor U4305 (N_4305,N_3991,N_3628);
nor U4306 (N_4306,N_2336,N_3951);
nand U4307 (N_4307,N_3821,N_2882);
nor U4308 (N_4308,N_3918,N_3393);
nand U4309 (N_4309,N_2708,N_3274);
nand U4310 (N_4310,N_3152,N_3504);
and U4311 (N_4311,N_3859,N_3250);
nand U4312 (N_4312,N_2546,N_3756);
or U4313 (N_4313,N_2435,N_3251);
nor U4314 (N_4314,N_3611,N_2013);
nand U4315 (N_4315,N_3074,N_3730);
or U4316 (N_4316,N_2848,N_2967);
nor U4317 (N_4317,N_3549,N_2291);
nor U4318 (N_4318,N_2592,N_3224);
nand U4319 (N_4319,N_2803,N_2677);
nand U4320 (N_4320,N_2650,N_2626);
and U4321 (N_4321,N_3259,N_3804);
nor U4322 (N_4322,N_2288,N_3646);
nor U4323 (N_4323,N_2758,N_3773);
and U4324 (N_4324,N_3554,N_2554);
nand U4325 (N_4325,N_2851,N_2783);
nor U4326 (N_4326,N_2865,N_3691);
nor U4327 (N_4327,N_3435,N_3940);
and U4328 (N_4328,N_2016,N_2653);
or U4329 (N_4329,N_3705,N_3452);
and U4330 (N_4330,N_3913,N_2196);
and U4331 (N_4331,N_2185,N_2557);
or U4332 (N_4332,N_2744,N_2749);
nand U4333 (N_4333,N_3533,N_3356);
and U4334 (N_4334,N_3348,N_3902);
and U4335 (N_4335,N_2269,N_2802);
nor U4336 (N_4336,N_2697,N_3811);
and U4337 (N_4337,N_3397,N_2041);
nand U4338 (N_4338,N_3137,N_2544);
or U4339 (N_4339,N_3893,N_2521);
or U4340 (N_4340,N_3290,N_3642);
and U4341 (N_4341,N_3697,N_2740);
nor U4342 (N_4342,N_2832,N_3102);
or U4343 (N_4343,N_2551,N_2822);
and U4344 (N_4344,N_2794,N_2573);
nor U4345 (N_4345,N_2405,N_3043);
nand U4346 (N_4346,N_3948,N_3381);
and U4347 (N_4347,N_2833,N_2159);
or U4348 (N_4348,N_2652,N_3419);
and U4349 (N_4349,N_3347,N_2055);
nor U4350 (N_4350,N_2037,N_2474);
or U4351 (N_4351,N_2450,N_3685);
xnor U4352 (N_4352,N_3413,N_2039);
and U4353 (N_4353,N_2693,N_3888);
and U4354 (N_4354,N_2831,N_3209);
or U4355 (N_4355,N_3514,N_2654);
and U4356 (N_4356,N_3922,N_3925);
or U4357 (N_4357,N_2687,N_2216);
and U4358 (N_4358,N_3791,N_2248);
and U4359 (N_4359,N_3683,N_2799);
xor U4360 (N_4360,N_2084,N_2528);
or U4361 (N_4361,N_2064,N_3754);
nor U4362 (N_4362,N_2207,N_3370);
and U4363 (N_4363,N_2562,N_2089);
nand U4364 (N_4364,N_2861,N_2328);
nand U4365 (N_4365,N_2502,N_2151);
and U4366 (N_4366,N_2853,N_2068);
or U4367 (N_4367,N_3740,N_3412);
nor U4368 (N_4368,N_3736,N_3379);
or U4369 (N_4369,N_2598,N_2778);
and U4370 (N_4370,N_2215,N_3174);
or U4371 (N_4371,N_2841,N_3025);
nand U4372 (N_4372,N_2320,N_3840);
nor U4373 (N_4373,N_3165,N_3524);
and U4374 (N_4374,N_2102,N_2712);
and U4375 (N_4375,N_2684,N_3759);
or U4376 (N_4376,N_2533,N_2259);
and U4377 (N_4377,N_2685,N_2462);
and U4378 (N_4378,N_2820,N_2958);
nor U4379 (N_4379,N_3936,N_3852);
and U4380 (N_4380,N_3513,N_3002);
and U4381 (N_4381,N_2532,N_3706);
and U4382 (N_4382,N_3421,N_3739);
or U4383 (N_4383,N_3018,N_2510);
nand U4384 (N_4384,N_3901,N_3005);
nand U4385 (N_4385,N_2666,N_3714);
and U4386 (N_4386,N_3307,N_2018);
and U4387 (N_4387,N_3503,N_2739);
and U4388 (N_4388,N_3033,N_2073);
and U4389 (N_4389,N_2234,N_2217);
and U4390 (N_4390,N_2738,N_3001);
nand U4391 (N_4391,N_3099,N_2258);
and U4392 (N_4392,N_3335,N_2032);
nor U4393 (N_4393,N_2776,N_2460);
nor U4394 (N_4394,N_3935,N_2111);
or U4395 (N_4395,N_2341,N_3483);
and U4396 (N_4396,N_3661,N_2926);
or U4397 (N_4397,N_2146,N_2077);
and U4398 (N_4398,N_2425,N_3064);
xor U4399 (N_4399,N_3557,N_2774);
or U4400 (N_4400,N_3622,N_2479);
or U4401 (N_4401,N_2368,N_2993);
nand U4402 (N_4402,N_2745,N_2021);
and U4403 (N_4403,N_2920,N_2946);
or U4404 (N_4404,N_3211,N_2819);
nand U4405 (N_4405,N_3625,N_2506);
or U4406 (N_4406,N_2499,N_3987);
nor U4407 (N_4407,N_2226,N_3090);
and U4408 (N_4408,N_3760,N_3055);
nor U4409 (N_4409,N_3273,N_2762);
and U4410 (N_4410,N_3401,N_3267);
and U4411 (N_4411,N_2296,N_3509);
or U4412 (N_4412,N_3943,N_2292);
nor U4413 (N_4413,N_3376,N_2274);
and U4414 (N_4414,N_3827,N_3056);
and U4415 (N_4415,N_3293,N_3737);
nor U4416 (N_4416,N_3696,N_2518);
nand U4417 (N_4417,N_2354,N_2953);
nor U4418 (N_4418,N_3998,N_3879);
nand U4419 (N_4419,N_2477,N_2097);
and U4420 (N_4420,N_2568,N_3885);
xnor U4421 (N_4421,N_3778,N_3285);
xnor U4422 (N_4422,N_2301,N_2957);
and U4423 (N_4423,N_2600,N_3131);
nand U4424 (N_4424,N_3608,N_2912);
and U4425 (N_4425,N_3098,N_3853);
nand U4426 (N_4426,N_2409,N_2854);
nor U4427 (N_4427,N_3302,N_3575);
nor U4428 (N_4428,N_3723,N_2194);
nor U4429 (N_4429,N_2035,N_3905);
and U4430 (N_4430,N_2295,N_2636);
nor U4431 (N_4431,N_3133,N_3422);
or U4432 (N_4432,N_3956,N_3303);
nand U4433 (N_4433,N_3655,N_3643);
and U4434 (N_4434,N_3605,N_2683);
and U4435 (N_4435,N_3287,N_3443);
or U4436 (N_4436,N_2628,N_3392);
nor U4437 (N_4437,N_3545,N_2707);
or U4438 (N_4438,N_2977,N_3995);
nand U4439 (N_4439,N_2095,N_3792);
nand U4440 (N_4440,N_3311,N_3400);
nor U4441 (N_4441,N_3871,N_2184);
or U4442 (N_4442,N_3831,N_3900);
nand U4443 (N_4443,N_2750,N_3981);
nor U4444 (N_4444,N_3684,N_2114);
nor U4445 (N_4445,N_3796,N_3100);
or U4446 (N_4446,N_3669,N_2898);
or U4447 (N_4447,N_2970,N_2691);
or U4448 (N_4448,N_2183,N_2983);
or U4449 (N_4449,N_2788,N_2072);
or U4450 (N_4450,N_3869,N_3542);
and U4451 (N_4451,N_2991,N_3799);
or U4452 (N_4452,N_3986,N_2143);
nor U4453 (N_4453,N_2923,N_3717);
or U4454 (N_4454,N_3526,N_3316);
nand U4455 (N_4455,N_3967,N_3227);
nand U4456 (N_4456,N_3380,N_2129);
nand U4457 (N_4457,N_3132,N_2153);
xor U4458 (N_4458,N_3887,N_3420);
nand U4459 (N_4459,N_3982,N_3635);
nand U4460 (N_4460,N_3121,N_3195);
or U4461 (N_4461,N_3540,N_2019);
nor U4462 (N_4462,N_2647,N_3774);
nand U4463 (N_4463,N_3573,N_3671);
nand U4464 (N_4464,N_3718,N_2012);
nor U4465 (N_4465,N_2118,N_2422);
nor U4466 (N_4466,N_2595,N_3011);
or U4467 (N_4467,N_2052,N_2961);
nor U4468 (N_4468,N_3515,N_3546);
or U4469 (N_4469,N_3354,N_3080);
and U4470 (N_4470,N_3518,N_2461);
or U4471 (N_4471,N_2305,N_3202);
or U4472 (N_4472,N_3410,N_3953);
nor U4473 (N_4473,N_2527,N_3992);
or U4474 (N_4474,N_3187,N_2878);
or U4475 (N_4475,N_3701,N_3120);
nor U4476 (N_4476,N_2244,N_2495);
and U4477 (N_4477,N_3969,N_3372);
and U4478 (N_4478,N_2538,N_3587);
and U4479 (N_4479,N_2621,N_3660);
nand U4480 (N_4480,N_2727,N_2046);
nor U4481 (N_4481,N_2218,N_3365);
and U4482 (N_4482,N_2192,N_2091);
or U4483 (N_4483,N_3363,N_3028);
nand U4484 (N_4484,N_2866,N_2535);
nand U4485 (N_4485,N_2464,N_3979);
nand U4486 (N_4486,N_2508,N_3204);
nand U4487 (N_4487,N_2271,N_3283);
or U4488 (N_4488,N_3854,N_2556);
nor U4489 (N_4489,N_2195,N_3424);
nand U4490 (N_4490,N_3674,N_2658);
nand U4491 (N_4491,N_3466,N_3119);
nor U4492 (N_4492,N_3193,N_2793);
nand U4493 (N_4493,N_2604,N_3566);
and U4494 (N_4494,N_3829,N_2373);
nor U4495 (N_4495,N_3476,N_2597);
or U4496 (N_4496,N_2887,N_3279);
nand U4497 (N_4497,N_2287,N_3093);
nand U4498 (N_4498,N_2057,N_3013);
and U4499 (N_4499,N_3077,N_2416);
or U4500 (N_4500,N_3937,N_3065);
or U4501 (N_4501,N_2116,N_2660);
and U4502 (N_4502,N_2126,N_3837);
nand U4503 (N_4503,N_3637,N_2587);
nand U4504 (N_4504,N_2530,N_2265);
nor U4505 (N_4505,N_3075,N_2175);
or U4506 (N_4506,N_2080,N_2951);
and U4507 (N_4507,N_3108,N_2939);
nor U4508 (N_4508,N_2835,N_2385);
nand U4509 (N_4509,N_3818,N_2383);
or U4510 (N_4510,N_3698,N_3322);
nor U4511 (N_4511,N_2925,N_2005);
nand U4512 (N_4512,N_2444,N_3248);
nor U4513 (N_4513,N_2470,N_3648);
nand U4514 (N_4514,N_3781,N_2430);
nand U4515 (N_4515,N_2828,N_3014);
and U4516 (N_4516,N_2791,N_3809);
nand U4517 (N_4517,N_3980,N_3749);
nor U4518 (N_4518,N_3789,N_2813);
or U4519 (N_4519,N_3327,N_2672);
and U4520 (N_4520,N_2700,N_2306);
nor U4521 (N_4521,N_3072,N_3708);
nand U4522 (N_4522,N_2268,N_2388);
or U4523 (N_4523,N_3169,N_3988);
and U4524 (N_4524,N_3783,N_2576);
and U4525 (N_4525,N_3039,N_2486);
or U4526 (N_4526,N_3488,N_2001);
or U4527 (N_4527,N_2246,N_2601);
and U4528 (N_4528,N_2611,N_3965);
nor U4529 (N_4529,N_2901,N_2696);
nand U4530 (N_4530,N_2960,N_3298);
or U4531 (N_4531,N_2555,N_3306);
or U4532 (N_4532,N_3047,N_3067);
nor U4533 (N_4533,N_3221,N_2840);
xor U4534 (N_4534,N_2225,N_3581);
nor U4535 (N_4535,N_2826,N_2142);
or U4536 (N_4536,N_3962,N_2571);
and U4537 (N_4537,N_3358,N_2339);
and U4538 (N_4538,N_2468,N_3632);
and U4539 (N_4539,N_2902,N_3054);
or U4540 (N_4540,N_3295,N_3402);
or U4541 (N_4541,N_3768,N_3003);
nand U4542 (N_4542,N_3073,N_2821);
nand U4543 (N_4543,N_2706,N_2503);
and U4544 (N_4544,N_2475,N_2047);
and U4545 (N_4545,N_3578,N_3784);
and U4546 (N_4546,N_3725,N_2485);
and U4547 (N_4547,N_3836,N_2593);
or U4548 (N_4548,N_2702,N_2648);
and U4549 (N_4549,N_2423,N_3734);
nand U4550 (N_4550,N_2324,N_3173);
nand U4551 (N_4551,N_3384,N_3106);
nor U4552 (N_4552,N_2351,N_2272);
and U4553 (N_4553,N_2709,N_3141);
and U4554 (N_4554,N_2807,N_3242);
nand U4555 (N_4555,N_3323,N_2836);
nand U4556 (N_4556,N_2838,N_3024);
xnor U4557 (N_4557,N_2918,N_3235);
nand U4558 (N_4558,N_3923,N_2220);
and U4559 (N_4559,N_3957,N_2816);
nor U4560 (N_4560,N_2428,N_3710);
nand U4561 (N_4561,N_2138,N_3797);
and U4562 (N_4562,N_3928,N_3952);
nor U4563 (N_4563,N_3746,N_3265);
nand U4564 (N_4564,N_3716,N_2076);
and U4565 (N_4565,N_2536,N_3571);
and U4566 (N_4566,N_2056,N_3833);
and U4567 (N_4567,N_3479,N_2673);
and U4568 (N_4568,N_2065,N_3226);
nand U4569 (N_4569,N_2154,N_2733);
nand U4570 (N_4570,N_2131,N_3472);
or U4571 (N_4571,N_2877,N_3911);
nand U4572 (N_4572,N_2094,N_2105);
nand U4573 (N_4573,N_2896,N_2247);
and U4574 (N_4574,N_3742,N_2755);
nor U4575 (N_4575,N_3445,N_3162);
or U4576 (N_4576,N_3097,N_2980);
and U4577 (N_4577,N_2596,N_3525);
or U4578 (N_4578,N_3582,N_3343);
nor U4579 (N_4579,N_3668,N_3168);
or U4580 (N_4580,N_3592,N_3616);
nor U4581 (N_4581,N_3145,N_3200);
nand U4582 (N_4582,N_2318,N_2390);
nor U4583 (N_4583,N_2389,N_2850);
and U4584 (N_4584,N_3063,N_3184);
nand U4585 (N_4585,N_2623,N_3349);
nand U4586 (N_4586,N_2937,N_3798);
or U4587 (N_4587,N_3594,N_3337);
nor U4588 (N_4588,N_3627,N_3051);
nand U4589 (N_4589,N_2797,N_2384);
or U4590 (N_4590,N_2589,N_2311);
nand U4591 (N_4591,N_2906,N_3766);
nor U4592 (N_4592,N_3175,N_3636);
nand U4593 (N_4593,N_3297,N_2157);
or U4594 (N_4594,N_2622,N_2730);
nand U4595 (N_4595,N_3429,N_3874);
or U4596 (N_4596,N_3366,N_3359);
nand U4597 (N_4597,N_2459,N_2099);
or U4598 (N_4598,N_2811,N_3721);
nand U4599 (N_4599,N_2346,N_3478);
nor U4600 (N_4600,N_3387,N_3825);
or U4601 (N_4601,N_3599,N_2519);
and U4602 (N_4602,N_3107,N_3607);
and U4603 (N_4603,N_2302,N_3130);
and U4604 (N_4604,N_3216,N_2289);
and U4605 (N_4605,N_2033,N_2487);
nand U4606 (N_4606,N_2531,N_3404);
or U4607 (N_4607,N_3318,N_3999);
nand U4608 (N_4608,N_2407,N_2843);
nand U4609 (N_4609,N_3715,N_3008);
or U4610 (N_4610,N_2364,N_2050);
and U4611 (N_4611,N_2325,N_3597);
and U4612 (N_4612,N_3369,N_2698);
or U4613 (N_4613,N_3333,N_2227);
or U4614 (N_4614,N_2525,N_3461);
nor U4615 (N_4615,N_3208,N_3946);
nand U4616 (N_4616,N_3377,N_2729);
nand U4617 (N_4617,N_2469,N_2132);
and U4618 (N_4618,N_2962,N_3240);
and U4619 (N_4619,N_3496,N_2526);
nor U4620 (N_4620,N_3059,N_2210);
nor U4621 (N_4621,N_2233,N_2285);
nand U4622 (N_4622,N_3908,N_3517);
or U4623 (N_4623,N_3666,N_2294);
xor U4624 (N_4624,N_3576,N_2540);
nand U4625 (N_4625,N_3062,N_3041);
or U4626 (N_4626,N_2036,N_3865);
or U4627 (N_4627,N_2125,N_2680);
nand U4628 (N_4628,N_3699,N_3921);
nor U4629 (N_4629,N_2522,N_3574);
or U4630 (N_4630,N_3409,N_2731);
or U4631 (N_4631,N_3492,N_3939);
nand U4632 (N_4632,N_3663,N_3271);
nand U4633 (N_4633,N_3249,N_3045);
nor U4634 (N_4634,N_3128,N_3345);
and U4635 (N_4635,N_3206,N_2972);
nor U4636 (N_4636,N_3180,N_3475);
and U4637 (N_4637,N_2403,N_2030);
nand U4638 (N_4638,N_3673,N_2170);
nor U4639 (N_4639,N_2371,N_2643);
or U4640 (N_4640,N_2352,N_2280);
and U4641 (N_4641,N_2570,N_3793);
and U4642 (N_4642,N_2481,N_2379);
and U4643 (N_4643,N_2139,N_3338);
nor U4644 (N_4644,N_2645,N_2765);
nor U4645 (N_4645,N_2549,N_2859);
or U4646 (N_4646,N_3634,N_2667);
and U4647 (N_4647,N_2322,N_3621);
nor U4648 (N_4648,N_3930,N_3522);
nand U4649 (N_4649,N_3919,N_3505);
nor U4650 (N_4650,N_2347,N_3088);
nor U4651 (N_4651,N_3929,N_2071);
nand U4652 (N_4652,N_3367,N_3341);
nand U4653 (N_4653,N_2156,N_2775);
or U4654 (N_4654,N_3344,N_2656);
and U4655 (N_4655,N_3118,N_2545);
or U4656 (N_4656,N_3903,N_2038);
or U4657 (N_4657,N_3764,N_2362);
or U4658 (N_4658,N_3382,N_3695);
nor U4659 (N_4659,N_2769,N_3989);
or U4660 (N_4660,N_3434,N_2704);
nand U4661 (N_4661,N_3700,N_3974);
nor U4662 (N_4662,N_3456,N_3950);
nand U4663 (N_4663,N_2501,N_3752);
or U4664 (N_4664,N_2358,N_2439);
and U4665 (N_4665,N_3061,N_3618);
and U4666 (N_4666,N_2067,N_3060);
nor U4667 (N_4667,N_3531,N_3142);
nand U4668 (N_4668,N_2350,N_3713);
and U4669 (N_4669,N_3711,N_2837);
nand U4670 (N_4670,N_2202,N_2523);
and U4671 (N_4671,N_2931,N_3219);
nor U4672 (N_4672,N_3848,N_2083);
nor U4673 (N_4673,N_2307,N_3610);
nor U4674 (N_4674,N_3527,N_2873);
and U4675 (N_4675,N_3771,N_2069);
and U4676 (N_4676,N_2161,N_3807);
nand U4677 (N_4677,N_2858,N_3423);
nor U4678 (N_4678,N_2177,N_3190);
and U4679 (N_4679,N_3310,N_2517);
xnor U4680 (N_4680,N_3977,N_2842);
nand U4681 (N_4681,N_2326,N_3727);
nor U4682 (N_4682,N_2438,N_2705);
nor U4683 (N_4683,N_2342,N_3052);
nor U4684 (N_4684,N_3569,N_2617);
nor U4685 (N_4685,N_3955,N_2786);
and U4686 (N_4686,N_2947,N_2110);
nor U4687 (N_4687,N_2317,N_2174);
and U4688 (N_4688,N_2829,N_3425);
or U4689 (N_4689,N_3246,N_3192);
nand U4690 (N_4690,N_3757,N_3436);
and U4691 (N_4691,N_3785,N_2000);
nor U4692 (N_4692,N_2204,N_2445);
and U4693 (N_4693,N_2182,N_2550);
and U4694 (N_4694,N_2635,N_2480);
and U4695 (N_4695,N_2577,N_2614);
or U4696 (N_4696,N_3458,N_2206);
and U4697 (N_4697,N_3012,N_2606);
nand U4698 (N_4698,N_3547,N_2315);
or U4699 (N_4699,N_2370,N_2100);
and U4700 (N_4700,N_3449,N_3814);
and U4701 (N_4701,N_2028,N_3115);
nand U4702 (N_4702,N_2335,N_3832);
nor U4703 (N_4703,N_2884,N_2167);
xor U4704 (N_4704,N_3529,N_3494);
nand U4705 (N_4705,N_3688,N_2928);
and U4706 (N_4706,N_3966,N_3006);
nand U4707 (N_4707,N_3364,N_2345);
or U4708 (N_4708,N_3653,N_2449);
and U4709 (N_4709,N_2605,N_2795);
and U4710 (N_4710,N_3411,N_2948);
and U4711 (N_4711,N_3046,N_2631);
or U4712 (N_4712,N_3159,N_3305);
or U4713 (N_4713,N_2392,N_2007);
and U4714 (N_4714,N_2415,N_3640);
nor U4715 (N_4715,N_2134,N_3841);
or U4716 (N_4716,N_3748,N_3282);
nor U4717 (N_4717,N_2539,N_3407);
and U4718 (N_4718,N_2936,N_3769);
nor U4719 (N_4719,N_2757,N_2649);
nor U4720 (N_4720,N_3767,N_3638);
and U4721 (N_4721,N_3731,N_3850);
nor U4722 (N_4722,N_3613,N_2963);
or U4723 (N_4723,N_2429,N_3189);
or U4724 (N_4724,N_3667,N_2801);
and U4725 (N_4725,N_2203,N_2136);
or U4726 (N_4726,N_2728,N_2417);
nand U4727 (N_4727,N_2905,N_3844);
and U4728 (N_4728,N_2144,N_2048);
or U4729 (N_4729,N_3247,N_2197);
or U4730 (N_4730,N_3010,N_2964);
nor U4731 (N_4731,N_2711,N_2222);
and U4732 (N_4732,N_3467,N_3704);
nor U4733 (N_4733,N_2818,N_2699);
and U4734 (N_4734,N_3722,N_2176);
nand U4735 (N_4735,N_2892,N_3284);
and U4736 (N_4736,N_3960,N_2781);
nor U4737 (N_4737,N_3291,N_3493);
and U4738 (N_4738,N_3828,N_3543);
nor U4739 (N_4739,N_3882,N_3491);
or U4740 (N_4740,N_3558,N_3127);
or U4741 (N_4741,N_2695,N_2173);
nor U4742 (N_4742,N_2989,N_2205);
nor U4743 (N_4743,N_2511,N_2764);
and U4744 (N_4744,N_3846,N_3182);
and U4745 (N_4745,N_3469,N_3229);
or U4746 (N_4746,N_2353,N_2079);
and U4747 (N_4747,N_2378,N_3823);
or U4748 (N_4748,N_3623,N_3017);
nand U4749 (N_4749,N_3912,N_3191);
nor U4750 (N_4750,N_3664,N_2045);
nand U4751 (N_4751,N_2867,N_3747);
nand U4752 (N_4752,N_2971,N_2513);
and U4753 (N_4753,N_3399,N_3604);
and U4754 (N_4754,N_3866,N_3406);
or U4755 (N_4755,N_2424,N_3329);
nand U4756 (N_4756,N_3891,N_3872);
nor U4757 (N_4757,N_2223,N_3177);
nor U4758 (N_4758,N_2921,N_2718);
nand U4759 (N_4759,N_2747,N_3898);
nand U4760 (N_4760,N_3326,N_2299);
nand U4761 (N_4761,N_2418,N_2230);
and U4762 (N_4762,N_2585,N_3252);
or U4763 (N_4763,N_2243,N_2864);
nor U4764 (N_4764,N_3944,N_2534);
and U4765 (N_4765,N_3938,N_3020);
or U4766 (N_4766,N_2945,N_2903);
or U4767 (N_4767,N_2959,N_2212);
nand U4768 (N_4768,N_2988,N_2059);
or U4769 (N_4769,N_3277,N_2284);
or U4770 (N_4770,N_3138,N_2688);
nand U4771 (N_4771,N_2640,N_3140);
nand U4772 (N_4772,N_2376,N_2277);
and U4773 (N_4773,N_3082,N_2239);
and U4774 (N_4774,N_2974,N_2520);
and U4775 (N_4775,N_2500,N_3690);
or U4776 (N_4776,N_2498,N_3942);
nor U4777 (N_4777,N_2924,N_3631);
and U4778 (N_4778,N_3447,N_2910);
nand U4779 (N_4779,N_3317,N_2031);
nor U4780 (N_4780,N_2249,N_3855);
nand U4781 (N_4781,N_2548,N_3147);
nor U4782 (N_4782,N_2661,N_3719);
and U4783 (N_4783,N_2847,N_2241);
or U4784 (N_4784,N_2927,N_3084);
and U4785 (N_4785,N_3378,N_2087);
nand U4786 (N_4786,N_2456,N_3958);
or U4787 (N_4787,N_3086,N_3868);
xor U4788 (N_4788,N_3103,N_3321);
nand U4789 (N_4789,N_3122,N_2978);
nor U4790 (N_4790,N_2187,N_3225);
nor U4791 (N_4791,N_3239,N_3561);
and U4792 (N_4792,N_3300,N_2874);
nor U4793 (N_4793,N_3858,N_3896);
nor U4794 (N_4794,N_2171,N_2760);
or U4795 (N_4795,N_2560,N_2011);
and U4796 (N_4796,N_3276,N_2845);
or U4797 (N_4797,N_2219,N_2938);
nand U4798 (N_4798,N_3593,N_3164);
nor U4799 (N_4799,N_3758,N_3551);
or U4800 (N_4800,N_2772,N_2830);
and U4801 (N_4801,N_2986,N_3053);
or U4802 (N_4802,N_2992,N_3886);
nor U4803 (N_4803,N_3357,N_3263);
nor U4804 (N_4804,N_3782,N_3724);
nand U4805 (N_4805,N_3315,N_2736);
nand U4806 (N_4806,N_3042,N_2889);
nor U4807 (N_4807,N_2615,N_2489);
nand U4808 (N_4808,N_2127,N_2922);
xor U4809 (N_4809,N_3486,N_3129);
and U4810 (N_4810,N_2208,N_3847);
nor U4811 (N_4811,N_2871,N_2090);
nor U4812 (N_4812,N_3537,N_2932);
or U4813 (N_4813,N_3806,N_2789);
nand U4814 (N_4814,N_2897,N_3136);
nor U4815 (N_4815,N_2123,N_3862);
nor U4816 (N_4816,N_2040,N_3559);
nor U4817 (N_4817,N_2824,N_2900);
nand U4818 (N_4818,N_2671,N_2999);
nor U4819 (N_4819,N_2827,N_2982);
nor U4820 (N_4820,N_3070,N_3880);
nand U4821 (N_4821,N_3899,N_2725);
nor U4822 (N_4822,N_2365,N_3567);
nand U4823 (N_4823,N_2419,N_3016);
nor U4824 (N_4824,N_2609,N_2586);
nand U4825 (N_4825,N_3457,N_2723);
nand U4826 (N_4826,N_3815,N_2669);
nand U4827 (N_4827,N_2108,N_2310);
nand U4828 (N_4828,N_3171,N_3031);
nor U4829 (N_4829,N_3105,N_2363);
or U4830 (N_4830,N_2254,N_3641);
xor U4831 (N_4831,N_2933,N_3143);
and U4832 (N_4832,N_2668,N_2427);
nand U4833 (N_4833,N_2894,N_3331);
nand U4834 (N_4834,N_3030,N_3021);
or U4835 (N_4835,N_3589,N_3647);
nor U4836 (N_4836,N_3520,N_2682);
or U4837 (N_4837,N_2583,N_3176);
and U4838 (N_4838,N_2283,N_2319);
and U4839 (N_4839,N_2141,N_3431);
nor U4840 (N_4840,N_3463,N_2965);
and U4841 (N_4841,N_2166,N_3539);
and U4842 (N_4842,N_3860,N_3538);
and U4843 (N_4843,N_3720,N_3670);
and U4844 (N_4844,N_3975,N_3630);
xnor U4845 (N_4845,N_2276,N_3934);
or U4846 (N_4846,N_2458,N_3166);
and U4847 (N_4847,N_2637,N_2743);
nand U4848 (N_4848,N_2431,N_2463);
or U4849 (N_4849,N_3816,N_3213);
nor U4850 (N_4850,N_3383,N_3113);
nand U4851 (N_4851,N_2612,N_3038);
nand U4852 (N_4852,N_2042,N_3910);
and U4853 (N_4853,N_3353,N_2180);
nor U4854 (N_4854,N_2323,N_3198);
and U4855 (N_4855,N_3536,N_2741);
and U4856 (N_4856,N_2629,N_3455);
nand U4857 (N_4857,N_3101,N_2401);
nor U4858 (N_4858,N_3550,N_3954);
nor U4859 (N_4859,N_2026,N_3126);
or U4860 (N_4860,N_2608,N_3532);
or U4861 (N_4861,N_3112,N_2359);
and U4862 (N_4862,N_3264,N_2251);
nand U4863 (N_4863,N_2777,N_2104);
and U4864 (N_4864,N_3512,N_3057);
nand U4865 (N_4865,N_3149,N_2868);
nor U4866 (N_4866,N_3591,N_2446);
nor U4867 (N_4867,N_3535,N_3440);
and U4868 (N_4868,N_3015,N_3873);
nor U4869 (N_4869,N_2476,N_3665);
nand U4870 (N_4870,N_3019,N_2124);
nor U4871 (N_4871,N_3924,N_2782);
nand U4872 (N_4872,N_3330,N_3729);
and U4873 (N_4873,N_2857,N_2092);
or U4874 (N_4874,N_3438,N_3066);
or U4875 (N_4875,N_2529,N_3626);
and U4876 (N_4876,N_2147,N_3777);
or U4877 (N_4877,N_2591,N_2466);
nor U4878 (N_4878,N_3441,N_3732);
nor U4879 (N_4879,N_3834,N_3530);
and U4880 (N_4880,N_3234,N_3650);
or U4881 (N_4881,N_3805,N_3693);
or U4882 (N_4882,N_2804,N_3161);
nor U4883 (N_4883,N_2642,N_2025);
and U4884 (N_4884,N_2490,N_3501);
or U4885 (N_4885,N_2966,N_3268);
or U4886 (N_4886,N_2710,N_2078);
nor U4887 (N_4887,N_3889,N_2380);
or U4888 (N_4888,N_3292,N_3450);
or U4889 (N_4889,N_3601,N_2221);
nor U4890 (N_4890,N_2488,N_3416);
nand U4891 (N_4891,N_2049,N_3808);
and U4892 (N_4892,N_2150,N_2261);
and U4893 (N_4893,N_3817,N_3294);
or U4894 (N_4894,N_2880,N_2201);
and U4895 (N_4895,N_2257,N_2638);
and U4896 (N_4896,N_3253,N_2165);
nor U4897 (N_4897,N_3095,N_3534);
nand U4898 (N_4898,N_3403,N_3123);
nand U4899 (N_4899,N_3186,N_3299);
and U4900 (N_4900,N_2996,N_3261);
nand U4901 (N_4901,N_3728,N_2720);
nor U4902 (N_4902,N_2751,N_2122);
nand U4903 (N_4903,N_3580,N_3916);
or U4904 (N_4904,N_2581,N_2784);
nand U4905 (N_4905,N_3651,N_3426);
and U4906 (N_4906,N_3238,N_3572);
nand U4907 (N_4907,N_2093,N_2834);
nand U4908 (N_4908,N_2885,N_3484);
nor U4909 (N_4909,N_2120,N_3917);
or U4910 (N_4910,N_3649,N_3430);
nor U4911 (N_4911,N_3022,N_2349);
or U4912 (N_4912,N_2504,N_2875);
xor U4913 (N_4913,N_2343,N_2748);
and U4914 (N_4914,N_3050,N_3026);
and U4915 (N_4915,N_2976,N_3355);
nor U4916 (N_4916,N_3437,N_3800);
and U4917 (N_4917,N_2930,N_2919);
or U4918 (N_4918,N_2229,N_3932);
or U4919 (N_4919,N_2815,N_3260);
or U4920 (N_4920,N_3480,N_2484);
nor U4921 (N_4921,N_3931,N_3000);
nand U4922 (N_4922,N_3304,N_3712);
nor U4923 (N_4923,N_3368,N_3511);
and U4924 (N_4924,N_2262,N_3680);
nor U4925 (N_4925,N_2941,N_2178);
and U4926 (N_4926,N_3083,N_3686);
nand U4927 (N_4927,N_3309,N_2421);
and U4928 (N_4928,N_3361,N_3762);
nor U4929 (N_4929,N_3477,N_3071);
or U4930 (N_4930,N_2870,N_3544);
or U4931 (N_4931,N_2075,N_2737);
nor U4932 (N_4932,N_2975,N_3352);
and U4933 (N_4933,N_3109,N_2825);
or U4934 (N_4934,N_3037,N_2541);
nor U4935 (N_4935,N_3619,N_3027);
or U4936 (N_4936,N_3741,N_2340);
nand U4937 (N_4937,N_3672,N_3508);
and U4938 (N_4938,N_2240,N_3048);
or U4939 (N_4939,N_2314,N_2689);
nand U4940 (N_4940,N_2943,N_2014);
nor U4941 (N_4941,N_3312,N_3763);
or U4942 (N_4942,N_2879,N_3096);
or U4943 (N_4943,N_2329,N_2179);
and U4944 (N_4944,N_2726,N_3398);
nor U4945 (N_4945,N_2664,N_2817);
and U4946 (N_4946,N_2968,N_2273);
xnor U4947 (N_4947,N_3990,N_3775);
and U4948 (N_4948,N_3433,N_2213);
or U4949 (N_4949,N_2565,N_3617);
nor U4950 (N_4950,N_3738,N_3262);
or U4951 (N_4951,N_2984,N_3615);
nand U4952 (N_4952,N_3023,N_3839);
or U4953 (N_4953,N_3895,N_3432);
or U4954 (N_4954,N_2665,N_2681);
or U4955 (N_4955,N_2771,N_3134);
nor U4956 (N_4956,N_2552,N_2911);
nand U4957 (N_4957,N_3676,N_2715);
nor U4958 (N_4958,N_2149,N_2085);
nor U4959 (N_4959,N_2566,N_2944);
or U4960 (N_4960,N_3677,N_3408);
and U4961 (N_4961,N_3156,N_2051);
nand U4962 (N_4962,N_2679,N_3217);
nor U4963 (N_4963,N_2856,N_3009);
and U4964 (N_4964,N_2330,N_2034);
nand U4965 (N_4965,N_2624,N_2321);
or U4966 (N_4966,N_2692,N_2010);
and U4967 (N_4967,N_2659,N_2721);
nand U4968 (N_4968,N_3810,N_3414);
or U4969 (N_4969,N_2408,N_3909);
nor U4970 (N_4970,N_3485,N_2467);
or U4971 (N_4971,N_3978,N_2580);
nor U4972 (N_4972,N_3155,N_2613);
nand U4973 (N_4973,N_3826,N_2759);
nor U4974 (N_4974,N_2260,N_3894);
and U4975 (N_4975,N_3682,N_2333);
or U4976 (N_4976,N_2768,N_2844);
nor U4977 (N_4977,N_2558,N_2872);
nor U4978 (N_4978,N_3181,N_2773);
nor U4979 (N_4979,N_3468,N_3442);
nand U4980 (N_4980,N_2881,N_3201);
nand U4981 (N_4981,N_2454,N_3004);
nand U4982 (N_4982,N_2752,N_3391);
nor U4983 (N_4983,N_3933,N_2561);
or U4984 (N_4984,N_3972,N_3614);
and U4985 (N_4985,N_2756,N_3961);
and U4986 (N_4986,N_2620,N_2024);
or U4987 (N_4987,N_3703,N_3875);
or U4988 (N_4988,N_2627,N_3418);
nand U4989 (N_4989,N_3564,N_3314);
nand U4990 (N_4990,N_2074,N_2263);
nand U4991 (N_4991,N_3332,N_3157);
or U4992 (N_4992,N_3188,N_3915);
or U4993 (N_4993,N_2746,N_2473);
nand U4994 (N_4994,N_2441,N_3163);
or U4995 (N_4995,N_3034,N_3904);
nand U4996 (N_4996,N_3148,N_3845);
nor U4997 (N_4997,N_2096,N_3506);
nor U4998 (N_4998,N_2377,N_3389);
nor U4999 (N_4999,N_2734,N_2716);
or U5000 (N_5000,N_2158,N_3863);
xnor U5001 (N_5001,N_3722,N_3184);
nor U5002 (N_5002,N_3268,N_3064);
nand U5003 (N_5003,N_2234,N_2878);
and U5004 (N_5004,N_3097,N_3285);
nor U5005 (N_5005,N_2915,N_3640);
nor U5006 (N_5006,N_3416,N_3066);
nor U5007 (N_5007,N_2488,N_2939);
and U5008 (N_5008,N_3629,N_2450);
and U5009 (N_5009,N_2254,N_3779);
nand U5010 (N_5010,N_3806,N_3111);
and U5011 (N_5011,N_2799,N_2029);
nor U5012 (N_5012,N_3212,N_3876);
and U5013 (N_5013,N_2408,N_3277);
nand U5014 (N_5014,N_2232,N_3280);
nor U5015 (N_5015,N_2723,N_2293);
and U5016 (N_5016,N_2447,N_3498);
or U5017 (N_5017,N_3372,N_3018);
nand U5018 (N_5018,N_3861,N_3683);
and U5019 (N_5019,N_2407,N_3898);
or U5020 (N_5020,N_3045,N_2498);
or U5021 (N_5021,N_2611,N_3748);
nor U5022 (N_5022,N_2325,N_3704);
or U5023 (N_5023,N_3222,N_3242);
or U5024 (N_5024,N_3748,N_2701);
or U5025 (N_5025,N_3774,N_3601);
nor U5026 (N_5026,N_3595,N_3166);
or U5027 (N_5027,N_2215,N_2713);
nor U5028 (N_5028,N_2066,N_2938);
nor U5029 (N_5029,N_2723,N_3003);
nor U5030 (N_5030,N_3378,N_3801);
nor U5031 (N_5031,N_3771,N_3328);
nor U5032 (N_5032,N_2500,N_2687);
or U5033 (N_5033,N_2486,N_2679);
nor U5034 (N_5034,N_2403,N_3333);
or U5035 (N_5035,N_2438,N_2658);
nor U5036 (N_5036,N_2756,N_3453);
or U5037 (N_5037,N_3756,N_2374);
and U5038 (N_5038,N_2022,N_3322);
nor U5039 (N_5039,N_3042,N_3558);
nor U5040 (N_5040,N_2864,N_2481);
nand U5041 (N_5041,N_2598,N_2493);
nor U5042 (N_5042,N_2350,N_2664);
nand U5043 (N_5043,N_2516,N_3660);
nand U5044 (N_5044,N_2868,N_2863);
nand U5045 (N_5045,N_3498,N_2520);
and U5046 (N_5046,N_3374,N_3963);
and U5047 (N_5047,N_3274,N_3750);
nand U5048 (N_5048,N_3848,N_3171);
nor U5049 (N_5049,N_2761,N_2470);
nand U5050 (N_5050,N_2828,N_2891);
or U5051 (N_5051,N_2660,N_2924);
nor U5052 (N_5052,N_3906,N_2188);
and U5053 (N_5053,N_2874,N_2258);
nand U5054 (N_5054,N_3079,N_3291);
nand U5055 (N_5055,N_2534,N_3102);
nand U5056 (N_5056,N_2374,N_2975);
and U5057 (N_5057,N_2941,N_2545);
and U5058 (N_5058,N_3890,N_2024);
nand U5059 (N_5059,N_2742,N_2050);
and U5060 (N_5060,N_3598,N_3153);
and U5061 (N_5061,N_3959,N_2961);
nand U5062 (N_5062,N_2365,N_3786);
and U5063 (N_5063,N_3615,N_2315);
nand U5064 (N_5064,N_3702,N_3747);
or U5065 (N_5065,N_3200,N_3442);
nand U5066 (N_5066,N_2294,N_3881);
or U5067 (N_5067,N_3679,N_3646);
nor U5068 (N_5068,N_2428,N_2788);
and U5069 (N_5069,N_3511,N_2659);
nand U5070 (N_5070,N_3275,N_3025);
nand U5071 (N_5071,N_3113,N_3262);
nor U5072 (N_5072,N_3105,N_3389);
or U5073 (N_5073,N_2062,N_2548);
or U5074 (N_5074,N_2039,N_2555);
and U5075 (N_5075,N_3165,N_2618);
nand U5076 (N_5076,N_2585,N_3385);
nor U5077 (N_5077,N_2380,N_2227);
nor U5078 (N_5078,N_2380,N_2924);
nor U5079 (N_5079,N_2145,N_2910);
nand U5080 (N_5080,N_3069,N_2456);
nor U5081 (N_5081,N_2667,N_3696);
and U5082 (N_5082,N_3905,N_3120);
or U5083 (N_5083,N_2053,N_2564);
or U5084 (N_5084,N_3778,N_2948);
nand U5085 (N_5085,N_3342,N_2163);
nor U5086 (N_5086,N_2805,N_3518);
and U5087 (N_5087,N_3430,N_2751);
or U5088 (N_5088,N_3162,N_2884);
nand U5089 (N_5089,N_3507,N_3134);
or U5090 (N_5090,N_2207,N_2877);
or U5091 (N_5091,N_3980,N_3675);
nand U5092 (N_5092,N_2601,N_2643);
nand U5093 (N_5093,N_2780,N_2978);
nor U5094 (N_5094,N_2425,N_2828);
nor U5095 (N_5095,N_3244,N_2795);
nor U5096 (N_5096,N_2431,N_3256);
xor U5097 (N_5097,N_2740,N_3704);
nor U5098 (N_5098,N_3965,N_2930);
and U5099 (N_5099,N_3938,N_2453);
nand U5100 (N_5100,N_3981,N_3505);
nand U5101 (N_5101,N_3882,N_3046);
or U5102 (N_5102,N_2617,N_3089);
or U5103 (N_5103,N_2473,N_2656);
or U5104 (N_5104,N_3286,N_2033);
and U5105 (N_5105,N_3132,N_2117);
or U5106 (N_5106,N_3922,N_2231);
nor U5107 (N_5107,N_3226,N_2344);
nand U5108 (N_5108,N_3826,N_2814);
nor U5109 (N_5109,N_3595,N_3308);
nand U5110 (N_5110,N_2731,N_3135);
nand U5111 (N_5111,N_3756,N_3986);
and U5112 (N_5112,N_2632,N_2820);
or U5113 (N_5113,N_3773,N_3170);
nor U5114 (N_5114,N_3301,N_3173);
or U5115 (N_5115,N_3035,N_3988);
nor U5116 (N_5116,N_3074,N_2567);
or U5117 (N_5117,N_2872,N_2208);
or U5118 (N_5118,N_2816,N_2549);
or U5119 (N_5119,N_3888,N_2141);
nand U5120 (N_5120,N_3484,N_2176);
nand U5121 (N_5121,N_3429,N_2467);
nor U5122 (N_5122,N_3871,N_3912);
and U5123 (N_5123,N_3857,N_2756);
or U5124 (N_5124,N_2181,N_2250);
and U5125 (N_5125,N_2794,N_3215);
or U5126 (N_5126,N_2608,N_3195);
nand U5127 (N_5127,N_2080,N_2304);
or U5128 (N_5128,N_2784,N_2262);
nand U5129 (N_5129,N_2338,N_3017);
or U5130 (N_5130,N_3798,N_3228);
or U5131 (N_5131,N_3234,N_3116);
nand U5132 (N_5132,N_2009,N_2374);
nand U5133 (N_5133,N_2237,N_2379);
or U5134 (N_5134,N_2737,N_2375);
and U5135 (N_5135,N_2169,N_3763);
and U5136 (N_5136,N_2734,N_3984);
and U5137 (N_5137,N_3700,N_2332);
nand U5138 (N_5138,N_2245,N_3392);
and U5139 (N_5139,N_2233,N_3801);
or U5140 (N_5140,N_3636,N_2552);
nor U5141 (N_5141,N_3599,N_3572);
nand U5142 (N_5142,N_2646,N_3247);
nand U5143 (N_5143,N_2506,N_3543);
and U5144 (N_5144,N_2313,N_2554);
and U5145 (N_5145,N_3548,N_3377);
nor U5146 (N_5146,N_2033,N_2394);
nand U5147 (N_5147,N_3178,N_2000);
nand U5148 (N_5148,N_2083,N_3053);
nand U5149 (N_5149,N_2900,N_2101);
nor U5150 (N_5150,N_2216,N_2619);
or U5151 (N_5151,N_2214,N_3786);
nor U5152 (N_5152,N_3816,N_2718);
or U5153 (N_5153,N_2328,N_2252);
or U5154 (N_5154,N_2372,N_2819);
or U5155 (N_5155,N_2066,N_3465);
or U5156 (N_5156,N_2886,N_3431);
and U5157 (N_5157,N_2381,N_3807);
or U5158 (N_5158,N_2655,N_2334);
nand U5159 (N_5159,N_2180,N_2250);
nor U5160 (N_5160,N_3529,N_2787);
nand U5161 (N_5161,N_2329,N_2707);
and U5162 (N_5162,N_3819,N_2820);
nor U5163 (N_5163,N_3986,N_3419);
nand U5164 (N_5164,N_2129,N_3240);
and U5165 (N_5165,N_2545,N_3835);
nand U5166 (N_5166,N_2336,N_3571);
or U5167 (N_5167,N_3550,N_2592);
nand U5168 (N_5168,N_2109,N_3584);
and U5169 (N_5169,N_3813,N_3852);
xor U5170 (N_5170,N_2048,N_2000);
and U5171 (N_5171,N_3180,N_3085);
and U5172 (N_5172,N_2983,N_3838);
nor U5173 (N_5173,N_3305,N_3806);
nand U5174 (N_5174,N_2326,N_2302);
or U5175 (N_5175,N_2560,N_2168);
nand U5176 (N_5176,N_3061,N_3158);
or U5177 (N_5177,N_3042,N_3229);
nand U5178 (N_5178,N_3396,N_2873);
or U5179 (N_5179,N_3949,N_2796);
nor U5180 (N_5180,N_3796,N_2431);
nand U5181 (N_5181,N_3161,N_2174);
and U5182 (N_5182,N_2972,N_3671);
nand U5183 (N_5183,N_3844,N_3300);
and U5184 (N_5184,N_2124,N_2301);
and U5185 (N_5185,N_3582,N_3483);
and U5186 (N_5186,N_2196,N_2247);
and U5187 (N_5187,N_2103,N_3237);
nor U5188 (N_5188,N_3174,N_2856);
or U5189 (N_5189,N_2614,N_2275);
or U5190 (N_5190,N_3100,N_2710);
and U5191 (N_5191,N_2073,N_2608);
nor U5192 (N_5192,N_2313,N_2546);
and U5193 (N_5193,N_2375,N_2369);
or U5194 (N_5194,N_3198,N_3165);
nor U5195 (N_5195,N_3822,N_2704);
nand U5196 (N_5196,N_2831,N_3085);
and U5197 (N_5197,N_2852,N_2599);
nand U5198 (N_5198,N_3408,N_2003);
nor U5199 (N_5199,N_3584,N_2655);
nand U5200 (N_5200,N_2243,N_3472);
or U5201 (N_5201,N_2477,N_3528);
or U5202 (N_5202,N_3870,N_3355);
nand U5203 (N_5203,N_2703,N_2232);
nor U5204 (N_5204,N_2427,N_3162);
and U5205 (N_5205,N_3905,N_3101);
and U5206 (N_5206,N_3834,N_2852);
nand U5207 (N_5207,N_2764,N_3963);
nor U5208 (N_5208,N_3557,N_3961);
or U5209 (N_5209,N_3569,N_3658);
nor U5210 (N_5210,N_2864,N_3509);
xnor U5211 (N_5211,N_2906,N_3690);
and U5212 (N_5212,N_2016,N_2536);
and U5213 (N_5213,N_2583,N_3941);
xor U5214 (N_5214,N_2378,N_2046);
and U5215 (N_5215,N_2900,N_2815);
or U5216 (N_5216,N_2410,N_2277);
nor U5217 (N_5217,N_2675,N_2784);
nand U5218 (N_5218,N_3698,N_2584);
nand U5219 (N_5219,N_2599,N_2525);
or U5220 (N_5220,N_2513,N_2652);
nor U5221 (N_5221,N_2406,N_3667);
and U5222 (N_5222,N_2727,N_2368);
and U5223 (N_5223,N_3663,N_2481);
or U5224 (N_5224,N_3395,N_3245);
nor U5225 (N_5225,N_2885,N_2147);
and U5226 (N_5226,N_3127,N_3836);
nor U5227 (N_5227,N_2504,N_3572);
and U5228 (N_5228,N_3695,N_2547);
or U5229 (N_5229,N_3584,N_3337);
and U5230 (N_5230,N_3264,N_2311);
or U5231 (N_5231,N_2023,N_3114);
nor U5232 (N_5232,N_2277,N_2909);
nand U5233 (N_5233,N_3540,N_2532);
or U5234 (N_5234,N_2485,N_2091);
and U5235 (N_5235,N_2076,N_3137);
or U5236 (N_5236,N_2161,N_3794);
and U5237 (N_5237,N_2901,N_2253);
nor U5238 (N_5238,N_2142,N_2872);
nor U5239 (N_5239,N_3006,N_2991);
nor U5240 (N_5240,N_3591,N_2860);
nor U5241 (N_5241,N_2596,N_2984);
nor U5242 (N_5242,N_2088,N_2030);
or U5243 (N_5243,N_2393,N_2936);
or U5244 (N_5244,N_2026,N_3953);
nor U5245 (N_5245,N_2828,N_3271);
or U5246 (N_5246,N_2093,N_2391);
or U5247 (N_5247,N_2215,N_2423);
nand U5248 (N_5248,N_2514,N_3818);
or U5249 (N_5249,N_3540,N_3380);
or U5250 (N_5250,N_3874,N_3553);
or U5251 (N_5251,N_2592,N_3719);
nor U5252 (N_5252,N_2805,N_2942);
or U5253 (N_5253,N_2272,N_3033);
or U5254 (N_5254,N_3530,N_2077);
and U5255 (N_5255,N_3519,N_2369);
nor U5256 (N_5256,N_2610,N_2809);
nor U5257 (N_5257,N_2896,N_3982);
and U5258 (N_5258,N_3319,N_3511);
nand U5259 (N_5259,N_3008,N_3905);
nand U5260 (N_5260,N_2154,N_3765);
nor U5261 (N_5261,N_3574,N_3098);
and U5262 (N_5262,N_3122,N_2047);
and U5263 (N_5263,N_3762,N_2289);
or U5264 (N_5264,N_3691,N_2853);
or U5265 (N_5265,N_3866,N_2193);
and U5266 (N_5266,N_2049,N_2814);
and U5267 (N_5267,N_2754,N_3434);
nor U5268 (N_5268,N_3725,N_2417);
and U5269 (N_5269,N_3009,N_2120);
nor U5270 (N_5270,N_3742,N_3633);
nor U5271 (N_5271,N_2002,N_2800);
nor U5272 (N_5272,N_3673,N_3067);
or U5273 (N_5273,N_2714,N_2827);
nor U5274 (N_5274,N_3096,N_3698);
nor U5275 (N_5275,N_2384,N_3007);
nor U5276 (N_5276,N_3605,N_2836);
nand U5277 (N_5277,N_3579,N_3214);
or U5278 (N_5278,N_3944,N_2854);
nand U5279 (N_5279,N_3087,N_2905);
nor U5280 (N_5280,N_2058,N_2333);
nand U5281 (N_5281,N_3742,N_3805);
nor U5282 (N_5282,N_2807,N_2706);
nand U5283 (N_5283,N_2834,N_2648);
or U5284 (N_5284,N_2888,N_2776);
nor U5285 (N_5285,N_2174,N_3793);
nand U5286 (N_5286,N_3786,N_2439);
or U5287 (N_5287,N_3113,N_2654);
xor U5288 (N_5288,N_3173,N_3401);
nand U5289 (N_5289,N_3627,N_3864);
or U5290 (N_5290,N_3496,N_3531);
or U5291 (N_5291,N_2103,N_2590);
nand U5292 (N_5292,N_2274,N_2919);
or U5293 (N_5293,N_2005,N_3264);
nor U5294 (N_5294,N_2063,N_3758);
nand U5295 (N_5295,N_3660,N_3102);
and U5296 (N_5296,N_3147,N_3629);
or U5297 (N_5297,N_2226,N_2409);
or U5298 (N_5298,N_3991,N_3547);
nand U5299 (N_5299,N_3139,N_3862);
and U5300 (N_5300,N_3488,N_2904);
and U5301 (N_5301,N_2250,N_2488);
and U5302 (N_5302,N_3420,N_3739);
nand U5303 (N_5303,N_2548,N_2956);
and U5304 (N_5304,N_2881,N_2251);
or U5305 (N_5305,N_2988,N_2090);
nand U5306 (N_5306,N_3849,N_2955);
and U5307 (N_5307,N_3262,N_3598);
nand U5308 (N_5308,N_2119,N_2205);
nor U5309 (N_5309,N_2874,N_3762);
nor U5310 (N_5310,N_2127,N_2985);
or U5311 (N_5311,N_3303,N_2629);
and U5312 (N_5312,N_3080,N_3541);
or U5313 (N_5313,N_3891,N_2211);
nand U5314 (N_5314,N_2951,N_3195);
or U5315 (N_5315,N_2187,N_3801);
nor U5316 (N_5316,N_2105,N_2394);
nor U5317 (N_5317,N_3336,N_3440);
and U5318 (N_5318,N_2179,N_3310);
nor U5319 (N_5319,N_3789,N_2209);
nor U5320 (N_5320,N_2209,N_2899);
nor U5321 (N_5321,N_3861,N_2523);
nor U5322 (N_5322,N_2215,N_2669);
xnor U5323 (N_5323,N_3553,N_2297);
nor U5324 (N_5324,N_2637,N_3056);
nor U5325 (N_5325,N_2116,N_2486);
or U5326 (N_5326,N_3869,N_3390);
nand U5327 (N_5327,N_3122,N_2766);
nor U5328 (N_5328,N_3305,N_3720);
or U5329 (N_5329,N_3502,N_3004);
and U5330 (N_5330,N_3644,N_2071);
or U5331 (N_5331,N_2003,N_2757);
and U5332 (N_5332,N_2669,N_2186);
nor U5333 (N_5333,N_3852,N_3935);
or U5334 (N_5334,N_3890,N_3946);
nand U5335 (N_5335,N_2331,N_2645);
nand U5336 (N_5336,N_2871,N_3378);
or U5337 (N_5337,N_2231,N_3148);
nand U5338 (N_5338,N_3554,N_2094);
nor U5339 (N_5339,N_3979,N_2582);
nand U5340 (N_5340,N_3424,N_3957);
and U5341 (N_5341,N_3407,N_3850);
or U5342 (N_5342,N_2209,N_3848);
nand U5343 (N_5343,N_2464,N_3342);
and U5344 (N_5344,N_3772,N_3862);
nand U5345 (N_5345,N_3448,N_2931);
nor U5346 (N_5346,N_3630,N_3109);
or U5347 (N_5347,N_3221,N_2340);
nor U5348 (N_5348,N_3356,N_3207);
nand U5349 (N_5349,N_2516,N_2555);
and U5350 (N_5350,N_3266,N_3714);
nand U5351 (N_5351,N_2598,N_2880);
or U5352 (N_5352,N_2707,N_2725);
nor U5353 (N_5353,N_3254,N_2407);
nand U5354 (N_5354,N_2448,N_3873);
nand U5355 (N_5355,N_2874,N_3087);
and U5356 (N_5356,N_2971,N_3762);
or U5357 (N_5357,N_2428,N_2672);
nand U5358 (N_5358,N_3824,N_2251);
or U5359 (N_5359,N_2817,N_3201);
nor U5360 (N_5360,N_3699,N_3829);
nand U5361 (N_5361,N_3253,N_3751);
or U5362 (N_5362,N_2377,N_2246);
nand U5363 (N_5363,N_3641,N_3505);
nor U5364 (N_5364,N_2511,N_3652);
or U5365 (N_5365,N_3098,N_2013);
nor U5366 (N_5366,N_2608,N_2296);
nand U5367 (N_5367,N_3952,N_2880);
nand U5368 (N_5368,N_3873,N_3744);
and U5369 (N_5369,N_3169,N_2703);
or U5370 (N_5370,N_2846,N_3444);
or U5371 (N_5371,N_3302,N_3929);
nand U5372 (N_5372,N_3685,N_3587);
nand U5373 (N_5373,N_2912,N_3881);
nand U5374 (N_5374,N_3697,N_3589);
and U5375 (N_5375,N_2372,N_3653);
and U5376 (N_5376,N_3653,N_3271);
nand U5377 (N_5377,N_3473,N_3806);
or U5378 (N_5378,N_3769,N_3536);
nor U5379 (N_5379,N_3363,N_3254);
nor U5380 (N_5380,N_2754,N_2684);
or U5381 (N_5381,N_2962,N_3124);
nor U5382 (N_5382,N_3002,N_3872);
nor U5383 (N_5383,N_3875,N_3459);
nand U5384 (N_5384,N_2235,N_3757);
and U5385 (N_5385,N_3425,N_3853);
nand U5386 (N_5386,N_2144,N_2030);
or U5387 (N_5387,N_2152,N_3377);
or U5388 (N_5388,N_3837,N_3425);
and U5389 (N_5389,N_3604,N_3671);
and U5390 (N_5390,N_2783,N_2512);
or U5391 (N_5391,N_3533,N_3710);
nand U5392 (N_5392,N_2754,N_3062);
nand U5393 (N_5393,N_3152,N_3371);
and U5394 (N_5394,N_3988,N_3716);
nand U5395 (N_5395,N_2335,N_2705);
xor U5396 (N_5396,N_2096,N_3406);
nor U5397 (N_5397,N_3025,N_2063);
and U5398 (N_5398,N_2247,N_2118);
and U5399 (N_5399,N_2801,N_2488);
or U5400 (N_5400,N_2245,N_3525);
nand U5401 (N_5401,N_3622,N_2612);
or U5402 (N_5402,N_3930,N_3558);
nand U5403 (N_5403,N_3406,N_2806);
nand U5404 (N_5404,N_3033,N_3737);
and U5405 (N_5405,N_2265,N_3098);
nor U5406 (N_5406,N_2893,N_3470);
or U5407 (N_5407,N_3719,N_2612);
and U5408 (N_5408,N_2266,N_2935);
nand U5409 (N_5409,N_3942,N_2609);
or U5410 (N_5410,N_3764,N_3521);
nor U5411 (N_5411,N_2505,N_2493);
or U5412 (N_5412,N_2941,N_2243);
and U5413 (N_5413,N_3081,N_3880);
or U5414 (N_5414,N_2123,N_2611);
or U5415 (N_5415,N_2820,N_3464);
or U5416 (N_5416,N_2004,N_3196);
nor U5417 (N_5417,N_2653,N_3480);
and U5418 (N_5418,N_2193,N_2889);
nand U5419 (N_5419,N_3498,N_2950);
and U5420 (N_5420,N_2146,N_2521);
nand U5421 (N_5421,N_3868,N_3888);
nor U5422 (N_5422,N_3735,N_3682);
nor U5423 (N_5423,N_2527,N_3132);
and U5424 (N_5424,N_3972,N_2957);
nor U5425 (N_5425,N_3925,N_2380);
or U5426 (N_5426,N_2730,N_2980);
nand U5427 (N_5427,N_3906,N_3064);
and U5428 (N_5428,N_2557,N_3458);
nand U5429 (N_5429,N_3441,N_2037);
and U5430 (N_5430,N_3836,N_2297);
and U5431 (N_5431,N_3909,N_3429);
nor U5432 (N_5432,N_3151,N_2906);
or U5433 (N_5433,N_3826,N_3888);
or U5434 (N_5434,N_3388,N_2580);
and U5435 (N_5435,N_3076,N_2950);
nor U5436 (N_5436,N_2961,N_3028);
or U5437 (N_5437,N_2045,N_3706);
nand U5438 (N_5438,N_3123,N_3512);
nand U5439 (N_5439,N_2800,N_2738);
nand U5440 (N_5440,N_2684,N_3883);
or U5441 (N_5441,N_3497,N_3523);
or U5442 (N_5442,N_2948,N_2709);
or U5443 (N_5443,N_3543,N_3615);
nor U5444 (N_5444,N_2855,N_3221);
and U5445 (N_5445,N_3782,N_3518);
nand U5446 (N_5446,N_2544,N_3219);
nand U5447 (N_5447,N_2753,N_3595);
nor U5448 (N_5448,N_2997,N_2180);
or U5449 (N_5449,N_3529,N_3843);
or U5450 (N_5450,N_2637,N_3637);
nor U5451 (N_5451,N_3483,N_2199);
and U5452 (N_5452,N_2383,N_3062);
or U5453 (N_5453,N_2454,N_2748);
nand U5454 (N_5454,N_2028,N_2844);
nand U5455 (N_5455,N_3467,N_2272);
or U5456 (N_5456,N_2978,N_3034);
nor U5457 (N_5457,N_3155,N_2412);
nor U5458 (N_5458,N_2029,N_2952);
nand U5459 (N_5459,N_2290,N_2232);
or U5460 (N_5460,N_3621,N_2589);
nand U5461 (N_5461,N_2273,N_2000);
and U5462 (N_5462,N_3433,N_3297);
and U5463 (N_5463,N_2412,N_2921);
nand U5464 (N_5464,N_3561,N_2368);
and U5465 (N_5465,N_2128,N_3749);
nand U5466 (N_5466,N_3982,N_3529);
and U5467 (N_5467,N_3831,N_2959);
or U5468 (N_5468,N_3883,N_3859);
and U5469 (N_5469,N_3746,N_3593);
or U5470 (N_5470,N_3967,N_2913);
or U5471 (N_5471,N_3046,N_2219);
or U5472 (N_5472,N_3859,N_2806);
nor U5473 (N_5473,N_2068,N_3206);
nand U5474 (N_5474,N_2919,N_2618);
and U5475 (N_5475,N_3450,N_3590);
nand U5476 (N_5476,N_3397,N_2931);
or U5477 (N_5477,N_3851,N_3911);
and U5478 (N_5478,N_2289,N_3248);
nor U5479 (N_5479,N_2984,N_2942);
nor U5480 (N_5480,N_2951,N_2798);
nand U5481 (N_5481,N_2026,N_2267);
and U5482 (N_5482,N_2474,N_3329);
and U5483 (N_5483,N_2197,N_3161);
and U5484 (N_5484,N_3287,N_2541);
nand U5485 (N_5485,N_3308,N_2000);
or U5486 (N_5486,N_2032,N_3849);
nand U5487 (N_5487,N_2300,N_3285);
or U5488 (N_5488,N_2205,N_2384);
or U5489 (N_5489,N_2403,N_2321);
and U5490 (N_5490,N_2074,N_2140);
nor U5491 (N_5491,N_2623,N_3420);
nand U5492 (N_5492,N_2207,N_3530);
or U5493 (N_5493,N_2531,N_2927);
or U5494 (N_5494,N_3900,N_2951);
nor U5495 (N_5495,N_2404,N_2050);
nor U5496 (N_5496,N_2175,N_2482);
and U5497 (N_5497,N_3574,N_3556);
or U5498 (N_5498,N_3330,N_2529);
and U5499 (N_5499,N_3084,N_2964);
and U5500 (N_5500,N_2883,N_2814);
nor U5501 (N_5501,N_2976,N_3983);
nand U5502 (N_5502,N_3825,N_2677);
and U5503 (N_5503,N_3455,N_2443);
nand U5504 (N_5504,N_2812,N_2434);
or U5505 (N_5505,N_3331,N_3775);
or U5506 (N_5506,N_2841,N_2755);
nand U5507 (N_5507,N_3339,N_2840);
or U5508 (N_5508,N_3830,N_2061);
nor U5509 (N_5509,N_3237,N_3498);
and U5510 (N_5510,N_3181,N_2641);
nor U5511 (N_5511,N_3975,N_3608);
nor U5512 (N_5512,N_2976,N_3344);
nand U5513 (N_5513,N_3384,N_2070);
nand U5514 (N_5514,N_2652,N_3421);
nor U5515 (N_5515,N_2118,N_2236);
or U5516 (N_5516,N_2945,N_2689);
or U5517 (N_5517,N_2755,N_3793);
nand U5518 (N_5518,N_2266,N_2657);
nor U5519 (N_5519,N_2748,N_2177);
nand U5520 (N_5520,N_3465,N_2926);
or U5521 (N_5521,N_3567,N_3252);
and U5522 (N_5522,N_2779,N_2814);
or U5523 (N_5523,N_2517,N_2001);
nor U5524 (N_5524,N_2785,N_3020);
or U5525 (N_5525,N_2736,N_3402);
or U5526 (N_5526,N_2586,N_3207);
or U5527 (N_5527,N_2683,N_2459);
nand U5528 (N_5528,N_3837,N_3016);
or U5529 (N_5529,N_3737,N_3073);
nor U5530 (N_5530,N_3227,N_2594);
and U5531 (N_5531,N_3541,N_3969);
and U5532 (N_5532,N_3316,N_3489);
nor U5533 (N_5533,N_2383,N_3816);
or U5534 (N_5534,N_3841,N_3360);
nand U5535 (N_5535,N_2982,N_3487);
and U5536 (N_5536,N_3406,N_3947);
and U5537 (N_5537,N_2423,N_3112);
and U5538 (N_5538,N_2944,N_3039);
or U5539 (N_5539,N_3952,N_3668);
or U5540 (N_5540,N_3019,N_2872);
or U5541 (N_5541,N_2064,N_2136);
nand U5542 (N_5542,N_3220,N_3376);
or U5543 (N_5543,N_2904,N_3876);
or U5544 (N_5544,N_3438,N_2446);
or U5545 (N_5545,N_3690,N_3570);
nand U5546 (N_5546,N_3797,N_2422);
or U5547 (N_5547,N_3146,N_3164);
and U5548 (N_5548,N_3839,N_2002);
nor U5549 (N_5549,N_3944,N_2690);
nand U5550 (N_5550,N_2497,N_3305);
or U5551 (N_5551,N_3960,N_3518);
or U5552 (N_5552,N_3475,N_3028);
nand U5553 (N_5553,N_2414,N_3587);
and U5554 (N_5554,N_2258,N_3767);
or U5555 (N_5555,N_3619,N_2169);
or U5556 (N_5556,N_2854,N_2882);
nand U5557 (N_5557,N_3862,N_3070);
nor U5558 (N_5558,N_3207,N_3518);
nor U5559 (N_5559,N_3785,N_3430);
and U5560 (N_5560,N_2154,N_3239);
or U5561 (N_5561,N_2663,N_3727);
nor U5562 (N_5562,N_2557,N_3237);
nand U5563 (N_5563,N_3719,N_3997);
nand U5564 (N_5564,N_2398,N_2737);
and U5565 (N_5565,N_2335,N_2200);
nand U5566 (N_5566,N_2400,N_3597);
and U5567 (N_5567,N_2440,N_2427);
nand U5568 (N_5568,N_3039,N_2835);
and U5569 (N_5569,N_3631,N_2942);
or U5570 (N_5570,N_2393,N_2823);
nor U5571 (N_5571,N_2602,N_2986);
or U5572 (N_5572,N_2105,N_3699);
or U5573 (N_5573,N_2111,N_3510);
nand U5574 (N_5574,N_2283,N_2046);
nand U5575 (N_5575,N_3327,N_2687);
and U5576 (N_5576,N_2697,N_2957);
nor U5577 (N_5577,N_3066,N_2581);
and U5578 (N_5578,N_2733,N_2110);
nor U5579 (N_5579,N_3053,N_3317);
nor U5580 (N_5580,N_2803,N_3957);
nor U5581 (N_5581,N_2860,N_3991);
nand U5582 (N_5582,N_3818,N_3088);
and U5583 (N_5583,N_3934,N_3224);
nand U5584 (N_5584,N_2712,N_2629);
nor U5585 (N_5585,N_2841,N_3053);
nand U5586 (N_5586,N_3824,N_2412);
nand U5587 (N_5587,N_3216,N_2746);
or U5588 (N_5588,N_3352,N_3865);
and U5589 (N_5589,N_2851,N_3017);
and U5590 (N_5590,N_3977,N_2944);
nand U5591 (N_5591,N_3635,N_2500);
nor U5592 (N_5592,N_3192,N_3891);
nor U5593 (N_5593,N_2920,N_2038);
or U5594 (N_5594,N_2496,N_3455);
and U5595 (N_5595,N_3417,N_2672);
and U5596 (N_5596,N_2480,N_3760);
and U5597 (N_5597,N_3006,N_2474);
or U5598 (N_5598,N_3963,N_2883);
or U5599 (N_5599,N_2175,N_2854);
and U5600 (N_5600,N_2385,N_3851);
or U5601 (N_5601,N_3443,N_3676);
nand U5602 (N_5602,N_2072,N_2355);
or U5603 (N_5603,N_2986,N_3849);
and U5604 (N_5604,N_2523,N_3433);
nand U5605 (N_5605,N_2814,N_3859);
and U5606 (N_5606,N_2319,N_2069);
and U5607 (N_5607,N_3605,N_2415);
or U5608 (N_5608,N_2479,N_3413);
nor U5609 (N_5609,N_2937,N_2720);
or U5610 (N_5610,N_3964,N_3742);
nand U5611 (N_5611,N_2898,N_2774);
nor U5612 (N_5612,N_3950,N_2509);
nand U5613 (N_5613,N_3477,N_2744);
nand U5614 (N_5614,N_2830,N_2734);
nand U5615 (N_5615,N_2548,N_3236);
or U5616 (N_5616,N_3814,N_2442);
and U5617 (N_5617,N_3433,N_3861);
xor U5618 (N_5618,N_2785,N_2683);
xnor U5619 (N_5619,N_3989,N_3378);
nand U5620 (N_5620,N_2761,N_2244);
nor U5621 (N_5621,N_2891,N_2372);
nor U5622 (N_5622,N_2399,N_2863);
nor U5623 (N_5623,N_2077,N_3046);
or U5624 (N_5624,N_3609,N_2098);
or U5625 (N_5625,N_3189,N_2993);
or U5626 (N_5626,N_3571,N_2958);
and U5627 (N_5627,N_2660,N_2005);
and U5628 (N_5628,N_3034,N_3479);
nor U5629 (N_5629,N_2660,N_2975);
nor U5630 (N_5630,N_3676,N_3501);
nand U5631 (N_5631,N_2392,N_3540);
and U5632 (N_5632,N_3844,N_3825);
nand U5633 (N_5633,N_3723,N_2187);
or U5634 (N_5634,N_2361,N_3353);
or U5635 (N_5635,N_3408,N_2694);
nor U5636 (N_5636,N_3356,N_2490);
or U5637 (N_5637,N_3608,N_3798);
or U5638 (N_5638,N_2066,N_2367);
nand U5639 (N_5639,N_2028,N_3157);
nand U5640 (N_5640,N_3710,N_2260);
nand U5641 (N_5641,N_3269,N_2210);
nor U5642 (N_5642,N_2901,N_3296);
and U5643 (N_5643,N_3549,N_3469);
or U5644 (N_5644,N_2515,N_2284);
nor U5645 (N_5645,N_2746,N_3587);
and U5646 (N_5646,N_3215,N_2293);
nand U5647 (N_5647,N_2825,N_3768);
nor U5648 (N_5648,N_3188,N_3859);
nand U5649 (N_5649,N_2051,N_2302);
nand U5650 (N_5650,N_3114,N_3702);
nor U5651 (N_5651,N_3638,N_3334);
nand U5652 (N_5652,N_2209,N_2506);
and U5653 (N_5653,N_3777,N_2458);
or U5654 (N_5654,N_3518,N_2641);
nand U5655 (N_5655,N_2156,N_3091);
and U5656 (N_5656,N_3408,N_3554);
and U5657 (N_5657,N_3596,N_2935);
nor U5658 (N_5658,N_3151,N_2249);
and U5659 (N_5659,N_3079,N_2221);
nor U5660 (N_5660,N_2479,N_3313);
and U5661 (N_5661,N_3371,N_3433);
or U5662 (N_5662,N_2398,N_2913);
nor U5663 (N_5663,N_2441,N_2958);
or U5664 (N_5664,N_3068,N_3163);
nor U5665 (N_5665,N_2282,N_3197);
or U5666 (N_5666,N_3316,N_3166);
and U5667 (N_5667,N_2458,N_2991);
nor U5668 (N_5668,N_3386,N_2866);
and U5669 (N_5669,N_2386,N_3806);
or U5670 (N_5670,N_3317,N_3208);
nand U5671 (N_5671,N_3359,N_3806);
or U5672 (N_5672,N_2995,N_2112);
and U5673 (N_5673,N_3377,N_3700);
nor U5674 (N_5674,N_3415,N_2417);
or U5675 (N_5675,N_3284,N_3247);
or U5676 (N_5676,N_3407,N_2107);
and U5677 (N_5677,N_3691,N_2508);
xnor U5678 (N_5678,N_3696,N_3849);
nor U5679 (N_5679,N_3339,N_3437);
and U5680 (N_5680,N_2622,N_2222);
or U5681 (N_5681,N_3225,N_2858);
and U5682 (N_5682,N_2150,N_3123);
or U5683 (N_5683,N_2512,N_3108);
nor U5684 (N_5684,N_2921,N_3011);
nand U5685 (N_5685,N_3301,N_2168);
nand U5686 (N_5686,N_2473,N_2661);
nor U5687 (N_5687,N_3413,N_3940);
or U5688 (N_5688,N_2084,N_3637);
nor U5689 (N_5689,N_2974,N_3275);
or U5690 (N_5690,N_3313,N_3822);
or U5691 (N_5691,N_2879,N_3526);
and U5692 (N_5692,N_3780,N_2615);
or U5693 (N_5693,N_2929,N_2023);
nand U5694 (N_5694,N_3666,N_2207);
nor U5695 (N_5695,N_2489,N_3438);
nor U5696 (N_5696,N_3375,N_3905);
and U5697 (N_5697,N_2435,N_2794);
or U5698 (N_5698,N_3335,N_3358);
nand U5699 (N_5699,N_3707,N_3581);
or U5700 (N_5700,N_2905,N_3308);
nor U5701 (N_5701,N_3093,N_2672);
or U5702 (N_5702,N_3164,N_3624);
nor U5703 (N_5703,N_2327,N_3755);
nor U5704 (N_5704,N_3478,N_3543);
nand U5705 (N_5705,N_3904,N_3315);
or U5706 (N_5706,N_3835,N_3308);
nor U5707 (N_5707,N_2762,N_2366);
or U5708 (N_5708,N_3260,N_3201);
or U5709 (N_5709,N_2115,N_2761);
nor U5710 (N_5710,N_3707,N_2005);
or U5711 (N_5711,N_3464,N_2161);
nand U5712 (N_5712,N_3429,N_2220);
nand U5713 (N_5713,N_2621,N_2931);
nand U5714 (N_5714,N_2090,N_3442);
nor U5715 (N_5715,N_3969,N_2145);
nor U5716 (N_5716,N_2355,N_3241);
or U5717 (N_5717,N_3288,N_2827);
or U5718 (N_5718,N_2544,N_2521);
nor U5719 (N_5719,N_2428,N_3286);
nor U5720 (N_5720,N_3366,N_3287);
nand U5721 (N_5721,N_3396,N_3358);
or U5722 (N_5722,N_3894,N_2180);
or U5723 (N_5723,N_2523,N_3667);
or U5724 (N_5724,N_3651,N_3167);
and U5725 (N_5725,N_2823,N_2349);
nand U5726 (N_5726,N_3205,N_2615);
xor U5727 (N_5727,N_3224,N_2587);
nor U5728 (N_5728,N_2498,N_2149);
and U5729 (N_5729,N_3738,N_2690);
and U5730 (N_5730,N_2822,N_2289);
or U5731 (N_5731,N_3114,N_2958);
and U5732 (N_5732,N_2320,N_2922);
nor U5733 (N_5733,N_2806,N_2625);
or U5734 (N_5734,N_3389,N_3589);
or U5735 (N_5735,N_3702,N_2517);
or U5736 (N_5736,N_2926,N_2768);
nor U5737 (N_5737,N_2214,N_2973);
and U5738 (N_5738,N_2408,N_3071);
or U5739 (N_5739,N_2161,N_2727);
nor U5740 (N_5740,N_3102,N_3427);
nor U5741 (N_5741,N_2583,N_2789);
or U5742 (N_5742,N_2561,N_2049);
and U5743 (N_5743,N_3695,N_2765);
and U5744 (N_5744,N_3904,N_2463);
and U5745 (N_5745,N_3522,N_2438);
nand U5746 (N_5746,N_3667,N_2241);
and U5747 (N_5747,N_2281,N_3711);
or U5748 (N_5748,N_2317,N_2905);
nor U5749 (N_5749,N_2232,N_2866);
and U5750 (N_5750,N_2519,N_2129);
nor U5751 (N_5751,N_3490,N_3445);
nor U5752 (N_5752,N_2302,N_2220);
and U5753 (N_5753,N_3922,N_2238);
nor U5754 (N_5754,N_3461,N_2613);
or U5755 (N_5755,N_3229,N_3792);
nand U5756 (N_5756,N_3252,N_2670);
and U5757 (N_5757,N_3603,N_3103);
nand U5758 (N_5758,N_3143,N_2125);
and U5759 (N_5759,N_3590,N_3407);
nand U5760 (N_5760,N_2903,N_3583);
or U5761 (N_5761,N_2474,N_2079);
and U5762 (N_5762,N_2058,N_3281);
nand U5763 (N_5763,N_2830,N_3698);
and U5764 (N_5764,N_3308,N_3284);
nand U5765 (N_5765,N_2940,N_3136);
or U5766 (N_5766,N_2578,N_3897);
nand U5767 (N_5767,N_2939,N_2044);
and U5768 (N_5768,N_2484,N_3079);
and U5769 (N_5769,N_2061,N_2724);
nand U5770 (N_5770,N_3801,N_2956);
nand U5771 (N_5771,N_3316,N_3767);
or U5772 (N_5772,N_3722,N_3897);
and U5773 (N_5773,N_3387,N_3871);
and U5774 (N_5774,N_2354,N_3549);
nand U5775 (N_5775,N_3554,N_2664);
xor U5776 (N_5776,N_3891,N_2262);
nand U5777 (N_5777,N_2886,N_3856);
or U5778 (N_5778,N_2103,N_2798);
nand U5779 (N_5779,N_3166,N_3593);
nor U5780 (N_5780,N_3989,N_2966);
and U5781 (N_5781,N_3232,N_3524);
nand U5782 (N_5782,N_3265,N_2116);
or U5783 (N_5783,N_2541,N_3576);
or U5784 (N_5784,N_2233,N_2373);
or U5785 (N_5785,N_3265,N_2888);
or U5786 (N_5786,N_2824,N_2288);
or U5787 (N_5787,N_3683,N_2473);
and U5788 (N_5788,N_3218,N_2262);
nand U5789 (N_5789,N_2174,N_3812);
or U5790 (N_5790,N_2643,N_3349);
and U5791 (N_5791,N_2402,N_2521);
and U5792 (N_5792,N_3572,N_2238);
or U5793 (N_5793,N_2248,N_3805);
nand U5794 (N_5794,N_2509,N_3754);
nor U5795 (N_5795,N_2301,N_2542);
nor U5796 (N_5796,N_2273,N_2539);
nand U5797 (N_5797,N_3353,N_2072);
or U5798 (N_5798,N_3593,N_2877);
and U5799 (N_5799,N_3696,N_3787);
or U5800 (N_5800,N_3257,N_3915);
or U5801 (N_5801,N_2104,N_2911);
xnor U5802 (N_5802,N_2730,N_3141);
nand U5803 (N_5803,N_2462,N_2180);
or U5804 (N_5804,N_2339,N_2320);
nor U5805 (N_5805,N_2113,N_3772);
nand U5806 (N_5806,N_3278,N_2256);
or U5807 (N_5807,N_2442,N_2662);
or U5808 (N_5808,N_2889,N_3441);
nand U5809 (N_5809,N_3412,N_2130);
nand U5810 (N_5810,N_3813,N_3150);
nor U5811 (N_5811,N_3070,N_3677);
nor U5812 (N_5812,N_2957,N_3038);
or U5813 (N_5813,N_3508,N_3303);
nand U5814 (N_5814,N_3901,N_3313);
nor U5815 (N_5815,N_3000,N_3838);
nand U5816 (N_5816,N_3185,N_3032);
nor U5817 (N_5817,N_3670,N_2410);
nor U5818 (N_5818,N_3046,N_2440);
or U5819 (N_5819,N_2408,N_2841);
and U5820 (N_5820,N_3135,N_2212);
nor U5821 (N_5821,N_2297,N_3120);
nor U5822 (N_5822,N_3094,N_2098);
xor U5823 (N_5823,N_3334,N_3461);
nor U5824 (N_5824,N_3539,N_3951);
nor U5825 (N_5825,N_3998,N_2025);
or U5826 (N_5826,N_3301,N_2011);
or U5827 (N_5827,N_3759,N_3017);
nand U5828 (N_5828,N_3427,N_3238);
nand U5829 (N_5829,N_2100,N_3533);
or U5830 (N_5830,N_2510,N_3851);
nand U5831 (N_5831,N_2697,N_2349);
nor U5832 (N_5832,N_3399,N_3822);
and U5833 (N_5833,N_3374,N_2585);
or U5834 (N_5834,N_3547,N_2086);
nor U5835 (N_5835,N_2530,N_3602);
nand U5836 (N_5836,N_2569,N_2490);
nand U5837 (N_5837,N_3381,N_2177);
and U5838 (N_5838,N_2317,N_2185);
and U5839 (N_5839,N_2723,N_3031);
nand U5840 (N_5840,N_2057,N_3558);
and U5841 (N_5841,N_2908,N_2681);
nor U5842 (N_5842,N_2091,N_2941);
and U5843 (N_5843,N_3824,N_3538);
or U5844 (N_5844,N_2207,N_2034);
and U5845 (N_5845,N_2253,N_2147);
nand U5846 (N_5846,N_3298,N_3613);
and U5847 (N_5847,N_3517,N_2955);
or U5848 (N_5848,N_3221,N_2104);
nor U5849 (N_5849,N_3402,N_2929);
nor U5850 (N_5850,N_3081,N_3067);
nor U5851 (N_5851,N_2549,N_3128);
or U5852 (N_5852,N_3186,N_2798);
and U5853 (N_5853,N_2024,N_2025);
nor U5854 (N_5854,N_2242,N_3036);
nand U5855 (N_5855,N_2284,N_3702);
xnor U5856 (N_5856,N_2416,N_2123);
or U5857 (N_5857,N_2260,N_3809);
nor U5858 (N_5858,N_2892,N_3119);
nor U5859 (N_5859,N_3706,N_2381);
and U5860 (N_5860,N_2164,N_2380);
nand U5861 (N_5861,N_2538,N_2063);
and U5862 (N_5862,N_3841,N_3837);
and U5863 (N_5863,N_3911,N_2658);
nor U5864 (N_5864,N_2231,N_2166);
nor U5865 (N_5865,N_3490,N_3321);
nand U5866 (N_5866,N_2146,N_3090);
nor U5867 (N_5867,N_3641,N_2064);
and U5868 (N_5868,N_3487,N_3591);
nand U5869 (N_5869,N_3802,N_2980);
nor U5870 (N_5870,N_3458,N_2453);
or U5871 (N_5871,N_2823,N_3531);
nor U5872 (N_5872,N_3916,N_2540);
or U5873 (N_5873,N_2132,N_2681);
and U5874 (N_5874,N_2712,N_2525);
and U5875 (N_5875,N_2406,N_2716);
or U5876 (N_5876,N_2669,N_3364);
nor U5877 (N_5877,N_2240,N_3772);
nand U5878 (N_5878,N_2463,N_2438);
nor U5879 (N_5879,N_3777,N_3710);
nor U5880 (N_5880,N_2623,N_3319);
and U5881 (N_5881,N_2356,N_3082);
and U5882 (N_5882,N_2934,N_3303);
or U5883 (N_5883,N_2849,N_2641);
or U5884 (N_5884,N_2685,N_2575);
or U5885 (N_5885,N_2015,N_3606);
nor U5886 (N_5886,N_2327,N_2939);
nor U5887 (N_5887,N_2050,N_2426);
or U5888 (N_5888,N_2378,N_3853);
and U5889 (N_5889,N_3951,N_3976);
nand U5890 (N_5890,N_3552,N_2984);
and U5891 (N_5891,N_3749,N_3064);
nand U5892 (N_5892,N_3660,N_2470);
or U5893 (N_5893,N_3918,N_2925);
nand U5894 (N_5894,N_3935,N_3807);
nor U5895 (N_5895,N_3349,N_2458);
nor U5896 (N_5896,N_3944,N_3207);
nor U5897 (N_5897,N_3682,N_3394);
and U5898 (N_5898,N_3198,N_2641);
nor U5899 (N_5899,N_2962,N_2208);
nand U5900 (N_5900,N_3923,N_2313);
or U5901 (N_5901,N_2145,N_3578);
nand U5902 (N_5902,N_3246,N_2332);
or U5903 (N_5903,N_2489,N_3399);
and U5904 (N_5904,N_2714,N_3816);
nand U5905 (N_5905,N_3896,N_3543);
or U5906 (N_5906,N_3121,N_2737);
nor U5907 (N_5907,N_3869,N_2118);
nor U5908 (N_5908,N_3181,N_3221);
or U5909 (N_5909,N_2412,N_3436);
or U5910 (N_5910,N_2223,N_2661);
and U5911 (N_5911,N_3790,N_3319);
and U5912 (N_5912,N_3302,N_2040);
nand U5913 (N_5913,N_2909,N_3523);
or U5914 (N_5914,N_2946,N_3997);
or U5915 (N_5915,N_3740,N_2549);
or U5916 (N_5916,N_2875,N_2136);
or U5917 (N_5917,N_3083,N_2411);
nand U5918 (N_5918,N_3216,N_2942);
or U5919 (N_5919,N_2529,N_3670);
nand U5920 (N_5920,N_2541,N_3053);
nand U5921 (N_5921,N_2414,N_3011);
or U5922 (N_5922,N_3491,N_3958);
and U5923 (N_5923,N_2928,N_3926);
nor U5924 (N_5924,N_3565,N_2222);
and U5925 (N_5925,N_3602,N_3550);
nand U5926 (N_5926,N_3571,N_3838);
nor U5927 (N_5927,N_2743,N_3534);
nor U5928 (N_5928,N_2570,N_3691);
nor U5929 (N_5929,N_3401,N_2218);
nand U5930 (N_5930,N_2381,N_2443);
nor U5931 (N_5931,N_2221,N_2669);
nand U5932 (N_5932,N_3149,N_3838);
nor U5933 (N_5933,N_3693,N_2054);
nand U5934 (N_5934,N_2924,N_3207);
nand U5935 (N_5935,N_3849,N_2210);
and U5936 (N_5936,N_2207,N_3000);
nor U5937 (N_5937,N_3962,N_2309);
nand U5938 (N_5938,N_2570,N_3780);
and U5939 (N_5939,N_2199,N_3482);
and U5940 (N_5940,N_3407,N_3715);
or U5941 (N_5941,N_3597,N_2123);
nor U5942 (N_5942,N_3221,N_3423);
or U5943 (N_5943,N_2557,N_2234);
or U5944 (N_5944,N_3023,N_3928);
nor U5945 (N_5945,N_3172,N_3110);
and U5946 (N_5946,N_3637,N_3425);
and U5947 (N_5947,N_3107,N_3175);
nand U5948 (N_5948,N_3729,N_2328);
and U5949 (N_5949,N_3107,N_2997);
or U5950 (N_5950,N_3662,N_3422);
and U5951 (N_5951,N_2199,N_2033);
nor U5952 (N_5952,N_3078,N_2615);
or U5953 (N_5953,N_3527,N_2582);
and U5954 (N_5954,N_3114,N_3773);
and U5955 (N_5955,N_3448,N_2596);
nor U5956 (N_5956,N_3335,N_3339);
and U5957 (N_5957,N_2510,N_3256);
or U5958 (N_5958,N_3919,N_3796);
and U5959 (N_5959,N_3991,N_2292);
nor U5960 (N_5960,N_2620,N_3885);
or U5961 (N_5961,N_2151,N_2912);
nor U5962 (N_5962,N_2552,N_2985);
and U5963 (N_5963,N_2764,N_3665);
and U5964 (N_5964,N_3157,N_3230);
and U5965 (N_5965,N_2260,N_3571);
or U5966 (N_5966,N_3670,N_3460);
nand U5967 (N_5967,N_2719,N_2863);
and U5968 (N_5968,N_2777,N_3582);
nand U5969 (N_5969,N_2746,N_2296);
nor U5970 (N_5970,N_2267,N_2331);
nor U5971 (N_5971,N_2504,N_2420);
nor U5972 (N_5972,N_2905,N_2906);
nor U5973 (N_5973,N_3392,N_3571);
nand U5974 (N_5974,N_2853,N_2121);
nor U5975 (N_5975,N_3307,N_2450);
or U5976 (N_5976,N_3520,N_2655);
nor U5977 (N_5977,N_2681,N_2314);
or U5978 (N_5978,N_3542,N_3136);
nor U5979 (N_5979,N_3147,N_3644);
or U5980 (N_5980,N_2879,N_3549);
nand U5981 (N_5981,N_2052,N_2227);
and U5982 (N_5982,N_3884,N_2847);
and U5983 (N_5983,N_2109,N_2622);
nand U5984 (N_5984,N_2282,N_3079);
nor U5985 (N_5985,N_3807,N_2544);
nor U5986 (N_5986,N_3406,N_3597);
or U5987 (N_5987,N_2041,N_2485);
or U5988 (N_5988,N_3951,N_2036);
or U5989 (N_5989,N_3465,N_3102);
or U5990 (N_5990,N_3601,N_2454);
nor U5991 (N_5991,N_2557,N_2475);
nand U5992 (N_5992,N_2216,N_2591);
nor U5993 (N_5993,N_3884,N_3724);
and U5994 (N_5994,N_3077,N_2778);
nor U5995 (N_5995,N_2127,N_3146);
or U5996 (N_5996,N_3969,N_3058);
and U5997 (N_5997,N_2382,N_3888);
nor U5998 (N_5998,N_3146,N_2913);
and U5999 (N_5999,N_2417,N_3083);
and U6000 (N_6000,N_4292,N_5648);
or U6001 (N_6001,N_4969,N_5313);
nand U6002 (N_6002,N_4789,N_4771);
nand U6003 (N_6003,N_5651,N_4516);
nor U6004 (N_6004,N_5245,N_5251);
nand U6005 (N_6005,N_5471,N_4370);
nor U6006 (N_6006,N_4564,N_4556);
nor U6007 (N_6007,N_5608,N_5791);
and U6008 (N_6008,N_5224,N_4888);
nand U6009 (N_6009,N_5529,N_5719);
and U6010 (N_6010,N_4599,N_4884);
nand U6011 (N_6011,N_4245,N_5149);
nand U6012 (N_6012,N_4592,N_4151);
and U6013 (N_6013,N_5188,N_5318);
nand U6014 (N_6014,N_5894,N_4800);
and U6015 (N_6015,N_5602,N_5732);
or U6016 (N_6016,N_5514,N_4179);
or U6017 (N_6017,N_5959,N_5876);
nor U6018 (N_6018,N_4666,N_5053);
and U6019 (N_6019,N_5988,N_5438);
or U6020 (N_6020,N_5232,N_5717);
or U6021 (N_6021,N_4461,N_5343);
or U6022 (N_6022,N_5002,N_5384);
and U6023 (N_6023,N_4918,N_4723);
and U6024 (N_6024,N_4540,N_4144);
nand U6025 (N_6025,N_5410,N_4428);
or U6026 (N_6026,N_5526,N_4215);
nand U6027 (N_6027,N_5391,N_4099);
nor U6028 (N_6028,N_4464,N_5065);
or U6029 (N_6029,N_5129,N_4646);
or U6030 (N_6030,N_4724,N_4819);
nor U6031 (N_6031,N_5385,N_4773);
and U6032 (N_6032,N_5699,N_5104);
nor U6033 (N_6033,N_4930,N_5944);
and U6034 (N_6034,N_4463,N_4020);
nand U6035 (N_6035,N_4212,N_5214);
nor U6036 (N_6036,N_4224,N_5409);
and U6037 (N_6037,N_5893,N_4696);
or U6038 (N_6038,N_5766,N_4010);
nand U6039 (N_6039,N_5741,N_4260);
nand U6040 (N_6040,N_5051,N_5965);
nand U6041 (N_6041,N_5390,N_5223);
nand U6042 (N_6042,N_4108,N_4268);
or U6043 (N_6043,N_5654,N_4741);
nand U6044 (N_6044,N_4955,N_4862);
nor U6045 (N_6045,N_4319,N_5094);
or U6046 (N_6046,N_4748,N_4860);
nor U6047 (N_6047,N_4347,N_5307);
or U6048 (N_6048,N_5895,N_5992);
nand U6049 (N_6049,N_4112,N_5942);
nor U6050 (N_6050,N_5818,N_5281);
and U6051 (N_6051,N_4587,N_5675);
nand U6052 (N_6052,N_5729,N_5364);
nand U6053 (N_6053,N_5023,N_5138);
nor U6054 (N_6054,N_4826,N_5263);
or U6055 (N_6055,N_4547,N_5600);
or U6056 (N_6056,N_4417,N_5649);
nor U6057 (N_6057,N_4238,N_4273);
nand U6058 (N_6058,N_5287,N_5258);
and U6059 (N_6059,N_4595,N_5153);
nor U6060 (N_6060,N_4700,N_4082);
nand U6061 (N_6061,N_4406,N_4375);
nor U6062 (N_6062,N_4174,N_4439);
and U6063 (N_6063,N_5453,N_4118);
nor U6064 (N_6064,N_4690,N_4585);
and U6065 (N_6065,N_4834,N_4494);
nand U6066 (N_6066,N_5580,N_4294);
nand U6067 (N_6067,N_5720,N_4021);
and U6068 (N_6068,N_4757,N_4920);
or U6069 (N_6069,N_4577,N_4380);
nor U6070 (N_6070,N_4244,N_5977);
or U6071 (N_6071,N_5493,N_4777);
nor U6072 (N_6072,N_5742,N_5797);
and U6073 (N_6073,N_4345,N_4162);
nand U6074 (N_6074,N_5069,N_4673);
nor U6075 (N_6075,N_5745,N_5465);
or U6076 (N_6076,N_5925,N_5664);
nor U6077 (N_6077,N_4557,N_5292);
nor U6078 (N_6078,N_5557,N_4891);
or U6079 (N_6079,N_4833,N_4953);
or U6080 (N_6080,N_5770,N_4002);
nor U6081 (N_6081,N_4173,N_4402);
nand U6082 (N_6082,N_5508,N_5411);
nand U6083 (N_6083,N_4382,N_5363);
nor U6084 (N_6084,N_4308,N_4498);
nand U6085 (N_6085,N_5619,N_5632);
and U6086 (N_6086,N_5111,N_5016);
nand U6087 (N_6087,N_4994,N_5277);
or U6088 (N_6088,N_5290,N_5034);
nand U6089 (N_6089,N_5670,N_4869);
nor U6090 (N_6090,N_5640,N_5194);
or U6091 (N_6091,N_5131,N_5377);
nor U6092 (N_6092,N_4110,N_5617);
and U6093 (N_6093,N_4885,N_4671);
nor U6094 (N_6094,N_4986,N_5687);
or U6095 (N_6095,N_4535,N_4353);
nand U6096 (N_6096,N_5203,N_4900);
and U6097 (N_6097,N_5774,N_4289);
and U6098 (N_6098,N_5999,N_5451);
and U6099 (N_6099,N_4870,N_4471);
nand U6100 (N_6100,N_4205,N_5354);
nand U6101 (N_6101,N_5040,N_5714);
nor U6102 (N_6102,N_5512,N_5433);
nand U6103 (N_6103,N_4803,N_5859);
or U6104 (N_6104,N_5124,N_5161);
and U6105 (N_6105,N_5630,N_5744);
nand U6106 (N_6106,N_4430,N_4802);
nor U6107 (N_6107,N_4638,N_5436);
nand U6108 (N_6108,N_4662,N_4692);
nor U6109 (N_6109,N_5595,N_4753);
nand U6110 (N_6110,N_5958,N_4688);
nor U6111 (N_6111,N_4652,N_5884);
nor U6112 (N_6112,N_4519,N_5540);
and U6113 (N_6113,N_4137,N_4015);
and U6114 (N_6114,N_4602,N_4365);
nand U6115 (N_6115,N_4225,N_4706);
or U6116 (N_6116,N_4455,N_5303);
nor U6117 (N_6117,N_4114,N_5692);
nor U6118 (N_6118,N_5388,N_4343);
nor U6119 (N_6119,N_5082,N_4069);
or U6120 (N_6120,N_5042,N_4991);
and U6121 (N_6121,N_5836,N_5177);
or U6122 (N_6122,N_4668,N_4605);
nor U6123 (N_6123,N_4210,N_5015);
and U6124 (N_6124,N_4187,N_4873);
nand U6125 (N_6125,N_5850,N_4642);
nor U6126 (N_6126,N_5254,N_5284);
nand U6127 (N_6127,N_5817,N_4189);
nand U6128 (N_6128,N_5725,N_5355);
nand U6129 (N_6129,N_5353,N_5728);
and U6130 (N_6130,N_4880,N_5696);
or U6131 (N_6131,N_5046,N_5607);
nor U6132 (N_6132,N_4130,N_4946);
or U6133 (N_6133,N_5319,N_5505);
nand U6134 (N_6134,N_4124,N_5734);
nand U6135 (N_6135,N_5446,N_5765);
or U6136 (N_6136,N_4686,N_4395);
and U6137 (N_6137,N_4056,N_4877);
or U6138 (N_6138,N_5571,N_5936);
nor U6139 (N_6139,N_4301,N_4752);
nor U6140 (N_6140,N_4734,N_4102);
and U6141 (N_6141,N_5616,N_4221);
and U6142 (N_6142,N_5427,N_5459);
nand U6143 (N_6143,N_4483,N_5558);
xnor U6144 (N_6144,N_5101,N_4565);
or U6145 (N_6145,N_4135,N_4368);
nor U6146 (N_6146,N_5569,N_4336);
nor U6147 (N_6147,N_5775,N_4964);
nor U6148 (N_6148,N_4397,N_4160);
nand U6149 (N_6149,N_4447,N_4222);
nand U6150 (N_6150,N_5199,N_4335);
nor U6151 (N_6151,N_4934,N_5285);
xnor U6152 (N_6152,N_4188,N_5211);
nor U6153 (N_6153,N_5941,N_5230);
nor U6154 (N_6154,N_4396,N_5998);
and U6155 (N_6155,N_4051,N_5657);
nor U6156 (N_6156,N_5899,N_5268);
nor U6157 (N_6157,N_5969,N_4213);
or U6158 (N_6158,N_5423,N_5402);
and U6159 (N_6159,N_5227,N_5584);
or U6160 (N_6160,N_5927,N_5976);
or U6161 (N_6161,N_4278,N_5389);
nand U6162 (N_6162,N_4917,N_4959);
or U6163 (N_6163,N_5464,N_5394);
and U6164 (N_6164,N_5907,N_4825);
nor U6165 (N_6165,N_4563,N_5854);
and U6166 (N_6166,N_5458,N_5024);
or U6167 (N_6167,N_5869,N_4522);
nand U6168 (N_6168,N_5049,N_4941);
and U6169 (N_6169,N_4444,N_5887);
nor U6170 (N_6170,N_4903,N_5706);
nor U6171 (N_6171,N_5740,N_4579);
and U6172 (N_6172,N_4109,N_4630);
or U6173 (N_6173,N_4663,N_4156);
and U6174 (N_6174,N_5496,N_4526);
and U6175 (N_6175,N_4237,N_5321);
nand U6176 (N_6176,N_5064,N_4598);
nor U6177 (N_6177,N_4176,N_4229);
nor U6178 (N_6178,N_5231,N_5813);
nor U6179 (N_6179,N_4363,N_4525);
nor U6180 (N_6180,N_4474,N_4100);
nand U6181 (N_6181,N_4768,N_4867);
nand U6182 (N_6182,N_4352,N_4331);
nand U6183 (N_6183,N_5957,N_4028);
or U6184 (N_6184,N_4658,N_5066);
and U6185 (N_6185,N_4321,N_5076);
or U6186 (N_6186,N_4866,N_5542);
or U6187 (N_6187,N_4373,N_5297);
nand U6188 (N_6188,N_4208,N_4147);
nand U6189 (N_6189,N_5819,N_4501);
or U6190 (N_6190,N_4159,N_4705);
or U6191 (N_6191,N_4544,N_4383);
nor U6192 (N_6192,N_5244,N_5345);
and U6193 (N_6193,N_5135,N_5162);
and U6194 (N_6194,N_5862,N_4635);
and U6195 (N_6195,N_5786,N_5554);
and U6196 (N_6196,N_5803,N_5327);
nor U6197 (N_6197,N_4636,N_4687);
and U6198 (N_6198,N_4193,N_4664);
nand U6199 (N_6199,N_5329,N_4931);
nand U6200 (N_6200,N_5904,N_5515);
nand U6201 (N_6201,N_4209,N_4644);
or U6202 (N_6202,N_5431,N_4017);
nor U6203 (N_6203,N_5440,N_4923);
and U6204 (N_6204,N_5623,N_4703);
or U6205 (N_6205,N_5739,N_4327);
nand U6206 (N_6206,N_5946,N_4532);
nor U6207 (N_6207,N_4451,N_5840);
and U6208 (N_6208,N_4622,N_5020);
and U6209 (N_6209,N_5886,N_4496);
nand U6210 (N_6210,N_4812,N_5011);
and U6211 (N_6211,N_4702,N_5098);
nor U6212 (N_6212,N_5494,N_4165);
or U6213 (N_6213,N_4822,N_5748);
nand U6214 (N_6214,N_4035,N_4284);
nor U6215 (N_6215,N_4460,N_5676);
nand U6216 (N_6216,N_5337,N_4943);
or U6217 (N_6217,N_5374,N_5105);
or U6218 (N_6218,N_4276,N_5047);
nor U6219 (N_6219,N_4886,N_5634);
and U6220 (N_6220,N_5168,N_5532);
or U6221 (N_6221,N_5918,N_5057);
nand U6222 (N_6222,N_5003,N_5782);
and U6223 (N_6223,N_5274,N_5008);
nand U6224 (N_6224,N_5289,N_4072);
nand U6225 (N_6225,N_5638,N_5122);
or U6226 (N_6226,N_4066,N_5430);
nor U6227 (N_6227,N_5084,N_5302);
nand U6228 (N_6228,N_5982,N_5222);
and U6229 (N_6229,N_4486,N_4256);
or U6230 (N_6230,N_4307,N_4078);
or U6231 (N_6231,N_5609,N_5265);
nor U6232 (N_6232,N_5916,N_4408);
or U6233 (N_6233,N_4511,N_4259);
nor U6234 (N_6234,N_4361,N_4329);
nand U6235 (N_6235,N_5221,N_5789);
nor U6236 (N_6236,N_4197,N_5650);
nor U6237 (N_6237,N_4034,N_5983);
and U6238 (N_6238,N_4458,N_4824);
and U6239 (N_6239,N_5144,N_4710);
and U6240 (N_6240,N_4899,N_4914);
or U6241 (N_6241,N_4037,N_4123);
nand U6242 (N_6242,N_5680,N_5005);
nor U6243 (N_6243,N_4133,N_5644);
nor U6244 (N_6244,N_4263,N_5127);
and U6245 (N_6245,N_4280,N_5175);
or U6246 (N_6246,N_4154,N_4153);
nand U6247 (N_6247,N_4413,N_5039);
nand U6248 (N_6248,N_4846,N_4507);
nand U6249 (N_6249,N_4076,N_5647);
or U6250 (N_6250,N_5033,N_4104);
and U6251 (N_6251,N_5738,N_4003);
or U6252 (N_6252,N_4962,N_4876);
nor U6253 (N_6253,N_4929,N_5968);
nor U6254 (N_6254,N_4061,N_5404);
nor U6255 (N_6255,N_4033,N_5553);
nor U6256 (N_6256,N_4623,N_5063);
and U6257 (N_6257,N_5928,N_5160);
or U6258 (N_6258,N_4029,N_5723);
nor U6259 (N_6259,N_5943,N_4626);
nor U6260 (N_6260,N_5397,N_4290);
nor U6261 (N_6261,N_5294,N_5314);
or U6262 (N_6262,N_5460,N_4325);
nand U6263 (N_6263,N_5981,N_4401);
nor U6264 (N_6264,N_4332,N_4714);
nor U6265 (N_6265,N_5578,N_4012);
nor U6266 (N_6266,N_5419,N_5366);
and U6267 (N_6267,N_4954,N_4048);
nand U6268 (N_6268,N_4597,N_4951);
and U6269 (N_6269,N_4933,N_4407);
nor U6270 (N_6270,N_4218,N_5856);
nor U6271 (N_6271,N_5780,N_5615);
nor U6272 (N_6272,N_5116,N_4203);
and U6273 (N_6273,N_4310,N_5953);
and U6274 (N_6274,N_4973,N_5912);
nand U6275 (N_6275,N_4311,N_4369);
nand U6276 (N_6276,N_4235,N_5798);
nor U6277 (N_6277,N_4480,N_5858);
or U6278 (N_6278,N_5155,N_5257);
or U6279 (N_6279,N_5762,N_5035);
nor U6280 (N_6280,N_5031,N_4404);
nor U6281 (N_6281,N_4729,N_4279);
nand U6282 (N_6282,N_4359,N_5352);
nor U6283 (N_6283,N_4610,N_4845);
nor U6284 (N_6284,N_4791,N_4393);
nand U6285 (N_6285,N_5785,N_5506);
nand U6286 (N_6286,N_4233,N_5420);
and U6287 (N_6287,N_5189,N_4770);
nand U6288 (N_6288,N_5213,N_5087);
xor U6289 (N_6289,N_5022,N_5825);
nand U6290 (N_6290,N_5338,N_5081);
nor U6291 (N_6291,N_5191,N_4713);
and U6292 (N_6292,N_4682,N_4960);
or U6293 (N_6293,N_4220,N_5528);
or U6294 (N_6294,N_5585,N_4491);
nand U6295 (N_6295,N_5123,N_4913);
and U6296 (N_6296,N_5248,N_4848);
nor U6297 (N_6297,N_5658,N_5807);
nand U6298 (N_6298,N_4465,N_4739);
or U6299 (N_6299,N_5688,N_5761);
and U6300 (N_6300,N_4249,N_5448);
nand U6301 (N_6301,N_4574,N_5172);
and U6302 (N_6302,N_5684,N_5660);
and U6303 (N_6303,N_5639,N_4707);
or U6304 (N_6304,N_4691,N_4504);
or U6305 (N_6305,N_4423,N_4985);
nor U6306 (N_6306,N_5629,N_5896);
nand U6307 (N_6307,N_4517,N_4390);
or U6308 (N_6308,N_4889,N_4575);
and U6309 (N_6309,N_4792,N_4182);
or U6310 (N_6310,N_4409,N_5103);
nand U6311 (N_6311,N_4527,N_4115);
or U6312 (N_6312,N_5426,N_5048);
nand U6313 (N_6313,N_4730,N_5183);
nor U6314 (N_6314,N_5737,N_4919);
nor U6315 (N_6315,N_5661,N_5091);
and U6316 (N_6316,N_4853,N_5073);
or U6317 (N_6317,N_4489,N_5370);
and U6318 (N_6318,N_4436,N_4354);
and U6319 (N_6319,N_4795,N_4787);
nand U6320 (N_6320,N_4357,N_4841);
nand U6321 (N_6321,N_4419,N_4944);
or U6322 (N_6322,N_4031,N_4531);
nor U6323 (N_6323,N_5163,N_4788);
or U6324 (N_6324,N_5356,N_5822);
and U6325 (N_6325,N_5241,N_5266);
nor U6326 (N_6326,N_4910,N_5253);
nor U6327 (N_6327,N_4759,N_4871);
or U6328 (N_6328,N_5443,N_5567);
nand U6329 (N_6329,N_4470,N_4616);
nor U6330 (N_6330,N_5286,N_4588);
or U6331 (N_6331,N_5697,N_5546);
or U6332 (N_6332,N_4101,N_4288);
nor U6333 (N_6333,N_5837,N_5242);
nand U6334 (N_6334,N_4448,N_4855);
nand U6335 (N_6335,N_5962,N_4672);
nor U6336 (N_6336,N_5966,N_4183);
nand U6337 (N_6337,N_4851,N_4879);
nand U6338 (N_6338,N_4590,N_5824);
nand U6339 (N_6339,N_4667,N_5470);
nand U6340 (N_6340,N_5300,N_4651);
and U6341 (N_6341,N_5435,N_4231);
nand U6342 (N_6342,N_5061,N_5642);
and U6343 (N_6343,N_5335,N_4815);
and U6344 (N_6344,N_4685,N_4537);
nand U6345 (N_6345,N_4181,N_5502);
and U6346 (N_6346,N_4897,N_4117);
nor U6347 (N_6347,N_5849,N_5985);
nand U6348 (N_6348,N_4798,N_4157);
nand U6349 (N_6349,N_5756,N_5246);
nor U6350 (N_6350,N_4505,N_4661);
and U6351 (N_6351,N_5141,N_4150);
and U6352 (N_6352,N_5677,N_4026);
or U6353 (N_6353,N_5673,N_4405);
and U6354 (N_6354,N_5403,N_5413);
or U6355 (N_6355,N_5262,N_5897);
or U6356 (N_6356,N_5527,N_5442);
or U6357 (N_6357,N_4217,N_4950);
nand U6358 (N_6358,N_4184,N_5336);
or U6359 (N_6359,N_4230,N_4939);
nand U6360 (N_6360,N_4980,N_4472);
xnor U6361 (N_6361,N_4836,N_5873);
or U6362 (N_6362,N_5573,N_5783);
and U6363 (N_6363,N_5306,N_4457);
nor U6364 (N_6364,N_5703,N_4573);
and U6365 (N_6365,N_5273,N_5831);
nor U6366 (N_6366,N_4062,N_5679);
nor U6367 (N_6367,N_5523,N_5143);
nand U6368 (N_6368,N_5169,N_4570);
or U6369 (N_6369,N_4346,N_4640);
and U6370 (N_6370,N_5414,N_4119);
or U6371 (N_6371,N_5109,N_5216);
nand U6372 (N_6372,N_5513,N_4198);
or U6373 (N_6373,N_5624,N_4793);
nor U6374 (N_6374,N_4442,N_4993);
and U6375 (N_6375,N_4426,N_5823);
nor U6376 (N_6376,N_5806,N_4216);
and U6377 (N_6377,N_4418,N_4747);
nor U6378 (N_6378,N_4328,N_4271);
nand U6379 (N_6379,N_4978,N_5534);
nand U6380 (N_6380,N_4783,N_5373);
nor U6381 (N_6381,N_5683,N_4764);
nand U6382 (N_6382,N_4859,N_4424);
nand U6383 (N_6383,N_4997,N_4887);
nand U6384 (N_6384,N_4659,N_4786);
or U6385 (N_6385,N_4872,N_4136);
or U6386 (N_6386,N_5137,N_4578);
nor U6387 (N_6387,N_5256,N_5067);
or U6388 (N_6388,N_4297,N_4776);
or U6389 (N_6389,N_4735,N_5754);
nand U6390 (N_6390,N_4655,N_4949);
and U6391 (N_6391,N_4333,N_5967);
or U6392 (N_6392,N_4603,N_4890);
and U6393 (N_6393,N_4701,N_5272);
and U6394 (N_6394,N_4161,N_5767);
and U6395 (N_6395,N_4670,N_5462);
or U6396 (N_6396,N_5054,N_4064);
xnor U6397 (N_6397,N_5312,N_5056);
nand U6398 (N_6398,N_5583,N_4559);
nor U6399 (N_6399,N_4782,N_4170);
and U6400 (N_6400,N_4163,N_4742);
nand U6401 (N_6401,N_5857,N_4695);
and U6402 (N_6402,N_5827,N_5535);
and U6403 (N_6403,N_4657,N_5901);
or U6404 (N_6404,N_4234,N_5746);
and U6405 (N_6405,N_5694,N_5062);
or U6406 (N_6406,N_5950,N_4740);
nor U6407 (N_6407,N_4358,N_5233);
nand U6408 (N_6408,N_5628,N_5974);
nor U6409 (N_6409,N_5777,N_4269);
or U6410 (N_6410,N_5800,N_5551);
nand U6411 (N_6411,N_5814,N_4591);
or U6412 (N_6412,N_4817,N_4554);
or U6413 (N_6413,N_5150,N_4774);
nand U6414 (N_6414,N_4906,N_5592);
or U6415 (N_6415,N_4689,N_5010);
or U6416 (N_6416,N_5304,N_4716);
or U6417 (N_6417,N_5293,N_5167);
nor U6418 (N_6418,N_4192,N_4813);
nand U6419 (N_6419,N_5269,N_4582);
or U6420 (N_6420,N_4733,N_5705);
and U6421 (N_6421,N_5547,N_4190);
nand U6422 (N_6422,N_5951,N_5429);
nand U6423 (N_6423,N_5089,N_5587);
and U6424 (N_6424,N_4096,N_5112);
and U6425 (N_6425,N_4084,N_5483);
nand U6426 (N_6426,N_5905,N_4415);
or U6427 (N_6427,N_4175,N_5524);
nand U6428 (N_6428,N_4970,N_4625);
or U6429 (N_6429,N_5455,N_4374);
nand U6430 (N_6430,N_4024,N_5915);
and U6431 (N_6431,N_4720,N_4027);
nand U6432 (N_6432,N_4113,N_4966);
nor U6433 (N_6433,N_5668,N_4738);
nor U6434 (N_6434,N_5171,N_5898);
or U6435 (N_6435,N_4633,N_4987);
and U6436 (N_6436,N_4749,N_4172);
and U6437 (N_6437,N_5301,N_4767);
and U6438 (N_6438,N_4009,N_5317);
or U6439 (N_6439,N_5769,N_4000);
and U6440 (N_6440,N_5360,N_5669);
or U6441 (N_6441,N_4087,N_5633);
nor U6442 (N_6442,N_4487,N_5666);
or U6443 (N_6443,N_5522,N_5450);
or U6444 (N_6444,N_5090,N_4704);
nand U6445 (N_6445,N_4555,N_5764);
nor U6446 (N_6446,N_4907,N_5249);
nand U6447 (N_6447,N_4521,N_4433);
nand U6448 (N_6448,N_5621,N_5636);
and U6449 (N_6449,N_5146,N_4761);
nor U6450 (N_6450,N_5880,N_5727);
nor U6451 (N_6451,N_4828,N_5398);
and U6452 (N_6452,N_5136,N_4312);
and U6453 (N_6453,N_4728,N_5481);
nand U6454 (N_6454,N_4639,N_4398);
or U6455 (N_6455,N_4979,N_5971);
nand U6456 (N_6456,N_5499,N_4152);
nor U6457 (N_6457,N_5844,N_5845);
and U6458 (N_6458,N_5487,N_4837);
nor U6459 (N_6459,N_4892,N_4274);
and U6460 (N_6460,N_5201,N_5349);
or U6461 (N_6461,N_5026,N_5718);
and U6462 (N_6462,N_4275,N_5736);
nor U6463 (N_6463,N_5888,N_5559);
and U6464 (N_6464,N_4924,N_4344);
or U6465 (N_6465,N_5165,N_4006);
nand U6466 (N_6466,N_5288,N_5068);
nand U6467 (N_6467,N_5151,N_5472);
nor U6468 (N_6468,N_4830,N_5393);
or U6469 (N_6469,N_5325,N_5267);
nor U6470 (N_6470,N_4482,N_4131);
and U6471 (N_6471,N_4059,N_5986);
nand U6472 (N_6472,N_4403,N_5842);
nor U6473 (N_6473,N_5802,N_5461);
nand U6474 (N_6474,N_4469,N_4512);
nor U6475 (N_6475,N_4242,N_4057);
nor U6476 (N_6476,N_4901,N_4098);
or U6477 (N_6477,N_4684,N_4542);
nand U6478 (N_6478,N_5626,N_4604);
nor U6479 (N_6479,N_5291,N_5358);
or U6480 (N_6480,N_4778,N_4141);
and U6481 (N_6481,N_5948,N_4902);
nor U6482 (N_6482,N_5456,N_4434);
nand U6483 (N_6483,N_5596,N_4932);
nor U6484 (N_6484,N_5715,N_4937);
nor U6485 (N_6485,N_5204,N_5340);
and U6486 (N_6486,N_5790,N_4552);
nand U6487 (N_6487,N_5710,N_4553);
and U6488 (N_6488,N_5605,N_4041);
nor U6489 (N_6489,N_5846,N_5519);
and U6490 (N_6490,N_4410,N_5305);
or U6491 (N_6491,N_5804,N_4536);
nand U6492 (N_6492,N_5334,N_5516);
nor U6493 (N_6493,N_4818,N_5000);
and U6494 (N_6494,N_5331,N_5179);
or U6495 (N_6495,N_4617,N_4807);
nand U6496 (N_6496,N_4011,N_4619);
nor U6497 (N_6497,N_4840,N_4202);
or U6498 (N_6498,N_5295,N_5280);
nor U6499 (N_6499,N_5341,N_4298);
nand U6500 (N_6500,N_4372,N_4518);
nand U6501 (N_6501,N_4385,N_4223);
or U6502 (N_6502,N_5195,N_5326);
and U6503 (N_6503,N_4865,N_5938);
and U6504 (N_6504,N_4453,N_4111);
or U6505 (N_6505,N_5730,N_5815);
nand U6506 (N_6506,N_4925,N_5164);
or U6507 (N_6507,N_4534,N_5247);
nor U6508 (N_6508,N_5013,N_4529);
nor U6509 (N_6509,N_4106,N_5731);
or U6510 (N_6510,N_5611,N_5126);
nand U6511 (N_6511,N_5415,N_4264);
and U6512 (N_6512,N_5539,N_5663);
nand U6513 (N_6513,N_4351,N_5296);
or U6514 (N_6514,N_4255,N_4799);
nor U6515 (N_6515,N_4513,N_5120);
or U6516 (N_6516,N_5028,N_4005);
or U6517 (N_6517,N_4550,N_4942);
and U6518 (N_6518,N_5032,N_5085);
and U6519 (N_6519,N_5900,N_5987);
or U6520 (N_6520,N_4341,N_5434);
nand U6521 (N_6521,N_5879,N_4606);
nand U6522 (N_6522,N_4854,N_5635);
and U6523 (N_6523,N_5695,N_4567);
or U6524 (N_6524,N_5816,N_5102);
and U6525 (N_6525,N_4095,N_5919);
or U6526 (N_6526,N_5202,N_5488);
nand U6527 (N_6527,N_4744,N_5174);
nor U6528 (N_6528,N_5758,N_5781);
nand U6529 (N_6529,N_4806,N_4971);
or U6530 (N_6530,N_5041,N_5652);
nand U6531 (N_6531,N_4116,N_4694);
and U6532 (N_6532,N_4476,N_4990);
and U6533 (N_6533,N_5372,N_5252);
nand U6534 (N_6534,N_4790,N_4989);
xnor U6535 (N_6535,N_4304,N_4581);
nand U6536 (N_6536,N_5132,N_5468);
and U6537 (N_6537,N_5342,N_5829);
nor U6538 (N_6538,N_5989,N_5747);
nor U6539 (N_6539,N_4167,N_4725);
and U6540 (N_6540,N_5096,N_4196);
nor U6541 (N_6541,N_4431,N_5348);
nor U6542 (N_6542,N_5952,N_5079);
and U6543 (N_6543,N_4940,N_5591);
nor U6544 (N_6544,N_5083,N_5332);
and U6545 (N_6545,N_5631,N_5119);
and U6546 (N_6546,N_5387,N_5541);
or U6547 (N_6547,N_5560,N_5838);
nand U6548 (N_6548,N_5469,N_5793);
nand U6549 (N_6549,N_5550,N_5218);
or U6550 (N_6550,N_4750,N_4070);
or U6551 (N_6551,N_4645,N_4832);
or U6552 (N_6552,N_4722,N_5344);
nand U6553 (N_6553,N_4811,N_5324);
or U6554 (N_6554,N_5978,N_5796);
nand U6555 (N_6555,N_5543,N_5937);
and U6556 (N_6556,N_4765,N_4983);
nand U6557 (N_6557,N_4754,N_4340);
or U6558 (N_6558,N_5521,N_4416);
nor U6559 (N_6559,N_4243,N_5545);
nand U6560 (N_6560,N_4601,N_4756);
or U6561 (N_6561,N_4656,N_4318);
nor U6562 (N_6562,N_4267,N_4211);
and U6563 (N_6563,N_5810,N_4322);
nand U6564 (N_6564,N_5812,N_4050);
and U6565 (N_6565,N_5601,N_5361);
nand U6566 (N_6566,N_4326,N_4240);
nor U6567 (N_6567,N_4252,N_4206);
nand U6568 (N_6568,N_4620,N_4400);
and U6569 (N_6569,N_5475,N_5995);
or U6570 (N_6570,N_4166,N_5238);
nor U6571 (N_6571,N_4755,N_4088);
nor U6572 (N_6572,N_5490,N_4085);
and U6573 (N_6573,N_5713,N_5416);
or U6574 (N_6574,N_4775,N_4299);
or U6575 (N_6575,N_5622,N_5125);
nor U6576 (N_6576,N_5892,N_5315);
and U6577 (N_6577,N_4334,N_4982);
nor U6578 (N_6578,N_4816,N_4239);
nor U6579 (N_6579,N_5643,N_4467);
nor U6580 (N_6580,N_5614,N_5072);
nand U6581 (N_6581,N_4503,N_4381);
nand U6582 (N_6582,N_4497,N_4936);
nand U6583 (N_6583,N_5667,N_5250);
or U6584 (N_6584,N_5474,N_5186);
and U6585 (N_6585,N_4339,N_4999);
nand U6586 (N_6586,N_4984,N_5128);
nand U6587 (N_6587,N_4073,N_5940);
and U6588 (N_6588,N_4364,N_5240);
or U6589 (N_6589,N_5702,N_4679);
and U6590 (N_6590,N_4829,N_4612);
and U6591 (N_6591,N_4571,N_5444);
or U6592 (N_6592,N_5808,N_4814);
or U6593 (N_6593,N_5525,N_5597);
nor U6594 (N_6594,N_4105,N_4277);
nor U6595 (N_6595,N_4810,N_4916);
or U6596 (N_6596,N_5834,N_5359);
nor U6597 (N_6597,N_5574,N_5653);
or U6598 (N_6598,N_5779,N_4697);
or U6599 (N_6599,N_5130,N_4246);
nor U6600 (N_6600,N_5572,N_4081);
nor U6601 (N_6601,N_5577,N_5159);
nand U6602 (N_6602,N_5365,N_5964);
and U6603 (N_6603,N_4143,N_5832);
or U6604 (N_6604,N_5392,N_4882);
nand U6605 (N_6605,N_5092,N_5417);
or U6606 (N_6606,N_4562,N_4731);
and U6607 (N_6607,N_4195,N_4998);
nor U6608 (N_6608,N_5922,N_5707);
and U6609 (N_6609,N_4712,N_4360);
and U6610 (N_6610,N_5107,N_5841);
and U6611 (N_6611,N_5801,N_5001);
or U6612 (N_6612,N_5424,N_4607);
nand U6613 (N_6613,N_5264,N_5339);
nor U6614 (N_6614,N_5382,N_5428);
and U6615 (N_6615,N_4842,N_5030);
or U6616 (N_6616,N_5371,N_5552);
and U6617 (N_6617,N_4387,N_5828);
xor U6618 (N_6618,N_4908,N_5115);
or U6619 (N_6619,N_4628,N_5870);
or U6620 (N_6620,N_4875,N_4435);
and U6621 (N_6621,N_5544,N_5439);
nand U6622 (N_6622,N_5278,N_4743);
and U6623 (N_6623,N_4286,N_4805);
and U6624 (N_6624,N_4947,N_4769);
nand U6625 (N_6625,N_5963,N_4796);
nand U6626 (N_6626,N_5106,N_4568);
nor U6627 (N_6627,N_5934,N_5215);
and U6628 (N_6628,N_5691,N_5701);
or U6629 (N_6629,N_5362,N_5055);
or U6630 (N_6630,N_5311,N_5755);
nand U6631 (N_6631,N_4459,N_4847);
nor U6632 (N_6632,N_4120,N_4258);
or U6633 (N_6633,N_5205,N_5408);
or U6634 (N_6634,N_4261,N_4727);
and U6635 (N_6635,N_5561,N_5484);
and U6636 (N_6636,N_5449,N_4194);
and U6637 (N_6637,N_5889,N_4838);
nand U6638 (N_6638,N_5996,N_5478);
and U6639 (N_6639,N_5590,N_5973);
and U6640 (N_6640,N_5038,N_5333);
nand U6641 (N_6641,N_4456,N_5993);
nand U6642 (N_6642,N_4449,N_4052);
nand U6643 (N_6643,N_4926,N_4935);
and U6644 (N_6644,N_5871,N_5980);
or U6645 (N_6645,N_5347,N_5913);
and U6646 (N_6646,N_5923,N_5787);
nand U6647 (N_6647,N_5320,N_5396);
or U6648 (N_6648,N_4036,N_5099);
or U6649 (N_6649,N_5504,N_5768);
or U6650 (N_6650,N_4611,N_4291);
nand U6651 (N_6651,N_5708,N_4414);
or U6652 (N_6652,N_4077,N_5997);
nor U6653 (N_6653,N_4450,N_5627);
and U6654 (N_6654,N_5612,N_4647);
or U6655 (N_6655,N_5581,N_4250);
and U6656 (N_6656,N_4178,N_5509);
xnor U6657 (N_6657,N_4241,N_5848);
nor U6658 (N_6658,N_4219,N_5589);
or U6659 (N_6659,N_4797,N_5861);
and U6660 (N_6660,N_5145,N_5009);
nor U6661 (N_6661,N_5412,N_4377);
or U6662 (N_6662,N_5637,N_4479);
or U6663 (N_6663,N_5275,N_5316);
nor U6664 (N_6664,N_5751,N_5322);
and U6665 (N_6665,N_5491,N_5452);
nand U6666 (N_6666,N_5750,N_4569);
nor U6667 (N_6667,N_4624,N_5865);
nand U6668 (N_6668,N_4389,N_5473);
or U6669 (N_6669,N_5236,N_5234);
or U6670 (N_6670,N_4721,N_4254);
nor U6671 (N_6671,N_4745,N_5113);
nor U6672 (N_6672,N_5722,N_4063);
nor U6673 (N_6673,N_5752,N_4593);
nand U6674 (N_6674,N_5432,N_5197);
or U6675 (N_6675,N_5878,N_4893);
or U6676 (N_6676,N_4618,N_5270);
nor U6677 (N_6677,N_4122,N_5375);
nand U6678 (N_6678,N_4632,N_5479);
xnor U6679 (N_6679,N_4648,N_4948);
nor U6680 (N_6680,N_4008,N_5058);
nor U6681 (N_6681,N_5564,N_5743);
or U6682 (N_6682,N_5733,N_4018);
or U6683 (N_6683,N_4475,N_5721);
nor U6684 (N_6684,N_5579,N_4839);
nor U6685 (N_6685,N_5097,N_5309);
nand U6686 (N_6686,N_4683,N_5209);
nor U6687 (N_6687,N_4762,N_4967);
nor U6688 (N_6688,N_4452,N_4650);
nand U6689 (N_6689,N_4746,N_4065);
or U6690 (N_6690,N_4420,N_5610);
and U6691 (N_6691,N_4466,N_5685);
or U6692 (N_6692,N_5839,N_4583);
nand U6693 (N_6693,N_4199,N_5050);
nand U6694 (N_6694,N_5386,N_5157);
nor U6695 (N_6695,N_5480,N_5598);
or U6696 (N_6696,N_4060,N_4228);
nand U6697 (N_6697,N_4961,N_5517);
nand U6698 (N_6698,N_5088,N_4324);
nor U6699 (N_6699,N_5704,N_5225);
and U6700 (N_6700,N_5932,N_4007);
nor U6701 (N_6701,N_5909,N_4158);
nor U6702 (N_6702,N_4523,N_4251);
nor U6703 (N_6703,N_5681,N_5004);
nand U6704 (N_6704,N_5466,N_4490);
and U6705 (N_6705,N_5735,N_5029);
and U6706 (N_6706,N_5027,N_5226);
or U6707 (N_6707,N_4337,N_5014);
and U6708 (N_6708,N_4493,N_5792);
nand U6709 (N_6709,N_4809,N_4438);
and U6710 (N_6710,N_4495,N_4693);
nand U6711 (N_6711,N_4185,N_5310);
and U6712 (N_6712,N_5298,N_4053);
and U6713 (N_6713,N_4766,N_4589);
nand U6714 (N_6714,N_5019,N_4412);
nor U6715 (N_6715,N_4093,N_5548);
and U6716 (N_6716,N_4868,N_5776);
nor U6717 (N_6717,N_4560,N_5877);
nand U6718 (N_6718,N_5860,N_4758);
nand U6719 (N_6719,N_5261,N_4134);
nor U6720 (N_6720,N_5911,N_5118);
xnor U6721 (N_6721,N_4171,N_4388);
nor U6722 (N_6722,N_5100,N_5259);
nand U6723 (N_6723,N_4711,N_5229);
and U6724 (N_6724,N_4266,N_5075);
nor U6725 (N_6725,N_5712,N_5217);
and U6726 (N_6726,N_5152,N_4032);
or U6727 (N_6727,N_5613,N_5902);
nor U6728 (N_6728,N_5193,N_5947);
and U6729 (N_6729,N_4772,N_5243);
nand U6730 (N_6730,N_4481,N_4677);
nor U6731 (N_6731,N_5778,N_4366);
and U6732 (N_6732,N_4874,N_4981);
or U6733 (N_6733,N_4596,N_5093);
nand U6734 (N_6734,N_4678,N_4399);
and U6735 (N_6735,N_4548,N_5820);
and U6736 (N_6736,N_4976,N_5220);
or U6737 (N_6737,N_4992,N_5530);
and U6738 (N_6738,N_4821,N_5891);
or U6739 (N_6739,N_5485,N_4956);
or U6740 (N_6740,N_5863,N_4996);
nor U6741 (N_6741,N_4080,N_4878);
nand U6742 (N_6742,N_4168,N_4058);
and U6743 (N_6743,N_5763,N_4468);
and U6744 (N_6744,N_4751,N_5139);
and U6745 (N_6745,N_5173,N_5021);
nor U6746 (N_6746,N_4149,N_5176);
and U6747 (N_6747,N_5074,N_5855);
nand U6748 (N_6748,N_4313,N_5182);
nor U6749 (N_6749,N_4801,N_4509);
nand U6750 (N_6750,N_4576,N_5196);
and U6751 (N_6751,N_4349,N_5235);
nor U6752 (N_6752,N_5979,N_5575);
nand U6753 (N_6753,N_5467,N_4317);
or U6754 (N_6754,N_5700,N_4265);
and U6755 (N_6755,N_4394,N_5346);
and U6756 (N_6756,N_4049,N_4075);
nand U6757 (N_6757,N_5043,N_5709);
or U6758 (N_6758,N_5537,N_4362);
nand U6759 (N_6759,N_4510,N_4835);
nand U6760 (N_6760,N_4905,N_4040);
nor U6761 (N_6761,N_4309,N_5166);
and U6762 (N_6762,N_4022,N_4145);
nand U6763 (N_6763,N_4898,N_5184);
nand U6764 (N_6764,N_5108,N_4392);
and U6765 (N_6765,N_5955,N_4427);
nand U6766 (N_6766,N_5418,N_4586);
nand U6767 (N_6767,N_4492,N_4440);
and U6768 (N_6768,N_4132,N_4200);
nor U6769 (N_6769,N_5903,N_5181);
and U6770 (N_6770,N_5593,N_4054);
or U6771 (N_6771,N_5447,N_4086);
or U6772 (N_6772,N_4584,N_5984);
nand U6773 (N_6773,N_4641,N_4107);
nand U6774 (N_6774,N_4247,N_4039);
nor U6775 (N_6775,N_4484,N_4784);
or U6776 (N_6776,N_5192,N_4091);
or U6777 (N_6777,N_4478,N_5401);
or U6778 (N_6778,N_5457,N_4316);
or U6779 (N_6779,N_4609,N_4293);
nand U6780 (N_6780,N_4074,N_5686);
nor U6781 (N_6781,N_5949,N_5437);
nand U6782 (N_6782,N_4631,N_4637);
or U6783 (N_6783,N_4214,N_4043);
or U6784 (N_6784,N_4314,N_4718);
nor U6785 (N_6785,N_4038,N_5228);
and U6786 (N_6786,N_4356,N_5549);
or U6787 (N_6787,N_4621,N_4445);
and U6788 (N_6788,N_5588,N_5868);
nand U6789 (N_6789,N_4128,N_4090);
nor U6790 (N_6790,N_4653,N_5299);
nand U6791 (N_6791,N_4384,N_5711);
and U6792 (N_6792,N_4083,N_4995);
nor U6793 (N_6793,N_4437,N_5603);
xnor U6794 (N_6794,N_5835,N_5656);
nand U6795 (N_6795,N_5180,N_5566);
nand U6796 (N_6796,N_5975,N_4615);
nand U6797 (N_6797,N_4600,N_4425);
nor U6798 (N_6798,N_5843,N_5939);
nor U6799 (N_6799,N_4763,N_4300);
nor U6800 (N_6800,N_4047,N_5463);
nor U6801 (N_6801,N_4699,N_5501);
and U6802 (N_6802,N_5929,N_5395);
or U6803 (N_6803,N_5350,N_5381);
and U6804 (N_6804,N_4780,N_5674);
nor U6805 (N_6805,N_5935,N_4285);
nand U6806 (N_6806,N_5117,N_4046);
or U6807 (N_6807,N_5059,N_5187);
nand U6808 (N_6808,N_5271,N_5219);
and U6809 (N_6809,N_5659,N_4226);
xnor U6810 (N_6810,N_4515,N_4025);
nand U6811 (N_6811,N_5771,N_4379);
and U6812 (N_6812,N_5960,N_4191);
nand U6813 (N_6813,N_4675,N_4227);
or U6814 (N_6814,N_5283,N_4421);
nand U6815 (N_6815,N_4454,N_5945);
and U6816 (N_6816,N_4975,N_5421);
or U6817 (N_6817,N_4169,N_4127);
nand U6818 (N_6818,N_4634,N_5682);
nor U6819 (N_6819,N_4895,N_5784);
or U6820 (N_6820,N_5753,N_4262);
or U6821 (N_6821,N_4963,N_4295);
nand U6822 (N_6822,N_4928,N_5380);
nor U6823 (N_6823,N_5045,N_4922);
or U6824 (N_6824,N_4338,N_4945);
nand U6825 (N_6825,N_5095,N_4528);
nor U6826 (N_6826,N_5520,N_4681);
or U6827 (N_6827,N_4079,N_5618);
and U6828 (N_6828,N_4138,N_4330);
and U6829 (N_6829,N_4977,N_4972);
nor U6830 (N_6830,N_4785,N_4843);
nor U6831 (N_6831,N_5693,N_4958);
and U6832 (N_6832,N_4140,N_4236);
and U6833 (N_6833,N_4023,N_4303);
nand U6834 (N_6834,N_4863,N_5805);
or U6835 (N_6835,N_5279,N_4514);
and U6836 (N_6836,N_5495,N_4092);
or U6837 (N_6837,N_5492,N_4857);
or U6838 (N_6838,N_5323,N_5036);
and U6839 (N_6839,N_4441,N_5148);
and U6840 (N_6840,N_5749,N_5874);
nand U6841 (N_6841,N_5134,N_4551);
nor U6842 (N_6842,N_4546,N_5140);
or U6843 (N_6843,N_4726,N_5060);
nand U6844 (N_6844,N_4030,N_5052);
and U6845 (N_6845,N_5511,N_4257);
nor U6846 (N_6846,N_4477,N_5477);
nor U6847 (N_6847,N_4281,N_4827);
or U6848 (N_6848,N_5376,N_5678);
or U6849 (N_6849,N_4524,N_5518);
or U6850 (N_6850,N_4629,N_4067);
or U6851 (N_6851,N_4530,N_5641);
nand U6852 (N_6852,N_4320,N_5568);
nand U6853 (N_6853,N_5799,N_4779);
nor U6854 (N_6854,N_5556,N_4594);
nor U6855 (N_6855,N_4391,N_5400);
nor U6856 (N_6856,N_5933,N_5190);
or U6857 (N_6857,N_4654,N_4896);
nand U6858 (N_6858,N_4561,N_4068);
nor U6859 (N_6859,N_4820,N_4155);
nor U6860 (N_6860,N_4323,N_5882);
nand U6861 (N_6861,N_4355,N_5282);
nand U6862 (N_6862,N_4539,N_5121);
nand U6863 (N_6863,N_5086,N_5991);
nand U6864 (N_6864,N_5454,N_5489);
and U6865 (N_6865,N_5507,N_4386);
or U6866 (N_6866,N_4055,N_5794);
nand U6867 (N_6867,N_5671,N_5498);
nand U6868 (N_6868,N_5864,N_4506);
nor U6869 (N_6869,N_4432,N_4558);
nor U6870 (N_6870,N_4760,N_4852);
or U6871 (N_6871,N_4864,N_4894);
or U6872 (N_6872,N_4488,N_5533);
or U6873 (N_6873,N_4350,N_5866);
nor U6874 (N_6874,N_4473,N_4207);
nand U6875 (N_6875,N_5170,N_4253);
nand U6876 (N_6876,N_5881,N_5422);
nor U6877 (N_6877,N_4177,N_5018);
xnor U6878 (N_6878,N_5441,N_5133);
nand U6879 (N_6879,N_4858,N_5555);
nand U6880 (N_6880,N_4094,N_5239);
nand U6881 (N_6881,N_5689,N_5830);
nor U6882 (N_6882,N_4014,N_4044);
nor U6883 (N_6883,N_5867,N_5809);
or U6884 (N_6884,N_5662,N_5276);
and U6885 (N_6885,N_4915,N_5007);
nand U6886 (N_6886,N_5852,N_5497);
nor U6887 (N_6887,N_5037,N_5811);
and U6888 (N_6888,N_5833,N_5924);
nor U6889 (N_6889,N_5646,N_5576);
nand U6890 (N_6890,N_4909,N_4342);
nand U6891 (N_6891,N_5531,N_5482);
or U6892 (N_6892,N_4004,N_5926);
nand U6893 (N_6893,N_4502,N_5405);
nor U6894 (N_6894,N_5914,N_4856);
and U6895 (N_6895,N_5760,N_5921);
or U6896 (N_6896,N_4921,N_4883);
nand U6897 (N_6897,N_4411,N_4974);
and U6898 (N_6898,N_5308,N_4794);
nand U6899 (N_6899,N_5994,N_4013);
or U6900 (N_6900,N_4306,N_4443);
nand U6901 (N_6901,N_5255,N_4781);
nor U6902 (N_6902,N_5772,N_5970);
or U6903 (N_6903,N_4904,N_5961);
or U6904 (N_6904,N_5563,N_5906);
nor U6905 (N_6905,N_4680,N_5476);
xor U6906 (N_6906,N_5759,N_5445);
and U6907 (N_6907,N_4180,N_4627);
nor U6908 (N_6908,N_4808,N_4302);
and U6909 (N_6909,N_5399,N_5425);
nor U6910 (N_6910,N_4572,N_4968);
or U6911 (N_6911,N_4305,N_4103);
nor U6912 (N_6912,N_5212,N_4541);
nand U6913 (N_6913,N_4533,N_5237);
or U6914 (N_6914,N_4608,N_5158);
nor U6915 (N_6915,N_5990,N_5200);
and U6916 (N_6916,N_5606,N_4566);
nor U6917 (N_6917,N_5851,N_5757);
and U6918 (N_6918,N_5077,N_5908);
nand U6919 (N_6919,N_4376,N_5672);
nor U6920 (N_6920,N_4698,N_5357);
or U6921 (N_6921,N_5956,N_4348);
xor U6922 (N_6922,N_4282,N_5795);
or U6923 (N_6923,N_5788,N_4287);
nand U6924 (N_6924,N_5872,N_4139);
nor U6925 (N_6925,N_4676,N_5885);
nand U6926 (N_6926,N_4614,N_4001);
nand U6927 (N_6927,N_5407,N_4499);
and U6928 (N_6928,N_5500,N_4669);
or U6929 (N_6929,N_4719,N_5565);
nand U6930 (N_6930,N_4248,N_5954);
and U6931 (N_6931,N_5570,N_5328);
nand U6932 (N_6932,N_5698,N_4204);
xor U6933 (N_6933,N_5599,N_4717);
nand U6934 (N_6934,N_5198,N_5351);
and U6935 (N_6935,N_4927,N_5604);
nand U6936 (N_6936,N_4097,N_4823);
nor U6937 (N_6937,N_5582,N_4545);
or U6938 (N_6938,N_5875,N_5586);
nor U6939 (N_6939,N_5156,N_5207);
nand U6940 (N_6940,N_5368,N_4121);
nor U6941 (N_6941,N_5486,N_5330);
nand U6942 (N_6942,N_5847,N_5110);
nor U6943 (N_6943,N_4715,N_5645);
xnor U6944 (N_6944,N_4643,N_5260);
and U6945 (N_6945,N_4736,N_5726);
nand U6946 (N_6946,N_4660,N_4016);
or U6947 (N_6947,N_5208,N_4508);
nand U6948 (N_6948,N_5080,N_5071);
and U6949 (N_6949,N_5625,N_5826);
nand U6950 (N_6950,N_4378,N_4844);
and U6951 (N_6951,N_4089,N_4129);
nand U6952 (N_6952,N_4201,N_4649);
and U6953 (N_6953,N_5510,N_4164);
nor U6954 (N_6954,N_4462,N_5594);
or U6955 (N_6955,N_5773,N_4538);
nor U6956 (N_6956,N_5724,N_5920);
nor U6957 (N_6957,N_4912,N_5070);
nand U6958 (N_6958,N_4272,N_4019);
or U6959 (N_6959,N_4831,N_5154);
and U6960 (N_6960,N_4146,N_5006);
and U6961 (N_6961,N_5210,N_5716);
and U6962 (N_6962,N_4861,N_4911);
or U6963 (N_6963,N_4881,N_4737);
and U6964 (N_6964,N_4952,N_4957);
or U6965 (N_6965,N_5665,N_5369);
nand U6966 (N_6966,N_5185,N_5890);
or U6967 (N_6967,N_5406,N_5078);
nor U6968 (N_6968,N_4580,N_4665);
nand U6969 (N_6969,N_4850,N_4126);
and U6970 (N_6970,N_5620,N_4422);
nand U6971 (N_6971,N_4549,N_5917);
or U6972 (N_6972,N_5536,N_4485);
or U6973 (N_6973,N_5972,N_4938);
and U6974 (N_6974,N_4543,N_5538);
and U6975 (N_6975,N_4125,N_4849);
and U6976 (N_6976,N_4283,N_4071);
nand U6977 (N_6977,N_4148,N_5910);
nor U6978 (N_6978,N_5383,N_4232);
and U6979 (N_6979,N_5379,N_5017);
nand U6980 (N_6980,N_4429,N_5821);
and U6981 (N_6981,N_4367,N_5931);
and U6982 (N_6982,N_5044,N_5562);
or U6983 (N_6983,N_4709,N_4315);
or U6984 (N_6984,N_5378,N_5114);
or U6985 (N_6985,N_4708,N_5178);
or U6986 (N_6986,N_4804,N_4674);
nor U6987 (N_6987,N_5025,N_4520);
nor U6988 (N_6988,N_4371,N_5367);
and U6989 (N_6989,N_4186,N_4270);
or U6990 (N_6990,N_4142,N_4446);
or U6991 (N_6991,N_5690,N_5655);
and U6992 (N_6992,N_5012,N_4613);
nand U6993 (N_6993,N_5503,N_5147);
nor U6994 (N_6994,N_5142,N_4988);
and U6995 (N_6995,N_5883,N_4965);
and U6996 (N_6996,N_4296,N_4045);
nand U6997 (N_6997,N_5930,N_4042);
nor U6998 (N_6998,N_5206,N_4732);
and U6999 (N_6999,N_5853,N_4500);
or U7000 (N_7000,N_4745,N_4077);
nor U7001 (N_7001,N_5991,N_4592);
or U7002 (N_7002,N_5776,N_4225);
or U7003 (N_7003,N_4033,N_4130);
nand U7004 (N_7004,N_5386,N_5847);
or U7005 (N_7005,N_5604,N_5920);
or U7006 (N_7006,N_4536,N_5726);
or U7007 (N_7007,N_4205,N_4275);
nand U7008 (N_7008,N_5869,N_5931);
nor U7009 (N_7009,N_4376,N_5328);
and U7010 (N_7010,N_4099,N_4930);
nor U7011 (N_7011,N_5625,N_5278);
nor U7012 (N_7012,N_5264,N_4669);
nand U7013 (N_7013,N_5710,N_5988);
and U7014 (N_7014,N_4101,N_4291);
and U7015 (N_7015,N_5897,N_5525);
nand U7016 (N_7016,N_5978,N_5831);
and U7017 (N_7017,N_5697,N_4083);
and U7018 (N_7018,N_4713,N_5636);
or U7019 (N_7019,N_4162,N_5414);
or U7020 (N_7020,N_5792,N_4113);
nand U7021 (N_7021,N_4842,N_4332);
and U7022 (N_7022,N_4833,N_4416);
or U7023 (N_7023,N_4686,N_4147);
and U7024 (N_7024,N_4577,N_4101);
nor U7025 (N_7025,N_4131,N_5800);
nand U7026 (N_7026,N_4747,N_4202);
xnor U7027 (N_7027,N_4085,N_5740);
nand U7028 (N_7028,N_4909,N_5659);
nand U7029 (N_7029,N_4996,N_4111);
and U7030 (N_7030,N_4129,N_5552);
and U7031 (N_7031,N_5026,N_5626);
nand U7032 (N_7032,N_4460,N_5576);
nand U7033 (N_7033,N_5892,N_4009);
nor U7034 (N_7034,N_4521,N_4701);
and U7035 (N_7035,N_4247,N_5796);
nand U7036 (N_7036,N_5341,N_5676);
and U7037 (N_7037,N_5030,N_5493);
and U7038 (N_7038,N_5560,N_5534);
nand U7039 (N_7039,N_5801,N_5524);
nor U7040 (N_7040,N_5395,N_5603);
nand U7041 (N_7041,N_5519,N_4947);
and U7042 (N_7042,N_5645,N_5424);
nand U7043 (N_7043,N_5126,N_5113);
nand U7044 (N_7044,N_5616,N_4295);
nand U7045 (N_7045,N_4269,N_4936);
nor U7046 (N_7046,N_4945,N_4661);
or U7047 (N_7047,N_4028,N_5200);
nor U7048 (N_7048,N_5893,N_5454);
nor U7049 (N_7049,N_5901,N_4303);
nor U7050 (N_7050,N_5801,N_5458);
or U7051 (N_7051,N_4329,N_4779);
and U7052 (N_7052,N_4394,N_5919);
and U7053 (N_7053,N_5069,N_4639);
or U7054 (N_7054,N_4380,N_5708);
nor U7055 (N_7055,N_5761,N_5776);
and U7056 (N_7056,N_5014,N_5264);
nand U7057 (N_7057,N_4060,N_5081);
and U7058 (N_7058,N_5789,N_5862);
nand U7059 (N_7059,N_4883,N_4344);
nor U7060 (N_7060,N_5567,N_5551);
and U7061 (N_7061,N_4873,N_4346);
nor U7062 (N_7062,N_4459,N_5088);
and U7063 (N_7063,N_4642,N_5050);
and U7064 (N_7064,N_5286,N_5681);
nand U7065 (N_7065,N_5850,N_5405);
nand U7066 (N_7066,N_4205,N_4374);
or U7067 (N_7067,N_5518,N_5840);
nand U7068 (N_7068,N_4821,N_5741);
nand U7069 (N_7069,N_5879,N_4871);
nor U7070 (N_7070,N_4896,N_5995);
or U7071 (N_7071,N_5336,N_4473);
nor U7072 (N_7072,N_5923,N_5455);
nor U7073 (N_7073,N_5076,N_5327);
nor U7074 (N_7074,N_4709,N_5961);
or U7075 (N_7075,N_4663,N_4590);
nor U7076 (N_7076,N_5714,N_5739);
nor U7077 (N_7077,N_5874,N_4443);
nor U7078 (N_7078,N_4957,N_4242);
or U7079 (N_7079,N_4480,N_4245);
or U7080 (N_7080,N_4888,N_5915);
nand U7081 (N_7081,N_5210,N_5848);
nand U7082 (N_7082,N_4332,N_4031);
nand U7083 (N_7083,N_4132,N_4854);
and U7084 (N_7084,N_5589,N_4646);
and U7085 (N_7085,N_5227,N_5196);
or U7086 (N_7086,N_5040,N_4499);
or U7087 (N_7087,N_4871,N_5394);
nand U7088 (N_7088,N_5306,N_4150);
nor U7089 (N_7089,N_4301,N_4019);
nand U7090 (N_7090,N_5305,N_5177);
and U7091 (N_7091,N_4514,N_4040);
nor U7092 (N_7092,N_4060,N_4892);
and U7093 (N_7093,N_4165,N_5061);
or U7094 (N_7094,N_5953,N_4244);
nor U7095 (N_7095,N_4988,N_5935);
or U7096 (N_7096,N_4725,N_4826);
nor U7097 (N_7097,N_4702,N_5737);
nand U7098 (N_7098,N_5163,N_5517);
and U7099 (N_7099,N_4736,N_4435);
nor U7100 (N_7100,N_5208,N_4352);
or U7101 (N_7101,N_5089,N_5021);
or U7102 (N_7102,N_5206,N_5934);
and U7103 (N_7103,N_4540,N_4007);
and U7104 (N_7104,N_5299,N_5239);
or U7105 (N_7105,N_5686,N_5300);
or U7106 (N_7106,N_4704,N_4189);
nand U7107 (N_7107,N_5480,N_4184);
nand U7108 (N_7108,N_4558,N_4632);
and U7109 (N_7109,N_4763,N_5283);
and U7110 (N_7110,N_5424,N_4710);
nor U7111 (N_7111,N_5841,N_5612);
or U7112 (N_7112,N_5332,N_4792);
nor U7113 (N_7113,N_4043,N_5995);
and U7114 (N_7114,N_4291,N_5692);
nor U7115 (N_7115,N_5213,N_4520);
or U7116 (N_7116,N_4056,N_4995);
or U7117 (N_7117,N_5784,N_4966);
nand U7118 (N_7118,N_5191,N_4153);
and U7119 (N_7119,N_4972,N_4845);
nor U7120 (N_7120,N_4214,N_5623);
or U7121 (N_7121,N_5851,N_5148);
and U7122 (N_7122,N_5506,N_5683);
or U7123 (N_7123,N_4349,N_4228);
and U7124 (N_7124,N_4656,N_4842);
nand U7125 (N_7125,N_4528,N_5765);
and U7126 (N_7126,N_4841,N_5152);
and U7127 (N_7127,N_4795,N_4736);
nand U7128 (N_7128,N_4350,N_5618);
and U7129 (N_7129,N_5109,N_4932);
nand U7130 (N_7130,N_5175,N_4614);
or U7131 (N_7131,N_5202,N_5014);
nand U7132 (N_7132,N_5487,N_4148);
nor U7133 (N_7133,N_4769,N_4790);
nor U7134 (N_7134,N_4401,N_4510);
nand U7135 (N_7135,N_5795,N_4103);
or U7136 (N_7136,N_5506,N_5304);
or U7137 (N_7137,N_5513,N_4149);
and U7138 (N_7138,N_4484,N_4244);
nor U7139 (N_7139,N_5773,N_4942);
and U7140 (N_7140,N_5902,N_4635);
and U7141 (N_7141,N_4747,N_4682);
and U7142 (N_7142,N_5932,N_4951);
nand U7143 (N_7143,N_5760,N_4531);
and U7144 (N_7144,N_4812,N_5766);
nor U7145 (N_7145,N_4066,N_5959);
and U7146 (N_7146,N_5549,N_5531);
and U7147 (N_7147,N_4226,N_5549);
nor U7148 (N_7148,N_5246,N_5952);
nor U7149 (N_7149,N_5578,N_5601);
or U7150 (N_7150,N_5782,N_4320);
nand U7151 (N_7151,N_4270,N_5581);
nand U7152 (N_7152,N_5523,N_4953);
and U7153 (N_7153,N_4561,N_5309);
and U7154 (N_7154,N_4649,N_4697);
nand U7155 (N_7155,N_5401,N_4917);
nand U7156 (N_7156,N_4943,N_5152);
nor U7157 (N_7157,N_5031,N_4183);
and U7158 (N_7158,N_5663,N_4600);
and U7159 (N_7159,N_4504,N_4571);
and U7160 (N_7160,N_5218,N_4854);
nor U7161 (N_7161,N_5079,N_4486);
nor U7162 (N_7162,N_4727,N_5747);
nor U7163 (N_7163,N_4071,N_5780);
nor U7164 (N_7164,N_5174,N_4880);
nand U7165 (N_7165,N_4864,N_5089);
and U7166 (N_7166,N_4830,N_5074);
nor U7167 (N_7167,N_5925,N_4100);
or U7168 (N_7168,N_4853,N_4490);
and U7169 (N_7169,N_4589,N_5260);
and U7170 (N_7170,N_4421,N_4574);
or U7171 (N_7171,N_4152,N_5954);
nand U7172 (N_7172,N_5319,N_5384);
and U7173 (N_7173,N_5976,N_5912);
and U7174 (N_7174,N_4261,N_5418);
nor U7175 (N_7175,N_4737,N_5892);
or U7176 (N_7176,N_4510,N_5710);
or U7177 (N_7177,N_5134,N_4078);
or U7178 (N_7178,N_5868,N_5274);
or U7179 (N_7179,N_5192,N_5217);
and U7180 (N_7180,N_4773,N_4042);
or U7181 (N_7181,N_4592,N_4419);
nand U7182 (N_7182,N_4996,N_4135);
and U7183 (N_7183,N_4303,N_4815);
nor U7184 (N_7184,N_5272,N_4766);
nor U7185 (N_7185,N_5539,N_4398);
or U7186 (N_7186,N_4673,N_4491);
or U7187 (N_7187,N_5026,N_5765);
and U7188 (N_7188,N_4433,N_4752);
nor U7189 (N_7189,N_5352,N_4973);
or U7190 (N_7190,N_5912,N_4140);
nor U7191 (N_7191,N_5971,N_5948);
or U7192 (N_7192,N_5758,N_4488);
or U7193 (N_7193,N_5384,N_4968);
or U7194 (N_7194,N_4820,N_5144);
or U7195 (N_7195,N_4291,N_4636);
and U7196 (N_7196,N_5972,N_4955);
nor U7197 (N_7197,N_4419,N_5259);
xor U7198 (N_7198,N_5018,N_4304);
and U7199 (N_7199,N_4997,N_5795);
nor U7200 (N_7200,N_4831,N_5159);
and U7201 (N_7201,N_5613,N_4550);
or U7202 (N_7202,N_4472,N_4696);
nor U7203 (N_7203,N_5949,N_5056);
and U7204 (N_7204,N_4500,N_4394);
nand U7205 (N_7205,N_5040,N_4787);
nand U7206 (N_7206,N_5175,N_4321);
nor U7207 (N_7207,N_4630,N_4365);
and U7208 (N_7208,N_4572,N_4876);
nand U7209 (N_7209,N_5001,N_4707);
and U7210 (N_7210,N_4649,N_5510);
and U7211 (N_7211,N_4842,N_4249);
xor U7212 (N_7212,N_4096,N_4300);
nand U7213 (N_7213,N_4514,N_4635);
nand U7214 (N_7214,N_4743,N_5977);
nand U7215 (N_7215,N_5071,N_5273);
nand U7216 (N_7216,N_5040,N_5831);
nor U7217 (N_7217,N_4695,N_5659);
nor U7218 (N_7218,N_4654,N_4258);
nor U7219 (N_7219,N_4288,N_4268);
nor U7220 (N_7220,N_5330,N_4013);
nand U7221 (N_7221,N_5294,N_4468);
and U7222 (N_7222,N_4377,N_4738);
nand U7223 (N_7223,N_4544,N_5009);
nor U7224 (N_7224,N_5764,N_4724);
nor U7225 (N_7225,N_5749,N_5146);
and U7226 (N_7226,N_5095,N_5472);
or U7227 (N_7227,N_5420,N_5672);
and U7228 (N_7228,N_4294,N_5375);
nand U7229 (N_7229,N_5399,N_5904);
and U7230 (N_7230,N_5669,N_5840);
nand U7231 (N_7231,N_5809,N_4277);
and U7232 (N_7232,N_4843,N_5092);
nand U7233 (N_7233,N_5556,N_5324);
nor U7234 (N_7234,N_5274,N_5581);
nor U7235 (N_7235,N_4142,N_5727);
nor U7236 (N_7236,N_5170,N_5339);
nor U7237 (N_7237,N_4272,N_4530);
nor U7238 (N_7238,N_4908,N_4280);
or U7239 (N_7239,N_4578,N_4570);
and U7240 (N_7240,N_5481,N_4331);
nand U7241 (N_7241,N_4869,N_5714);
or U7242 (N_7242,N_5132,N_4526);
or U7243 (N_7243,N_4632,N_4694);
and U7244 (N_7244,N_5848,N_4622);
nor U7245 (N_7245,N_5320,N_4289);
nor U7246 (N_7246,N_4051,N_4806);
and U7247 (N_7247,N_4606,N_4289);
and U7248 (N_7248,N_4231,N_4948);
and U7249 (N_7249,N_5788,N_5345);
nand U7250 (N_7250,N_4422,N_5158);
nor U7251 (N_7251,N_5680,N_5309);
nor U7252 (N_7252,N_5929,N_5997);
or U7253 (N_7253,N_4936,N_4274);
and U7254 (N_7254,N_5227,N_5694);
nor U7255 (N_7255,N_5699,N_4227);
nor U7256 (N_7256,N_5085,N_5363);
and U7257 (N_7257,N_4359,N_5414);
and U7258 (N_7258,N_5295,N_4226);
nor U7259 (N_7259,N_5673,N_5026);
and U7260 (N_7260,N_5018,N_4794);
and U7261 (N_7261,N_5795,N_4632);
nand U7262 (N_7262,N_5398,N_5152);
nand U7263 (N_7263,N_4593,N_4033);
nor U7264 (N_7264,N_5307,N_5002);
nand U7265 (N_7265,N_4238,N_5887);
and U7266 (N_7266,N_5760,N_5597);
and U7267 (N_7267,N_5756,N_4583);
nor U7268 (N_7268,N_5892,N_5572);
nor U7269 (N_7269,N_4139,N_5919);
nor U7270 (N_7270,N_4013,N_5988);
nor U7271 (N_7271,N_4008,N_4645);
nor U7272 (N_7272,N_5899,N_5800);
xnor U7273 (N_7273,N_4898,N_5904);
nand U7274 (N_7274,N_5421,N_4472);
or U7275 (N_7275,N_5264,N_4660);
and U7276 (N_7276,N_5107,N_4242);
or U7277 (N_7277,N_5045,N_4416);
nor U7278 (N_7278,N_5388,N_5949);
nand U7279 (N_7279,N_5489,N_4875);
nor U7280 (N_7280,N_4071,N_5737);
nor U7281 (N_7281,N_4518,N_4273);
and U7282 (N_7282,N_4562,N_4107);
and U7283 (N_7283,N_5960,N_4329);
and U7284 (N_7284,N_4487,N_4059);
nor U7285 (N_7285,N_4277,N_4356);
and U7286 (N_7286,N_5360,N_4621);
nand U7287 (N_7287,N_4708,N_4301);
and U7288 (N_7288,N_5798,N_5007);
nand U7289 (N_7289,N_5172,N_5728);
nor U7290 (N_7290,N_5747,N_4051);
and U7291 (N_7291,N_5748,N_4008);
and U7292 (N_7292,N_4878,N_4864);
and U7293 (N_7293,N_4447,N_4187);
nor U7294 (N_7294,N_4568,N_5293);
nor U7295 (N_7295,N_4783,N_5844);
or U7296 (N_7296,N_5979,N_4346);
or U7297 (N_7297,N_4403,N_5061);
and U7298 (N_7298,N_5975,N_4827);
nor U7299 (N_7299,N_4873,N_4334);
nand U7300 (N_7300,N_4998,N_4790);
and U7301 (N_7301,N_4943,N_5384);
or U7302 (N_7302,N_4699,N_4883);
and U7303 (N_7303,N_4433,N_4858);
nand U7304 (N_7304,N_4683,N_4602);
and U7305 (N_7305,N_4968,N_5772);
xor U7306 (N_7306,N_4290,N_4380);
and U7307 (N_7307,N_4054,N_4139);
nand U7308 (N_7308,N_4310,N_4254);
or U7309 (N_7309,N_5700,N_4961);
xnor U7310 (N_7310,N_5888,N_4128);
nor U7311 (N_7311,N_4128,N_4722);
and U7312 (N_7312,N_5751,N_4623);
and U7313 (N_7313,N_4770,N_4885);
and U7314 (N_7314,N_5571,N_5454);
nor U7315 (N_7315,N_4382,N_5272);
or U7316 (N_7316,N_5003,N_4291);
and U7317 (N_7317,N_5242,N_4937);
and U7318 (N_7318,N_5576,N_4441);
or U7319 (N_7319,N_5085,N_5358);
nor U7320 (N_7320,N_4498,N_4111);
and U7321 (N_7321,N_5926,N_5917);
and U7322 (N_7322,N_5323,N_4315);
or U7323 (N_7323,N_5898,N_5295);
or U7324 (N_7324,N_5942,N_4240);
nor U7325 (N_7325,N_5879,N_5381);
and U7326 (N_7326,N_4258,N_4440);
and U7327 (N_7327,N_5710,N_5293);
nor U7328 (N_7328,N_4954,N_5929);
nand U7329 (N_7329,N_5085,N_5619);
nor U7330 (N_7330,N_5010,N_4717);
nor U7331 (N_7331,N_4081,N_5235);
or U7332 (N_7332,N_4137,N_5507);
and U7333 (N_7333,N_5054,N_5595);
or U7334 (N_7334,N_5627,N_4529);
or U7335 (N_7335,N_4076,N_5855);
nand U7336 (N_7336,N_5048,N_4740);
or U7337 (N_7337,N_4784,N_4864);
or U7338 (N_7338,N_4313,N_4432);
nor U7339 (N_7339,N_4697,N_4321);
or U7340 (N_7340,N_4345,N_5126);
nor U7341 (N_7341,N_4344,N_4043);
and U7342 (N_7342,N_4222,N_5550);
nor U7343 (N_7343,N_4466,N_5975);
and U7344 (N_7344,N_4910,N_5711);
or U7345 (N_7345,N_5915,N_4343);
nand U7346 (N_7346,N_4343,N_5872);
and U7347 (N_7347,N_4313,N_5123);
and U7348 (N_7348,N_5107,N_5292);
nor U7349 (N_7349,N_4555,N_4385);
nand U7350 (N_7350,N_4863,N_4183);
nand U7351 (N_7351,N_4074,N_4882);
nor U7352 (N_7352,N_5420,N_5916);
nor U7353 (N_7353,N_4075,N_4345);
nand U7354 (N_7354,N_5056,N_4045);
nor U7355 (N_7355,N_5071,N_5320);
and U7356 (N_7356,N_4495,N_4558);
nor U7357 (N_7357,N_4505,N_4474);
and U7358 (N_7358,N_5546,N_4783);
nand U7359 (N_7359,N_4262,N_4476);
nor U7360 (N_7360,N_4741,N_4770);
nand U7361 (N_7361,N_4374,N_5091);
and U7362 (N_7362,N_5673,N_4639);
nand U7363 (N_7363,N_5069,N_5654);
and U7364 (N_7364,N_5479,N_5466);
and U7365 (N_7365,N_4938,N_4120);
nor U7366 (N_7366,N_5675,N_5964);
nand U7367 (N_7367,N_4346,N_5063);
nor U7368 (N_7368,N_4256,N_5330);
and U7369 (N_7369,N_4425,N_4950);
nor U7370 (N_7370,N_4774,N_5931);
and U7371 (N_7371,N_4527,N_4326);
and U7372 (N_7372,N_5678,N_5091);
nor U7373 (N_7373,N_4101,N_4474);
nand U7374 (N_7374,N_4988,N_5841);
or U7375 (N_7375,N_4132,N_5928);
and U7376 (N_7376,N_4255,N_5498);
nor U7377 (N_7377,N_5240,N_4135);
or U7378 (N_7378,N_5263,N_5204);
and U7379 (N_7379,N_4553,N_4598);
nor U7380 (N_7380,N_5752,N_4058);
and U7381 (N_7381,N_4362,N_5849);
nand U7382 (N_7382,N_4819,N_4917);
and U7383 (N_7383,N_5031,N_5102);
or U7384 (N_7384,N_5221,N_4734);
or U7385 (N_7385,N_5947,N_5743);
or U7386 (N_7386,N_5535,N_4469);
nor U7387 (N_7387,N_4190,N_5550);
nand U7388 (N_7388,N_4394,N_4588);
nand U7389 (N_7389,N_5369,N_5252);
or U7390 (N_7390,N_5261,N_5216);
nor U7391 (N_7391,N_4158,N_5069);
and U7392 (N_7392,N_5917,N_5034);
nand U7393 (N_7393,N_5177,N_5852);
nor U7394 (N_7394,N_5820,N_4814);
or U7395 (N_7395,N_4780,N_4660);
and U7396 (N_7396,N_4265,N_4624);
nor U7397 (N_7397,N_4625,N_4473);
nor U7398 (N_7398,N_4574,N_5981);
and U7399 (N_7399,N_4376,N_4919);
and U7400 (N_7400,N_4397,N_5136);
or U7401 (N_7401,N_4446,N_5220);
nand U7402 (N_7402,N_5416,N_5261);
nand U7403 (N_7403,N_4204,N_4883);
or U7404 (N_7404,N_4788,N_5010);
and U7405 (N_7405,N_5866,N_5125);
nand U7406 (N_7406,N_4749,N_4096);
or U7407 (N_7407,N_4026,N_4380);
nand U7408 (N_7408,N_5797,N_5168);
or U7409 (N_7409,N_5586,N_4716);
or U7410 (N_7410,N_4906,N_4723);
or U7411 (N_7411,N_5561,N_5910);
nor U7412 (N_7412,N_5631,N_4515);
or U7413 (N_7413,N_4973,N_4537);
or U7414 (N_7414,N_4174,N_5539);
nand U7415 (N_7415,N_4665,N_4036);
nand U7416 (N_7416,N_5815,N_4461);
nor U7417 (N_7417,N_4413,N_4349);
nor U7418 (N_7418,N_4550,N_5919);
and U7419 (N_7419,N_4657,N_5725);
and U7420 (N_7420,N_5860,N_4901);
or U7421 (N_7421,N_5574,N_5800);
nor U7422 (N_7422,N_4000,N_4750);
and U7423 (N_7423,N_5639,N_4211);
or U7424 (N_7424,N_5475,N_4181);
or U7425 (N_7425,N_5183,N_4901);
nand U7426 (N_7426,N_5792,N_4902);
or U7427 (N_7427,N_4925,N_4969);
nand U7428 (N_7428,N_4689,N_5191);
nor U7429 (N_7429,N_5615,N_5286);
nor U7430 (N_7430,N_4434,N_5607);
and U7431 (N_7431,N_4170,N_4861);
nor U7432 (N_7432,N_5491,N_4332);
or U7433 (N_7433,N_5004,N_5862);
or U7434 (N_7434,N_4330,N_4290);
nor U7435 (N_7435,N_5144,N_5241);
nand U7436 (N_7436,N_4936,N_5349);
or U7437 (N_7437,N_4824,N_5200);
nor U7438 (N_7438,N_4691,N_4479);
or U7439 (N_7439,N_5034,N_5070);
nor U7440 (N_7440,N_4938,N_4203);
nand U7441 (N_7441,N_5593,N_5680);
nor U7442 (N_7442,N_5720,N_4743);
and U7443 (N_7443,N_4136,N_5896);
nand U7444 (N_7444,N_4704,N_4300);
and U7445 (N_7445,N_4470,N_5773);
or U7446 (N_7446,N_4978,N_5577);
and U7447 (N_7447,N_4794,N_4781);
and U7448 (N_7448,N_5484,N_5812);
nor U7449 (N_7449,N_5259,N_5518);
nor U7450 (N_7450,N_4612,N_4533);
nor U7451 (N_7451,N_4195,N_5523);
nand U7452 (N_7452,N_5019,N_5268);
or U7453 (N_7453,N_4796,N_4735);
nor U7454 (N_7454,N_4859,N_4431);
nand U7455 (N_7455,N_5255,N_5439);
xnor U7456 (N_7456,N_5264,N_4612);
or U7457 (N_7457,N_4935,N_5568);
nand U7458 (N_7458,N_4894,N_4512);
nand U7459 (N_7459,N_4408,N_4653);
and U7460 (N_7460,N_5321,N_5182);
nand U7461 (N_7461,N_4148,N_4210);
nand U7462 (N_7462,N_5760,N_5910);
nor U7463 (N_7463,N_5587,N_4956);
or U7464 (N_7464,N_5004,N_4481);
and U7465 (N_7465,N_4239,N_5270);
nand U7466 (N_7466,N_5267,N_5896);
or U7467 (N_7467,N_4287,N_4003);
nand U7468 (N_7468,N_5826,N_4106);
nand U7469 (N_7469,N_4676,N_5698);
or U7470 (N_7470,N_4409,N_4833);
and U7471 (N_7471,N_5219,N_5025);
and U7472 (N_7472,N_4249,N_4088);
and U7473 (N_7473,N_5080,N_4499);
or U7474 (N_7474,N_5535,N_5675);
nand U7475 (N_7475,N_5554,N_5307);
or U7476 (N_7476,N_4653,N_5113);
nand U7477 (N_7477,N_5866,N_4542);
or U7478 (N_7478,N_4362,N_4997);
and U7479 (N_7479,N_5491,N_4545);
and U7480 (N_7480,N_4389,N_5007);
and U7481 (N_7481,N_4800,N_5232);
or U7482 (N_7482,N_4842,N_4254);
or U7483 (N_7483,N_5300,N_4235);
nor U7484 (N_7484,N_4410,N_4181);
nand U7485 (N_7485,N_4502,N_5580);
and U7486 (N_7486,N_4527,N_4209);
or U7487 (N_7487,N_4599,N_4281);
or U7488 (N_7488,N_5350,N_5884);
nor U7489 (N_7489,N_5331,N_5094);
nand U7490 (N_7490,N_4022,N_5093);
nor U7491 (N_7491,N_4152,N_4942);
and U7492 (N_7492,N_5320,N_4905);
or U7493 (N_7493,N_4372,N_4395);
and U7494 (N_7494,N_5296,N_4281);
nor U7495 (N_7495,N_5295,N_4753);
or U7496 (N_7496,N_4427,N_5043);
nand U7497 (N_7497,N_4901,N_5636);
nor U7498 (N_7498,N_5124,N_4084);
and U7499 (N_7499,N_5550,N_4674);
nor U7500 (N_7500,N_5559,N_4806);
nor U7501 (N_7501,N_5373,N_4804);
and U7502 (N_7502,N_5242,N_5754);
nand U7503 (N_7503,N_5891,N_4579);
nor U7504 (N_7504,N_4472,N_5649);
nor U7505 (N_7505,N_5143,N_4130);
or U7506 (N_7506,N_4456,N_4655);
and U7507 (N_7507,N_4434,N_4191);
or U7508 (N_7508,N_5474,N_5603);
nand U7509 (N_7509,N_5211,N_4116);
and U7510 (N_7510,N_4764,N_4533);
nand U7511 (N_7511,N_5318,N_4917);
nor U7512 (N_7512,N_5493,N_4344);
nor U7513 (N_7513,N_5592,N_4844);
and U7514 (N_7514,N_4122,N_4395);
nand U7515 (N_7515,N_5846,N_4677);
nor U7516 (N_7516,N_5238,N_5449);
and U7517 (N_7517,N_5040,N_5399);
nor U7518 (N_7518,N_5431,N_4192);
and U7519 (N_7519,N_5323,N_5747);
and U7520 (N_7520,N_5502,N_5622);
nand U7521 (N_7521,N_4101,N_4365);
nand U7522 (N_7522,N_5030,N_5273);
nor U7523 (N_7523,N_5805,N_4972);
and U7524 (N_7524,N_5086,N_4004);
or U7525 (N_7525,N_4788,N_5870);
and U7526 (N_7526,N_5620,N_5221);
and U7527 (N_7527,N_5906,N_5660);
and U7528 (N_7528,N_4837,N_4166);
nand U7529 (N_7529,N_4192,N_5564);
and U7530 (N_7530,N_5413,N_4027);
or U7531 (N_7531,N_5999,N_5661);
nand U7532 (N_7532,N_4512,N_5060);
nand U7533 (N_7533,N_5143,N_5312);
nor U7534 (N_7534,N_5611,N_4351);
and U7535 (N_7535,N_4065,N_4988);
nor U7536 (N_7536,N_4294,N_4559);
nor U7537 (N_7537,N_5499,N_5282);
and U7538 (N_7538,N_4833,N_4858);
nor U7539 (N_7539,N_5393,N_4089);
nor U7540 (N_7540,N_4728,N_4441);
nor U7541 (N_7541,N_4629,N_5621);
nor U7542 (N_7542,N_4887,N_4691);
nand U7543 (N_7543,N_5554,N_5365);
and U7544 (N_7544,N_4583,N_4436);
nand U7545 (N_7545,N_5653,N_4711);
nand U7546 (N_7546,N_4561,N_4057);
and U7547 (N_7547,N_4902,N_4686);
nand U7548 (N_7548,N_5400,N_4426);
or U7549 (N_7549,N_4627,N_4092);
and U7550 (N_7550,N_5618,N_4009);
or U7551 (N_7551,N_4307,N_5328);
and U7552 (N_7552,N_4473,N_4918);
or U7553 (N_7553,N_5205,N_4638);
nor U7554 (N_7554,N_4222,N_4243);
nor U7555 (N_7555,N_4192,N_5797);
nand U7556 (N_7556,N_4210,N_5275);
nand U7557 (N_7557,N_4555,N_4898);
nor U7558 (N_7558,N_4564,N_4468);
or U7559 (N_7559,N_4516,N_4912);
and U7560 (N_7560,N_5517,N_5812);
nor U7561 (N_7561,N_5542,N_4974);
nand U7562 (N_7562,N_5973,N_5806);
and U7563 (N_7563,N_5074,N_5203);
nor U7564 (N_7564,N_5957,N_5900);
nand U7565 (N_7565,N_4910,N_4485);
nand U7566 (N_7566,N_4361,N_4881);
nor U7567 (N_7567,N_5367,N_4799);
or U7568 (N_7568,N_5883,N_4935);
or U7569 (N_7569,N_5034,N_5822);
nand U7570 (N_7570,N_5673,N_4340);
nor U7571 (N_7571,N_5193,N_4527);
nand U7572 (N_7572,N_4374,N_5429);
nand U7573 (N_7573,N_5623,N_5443);
nor U7574 (N_7574,N_4255,N_4903);
and U7575 (N_7575,N_4667,N_5864);
and U7576 (N_7576,N_4003,N_5561);
or U7577 (N_7577,N_4669,N_4309);
nand U7578 (N_7578,N_4819,N_5028);
nor U7579 (N_7579,N_5597,N_5337);
or U7580 (N_7580,N_4836,N_5334);
and U7581 (N_7581,N_5718,N_5546);
or U7582 (N_7582,N_5227,N_4698);
and U7583 (N_7583,N_5040,N_4963);
or U7584 (N_7584,N_4281,N_4847);
nand U7585 (N_7585,N_5996,N_4208);
or U7586 (N_7586,N_4670,N_5029);
nand U7587 (N_7587,N_5809,N_5978);
and U7588 (N_7588,N_5325,N_4484);
nand U7589 (N_7589,N_5765,N_4398);
nand U7590 (N_7590,N_4965,N_5455);
or U7591 (N_7591,N_4352,N_4856);
and U7592 (N_7592,N_5634,N_5482);
nor U7593 (N_7593,N_4221,N_4658);
and U7594 (N_7594,N_4504,N_5495);
nor U7595 (N_7595,N_5722,N_4922);
nand U7596 (N_7596,N_4640,N_5289);
nand U7597 (N_7597,N_5296,N_5223);
nand U7598 (N_7598,N_5589,N_5058);
nor U7599 (N_7599,N_5417,N_5546);
nand U7600 (N_7600,N_5748,N_4803);
xor U7601 (N_7601,N_4542,N_5388);
or U7602 (N_7602,N_4076,N_4566);
nand U7603 (N_7603,N_5872,N_5987);
or U7604 (N_7604,N_4546,N_4697);
or U7605 (N_7605,N_5661,N_5173);
and U7606 (N_7606,N_4770,N_4160);
or U7607 (N_7607,N_5908,N_5338);
and U7608 (N_7608,N_5921,N_4557);
or U7609 (N_7609,N_4613,N_4074);
or U7610 (N_7610,N_4714,N_5400);
or U7611 (N_7611,N_5896,N_4082);
and U7612 (N_7612,N_4651,N_4143);
or U7613 (N_7613,N_5445,N_4621);
and U7614 (N_7614,N_5358,N_4432);
or U7615 (N_7615,N_5094,N_4937);
and U7616 (N_7616,N_4949,N_4179);
nor U7617 (N_7617,N_5739,N_5660);
and U7618 (N_7618,N_5414,N_4593);
nor U7619 (N_7619,N_5368,N_4769);
and U7620 (N_7620,N_4925,N_5529);
or U7621 (N_7621,N_5375,N_5303);
or U7622 (N_7622,N_5528,N_4755);
and U7623 (N_7623,N_4954,N_4712);
nor U7624 (N_7624,N_5038,N_4180);
nor U7625 (N_7625,N_5695,N_5099);
nor U7626 (N_7626,N_5354,N_4540);
or U7627 (N_7627,N_4551,N_5224);
nor U7628 (N_7628,N_5557,N_4402);
nand U7629 (N_7629,N_5458,N_4245);
nand U7630 (N_7630,N_5145,N_4046);
nand U7631 (N_7631,N_4058,N_5760);
or U7632 (N_7632,N_5087,N_4805);
nor U7633 (N_7633,N_5600,N_4421);
nor U7634 (N_7634,N_4762,N_5137);
and U7635 (N_7635,N_4773,N_5966);
nor U7636 (N_7636,N_4706,N_4921);
xnor U7637 (N_7637,N_5042,N_5789);
nor U7638 (N_7638,N_4375,N_4784);
nand U7639 (N_7639,N_4858,N_5230);
or U7640 (N_7640,N_4608,N_4537);
nor U7641 (N_7641,N_4301,N_4119);
and U7642 (N_7642,N_4929,N_5361);
nor U7643 (N_7643,N_4705,N_5139);
nor U7644 (N_7644,N_5857,N_4010);
nor U7645 (N_7645,N_4923,N_5824);
nand U7646 (N_7646,N_4176,N_4009);
and U7647 (N_7647,N_5675,N_4438);
or U7648 (N_7648,N_5419,N_4966);
nand U7649 (N_7649,N_5803,N_5200);
nand U7650 (N_7650,N_5180,N_4616);
and U7651 (N_7651,N_4302,N_4564);
nand U7652 (N_7652,N_4518,N_5276);
nor U7653 (N_7653,N_4901,N_5306);
nor U7654 (N_7654,N_5790,N_5379);
or U7655 (N_7655,N_5182,N_4037);
or U7656 (N_7656,N_5972,N_5722);
or U7657 (N_7657,N_5177,N_5436);
nand U7658 (N_7658,N_5354,N_5007);
or U7659 (N_7659,N_4194,N_5109);
nand U7660 (N_7660,N_5122,N_4984);
and U7661 (N_7661,N_4301,N_4103);
and U7662 (N_7662,N_5035,N_5839);
xnor U7663 (N_7663,N_5510,N_5318);
or U7664 (N_7664,N_5992,N_4611);
nand U7665 (N_7665,N_5764,N_4173);
and U7666 (N_7666,N_5890,N_4059);
or U7667 (N_7667,N_5964,N_4359);
or U7668 (N_7668,N_4539,N_5611);
nor U7669 (N_7669,N_4011,N_5609);
nand U7670 (N_7670,N_4652,N_4796);
nand U7671 (N_7671,N_4532,N_4891);
nor U7672 (N_7672,N_5337,N_4641);
or U7673 (N_7673,N_4539,N_4477);
nand U7674 (N_7674,N_5897,N_4964);
nand U7675 (N_7675,N_4277,N_4720);
xor U7676 (N_7676,N_4937,N_5216);
or U7677 (N_7677,N_4545,N_5090);
nand U7678 (N_7678,N_5103,N_4603);
nand U7679 (N_7679,N_5698,N_5730);
nand U7680 (N_7680,N_4500,N_5227);
and U7681 (N_7681,N_4534,N_5222);
and U7682 (N_7682,N_4079,N_5134);
nor U7683 (N_7683,N_5890,N_4573);
or U7684 (N_7684,N_4986,N_5781);
and U7685 (N_7685,N_5274,N_4397);
nor U7686 (N_7686,N_4159,N_4412);
nor U7687 (N_7687,N_5784,N_4700);
nor U7688 (N_7688,N_4646,N_5784);
nand U7689 (N_7689,N_4516,N_5730);
nor U7690 (N_7690,N_4245,N_4035);
or U7691 (N_7691,N_5063,N_5949);
nor U7692 (N_7692,N_5301,N_4188);
nand U7693 (N_7693,N_5510,N_5322);
nor U7694 (N_7694,N_5405,N_5752);
nand U7695 (N_7695,N_4385,N_5318);
or U7696 (N_7696,N_5416,N_5338);
nor U7697 (N_7697,N_4388,N_4789);
and U7698 (N_7698,N_4553,N_5581);
or U7699 (N_7699,N_5190,N_5133);
nand U7700 (N_7700,N_5033,N_4653);
nand U7701 (N_7701,N_5795,N_5393);
nor U7702 (N_7702,N_5741,N_5426);
nand U7703 (N_7703,N_4027,N_5288);
and U7704 (N_7704,N_4591,N_4960);
and U7705 (N_7705,N_5306,N_4228);
nor U7706 (N_7706,N_4631,N_4823);
nor U7707 (N_7707,N_4151,N_4656);
and U7708 (N_7708,N_4603,N_5891);
and U7709 (N_7709,N_4623,N_5359);
nor U7710 (N_7710,N_4175,N_4671);
nand U7711 (N_7711,N_5123,N_5543);
or U7712 (N_7712,N_5547,N_4475);
or U7713 (N_7713,N_4490,N_4092);
nor U7714 (N_7714,N_5666,N_4767);
nor U7715 (N_7715,N_5759,N_5516);
or U7716 (N_7716,N_5515,N_4107);
nand U7717 (N_7717,N_5123,N_5898);
nor U7718 (N_7718,N_4429,N_5390);
xor U7719 (N_7719,N_4988,N_5326);
or U7720 (N_7720,N_4357,N_4441);
or U7721 (N_7721,N_5864,N_5802);
or U7722 (N_7722,N_4440,N_4804);
nor U7723 (N_7723,N_5078,N_4082);
or U7724 (N_7724,N_5885,N_5577);
nor U7725 (N_7725,N_4667,N_4901);
and U7726 (N_7726,N_5465,N_5107);
nand U7727 (N_7727,N_5711,N_4979);
and U7728 (N_7728,N_4230,N_5548);
nand U7729 (N_7729,N_5538,N_4427);
nor U7730 (N_7730,N_5293,N_4165);
nand U7731 (N_7731,N_5310,N_4312);
and U7732 (N_7732,N_5540,N_5056);
nor U7733 (N_7733,N_4470,N_5729);
and U7734 (N_7734,N_5756,N_5453);
and U7735 (N_7735,N_5698,N_5872);
and U7736 (N_7736,N_5362,N_5835);
or U7737 (N_7737,N_5341,N_4173);
nand U7738 (N_7738,N_4522,N_4177);
and U7739 (N_7739,N_4590,N_5712);
nand U7740 (N_7740,N_4177,N_4894);
nor U7741 (N_7741,N_4598,N_5570);
nor U7742 (N_7742,N_4749,N_5674);
nor U7743 (N_7743,N_5121,N_4661);
nand U7744 (N_7744,N_5783,N_4191);
nor U7745 (N_7745,N_4259,N_4984);
or U7746 (N_7746,N_4316,N_4171);
nand U7747 (N_7747,N_4302,N_5974);
and U7748 (N_7748,N_4606,N_4625);
and U7749 (N_7749,N_5163,N_4877);
nand U7750 (N_7750,N_4858,N_4172);
and U7751 (N_7751,N_5202,N_5035);
and U7752 (N_7752,N_5616,N_5700);
nand U7753 (N_7753,N_5558,N_5199);
nor U7754 (N_7754,N_5292,N_5350);
and U7755 (N_7755,N_4940,N_5517);
or U7756 (N_7756,N_5079,N_5582);
nor U7757 (N_7757,N_5194,N_5485);
nand U7758 (N_7758,N_4036,N_4369);
or U7759 (N_7759,N_5986,N_5588);
nand U7760 (N_7760,N_5141,N_4502);
and U7761 (N_7761,N_4302,N_4442);
xor U7762 (N_7762,N_5950,N_4425);
or U7763 (N_7763,N_4643,N_5427);
nor U7764 (N_7764,N_5555,N_4009);
nor U7765 (N_7765,N_5519,N_5260);
and U7766 (N_7766,N_4052,N_5219);
and U7767 (N_7767,N_5427,N_5682);
or U7768 (N_7768,N_5878,N_5449);
xor U7769 (N_7769,N_5731,N_4164);
nand U7770 (N_7770,N_4144,N_4071);
nor U7771 (N_7771,N_4912,N_4140);
nor U7772 (N_7772,N_5141,N_5925);
nor U7773 (N_7773,N_4957,N_5261);
nor U7774 (N_7774,N_5002,N_5733);
nand U7775 (N_7775,N_5876,N_5689);
and U7776 (N_7776,N_4604,N_5233);
and U7777 (N_7777,N_4663,N_5033);
nor U7778 (N_7778,N_4412,N_5857);
and U7779 (N_7779,N_4520,N_5792);
or U7780 (N_7780,N_5986,N_4917);
and U7781 (N_7781,N_5979,N_4653);
and U7782 (N_7782,N_4487,N_5931);
and U7783 (N_7783,N_5380,N_5523);
nand U7784 (N_7784,N_5267,N_4170);
nand U7785 (N_7785,N_4161,N_5922);
or U7786 (N_7786,N_5281,N_5787);
nor U7787 (N_7787,N_5832,N_4274);
and U7788 (N_7788,N_4669,N_4736);
and U7789 (N_7789,N_4219,N_4595);
nor U7790 (N_7790,N_5159,N_4642);
or U7791 (N_7791,N_5634,N_4003);
nand U7792 (N_7792,N_4394,N_4396);
and U7793 (N_7793,N_4396,N_5932);
nand U7794 (N_7794,N_4869,N_5550);
nand U7795 (N_7795,N_5296,N_5084);
nor U7796 (N_7796,N_5729,N_4248);
xor U7797 (N_7797,N_5184,N_5220);
and U7798 (N_7798,N_5491,N_4937);
nor U7799 (N_7799,N_4309,N_5681);
nand U7800 (N_7800,N_4882,N_4858);
nand U7801 (N_7801,N_5975,N_4983);
and U7802 (N_7802,N_4026,N_4594);
or U7803 (N_7803,N_4979,N_5584);
and U7804 (N_7804,N_4872,N_5105);
or U7805 (N_7805,N_4118,N_4082);
and U7806 (N_7806,N_4444,N_5304);
nor U7807 (N_7807,N_5398,N_5661);
or U7808 (N_7808,N_5207,N_4551);
xor U7809 (N_7809,N_4191,N_4674);
or U7810 (N_7810,N_4704,N_5272);
nand U7811 (N_7811,N_4037,N_4005);
nor U7812 (N_7812,N_4251,N_5169);
nand U7813 (N_7813,N_5388,N_4667);
and U7814 (N_7814,N_4448,N_5857);
or U7815 (N_7815,N_4893,N_4414);
nor U7816 (N_7816,N_5571,N_5352);
nand U7817 (N_7817,N_5947,N_5150);
or U7818 (N_7818,N_5928,N_4092);
nand U7819 (N_7819,N_4293,N_4174);
or U7820 (N_7820,N_4605,N_4842);
nand U7821 (N_7821,N_4482,N_4673);
nand U7822 (N_7822,N_5473,N_4030);
and U7823 (N_7823,N_5833,N_5402);
or U7824 (N_7824,N_4735,N_4178);
or U7825 (N_7825,N_4791,N_4100);
nand U7826 (N_7826,N_5511,N_5557);
or U7827 (N_7827,N_5085,N_4545);
and U7828 (N_7828,N_5091,N_5191);
nor U7829 (N_7829,N_4960,N_5370);
and U7830 (N_7830,N_5120,N_5876);
nand U7831 (N_7831,N_5443,N_5021);
or U7832 (N_7832,N_5162,N_5934);
xnor U7833 (N_7833,N_4104,N_4291);
or U7834 (N_7834,N_5234,N_5625);
nor U7835 (N_7835,N_5371,N_5823);
or U7836 (N_7836,N_4492,N_5962);
nor U7837 (N_7837,N_5399,N_5135);
or U7838 (N_7838,N_5310,N_5802);
or U7839 (N_7839,N_4841,N_4304);
nand U7840 (N_7840,N_4286,N_5108);
or U7841 (N_7841,N_4638,N_5199);
nand U7842 (N_7842,N_5311,N_4825);
nor U7843 (N_7843,N_4256,N_5097);
and U7844 (N_7844,N_5747,N_4913);
and U7845 (N_7845,N_5495,N_4181);
nor U7846 (N_7846,N_5300,N_4961);
nand U7847 (N_7847,N_4885,N_4107);
nor U7848 (N_7848,N_5211,N_4919);
and U7849 (N_7849,N_5220,N_5237);
and U7850 (N_7850,N_5127,N_5312);
nand U7851 (N_7851,N_5080,N_5811);
nor U7852 (N_7852,N_4567,N_4316);
nand U7853 (N_7853,N_5980,N_5499);
and U7854 (N_7854,N_5960,N_5882);
or U7855 (N_7855,N_5702,N_4744);
and U7856 (N_7856,N_5964,N_4986);
and U7857 (N_7857,N_5764,N_4540);
and U7858 (N_7858,N_4864,N_4058);
nor U7859 (N_7859,N_5323,N_5529);
nand U7860 (N_7860,N_4149,N_5206);
and U7861 (N_7861,N_4336,N_4486);
nand U7862 (N_7862,N_4566,N_5211);
nand U7863 (N_7863,N_4733,N_4218);
and U7864 (N_7864,N_4341,N_4277);
nand U7865 (N_7865,N_5869,N_5782);
or U7866 (N_7866,N_5353,N_4114);
nor U7867 (N_7867,N_5182,N_5100);
and U7868 (N_7868,N_4582,N_4238);
or U7869 (N_7869,N_4050,N_5217);
or U7870 (N_7870,N_5552,N_4643);
or U7871 (N_7871,N_4899,N_5214);
nand U7872 (N_7872,N_4500,N_5173);
or U7873 (N_7873,N_5314,N_5002);
nor U7874 (N_7874,N_4263,N_5329);
nand U7875 (N_7875,N_5460,N_4674);
nand U7876 (N_7876,N_4546,N_5389);
and U7877 (N_7877,N_5393,N_4355);
and U7878 (N_7878,N_5593,N_4312);
nand U7879 (N_7879,N_4744,N_4112);
nand U7880 (N_7880,N_4927,N_5820);
and U7881 (N_7881,N_5127,N_4953);
nand U7882 (N_7882,N_5488,N_5707);
or U7883 (N_7883,N_5547,N_5182);
or U7884 (N_7884,N_5430,N_4046);
nand U7885 (N_7885,N_4057,N_4722);
nand U7886 (N_7886,N_4457,N_4662);
nor U7887 (N_7887,N_5385,N_4865);
and U7888 (N_7888,N_4485,N_5816);
nand U7889 (N_7889,N_5458,N_5571);
and U7890 (N_7890,N_4926,N_5835);
and U7891 (N_7891,N_4931,N_4073);
nor U7892 (N_7892,N_4260,N_5933);
and U7893 (N_7893,N_4226,N_5173);
nor U7894 (N_7894,N_4309,N_5102);
or U7895 (N_7895,N_5635,N_4508);
or U7896 (N_7896,N_4330,N_5356);
nor U7897 (N_7897,N_5151,N_5183);
nor U7898 (N_7898,N_5368,N_5041);
nor U7899 (N_7899,N_4670,N_4767);
nand U7900 (N_7900,N_5833,N_4892);
nor U7901 (N_7901,N_5813,N_4939);
nor U7902 (N_7902,N_5731,N_5635);
or U7903 (N_7903,N_4770,N_5913);
nor U7904 (N_7904,N_5709,N_5463);
and U7905 (N_7905,N_5171,N_4363);
nor U7906 (N_7906,N_5559,N_5768);
nor U7907 (N_7907,N_4281,N_4952);
or U7908 (N_7908,N_5929,N_5809);
nand U7909 (N_7909,N_4198,N_4163);
nand U7910 (N_7910,N_5880,N_5272);
nor U7911 (N_7911,N_4713,N_5122);
nand U7912 (N_7912,N_5671,N_5998);
and U7913 (N_7913,N_4407,N_4842);
nand U7914 (N_7914,N_4974,N_5952);
nor U7915 (N_7915,N_5981,N_4502);
or U7916 (N_7916,N_5033,N_4361);
nand U7917 (N_7917,N_4332,N_5949);
nor U7918 (N_7918,N_4345,N_4317);
nand U7919 (N_7919,N_4165,N_4219);
nand U7920 (N_7920,N_4400,N_4532);
nor U7921 (N_7921,N_5790,N_4398);
nand U7922 (N_7922,N_4550,N_5847);
or U7923 (N_7923,N_5155,N_5059);
or U7924 (N_7924,N_5395,N_4653);
nor U7925 (N_7925,N_4588,N_4277);
and U7926 (N_7926,N_4365,N_4392);
or U7927 (N_7927,N_5655,N_5145);
and U7928 (N_7928,N_5105,N_4519);
and U7929 (N_7929,N_5946,N_5959);
nor U7930 (N_7930,N_4992,N_5622);
and U7931 (N_7931,N_5763,N_5691);
or U7932 (N_7932,N_5210,N_5025);
or U7933 (N_7933,N_4030,N_5798);
and U7934 (N_7934,N_5251,N_4818);
nor U7935 (N_7935,N_4813,N_5362);
nor U7936 (N_7936,N_4066,N_4062);
or U7937 (N_7937,N_5800,N_4922);
nor U7938 (N_7938,N_4547,N_4936);
or U7939 (N_7939,N_5179,N_4507);
nand U7940 (N_7940,N_4461,N_4536);
or U7941 (N_7941,N_5696,N_5937);
or U7942 (N_7942,N_4749,N_5068);
or U7943 (N_7943,N_5345,N_5292);
nand U7944 (N_7944,N_5657,N_5039);
or U7945 (N_7945,N_5465,N_5568);
nand U7946 (N_7946,N_5548,N_4169);
or U7947 (N_7947,N_4796,N_4723);
nor U7948 (N_7948,N_4545,N_5852);
and U7949 (N_7949,N_5689,N_4330);
or U7950 (N_7950,N_5404,N_4078);
nor U7951 (N_7951,N_4472,N_5317);
nor U7952 (N_7952,N_5502,N_5119);
or U7953 (N_7953,N_5760,N_5445);
or U7954 (N_7954,N_4328,N_5581);
nor U7955 (N_7955,N_4176,N_4161);
and U7956 (N_7956,N_4422,N_5337);
xor U7957 (N_7957,N_5385,N_4603);
nor U7958 (N_7958,N_4949,N_5959);
nand U7959 (N_7959,N_5498,N_5934);
nor U7960 (N_7960,N_5555,N_4683);
nor U7961 (N_7961,N_5355,N_5412);
and U7962 (N_7962,N_5894,N_5347);
or U7963 (N_7963,N_4947,N_5163);
and U7964 (N_7964,N_4313,N_4434);
nor U7965 (N_7965,N_5695,N_5984);
nand U7966 (N_7966,N_4378,N_5411);
or U7967 (N_7967,N_5557,N_4415);
nand U7968 (N_7968,N_5011,N_5338);
nand U7969 (N_7969,N_5150,N_4265);
nor U7970 (N_7970,N_4231,N_4802);
and U7971 (N_7971,N_4829,N_5128);
nor U7972 (N_7972,N_4805,N_5567);
nand U7973 (N_7973,N_5060,N_5746);
nor U7974 (N_7974,N_5266,N_4378);
nor U7975 (N_7975,N_4592,N_5302);
and U7976 (N_7976,N_4049,N_4358);
and U7977 (N_7977,N_4704,N_4167);
nor U7978 (N_7978,N_5146,N_5177);
nand U7979 (N_7979,N_5829,N_4053);
nand U7980 (N_7980,N_5976,N_4012);
nand U7981 (N_7981,N_5854,N_5702);
nand U7982 (N_7982,N_5022,N_4283);
nand U7983 (N_7983,N_5995,N_4667);
nand U7984 (N_7984,N_4815,N_5057);
nand U7985 (N_7985,N_5457,N_4481);
and U7986 (N_7986,N_5465,N_4546);
or U7987 (N_7987,N_4353,N_4377);
nor U7988 (N_7988,N_5579,N_4996);
nand U7989 (N_7989,N_4921,N_4801);
nand U7990 (N_7990,N_5853,N_5320);
nor U7991 (N_7991,N_5129,N_5036);
or U7992 (N_7992,N_5687,N_4566);
and U7993 (N_7993,N_5904,N_5130);
xnor U7994 (N_7994,N_4027,N_4696);
nor U7995 (N_7995,N_5687,N_5352);
or U7996 (N_7996,N_4539,N_4401);
nand U7997 (N_7997,N_5575,N_4633);
or U7998 (N_7998,N_5608,N_4303);
nand U7999 (N_7999,N_5817,N_4501);
or U8000 (N_8000,N_7891,N_7388);
and U8001 (N_8001,N_6227,N_6944);
or U8002 (N_8002,N_7214,N_6546);
nand U8003 (N_8003,N_7673,N_6143);
or U8004 (N_8004,N_7333,N_6484);
or U8005 (N_8005,N_6213,N_6324);
and U8006 (N_8006,N_7749,N_6666);
or U8007 (N_8007,N_6351,N_6783);
or U8008 (N_8008,N_7703,N_7476);
nor U8009 (N_8009,N_7776,N_7087);
and U8010 (N_8010,N_6295,N_7288);
and U8011 (N_8011,N_7147,N_6681);
nand U8012 (N_8012,N_6799,N_6385);
nor U8013 (N_8013,N_6990,N_7195);
nor U8014 (N_8014,N_7565,N_6617);
and U8015 (N_8015,N_7132,N_6129);
and U8016 (N_8016,N_6564,N_6019);
nor U8017 (N_8017,N_6474,N_6517);
or U8018 (N_8018,N_7734,N_7173);
nor U8019 (N_8019,N_7268,N_7468);
nand U8020 (N_8020,N_6195,N_7904);
and U8021 (N_8021,N_7228,N_6752);
and U8022 (N_8022,N_6225,N_6728);
nor U8023 (N_8023,N_6076,N_7366);
and U8024 (N_8024,N_6429,N_7786);
nand U8025 (N_8025,N_7047,N_7923);
and U8026 (N_8026,N_7907,N_7062);
nor U8027 (N_8027,N_7315,N_7737);
and U8028 (N_8028,N_6203,N_7984);
and U8029 (N_8029,N_6999,N_6470);
xor U8030 (N_8030,N_7157,N_6138);
and U8031 (N_8031,N_7005,N_7819);
nor U8032 (N_8032,N_6508,N_7112);
nor U8033 (N_8033,N_6568,N_6284);
nor U8034 (N_8034,N_6023,N_7068);
and U8035 (N_8035,N_6430,N_6722);
or U8036 (N_8036,N_6081,N_6342);
or U8037 (N_8037,N_7630,N_7202);
and U8038 (N_8038,N_6184,N_7402);
nand U8039 (N_8039,N_7219,N_7508);
and U8040 (N_8040,N_6476,N_6045);
and U8041 (N_8041,N_6208,N_7263);
and U8042 (N_8042,N_6473,N_6460);
nor U8043 (N_8043,N_6620,N_6742);
or U8044 (N_8044,N_6587,N_7486);
nand U8045 (N_8045,N_6632,N_7296);
nor U8046 (N_8046,N_7572,N_7139);
and U8047 (N_8047,N_6581,N_6247);
nand U8048 (N_8048,N_6610,N_7148);
nand U8049 (N_8049,N_7206,N_6601);
and U8050 (N_8050,N_7729,N_6072);
nor U8051 (N_8051,N_6827,N_7085);
or U8052 (N_8052,N_6882,N_7986);
nor U8053 (N_8053,N_6588,N_6891);
or U8054 (N_8054,N_7006,N_7467);
nor U8055 (N_8055,N_6008,N_7599);
nor U8056 (N_8056,N_7817,N_6472);
and U8057 (N_8057,N_6895,N_7763);
or U8058 (N_8058,N_6776,N_7616);
or U8059 (N_8059,N_7016,N_6679);
nor U8060 (N_8060,N_7118,N_7973);
nor U8061 (N_8061,N_7646,N_7213);
nand U8062 (N_8062,N_6044,N_7444);
or U8063 (N_8063,N_6572,N_6505);
and U8064 (N_8064,N_6626,N_7610);
nor U8065 (N_8065,N_7951,N_6277);
nand U8066 (N_8066,N_7620,N_7253);
and U8067 (N_8067,N_6786,N_6466);
and U8068 (N_8068,N_7832,N_6443);
nand U8069 (N_8069,N_6793,N_7879);
nand U8070 (N_8070,N_7298,N_7856);
nor U8071 (N_8071,N_6604,N_7196);
and U8072 (N_8072,N_6199,N_7496);
and U8073 (N_8073,N_7245,N_7593);
and U8074 (N_8074,N_7474,N_7691);
nand U8075 (N_8075,N_6426,N_7320);
nor U8076 (N_8076,N_7696,N_6721);
or U8077 (N_8077,N_6964,N_7928);
and U8078 (N_8078,N_6532,N_7617);
nor U8079 (N_8079,N_7700,N_6688);
and U8080 (N_8080,N_7961,N_7479);
and U8081 (N_8081,N_6229,N_6988);
or U8082 (N_8082,N_6034,N_6654);
or U8083 (N_8083,N_6198,N_6383);
nand U8084 (N_8084,N_6265,N_7080);
or U8085 (N_8085,N_6984,N_6100);
nand U8086 (N_8086,N_6297,N_7101);
and U8087 (N_8087,N_7433,N_7520);
nor U8088 (N_8088,N_6362,N_6387);
nand U8089 (N_8089,N_7127,N_7732);
and U8090 (N_8090,N_6368,N_7241);
or U8091 (N_8091,N_7741,N_7609);
and U8092 (N_8092,N_6823,N_6515);
nand U8093 (N_8093,N_7347,N_6040);
or U8094 (N_8094,N_7871,N_6553);
nor U8095 (N_8095,N_6866,N_7850);
nand U8096 (N_8096,N_7415,N_7330);
nor U8097 (N_8097,N_6734,N_7262);
and U8098 (N_8098,N_6500,N_6145);
nor U8099 (N_8099,N_6210,N_7054);
or U8100 (N_8100,N_7019,N_6569);
nand U8101 (N_8101,N_6105,N_6375);
nor U8102 (N_8102,N_6586,N_6236);
or U8103 (N_8103,N_7611,N_7070);
nand U8104 (N_8104,N_6746,N_7563);
nand U8105 (N_8105,N_7038,N_6260);
nor U8106 (N_8106,N_6312,N_7314);
nand U8107 (N_8107,N_7652,N_7257);
xnor U8108 (N_8108,N_6118,N_6937);
nand U8109 (N_8109,N_6186,N_7635);
or U8110 (N_8110,N_6615,N_6200);
or U8111 (N_8111,N_6938,N_7506);
and U8112 (N_8112,N_6552,N_6951);
or U8113 (N_8113,N_6712,N_7002);
nor U8114 (N_8114,N_7152,N_7411);
nand U8115 (N_8115,N_7276,N_7647);
nand U8116 (N_8116,N_6444,N_6415);
and U8117 (N_8117,N_7715,N_6458);
nand U8118 (N_8118,N_7892,N_7915);
or U8119 (N_8119,N_7397,N_6378);
nand U8120 (N_8120,N_7924,N_6989);
nor U8121 (N_8121,N_6903,N_7799);
nor U8122 (N_8122,N_6413,N_7642);
or U8123 (N_8123,N_7072,N_6218);
or U8124 (N_8124,N_6773,N_6491);
and U8125 (N_8125,N_7418,N_7727);
nor U8126 (N_8126,N_7194,N_7551);
nand U8127 (N_8127,N_7004,N_6402);
or U8128 (N_8128,N_6598,N_7857);
or U8129 (N_8129,N_7665,N_6097);
nand U8130 (N_8130,N_6052,N_6391);
nor U8131 (N_8131,N_7930,N_7510);
and U8132 (N_8132,N_6162,N_7143);
nand U8133 (N_8133,N_7706,N_7485);
or U8134 (N_8134,N_6871,N_7334);
or U8135 (N_8135,N_6315,N_6669);
nor U8136 (N_8136,N_6778,N_7462);
or U8137 (N_8137,N_7403,N_7406);
or U8138 (N_8138,N_7759,N_6910);
and U8139 (N_8139,N_6879,N_7839);
nand U8140 (N_8140,N_6949,N_6696);
nor U8141 (N_8141,N_7654,N_6738);
nand U8142 (N_8142,N_7104,N_7949);
or U8143 (N_8143,N_7633,N_6830);
xor U8144 (N_8144,N_7882,N_7775);
or U8145 (N_8145,N_6004,N_7632);
xnor U8146 (N_8146,N_6445,N_7414);
nor U8147 (N_8147,N_6787,N_6541);
nor U8148 (N_8148,N_7483,N_7061);
or U8149 (N_8149,N_7575,N_6176);
and U8150 (N_8150,N_6743,N_6220);
or U8151 (N_8151,N_7178,N_7271);
nor U8152 (N_8152,N_6908,N_6056);
nor U8153 (N_8153,N_7046,N_6255);
nor U8154 (N_8154,N_6573,N_7344);
or U8155 (N_8155,N_6675,N_7625);
nor U8156 (N_8156,N_7941,N_6073);
nand U8157 (N_8157,N_7735,N_7313);
nor U8158 (N_8158,N_6887,N_6447);
xor U8159 (N_8159,N_7730,N_6843);
xor U8160 (N_8160,N_6884,N_6400);
and U8161 (N_8161,N_7461,N_6239);
nand U8162 (N_8162,N_6453,N_6619);
and U8163 (N_8163,N_7578,N_6616);
or U8164 (N_8164,N_6739,N_6465);
and U8165 (N_8165,N_7149,N_7203);
and U8166 (N_8166,N_7509,N_7866);
xor U8167 (N_8167,N_7182,N_6668);
nand U8168 (N_8168,N_7186,N_7355);
nand U8169 (N_8169,N_6369,N_7223);
nor U8170 (N_8170,N_7480,N_6256);
and U8171 (N_8171,N_6270,N_7874);
or U8172 (N_8172,N_6149,N_7844);
nand U8173 (N_8173,N_7784,N_6597);
nand U8174 (N_8174,N_7400,N_7726);
or U8175 (N_8175,N_6772,N_6510);
nand U8176 (N_8176,N_7723,N_7371);
nor U8177 (N_8177,N_6958,N_6857);
nor U8178 (N_8178,N_7064,N_6554);
and U8179 (N_8179,N_7111,N_6856);
nor U8180 (N_8180,N_6818,N_6766);
nor U8181 (N_8181,N_7438,N_6602);
nand U8182 (N_8182,N_7770,N_6334);
nor U8183 (N_8183,N_6091,N_7121);
and U8184 (N_8184,N_6412,N_6689);
nand U8185 (N_8185,N_6906,N_7192);
or U8186 (N_8186,N_7096,N_6985);
and U8187 (N_8187,N_7693,N_6529);
and U8188 (N_8188,N_7059,N_6448);
nand U8189 (N_8189,N_6749,N_7995);
and U8190 (N_8190,N_6955,N_7933);
or U8191 (N_8191,N_7683,N_6457);
or U8192 (N_8192,N_6607,N_6132);
nor U8193 (N_8193,N_7685,N_7015);
or U8194 (N_8194,N_7908,N_7686);
and U8195 (N_8195,N_6211,N_7052);
nand U8196 (N_8196,N_6242,N_7237);
or U8197 (N_8197,N_6685,N_7757);
nor U8198 (N_8198,N_7695,N_7848);
or U8199 (N_8199,N_7238,N_7106);
nor U8200 (N_8200,N_7247,N_6889);
or U8201 (N_8201,N_6074,N_6841);
or U8202 (N_8202,N_7130,N_7272);
nor U8203 (N_8203,N_6165,N_6068);
nor U8204 (N_8204,N_6104,N_7164);
or U8205 (N_8205,N_6405,N_6011);
nor U8206 (N_8206,N_6237,N_7780);
and U8207 (N_8207,N_6299,N_6409);
nor U8208 (N_8208,N_6219,N_6950);
nand U8209 (N_8209,N_7615,N_7525);
and U8210 (N_8210,N_6563,N_6677);
and U8211 (N_8211,N_6902,N_6847);
or U8212 (N_8212,N_6396,N_7275);
or U8213 (N_8213,N_7240,N_7678);
nor U8214 (N_8214,N_7634,N_6253);
nor U8215 (N_8215,N_7287,N_6087);
nor U8216 (N_8216,N_7138,N_6125);
nor U8217 (N_8217,N_7000,N_6539);
and U8218 (N_8218,N_6590,N_6966);
nand U8219 (N_8219,N_7699,N_7657);
nor U8220 (N_8220,N_6877,N_6838);
nor U8221 (N_8221,N_7837,N_7714);
nor U8222 (N_8222,N_6854,N_6451);
nor U8223 (N_8223,N_6657,N_6488);
and U8224 (N_8224,N_7207,N_7492);
nand U8225 (N_8225,N_7976,N_7945);
or U8226 (N_8226,N_6029,N_7583);
nand U8227 (N_8227,N_7449,N_6380);
and U8228 (N_8228,N_7339,N_6306);
and U8229 (N_8229,N_6280,N_7389);
nor U8230 (N_8230,N_6631,N_6028);
or U8231 (N_8231,N_6965,N_7140);
or U8232 (N_8232,N_7988,N_7867);
nor U8233 (N_8233,N_6996,N_7938);
or U8234 (N_8234,N_7055,N_7208);
nand U8235 (N_8235,N_6422,N_6069);
and U8236 (N_8236,N_6623,N_7649);
nand U8237 (N_8237,N_7382,N_7133);
nor U8238 (N_8238,N_6649,N_7364);
and U8239 (N_8239,N_6873,N_7564);
nand U8240 (N_8240,N_6355,N_6578);
xor U8241 (N_8241,N_7932,N_6924);
nor U8242 (N_8242,N_7889,N_7943);
nor U8243 (N_8243,N_7264,N_6423);
nor U8244 (N_8244,N_7399,N_7821);
and U8245 (N_8245,N_7802,N_6531);
and U8246 (N_8246,N_6092,N_6379);
nor U8247 (N_8247,N_6796,N_6454);
or U8248 (N_8248,N_7656,N_7550);
nor U8249 (N_8249,N_6030,N_7225);
nand U8250 (N_8250,N_6931,N_7746);
and U8251 (N_8251,N_6090,N_6916);
or U8252 (N_8252,N_7032,N_7128);
and U8253 (N_8253,N_6540,N_6702);
and U8254 (N_8254,N_6436,N_6262);
nand U8255 (N_8255,N_6042,N_6945);
and U8256 (N_8256,N_7120,N_7705);
or U8257 (N_8257,N_6263,N_6751);
nand U8258 (N_8258,N_6067,N_7664);
and U8259 (N_8259,N_6725,N_6706);
nand U8260 (N_8260,N_6645,N_7316);
nand U8261 (N_8261,N_7585,N_6852);
and U8262 (N_8262,N_6711,N_7155);
or U8263 (N_8263,N_6930,N_6957);
and U8264 (N_8264,N_7341,N_7342);
nand U8265 (N_8265,N_6868,N_7567);
or U8266 (N_8266,N_6462,N_7459);
and U8267 (N_8267,N_7612,N_7830);
and U8268 (N_8268,N_6126,N_6456);
and U8269 (N_8269,N_7299,N_6980);
or U8270 (N_8270,N_6635,N_6167);
or U8271 (N_8271,N_7081,N_6490);
or U8272 (N_8272,N_6226,N_7872);
nor U8273 (N_8273,N_6947,N_7346);
nor U8274 (N_8274,N_7547,N_6151);
and U8275 (N_8275,N_6278,N_6007);
and U8276 (N_8276,N_7211,N_7868);
nor U8277 (N_8277,N_7660,N_6566);
nor U8278 (N_8278,N_7498,N_6939);
and U8279 (N_8279,N_6459,N_7343);
and U8280 (N_8280,N_7336,N_6603);
nand U8281 (N_8281,N_7190,N_6538);
and U8282 (N_8282,N_7968,N_6340);
nand U8283 (N_8283,N_7852,N_7880);
or U8284 (N_8284,N_6562,N_7541);
nand U8285 (N_8285,N_6037,N_6522);
and U8286 (N_8286,N_6833,N_6812);
and U8287 (N_8287,N_7952,N_7845);
nand U8288 (N_8288,N_7589,N_6249);
and U8289 (N_8289,N_6960,N_7269);
nor U8290 (N_8290,N_6006,N_6479);
or U8291 (N_8291,N_6723,N_6550);
nand U8292 (N_8292,N_7326,N_7374);
and U8293 (N_8293,N_7380,N_6813);
xor U8294 (N_8294,N_6349,N_7381);
or U8295 (N_8295,N_6690,N_6374);
or U8296 (N_8296,N_6808,N_7917);
or U8297 (N_8297,N_6373,N_6494);
or U8298 (N_8298,N_6428,N_7452);
nor U8299 (N_8299,N_6653,N_6173);
and U8300 (N_8300,N_6478,N_6050);
nor U8301 (N_8301,N_6815,N_7289);
nand U8302 (N_8302,N_7216,N_6560);
and U8303 (N_8303,N_7922,N_7325);
nor U8304 (N_8304,N_6504,N_7690);
and U8305 (N_8305,N_7293,N_6820);
and U8306 (N_8306,N_7849,N_6968);
or U8307 (N_8307,N_6502,N_7692);
and U8308 (N_8308,N_6883,N_7742);
or U8309 (N_8309,N_6112,N_6507);
nor U8310 (N_8310,N_7591,N_6775);
or U8311 (N_8311,N_6322,N_6923);
and U8312 (N_8312,N_6078,N_6790);
or U8313 (N_8313,N_6797,N_6760);
nand U8314 (N_8314,N_6970,N_7358);
or U8315 (N_8315,N_6648,N_6302);
nor U8316 (N_8316,N_7230,N_6952);
nand U8317 (N_8317,N_7417,N_7179);
nand U8318 (N_8318,N_6670,N_6605);
or U8319 (N_8319,N_6464,N_7026);
nor U8320 (N_8320,N_7533,N_6733);
or U8321 (N_8321,N_6977,N_7250);
nand U8322 (N_8322,N_6983,N_7621);
nand U8323 (N_8323,N_7154,N_7445);
and U8324 (N_8324,N_6463,N_6650);
nor U8325 (N_8325,N_7827,N_7761);
and U8326 (N_8326,N_7905,N_6316);
nand U8327 (N_8327,N_7448,N_7752);
and U8328 (N_8328,N_7345,N_6655);
or U8329 (N_8329,N_6013,N_6513);
or U8330 (N_8330,N_7540,N_7259);
nor U8331 (N_8331,N_7513,N_6535);
nand U8332 (N_8332,N_6661,N_6741);
and U8333 (N_8333,N_7393,N_7489);
and U8334 (N_8334,N_7153,N_7764);
nand U8335 (N_8335,N_6424,N_6487);
or U8336 (N_8336,N_7925,N_6821);
or U8337 (N_8337,N_6840,N_7035);
nand U8338 (N_8338,N_7544,N_7451);
nor U8339 (N_8339,N_6274,N_7359);
nor U8340 (N_8340,N_7161,N_7176);
nand U8341 (N_8341,N_7787,N_6286);
and U8342 (N_8342,N_6320,N_7043);
nor U8343 (N_8343,N_7457,N_6356);
and U8344 (N_8344,N_6810,N_7888);
nor U8345 (N_8345,N_6111,N_7370);
xnor U8346 (N_8346,N_6010,N_6547);
nand U8347 (N_8347,N_7719,N_6730);
or U8348 (N_8348,N_6969,N_6561);
and U8349 (N_8349,N_7772,N_7955);
or U8350 (N_8350,N_6680,N_6664);
and U8351 (N_8351,N_7996,N_7440);
and U8352 (N_8352,N_7372,N_6471);
nand U8353 (N_8353,N_6285,N_7768);
or U8354 (N_8354,N_6155,N_7390);
or U8355 (N_8355,N_6043,N_7739);
and U8356 (N_8356,N_6051,N_6867);
or U8357 (N_8357,N_7204,N_6057);
and U8358 (N_8358,N_7170,N_6215);
nor U8359 (N_8359,N_7846,N_7765);
nand U8360 (N_8360,N_7584,N_7684);
or U8361 (N_8361,N_6026,N_6367);
nor U8362 (N_8362,N_6524,N_7638);
nand U8363 (N_8363,N_7185,N_7965);
and U8364 (N_8364,N_7524,N_6736);
or U8365 (N_8365,N_7265,N_7303);
or U8366 (N_8366,N_7701,N_6414);
and U8367 (N_8367,N_7012,N_7137);
or U8368 (N_8368,N_6089,N_6254);
nand U8369 (N_8369,N_7095,N_7721);
and U8370 (N_8370,N_6880,N_7651);
nor U8371 (N_8371,N_6503,N_7893);
and U8372 (N_8372,N_6703,N_6235);
nand U8373 (N_8373,N_6330,N_6558);
nor U8374 (N_8374,N_7713,N_6953);
nor U8375 (N_8375,N_6031,N_6501);
nor U8376 (N_8376,N_7171,N_7515);
or U8377 (N_8377,N_7626,N_6577);
and U8378 (N_8378,N_7362,N_6994);
and U8379 (N_8379,N_7861,N_7720);
or U8380 (N_8380,N_7782,N_6183);
nand U8381 (N_8381,N_6606,N_7385);
and U8382 (N_8382,N_7663,N_6000);
or U8383 (N_8383,N_6544,N_6233);
and U8384 (N_8384,N_7180,N_7779);
nand U8385 (N_8385,N_6727,N_6963);
nand U8386 (N_8386,N_6272,N_7159);
nand U8387 (N_8387,N_6644,N_6836);
xnor U8388 (N_8388,N_7235,N_6296);
nand U8389 (N_8389,N_7841,N_7075);
nand U8390 (N_8390,N_6257,N_7490);
and U8391 (N_8391,N_6663,N_6058);
and U8392 (N_8392,N_7790,N_7831);
or U8393 (N_8393,N_7982,N_6897);
nand U8394 (N_8394,N_7586,N_7937);
nor U8395 (N_8395,N_7156,N_6314);
nor U8396 (N_8396,N_7698,N_7579);
or U8397 (N_8397,N_7931,N_7048);
or U8398 (N_8398,N_7640,N_7375);
and U8399 (N_8399,N_6169,N_7484);
and U8400 (N_8400,N_7007,N_7057);
and U8401 (N_8401,N_6376,N_6925);
or U8402 (N_8402,N_6191,N_7967);
and U8403 (N_8403,N_6292,N_7789);
nand U8404 (N_8404,N_6716,N_7974);
and U8405 (N_8405,N_7368,N_6442);
and U8406 (N_8406,N_6918,N_6357);
nand U8407 (N_8407,N_6846,N_6894);
or U8408 (N_8408,N_6673,N_6325);
xor U8409 (N_8409,N_7274,N_7637);
and U8410 (N_8410,N_6305,N_7447);
nor U8411 (N_8411,N_6021,N_6303);
nor U8412 (N_8412,N_6731,N_6932);
nand U8413 (N_8413,N_7425,N_7103);
nor U8414 (N_8414,N_7220,N_6360);
and U8415 (N_8415,N_6735,N_7512);
or U8416 (N_8416,N_7800,N_6117);
and U8417 (N_8417,N_7530,N_6845);
and U8418 (N_8418,N_7266,N_7184);
nand U8419 (N_8419,N_7576,N_6079);
nor U8420 (N_8420,N_6403,N_7473);
or U8421 (N_8421,N_7901,N_6063);
and U8422 (N_8422,N_6196,N_6217);
or U8423 (N_8423,N_6638,N_6344);
and U8424 (N_8424,N_6826,N_7422);
nand U8425 (N_8425,N_6108,N_7903);
nand U8426 (N_8426,N_6482,N_7788);
and U8427 (N_8427,N_7569,N_6483);
and U8428 (N_8428,N_7919,N_7875);
nand U8429 (N_8429,N_6130,N_6506);
and U8430 (N_8430,N_6288,N_7323);
or U8431 (N_8431,N_7519,N_6758);
nor U8432 (N_8432,N_7722,N_6627);
or U8433 (N_8433,N_7442,N_6801);
nor U8434 (N_8434,N_7009,N_6480);
nand U8435 (N_8435,N_6300,N_7518);
nor U8436 (N_8436,N_7307,N_6318);
or U8437 (N_8437,N_7959,N_6495);
and U8438 (N_8438,N_6364,N_7668);
nand U8439 (N_8439,N_7758,N_6863);
or U8440 (N_8440,N_7441,N_6441);
nor U8441 (N_8441,N_6224,N_6579);
or U8442 (N_8442,N_7309,N_7731);
nor U8443 (N_8443,N_6033,N_6608);
and U8444 (N_8444,N_7934,N_7407);
nand U8445 (N_8445,N_7535,N_6240);
nand U8446 (N_8446,N_7376,N_6595);
or U8447 (N_8447,N_6452,N_6401);
nand U8448 (N_8448,N_6518,N_7793);
or U8449 (N_8449,N_7834,N_6201);
nand U8450 (N_8450,N_6684,N_6973);
nand U8451 (N_8451,N_7123,N_7962);
or U8452 (N_8452,N_6520,N_6956);
or U8453 (N_8453,N_6915,N_7702);
or U8454 (N_8454,N_6946,N_6971);
nand U8455 (N_8455,N_6770,N_7471);
nand U8456 (N_8456,N_6060,N_6848);
and U8457 (N_8457,N_6982,N_6744);
xnor U8458 (N_8458,N_6571,N_6621);
nor U8459 (N_8459,N_7991,N_7682);
nand U8460 (N_8460,N_7039,N_6082);
nor U8461 (N_8461,N_7091,N_6714);
and U8462 (N_8462,N_6389,N_6001);
nand U8463 (N_8463,N_6266,N_7818);
nand U8464 (N_8464,N_6636,N_7936);
or U8465 (N_8465,N_6064,N_6197);
nand U8466 (N_8466,N_6194,N_6086);
and U8467 (N_8467,N_7248,N_6781);
and U8468 (N_8468,N_6726,N_7975);
or U8469 (N_8469,N_6530,N_6851);
or U8470 (N_8470,N_6614,N_7114);
or U8471 (N_8471,N_6204,N_6585);
nor U8472 (N_8472,N_7662,N_6811);
nand U8473 (N_8473,N_6083,N_6695);
nand U8474 (N_8474,N_7408,N_6917);
nor U8475 (N_8475,N_7013,N_6435);
nor U8476 (N_8476,N_7950,N_7387);
nor U8477 (N_8477,N_7082,N_7285);
nand U8478 (N_8478,N_7824,N_7843);
and U8479 (N_8479,N_6241,N_7553);
or U8480 (N_8480,N_7079,N_6881);
nor U8481 (N_8481,N_6345,N_7360);
and U8482 (N_8482,N_6934,N_7317);
and U8483 (N_8483,N_7436,N_6046);
and U8484 (N_8484,N_6071,N_7210);
xor U8485 (N_8485,N_7753,N_7260);
and U8486 (N_8486,N_7828,N_7246);
nor U8487 (N_8487,N_6185,N_7308);
and U8488 (N_8488,N_7177,N_6574);
or U8489 (N_8489,N_7332,N_7588);
and U8490 (N_8490,N_6637,N_7767);
and U8491 (N_8491,N_7413,N_7044);
nand U8492 (N_8492,N_7040,N_6408);
or U8493 (N_8493,N_6816,N_7434);
or U8494 (N_8494,N_7231,N_7398);
nor U8495 (N_8495,N_7354,N_7378);
nand U8496 (N_8496,N_6323,N_6600);
or U8497 (N_8497,N_6913,N_7909);
nand U8498 (N_8498,N_6489,N_7851);
and U8499 (N_8499,N_7501,N_7067);
nand U8500 (N_8500,N_7136,N_7914);
xor U8501 (N_8501,N_7885,N_7792);
and U8502 (N_8502,N_6486,N_6921);
and U8503 (N_8503,N_6193,N_6774);
and U8504 (N_8504,N_7724,N_6549);
nand U8505 (N_8505,N_7083,N_7750);
or U8506 (N_8506,N_7801,N_7078);
and U8507 (N_8507,N_7141,N_6307);
nor U8508 (N_8508,N_7674,N_6780);
and U8509 (N_8509,N_7302,N_7466);
or U8510 (N_8510,N_7605,N_7598);
nor U8511 (N_8511,N_7056,N_6461);
and U8512 (N_8512,N_6206,N_7527);
nor U8513 (N_8513,N_6358,N_6656);
nand U8514 (N_8514,N_7816,N_6519);
nand U8515 (N_8515,N_7197,N_7558);
nand U8516 (N_8516,N_6699,N_6346);
nor U8517 (N_8517,N_7167,N_7717);
nand U8518 (N_8518,N_6337,N_6232);
nor U8519 (N_8519,N_6942,N_7409);
nand U8520 (N_8520,N_6729,N_6234);
or U8521 (N_8521,N_6618,N_6174);
and U8522 (N_8522,N_7337,N_7312);
or U8523 (N_8523,N_7906,N_7958);
and U8524 (N_8524,N_6898,N_6294);
nand U8525 (N_8525,N_6869,N_6831);
and U8526 (N_8526,N_6095,N_7494);
and U8527 (N_8527,N_7045,N_7677);
nor U8528 (N_8528,N_6384,N_6187);
nor U8529 (N_8529,N_7883,N_7107);
and U8530 (N_8530,N_6139,N_6805);
and U8531 (N_8531,N_6628,N_7116);
or U8532 (N_8532,N_6803,N_6152);
nor U8533 (N_8533,N_6639,N_6527);
and U8534 (N_8534,N_6768,N_7146);
nor U8535 (N_8535,N_7430,N_7971);
and U8536 (N_8536,N_6014,N_6765);
or U8537 (N_8537,N_6137,N_7488);
nor U8538 (N_8538,N_7267,N_6273);
or U8539 (N_8539,N_7124,N_7187);
and U8540 (N_8540,N_6406,N_7163);
and U8541 (N_8541,N_7511,N_6771);
or U8542 (N_8542,N_6099,N_7014);
or U8543 (N_8543,N_6327,N_6371);
and U8544 (N_8544,N_6672,N_7556);
nor U8545 (N_8545,N_7884,N_7733);
and U8546 (N_8546,N_7008,N_6313);
nand U8547 (N_8547,N_6041,N_7356);
or U8548 (N_8548,N_6172,N_7549);
xor U8549 (N_8549,N_6496,N_7560);
or U8550 (N_8550,N_7822,N_7162);
and U8551 (N_8551,N_6009,N_6419);
nand U8552 (N_8552,N_7281,N_6724);
nor U8553 (N_8553,N_7165,N_7956);
or U8554 (N_8554,N_7310,N_7804);
and U8555 (N_8555,N_7352,N_6437);
nand U8556 (N_8556,N_6148,N_7249);
and U8557 (N_8557,N_6311,N_6115);
nor U8558 (N_8558,N_6146,N_7126);
and U8559 (N_8559,N_7840,N_6817);
or U8560 (N_8560,N_6431,N_7348);
or U8561 (N_8561,N_6150,N_7963);
and U8562 (N_8562,N_7797,N_6974);
nor U8563 (N_8563,N_7244,N_7623);
or U8564 (N_8564,N_7188,N_6163);
xnor U8565 (N_8565,N_7989,N_7887);
or U8566 (N_8566,N_6686,N_6710);
nor U8567 (N_8567,N_7778,N_7537);
or U8568 (N_8568,N_7301,N_7688);
and U8569 (N_8569,N_7532,N_7985);
or U8570 (N_8570,N_7571,N_7862);
and U8571 (N_8571,N_6276,N_7027);
nand U8572 (N_8572,N_6593,N_7526);
nor U8573 (N_8573,N_6120,N_7439);
or U8574 (N_8574,N_6589,N_6624);
or U8575 (N_8575,N_7108,N_6660);
or U8576 (N_8576,N_6893,N_6251);
or U8577 (N_8577,N_6640,N_6439);
and U8578 (N_8578,N_7771,N_6962);
or U8579 (N_8579,N_7600,N_7648);
nand U8580 (N_8580,N_6864,N_7036);
or U8581 (N_8581,N_6410,N_6003);
nand U8582 (N_8582,N_7495,N_7117);
nor U8583 (N_8583,N_6109,N_6250);
nor U8584 (N_8584,N_7847,N_7311);
or U8585 (N_8585,N_6718,N_7340);
and U8586 (N_8586,N_7331,N_6395);
and U8587 (N_8587,N_6878,N_7189);
or U8588 (N_8588,N_6350,N_7523);
and U8589 (N_8589,N_6434,N_6759);
nor U8590 (N_8590,N_6222,N_7855);
and U8591 (N_8591,N_6829,N_7859);
and U8592 (N_8592,N_7423,N_7954);
or U8593 (N_8593,N_6807,N_6622);
nor U8594 (N_8594,N_7094,N_7670);
and U8595 (N_8595,N_7666,N_6753);
nand U8596 (N_8596,N_7029,N_7707);
and U8597 (N_8597,N_6542,N_7725);
and U8598 (N_8598,N_6025,N_7412);
nand U8599 (N_8599,N_6643,N_6416);
or U8600 (N_8600,N_7740,N_6936);
nor U8601 (N_8601,N_7215,N_7631);
nand U8602 (N_8602,N_7601,N_7115);
nor U8603 (N_8603,N_7773,N_7505);
and U8604 (N_8604,N_7041,N_6331);
and U8605 (N_8605,N_6886,N_6053);
and U8606 (N_8606,N_7997,N_6261);
and U8607 (N_8607,N_7424,N_6212);
or U8608 (N_8608,N_7318,N_7500);
or U8609 (N_8609,N_7920,N_6678);
nor U8610 (N_8610,N_7858,N_6551);
nand U8611 (N_8611,N_7983,N_7838);
nand U8612 (N_8612,N_7377,N_6121);
or U8613 (N_8613,N_7367,N_6388);
or U8614 (N_8614,N_6763,N_7383);
or U8615 (N_8615,N_7675,N_6777);
nor U8616 (N_8616,N_7546,N_7644);
nor U8617 (N_8617,N_7455,N_6609);
or U8618 (N_8618,N_7010,N_7814);
xnor U8619 (N_8619,N_6166,N_6748);
or U8620 (N_8620,N_6526,N_7863);
nand U8621 (N_8621,N_6769,N_6096);
and U8622 (N_8622,N_6264,N_6170);
nor U8623 (N_8623,N_7559,N_6909);
nand U8624 (N_8624,N_7680,N_7711);
nand U8625 (N_8625,N_6246,N_6157);
nor U8626 (N_8626,N_6580,N_6417);
and U8627 (N_8627,N_7291,N_7566);
or U8628 (N_8628,N_7785,N_7454);
nand U8629 (N_8629,N_7273,N_6433);
nor U8630 (N_8630,N_6998,N_6175);
and U8631 (N_8631,N_7338,N_7077);
nand U8632 (N_8632,N_6039,N_6647);
and U8633 (N_8633,N_6216,N_6283);
or U8634 (N_8634,N_6785,N_7658);
nor U8635 (N_8635,N_7493,N_7810);
nand U8636 (N_8636,N_6565,N_7998);
nor U8637 (N_8637,N_7066,N_7357);
or U8638 (N_8638,N_7916,N_6583);
and U8639 (N_8639,N_7681,N_7645);
nand U8640 (N_8640,N_7873,N_7661);
nor U8641 (N_8641,N_7708,N_7745);
and U8642 (N_8642,N_7960,N_7456);
and U8643 (N_8643,N_6022,N_6077);
nand U8644 (N_8644,N_7294,N_6047);
nor U8645 (N_8645,N_6298,N_6819);
and U8646 (N_8646,N_6098,N_7545);
nor U8647 (N_8647,N_6243,N_7570);
nand U8648 (N_8648,N_6189,N_6475);
and U8649 (N_8649,N_6641,N_6339);
nand U8650 (N_8650,N_6370,N_6704);
or U8651 (N_8651,N_7193,N_6158);
or U8652 (N_8652,N_7596,N_7481);
nor U8653 (N_8653,N_7534,N_6421);
or U8654 (N_8654,N_6865,N_6188);
and U8655 (N_8655,N_7384,N_7636);
nand U8656 (N_8656,N_7217,N_6427);
nand U8657 (N_8657,N_6352,N_6065);
nor U8658 (N_8658,N_6289,N_7306);
nand U8659 (N_8659,N_7929,N_6179);
nand U8660 (N_8660,N_6275,N_7410);
nand U8661 (N_8661,N_6806,N_7232);
and U8662 (N_8662,N_6267,N_6928);
nor U8663 (N_8663,N_7234,N_7503);
and U8664 (N_8664,N_7158,N_7463);
nor U8665 (N_8665,N_6694,N_7175);
nand U8666 (N_8666,N_6070,N_6832);
nor U8667 (N_8667,N_6244,N_6161);
nor U8668 (N_8668,N_6905,N_7944);
nand U8669 (N_8669,N_6548,N_6363);
and U8670 (N_8670,N_7297,N_7899);
and U8671 (N_8671,N_7864,N_7940);
nor U8672 (N_8672,N_6122,N_6700);
or U8673 (N_8673,N_6896,N_7653);
nand U8674 (N_8674,N_6683,N_6116);
xor U8675 (N_8675,N_7536,N_7710);
nand U8676 (N_8676,N_6521,N_6135);
and U8677 (N_8677,N_6024,N_7142);
nand U8678 (N_8678,N_7756,N_7811);
nand U8679 (N_8679,N_7603,N_6038);
nor U8680 (N_8680,N_7098,N_6667);
xor U8681 (N_8681,N_7351,N_6858);
nor U8682 (N_8682,N_7460,N_6366);
and U8683 (N_8683,N_6027,N_6114);
and U8684 (N_8684,N_7102,N_6533);
and U8685 (N_8685,N_7689,N_6691);
nand U8686 (N_8686,N_6511,N_7392);
or U8687 (N_8687,N_7295,N_6418);
or U8688 (N_8688,N_7349,N_7910);
nor U8689 (N_8689,N_6449,N_7539);
and U8690 (N_8690,N_6567,N_6922);
and U8691 (N_8691,N_7978,N_7003);
nand U8692 (N_8692,N_7900,N_7218);
and U8693 (N_8693,N_6245,N_6659);
or U8694 (N_8694,N_7529,N_6555);
and U8695 (N_8695,N_7428,N_6066);
and U8696 (N_8696,N_7835,N_6570);
and U8697 (N_8697,N_6192,N_6582);
nor U8698 (N_8698,N_7966,N_7592);
nor U8699 (N_8699,N_6892,N_7531);
or U8700 (N_8700,N_6764,N_6361);
xor U8701 (N_8701,N_7361,N_7491);
nand U8702 (N_8702,N_7369,N_6682);
or U8703 (N_8703,N_6814,N_6676);
xnor U8704 (N_8704,N_7641,N_7813);
and U8705 (N_8705,N_7300,N_7894);
nand U8706 (N_8706,N_6085,N_7290);
nor U8707 (N_8707,N_6398,N_6850);
nor U8708 (N_8708,N_7166,N_6708);
or U8709 (N_8709,N_6862,N_6207);
nand U8710 (N_8710,N_7574,N_7429);
or U8711 (N_8711,N_7748,N_6230);
nand U8712 (N_8712,N_7659,N_6497);
or U8713 (N_8713,N_7198,N_6611);
and U8714 (N_8714,N_6055,N_6979);
or U8715 (N_8715,N_6975,N_7458);
or U8716 (N_8716,N_7305,N_7783);
nor U8717 (N_8717,N_6252,N_6633);
and U8718 (N_8718,N_6438,N_6420);
and U8719 (N_8719,N_7798,N_7687);
nor U8720 (N_8720,N_6336,N_6002);
nand U8721 (N_8721,N_6492,N_7034);
or U8722 (N_8722,N_6178,N_6556);
nand U8723 (N_8723,N_6329,N_7063);
nand U8724 (N_8724,N_7522,N_7497);
nor U8725 (N_8725,N_7037,N_6259);
nand U8726 (N_8726,N_6919,N_6646);
and U8727 (N_8727,N_7627,N_7671);
or U8728 (N_8728,N_7927,N_6692);
nand U8729 (N_8729,N_6849,N_6720);
nand U8730 (N_8730,N_6855,N_7619);
and U8731 (N_8731,N_6128,N_7581);
or U8732 (N_8732,N_6477,N_6757);
nand U8733 (N_8733,N_7286,N_7239);
or U8734 (N_8734,N_7568,N_6929);
or U8735 (N_8735,N_6876,N_6177);
nand U8736 (N_8736,N_6625,N_7254);
and U8737 (N_8737,N_7806,N_7577);
nor U8738 (N_8738,N_7912,N_7878);
nand U8739 (N_8739,N_6354,N_7419);
nor U8740 (N_8740,N_7898,N_7292);
nor U8741 (N_8741,N_7921,N_7833);
or U8742 (N_8742,N_6036,N_6332);
nor U8743 (N_8743,N_7097,N_6168);
nor U8744 (N_8744,N_6839,N_7516);
or U8745 (N_8745,N_6756,N_6927);
or U8746 (N_8746,N_6317,N_7199);
or U8747 (N_8747,N_7870,N_7209);
or U8748 (N_8748,N_6258,N_7482);
nor U8749 (N_8749,N_6101,N_7953);
nand U8750 (N_8750,N_6016,N_7395);
and U8751 (N_8751,N_7980,N_6613);
nor U8752 (N_8752,N_6804,N_6269);
or U8753 (N_8753,N_7796,N_7221);
nor U8754 (N_8754,N_7613,N_7744);
or U8755 (N_8755,N_7401,N_6612);
and U8756 (N_8756,N_7023,N_7794);
and U8757 (N_8757,N_7994,N_6310);
nor U8758 (N_8758,N_7477,N_7431);
or U8759 (N_8759,N_7319,N_7791);
and U8760 (N_8760,N_6509,N_7886);
and U8761 (N_8761,N_6328,N_6214);
nand U8762 (N_8762,N_7183,N_6875);
nand U8763 (N_8763,N_7979,N_7608);
or U8764 (N_8764,N_7089,N_7595);
or U8765 (N_8765,N_7981,N_6156);
or U8766 (N_8766,N_7947,N_7504);
nand U8767 (N_8767,N_7964,N_7131);
nor U8768 (N_8768,N_7243,N_6557);
nand U8769 (N_8769,N_7672,N_7446);
and U8770 (N_8770,N_7327,N_6467);
nand U8771 (N_8771,N_7805,N_7021);
nand U8772 (N_8772,N_6159,N_6842);
nor U8773 (N_8773,N_6629,N_7760);
and U8774 (N_8774,N_6658,N_7557);
or U8775 (N_8775,N_6499,N_7283);
or U8776 (N_8776,N_6171,N_6020);
and U8777 (N_8777,N_6872,N_6750);
and U8778 (N_8778,N_6576,N_6824);
nor U8779 (N_8779,N_7018,N_6943);
nor U8780 (N_8780,N_7881,N_7853);
nor U8781 (N_8781,N_6291,N_7561);
or U8782 (N_8782,N_7977,N_7144);
and U8783 (N_8783,N_6123,N_6113);
and U8784 (N_8784,N_7548,N_6662);
or U8785 (N_8785,N_6093,N_6907);
and U8786 (N_8786,N_7826,N_6338);
nor U8787 (N_8787,N_7487,N_7781);
and U8788 (N_8788,N_6870,N_6941);
and U8789 (N_8789,N_7475,N_6732);
or U8790 (N_8790,N_7050,N_7233);
and U8791 (N_8791,N_6802,N_6634);
nand U8792 (N_8792,N_6584,N_7594);
or U8793 (N_8793,N_6707,N_6992);
and U8794 (N_8794,N_7145,N_7453);
or U8795 (N_8795,N_6697,N_7622);
or U8796 (N_8796,N_7437,N_6795);
nand U8797 (N_8797,N_6594,N_7051);
nand U8798 (N_8798,N_6248,N_7172);
nor U8799 (N_8799,N_6372,N_7277);
nor U8800 (N_8800,N_6834,N_6935);
nand U8801 (N_8801,N_7865,N_6231);
nand U8802 (N_8802,N_7105,N_7024);
nor U8803 (N_8803,N_7261,N_6333);
or U8804 (N_8804,N_6075,N_7226);
and U8805 (N_8805,N_7562,N_7020);
or U8806 (N_8806,N_7716,N_6717);
nand U8807 (N_8807,N_7450,N_7517);
and U8808 (N_8808,N_7469,N_6701);
or U8809 (N_8809,N_7069,N_7420);
and U8810 (N_8810,N_6205,N_7624);
nor U8811 (N_8811,N_7270,N_7842);
nand U8812 (N_8812,N_6319,N_7074);
nor U8813 (N_8813,N_7769,N_7435);
or U8814 (N_8814,N_7134,N_7280);
nand U8815 (N_8815,N_7200,N_7538);
or U8816 (N_8816,N_6119,N_7972);
or U8817 (N_8817,N_6713,N_6693);
and U8818 (N_8818,N_6153,N_7942);
or U8819 (N_8819,N_7829,N_7099);
nor U8820 (N_8820,N_7602,N_6160);
nor U8821 (N_8821,N_7322,N_6164);
nand U8822 (N_8822,N_7443,N_7465);
and U8823 (N_8823,N_6238,N_6888);
or U8824 (N_8824,N_7135,N_7113);
or U8825 (N_8825,N_7897,N_6912);
nor U8826 (N_8826,N_6142,N_6018);
and U8827 (N_8827,N_6959,N_6144);
nand U8828 (N_8828,N_6809,N_7667);
or U8829 (N_8829,N_6525,N_6180);
and U8830 (N_8830,N_6523,N_6440);
nor U8831 (N_8831,N_7224,N_6698);
nor U8832 (N_8832,N_7404,N_7090);
nand U8833 (N_8833,N_6394,N_6308);
or U8834 (N_8834,N_6987,N_7022);
and U8835 (N_8835,N_6995,N_6382);
and U8836 (N_8836,N_7582,N_6110);
or U8837 (N_8837,N_7353,N_6767);
or U8838 (N_8838,N_7031,N_7125);
or U8839 (N_8839,N_6972,N_6859);
nor U8840 (N_8840,N_6293,N_7391);
nor U8841 (N_8841,N_7328,N_7470);
or U8842 (N_8842,N_6353,N_7304);
and U8843 (N_8843,N_7807,N_6792);
nor U8844 (N_8844,N_7350,N_6844);
xnor U8845 (N_8845,N_6048,N_6512);
nand U8846 (N_8846,N_6800,N_6926);
nor U8847 (N_8847,N_7948,N_7877);
nor U8848 (N_8848,N_6049,N_6754);
or U8849 (N_8849,N_6469,N_7017);
nor U8850 (N_8850,N_6493,N_7084);
nor U8851 (N_8851,N_6537,N_6687);
and U8852 (N_8852,N_6545,N_6136);
nand U8853 (N_8853,N_7990,N_6592);
or U8854 (N_8854,N_6347,N_6993);
nor U8855 (N_8855,N_6791,N_6446);
nor U8856 (N_8856,N_7896,N_7825);
and U8857 (N_8857,N_6377,N_7694);
nor U8858 (N_8858,N_6032,N_6381);
and U8859 (N_8859,N_6481,N_6059);
and U8860 (N_8860,N_7957,N_7999);
and U8861 (N_8861,N_7521,N_7747);
or U8862 (N_8862,N_6798,N_7712);
or U8863 (N_8863,N_7122,N_7655);
or U8864 (N_8864,N_6485,N_6399);
nand U8865 (N_8865,N_6054,N_6737);
or U8866 (N_8866,N_7736,N_6528);
and U8867 (N_8867,N_7365,N_7242);
and U8868 (N_8868,N_6835,N_6035);
nand U8869 (N_8869,N_6591,N_7795);
and U8870 (N_8870,N_7073,N_6860);
nand U8871 (N_8871,N_6131,N_6788);
nor U8872 (N_8872,N_7650,N_7150);
or U8873 (N_8873,N_6761,N_6705);
and U8874 (N_8874,N_6304,N_7058);
and U8875 (N_8875,N_6432,N_7042);
and U8876 (N_8876,N_7618,N_6450);
and U8877 (N_8877,N_6961,N_6940);
or U8878 (N_8878,N_6991,N_6103);
nand U8879 (N_8879,N_7992,N_7587);
or U8880 (N_8880,N_7629,N_7212);
and U8881 (N_8881,N_7607,N_6080);
or U8882 (N_8882,N_6630,N_6933);
nor U8883 (N_8883,N_7405,N_6335);
or U8884 (N_8884,N_6321,N_7174);
nor U8885 (N_8885,N_7993,N_6202);
nand U8886 (N_8886,N_6134,N_6468);
and U8887 (N_8887,N_6182,N_7606);
nand U8888 (N_8888,N_7777,N_7628);
nor U8889 (N_8889,N_7643,N_7935);
and U8890 (N_8890,N_7514,N_6978);
nand U8891 (N_8891,N_6390,N_6124);
nand U8892 (N_8892,N_6904,N_6745);
nand U8893 (N_8893,N_7815,N_6393);
and U8894 (N_8894,N_7709,N_7472);
nand U8895 (N_8895,N_7969,N_7001);
and U8896 (N_8896,N_6740,N_6094);
nand U8897 (N_8897,N_7774,N_7507);
xnor U8898 (N_8898,N_6789,N_7033);
and U8899 (N_8899,N_7229,N_7432);
or U8900 (N_8900,N_7256,N_7416);
nand U8901 (N_8901,N_7076,N_7573);
or U8902 (N_8902,N_6005,N_7946);
and U8903 (N_8903,N_6279,N_7543);
and U8904 (N_8904,N_7854,N_7093);
and U8905 (N_8905,N_7836,N_7580);
or U8906 (N_8906,N_7100,N_7427);
or U8907 (N_8907,N_7205,N_7426);
or U8908 (N_8908,N_6719,N_6228);
or U8909 (N_8909,N_6012,N_7421);
or U8910 (N_8910,N_7895,N_7542);
nor U8911 (N_8911,N_6084,N_7869);
or U8912 (N_8912,N_7743,N_6747);
nor U8913 (N_8913,N_7025,N_6674);
and U8914 (N_8914,N_6779,N_6665);
or U8915 (N_8915,N_6762,N_6223);
nand U8916 (N_8916,N_7065,N_7755);
and U8917 (N_8917,N_6407,N_7911);
nand U8918 (N_8918,N_6404,N_6359);
nor U8919 (N_8919,N_6341,N_7278);
nand U8920 (N_8920,N_7808,N_6392);
and U8921 (N_8921,N_7373,N_6920);
and U8922 (N_8922,N_7252,N_6853);
or U8923 (N_8923,N_6755,N_6543);
or U8924 (N_8924,N_7669,N_6911);
or U8925 (N_8925,N_7110,N_7552);
nand U8926 (N_8926,N_7918,N_6651);
or U8927 (N_8927,N_7499,N_7386);
nand U8928 (N_8928,N_6536,N_7258);
nor U8929 (N_8929,N_6455,N_7766);
and U8930 (N_8930,N_6715,N_6794);
nand U8931 (N_8931,N_6147,N_6981);
nor U8932 (N_8932,N_7913,N_7876);
nor U8933 (N_8933,N_6365,N_7614);
and U8934 (N_8934,N_7639,N_7478);
or U8935 (N_8935,N_7738,N_6967);
xor U8936 (N_8936,N_6885,N_7987);
nor U8937 (N_8937,N_7251,N_7590);
nor U8938 (N_8938,N_7890,N_7394);
and U8939 (N_8939,N_6154,N_7109);
and U8940 (N_8940,N_7227,N_6106);
nand U8941 (N_8941,N_6534,N_7236);
nand U8942 (N_8942,N_7820,N_6822);
and U8943 (N_8943,N_6107,N_7222);
and U8944 (N_8944,N_6861,N_7860);
and U8945 (N_8945,N_7088,N_7284);
or U8946 (N_8946,N_7812,N_6709);
and U8947 (N_8947,N_6784,N_7169);
and U8948 (N_8948,N_6343,N_6425);
nor U8949 (N_8949,N_7191,N_7049);
and U8950 (N_8950,N_7728,N_6326);
nor U8951 (N_8951,N_6596,N_6948);
nor U8952 (N_8952,N_6397,N_6914);
nor U8953 (N_8953,N_7379,N_6017);
nor U8954 (N_8954,N_7555,N_6088);
nand U8955 (N_8955,N_6282,N_6516);
nand U8956 (N_8956,N_7809,N_6498);
nor U8957 (N_8957,N_6181,N_6825);
nor U8958 (N_8958,N_6599,N_6828);
xnor U8959 (N_8959,N_7803,N_6140);
nor U8960 (N_8960,N_6015,N_7762);
and U8961 (N_8961,N_7030,N_6290);
or U8962 (N_8962,N_7704,N_7679);
nand U8963 (N_8963,N_6301,N_6061);
and U8964 (N_8964,N_7011,N_6209);
nor U8965 (N_8965,N_6782,N_6954);
nand U8966 (N_8966,N_7151,N_7970);
nand U8967 (N_8967,N_7718,N_7160);
nand U8968 (N_8968,N_6309,N_7751);
nor U8969 (N_8969,N_6976,N_6127);
nor U8970 (N_8970,N_7279,N_7282);
nand U8971 (N_8971,N_6271,N_7926);
and U8972 (N_8972,N_6190,N_7502);
and U8973 (N_8973,N_6575,N_6102);
nor U8974 (N_8974,N_6986,N_6411);
and U8975 (N_8975,N_7902,N_6642);
nand U8976 (N_8976,N_6671,N_7396);
nor U8977 (N_8977,N_7464,N_6348);
and U8978 (N_8978,N_6281,N_6062);
or U8979 (N_8979,N_7823,N_7363);
nand U8980 (N_8980,N_6514,N_7086);
nand U8981 (N_8981,N_6900,N_6901);
and U8982 (N_8982,N_7335,N_7028);
nand U8983 (N_8983,N_7060,N_6221);
and U8984 (N_8984,N_7528,N_7324);
nor U8985 (N_8985,N_7597,N_7129);
nor U8986 (N_8986,N_6287,N_6874);
and U8987 (N_8987,N_7255,N_6890);
and U8988 (N_8988,N_7201,N_6652);
and U8989 (N_8989,N_7053,N_6997);
or U8990 (N_8990,N_7604,N_7092);
nor U8991 (N_8991,N_7697,N_6837);
xnor U8992 (N_8992,N_7329,N_6899);
and U8993 (N_8993,N_6386,N_6268);
or U8994 (N_8994,N_6559,N_7071);
nor U8995 (N_8995,N_7939,N_7676);
nor U8996 (N_8996,N_6133,N_7754);
nor U8997 (N_8997,N_7168,N_7181);
nand U8998 (N_8998,N_7321,N_7554);
and U8999 (N_8999,N_7119,N_6141);
nor U9000 (N_9000,N_7331,N_7353);
nand U9001 (N_9001,N_6850,N_6313);
or U9002 (N_9002,N_6108,N_7141);
nor U9003 (N_9003,N_7756,N_6559);
and U9004 (N_9004,N_6568,N_7881);
and U9005 (N_9005,N_6900,N_6652);
and U9006 (N_9006,N_6676,N_6830);
nor U9007 (N_9007,N_7009,N_7587);
or U9008 (N_9008,N_6798,N_7959);
and U9009 (N_9009,N_6119,N_6998);
nor U9010 (N_9010,N_6500,N_6826);
or U9011 (N_9011,N_6224,N_6782);
nand U9012 (N_9012,N_7956,N_7981);
and U9013 (N_9013,N_7687,N_6094);
and U9014 (N_9014,N_6941,N_6939);
or U9015 (N_9015,N_7600,N_6304);
nor U9016 (N_9016,N_6825,N_6693);
nand U9017 (N_9017,N_6030,N_7017);
or U9018 (N_9018,N_7981,N_7927);
nor U9019 (N_9019,N_6589,N_6114);
nor U9020 (N_9020,N_6453,N_7765);
or U9021 (N_9021,N_6494,N_7311);
and U9022 (N_9022,N_7076,N_6617);
and U9023 (N_9023,N_7705,N_6743);
or U9024 (N_9024,N_6113,N_7797);
and U9025 (N_9025,N_7569,N_7781);
and U9026 (N_9026,N_7400,N_6642);
and U9027 (N_9027,N_7529,N_6113);
and U9028 (N_9028,N_6859,N_6322);
nand U9029 (N_9029,N_6463,N_7079);
and U9030 (N_9030,N_6936,N_6116);
nand U9031 (N_9031,N_6200,N_7923);
nor U9032 (N_9032,N_6606,N_6286);
nand U9033 (N_9033,N_7784,N_7210);
nor U9034 (N_9034,N_7106,N_6796);
or U9035 (N_9035,N_6594,N_6691);
nor U9036 (N_9036,N_7741,N_7310);
or U9037 (N_9037,N_6068,N_7027);
and U9038 (N_9038,N_6525,N_6024);
or U9039 (N_9039,N_7195,N_6171);
and U9040 (N_9040,N_7517,N_7411);
and U9041 (N_9041,N_6751,N_7960);
and U9042 (N_9042,N_6334,N_6210);
and U9043 (N_9043,N_6904,N_7264);
or U9044 (N_9044,N_6232,N_6357);
or U9045 (N_9045,N_7891,N_6856);
nor U9046 (N_9046,N_7614,N_7564);
nor U9047 (N_9047,N_7599,N_6620);
and U9048 (N_9048,N_6289,N_6988);
nor U9049 (N_9049,N_7076,N_6508);
or U9050 (N_9050,N_6414,N_6686);
and U9051 (N_9051,N_7549,N_6838);
nand U9052 (N_9052,N_7398,N_6043);
or U9053 (N_9053,N_7059,N_6382);
nor U9054 (N_9054,N_6921,N_6452);
or U9055 (N_9055,N_7030,N_7761);
and U9056 (N_9056,N_7118,N_7373);
and U9057 (N_9057,N_6695,N_7301);
nand U9058 (N_9058,N_6174,N_6729);
and U9059 (N_9059,N_6682,N_7880);
or U9060 (N_9060,N_6283,N_6732);
or U9061 (N_9061,N_7089,N_6681);
nand U9062 (N_9062,N_6995,N_7467);
nor U9063 (N_9063,N_7111,N_6813);
or U9064 (N_9064,N_6638,N_7297);
nand U9065 (N_9065,N_6413,N_6683);
or U9066 (N_9066,N_6694,N_6403);
or U9067 (N_9067,N_6444,N_6563);
and U9068 (N_9068,N_6954,N_7003);
and U9069 (N_9069,N_6932,N_6810);
and U9070 (N_9070,N_6766,N_6299);
and U9071 (N_9071,N_7947,N_6550);
and U9072 (N_9072,N_7266,N_6467);
or U9073 (N_9073,N_7123,N_7148);
nor U9074 (N_9074,N_6699,N_6056);
nand U9075 (N_9075,N_7004,N_6192);
or U9076 (N_9076,N_7354,N_7572);
or U9077 (N_9077,N_6695,N_7835);
nor U9078 (N_9078,N_6081,N_7842);
and U9079 (N_9079,N_6096,N_6917);
nand U9080 (N_9080,N_7422,N_6596);
or U9081 (N_9081,N_6733,N_6193);
or U9082 (N_9082,N_6836,N_7472);
and U9083 (N_9083,N_6264,N_7902);
or U9084 (N_9084,N_6158,N_7721);
nand U9085 (N_9085,N_7996,N_6459);
nor U9086 (N_9086,N_7854,N_6656);
nor U9087 (N_9087,N_6762,N_6696);
or U9088 (N_9088,N_6298,N_7147);
nand U9089 (N_9089,N_7754,N_7582);
and U9090 (N_9090,N_7659,N_6811);
nor U9091 (N_9091,N_7760,N_6214);
nor U9092 (N_9092,N_7286,N_6984);
nand U9093 (N_9093,N_7983,N_7348);
and U9094 (N_9094,N_6155,N_6774);
or U9095 (N_9095,N_7464,N_6235);
nor U9096 (N_9096,N_6742,N_7507);
nor U9097 (N_9097,N_7573,N_7552);
xor U9098 (N_9098,N_7899,N_7076);
nor U9099 (N_9099,N_6075,N_7942);
and U9100 (N_9100,N_6089,N_6799);
nor U9101 (N_9101,N_7601,N_7573);
and U9102 (N_9102,N_7795,N_7849);
nor U9103 (N_9103,N_6651,N_6585);
or U9104 (N_9104,N_7179,N_7305);
and U9105 (N_9105,N_7686,N_7118);
or U9106 (N_9106,N_7294,N_7397);
or U9107 (N_9107,N_6023,N_6768);
or U9108 (N_9108,N_7809,N_7787);
and U9109 (N_9109,N_6894,N_6349);
nor U9110 (N_9110,N_6367,N_6886);
or U9111 (N_9111,N_7013,N_7177);
and U9112 (N_9112,N_7535,N_7581);
and U9113 (N_9113,N_6334,N_7644);
nor U9114 (N_9114,N_7518,N_7041);
and U9115 (N_9115,N_6897,N_6508);
nor U9116 (N_9116,N_7981,N_7972);
and U9117 (N_9117,N_6616,N_6797);
nor U9118 (N_9118,N_6918,N_7399);
nor U9119 (N_9119,N_6481,N_7581);
nand U9120 (N_9120,N_7416,N_6150);
nand U9121 (N_9121,N_7136,N_7803);
nor U9122 (N_9122,N_7683,N_7438);
and U9123 (N_9123,N_6284,N_6952);
nand U9124 (N_9124,N_6977,N_6882);
nand U9125 (N_9125,N_7146,N_6445);
nor U9126 (N_9126,N_6074,N_7871);
nand U9127 (N_9127,N_7401,N_7838);
or U9128 (N_9128,N_7530,N_7755);
nor U9129 (N_9129,N_7029,N_7493);
nor U9130 (N_9130,N_7781,N_7116);
nor U9131 (N_9131,N_7845,N_6286);
and U9132 (N_9132,N_7984,N_7396);
or U9133 (N_9133,N_7821,N_6317);
nand U9134 (N_9134,N_7371,N_6096);
and U9135 (N_9135,N_6333,N_6547);
and U9136 (N_9136,N_6336,N_6378);
nand U9137 (N_9137,N_6579,N_7336);
nor U9138 (N_9138,N_7211,N_6204);
nand U9139 (N_9139,N_6980,N_6246);
nand U9140 (N_9140,N_7175,N_6863);
and U9141 (N_9141,N_7484,N_7952);
and U9142 (N_9142,N_7407,N_7747);
nor U9143 (N_9143,N_6036,N_6708);
and U9144 (N_9144,N_7413,N_7608);
nand U9145 (N_9145,N_6975,N_6528);
and U9146 (N_9146,N_7971,N_7788);
nor U9147 (N_9147,N_6775,N_7965);
or U9148 (N_9148,N_7633,N_6841);
or U9149 (N_9149,N_6182,N_7939);
or U9150 (N_9150,N_7256,N_6381);
and U9151 (N_9151,N_6705,N_7852);
and U9152 (N_9152,N_6303,N_6120);
nor U9153 (N_9153,N_6853,N_6557);
nor U9154 (N_9154,N_6907,N_7085);
and U9155 (N_9155,N_6851,N_6878);
and U9156 (N_9156,N_7167,N_7091);
nor U9157 (N_9157,N_6941,N_6893);
or U9158 (N_9158,N_6480,N_6332);
nand U9159 (N_9159,N_6295,N_6563);
nand U9160 (N_9160,N_6045,N_6339);
nand U9161 (N_9161,N_7369,N_6936);
and U9162 (N_9162,N_6077,N_7522);
nor U9163 (N_9163,N_7003,N_6360);
and U9164 (N_9164,N_6496,N_6222);
or U9165 (N_9165,N_6529,N_6243);
nor U9166 (N_9166,N_7587,N_6541);
nand U9167 (N_9167,N_7653,N_7828);
or U9168 (N_9168,N_7379,N_6229);
nor U9169 (N_9169,N_6392,N_6063);
nand U9170 (N_9170,N_7132,N_6812);
nor U9171 (N_9171,N_7911,N_7983);
nor U9172 (N_9172,N_7814,N_6856);
nand U9173 (N_9173,N_6951,N_6357);
or U9174 (N_9174,N_7111,N_7077);
and U9175 (N_9175,N_6199,N_7891);
and U9176 (N_9176,N_7734,N_7902);
nor U9177 (N_9177,N_6510,N_7042);
and U9178 (N_9178,N_7626,N_6290);
nand U9179 (N_9179,N_6533,N_6938);
nor U9180 (N_9180,N_7200,N_7594);
or U9181 (N_9181,N_6375,N_6036);
nor U9182 (N_9182,N_7471,N_7240);
or U9183 (N_9183,N_6610,N_7655);
or U9184 (N_9184,N_6761,N_7492);
and U9185 (N_9185,N_6394,N_7439);
or U9186 (N_9186,N_6322,N_7966);
nor U9187 (N_9187,N_7886,N_7906);
and U9188 (N_9188,N_7800,N_7443);
nor U9189 (N_9189,N_6122,N_7313);
and U9190 (N_9190,N_6982,N_7578);
or U9191 (N_9191,N_6441,N_7777);
and U9192 (N_9192,N_7492,N_6967);
nand U9193 (N_9193,N_6990,N_7239);
nand U9194 (N_9194,N_6169,N_6534);
nand U9195 (N_9195,N_7536,N_7802);
and U9196 (N_9196,N_7603,N_7060);
or U9197 (N_9197,N_6426,N_7829);
and U9198 (N_9198,N_7285,N_7312);
nand U9199 (N_9199,N_7118,N_6087);
nor U9200 (N_9200,N_7443,N_6682);
nor U9201 (N_9201,N_7726,N_6850);
nor U9202 (N_9202,N_6177,N_7897);
and U9203 (N_9203,N_7461,N_7918);
xnor U9204 (N_9204,N_6005,N_6586);
or U9205 (N_9205,N_7103,N_7831);
nand U9206 (N_9206,N_7750,N_7813);
or U9207 (N_9207,N_7558,N_6905);
nand U9208 (N_9208,N_6757,N_6359);
nor U9209 (N_9209,N_7103,N_6687);
or U9210 (N_9210,N_6360,N_6821);
or U9211 (N_9211,N_7337,N_6850);
nor U9212 (N_9212,N_7669,N_6789);
and U9213 (N_9213,N_6106,N_7565);
or U9214 (N_9214,N_6108,N_7367);
nand U9215 (N_9215,N_7504,N_7455);
nor U9216 (N_9216,N_6637,N_6838);
nor U9217 (N_9217,N_6591,N_6099);
nor U9218 (N_9218,N_7769,N_6063);
nand U9219 (N_9219,N_6876,N_6946);
nand U9220 (N_9220,N_7597,N_6067);
and U9221 (N_9221,N_7300,N_6291);
nand U9222 (N_9222,N_7852,N_6287);
and U9223 (N_9223,N_7756,N_6710);
and U9224 (N_9224,N_6704,N_7313);
nor U9225 (N_9225,N_6238,N_7748);
xnor U9226 (N_9226,N_7634,N_6364);
or U9227 (N_9227,N_7140,N_7257);
or U9228 (N_9228,N_7558,N_7994);
nor U9229 (N_9229,N_7147,N_6717);
nor U9230 (N_9230,N_7126,N_6560);
or U9231 (N_9231,N_6656,N_6624);
or U9232 (N_9232,N_7275,N_7233);
and U9233 (N_9233,N_6788,N_6137);
nor U9234 (N_9234,N_7739,N_6446);
or U9235 (N_9235,N_7827,N_7149);
nor U9236 (N_9236,N_7995,N_6319);
nand U9237 (N_9237,N_7471,N_7321);
nor U9238 (N_9238,N_7517,N_7396);
nand U9239 (N_9239,N_7356,N_6444);
nor U9240 (N_9240,N_7397,N_7886);
nand U9241 (N_9241,N_6384,N_6603);
and U9242 (N_9242,N_7552,N_7948);
and U9243 (N_9243,N_7951,N_7248);
or U9244 (N_9244,N_7400,N_7485);
nor U9245 (N_9245,N_6641,N_6414);
and U9246 (N_9246,N_6306,N_7013);
nor U9247 (N_9247,N_7157,N_6480);
and U9248 (N_9248,N_6387,N_7793);
and U9249 (N_9249,N_6727,N_7447);
nor U9250 (N_9250,N_7977,N_6166);
and U9251 (N_9251,N_7668,N_6837);
nand U9252 (N_9252,N_6073,N_7472);
nand U9253 (N_9253,N_7878,N_7012);
nor U9254 (N_9254,N_7647,N_6513);
or U9255 (N_9255,N_6657,N_6534);
or U9256 (N_9256,N_6434,N_6745);
nand U9257 (N_9257,N_7787,N_6004);
nand U9258 (N_9258,N_7785,N_7907);
and U9259 (N_9259,N_6215,N_6553);
nand U9260 (N_9260,N_6597,N_7570);
and U9261 (N_9261,N_7438,N_6903);
and U9262 (N_9262,N_7621,N_6640);
or U9263 (N_9263,N_7149,N_7950);
nor U9264 (N_9264,N_6443,N_6679);
nand U9265 (N_9265,N_7716,N_6015);
or U9266 (N_9266,N_7671,N_7919);
or U9267 (N_9267,N_7070,N_7003);
and U9268 (N_9268,N_7138,N_7686);
or U9269 (N_9269,N_7441,N_7956);
and U9270 (N_9270,N_6203,N_6389);
or U9271 (N_9271,N_7476,N_6176);
nor U9272 (N_9272,N_7744,N_7960);
nor U9273 (N_9273,N_6612,N_7970);
nor U9274 (N_9274,N_7502,N_6317);
or U9275 (N_9275,N_6903,N_6762);
nor U9276 (N_9276,N_6994,N_6867);
nor U9277 (N_9277,N_6802,N_6204);
nor U9278 (N_9278,N_6326,N_7962);
xor U9279 (N_9279,N_6244,N_6421);
and U9280 (N_9280,N_7840,N_6141);
nor U9281 (N_9281,N_6908,N_6179);
nand U9282 (N_9282,N_7350,N_7445);
nor U9283 (N_9283,N_7540,N_7378);
nor U9284 (N_9284,N_6376,N_7577);
and U9285 (N_9285,N_6317,N_6440);
or U9286 (N_9286,N_6278,N_6098);
and U9287 (N_9287,N_7348,N_7252);
nor U9288 (N_9288,N_6323,N_7456);
and U9289 (N_9289,N_7633,N_6735);
or U9290 (N_9290,N_6337,N_7313);
nand U9291 (N_9291,N_6354,N_7957);
or U9292 (N_9292,N_7118,N_7874);
or U9293 (N_9293,N_6869,N_6007);
or U9294 (N_9294,N_6997,N_7097);
or U9295 (N_9295,N_6122,N_7526);
or U9296 (N_9296,N_7094,N_7170);
and U9297 (N_9297,N_6327,N_7953);
nor U9298 (N_9298,N_6676,N_7091);
nor U9299 (N_9299,N_7301,N_6017);
or U9300 (N_9300,N_7604,N_7800);
and U9301 (N_9301,N_6147,N_7640);
nand U9302 (N_9302,N_7469,N_6269);
and U9303 (N_9303,N_7816,N_6326);
and U9304 (N_9304,N_7438,N_6197);
xnor U9305 (N_9305,N_6756,N_7413);
nor U9306 (N_9306,N_6128,N_6270);
or U9307 (N_9307,N_6338,N_7772);
and U9308 (N_9308,N_6139,N_6393);
and U9309 (N_9309,N_6314,N_6158);
nand U9310 (N_9310,N_7534,N_6255);
nor U9311 (N_9311,N_6957,N_7182);
and U9312 (N_9312,N_7511,N_6966);
or U9313 (N_9313,N_7577,N_6035);
or U9314 (N_9314,N_6798,N_6128);
nand U9315 (N_9315,N_7487,N_7395);
nand U9316 (N_9316,N_6748,N_7616);
nor U9317 (N_9317,N_7199,N_7631);
or U9318 (N_9318,N_6463,N_7178);
nand U9319 (N_9319,N_6729,N_7799);
nor U9320 (N_9320,N_6550,N_6143);
nand U9321 (N_9321,N_6544,N_6092);
nor U9322 (N_9322,N_6261,N_6373);
or U9323 (N_9323,N_7732,N_6153);
nor U9324 (N_9324,N_7651,N_7832);
and U9325 (N_9325,N_7632,N_6186);
or U9326 (N_9326,N_6677,N_7804);
and U9327 (N_9327,N_6854,N_6836);
nor U9328 (N_9328,N_6596,N_7958);
nor U9329 (N_9329,N_7523,N_7936);
nor U9330 (N_9330,N_6970,N_6760);
nand U9331 (N_9331,N_7886,N_6515);
nor U9332 (N_9332,N_7796,N_6512);
nor U9333 (N_9333,N_6752,N_6036);
nor U9334 (N_9334,N_6767,N_7937);
nand U9335 (N_9335,N_6395,N_7392);
and U9336 (N_9336,N_6335,N_7828);
nand U9337 (N_9337,N_7057,N_6600);
and U9338 (N_9338,N_7366,N_6386);
and U9339 (N_9339,N_6250,N_7756);
nor U9340 (N_9340,N_7933,N_6618);
nand U9341 (N_9341,N_6133,N_6455);
nand U9342 (N_9342,N_7510,N_6526);
nand U9343 (N_9343,N_6717,N_6178);
and U9344 (N_9344,N_6067,N_7325);
nand U9345 (N_9345,N_7257,N_6499);
nor U9346 (N_9346,N_6687,N_7838);
nor U9347 (N_9347,N_6565,N_7062);
nor U9348 (N_9348,N_6760,N_7026);
and U9349 (N_9349,N_6722,N_7843);
nor U9350 (N_9350,N_6196,N_7380);
nor U9351 (N_9351,N_7339,N_6059);
nand U9352 (N_9352,N_6453,N_6066);
nand U9353 (N_9353,N_7870,N_7336);
nor U9354 (N_9354,N_7862,N_7488);
or U9355 (N_9355,N_6069,N_7474);
nand U9356 (N_9356,N_7928,N_7326);
nand U9357 (N_9357,N_7012,N_6390);
nand U9358 (N_9358,N_7780,N_7734);
nand U9359 (N_9359,N_7528,N_7792);
and U9360 (N_9360,N_6624,N_7374);
nor U9361 (N_9361,N_6802,N_6241);
nand U9362 (N_9362,N_7545,N_6248);
and U9363 (N_9363,N_7754,N_6611);
and U9364 (N_9364,N_6892,N_6871);
or U9365 (N_9365,N_7903,N_7692);
nor U9366 (N_9366,N_7343,N_7636);
nand U9367 (N_9367,N_6964,N_6866);
or U9368 (N_9368,N_7880,N_6135);
nor U9369 (N_9369,N_7423,N_7177);
nand U9370 (N_9370,N_6086,N_6717);
nand U9371 (N_9371,N_6769,N_7016);
nor U9372 (N_9372,N_7024,N_7216);
nor U9373 (N_9373,N_6946,N_7360);
nor U9374 (N_9374,N_7145,N_7974);
and U9375 (N_9375,N_6755,N_6848);
or U9376 (N_9376,N_6035,N_6600);
or U9377 (N_9377,N_7509,N_7649);
or U9378 (N_9378,N_7096,N_6508);
nor U9379 (N_9379,N_6165,N_6865);
nor U9380 (N_9380,N_6561,N_6660);
nand U9381 (N_9381,N_6635,N_7270);
and U9382 (N_9382,N_6416,N_6561);
nor U9383 (N_9383,N_7249,N_7209);
nor U9384 (N_9384,N_7429,N_6286);
nor U9385 (N_9385,N_7504,N_6747);
or U9386 (N_9386,N_6412,N_7370);
nor U9387 (N_9387,N_7192,N_7904);
and U9388 (N_9388,N_7442,N_6856);
nor U9389 (N_9389,N_7811,N_6473);
nand U9390 (N_9390,N_7687,N_7142);
or U9391 (N_9391,N_6925,N_7633);
or U9392 (N_9392,N_6175,N_7874);
and U9393 (N_9393,N_6829,N_7774);
nor U9394 (N_9394,N_7795,N_7705);
nor U9395 (N_9395,N_7513,N_7832);
or U9396 (N_9396,N_7933,N_7641);
or U9397 (N_9397,N_6558,N_7905);
and U9398 (N_9398,N_6579,N_7184);
or U9399 (N_9399,N_6632,N_7111);
or U9400 (N_9400,N_6452,N_6545);
and U9401 (N_9401,N_6238,N_7598);
nand U9402 (N_9402,N_7439,N_6575);
nor U9403 (N_9403,N_7324,N_7246);
and U9404 (N_9404,N_6103,N_6170);
nand U9405 (N_9405,N_6782,N_7765);
nor U9406 (N_9406,N_7276,N_7176);
or U9407 (N_9407,N_6411,N_7022);
nand U9408 (N_9408,N_6365,N_7074);
nor U9409 (N_9409,N_6706,N_6391);
nor U9410 (N_9410,N_7389,N_7501);
and U9411 (N_9411,N_6517,N_7543);
and U9412 (N_9412,N_6255,N_6908);
nand U9413 (N_9413,N_7719,N_7583);
and U9414 (N_9414,N_7392,N_6964);
or U9415 (N_9415,N_6683,N_6874);
or U9416 (N_9416,N_7864,N_7392);
nand U9417 (N_9417,N_6567,N_6499);
and U9418 (N_9418,N_6372,N_6770);
nor U9419 (N_9419,N_6359,N_6686);
and U9420 (N_9420,N_7492,N_6496);
and U9421 (N_9421,N_7818,N_6504);
or U9422 (N_9422,N_6394,N_7902);
nor U9423 (N_9423,N_7878,N_6236);
nor U9424 (N_9424,N_7843,N_7181);
nor U9425 (N_9425,N_7325,N_7613);
nand U9426 (N_9426,N_6786,N_7657);
nand U9427 (N_9427,N_6478,N_7097);
and U9428 (N_9428,N_7429,N_7911);
nand U9429 (N_9429,N_6912,N_6252);
and U9430 (N_9430,N_7556,N_7792);
and U9431 (N_9431,N_6064,N_6761);
or U9432 (N_9432,N_6232,N_7167);
and U9433 (N_9433,N_7053,N_6365);
or U9434 (N_9434,N_7180,N_7062);
and U9435 (N_9435,N_7260,N_7629);
nor U9436 (N_9436,N_6079,N_6978);
nor U9437 (N_9437,N_6449,N_6870);
and U9438 (N_9438,N_7485,N_7437);
nand U9439 (N_9439,N_7268,N_6654);
and U9440 (N_9440,N_7185,N_6512);
nand U9441 (N_9441,N_7857,N_6460);
or U9442 (N_9442,N_6293,N_7939);
nor U9443 (N_9443,N_6308,N_6298);
and U9444 (N_9444,N_6958,N_7542);
nand U9445 (N_9445,N_6314,N_6402);
or U9446 (N_9446,N_7906,N_6584);
nand U9447 (N_9447,N_6811,N_7111);
nand U9448 (N_9448,N_7169,N_7283);
and U9449 (N_9449,N_6406,N_6228);
nor U9450 (N_9450,N_6589,N_7750);
and U9451 (N_9451,N_6898,N_6415);
nand U9452 (N_9452,N_7912,N_7058);
nand U9453 (N_9453,N_6134,N_6894);
and U9454 (N_9454,N_7885,N_7679);
and U9455 (N_9455,N_6045,N_6384);
nor U9456 (N_9456,N_6014,N_6215);
and U9457 (N_9457,N_6083,N_7743);
and U9458 (N_9458,N_7078,N_6421);
and U9459 (N_9459,N_7999,N_6823);
nand U9460 (N_9460,N_7424,N_7736);
nand U9461 (N_9461,N_7497,N_6661);
and U9462 (N_9462,N_6245,N_7675);
nor U9463 (N_9463,N_7941,N_7078);
nand U9464 (N_9464,N_7493,N_7333);
and U9465 (N_9465,N_6860,N_6083);
or U9466 (N_9466,N_7743,N_7390);
nor U9467 (N_9467,N_6595,N_6644);
nor U9468 (N_9468,N_6109,N_7345);
and U9469 (N_9469,N_6283,N_6169);
nor U9470 (N_9470,N_6599,N_6615);
or U9471 (N_9471,N_7392,N_7248);
or U9472 (N_9472,N_7941,N_7856);
nor U9473 (N_9473,N_7500,N_6594);
and U9474 (N_9474,N_7803,N_7178);
nor U9475 (N_9475,N_6902,N_7232);
nor U9476 (N_9476,N_6873,N_6672);
nand U9477 (N_9477,N_6061,N_6236);
and U9478 (N_9478,N_6911,N_6902);
or U9479 (N_9479,N_7685,N_6552);
and U9480 (N_9480,N_6251,N_7721);
nand U9481 (N_9481,N_7286,N_7287);
nor U9482 (N_9482,N_6288,N_7611);
nor U9483 (N_9483,N_7027,N_6738);
nand U9484 (N_9484,N_7404,N_7678);
nand U9485 (N_9485,N_7291,N_6328);
and U9486 (N_9486,N_6612,N_7592);
and U9487 (N_9487,N_6685,N_7043);
or U9488 (N_9488,N_6183,N_7691);
or U9489 (N_9489,N_7901,N_6757);
xor U9490 (N_9490,N_6641,N_7064);
nor U9491 (N_9491,N_7936,N_6532);
nand U9492 (N_9492,N_7189,N_6448);
and U9493 (N_9493,N_7251,N_7133);
or U9494 (N_9494,N_7559,N_6972);
or U9495 (N_9495,N_7287,N_6481);
nor U9496 (N_9496,N_6475,N_6926);
and U9497 (N_9497,N_6671,N_7263);
or U9498 (N_9498,N_7705,N_7352);
and U9499 (N_9499,N_7841,N_6221);
nand U9500 (N_9500,N_7266,N_7038);
nor U9501 (N_9501,N_7663,N_6721);
and U9502 (N_9502,N_6733,N_7773);
and U9503 (N_9503,N_7526,N_7292);
nand U9504 (N_9504,N_7230,N_7482);
nor U9505 (N_9505,N_7276,N_6079);
nand U9506 (N_9506,N_6623,N_6624);
nor U9507 (N_9507,N_7295,N_6511);
or U9508 (N_9508,N_6825,N_7340);
nor U9509 (N_9509,N_7037,N_6969);
or U9510 (N_9510,N_6501,N_7604);
or U9511 (N_9511,N_6522,N_7406);
nand U9512 (N_9512,N_6289,N_7234);
and U9513 (N_9513,N_6648,N_7401);
and U9514 (N_9514,N_6777,N_6184);
and U9515 (N_9515,N_6048,N_7344);
nor U9516 (N_9516,N_7372,N_7096);
or U9517 (N_9517,N_6017,N_7259);
nor U9518 (N_9518,N_7362,N_6321);
or U9519 (N_9519,N_7380,N_7407);
nand U9520 (N_9520,N_6298,N_7458);
nor U9521 (N_9521,N_7707,N_6143);
and U9522 (N_9522,N_7320,N_7631);
or U9523 (N_9523,N_6176,N_7181);
or U9524 (N_9524,N_6462,N_6294);
nand U9525 (N_9525,N_7762,N_7947);
nor U9526 (N_9526,N_7295,N_6501);
and U9527 (N_9527,N_7798,N_6854);
nand U9528 (N_9528,N_6606,N_7755);
or U9529 (N_9529,N_6526,N_7654);
and U9530 (N_9530,N_7801,N_6395);
nand U9531 (N_9531,N_6561,N_6677);
nand U9532 (N_9532,N_6472,N_7236);
and U9533 (N_9533,N_6438,N_7221);
nand U9534 (N_9534,N_6759,N_7158);
or U9535 (N_9535,N_7923,N_6609);
nor U9536 (N_9536,N_6275,N_6647);
nand U9537 (N_9537,N_7187,N_7174);
and U9538 (N_9538,N_7140,N_7087);
nand U9539 (N_9539,N_6962,N_7554);
or U9540 (N_9540,N_7906,N_7613);
and U9541 (N_9541,N_6877,N_7742);
nand U9542 (N_9542,N_7273,N_7980);
or U9543 (N_9543,N_7179,N_7805);
nor U9544 (N_9544,N_7476,N_7852);
and U9545 (N_9545,N_6717,N_6312);
nand U9546 (N_9546,N_7370,N_7532);
nand U9547 (N_9547,N_7443,N_6127);
or U9548 (N_9548,N_6212,N_6149);
and U9549 (N_9549,N_7786,N_7455);
nor U9550 (N_9550,N_7558,N_7453);
or U9551 (N_9551,N_6273,N_6923);
nand U9552 (N_9552,N_7009,N_6846);
nand U9553 (N_9553,N_6123,N_7428);
or U9554 (N_9554,N_6514,N_7396);
nand U9555 (N_9555,N_7168,N_6435);
or U9556 (N_9556,N_6241,N_7113);
nand U9557 (N_9557,N_7227,N_6505);
nor U9558 (N_9558,N_6797,N_6669);
and U9559 (N_9559,N_6772,N_7715);
and U9560 (N_9560,N_6248,N_6302);
nand U9561 (N_9561,N_6238,N_6933);
nand U9562 (N_9562,N_7286,N_6668);
or U9563 (N_9563,N_7579,N_7335);
nand U9564 (N_9564,N_7703,N_6101);
or U9565 (N_9565,N_6629,N_6428);
nor U9566 (N_9566,N_7793,N_6930);
nand U9567 (N_9567,N_6683,N_6977);
nand U9568 (N_9568,N_6101,N_7460);
or U9569 (N_9569,N_7625,N_6849);
nor U9570 (N_9570,N_7642,N_7464);
or U9571 (N_9571,N_6378,N_6830);
nand U9572 (N_9572,N_7004,N_7582);
nor U9573 (N_9573,N_7696,N_6034);
and U9574 (N_9574,N_6208,N_6565);
or U9575 (N_9575,N_6214,N_7234);
nand U9576 (N_9576,N_7847,N_7677);
and U9577 (N_9577,N_7620,N_7464);
and U9578 (N_9578,N_6051,N_6340);
or U9579 (N_9579,N_7172,N_6192);
nand U9580 (N_9580,N_7618,N_6706);
and U9581 (N_9581,N_7466,N_6610);
or U9582 (N_9582,N_7327,N_7297);
nand U9583 (N_9583,N_7437,N_7577);
nor U9584 (N_9584,N_6803,N_6337);
nor U9585 (N_9585,N_7615,N_6128);
or U9586 (N_9586,N_7031,N_7131);
nand U9587 (N_9587,N_7632,N_7762);
nor U9588 (N_9588,N_6371,N_6565);
nor U9589 (N_9589,N_6760,N_7841);
and U9590 (N_9590,N_6418,N_6211);
xor U9591 (N_9591,N_7235,N_6487);
nand U9592 (N_9592,N_6338,N_7639);
or U9593 (N_9593,N_6667,N_7041);
and U9594 (N_9594,N_7535,N_6787);
and U9595 (N_9595,N_6260,N_6719);
nand U9596 (N_9596,N_7846,N_6121);
nand U9597 (N_9597,N_7763,N_6927);
or U9598 (N_9598,N_6335,N_6159);
nor U9599 (N_9599,N_6598,N_7570);
nor U9600 (N_9600,N_7937,N_6397);
nand U9601 (N_9601,N_6542,N_7662);
nand U9602 (N_9602,N_6288,N_6432);
or U9603 (N_9603,N_7088,N_6662);
nand U9604 (N_9604,N_6619,N_7980);
nand U9605 (N_9605,N_6621,N_7442);
nand U9606 (N_9606,N_7809,N_6960);
nand U9607 (N_9607,N_7521,N_6120);
or U9608 (N_9608,N_7954,N_7821);
or U9609 (N_9609,N_6401,N_6766);
or U9610 (N_9610,N_7931,N_7849);
nand U9611 (N_9611,N_7053,N_6285);
nand U9612 (N_9612,N_6211,N_7463);
xor U9613 (N_9613,N_6285,N_6538);
xor U9614 (N_9614,N_7566,N_7011);
and U9615 (N_9615,N_7238,N_7059);
nor U9616 (N_9616,N_7232,N_6327);
nor U9617 (N_9617,N_7676,N_6227);
or U9618 (N_9618,N_7995,N_7780);
and U9619 (N_9619,N_7818,N_7922);
or U9620 (N_9620,N_7882,N_6122);
or U9621 (N_9621,N_7009,N_6194);
or U9622 (N_9622,N_7243,N_7956);
nor U9623 (N_9623,N_7736,N_6668);
nand U9624 (N_9624,N_6424,N_7609);
nor U9625 (N_9625,N_6748,N_7543);
nand U9626 (N_9626,N_7977,N_7659);
or U9627 (N_9627,N_6218,N_6311);
nand U9628 (N_9628,N_7453,N_7436);
and U9629 (N_9629,N_7602,N_6661);
or U9630 (N_9630,N_7236,N_7369);
nand U9631 (N_9631,N_7769,N_6160);
or U9632 (N_9632,N_6515,N_6310);
and U9633 (N_9633,N_7638,N_7087);
or U9634 (N_9634,N_7869,N_7674);
nor U9635 (N_9635,N_6696,N_6938);
or U9636 (N_9636,N_7123,N_7184);
nand U9637 (N_9637,N_7533,N_6864);
nand U9638 (N_9638,N_7055,N_6697);
or U9639 (N_9639,N_6065,N_6513);
or U9640 (N_9640,N_6742,N_7063);
and U9641 (N_9641,N_7689,N_7828);
xor U9642 (N_9642,N_6678,N_6257);
or U9643 (N_9643,N_7599,N_7109);
or U9644 (N_9644,N_6564,N_6646);
xor U9645 (N_9645,N_6627,N_6643);
nand U9646 (N_9646,N_6392,N_7672);
or U9647 (N_9647,N_6849,N_7395);
and U9648 (N_9648,N_7354,N_6186);
and U9649 (N_9649,N_6961,N_6308);
or U9650 (N_9650,N_6085,N_6389);
or U9651 (N_9651,N_7256,N_7842);
nand U9652 (N_9652,N_6873,N_7361);
nand U9653 (N_9653,N_7388,N_7077);
nor U9654 (N_9654,N_6105,N_7216);
nor U9655 (N_9655,N_7414,N_7346);
nor U9656 (N_9656,N_7818,N_7816);
or U9657 (N_9657,N_6211,N_7737);
nor U9658 (N_9658,N_6401,N_6488);
nand U9659 (N_9659,N_6506,N_7561);
nor U9660 (N_9660,N_7976,N_7218);
nand U9661 (N_9661,N_6032,N_7193);
or U9662 (N_9662,N_6213,N_6718);
nor U9663 (N_9663,N_6324,N_6370);
nand U9664 (N_9664,N_6533,N_6088);
nor U9665 (N_9665,N_6201,N_7881);
nand U9666 (N_9666,N_6577,N_7124);
nand U9667 (N_9667,N_7487,N_7840);
or U9668 (N_9668,N_6809,N_6374);
nor U9669 (N_9669,N_6835,N_6842);
nand U9670 (N_9670,N_7964,N_7585);
nor U9671 (N_9671,N_7705,N_6651);
and U9672 (N_9672,N_6944,N_6690);
nor U9673 (N_9673,N_7589,N_7147);
or U9674 (N_9674,N_6391,N_7951);
nor U9675 (N_9675,N_6726,N_6941);
and U9676 (N_9676,N_6699,N_7959);
nor U9677 (N_9677,N_6443,N_6567);
or U9678 (N_9678,N_6967,N_7260);
nand U9679 (N_9679,N_7035,N_6155);
nor U9680 (N_9680,N_7311,N_6911);
nor U9681 (N_9681,N_6779,N_6341);
or U9682 (N_9682,N_7718,N_7538);
or U9683 (N_9683,N_6949,N_7245);
nor U9684 (N_9684,N_7116,N_6589);
nor U9685 (N_9685,N_6762,N_6067);
and U9686 (N_9686,N_6156,N_6774);
and U9687 (N_9687,N_6845,N_7958);
or U9688 (N_9688,N_7674,N_7950);
or U9689 (N_9689,N_6910,N_7328);
nand U9690 (N_9690,N_6270,N_7418);
or U9691 (N_9691,N_6435,N_6943);
nand U9692 (N_9692,N_6429,N_7459);
nor U9693 (N_9693,N_7470,N_7823);
and U9694 (N_9694,N_6255,N_7610);
or U9695 (N_9695,N_6517,N_6999);
or U9696 (N_9696,N_6460,N_6511);
nand U9697 (N_9697,N_6833,N_6577);
nand U9698 (N_9698,N_6595,N_6818);
or U9699 (N_9699,N_6354,N_7802);
or U9700 (N_9700,N_7972,N_6589);
nand U9701 (N_9701,N_7246,N_7549);
nor U9702 (N_9702,N_6392,N_6601);
and U9703 (N_9703,N_6581,N_6768);
and U9704 (N_9704,N_6870,N_6736);
and U9705 (N_9705,N_7856,N_7418);
or U9706 (N_9706,N_6564,N_7437);
nand U9707 (N_9707,N_6771,N_6483);
xor U9708 (N_9708,N_7717,N_6348);
and U9709 (N_9709,N_7476,N_7666);
nand U9710 (N_9710,N_6338,N_6337);
and U9711 (N_9711,N_7796,N_7637);
nand U9712 (N_9712,N_7683,N_6120);
or U9713 (N_9713,N_6682,N_6217);
and U9714 (N_9714,N_6720,N_7360);
nand U9715 (N_9715,N_6833,N_7947);
nor U9716 (N_9716,N_6546,N_6886);
nor U9717 (N_9717,N_6980,N_6482);
and U9718 (N_9718,N_6075,N_7434);
and U9719 (N_9719,N_7326,N_7009);
and U9720 (N_9720,N_7870,N_7337);
and U9721 (N_9721,N_7204,N_6330);
nand U9722 (N_9722,N_7862,N_7741);
or U9723 (N_9723,N_7654,N_7643);
nor U9724 (N_9724,N_6401,N_7282);
nor U9725 (N_9725,N_6757,N_7347);
nand U9726 (N_9726,N_7790,N_6089);
nor U9727 (N_9727,N_7417,N_7858);
or U9728 (N_9728,N_6437,N_7774);
or U9729 (N_9729,N_6346,N_6269);
nor U9730 (N_9730,N_7730,N_7415);
and U9731 (N_9731,N_7434,N_7833);
nor U9732 (N_9732,N_6875,N_7266);
nor U9733 (N_9733,N_6841,N_7106);
and U9734 (N_9734,N_6736,N_7321);
nand U9735 (N_9735,N_7607,N_7031);
or U9736 (N_9736,N_7462,N_6483);
nor U9737 (N_9737,N_6245,N_7631);
and U9738 (N_9738,N_6101,N_6140);
and U9739 (N_9739,N_7740,N_6497);
and U9740 (N_9740,N_7414,N_7039);
nor U9741 (N_9741,N_7657,N_6751);
or U9742 (N_9742,N_7169,N_6362);
nor U9743 (N_9743,N_7144,N_6495);
or U9744 (N_9744,N_7732,N_6578);
and U9745 (N_9745,N_6217,N_6949);
nand U9746 (N_9746,N_6091,N_7295);
nor U9747 (N_9747,N_7001,N_7198);
nand U9748 (N_9748,N_7590,N_6220);
nor U9749 (N_9749,N_6932,N_7498);
nor U9750 (N_9750,N_6011,N_6706);
nand U9751 (N_9751,N_6009,N_7190);
nand U9752 (N_9752,N_6930,N_6730);
or U9753 (N_9753,N_7648,N_6300);
nand U9754 (N_9754,N_7215,N_6929);
nor U9755 (N_9755,N_7237,N_7981);
nor U9756 (N_9756,N_6144,N_7405);
or U9757 (N_9757,N_6949,N_7414);
nand U9758 (N_9758,N_7731,N_6207);
nor U9759 (N_9759,N_6688,N_6888);
nor U9760 (N_9760,N_6235,N_6078);
nor U9761 (N_9761,N_6620,N_7313);
and U9762 (N_9762,N_7524,N_6059);
and U9763 (N_9763,N_7623,N_7856);
nand U9764 (N_9764,N_6032,N_7839);
nor U9765 (N_9765,N_7095,N_6990);
nor U9766 (N_9766,N_6768,N_6618);
nor U9767 (N_9767,N_7983,N_6139);
or U9768 (N_9768,N_7744,N_6919);
nand U9769 (N_9769,N_6106,N_7410);
nor U9770 (N_9770,N_6099,N_7202);
nand U9771 (N_9771,N_7037,N_6561);
and U9772 (N_9772,N_6415,N_6207);
and U9773 (N_9773,N_6049,N_7737);
or U9774 (N_9774,N_7308,N_7384);
and U9775 (N_9775,N_7488,N_6306);
or U9776 (N_9776,N_7480,N_7836);
nand U9777 (N_9777,N_6775,N_6446);
and U9778 (N_9778,N_6128,N_6624);
or U9779 (N_9779,N_7201,N_6592);
and U9780 (N_9780,N_6651,N_6879);
nand U9781 (N_9781,N_6812,N_6787);
or U9782 (N_9782,N_7750,N_6175);
nand U9783 (N_9783,N_6329,N_6757);
or U9784 (N_9784,N_6314,N_7382);
or U9785 (N_9785,N_6870,N_7207);
nand U9786 (N_9786,N_6544,N_7818);
or U9787 (N_9787,N_7632,N_6331);
and U9788 (N_9788,N_7165,N_7839);
nor U9789 (N_9789,N_7062,N_6043);
and U9790 (N_9790,N_6932,N_6557);
nand U9791 (N_9791,N_6775,N_6810);
or U9792 (N_9792,N_7181,N_7553);
and U9793 (N_9793,N_7748,N_6183);
and U9794 (N_9794,N_6154,N_7121);
nand U9795 (N_9795,N_6170,N_6784);
or U9796 (N_9796,N_6289,N_7379);
or U9797 (N_9797,N_6474,N_6071);
or U9798 (N_9798,N_7961,N_6593);
nand U9799 (N_9799,N_7888,N_6583);
or U9800 (N_9800,N_6144,N_7912);
nand U9801 (N_9801,N_6297,N_7497);
nand U9802 (N_9802,N_6870,N_6360);
nand U9803 (N_9803,N_7157,N_7512);
and U9804 (N_9804,N_7409,N_7889);
or U9805 (N_9805,N_6933,N_7825);
and U9806 (N_9806,N_6445,N_7944);
or U9807 (N_9807,N_7476,N_7339);
nand U9808 (N_9808,N_7654,N_7876);
nor U9809 (N_9809,N_7271,N_7286);
nand U9810 (N_9810,N_6851,N_7074);
and U9811 (N_9811,N_6108,N_6819);
nand U9812 (N_9812,N_7751,N_6740);
and U9813 (N_9813,N_6439,N_6307);
nor U9814 (N_9814,N_6359,N_7980);
nor U9815 (N_9815,N_7938,N_6987);
nand U9816 (N_9816,N_6544,N_6442);
or U9817 (N_9817,N_6082,N_6323);
nand U9818 (N_9818,N_6278,N_7487);
nor U9819 (N_9819,N_6851,N_7860);
and U9820 (N_9820,N_6975,N_6108);
or U9821 (N_9821,N_6714,N_7472);
nand U9822 (N_9822,N_7060,N_6456);
and U9823 (N_9823,N_6658,N_7062);
nand U9824 (N_9824,N_7245,N_6205);
nand U9825 (N_9825,N_6379,N_7901);
or U9826 (N_9826,N_6359,N_6010);
and U9827 (N_9827,N_6232,N_7418);
or U9828 (N_9828,N_7829,N_7917);
or U9829 (N_9829,N_6717,N_6614);
and U9830 (N_9830,N_7529,N_6505);
or U9831 (N_9831,N_6667,N_7648);
nor U9832 (N_9832,N_6628,N_7631);
nand U9833 (N_9833,N_6697,N_7738);
or U9834 (N_9834,N_6542,N_6394);
and U9835 (N_9835,N_6366,N_6970);
and U9836 (N_9836,N_7487,N_6762);
and U9837 (N_9837,N_6913,N_6333);
or U9838 (N_9838,N_6815,N_7243);
and U9839 (N_9839,N_7848,N_7065);
nand U9840 (N_9840,N_6736,N_6029);
and U9841 (N_9841,N_6116,N_6692);
nand U9842 (N_9842,N_6049,N_6178);
nor U9843 (N_9843,N_7338,N_6705);
nand U9844 (N_9844,N_7464,N_7867);
nand U9845 (N_9845,N_7036,N_7503);
xor U9846 (N_9846,N_7767,N_6851);
nor U9847 (N_9847,N_6912,N_7543);
nand U9848 (N_9848,N_6153,N_6336);
or U9849 (N_9849,N_6688,N_7221);
and U9850 (N_9850,N_6211,N_7186);
nand U9851 (N_9851,N_6818,N_7211);
or U9852 (N_9852,N_6077,N_6382);
and U9853 (N_9853,N_6032,N_7620);
and U9854 (N_9854,N_6908,N_7594);
nand U9855 (N_9855,N_7918,N_7134);
nor U9856 (N_9856,N_6167,N_7556);
and U9857 (N_9857,N_7239,N_7250);
nand U9858 (N_9858,N_6288,N_6363);
nand U9859 (N_9859,N_6133,N_7723);
and U9860 (N_9860,N_6074,N_7974);
nor U9861 (N_9861,N_7102,N_7052);
and U9862 (N_9862,N_7084,N_7752);
or U9863 (N_9863,N_6817,N_7151);
or U9864 (N_9864,N_7698,N_6892);
and U9865 (N_9865,N_7655,N_7441);
nor U9866 (N_9866,N_7592,N_6243);
or U9867 (N_9867,N_6802,N_6912);
nor U9868 (N_9868,N_6631,N_6848);
nand U9869 (N_9869,N_6619,N_7317);
or U9870 (N_9870,N_6420,N_7942);
nand U9871 (N_9871,N_7748,N_6410);
nor U9872 (N_9872,N_6313,N_7556);
nand U9873 (N_9873,N_6669,N_7578);
and U9874 (N_9874,N_7769,N_6155);
nor U9875 (N_9875,N_6968,N_7791);
nand U9876 (N_9876,N_7395,N_6769);
or U9877 (N_9877,N_6055,N_6327);
or U9878 (N_9878,N_6001,N_6557);
nor U9879 (N_9879,N_6808,N_7424);
nor U9880 (N_9880,N_7214,N_6756);
and U9881 (N_9881,N_6613,N_6183);
nand U9882 (N_9882,N_7050,N_7639);
nor U9883 (N_9883,N_6468,N_6388);
and U9884 (N_9884,N_7753,N_6115);
nor U9885 (N_9885,N_6190,N_6352);
and U9886 (N_9886,N_6050,N_6468);
xor U9887 (N_9887,N_6964,N_7543);
and U9888 (N_9888,N_7334,N_7590);
or U9889 (N_9889,N_6967,N_6533);
nor U9890 (N_9890,N_6487,N_7536);
or U9891 (N_9891,N_6614,N_7258);
and U9892 (N_9892,N_7933,N_7036);
or U9893 (N_9893,N_7758,N_6008);
or U9894 (N_9894,N_6245,N_6809);
or U9895 (N_9895,N_7120,N_6452);
nand U9896 (N_9896,N_6614,N_7400);
nor U9897 (N_9897,N_6245,N_7517);
nor U9898 (N_9898,N_7902,N_6368);
nor U9899 (N_9899,N_6117,N_6780);
nand U9900 (N_9900,N_6717,N_6090);
nor U9901 (N_9901,N_7770,N_6408);
and U9902 (N_9902,N_6471,N_7942);
and U9903 (N_9903,N_7770,N_6353);
or U9904 (N_9904,N_7628,N_6341);
or U9905 (N_9905,N_6924,N_7248);
nand U9906 (N_9906,N_6953,N_6881);
nand U9907 (N_9907,N_6716,N_7911);
and U9908 (N_9908,N_7033,N_7567);
nor U9909 (N_9909,N_6703,N_7091);
nor U9910 (N_9910,N_7533,N_7017);
and U9911 (N_9911,N_7411,N_7772);
nand U9912 (N_9912,N_7483,N_7173);
and U9913 (N_9913,N_7293,N_6037);
nor U9914 (N_9914,N_7652,N_6256);
nor U9915 (N_9915,N_7663,N_6085);
and U9916 (N_9916,N_7761,N_7498);
nor U9917 (N_9917,N_7117,N_6861);
nor U9918 (N_9918,N_6912,N_6281);
and U9919 (N_9919,N_6879,N_7732);
nand U9920 (N_9920,N_7814,N_6115);
nand U9921 (N_9921,N_7566,N_6244);
or U9922 (N_9922,N_7978,N_7130);
xor U9923 (N_9923,N_7519,N_7445);
or U9924 (N_9924,N_7923,N_6446);
nor U9925 (N_9925,N_7951,N_7567);
or U9926 (N_9926,N_7292,N_6451);
or U9927 (N_9927,N_6249,N_7579);
nand U9928 (N_9928,N_6553,N_7086);
and U9929 (N_9929,N_7609,N_7523);
nor U9930 (N_9930,N_7470,N_6945);
or U9931 (N_9931,N_7386,N_7117);
and U9932 (N_9932,N_7065,N_7458);
and U9933 (N_9933,N_7323,N_7506);
nor U9934 (N_9934,N_6697,N_7329);
nor U9935 (N_9935,N_6220,N_7173);
nor U9936 (N_9936,N_6891,N_7594);
nand U9937 (N_9937,N_7758,N_7710);
or U9938 (N_9938,N_6487,N_6235);
nor U9939 (N_9939,N_6467,N_6113);
or U9940 (N_9940,N_7423,N_7971);
or U9941 (N_9941,N_6547,N_7398);
or U9942 (N_9942,N_6926,N_7000);
nor U9943 (N_9943,N_6738,N_6214);
or U9944 (N_9944,N_6582,N_7666);
and U9945 (N_9945,N_7153,N_6981);
nand U9946 (N_9946,N_7645,N_6487);
and U9947 (N_9947,N_6529,N_7911);
and U9948 (N_9948,N_7741,N_6791);
and U9949 (N_9949,N_7998,N_7393);
nand U9950 (N_9950,N_6104,N_7031);
or U9951 (N_9951,N_7847,N_6988);
nor U9952 (N_9952,N_6754,N_7913);
and U9953 (N_9953,N_7620,N_6124);
or U9954 (N_9954,N_6547,N_7204);
and U9955 (N_9955,N_6928,N_7679);
and U9956 (N_9956,N_6795,N_6327);
or U9957 (N_9957,N_6076,N_7262);
and U9958 (N_9958,N_7098,N_7275);
and U9959 (N_9959,N_7663,N_7595);
xor U9960 (N_9960,N_6306,N_7024);
or U9961 (N_9961,N_7709,N_6970);
nand U9962 (N_9962,N_6170,N_6071);
and U9963 (N_9963,N_7121,N_6903);
and U9964 (N_9964,N_7707,N_6203);
and U9965 (N_9965,N_7988,N_7230);
nand U9966 (N_9966,N_6531,N_7586);
nor U9967 (N_9967,N_6950,N_6621);
nand U9968 (N_9968,N_6238,N_6267);
nor U9969 (N_9969,N_7480,N_6807);
nor U9970 (N_9970,N_7990,N_7291);
nor U9971 (N_9971,N_7153,N_7660);
and U9972 (N_9972,N_7585,N_7419);
and U9973 (N_9973,N_6085,N_7828);
nand U9974 (N_9974,N_6989,N_6683);
or U9975 (N_9975,N_7990,N_6895);
nor U9976 (N_9976,N_7371,N_7872);
nand U9977 (N_9977,N_6247,N_6350);
nand U9978 (N_9978,N_6117,N_6790);
nor U9979 (N_9979,N_7166,N_6866);
and U9980 (N_9980,N_6699,N_6028);
or U9981 (N_9981,N_7517,N_6903);
and U9982 (N_9982,N_6468,N_6877);
nor U9983 (N_9983,N_7468,N_7023);
xor U9984 (N_9984,N_7955,N_7596);
or U9985 (N_9985,N_6349,N_7825);
nand U9986 (N_9986,N_6133,N_6773);
and U9987 (N_9987,N_6023,N_6919);
nor U9988 (N_9988,N_6938,N_6205);
nand U9989 (N_9989,N_6916,N_7814);
or U9990 (N_9990,N_7482,N_6109);
and U9991 (N_9991,N_7983,N_6674);
or U9992 (N_9992,N_7050,N_6421);
and U9993 (N_9993,N_6868,N_6904);
or U9994 (N_9994,N_7497,N_6200);
or U9995 (N_9995,N_7301,N_6440);
nand U9996 (N_9996,N_6117,N_7497);
nand U9997 (N_9997,N_6988,N_7483);
and U9998 (N_9998,N_6745,N_6175);
and U9999 (N_9999,N_6639,N_6348);
nand UO_0 (O_0,N_9602,N_9372);
and UO_1 (O_1,N_9288,N_8002);
or UO_2 (O_2,N_9180,N_8148);
or UO_3 (O_3,N_8205,N_8299);
and UO_4 (O_4,N_9743,N_8894);
nand UO_5 (O_5,N_8848,N_8158);
nand UO_6 (O_6,N_8572,N_8619);
and UO_7 (O_7,N_8945,N_8783);
and UO_8 (O_8,N_9851,N_8365);
nand UO_9 (O_9,N_9244,N_8076);
and UO_10 (O_10,N_9974,N_8310);
nor UO_11 (O_11,N_9558,N_8962);
and UO_12 (O_12,N_8160,N_8041);
xor UO_13 (O_13,N_9616,N_8057);
and UO_14 (O_14,N_9381,N_9234);
xor UO_15 (O_15,N_9487,N_8346);
or UO_16 (O_16,N_9919,N_9702);
or UO_17 (O_17,N_9018,N_9146);
nand UO_18 (O_18,N_9511,N_9868);
nand UO_19 (O_19,N_8523,N_8879);
and UO_20 (O_20,N_9296,N_8765);
nor UO_21 (O_21,N_9029,N_8941);
or UO_22 (O_22,N_9502,N_9371);
nand UO_23 (O_23,N_9541,N_9827);
or UO_24 (O_24,N_8627,N_9960);
nor UO_25 (O_25,N_8430,N_9788);
nor UO_26 (O_26,N_8670,N_9658);
nor UO_27 (O_27,N_8254,N_9102);
or UO_28 (O_28,N_9025,N_9678);
nor UO_29 (O_29,N_9545,N_9193);
nor UO_30 (O_30,N_8987,N_8729);
nor UO_31 (O_31,N_8671,N_9747);
and UO_32 (O_32,N_8676,N_8394);
and UO_33 (O_33,N_8469,N_9218);
nand UO_34 (O_34,N_9028,N_8610);
or UO_35 (O_35,N_9284,N_8015);
nand UO_36 (O_36,N_9515,N_8668);
nand UO_37 (O_37,N_9145,N_8171);
or UO_38 (O_38,N_8323,N_8536);
and UO_39 (O_39,N_9829,N_8681);
nand UO_40 (O_40,N_8471,N_9256);
and UO_41 (O_41,N_8716,N_8935);
nor UO_42 (O_42,N_8123,N_8480);
or UO_43 (O_43,N_9049,N_9163);
and UO_44 (O_44,N_8781,N_9937);
and UO_45 (O_45,N_8808,N_9473);
nand UO_46 (O_46,N_8195,N_8747);
or UO_47 (O_47,N_8576,N_9358);
nand UO_48 (O_48,N_9113,N_8278);
nor UO_49 (O_49,N_8376,N_8180);
nor UO_50 (O_50,N_9855,N_9507);
and UO_51 (O_51,N_8155,N_9043);
nand UO_52 (O_52,N_8340,N_8784);
nand UO_53 (O_53,N_9273,N_8512);
or UO_54 (O_54,N_9807,N_8801);
and UO_55 (O_55,N_9073,N_8897);
nor UO_56 (O_56,N_9739,N_9362);
nor UO_57 (O_57,N_8181,N_8882);
nand UO_58 (O_58,N_9825,N_8521);
and UO_59 (O_59,N_8113,N_9056);
and UO_60 (O_60,N_8886,N_9260);
and UO_61 (O_61,N_8359,N_9436);
and UO_62 (O_62,N_8549,N_8895);
nor UO_63 (O_63,N_8048,N_8552);
and UO_64 (O_64,N_8168,N_8728);
or UO_65 (O_65,N_9012,N_8199);
and UO_66 (O_66,N_9875,N_9732);
and UO_67 (O_67,N_8033,N_9759);
and UO_68 (O_68,N_9742,N_9482);
nor UO_69 (O_69,N_9815,N_9217);
nor UO_70 (O_70,N_9725,N_8562);
or UO_71 (O_71,N_8485,N_9166);
and UO_72 (O_72,N_9513,N_8596);
and UO_73 (O_73,N_9715,N_8734);
nor UO_74 (O_74,N_8755,N_8134);
and UO_75 (O_75,N_8042,N_9258);
or UO_76 (O_76,N_8216,N_9533);
or UO_77 (O_77,N_8061,N_9944);
nor UO_78 (O_78,N_8994,N_9156);
or UO_79 (O_79,N_8253,N_9448);
nand UO_80 (O_80,N_9719,N_8289);
or UO_81 (O_81,N_9740,N_8046);
nor UO_82 (O_82,N_8114,N_8420);
nor UO_83 (O_83,N_9775,N_9434);
and UO_84 (O_84,N_8331,N_9453);
nor UO_85 (O_85,N_8255,N_8878);
xnor UO_86 (O_86,N_9345,N_8145);
nor UO_87 (O_87,N_8974,N_8900);
and UO_88 (O_88,N_9925,N_8256);
nor UO_89 (O_89,N_8178,N_8482);
and UO_90 (O_90,N_8782,N_8544);
nand UO_91 (O_91,N_8044,N_8099);
nor UO_92 (O_92,N_9294,N_8301);
or UO_93 (O_93,N_9538,N_9312);
and UO_94 (O_94,N_9017,N_9269);
and UO_95 (O_95,N_8788,N_8964);
nor UO_96 (O_96,N_8581,N_9069);
nor UO_97 (O_97,N_8504,N_8856);
nor UO_98 (O_98,N_8029,N_9174);
or UO_99 (O_99,N_9540,N_8957);
nand UO_100 (O_100,N_8337,N_8436);
nor UO_101 (O_101,N_9902,N_9873);
nand UO_102 (O_102,N_8481,N_8919);
and UO_103 (O_103,N_8858,N_9886);
xnor UO_104 (O_104,N_9036,N_9070);
and UO_105 (O_105,N_8679,N_8266);
nand UO_106 (O_106,N_9407,N_8628);
nand UO_107 (O_107,N_9491,N_8131);
nor UO_108 (O_108,N_8021,N_8689);
nand UO_109 (O_109,N_8890,N_8772);
nor UO_110 (O_110,N_8785,N_9058);
nor UO_111 (O_111,N_8335,N_8379);
and UO_112 (O_112,N_8970,N_9211);
nand UO_113 (O_113,N_9741,N_9891);
nand UO_114 (O_114,N_9813,N_8479);
nand UO_115 (O_115,N_9999,N_9626);
or UO_116 (O_116,N_8972,N_8675);
nand UO_117 (O_117,N_8413,N_9645);
and UO_118 (O_118,N_9749,N_8857);
nor UO_119 (O_119,N_8654,N_9190);
nand UO_120 (O_120,N_8590,N_8949);
nor UO_121 (O_121,N_9450,N_9782);
nor UO_122 (O_122,N_8938,N_8827);
nor UO_123 (O_123,N_9208,N_9941);
nor UO_124 (O_124,N_9410,N_9798);
nor UO_125 (O_125,N_8718,N_8130);
nand UO_126 (O_126,N_8956,N_9054);
and UO_127 (O_127,N_8012,N_9561);
or UO_128 (O_128,N_9920,N_9975);
nor UO_129 (O_129,N_9657,N_9554);
and UO_130 (O_130,N_9360,N_8170);
and UO_131 (O_131,N_9903,N_8090);
nand UO_132 (O_132,N_9750,N_9659);
nand UO_133 (O_133,N_8969,N_8796);
nor UO_134 (O_134,N_8548,N_9006);
and UO_135 (O_135,N_9066,N_9929);
or UO_136 (O_136,N_9245,N_8721);
or UO_137 (O_137,N_8906,N_9316);
or UO_138 (O_138,N_8532,N_8460);
or UO_139 (O_139,N_8704,N_9132);
and UO_140 (O_140,N_8022,N_9323);
nand UO_141 (O_141,N_9774,N_9213);
nand UO_142 (O_142,N_8226,N_8363);
and UO_143 (O_143,N_9283,N_8541);
xnor UO_144 (O_144,N_9789,N_9388);
nor UO_145 (O_145,N_9641,N_9990);
nand UO_146 (O_146,N_8898,N_9050);
or UO_147 (O_147,N_9871,N_9035);
nor UO_148 (O_148,N_9821,N_8214);
nor UO_149 (O_149,N_9267,N_8739);
nor UO_150 (O_150,N_9475,N_8443);
nand UO_151 (O_151,N_8708,N_8334);
and UO_152 (O_152,N_9397,N_8140);
nor UO_153 (O_153,N_9246,N_9162);
nand UO_154 (O_154,N_9948,N_9242);
and UO_155 (O_155,N_9022,N_8494);
nor UO_156 (O_156,N_9860,N_8595);
nand UO_157 (O_157,N_9693,N_8756);
nor UO_158 (O_158,N_9441,N_8837);
nand UO_159 (O_159,N_8725,N_8092);
and UO_160 (O_160,N_9897,N_9008);
or UO_161 (O_161,N_9562,N_8866);
or UO_162 (O_162,N_8304,N_8281);
or UO_163 (O_163,N_9298,N_8865);
xnor UO_164 (O_164,N_9781,N_8792);
and UO_165 (O_165,N_9128,N_8556);
and UO_166 (O_166,N_9623,N_8237);
nor UO_167 (O_167,N_8010,N_8311);
nand UO_168 (O_168,N_8509,N_8003);
and UO_169 (O_169,N_9326,N_8881);
and UO_170 (O_170,N_8585,N_8350);
or UO_171 (O_171,N_9342,N_9532);
nor UO_172 (O_172,N_9062,N_9007);
and UO_173 (O_173,N_8356,N_8613);
or UO_174 (O_174,N_8682,N_8292);
nor UO_175 (O_175,N_9292,N_9227);
or UO_176 (O_176,N_8832,N_9764);
and UO_177 (O_177,N_9539,N_8876);
and UO_178 (O_178,N_8269,N_9862);
nor UO_179 (O_179,N_9885,N_9276);
and UO_180 (O_180,N_9431,N_8317);
nor UO_181 (O_181,N_9148,N_8518);
or UO_182 (O_182,N_8007,N_8799);
nand UO_183 (O_183,N_8452,N_9464);
and UO_184 (O_184,N_8445,N_8766);
nand UO_185 (O_185,N_9060,N_8902);
and UO_186 (O_186,N_8014,N_9013);
or UO_187 (O_187,N_9463,N_9998);
nor UO_188 (O_188,N_8825,N_9640);
and UO_189 (O_189,N_9557,N_9186);
nor UO_190 (O_190,N_8179,N_8789);
xnor UO_191 (O_191,N_8603,N_8844);
and UO_192 (O_192,N_9355,N_8803);
nand UO_193 (O_193,N_9026,N_8667);
or UO_194 (O_194,N_8072,N_8446);
and UO_195 (O_195,N_8280,N_9906);
nand UO_196 (O_196,N_9385,N_9194);
and UO_197 (O_197,N_8868,N_9196);
and UO_198 (O_198,N_8745,N_8615);
and UO_199 (O_199,N_8024,N_9956);
nand UO_200 (O_200,N_9814,N_9876);
and UO_201 (O_201,N_8045,N_9926);
nand UO_202 (O_202,N_8558,N_9403);
nor UO_203 (O_203,N_9783,N_8241);
nand UO_204 (O_204,N_9714,N_8129);
nor UO_205 (O_205,N_9380,N_9164);
or UO_206 (O_206,N_8203,N_8508);
nand UO_207 (O_207,N_9223,N_9248);
or UO_208 (O_208,N_8979,N_8672);
or UO_209 (O_209,N_8620,N_8539);
or UO_210 (O_210,N_9842,N_8923);
nor UO_211 (O_211,N_8475,N_8580);
nand UO_212 (O_212,N_9934,N_9099);
nand UO_213 (O_213,N_9843,N_9184);
nand UO_214 (O_214,N_8490,N_8319);
or UO_215 (O_215,N_8638,N_9303);
and UO_216 (O_216,N_8498,N_9176);
and UO_217 (O_217,N_9157,N_9278);
or UO_218 (O_218,N_9263,N_9953);
nand UO_219 (O_219,N_8678,N_8247);
nand UO_220 (O_220,N_8273,N_9898);
or UO_221 (O_221,N_9824,N_8097);
nand UO_222 (O_222,N_8493,N_9905);
and UO_223 (O_223,N_8710,N_9845);
nand UO_224 (O_224,N_9527,N_8393);
nand UO_225 (O_225,N_8488,N_9044);
nor UO_226 (O_226,N_9212,N_9422);
or UO_227 (O_227,N_9080,N_8373);
and UO_228 (O_228,N_8954,N_9899);
and UO_229 (O_229,N_9187,N_9675);
and UO_230 (O_230,N_8196,N_9155);
nor UO_231 (O_231,N_8946,N_9496);
nor UO_232 (O_232,N_8978,N_9379);
and UO_233 (O_233,N_8860,N_8143);
and UO_234 (O_234,N_8149,N_9467);
nor UO_235 (O_235,N_9247,N_9405);
nor UO_236 (O_236,N_8248,N_9309);
and UO_237 (O_237,N_8074,N_8732);
and UO_238 (O_238,N_8983,N_9993);
nor UO_239 (O_239,N_9266,N_8221);
nand UO_240 (O_240,N_9904,N_9404);
or UO_241 (O_241,N_8843,N_8395);
and UO_242 (O_242,N_8065,N_9858);
or UO_243 (O_243,N_8391,N_9817);
nor UO_244 (O_244,N_8028,N_9852);
nand UO_245 (O_245,N_9343,N_9844);
nor UO_246 (O_246,N_8588,N_9231);
or UO_247 (O_247,N_8757,N_9964);
or UO_248 (O_248,N_8940,N_8167);
nor UO_249 (O_249,N_9887,N_8333);
or UO_250 (O_250,N_9230,N_8050);
nor UO_251 (O_251,N_9350,N_9680);
nand UO_252 (O_252,N_8648,N_8545);
and UO_253 (O_253,N_8584,N_9220);
nand UO_254 (O_254,N_9888,N_8934);
or UO_255 (O_255,N_9650,N_8736);
nand UO_256 (O_256,N_9074,N_8250);
or UO_257 (O_257,N_9610,N_9285);
or UO_258 (O_258,N_9786,N_9517);
and UO_259 (O_259,N_9427,N_8093);
nor UO_260 (O_260,N_8327,N_8067);
and UO_261 (O_261,N_8016,N_8998);
and UO_262 (O_262,N_9712,N_9052);
nand UO_263 (O_263,N_8368,N_9133);
nor UO_264 (O_264,N_9051,N_8125);
and UO_265 (O_265,N_9098,N_8174);
nand UO_266 (O_266,N_9598,N_8727);
nor UO_267 (O_267,N_8230,N_8606);
nand UO_268 (O_268,N_9793,N_9976);
nand UO_269 (O_269,N_8371,N_8798);
nand UO_270 (O_270,N_8101,N_8888);
nor UO_271 (O_271,N_9563,N_9981);
nor UO_272 (O_272,N_9553,N_8884);
nand UO_273 (O_273,N_8840,N_9861);
and UO_274 (O_274,N_9512,N_8288);
or UO_275 (O_275,N_9571,N_9762);
or UO_276 (O_276,N_9606,N_9794);
xnor UO_277 (O_277,N_8328,N_9255);
or UO_278 (O_278,N_9418,N_9818);
nor UO_279 (O_279,N_8666,N_9141);
or UO_280 (O_280,N_9688,N_8794);
and UO_281 (O_281,N_9462,N_9895);
nand UO_282 (O_282,N_9978,N_8980);
nand UO_283 (O_283,N_8828,N_8127);
or UO_284 (O_284,N_8818,N_8064);
nand UO_285 (O_285,N_9315,N_8569);
or UO_286 (O_286,N_8950,N_9093);
nor UO_287 (O_287,N_9810,N_8385);
nand UO_288 (O_288,N_8960,N_8116);
nand UO_289 (O_289,N_9546,N_8054);
nand UO_290 (O_290,N_9210,N_8849);
nand UO_291 (O_291,N_8661,N_8444);
nand UO_292 (O_292,N_9081,N_8431);
and UO_293 (O_293,N_8455,N_9711);
and UO_294 (O_294,N_9932,N_8939);
nor UO_295 (O_295,N_9836,N_9279);
nor UO_296 (O_296,N_9835,N_8753);
nand UO_297 (O_297,N_9850,N_9703);
nand UO_298 (O_298,N_8822,N_9632);
and UO_299 (O_299,N_8202,N_9116);
nand UO_300 (O_300,N_9763,N_8187);
or UO_301 (O_301,N_8075,N_8663);
nand UO_302 (O_302,N_8624,N_8000);
or UO_303 (O_303,N_8309,N_8709);
or UO_304 (O_304,N_8147,N_8448);
nor UO_305 (O_305,N_9947,N_8403);
nor UO_306 (O_306,N_9795,N_9530);
and UO_307 (O_307,N_8733,N_8953);
and UO_308 (O_308,N_8920,N_8662);
nor UO_309 (O_309,N_9499,N_8501);
and UO_310 (O_310,N_9236,N_9391);
or UO_311 (O_311,N_8107,N_8870);
or UO_312 (O_312,N_9301,N_8495);
or UO_313 (O_313,N_8903,N_9444);
and UO_314 (O_314,N_8622,N_8514);
and UO_315 (O_315,N_8405,N_9869);
and UO_316 (O_316,N_9311,N_8457);
nand UO_317 (O_317,N_8239,N_9199);
nor UO_318 (O_318,N_8397,N_9100);
or UO_319 (O_319,N_8813,N_9957);
nand UO_320 (O_320,N_8804,N_8108);
nand UO_321 (O_321,N_9289,N_8749);
nor UO_322 (O_322,N_8821,N_8396);
nor UO_323 (O_323,N_9585,N_8573);
nor UO_324 (O_324,N_8565,N_9476);
and UO_325 (O_325,N_8916,N_8973);
nor UO_326 (O_326,N_9572,N_8197);
or UO_327 (O_327,N_8816,N_9834);
or UO_328 (O_328,N_9030,N_8442);
nand UO_329 (O_329,N_8102,N_8823);
nand UO_330 (O_330,N_8850,N_9609);
or UO_331 (O_331,N_9175,N_8451);
and UO_332 (O_332,N_9596,N_8347);
nor UO_333 (O_333,N_8218,N_9037);
nor UO_334 (O_334,N_9129,N_8246);
nand UO_335 (O_335,N_9647,N_9587);
nor UO_336 (O_336,N_8871,N_9819);
or UO_337 (O_337,N_8758,N_8971);
nand UO_338 (O_338,N_8128,N_9314);
nand UO_339 (O_339,N_8612,N_8705);
and UO_340 (O_340,N_9357,N_8811);
and UO_341 (O_341,N_9617,N_8831);
nor UO_342 (O_342,N_8060,N_8302);
nand UO_343 (O_343,N_8418,N_9579);
nand UO_344 (O_344,N_8982,N_9349);
and UO_345 (O_345,N_8839,N_9566);
or UO_346 (O_346,N_9353,N_8184);
and UO_347 (O_347,N_8262,N_8694);
xnor UO_348 (O_348,N_9119,N_8390);
nor UO_349 (O_349,N_9655,N_8657);
nand UO_350 (O_350,N_8917,N_8274);
nand UO_351 (O_351,N_9966,N_9880);
or UO_352 (O_352,N_8645,N_8408);
and UO_353 (O_353,N_8815,N_8547);
nand UO_354 (O_354,N_9560,N_8236);
or UO_355 (O_355,N_9972,N_8383);
nand UO_356 (O_356,N_9758,N_8440);
or UO_357 (O_357,N_8639,N_8688);
nand UO_358 (O_358,N_9633,N_8754);
nand UO_359 (O_359,N_9480,N_8105);
nand UO_360 (O_360,N_8511,N_9574);
or UO_361 (O_361,N_9677,N_9802);
or UO_362 (O_362,N_8575,N_9237);
nor UO_363 (O_363,N_9045,N_8561);
nor UO_364 (O_364,N_9826,N_8176);
nor UO_365 (O_365,N_8691,N_8425);
and UO_366 (O_366,N_9791,N_9833);
nor UO_367 (O_367,N_9139,N_9306);
xnor UO_368 (O_368,N_8122,N_9398);
and UO_369 (O_369,N_9692,N_8872);
nor UO_370 (O_370,N_8700,N_9639);
nand UO_371 (O_371,N_9986,N_8275);
nand UO_372 (O_372,N_8264,N_8392);
nand UO_373 (O_373,N_9325,N_8115);
nand UO_374 (O_374,N_8177,N_9063);
nor UO_375 (O_375,N_8263,N_9982);
and UO_376 (O_376,N_9032,N_9935);
nand UO_377 (O_377,N_9400,N_9921);
nand UO_378 (O_378,N_9117,N_8326);
and UO_379 (O_379,N_8929,N_8968);
or UO_380 (O_380,N_9951,N_8005);
nor UO_381 (O_381,N_8996,N_8009);
nand UO_382 (O_382,N_8535,N_8071);
nor UO_383 (O_383,N_9994,N_9652);
nand UO_384 (O_384,N_8805,N_9662);
nor UO_385 (O_385,N_9494,N_8988);
or UO_386 (O_386,N_8209,N_9454);
and UO_387 (O_387,N_8601,N_8877);
nand UO_388 (O_388,N_8767,N_8387);
nand UO_389 (O_389,N_8407,N_8557);
nand UO_390 (O_390,N_9351,N_9737);
or UO_391 (O_391,N_9332,N_9159);
xor UO_392 (O_392,N_8780,N_8642);
nand UO_393 (O_393,N_9295,N_8166);
or UO_394 (O_394,N_9165,N_8404);
nor UO_395 (O_395,N_9673,N_8141);
and UO_396 (O_396,N_9698,N_9254);
and UO_397 (O_397,N_9160,N_9300);
nor UO_398 (O_398,N_9277,N_9581);
nand UO_399 (O_399,N_9600,N_8159);
nand UO_400 (O_400,N_8993,N_9653);
or UO_401 (O_401,N_8659,N_9613);
nor UO_402 (O_402,N_9620,N_9930);
nand UO_403 (O_403,N_8438,N_9172);
nand UO_404 (O_404,N_8285,N_8293);
nand UO_405 (O_405,N_9514,N_9386);
nor UO_406 (O_406,N_9790,N_8077);
nor UO_407 (O_407,N_9634,N_8164);
nand UO_408 (O_408,N_8609,N_8693);
nand UO_409 (O_409,N_9250,N_8314);
nand UO_410 (O_410,N_9469,N_9946);
or UO_411 (O_411,N_8602,N_9161);
nor UO_412 (O_412,N_9654,N_9216);
nor UO_413 (O_413,N_9331,N_9979);
nand UO_414 (O_414,N_8206,N_9251);
nor UO_415 (O_415,N_8193,N_8646);
nor UO_416 (O_416,N_8103,N_9757);
nand UO_417 (O_417,N_8038,N_8519);
and UO_418 (O_418,N_9290,N_8905);
and UO_419 (O_419,N_9520,N_9023);
nand UO_420 (O_420,N_9382,N_9375);
nor UO_421 (O_421,N_9493,N_8043);
nand UO_422 (O_422,N_8154,N_8019);
or UO_423 (O_423,N_9126,N_8952);
or UO_424 (O_424,N_9082,N_8316);
and UO_425 (O_425,N_9430,N_9125);
and UO_426 (O_426,N_8673,N_8797);
or UO_427 (O_427,N_8052,N_8959);
nor UO_428 (O_428,N_8507,N_9735);
nand UO_429 (O_429,N_9171,N_8039);
or UO_430 (O_430,N_8303,N_8738);
nor UO_431 (O_431,N_9039,N_8465);
or UO_432 (O_432,N_9068,N_9812);
nor UO_433 (O_433,N_9578,N_8806);
and UO_434 (O_434,N_9849,N_9206);
and UO_435 (O_435,N_9287,N_9310);
nor UO_436 (O_436,N_9363,N_8722);
and UO_437 (O_437,N_9535,N_8658);
nor UO_438 (O_438,N_9866,N_9543);
or UO_439 (O_439,N_8887,N_9015);
or UO_440 (O_440,N_8354,N_8750);
nor UO_441 (O_441,N_8242,N_8428);
nand UO_442 (O_442,N_8406,N_8647);
and UO_443 (O_443,N_9729,N_9627);
and UO_444 (O_444,N_8775,N_9105);
nand UO_445 (O_445,N_8899,N_9995);
nor UO_446 (O_446,N_8910,N_8030);
or UO_447 (O_447,N_9805,N_9767);
nand UO_448 (O_448,N_9931,N_8069);
or UO_449 (O_449,N_9544,N_9151);
nor UO_450 (O_450,N_8423,N_9078);
and UO_451 (O_451,N_9718,N_8652);
and UO_452 (O_452,N_9809,N_9421);
and UO_453 (O_453,N_9313,N_8817);
nor UO_454 (O_454,N_8567,N_8424);
nand UO_455 (O_455,N_8070,N_9548);
nand UO_456 (O_456,N_8004,N_8104);
or UO_457 (O_457,N_9002,N_9106);
and UO_458 (O_458,N_9649,N_8235);
or UO_459 (O_459,N_9518,N_9091);
nand UO_460 (O_460,N_8464,N_8761);
nand UO_461 (O_461,N_8279,N_8163);
nand UO_462 (O_462,N_9034,N_9992);
or UO_463 (O_463,N_8332,N_9949);
nand UO_464 (O_464,N_8568,N_8220);
nand UO_465 (O_465,N_8621,N_9594);
nor UO_466 (O_466,N_9433,N_9577);
nor UO_467 (O_467,N_8677,N_8467);
or UO_468 (O_468,N_9359,N_8992);
nor UO_469 (O_469,N_8416,N_8847);
nand UO_470 (O_470,N_8560,N_8348);
and UO_471 (O_471,N_8928,N_8083);
nor UO_472 (O_472,N_8173,N_9768);
nand UO_473 (O_473,N_9134,N_8531);
nor UO_474 (O_474,N_8499,N_8315);
nor UO_475 (O_475,N_9985,N_9432);
nor UO_476 (O_476,N_9526,N_8618);
or UO_477 (O_477,N_9319,N_9751);
nand UO_478 (O_478,N_9615,N_9646);
and UO_479 (O_479,N_9676,N_8223);
or UO_480 (O_480,N_9754,N_9455);
nor UO_481 (O_481,N_9088,N_9478);
or UO_482 (O_482,N_9648,N_9318);
nor UO_483 (O_483,N_9396,N_8614);
or UO_484 (O_484,N_8414,N_9707);
nand UO_485 (O_485,N_9173,N_8812);
or UO_486 (O_486,N_9822,N_8433);
nor UO_487 (O_487,N_9604,N_9955);
and UO_488 (O_488,N_9806,N_8110);
nor UO_489 (O_489,N_8085,N_9521);
nand UO_490 (O_490,N_8948,N_9506);
nand UO_491 (O_491,N_8496,N_9529);
or UO_492 (O_492,N_8474,N_8295);
nand UO_493 (O_493,N_8358,N_9426);
and UO_494 (O_494,N_8377,N_8401);
and UO_495 (O_495,N_9716,N_8051);
and UO_496 (O_496,N_9341,N_8632);
nor UO_497 (O_497,N_9038,N_9477);
and UO_498 (O_498,N_8975,N_9731);
nand UO_499 (O_499,N_9390,N_8384);
or UO_500 (O_500,N_8810,N_8880);
nor UO_501 (O_501,N_8243,N_8298);
nor UO_502 (O_502,N_9440,N_9031);
or UO_503 (O_503,N_9590,N_8441);
nor UO_504 (O_504,N_9270,N_9962);
nand UO_505 (O_505,N_9547,N_9713);
nor UO_506 (O_506,N_9787,N_9340);
nand UO_507 (O_507,N_9003,N_8415);
and UO_508 (O_508,N_8769,N_8081);
nand UO_509 (O_509,N_9570,N_8814);
nand UO_510 (O_510,N_8611,N_8786);
or UO_511 (O_511,N_9564,N_9686);
or UO_512 (O_512,N_9451,N_9411);
nand UO_513 (O_513,N_9154,N_9987);
and UO_514 (O_514,N_8807,N_9784);
and UO_515 (O_515,N_9485,N_9912);
nor UO_516 (O_516,N_9077,N_9192);
nor UO_517 (O_517,N_9075,N_9235);
or UO_518 (O_518,N_9201,N_8047);
nand UO_519 (O_519,N_8859,N_8183);
nor UO_520 (O_520,N_8915,N_9980);
nor UO_521 (O_521,N_8597,N_9717);
or UO_522 (O_522,N_8896,N_8829);
and UO_523 (O_523,N_8995,N_8660);
or UO_524 (O_524,N_8257,N_8540);
nor UO_525 (O_525,N_9828,N_9595);
nor UO_526 (O_526,N_8737,N_8307);
nor UO_527 (O_527,N_8587,N_8926);
nor UO_528 (O_528,N_9364,N_8918);
and UO_529 (O_529,N_9439,N_9498);
nand UO_530 (O_530,N_9324,N_8426);
nor UO_531 (O_531,N_8483,N_8082);
and UO_532 (O_532,N_9147,N_8294);
or UO_533 (O_533,N_8516,N_8594);
or UO_534 (O_534,N_8665,N_8456);
or UO_535 (O_535,N_8955,N_9582);
or UO_536 (O_536,N_8219,N_8162);
nor UO_537 (O_537,N_9123,N_8018);
nand UO_538 (O_538,N_9667,N_8411);
and UO_539 (O_539,N_8381,N_8489);
or UO_540 (O_540,N_8720,N_9262);
and UO_541 (O_541,N_9470,N_8089);
nor UO_542 (O_542,N_8748,N_8889);
or UO_543 (O_543,N_9510,N_8095);
nand UO_544 (O_544,N_9568,N_9144);
and UO_545 (O_545,N_8864,N_9573);
and UO_546 (O_546,N_9872,N_8161);
and UO_547 (O_547,N_9090,N_9524);
nand UO_548 (O_548,N_9497,N_9072);
or UO_549 (O_549,N_9700,N_9370);
or UO_550 (O_550,N_9191,N_8706);
nand UO_551 (O_551,N_9638,N_9089);
nor UO_552 (O_552,N_8080,N_9001);
nand UO_553 (O_553,N_9778,N_9048);
or UO_554 (O_554,N_9084,N_8032);
nor UO_555 (O_555,N_9997,N_8773);
and UO_556 (O_556,N_8842,N_8389);
nor UO_557 (O_557,N_9000,N_8027);
nor UO_558 (O_558,N_8841,N_9228);
nand UO_559 (O_559,N_9519,N_9112);
and UO_560 (O_560,N_9505,N_8252);
or UO_561 (O_561,N_8228,N_8914);
or UO_562 (O_562,N_8937,N_9682);
or UO_563 (O_563,N_9495,N_9666);
nor UO_564 (O_564,N_9769,N_9651);
nand UO_565 (O_565,N_8977,N_9356);
nand UO_566 (O_566,N_8764,N_9321);
xor UO_567 (O_567,N_8599,N_9965);
or UO_568 (O_568,N_9489,N_9059);
or UO_569 (O_569,N_9083,N_9968);
nand UO_570 (O_570,N_8550,N_9456);
xnor UO_571 (O_571,N_8604,N_9232);
or UO_572 (O_572,N_8885,N_8686);
nor UO_573 (O_573,N_9214,N_8711);
and UO_574 (O_574,N_9724,N_8339);
nor UO_575 (O_575,N_9131,N_9954);
or UO_576 (O_576,N_8997,N_9138);
nor UO_577 (O_577,N_9471,N_8719);
or UO_578 (O_578,N_8593,N_9509);
nand UO_579 (O_579,N_9459,N_9720);
nor UO_580 (O_580,N_8925,N_9556);
nand UO_581 (O_581,N_8631,N_8752);
or UO_582 (O_582,N_8259,N_8517);
or UO_583 (O_583,N_9766,N_8459);
and UO_584 (O_584,N_8524,N_8136);
or UO_585 (O_585,N_9629,N_8976);
and UO_586 (O_586,N_8165,N_8869);
and UO_587 (O_587,N_9419,N_8286);
nand UO_588 (O_588,N_8435,N_8470);
nand UO_589 (O_589,N_8462,N_9847);
and UO_590 (O_590,N_8768,N_9501);
nand UO_591 (O_591,N_8084,N_8834);
nand UO_592 (O_592,N_8846,N_9399);
or UO_593 (O_593,N_9346,N_9021);
nand UO_594 (O_594,N_9352,N_9580);
or UO_595 (O_595,N_9863,N_8851);
or UO_596 (O_596,N_9221,N_8361);
and UO_597 (O_597,N_8500,N_9779);
nand UO_598 (O_598,N_9924,N_9593);
or UO_599 (O_599,N_8204,N_8374);
nor UO_600 (O_600,N_9484,N_8875);
nor UO_601 (O_601,N_9777,N_8553);
or UO_602 (O_602,N_8121,N_8190);
nor UO_603 (O_603,N_9504,N_9846);
or UO_604 (O_604,N_9752,N_9047);
nand UO_605 (O_605,N_8651,N_8922);
nand UO_606 (O_606,N_9189,N_9706);
nor UO_607 (O_607,N_9909,N_8484);
nor UO_608 (O_608,N_9663,N_8215);
nor UO_609 (O_609,N_8386,N_9168);
nor UO_610 (O_610,N_9761,N_8367);
or UO_611 (O_611,N_9689,N_9550);
or UO_612 (O_612,N_8351,N_8911);
nand UO_613 (O_613,N_8096,N_9339);
nor UO_614 (O_614,N_8227,N_8357);
or UO_615 (O_615,N_9760,N_8283);
nand UO_616 (O_616,N_9182,N_8762);
or UO_617 (O_617,N_9304,N_8571);
and UO_618 (O_618,N_8449,N_8763);
or UO_619 (O_619,N_9525,N_9865);
or UO_620 (O_620,N_8776,N_9366);
or UO_621 (O_621,N_8824,N_9797);
xor UO_622 (O_622,N_8853,N_9071);
nand UO_623 (O_623,N_8169,N_8826);
and UO_624 (O_624,N_9169,N_8261);
nand UO_625 (O_625,N_8746,N_8025);
or UO_626 (O_626,N_9608,N_9490);
and UO_627 (O_627,N_8726,N_9879);
nand UO_628 (O_628,N_8777,N_9691);
nand UO_629 (O_629,N_8313,N_9508);
and UO_630 (O_630,N_8927,N_9914);
nand UO_631 (O_631,N_9883,N_9753);
and UO_632 (O_632,N_9143,N_9726);
and UO_633 (O_633,N_9808,N_9841);
nand UO_634 (O_634,N_8244,N_8701);
nor UO_635 (O_635,N_9801,N_9033);
nor UO_636 (O_636,N_9205,N_8063);
and UO_637 (O_637,N_8378,N_8791);
and UO_638 (O_638,N_8538,N_8200);
or UO_639 (O_639,N_8240,N_8229);
nor UO_640 (O_640,N_9402,N_8522);
and UO_641 (O_641,N_8296,N_8510);
nor UO_642 (O_642,N_8731,N_9415);
or UO_643 (O_643,N_8437,N_8453);
and UO_644 (O_644,N_8861,N_8454);
nand UO_645 (O_645,N_8492,N_9005);
nand UO_646 (O_646,N_9927,N_8908);
and UO_647 (O_647,N_8191,N_8936);
nor UO_648 (O_648,N_9983,N_8478);
nand UO_649 (O_649,N_8087,N_9612);
nand UO_650 (O_650,N_8152,N_9465);
nand UO_651 (O_651,N_9016,N_8674);
and UO_652 (O_652,N_9474,N_9668);
nor UO_653 (O_653,N_8795,N_9274);
nand UO_654 (O_654,N_8233,N_9559);
nand UO_655 (O_655,N_9690,N_9040);
or UO_656 (O_656,N_9624,N_9970);
nand UO_657 (O_657,N_9466,N_8305);
and UO_658 (O_658,N_8399,N_8324);
nand UO_659 (O_659,N_9950,N_8582);
nor UO_660 (O_660,N_8276,N_8458);
nand UO_661 (O_661,N_9479,N_8109);
and UO_662 (O_662,N_9785,N_9486);
nand UO_663 (O_663,N_9445,N_9619);
nor UO_664 (O_664,N_9365,N_8210);
nand UO_665 (O_665,N_9928,N_8172);
nand UO_666 (O_666,N_9483,N_8717);
and UO_667 (O_667,N_8802,N_8779);
and UO_668 (O_668,N_8984,N_8011);
nand UO_669 (O_669,N_9307,N_9591);
xor UO_670 (O_670,N_8669,N_9625);
or UO_671 (O_671,N_9628,N_8608);
and UO_672 (O_672,N_9971,N_9643);
or UO_673 (O_673,N_9111,N_9733);
and UO_674 (O_674,N_9424,N_9977);
nand UO_675 (O_675,N_9257,N_9097);
nand UO_676 (O_676,N_9135,N_9942);
or UO_677 (O_677,N_9661,N_9181);
or UO_678 (O_678,N_8634,N_8124);
or UO_679 (O_679,N_8551,N_9603);
or UO_680 (O_680,N_9940,N_9115);
and UO_681 (O_681,N_8564,N_9209);
or UO_682 (O_682,N_8207,N_9756);
nand UO_683 (O_683,N_8636,N_9601);
or UO_684 (O_684,N_8330,N_8759);
or UO_685 (O_685,N_9414,N_9552);
nor UO_686 (O_686,N_9721,N_9457);
or UO_687 (O_687,N_9699,N_8735);
nor UO_688 (O_688,N_8135,N_8321);
nand UO_689 (O_689,N_9079,N_8526);
and UO_690 (O_690,N_8931,N_9299);
nand UO_691 (O_691,N_8751,N_9792);
nand UO_692 (O_692,N_8592,N_9118);
nand UO_693 (O_693,N_9780,N_9773);
nor UO_694 (O_694,N_9443,N_9710);
and UO_695 (O_695,N_9369,N_8655);
or UO_696 (O_696,N_8106,N_8186);
and UO_697 (O_697,N_9249,N_8644);
nor UO_698 (O_698,N_8447,N_9253);
nand UO_699 (O_699,N_9204,N_9020);
or UO_700 (O_700,N_8320,N_9799);
nor UO_701 (O_701,N_8893,N_8058);
nor UO_702 (O_702,N_9923,N_8417);
nand UO_703 (O_703,N_9969,N_9195);
nand UO_704 (O_704,N_9347,N_8410);
nor UO_705 (O_705,N_8098,N_8793);
nand UO_706 (O_706,N_8156,N_8059);
or UO_707 (O_707,N_8932,N_8656);
and UO_708 (O_708,N_9642,N_8515);
and UO_709 (O_709,N_8427,N_8372);
nor UO_710 (O_710,N_8370,N_8217);
nand UO_711 (O_711,N_9896,N_8873);
and UO_712 (O_712,N_8251,N_8863);
nand UO_713 (O_713,N_9406,N_9830);
and UO_714 (O_714,N_9637,N_8461);
nand UO_715 (O_715,N_8583,N_9389);
or UO_716 (O_716,N_8267,N_9107);
or UO_717 (O_717,N_8649,N_8188);
and UO_718 (O_718,N_9170,N_8224);
nor UO_719 (O_719,N_8318,N_8566);
nor UO_720 (O_720,N_9409,N_9738);
and UO_721 (O_721,N_9425,N_8684);
and UO_722 (O_722,N_8529,N_8380);
or UO_723 (O_723,N_9320,N_8563);
or UO_724 (O_724,N_8527,N_8616);
and UO_725 (O_725,N_8402,N_9621);
nor UO_726 (O_726,N_9734,N_9322);
nor UO_727 (O_727,N_9297,N_8698);
nand UO_728 (O_728,N_8343,N_9536);
and UO_729 (O_729,N_9264,N_9679);
and UO_730 (O_730,N_9607,N_8965);
or UO_731 (O_731,N_8913,N_8245);
nand UO_732 (O_732,N_9687,N_9933);
nand UO_733 (O_733,N_8153,N_9867);
nor UO_734 (O_734,N_9328,N_8157);
or UO_735 (O_735,N_8625,N_8643);
and UO_736 (O_736,N_8505,N_9660);
and UO_737 (O_737,N_8023,N_8741);
and UO_738 (O_738,N_9551,N_9669);
and UO_739 (O_739,N_8297,N_8137);
and UO_740 (O_740,N_8626,N_9611);
or UO_741 (O_741,N_9736,N_9428);
and UO_742 (O_742,N_9395,N_9804);
or UO_743 (O_743,N_9137,N_9271);
nor UO_744 (O_744,N_8637,N_8697);
nand UO_745 (O_745,N_9429,N_8743);
or UO_746 (O_746,N_8055,N_9127);
and UO_747 (O_747,N_8144,N_9701);
nor UO_748 (O_748,N_8502,N_8546);
and UO_749 (O_749,N_9408,N_8730);
and UO_750 (O_750,N_8382,N_8225);
nor UO_751 (O_751,N_9153,N_9848);
nand UO_752 (O_752,N_9420,N_9085);
or UO_753 (O_753,N_9882,N_9820);
nor UO_754 (O_754,N_8342,N_8633);
nor UO_755 (O_755,N_8486,N_9599);
nand UO_756 (O_756,N_9967,N_8683);
and UO_757 (O_757,N_9771,N_9435);
nand UO_758 (O_758,N_8353,N_9936);
nand UO_759 (O_759,N_8874,N_8439);
or UO_760 (O_760,N_9110,N_8053);
nand UO_761 (O_761,N_9286,N_9291);
and UO_762 (O_762,N_9354,N_9945);
nor UO_763 (O_763,N_8375,N_8198);
or UO_764 (O_764,N_9832,N_8400);
or UO_765 (O_765,N_9727,N_9586);
and UO_766 (O_766,N_9092,N_9528);
nand UO_767 (O_767,N_9442,N_9549);
and UO_768 (O_768,N_9302,N_8412);
and UO_769 (O_769,N_8040,N_8270);
or UO_770 (O_770,N_9697,N_8947);
nand UO_771 (O_771,N_9631,N_9665);
and UO_772 (O_772,N_9605,N_9412);
nand UO_773 (O_773,N_8472,N_9337);
and UO_774 (O_774,N_8664,N_9064);
nor UO_775 (O_775,N_8680,N_9114);
nor UO_776 (O_776,N_9917,N_8049);
nor UO_777 (O_777,N_8212,N_9413);
nor UO_778 (O_778,N_8629,N_9823);
nand UO_779 (O_779,N_8554,N_8213);
or UO_780 (O_780,N_9870,N_9446);
nor UO_781 (O_781,N_8707,N_9383);
xor UO_782 (O_782,N_8892,N_9958);
nand UO_783 (O_783,N_8617,N_8981);
nor UO_784 (O_784,N_9142,N_8013);
nor UO_785 (O_785,N_8986,N_9472);
and UO_786 (O_786,N_9449,N_9796);
or UO_787 (O_787,N_8600,N_9261);
or UO_788 (O_788,N_8774,N_8838);
or UO_789 (O_789,N_8506,N_8855);
nor UO_790 (O_790,N_8497,N_9584);
nand UO_791 (O_791,N_8787,N_9202);
or UO_792 (O_792,N_9252,N_9728);
nand UO_793 (O_793,N_8574,N_8883);
and UO_794 (O_794,N_9121,N_9889);
nor UO_795 (O_795,N_9024,N_8066);
nand UO_796 (O_796,N_9158,N_8867);
nor UO_797 (O_797,N_8771,N_9893);
or UO_798 (O_798,N_8513,N_8291);
and UO_799 (O_799,N_9630,N_9683);
and UO_800 (O_800,N_9305,N_9461);
or UO_801 (O_801,N_9109,N_8265);
nand UO_802 (O_802,N_9057,N_9329);
or UO_803 (O_803,N_8419,N_8473);
nor UO_804 (O_804,N_8422,N_8778);
or UO_805 (O_805,N_8714,N_9239);
or UO_806 (O_806,N_8534,N_9348);
nand UO_807 (O_807,N_9333,N_8477);
or UO_808 (O_808,N_9416,N_8819);
and UO_809 (O_809,N_9800,N_8909);
and UO_810 (O_810,N_8182,N_8138);
nor UO_811 (O_811,N_9226,N_9705);
and UO_812 (O_812,N_8341,N_9014);
and UO_813 (O_813,N_8189,N_8056);
and UO_814 (O_814,N_9452,N_9293);
or UO_815 (O_815,N_8537,N_8641);
or UO_816 (O_816,N_9061,N_8951);
and UO_817 (O_817,N_9330,N_8112);
or UO_818 (O_818,N_9911,N_9708);
or UO_819 (O_819,N_9438,N_8809);
nor UO_820 (O_820,N_9183,N_9086);
nor UO_821 (O_821,N_9565,N_8450);
and UO_822 (O_822,N_8921,N_8232);
nand UO_823 (O_823,N_9238,N_9401);
or UO_824 (O_824,N_8715,N_8234);
nand UO_825 (O_825,N_8907,N_9884);
or UO_826 (O_826,N_9065,N_9087);
or UO_827 (O_827,N_9770,N_9374);
nand UO_828 (O_828,N_9984,N_8312);
and UO_829 (O_829,N_9377,N_9597);
or UO_830 (O_830,N_9555,N_9881);
nor UO_831 (O_831,N_8491,N_8306);
or UO_832 (O_832,N_9745,N_9265);
nor UO_833 (O_833,N_8744,N_8852);
and UO_834 (O_834,N_9179,N_8830);
and UO_835 (O_835,N_8146,N_9894);
and UO_836 (O_836,N_8086,N_9938);
nor UO_837 (O_837,N_8100,N_9387);
nand UO_838 (O_838,N_9378,N_8272);
and UO_839 (O_839,N_9695,N_9916);
and UO_840 (O_840,N_8031,N_9857);
nand UO_841 (O_841,N_8238,N_8421);
nand UO_842 (O_842,N_8091,N_9222);
nor UO_843 (O_843,N_9224,N_8119);
nand UO_844 (O_844,N_9338,N_8942);
or UO_845 (O_845,N_9592,N_8476);
and UO_846 (O_846,N_8963,N_9027);
nand UO_847 (O_847,N_8901,N_8366);
nor UO_848 (O_848,N_8695,N_9636);
or UO_849 (O_849,N_9755,N_8990);
or UO_850 (O_850,N_8723,N_9963);
nor UO_851 (O_851,N_9334,N_9918);
nand UO_852 (O_852,N_9197,N_8271);
or UO_853 (O_853,N_8525,N_8338);
and UO_854 (O_854,N_8409,N_9384);
or UO_855 (O_855,N_9859,N_9854);
and UO_856 (O_856,N_9104,N_8434);
and UO_857 (O_857,N_9042,N_8349);
or UO_858 (O_858,N_8336,N_9460);
nand UO_859 (O_859,N_8924,N_9423);
nor UO_860 (O_860,N_9152,N_9877);
or UO_861 (O_861,N_8035,N_9094);
and UO_862 (O_862,N_9492,N_8277);
nor UO_863 (O_863,N_9537,N_9772);
nor UO_864 (O_864,N_9108,N_8845);
nor UO_865 (O_865,N_9892,N_9335);
nand UO_866 (O_866,N_8724,N_8006);
nor UO_867 (O_867,N_9367,N_8760);
or UO_868 (O_868,N_8201,N_8062);
nand UO_869 (O_869,N_8650,N_9913);
nand UO_870 (O_870,N_9468,N_8037);
and UO_871 (O_871,N_8742,N_8151);
nand UO_872 (O_872,N_9959,N_8133);
nand UO_873 (O_873,N_8713,N_9694);
nor UO_874 (O_874,N_8520,N_8605);
and UO_875 (O_875,N_8503,N_9583);
nor UO_876 (O_876,N_9280,N_8388);
nand UO_877 (O_877,N_8702,N_9730);
or UO_878 (O_878,N_9096,N_9672);
nor UO_879 (O_879,N_9837,N_8249);
nand UO_880 (O_880,N_9656,N_8068);
nor UO_881 (O_881,N_8933,N_8185);
or UO_882 (O_882,N_9055,N_8854);
nor UO_883 (O_883,N_9856,N_9458);
or UO_884 (O_884,N_8117,N_8194);
and UO_885 (O_885,N_9803,N_9952);
or UO_886 (O_886,N_8712,N_8991);
or UO_887 (O_887,N_9004,N_8891);
nand UO_888 (O_888,N_9901,N_9437);
nand UO_889 (O_889,N_9618,N_8094);
and UO_890 (O_890,N_9900,N_8543);
or UO_891 (O_891,N_8111,N_9101);
nor UO_892 (O_892,N_8820,N_9229);
nand UO_893 (O_893,N_9392,N_8578);
and UO_894 (O_894,N_9219,N_9053);
and UO_895 (O_895,N_9939,N_8862);
nor UO_896 (O_896,N_8528,N_8579);
xnor UO_897 (O_897,N_9915,N_9067);
or UO_898 (O_898,N_8088,N_9281);
nand UO_899 (O_899,N_9376,N_9765);
nand UO_900 (O_900,N_9744,N_8740);
nor UO_901 (O_901,N_9878,N_9722);
nor UO_902 (O_902,N_9200,N_9243);
nand UO_903 (O_903,N_9991,N_8912);
nor UO_904 (O_904,N_8345,N_8344);
nand UO_905 (O_905,N_8835,N_8699);
or UO_906 (O_906,N_9103,N_8985);
or UO_907 (O_907,N_9534,N_8653);
and UO_908 (O_908,N_9275,N_8463);
nor UO_909 (O_909,N_8175,N_9746);
nand UO_910 (O_910,N_9268,N_9531);
or UO_911 (O_911,N_8466,N_8329);
or UO_912 (O_912,N_8322,N_8589);
nand UO_913 (O_913,N_9569,N_8118);
nand UO_914 (O_914,N_9336,N_9225);
nor UO_915 (O_915,N_9167,N_8542);
or UO_916 (O_916,N_9696,N_9207);
and UO_917 (O_917,N_8355,N_8607);
nor UO_918 (O_918,N_8999,N_9622);
and UO_919 (O_919,N_8142,N_8268);
nand UO_920 (O_920,N_8591,N_8139);
nand UO_921 (O_921,N_8026,N_8944);
nand UO_922 (O_922,N_8530,N_9831);
and UO_923 (O_923,N_8282,N_8034);
nor UO_924 (O_924,N_9575,N_9259);
and UO_925 (O_925,N_8362,N_8073);
nand UO_926 (O_926,N_9709,N_9373);
or UO_927 (O_927,N_9010,N_8020);
or UO_928 (O_928,N_8211,N_8260);
nor UO_929 (O_929,N_8126,N_8630);
nor UO_930 (O_930,N_9394,N_8079);
and UO_931 (O_931,N_8967,N_8222);
nand UO_932 (O_932,N_9840,N_9973);
nor UO_933 (O_933,N_8533,N_9019);
or UO_934 (O_934,N_8836,N_8487);
nand UO_935 (O_935,N_9908,N_8001);
nor UO_936 (O_936,N_9198,N_9723);
nor UO_937 (O_937,N_9748,N_8364);
xnor UO_938 (O_938,N_8468,N_8120);
and UO_939 (O_939,N_9393,N_8258);
nor UO_940 (O_940,N_8352,N_9996);
nand UO_941 (O_941,N_8577,N_8555);
nor UO_942 (O_942,N_9864,N_9188);
nor UO_943 (O_943,N_9567,N_8036);
nand UO_944 (O_944,N_8208,N_8958);
or UO_945 (O_945,N_8078,N_9011);
nor UO_946 (O_946,N_8231,N_8696);
and UO_947 (O_947,N_9685,N_8623);
or UO_948 (O_948,N_8943,N_9522);
nand UO_949 (O_949,N_8192,N_8930);
or UO_950 (O_950,N_8770,N_8687);
nor UO_951 (O_951,N_9344,N_8017);
nand UO_952 (O_952,N_9241,N_9203);
nor UO_953 (O_953,N_9136,N_9185);
or UO_954 (O_954,N_9644,N_9989);
and UO_955 (O_955,N_9684,N_8703);
nand UO_956 (O_956,N_9130,N_9910);
and UO_957 (O_957,N_9240,N_8432);
and UO_958 (O_958,N_8685,N_9961);
and UO_959 (O_959,N_8325,N_8284);
nor UO_960 (O_960,N_9874,N_8640);
and UO_961 (O_961,N_8570,N_8690);
nor UO_962 (O_962,N_9177,N_9327);
nand UO_963 (O_963,N_8559,N_9839);
nor UO_964 (O_964,N_9576,N_9838);
nand UO_965 (O_965,N_9670,N_9816);
and UO_966 (O_966,N_9076,N_9417);
and UO_967 (O_967,N_9811,N_9488);
nor UO_968 (O_968,N_9523,N_9671);
or UO_969 (O_969,N_9890,N_8150);
nor UO_970 (O_970,N_9500,N_9124);
nor UO_971 (O_971,N_9317,N_8369);
or UO_972 (O_972,N_9635,N_8635);
and UO_973 (O_973,N_9282,N_9589);
and UO_974 (O_974,N_9272,N_8429);
or UO_975 (O_975,N_9922,N_8800);
nor UO_976 (O_976,N_9095,N_9776);
nor UO_977 (O_977,N_9361,N_9149);
xor UO_978 (O_978,N_9215,N_8989);
nand UO_979 (O_979,N_8966,N_9943);
or UO_980 (O_980,N_9447,N_8300);
and UO_981 (O_981,N_8290,N_9308);
nor UO_982 (O_982,N_8360,N_8692);
nor UO_983 (O_983,N_9614,N_9046);
and UO_984 (O_984,N_9481,N_8008);
nand UO_985 (O_985,N_9907,N_9503);
and UO_986 (O_986,N_9120,N_9681);
nor UO_987 (O_987,N_9704,N_9009);
or UO_988 (O_988,N_8586,N_9988);
or UO_989 (O_989,N_8132,N_9140);
nor UO_990 (O_990,N_8308,N_9853);
and UO_991 (O_991,N_9664,N_8598);
and UO_992 (O_992,N_9178,N_9542);
and UO_993 (O_993,N_9516,N_9368);
or UO_994 (O_994,N_8961,N_9122);
and UO_995 (O_995,N_8287,N_9233);
or UO_996 (O_996,N_9674,N_9041);
or UO_997 (O_997,N_8398,N_9588);
nand UO_998 (O_998,N_8904,N_9150);
nor UO_999 (O_999,N_8833,N_8790);
nand UO_1000 (O_1000,N_9681,N_8157);
nor UO_1001 (O_1001,N_9372,N_8493);
nand UO_1002 (O_1002,N_9238,N_9449);
or UO_1003 (O_1003,N_8662,N_8445);
nand UO_1004 (O_1004,N_9271,N_9443);
nor UO_1005 (O_1005,N_8760,N_8694);
or UO_1006 (O_1006,N_9367,N_8586);
nand UO_1007 (O_1007,N_8685,N_8908);
nand UO_1008 (O_1008,N_8505,N_9512);
nand UO_1009 (O_1009,N_9667,N_9477);
and UO_1010 (O_1010,N_9757,N_9738);
or UO_1011 (O_1011,N_9841,N_9787);
nor UO_1012 (O_1012,N_8903,N_9650);
nor UO_1013 (O_1013,N_8240,N_8728);
and UO_1014 (O_1014,N_8459,N_9056);
or UO_1015 (O_1015,N_9973,N_9230);
or UO_1016 (O_1016,N_9840,N_9725);
or UO_1017 (O_1017,N_9080,N_8518);
and UO_1018 (O_1018,N_9524,N_9186);
nand UO_1019 (O_1019,N_9943,N_9998);
nor UO_1020 (O_1020,N_8014,N_9706);
nor UO_1021 (O_1021,N_8495,N_9943);
and UO_1022 (O_1022,N_9205,N_9054);
or UO_1023 (O_1023,N_8076,N_9833);
and UO_1024 (O_1024,N_8171,N_9142);
and UO_1025 (O_1025,N_8247,N_9250);
nor UO_1026 (O_1026,N_8067,N_9349);
nand UO_1027 (O_1027,N_9919,N_9927);
and UO_1028 (O_1028,N_8997,N_8927);
and UO_1029 (O_1029,N_9486,N_9034);
and UO_1030 (O_1030,N_8201,N_9646);
or UO_1031 (O_1031,N_8147,N_8777);
and UO_1032 (O_1032,N_9851,N_8204);
nor UO_1033 (O_1033,N_8884,N_9747);
nor UO_1034 (O_1034,N_8516,N_8670);
or UO_1035 (O_1035,N_8033,N_8294);
or UO_1036 (O_1036,N_8715,N_9037);
nand UO_1037 (O_1037,N_9059,N_9132);
nand UO_1038 (O_1038,N_9685,N_8458);
or UO_1039 (O_1039,N_8229,N_9358);
or UO_1040 (O_1040,N_9981,N_8847);
nand UO_1041 (O_1041,N_8604,N_9804);
and UO_1042 (O_1042,N_8370,N_9603);
and UO_1043 (O_1043,N_9025,N_9669);
nand UO_1044 (O_1044,N_8281,N_8254);
or UO_1045 (O_1045,N_9076,N_8454);
nand UO_1046 (O_1046,N_8086,N_9009);
and UO_1047 (O_1047,N_8547,N_8681);
and UO_1048 (O_1048,N_8164,N_8045);
nand UO_1049 (O_1049,N_8076,N_8181);
nor UO_1050 (O_1050,N_9405,N_9516);
nand UO_1051 (O_1051,N_9128,N_8806);
nor UO_1052 (O_1052,N_9575,N_8574);
nand UO_1053 (O_1053,N_9848,N_8013);
or UO_1054 (O_1054,N_9273,N_8701);
and UO_1055 (O_1055,N_9495,N_9768);
and UO_1056 (O_1056,N_8232,N_9442);
and UO_1057 (O_1057,N_8457,N_9662);
nand UO_1058 (O_1058,N_8396,N_8905);
and UO_1059 (O_1059,N_8545,N_9085);
nor UO_1060 (O_1060,N_8308,N_8054);
nand UO_1061 (O_1061,N_8157,N_9205);
and UO_1062 (O_1062,N_9606,N_8098);
nand UO_1063 (O_1063,N_9994,N_9703);
or UO_1064 (O_1064,N_9689,N_8732);
nand UO_1065 (O_1065,N_8236,N_9314);
or UO_1066 (O_1066,N_8019,N_8650);
nand UO_1067 (O_1067,N_8022,N_8392);
or UO_1068 (O_1068,N_8641,N_9226);
and UO_1069 (O_1069,N_9571,N_8284);
or UO_1070 (O_1070,N_9343,N_9246);
or UO_1071 (O_1071,N_9822,N_8178);
or UO_1072 (O_1072,N_8896,N_9472);
nand UO_1073 (O_1073,N_8534,N_8342);
xor UO_1074 (O_1074,N_8116,N_8298);
nand UO_1075 (O_1075,N_9289,N_9338);
nor UO_1076 (O_1076,N_9279,N_8886);
or UO_1077 (O_1077,N_9607,N_8590);
nand UO_1078 (O_1078,N_8380,N_8634);
and UO_1079 (O_1079,N_9853,N_9422);
nand UO_1080 (O_1080,N_9365,N_9355);
xor UO_1081 (O_1081,N_8907,N_8066);
or UO_1082 (O_1082,N_8991,N_9661);
xnor UO_1083 (O_1083,N_8282,N_8628);
nor UO_1084 (O_1084,N_9050,N_8252);
nand UO_1085 (O_1085,N_9516,N_8485);
and UO_1086 (O_1086,N_9969,N_8337);
nor UO_1087 (O_1087,N_9354,N_9379);
or UO_1088 (O_1088,N_8044,N_9062);
nand UO_1089 (O_1089,N_9694,N_9566);
xnor UO_1090 (O_1090,N_9525,N_9720);
nor UO_1091 (O_1091,N_9719,N_9804);
and UO_1092 (O_1092,N_9011,N_8531);
nor UO_1093 (O_1093,N_9571,N_8335);
nand UO_1094 (O_1094,N_9734,N_9160);
and UO_1095 (O_1095,N_9045,N_9391);
nor UO_1096 (O_1096,N_9610,N_9123);
or UO_1097 (O_1097,N_8152,N_9364);
nor UO_1098 (O_1098,N_9523,N_8351);
or UO_1099 (O_1099,N_8225,N_8376);
and UO_1100 (O_1100,N_8383,N_9821);
nand UO_1101 (O_1101,N_9919,N_8960);
nand UO_1102 (O_1102,N_8779,N_9921);
and UO_1103 (O_1103,N_9716,N_8115);
nand UO_1104 (O_1104,N_9131,N_8289);
nand UO_1105 (O_1105,N_8003,N_8437);
or UO_1106 (O_1106,N_8993,N_9430);
and UO_1107 (O_1107,N_9859,N_9413);
nand UO_1108 (O_1108,N_8610,N_9828);
and UO_1109 (O_1109,N_8079,N_9103);
and UO_1110 (O_1110,N_9289,N_9135);
nor UO_1111 (O_1111,N_9658,N_8842);
and UO_1112 (O_1112,N_8716,N_9224);
or UO_1113 (O_1113,N_8286,N_9749);
nand UO_1114 (O_1114,N_9232,N_9088);
and UO_1115 (O_1115,N_9696,N_8887);
and UO_1116 (O_1116,N_9019,N_9447);
nor UO_1117 (O_1117,N_9725,N_9365);
nand UO_1118 (O_1118,N_9694,N_9005);
or UO_1119 (O_1119,N_9720,N_9864);
or UO_1120 (O_1120,N_8273,N_9839);
or UO_1121 (O_1121,N_8444,N_9531);
nor UO_1122 (O_1122,N_9068,N_8292);
and UO_1123 (O_1123,N_8461,N_8175);
or UO_1124 (O_1124,N_8915,N_8830);
or UO_1125 (O_1125,N_8989,N_8439);
nand UO_1126 (O_1126,N_9067,N_9514);
nor UO_1127 (O_1127,N_8904,N_9205);
or UO_1128 (O_1128,N_8611,N_9477);
and UO_1129 (O_1129,N_8832,N_9726);
nor UO_1130 (O_1130,N_8025,N_9968);
and UO_1131 (O_1131,N_9085,N_8169);
nand UO_1132 (O_1132,N_8981,N_9115);
and UO_1133 (O_1133,N_8176,N_8742);
nand UO_1134 (O_1134,N_8954,N_8888);
nor UO_1135 (O_1135,N_8107,N_8182);
nor UO_1136 (O_1136,N_9878,N_9588);
nand UO_1137 (O_1137,N_9510,N_8892);
and UO_1138 (O_1138,N_8042,N_8945);
and UO_1139 (O_1139,N_9094,N_9079);
nor UO_1140 (O_1140,N_8519,N_9013);
nand UO_1141 (O_1141,N_9909,N_9983);
nor UO_1142 (O_1142,N_9626,N_9394);
and UO_1143 (O_1143,N_9037,N_9756);
nor UO_1144 (O_1144,N_8168,N_9249);
or UO_1145 (O_1145,N_8763,N_8250);
nor UO_1146 (O_1146,N_8882,N_9916);
xor UO_1147 (O_1147,N_8189,N_9548);
nor UO_1148 (O_1148,N_9562,N_8675);
nor UO_1149 (O_1149,N_9265,N_9987);
nor UO_1150 (O_1150,N_9731,N_8034);
or UO_1151 (O_1151,N_9727,N_9736);
nand UO_1152 (O_1152,N_9910,N_9386);
and UO_1153 (O_1153,N_9730,N_8221);
or UO_1154 (O_1154,N_8477,N_8484);
nor UO_1155 (O_1155,N_9198,N_9829);
and UO_1156 (O_1156,N_8179,N_9640);
and UO_1157 (O_1157,N_9482,N_9565);
or UO_1158 (O_1158,N_9732,N_9853);
nor UO_1159 (O_1159,N_9259,N_8225);
and UO_1160 (O_1160,N_9641,N_9749);
nand UO_1161 (O_1161,N_9779,N_9314);
and UO_1162 (O_1162,N_8104,N_8563);
nor UO_1163 (O_1163,N_9874,N_8664);
or UO_1164 (O_1164,N_9378,N_8137);
nand UO_1165 (O_1165,N_9375,N_8082);
and UO_1166 (O_1166,N_9235,N_9677);
nor UO_1167 (O_1167,N_9925,N_9180);
nor UO_1168 (O_1168,N_9551,N_9289);
nand UO_1169 (O_1169,N_8097,N_8734);
nor UO_1170 (O_1170,N_9902,N_9966);
nor UO_1171 (O_1171,N_9534,N_9109);
and UO_1172 (O_1172,N_9373,N_8484);
nand UO_1173 (O_1173,N_8150,N_8657);
and UO_1174 (O_1174,N_8165,N_8661);
nand UO_1175 (O_1175,N_9193,N_9551);
nor UO_1176 (O_1176,N_8396,N_8716);
nand UO_1177 (O_1177,N_8135,N_9486);
and UO_1178 (O_1178,N_8738,N_8055);
nor UO_1179 (O_1179,N_8339,N_8802);
nor UO_1180 (O_1180,N_9299,N_9750);
or UO_1181 (O_1181,N_9865,N_9912);
nand UO_1182 (O_1182,N_8625,N_9571);
nor UO_1183 (O_1183,N_9383,N_9411);
nor UO_1184 (O_1184,N_8144,N_9997);
nand UO_1185 (O_1185,N_9047,N_8530);
nand UO_1186 (O_1186,N_9384,N_8991);
or UO_1187 (O_1187,N_8314,N_9007);
nor UO_1188 (O_1188,N_9052,N_9708);
nand UO_1189 (O_1189,N_9052,N_8583);
or UO_1190 (O_1190,N_8320,N_9749);
nand UO_1191 (O_1191,N_9005,N_8923);
nand UO_1192 (O_1192,N_9699,N_8681);
and UO_1193 (O_1193,N_8962,N_8548);
or UO_1194 (O_1194,N_8100,N_9155);
nand UO_1195 (O_1195,N_8819,N_9007);
nor UO_1196 (O_1196,N_8768,N_9900);
nor UO_1197 (O_1197,N_9469,N_9786);
or UO_1198 (O_1198,N_9607,N_9923);
and UO_1199 (O_1199,N_9513,N_8375);
nor UO_1200 (O_1200,N_8392,N_8386);
or UO_1201 (O_1201,N_9118,N_9971);
nor UO_1202 (O_1202,N_9543,N_8056);
or UO_1203 (O_1203,N_9837,N_9888);
nand UO_1204 (O_1204,N_9729,N_9953);
and UO_1205 (O_1205,N_8353,N_8863);
or UO_1206 (O_1206,N_9910,N_9847);
or UO_1207 (O_1207,N_9199,N_8859);
nor UO_1208 (O_1208,N_9394,N_8956);
nor UO_1209 (O_1209,N_8389,N_9010);
nor UO_1210 (O_1210,N_9302,N_8429);
and UO_1211 (O_1211,N_9181,N_9628);
and UO_1212 (O_1212,N_8036,N_8587);
or UO_1213 (O_1213,N_9756,N_9135);
nand UO_1214 (O_1214,N_8705,N_8080);
nor UO_1215 (O_1215,N_9347,N_8478);
and UO_1216 (O_1216,N_8204,N_9068);
nor UO_1217 (O_1217,N_9700,N_8497);
or UO_1218 (O_1218,N_8924,N_9079);
nor UO_1219 (O_1219,N_9786,N_9357);
or UO_1220 (O_1220,N_8578,N_8210);
nor UO_1221 (O_1221,N_8113,N_8727);
nand UO_1222 (O_1222,N_9717,N_8758);
nand UO_1223 (O_1223,N_9780,N_8204);
or UO_1224 (O_1224,N_9663,N_9704);
or UO_1225 (O_1225,N_9675,N_8127);
nor UO_1226 (O_1226,N_9173,N_8207);
nand UO_1227 (O_1227,N_9702,N_9503);
and UO_1228 (O_1228,N_8965,N_9242);
nand UO_1229 (O_1229,N_8591,N_8403);
and UO_1230 (O_1230,N_8385,N_8753);
nor UO_1231 (O_1231,N_9340,N_9985);
or UO_1232 (O_1232,N_8090,N_8004);
nand UO_1233 (O_1233,N_8047,N_9987);
or UO_1234 (O_1234,N_8559,N_8341);
or UO_1235 (O_1235,N_9325,N_8278);
nand UO_1236 (O_1236,N_9715,N_9980);
nand UO_1237 (O_1237,N_8021,N_9389);
or UO_1238 (O_1238,N_9144,N_8213);
nand UO_1239 (O_1239,N_9751,N_8556);
nand UO_1240 (O_1240,N_9018,N_8139);
nor UO_1241 (O_1241,N_9899,N_8865);
and UO_1242 (O_1242,N_8301,N_9226);
nor UO_1243 (O_1243,N_9697,N_8376);
and UO_1244 (O_1244,N_8208,N_9037);
nand UO_1245 (O_1245,N_8688,N_9025);
nand UO_1246 (O_1246,N_9363,N_9315);
nand UO_1247 (O_1247,N_8120,N_9018);
nand UO_1248 (O_1248,N_9729,N_8593);
and UO_1249 (O_1249,N_9281,N_8557);
nor UO_1250 (O_1250,N_9975,N_9661);
and UO_1251 (O_1251,N_8267,N_9039);
nand UO_1252 (O_1252,N_8693,N_8169);
and UO_1253 (O_1253,N_9667,N_8101);
nor UO_1254 (O_1254,N_9158,N_8748);
or UO_1255 (O_1255,N_9601,N_9051);
or UO_1256 (O_1256,N_8981,N_8782);
nand UO_1257 (O_1257,N_9570,N_8045);
and UO_1258 (O_1258,N_8800,N_8056);
nand UO_1259 (O_1259,N_8310,N_9086);
and UO_1260 (O_1260,N_8693,N_9163);
and UO_1261 (O_1261,N_9482,N_8384);
nand UO_1262 (O_1262,N_8019,N_8669);
or UO_1263 (O_1263,N_8633,N_8423);
nand UO_1264 (O_1264,N_8334,N_9643);
nor UO_1265 (O_1265,N_9771,N_9922);
and UO_1266 (O_1266,N_8979,N_8232);
nand UO_1267 (O_1267,N_9057,N_8297);
or UO_1268 (O_1268,N_8445,N_9073);
nand UO_1269 (O_1269,N_9912,N_9236);
nand UO_1270 (O_1270,N_9703,N_9931);
nand UO_1271 (O_1271,N_8034,N_8914);
or UO_1272 (O_1272,N_9249,N_9751);
nand UO_1273 (O_1273,N_9144,N_9763);
nor UO_1274 (O_1274,N_9931,N_8957);
nand UO_1275 (O_1275,N_8367,N_8289);
nand UO_1276 (O_1276,N_9533,N_9992);
nand UO_1277 (O_1277,N_8886,N_9307);
nor UO_1278 (O_1278,N_8993,N_8734);
and UO_1279 (O_1279,N_9737,N_9580);
or UO_1280 (O_1280,N_9562,N_8766);
or UO_1281 (O_1281,N_9622,N_8254);
and UO_1282 (O_1282,N_9011,N_9687);
and UO_1283 (O_1283,N_9230,N_9110);
nor UO_1284 (O_1284,N_8154,N_8549);
or UO_1285 (O_1285,N_9003,N_8306);
nor UO_1286 (O_1286,N_8266,N_9896);
nand UO_1287 (O_1287,N_8745,N_9233);
nand UO_1288 (O_1288,N_8173,N_8986);
nor UO_1289 (O_1289,N_8386,N_9932);
and UO_1290 (O_1290,N_9322,N_8687);
nand UO_1291 (O_1291,N_8774,N_8659);
or UO_1292 (O_1292,N_9443,N_8622);
and UO_1293 (O_1293,N_8028,N_8182);
nor UO_1294 (O_1294,N_8700,N_9865);
nor UO_1295 (O_1295,N_8921,N_8044);
and UO_1296 (O_1296,N_9990,N_9066);
nor UO_1297 (O_1297,N_8023,N_8747);
and UO_1298 (O_1298,N_9355,N_9875);
nor UO_1299 (O_1299,N_9899,N_8808);
nand UO_1300 (O_1300,N_8059,N_9608);
and UO_1301 (O_1301,N_9662,N_9818);
nand UO_1302 (O_1302,N_8260,N_9252);
and UO_1303 (O_1303,N_9792,N_9199);
nor UO_1304 (O_1304,N_8517,N_9935);
and UO_1305 (O_1305,N_8373,N_9194);
nand UO_1306 (O_1306,N_8108,N_8240);
nor UO_1307 (O_1307,N_8663,N_9705);
or UO_1308 (O_1308,N_8187,N_9103);
nand UO_1309 (O_1309,N_8201,N_9493);
and UO_1310 (O_1310,N_9015,N_9637);
or UO_1311 (O_1311,N_8606,N_9241);
or UO_1312 (O_1312,N_9409,N_8231);
nand UO_1313 (O_1313,N_8095,N_8737);
and UO_1314 (O_1314,N_8666,N_9283);
or UO_1315 (O_1315,N_8657,N_8077);
and UO_1316 (O_1316,N_8054,N_9699);
and UO_1317 (O_1317,N_8157,N_9839);
or UO_1318 (O_1318,N_9842,N_9028);
nand UO_1319 (O_1319,N_9699,N_9045);
or UO_1320 (O_1320,N_9759,N_9855);
or UO_1321 (O_1321,N_9610,N_8976);
nor UO_1322 (O_1322,N_9307,N_8150);
or UO_1323 (O_1323,N_9499,N_9383);
or UO_1324 (O_1324,N_8412,N_8984);
nor UO_1325 (O_1325,N_8318,N_8592);
nor UO_1326 (O_1326,N_8484,N_8428);
or UO_1327 (O_1327,N_8454,N_8305);
nor UO_1328 (O_1328,N_9423,N_8308);
nand UO_1329 (O_1329,N_9855,N_9567);
and UO_1330 (O_1330,N_8479,N_9413);
nor UO_1331 (O_1331,N_9687,N_8832);
nor UO_1332 (O_1332,N_9304,N_8361);
nor UO_1333 (O_1333,N_9916,N_8035);
and UO_1334 (O_1334,N_9006,N_8704);
nor UO_1335 (O_1335,N_9988,N_8143);
or UO_1336 (O_1336,N_8356,N_8211);
nand UO_1337 (O_1337,N_9611,N_8587);
or UO_1338 (O_1338,N_9915,N_8306);
or UO_1339 (O_1339,N_9380,N_9063);
nand UO_1340 (O_1340,N_9166,N_8950);
nor UO_1341 (O_1341,N_8251,N_8630);
nand UO_1342 (O_1342,N_8395,N_8464);
nand UO_1343 (O_1343,N_9663,N_8658);
nand UO_1344 (O_1344,N_9760,N_8779);
nor UO_1345 (O_1345,N_9380,N_8496);
nand UO_1346 (O_1346,N_8196,N_9878);
nor UO_1347 (O_1347,N_9500,N_9810);
nand UO_1348 (O_1348,N_8787,N_8059);
or UO_1349 (O_1349,N_8690,N_9485);
nor UO_1350 (O_1350,N_8424,N_9366);
and UO_1351 (O_1351,N_8758,N_9233);
nor UO_1352 (O_1352,N_9148,N_9911);
and UO_1353 (O_1353,N_9231,N_8341);
nor UO_1354 (O_1354,N_9879,N_8745);
and UO_1355 (O_1355,N_8592,N_8449);
or UO_1356 (O_1356,N_8302,N_9901);
and UO_1357 (O_1357,N_8465,N_8001);
and UO_1358 (O_1358,N_9830,N_8227);
nand UO_1359 (O_1359,N_9069,N_9779);
xnor UO_1360 (O_1360,N_9715,N_8440);
and UO_1361 (O_1361,N_9711,N_9680);
and UO_1362 (O_1362,N_8772,N_9762);
nand UO_1363 (O_1363,N_9387,N_8983);
or UO_1364 (O_1364,N_9947,N_8616);
nand UO_1365 (O_1365,N_8094,N_9043);
nor UO_1366 (O_1366,N_9558,N_9952);
and UO_1367 (O_1367,N_9902,N_8616);
or UO_1368 (O_1368,N_8440,N_8198);
nor UO_1369 (O_1369,N_8316,N_9733);
or UO_1370 (O_1370,N_9425,N_9846);
and UO_1371 (O_1371,N_9234,N_8074);
and UO_1372 (O_1372,N_9653,N_8388);
or UO_1373 (O_1373,N_8447,N_9966);
nor UO_1374 (O_1374,N_8921,N_9016);
nor UO_1375 (O_1375,N_8860,N_9226);
nor UO_1376 (O_1376,N_8425,N_9535);
nand UO_1377 (O_1377,N_9543,N_8616);
and UO_1378 (O_1378,N_8669,N_8323);
and UO_1379 (O_1379,N_9534,N_9919);
nor UO_1380 (O_1380,N_8979,N_8313);
or UO_1381 (O_1381,N_8433,N_8274);
nor UO_1382 (O_1382,N_9760,N_9041);
nand UO_1383 (O_1383,N_9759,N_9889);
and UO_1384 (O_1384,N_8806,N_8869);
and UO_1385 (O_1385,N_9756,N_8201);
or UO_1386 (O_1386,N_9250,N_9256);
and UO_1387 (O_1387,N_9405,N_9037);
and UO_1388 (O_1388,N_8597,N_9673);
nand UO_1389 (O_1389,N_8923,N_8387);
nor UO_1390 (O_1390,N_8966,N_9180);
and UO_1391 (O_1391,N_8036,N_8964);
or UO_1392 (O_1392,N_9783,N_9386);
nand UO_1393 (O_1393,N_9044,N_8593);
nor UO_1394 (O_1394,N_8753,N_9855);
nor UO_1395 (O_1395,N_9946,N_9358);
nand UO_1396 (O_1396,N_8043,N_9541);
and UO_1397 (O_1397,N_8274,N_8774);
xnor UO_1398 (O_1398,N_8182,N_8444);
nor UO_1399 (O_1399,N_8919,N_9193);
nor UO_1400 (O_1400,N_9753,N_9732);
or UO_1401 (O_1401,N_9915,N_8041);
or UO_1402 (O_1402,N_9781,N_8410);
and UO_1403 (O_1403,N_8412,N_8132);
and UO_1404 (O_1404,N_9857,N_8873);
and UO_1405 (O_1405,N_9180,N_9725);
and UO_1406 (O_1406,N_8449,N_9803);
nor UO_1407 (O_1407,N_9292,N_9145);
and UO_1408 (O_1408,N_8782,N_9592);
nor UO_1409 (O_1409,N_8046,N_8392);
nor UO_1410 (O_1410,N_8552,N_8936);
or UO_1411 (O_1411,N_9695,N_8046);
nor UO_1412 (O_1412,N_8304,N_9974);
nor UO_1413 (O_1413,N_9829,N_8120);
nor UO_1414 (O_1414,N_9732,N_8724);
and UO_1415 (O_1415,N_8470,N_9789);
or UO_1416 (O_1416,N_8759,N_8024);
nor UO_1417 (O_1417,N_9075,N_8371);
or UO_1418 (O_1418,N_8706,N_8601);
or UO_1419 (O_1419,N_8660,N_9756);
and UO_1420 (O_1420,N_9914,N_8168);
nand UO_1421 (O_1421,N_8121,N_8917);
nand UO_1422 (O_1422,N_8989,N_8297);
nand UO_1423 (O_1423,N_8323,N_8542);
nand UO_1424 (O_1424,N_8744,N_9073);
nor UO_1425 (O_1425,N_8686,N_8226);
and UO_1426 (O_1426,N_9560,N_9266);
or UO_1427 (O_1427,N_9483,N_8556);
nand UO_1428 (O_1428,N_9835,N_8960);
and UO_1429 (O_1429,N_8294,N_9014);
nand UO_1430 (O_1430,N_9292,N_8800);
or UO_1431 (O_1431,N_9325,N_9023);
or UO_1432 (O_1432,N_9355,N_9972);
nor UO_1433 (O_1433,N_8140,N_8692);
and UO_1434 (O_1434,N_9626,N_8773);
or UO_1435 (O_1435,N_8139,N_9134);
and UO_1436 (O_1436,N_9590,N_8131);
and UO_1437 (O_1437,N_9395,N_8408);
nand UO_1438 (O_1438,N_9787,N_9798);
nand UO_1439 (O_1439,N_9463,N_8904);
or UO_1440 (O_1440,N_8347,N_8337);
and UO_1441 (O_1441,N_8657,N_9554);
nor UO_1442 (O_1442,N_8186,N_8433);
nand UO_1443 (O_1443,N_8222,N_8256);
or UO_1444 (O_1444,N_8280,N_9475);
nand UO_1445 (O_1445,N_8368,N_8473);
and UO_1446 (O_1446,N_8975,N_9551);
and UO_1447 (O_1447,N_8401,N_8084);
or UO_1448 (O_1448,N_9992,N_9628);
nand UO_1449 (O_1449,N_8173,N_8121);
nand UO_1450 (O_1450,N_8046,N_8985);
nor UO_1451 (O_1451,N_8974,N_8004);
and UO_1452 (O_1452,N_9867,N_9304);
nor UO_1453 (O_1453,N_9284,N_9588);
nor UO_1454 (O_1454,N_9999,N_8403);
and UO_1455 (O_1455,N_9785,N_9355);
nor UO_1456 (O_1456,N_8898,N_8647);
and UO_1457 (O_1457,N_9487,N_9177);
or UO_1458 (O_1458,N_8328,N_9634);
or UO_1459 (O_1459,N_8282,N_8566);
or UO_1460 (O_1460,N_9451,N_9342);
nand UO_1461 (O_1461,N_8612,N_9193);
or UO_1462 (O_1462,N_9715,N_9860);
nor UO_1463 (O_1463,N_9556,N_9236);
or UO_1464 (O_1464,N_9240,N_9664);
and UO_1465 (O_1465,N_8824,N_8973);
and UO_1466 (O_1466,N_8354,N_8289);
and UO_1467 (O_1467,N_8049,N_9224);
and UO_1468 (O_1468,N_9300,N_8649);
and UO_1469 (O_1469,N_9186,N_9532);
or UO_1470 (O_1470,N_9509,N_8211);
nor UO_1471 (O_1471,N_8847,N_8236);
and UO_1472 (O_1472,N_8673,N_8077);
nor UO_1473 (O_1473,N_8723,N_9485);
and UO_1474 (O_1474,N_8529,N_8990);
and UO_1475 (O_1475,N_9805,N_9898);
nand UO_1476 (O_1476,N_8578,N_8849);
or UO_1477 (O_1477,N_8268,N_8709);
nand UO_1478 (O_1478,N_9332,N_9075);
or UO_1479 (O_1479,N_9103,N_9333);
nor UO_1480 (O_1480,N_9871,N_8982);
or UO_1481 (O_1481,N_8808,N_8688);
and UO_1482 (O_1482,N_9268,N_8368);
and UO_1483 (O_1483,N_9092,N_9663);
or UO_1484 (O_1484,N_9790,N_9582);
and UO_1485 (O_1485,N_8549,N_9394);
nand UO_1486 (O_1486,N_8523,N_8940);
xnor UO_1487 (O_1487,N_9773,N_9463);
and UO_1488 (O_1488,N_8256,N_8459);
nor UO_1489 (O_1489,N_8784,N_8430);
nand UO_1490 (O_1490,N_9183,N_9217);
nor UO_1491 (O_1491,N_9784,N_9073);
nand UO_1492 (O_1492,N_9361,N_9887);
nand UO_1493 (O_1493,N_8826,N_8233);
nand UO_1494 (O_1494,N_8599,N_9185);
and UO_1495 (O_1495,N_9105,N_8766);
or UO_1496 (O_1496,N_9960,N_8288);
nand UO_1497 (O_1497,N_8995,N_9929);
and UO_1498 (O_1498,N_9328,N_8432);
and UO_1499 (O_1499,N_9897,N_9667);
endmodule