module basic_3000_30000_3500_10_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2916,In_1535);
nand U1 (N_1,In_1959,In_652);
nand U2 (N_2,In_1313,In_1642);
nand U3 (N_3,In_243,In_1661);
or U4 (N_4,In_1629,In_2389);
and U5 (N_5,In_398,In_2705);
and U6 (N_6,In_1148,In_2503);
or U7 (N_7,In_2461,In_1391);
nor U8 (N_8,In_376,In_2100);
nor U9 (N_9,In_1737,In_2787);
xor U10 (N_10,In_2774,In_374);
nor U11 (N_11,In_1695,In_656);
and U12 (N_12,In_425,In_1668);
nor U13 (N_13,In_117,In_2020);
or U14 (N_14,In_2628,In_779);
nor U15 (N_15,In_1736,In_1281);
or U16 (N_16,In_1404,In_2475);
xor U17 (N_17,In_1303,In_483);
xnor U18 (N_18,In_1713,In_2026);
and U19 (N_19,In_513,In_1447);
xor U20 (N_20,In_2487,In_862);
or U21 (N_21,In_1178,In_2947);
nor U22 (N_22,In_2945,In_844);
nand U23 (N_23,In_2647,In_67);
nand U24 (N_24,In_409,In_90);
xnor U25 (N_25,In_172,In_2871);
or U26 (N_26,In_2108,In_944);
or U27 (N_27,In_2374,In_1788);
or U28 (N_28,In_2930,In_2239);
xnor U29 (N_29,In_1009,In_879);
or U30 (N_30,In_882,In_1089);
nor U31 (N_31,In_556,In_53);
and U32 (N_32,In_263,In_1314);
nand U33 (N_33,In_208,In_987);
and U34 (N_34,In_2229,In_1651);
and U35 (N_35,In_2394,In_1115);
and U36 (N_36,In_480,In_1613);
and U37 (N_37,In_1809,In_1222);
xor U38 (N_38,In_871,In_1674);
nor U39 (N_39,In_1769,In_996);
xnor U40 (N_40,In_337,In_2580);
nor U41 (N_41,In_519,In_2114);
nand U42 (N_42,In_2614,In_2941);
and U43 (N_43,In_2755,In_285);
nor U44 (N_44,In_1011,In_517);
nor U45 (N_45,In_1251,In_1531);
nand U46 (N_46,In_1263,In_1210);
or U47 (N_47,In_1658,In_123);
and U48 (N_48,In_2934,In_1026);
xnor U49 (N_49,In_2134,In_981);
nand U50 (N_50,In_258,In_2791);
xnor U51 (N_51,In_1446,In_2306);
and U52 (N_52,In_2967,In_651);
nand U53 (N_53,In_1854,In_2397);
and U54 (N_54,In_2135,In_1073);
and U55 (N_55,In_1352,In_38);
xor U56 (N_56,In_12,In_2595);
and U57 (N_57,In_2543,In_1338);
nor U58 (N_58,In_941,In_2081);
nand U59 (N_59,In_2340,In_709);
nor U60 (N_60,In_1064,In_649);
and U61 (N_61,In_2384,In_1364);
and U62 (N_62,In_1897,In_420);
xor U63 (N_63,In_2506,In_2619);
or U64 (N_64,In_1253,In_1509);
xor U65 (N_65,In_2055,In_288);
xnor U66 (N_66,In_643,In_1424);
nor U67 (N_67,In_2679,In_892);
and U68 (N_68,In_802,In_2817);
nor U69 (N_69,In_1866,In_2611);
nor U70 (N_70,In_1533,In_1716);
nor U71 (N_71,In_1728,In_771);
or U72 (N_72,In_973,In_1987);
nand U73 (N_73,In_1324,In_1955);
or U74 (N_74,In_2436,In_1905);
or U75 (N_75,In_590,In_2470);
or U76 (N_76,In_1259,In_2914);
and U77 (N_77,In_2594,In_1687);
nor U78 (N_78,In_2836,In_2039);
nor U79 (N_79,In_1326,In_1800);
nor U80 (N_80,In_1031,In_188);
or U81 (N_81,In_378,In_1407);
nand U82 (N_82,In_2865,In_1885);
and U83 (N_83,In_849,In_2471);
xor U84 (N_84,In_1903,In_2726);
and U85 (N_85,In_1135,In_2180);
or U86 (N_86,In_2280,In_1168);
nand U87 (N_87,In_1720,In_2735);
xor U88 (N_88,In_685,In_1308);
nor U89 (N_89,In_1577,In_502);
nor U90 (N_90,In_413,In_1305);
nand U91 (N_91,In_1467,In_1504);
nor U92 (N_92,In_2604,In_2783);
nand U93 (N_93,In_522,In_865);
xnor U94 (N_94,In_274,In_1193);
and U95 (N_95,In_2222,In_136);
xor U96 (N_96,In_16,In_536);
or U97 (N_97,In_2145,In_568);
nand U98 (N_98,In_195,In_562);
or U99 (N_99,In_782,In_2017);
or U100 (N_100,In_1244,In_2396);
xnor U101 (N_101,In_2237,In_2042);
or U102 (N_102,In_229,In_1553);
and U103 (N_103,In_106,In_1611);
or U104 (N_104,In_1512,In_1933);
nor U105 (N_105,In_881,In_2303);
xnor U106 (N_106,In_2953,In_1254);
and U107 (N_107,In_189,In_2191);
nor U108 (N_108,In_1798,In_2887);
or U109 (N_109,In_1237,In_1890);
nor U110 (N_110,In_2187,In_868);
nor U111 (N_111,In_2868,In_164);
or U112 (N_112,In_569,In_2944);
nand U113 (N_113,In_2313,In_564);
xor U114 (N_114,In_2176,In_1264);
nor U115 (N_115,In_1370,In_2546);
nand U116 (N_116,In_1057,In_610);
xnor U117 (N_117,In_2172,In_1335);
or U118 (N_118,In_1300,In_2109);
and U119 (N_119,In_873,In_63);
or U120 (N_120,In_1449,In_2927);
nand U121 (N_121,In_226,In_2491);
xor U122 (N_122,In_1302,In_1567);
and U123 (N_123,In_2955,In_2716);
xor U124 (N_124,In_1097,In_2830);
xor U125 (N_125,In_2202,In_1060);
and U126 (N_126,In_2124,In_88);
and U127 (N_127,In_283,In_1498);
nand U128 (N_128,In_877,In_746);
nand U129 (N_129,In_321,In_2008);
nand U130 (N_130,In_2365,In_410);
nand U131 (N_131,In_1102,In_487);
nor U132 (N_132,In_2300,In_1350);
nand U133 (N_133,In_199,In_516);
or U134 (N_134,In_2088,In_1831);
nor U135 (N_135,In_670,In_1018);
xnor U136 (N_136,In_352,In_560);
nand U137 (N_137,In_1765,In_1950);
xnor U138 (N_138,In_2906,In_870);
nand U139 (N_139,In_2210,In_2957);
nor U140 (N_140,In_2336,In_2304);
and U141 (N_141,In_1941,In_888);
nor U142 (N_142,In_1922,In_490);
or U143 (N_143,In_393,In_1956);
nand U144 (N_144,In_441,In_1960);
and U145 (N_145,In_626,In_295);
and U146 (N_146,In_2578,In_2096);
nor U147 (N_147,In_2767,In_2213);
and U148 (N_148,In_1369,In_2203);
xnor U149 (N_149,In_886,In_693);
nor U150 (N_150,In_1228,In_1319);
and U151 (N_151,In_170,In_24);
nand U152 (N_152,In_317,In_2810);
nand U153 (N_153,In_1667,In_676);
nor U154 (N_154,In_2666,In_1639);
nand U155 (N_155,In_2056,In_2936);
or U156 (N_156,In_132,In_1094);
or U157 (N_157,In_311,In_1562);
xor U158 (N_158,In_2035,In_2201);
or U159 (N_159,In_2334,In_2902);
nand U160 (N_160,In_2411,In_1571);
and U161 (N_161,In_765,In_1276);
xor U162 (N_162,In_201,In_2965);
or U163 (N_163,In_2282,In_1612);
nor U164 (N_164,In_1807,In_819);
or U165 (N_165,In_2036,In_2713);
or U166 (N_166,In_2922,In_2472);
or U167 (N_167,In_127,In_2601);
or U168 (N_168,In_2708,In_1721);
nor U169 (N_169,In_34,In_1939);
or U170 (N_170,In_234,In_237);
nand U171 (N_171,In_244,In_2691);
or U172 (N_172,In_2466,In_2177);
xor U173 (N_173,In_2861,In_1564);
xor U174 (N_174,In_2740,In_157);
or U175 (N_175,In_2241,In_1213);
nand U176 (N_176,In_2801,In_2525);
nand U177 (N_177,In_402,In_277);
and U178 (N_178,In_2169,In_1755);
and U179 (N_179,In_2577,In_1093);
xnor U180 (N_180,In_1828,In_2463);
or U181 (N_181,In_1545,In_783);
nor U182 (N_182,In_1005,In_1241);
or U183 (N_183,In_667,In_2084);
xor U184 (N_184,In_1991,In_354);
nand U185 (N_185,In_2523,In_322);
nor U186 (N_186,In_330,In_2478);
nand U187 (N_187,In_1332,In_1988);
nand U188 (N_188,In_1006,In_2949);
nand U189 (N_189,In_2845,In_2843);
or U190 (N_190,In_426,In_512);
xnor U191 (N_191,In_642,In_2984);
nor U192 (N_192,In_2058,In_1110);
nor U193 (N_193,In_1059,In_2481);
nor U194 (N_194,In_156,In_1621);
nand U195 (N_195,In_2698,In_1990);
nor U196 (N_196,In_1231,In_1707);
xnor U197 (N_197,In_1017,In_141);
and U198 (N_198,In_1596,In_1212);
or U199 (N_199,In_2988,In_2004);
xnor U200 (N_200,In_723,In_163);
and U201 (N_201,In_1749,In_2003);
nor U202 (N_202,In_2188,In_1678);
nor U203 (N_203,In_2414,In_436);
nor U204 (N_204,In_1969,In_2391);
and U205 (N_205,In_1069,In_1789);
or U206 (N_206,In_1206,In_2355);
nand U207 (N_207,In_460,In_1224);
nor U208 (N_208,In_366,In_1588);
and U209 (N_209,In_2428,In_242);
or U210 (N_210,In_1341,In_1365);
xor U211 (N_211,In_2924,In_2328);
and U212 (N_212,In_991,In_635);
or U213 (N_213,In_2321,In_2119);
xnor U214 (N_214,In_271,In_2551);
nor U215 (N_215,In_2590,In_1188);
and U216 (N_216,In_1908,In_2878);
xnor U217 (N_217,In_798,In_2370);
nand U218 (N_218,In_617,In_546);
and U219 (N_219,In_1310,In_2269);
xor U220 (N_220,In_2083,In_903);
xor U221 (N_221,In_2331,In_995);
nand U222 (N_222,In_2163,In_1655);
nand U223 (N_223,In_159,In_2676);
xnor U224 (N_224,In_843,In_1849);
nor U225 (N_225,In_2102,In_687);
xor U226 (N_226,In_1007,In_2009);
or U227 (N_227,In_1420,In_583);
nor U228 (N_228,In_857,In_2979);
nand U229 (N_229,In_1479,In_2970);
and U230 (N_230,In_1132,In_2447);
nor U231 (N_231,In_815,In_2655);
nor U232 (N_232,In_47,In_61);
and U233 (N_233,In_2013,In_2717);
nand U234 (N_234,In_1551,In_1899);
and U235 (N_235,In_1130,In_1992);
and U236 (N_236,In_2153,In_1438);
nor U237 (N_237,In_362,In_228);
xor U238 (N_238,In_2136,In_1848);
or U239 (N_239,In_1811,In_2405);
nor U240 (N_240,In_1693,In_35);
or U241 (N_241,In_30,In_457);
or U242 (N_242,In_1563,In_412);
nor U243 (N_243,In_2854,In_2996);
nor U244 (N_244,In_2521,In_2777);
and U245 (N_245,In_2443,In_1200);
and U246 (N_246,In_2657,In_1619);
or U247 (N_247,In_2950,In_262);
xor U248 (N_248,In_301,In_1714);
nand U249 (N_249,In_2693,In_2770);
nand U250 (N_250,In_1706,In_1403);
nand U251 (N_251,In_2120,In_2236);
and U252 (N_252,In_1247,In_2077);
and U253 (N_253,In_1123,In_1748);
or U254 (N_254,In_1850,In_668);
and U255 (N_255,In_98,In_853);
nor U256 (N_256,In_1670,In_2792);
and U257 (N_257,In_2536,In_1436);
and U258 (N_258,In_1902,In_1480);
or U259 (N_259,In_2294,In_2442);
nand U260 (N_260,In_1034,In_68);
nand U261 (N_261,In_2168,In_2759);
nand U262 (N_262,In_2274,In_1919);
nand U263 (N_263,In_681,In_2966);
nor U264 (N_264,In_922,In_2732);
and U265 (N_265,In_1785,In_2803);
and U266 (N_266,In_1511,In_138);
and U267 (N_267,In_920,In_1355);
nand U268 (N_268,In_909,In_83);
and U269 (N_269,In_2449,In_2508);
and U270 (N_270,In_1782,In_2040);
xnor U271 (N_271,In_2179,In_2681);
or U272 (N_272,In_2221,In_2931);
nand U273 (N_273,In_225,In_1245);
and U274 (N_274,In_1043,In_764);
xnor U275 (N_275,In_1208,In_2510);
and U276 (N_276,In_1382,In_145);
or U277 (N_277,In_606,In_2011);
nor U278 (N_278,In_2403,In_2060);
xor U279 (N_279,In_1151,In_1746);
nor U280 (N_280,In_461,In_1595);
nand U281 (N_281,In_2171,In_1537);
or U282 (N_282,In_2524,In_1523);
or U283 (N_283,In_2069,In_608);
xnor U284 (N_284,In_1426,In_1062);
nor U285 (N_285,In_674,In_925);
or U286 (N_286,In_1842,In_2633);
nor U287 (N_287,In_2502,In_2107);
xnor U288 (N_288,In_2653,In_1602);
xnor U289 (N_289,In_2820,In_2568);
or U290 (N_290,In_2976,In_2884);
or U291 (N_291,In_73,In_1176);
nand U292 (N_292,In_218,In_789);
and U293 (N_293,In_1121,In_291);
nand U294 (N_294,In_1218,In_1260);
nor U295 (N_295,In_1895,In_2634);
or U296 (N_296,In_206,In_1702);
or U297 (N_297,In_700,In_1004);
and U298 (N_298,In_767,In_496);
xnor U299 (N_299,In_718,In_2702);
xnor U300 (N_300,In_1569,In_497);
xor U301 (N_301,In_1593,In_2287);
or U302 (N_302,In_548,In_680);
nor U303 (N_303,In_2127,In_1656);
xnor U304 (N_304,In_2807,In_2562);
nand U305 (N_305,In_74,In_1943);
nor U306 (N_306,In_712,In_209);
nand U307 (N_307,In_846,In_1853);
and U308 (N_308,In_1764,In_278);
or U309 (N_309,In_2413,In_1934);
nor U310 (N_310,In_1843,In_1795);
and U311 (N_311,In_808,In_1700);
xor U312 (N_312,In_1677,In_2099);
xnor U313 (N_313,In_1050,In_81);
xor U314 (N_314,In_2962,In_2110);
or U315 (N_315,In_1106,In_761);
or U316 (N_316,In_1376,In_382);
nand U317 (N_317,In_251,In_2641);
or U318 (N_318,In_150,In_1835);
or U319 (N_319,In_1876,In_2790);
nor U320 (N_320,In_1672,In_272);
nor U321 (N_321,In_2369,In_1771);
nand U322 (N_322,In_1232,In_2105);
or U323 (N_323,In_1662,In_2122);
and U324 (N_324,In_2227,In_912);
or U325 (N_325,In_1779,In_600);
nor U326 (N_326,In_2245,In_1858);
and U327 (N_327,In_1035,In_2);
nor U328 (N_328,In_1286,In_1078);
nor U329 (N_329,In_683,In_1703);
xor U330 (N_330,In_1126,In_2046);
or U331 (N_331,In_2821,In_84);
xor U332 (N_332,In_40,In_596);
xnor U333 (N_333,In_193,In_439);
and U334 (N_334,In_2881,In_2349);
and U335 (N_335,In_1023,In_2812);
nand U336 (N_336,In_1780,In_1543);
and U337 (N_337,In_790,In_1174);
nor U338 (N_338,In_1267,In_2430);
xnor U339 (N_339,In_1898,In_986);
and U340 (N_340,In_840,In_1353);
or U341 (N_341,In_2452,In_1490);
xnor U342 (N_342,In_2637,In_1615);
nor U343 (N_343,In_2215,In_2429);
nor U344 (N_344,In_2724,In_889);
and U345 (N_345,In_1336,In_1143);
xor U346 (N_346,In_2768,In_694);
or U347 (N_347,In_2247,In_1647);
and U348 (N_348,In_1773,In_2322);
or U349 (N_349,In_954,In_452);
or U350 (N_350,In_1568,In_1565);
and U351 (N_351,In_1698,In_725);
and U352 (N_352,In_144,In_942);
and U353 (N_353,In_890,In_2549);
nor U354 (N_354,In_1650,In_324);
nand U355 (N_355,In_1405,In_17);
or U356 (N_356,In_264,In_2263);
and U357 (N_357,In_2901,In_983);
or U358 (N_358,In_1181,In_1603);
or U359 (N_359,In_2761,In_742);
or U360 (N_360,In_331,In_485);
or U361 (N_361,In_1972,In_1384);
and U362 (N_362,In_433,In_121);
and U363 (N_363,In_1673,In_1740);
xnor U364 (N_364,In_1195,In_2511);
and U365 (N_365,In_2174,In_137);
nor U366 (N_366,In_2123,In_1323);
or U367 (N_367,In_799,In_907);
or U368 (N_368,In_834,In_915);
and U369 (N_369,In_1989,In_508);
nor U370 (N_370,In_2029,In_2889);
nand U371 (N_371,In_1041,In_1327);
and U372 (N_372,In_155,In_589);
xor U373 (N_373,In_1344,In_2439);
xnor U374 (N_374,In_2454,In_1816);
and U375 (N_375,In_2231,In_148);
or U376 (N_376,In_2419,In_2954);
and U377 (N_377,In_259,In_974);
and U378 (N_378,In_151,In_2711);
nand U379 (N_379,In_1122,In_2893);
xor U380 (N_380,In_1648,In_1137);
xor U381 (N_381,In_1819,In_1817);
xnor U382 (N_382,In_268,In_1033);
xnor U383 (N_383,In_185,In_940);
xor U384 (N_384,In_917,In_514);
and U385 (N_385,In_2288,In_554);
and U386 (N_386,In_2599,In_1401);
and U387 (N_387,In_1024,In_2189);
nor U388 (N_388,In_133,In_1186);
xnor U389 (N_389,In_704,In_1844);
xnor U390 (N_390,In_2948,In_328);
nand U391 (N_391,In_1040,In_1362);
nand U392 (N_392,In_1832,In_221);
nand U393 (N_393,In_2353,In_1032);
and U394 (N_394,In_386,In_2271);
xor U395 (N_395,In_2886,In_1628);
nor U396 (N_396,In_2789,In_740);
nand U397 (N_397,In_2728,In_1464);
nor U398 (N_398,In_2857,In_2284);
and U399 (N_399,In_2410,In_1875);
nor U400 (N_400,In_2438,In_966);
and U401 (N_401,In_469,In_855);
xor U402 (N_402,In_1501,In_2087);
and U403 (N_403,In_650,In_22);
nor U404 (N_404,In_87,In_1730);
and U405 (N_405,In_355,In_970);
or U406 (N_406,In_1189,In_120);
and U407 (N_407,In_139,In_692);
nor U408 (N_408,In_1957,In_196);
xor U409 (N_409,In_2824,In_2279);
nor U410 (N_410,In_1869,In_1701);
or U411 (N_411,In_1010,In_171);
or U412 (N_412,In_55,In_2785);
and U413 (N_413,In_309,In_158);
nor U414 (N_414,In_1086,In_2943);
and U415 (N_415,In_2880,In_1691);
nand U416 (N_416,In_66,In_1521);
xor U417 (N_417,In_1469,In_609);
and U418 (N_418,In_1125,In_1081);
nor U419 (N_419,In_520,In_1830);
nor U420 (N_420,In_2904,In_975);
xor U421 (N_421,In_2827,In_0);
nand U422 (N_422,In_2952,In_182);
and U423 (N_423,In_2704,In_2507);
nor U424 (N_424,In_2217,In_2368);
and U425 (N_425,In_2618,In_1325);
or U426 (N_426,In_2129,In_1165);
nor U427 (N_427,In_1888,In_887);
xor U428 (N_428,In_774,In_766);
or U429 (N_429,In_1645,In_2675);
or U430 (N_430,In_2648,In_306);
nand U431 (N_431,In_1578,In_2686);
nand U432 (N_432,In_1552,In_1095);
nand U433 (N_433,In_2908,In_2453);
xor U434 (N_434,In_813,In_2951);
or U435 (N_435,In_1383,In_2106);
or U436 (N_436,In_2603,In_760);
xor U437 (N_437,In_584,In_2645);
or U438 (N_438,In_2341,In_2152);
nand U439 (N_439,In_1297,In_2866);
nand U440 (N_440,In_2720,In_678);
xor U441 (N_441,In_1710,In_1256);
xnor U442 (N_442,In_1643,In_1105);
xnor U443 (N_443,In_1725,In_821);
or U444 (N_444,In_607,In_1560);
or U445 (N_445,In_1731,In_1522);
nor U446 (N_446,In_817,In_1754);
nand U447 (N_447,In_2401,In_1907);
nand U448 (N_448,In_851,In_414);
xor U449 (N_449,In_1534,In_602);
xnor U450 (N_450,In_1374,In_1191);
xnor U451 (N_451,In_1952,In_2572);
nand U452 (N_452,In_464,In_679);
or U453 (N_453,In_1409,In_775);
xor U454 (N_454,In_473,In_1294);
or U455 (N_455,In_1851,In_2305);
or U456 (N_456,In_112,In_1282);
nand U457 (N_457,In_533,In_2598);
nand U458 (N_458,In_2513,In_95);
or U459 (N_459,In_2072,In_741);
and U460 (N_460,In_2367,In_1269);
or U461 (N_461,In_937,In_2778);
xnor U462 (N_462,In_2052,In_1676);
nor U463 (N_463,In_2905,In_1275);
nor U464 (N_464,In_270,In_1279);
or U465 (N_465,In_2261,In_2749);
xor U466 (N_466,In_1584,In_361);
nor U467 (N_467,In_1170,In_1995);
and U468 (N_468,In_1711,In_168);
nor U469 (N_469,In_421,In_273);
or U470 (N_470,In_1708,In_2170);
xor U471 (N_471,In_72,In_2900);
and U472 (N_472,In_178,In_2671);
xor U473 (N_473,In_2208,In_2356);
or U474 (N_474,In_26,In_282);
nor U475 (N_475,In_1145,In_1020);
or U476 (N_476,In_2547,In_1538);
xor U477 (N_477,In_1975,In_1088);
and U478 (N_478,In_686,In_856);
nand U479 (N_479,In_2157,In_1872);
nor U480 (N_480,In_192,In_2486);
or U481 (N_481,In_2347,In_754);
and U482 (N_482,In_347,In_978);
and U483 (N_483,In_2192,In_2677);
xnor U484 (N_484,In_1519,In_806);
xor U485 (N_485,In_1169,In_2381);
nor U486 (N_486,In_2346,In_1378);
nand U487 (N_487,In_729,In_919);
nor U488 (N_488,In_1961,In_1547);
nor U489 (N_489,In_861,In_2094);
or U490 (N_490,In_1753,In_875);
and U491 (N_491,In_2316,In_1823);
nand U492 (N_492,In_85,In_216);
nand U493 (N_493,In_1966,In_507);
nor U494 (N_494,In_2842,In_364);
and U495 (N_495,In_599,In_2876);
xor U496 (N_496,In_1249,In_2548);
nor U497 (N_497,In_2051,In_1164);
nor U498 (N_498,In_1894,In_854);
nand U499 (N_499,In_2998,In_2786);
and U500 (N_500,In_699,In_438);
and U501 (N_501,In_1483,In_567);
or U502 (N_502,In_2849,In_2493);
nor U503 (N_503,In_408,In_358);
xnor U504 (N_504,In_1075,In_2492);
and U505 (N_505,In_504,In_404);
xor U506 (N_506,In_238,In_2710);
xnor U507 (N_507,In_89,In_416);
and U508 (N_508,In_1309,In_2923);
or U509 (N_509,In_2186,In_491);
and U510 (N_510,In_988,In_2024);
xor U511 (N_511,In_800,In_175);
and U512 (N_512,In_211,In_2339);
or U513 (N_513,In_2632,In_1432);
xnor U514 (N_514,In_1421,In_344);
xor U515 (N_515,In_648,In_1320);
nor U516 (N_516,In_1932,In_1246);
and U517 (N_517,In_2065,In_1235);
xnor U518 (N_518,In_25,In_597);
and U519 (N_519,In_1915,In_2097);
and U520 (N_520,In_1312,In_918);
nor U521 (N_521,In_1532,In_757);
nor U522 (N_522,In_869,In_1390);
nand U523 (N_523,In_1864,In_2804);
and U524 (N_524,In_734,In_1394);
nand U525 (N_525,In_1455,In_2680);
nand U526 (N_526,In_2469,In_1167);
nand U527 (N_527,In_2223,In_1221);
nand U528 (N_528,In_2038,In_542);
and U529 (N_529,In_1462,In_1425);
nand U530 (N_530,In_1608,In_1722);
or U531 (N_531,In_2027,In_1794);
and U532 (N_532,In_302,In_129);
or U533 (N_533,In_1234,In_1417);
and U534 (N_534,In_2918,In_777);
nand U535 (N_535,In_2075,In_748);
xnor U536 (N_536,In_1014,In_1022);
nand U537 (N_537,In_99,In_1289);
nor U538 (N_538,In_1217,In_2850);
nand U539 (N_539,In_2654,In_2620);
or U540 (N_540,In_1496,In_2366);
xor U541 (N_541,In_2932,In_2023);
and U542 (N_542,In_1696,In_2561);
nand U543 (N_543,In_2813,In_1227);
and U544 (N_544,In_751,In_2407);
xnor U545 (N_545,In_2175,In_762);
and U546 (N_546,In_2769,In_743);
nand U547 (N_547,In_1739,In_2748);
and U548 (N_548,In_455,In_380);
and U549 (N_549,In_1723,In_2707);
xnor U550 (N_550,In_2393,In_2664);
xor U551 (N_551,In_1494,In_2142);
xor U552 (N_552,In_2352,In_479);
xnor U553 (N_553,In_2388,In_1630);
nor U554 (N_554,In_357,In_349);
or U555 (N_555,In_733,In_2883);
nand U556 (N_556,In_2545,In_2151);
nand U557 (N_557,In_1478,In_2797);
and U558 (N_558,In_10,In_1499);
nor U559 (N_559,In_621,In_695);
nor U560 (N_560,In_1389,In_1229);
xor U561 (N_561,In_1839,In_214);
and U562 (N_562,In_955,In_1986);
or U563 (N_563,In_2917,In_2616);
or U564 (N_564,In_629,In_1901);
xnor U565 (N_565,In_1160,In_2256);
and U566 (N_566,In_780,In_566);
xnor U567 (N_567,In_638,In_101);
nand U568 (N_568,In_2898,In_2007);
nand U569 (N_569,In_82,In_2053);
and U570 (N_570,In_1528,In_2362);
xor U571 (N_571,In_1859,In_1527);
or U572 (N_572,In_2556,In_2143);
xnor U573 (N_573,In_37,In_2412);
nor U574 (N_574,In_471,In_1318);
or U575 (N_575,In_1624,In_1171);
xnor U576 (N_576,In_2422,In_1127);
nor U577 (N_577,In_2101,In_493);
nand U578 (N_578,In_1418,In_280);
or U579 (N_579,In_1743,In_1813);
xnor U580 (N_580,In_2991,In_778);
xnor U581 (N_581,In_1845,In_64);
xnor U582 (N_582,In_2054,In_2833);
or U583 (N_583,In_2515,In_2141);
and U584 (N_584,In_1574,In_1556);
nor U585 (N_585,In_2435,In_721);
nor U586 (N_586,In_2650,In_57);
nor U587 (N_587,In_2621,In_763);
and U588 (N_588,In_2828,In_1985);
nand U589 (N_589,In_2037,In_1994);
or U590 (N_590,In_75,In_2796);
or U591 (N_591,In_669,In_2448);
nor U592 (N_592,In_2258,In_1087);
nor U593 (N_593,In_697,In_371);
or U594 (N_594,In_2385,In_1704);
and U595 (N_595,In_1393,In_671);
and U596 (N_596,In_575,In_1964);
nor U597 (N_597,In_2571,In_1451);
and U598 (N_598,In_339,In_1301);
nand U599 (N_599,In_104,In_2935);
xor U600 (N_600,In_558,In_1649);
and U601 (N_601,In_2763,In_858);
and U602 (N_602,In_230,In_2338);
nor U603 (N_603,In_1133,In_1640);
nor U604 (N_604,In_959,In_1453);
or U605 (N_605,In_1979,In_1042);
nand U606 (N_606,In_2089,In_967);
nor U607 (N_607,In_2154,In_1016);
nand U608 (N_608,In_2668,In_499);
nand U609 (N_609,In_2684,In_1997);
nand U610 (N_610,In_2126,In_2196);
xor U611 (N_611,In_2567,In_1573);
xor U612 (N_612,In_902,In_475);
xnor U613 (N_613,In_604,In_2111);
nor U614 (N_614,In_662,In_820);
nand U615 (N_615,In_422,In_1692);
and U616 (N_616,In_710,In_2489);
nand U617 (N_617,In_60,In_916);
xor U618 (N_618,In_832,In_2651);
and U619 (N_619,In_759,In_624);
xor U620 (N_620,In_2554,In_835);
or U621 (N_621,In_2592,In_1607);
and U622 (N_622,In_1358,In_1818);
nor U623 (N_623,In_794,In_615);
and U624 (N_624,In_1949,In_1502);
and U625 (N_625,In_1946,In_368);
and U626 (N_626,In_2333,In_2073);
or U627 (N_627,In_11,In_1146);
xnor U628 (N_628,In_247,In_565);
and U629 (N_629,In_2267,In_552);
and U630 (N_630,In_2532,In_1141);
nand U631 (N_631,In_2474,In_152);
and U632 (N_632,In_1156,In_2289);
nor U633 (N_633,In_1576,In_2257);
nand U634 (N_634,In_2831,In_1250);
nand U635 (N_635,In_323,In_2344);
nor U636 (N_636,In_360,In_2589);
and U637 (N_637,In_2613,In_842);
nand U638 (N_638,In_281,In_429);
nand U639 (N_639,In_660,In_2663);
xor U640 (N_640,In_1974,In_246);
xor U641 (N_641,In_1202,In_2315);
and U642 (N_642,In_1295,In_1416);
nor U643 (N_643,In_831,In_1774);
nor U644 (N_644,In_1154,In_1520);
nand U645 (N_645,In_2030,In_1508);
or U646 (N_646,In_2856,In_1359);
or U647 (N_647,In_928,In_2253);
xor U648 (N_648,In_948,In_666);
nand U649 (N_649,In_1970,In_2712);
and U650 (N_650,In_2399,In_367);
nor U651 (N_651,In_1665,In_644);
nand U652 (N_652,In_173,In_147);
nor U653 (N_653,In_2074,In_32);
xor U654 (N_654,In_1108,In_1284);
nand U655 (N_655,In_2776,In_1686);
nor U656 (N_656,In_165,In_2034);
nor U657 (N_657,In_1652,In_1192);
nand U658 (N_658,In_1161,In_982);
or U659 (N_659,In_14,In_1351);
or U660 (N_660,In_1277,In_2814);
nand U661 (N_661,In_207,In_2946);
nand U662 (N_662,In_639,In_2522);
or U663 (N_663,In_2882,In_1233);
nand U664 (N_664,In_2799,In_1278);
nor U665 (N_665,In_2093,In_1427);
and U666 (N_666,In_1570,In_2485);
nor U667 (N_667,In_2392,In_1287);
xor U668 (N_668,In_2354,In_2235);
xor U669 (N_669,In_2371,In_2584);
nand U670 (N_670,In_453,In_1450);
and U671 (N_671,In_1594,In_1635);
or U672 (N_672,In_2602,In_1239);
and U673 (N_673,In_2659,In_1079);
or U674 (N_674,In_1236,In_816);
and U675 (N_675,In_1548,In_2756);
nand U676 (N_676,In_1536,In_1);
and U677 (N_677,In_2535,In_2319);
nor U678 (N_678,In_319,In_2167);
nor U679 (N_679,In_1155,In_2760);
or U680 (N_680,In_2531,In_645);
xnor U681 (N_681,In_2538,In_407);
and U682 (N_682,In_998,In_142);
or U683 (N_683,In_1524,In_675);
and U684 (N_684,In_601,In_2907);
nor U685 (N_685,In_1912,In_1724);
nand U686 (N_686,In_91,In_585);
xor U687 (N_687,In_1271,In_2779);
xor U688 (N_688,In_23,In_2445);
and U689 (N_689,In_523,In_2387);
xor U690 (N_690,In_2190,In_1392);
nor U691 (N_691,In_1507,In_598);
and U692 (N_692,In_6,In_795);
and U693 (N_693,In_1460,In_2264);
nor U694 (N_694,In_2656,In_2376);
or U695 (N_695,In_279,In_1962);
nand U696 (N_696,In_1349,In_1646);
nor U697 (N_697,In_58,In_2085);
nor U698 (N_698,In_2643,In_1036);
and U699 (N_699,In_36,In_2327);
and U700 (N_700,In_929,In_2736);
nor U701 (N_701,In_2010,In_1921);
nor U702 (N_702,In_1802,In_797);
xnor U703 (N_703,In_2373,In_2853);
nor U704 (N_704,In_341,In_174);
nand U705 (N_705,In_1500,In_2498);
and U706 (N_706,In_859,In_111);
nor U707 (N_707,In_1113,In_895);
and U708 (N_708,In_50,In_672);
or U709 (N_709,In_2317,In_167);
xor U710 (N_710,In_2314,In_1579);
xor U711 (N_711,In_2214,In_921);
and U712 (N_712,In_2980,In_2216);
nor U713 (N_713,In_2739,In_1679);
and U714 (N_714,In_2690,In_333);
nor U715 (N_715,In_1262,In_1207);
or U716 (N_716,In_1971,In_2971);
nand U717 (N_717,In_2112,In_2432);
nand U718 (N_718,In_1185,In_1801);
xnor U719 (N_719,In_2985,In_1664);
nor U720 (N_720,In_588,In_2477);
or U721 (N_721,In_1751,In_2147);
xor U722 (N_722,In_1172,In_2500);
nand U723 (N_723,In_2612,In_1038);
nand U724 (N_724,In_2622,In_878);
nand U725 (N_725,In_935,In_1030);
nand U726 (N_726,In_505,In_1786);
and U727 (N_727,In_830,In_2624);
or U728 (N_728,In_2234,In_1793);
and U729 (N_729,In_2064,In_2915);
nor U730 (N_730,In_489,In_1398);
xor U731 (N_731,In_423,In_434);
nor U732 (N_732,In_124,In_1354);
xor U733 (N_733,In_1098,In_183);
or U734 (N_734,In_1182,In_2959);
nand U735 (N_735,In_1184,In_449);
xnor U736 (N_736,In_478,In_1732);
xnor U737 (N_737,In_1684,In_2563);
nor U738 (N_738,In_248,In_784);
nor U739 (N_739,In_2377,In_953);
nand U740 (N_740,In_2891,In_1909);
nand U741 (N_741,In_1806,In_913);
or U742 (N_742,In_2156,In_2183);
nand U743 (N_743,In_1272,In_2913);
xor U744 (N_744,In_1634,In_2669);
nand U745 (N_745,In_1804,In_993);
nor U746 (N_746,In_1926,In_1938);
xor U747 (N_747,In_2722,In_2533);
xnor U748 (N_748,In_1357,In_2128);
or U749 (N_749,In_2312,In_2742);
nand U750 (N_750,In_346,In_454);
nand U751 (N_751,In_70,In_149);
nor U752 (N_752,In_811,In_801);
nor U753 (N_753,In_574,In_792);
nand U754 (N_754,In_1348,In_1477);
nand U755 (N_755,In_1836,In_1689);
nand U756 (N_756,In_1947,In_1870);
xor U757 (N_757,In_2320,In_2863);
and U758 (N_758,In_571,In_1175);
and U759 (N_759,In_872,In_1541);
xnor U760 (N_760,In_2499,In_1910);
and U761 (N_761,In_1397,In_2888);
nand U762 (N_762,In_1837,In_1199);
xor U763 (N_763,In_2754,In_2063);
nand U764 (N_764,In_1680,In_1475);
or U765 (N_765,In_2864,In_2358);
nor U766 (N_766,In_377,In_1315);
or U767 (N_767,In_2784,In_1388);
nand U768 (N_768,In_2816,In_561);
nor U769 (N_769,In_2520,In_181);
or U770 (N_770,In_1637,In_1299);
nand U771 (N_771,In_1697,In_503);
or U772 (N_772,In_1683,In_1002);
and U773 (N_773,In_2897,In_2703);
or U774 (N_774,In_1265,In_1729);
and U775 (N_775,In_1605,In_2243);
xnor U776 (N_776,In_2002,In_1863);
and U777 (N_777,In_140,In_1413);
nor U778 (N_778,In_143,In_2255);
or U779 (N_779,In_2873,In_1505);
and U780 (N_780,In_1273,In_2459);
and U781 (N_781,In_1209,In_984);
or U782 (N_782,In_661,In_549);
nor U783 (N_783,In_1587,In_1942);
nand U784 (N_784,In_1826,In_2240);
or U785 (N_785,In_1622,In_1111);
nor U786 (N_786,In_2608,In_1738);
or U787 (N_787,In_1857,In_1402);
nor U788 (N_788,In_2514,In_1197);
nor U789 (N_789,In_2364,In_2835);
or U790 (N_790,In_961,In_2125);
nor U791 (N_791,In_1437,In_241);
nor U792 (N_792,In_1049,In_2348);
nor U793 (N_793,In_1471,In_2661);
or U794 (N_794,In_2068,In_2343);
nor U795 (N_795,In_1558,In_2375);
nor U796 (N_796,In_1381,In_1838);
and U797 (N_797,In_1825,In_71);
or U798 (N_798,In_1913,In_2800);
nor U799 (N_799,In_2721,In_2062);
nand U800 (N_800,In_1586,In_308);
nand U801 (N_801,In_2557,In_2625);
and U802 (N_802,In_122,In_1618);
or U803 (N_803,In_1484,In_949);
nand U804 (N_804,In_49,In_2526);
or U805 (N_805,In_582,In_1292);
and U806 (N_806,In_630,In_539);
xnor U807 (N_807,In_1395,In_2464);
or U808 (N_808,In_1530,In_619);
nand U809 (N_809,In_1747,In_2579);
nor U810 (N_810,In_2751,In_803);
and U811 (N_811,In_1880,In_2586);
xor U812 (N_812,In_1430,In_356);
nand U813 (N_813,In_1117,In_897);
nor U814 (N_814,In_1948,In_1296);
or U815 (N_815,In_231,In_2995);
nor U816 (N_816,In_2745,In_2350);
and U817 (N_817,In_1861,In_2846);
xnor U818 (N_818,In_451,In_506);
nand U819 (N_819,In_2875,In_977);
nor U820 (N_820,In_654,In_657);
nor U821 (N_821,In_2765,In_828);
or U822 (N_822,In_1757,In_256);
nand U823 (N_823,In_338,In_2226);
nand U824 (N_824,In_1561,In_1092);
and U825 (N_825,In_2148,In_1733);
xor U826 (N_826,In_2999,In_980);
or U827 (N_827,In_92,In_310);
or U828 (N_828,In_634,In_553);
nor U829 (N_829,In_1756,In_204);
xor U830 (N_830,In_125,In_786);
nor U831 (N_831,In_2242,In_391);
nor U832 (N_832,In_2246,In_28);
and U833 (N_833,In_2378,In_2788);
nand U834 (N_834,In_2155,In_2806);
or U835 (N_835,In_2859,In_94);
xor U836 (N_836,In_1422,In_1867);
and U837 (N_837,In_1008,In_205);
nand U838 (N_838,In_1372,In_1066);
nand U839 (N_839,In_1071,In_603);
xnor U840 (N_840,In_161,In_2673);
and U841 (N_841,In_1258,In_2173);
nor U842 (N_842,In_2150,In_110);
nand U843 (N_843,In_2091,In_2395);
nor U844 (N_844,In_7,In_2044);
xor U845 (N_845,In_2496,In_1796);
nand U846 (N_846,In_2457,In_898);
nand U847 (N_847,In_1666,In_1625);
xnor U848 (N_848,In_2379,In_605);
or U849 (N_849,In_215,In_1486);
and U850 (N_850,In_2437,In_1183);
xor U851 (N_851,In_107,In_528);
nand U852 (N_852,In_1433,In_791);
xnor U853 (N_853,In_1927,In_1784);
xor U854 (N_854,In_511,In_1840);
nand U855 (N_855,In_2139,In_2758);
nand U856 (N_856,In_3,In_1485);
nand U857 (N_857,In_2517,In_1623);
nor U858 (N_858,In_1163,In_1873);
xnor U859 (N_859,In_1718,In_2746);
nor U860 (N_860,In_2993,In_2290);
and U861 (N_861,In_1118,In_2990);
xnor U862 (N_862,In_345,In_1307);
nor U863 (N_863,In_254,In_593);
xor U864 (N_864,In_2228,In_550);
nand U865 (N_865,In_1954,In_960);
xor U866 (N_866,In_2497,In_392);
and U867 (N_867,In_1345,In_190);
and U868 (N_868,In_2165,In_836);
nor U869 (N_869,In_2542,In_728);
xor U870 (N_870,In_2079,In_939);
nor U871 (N_871,In_2879,In_1983);
nand U872 (N_872,In_773,In_2609);
nor U873 (N_873,In_481,In_2408);
or U874 (N_874,In_2926,In_1787);
and U875 (N_875,In_2185,In_2809);
nor U876 (N_876,In_1820,In_1572);
xor U877 (N_877,In_21,In_2640);
and U878 (N_878,In_2086,In_1019);
and U879 (N_879,In_730,In_8);
xor U880 (N_880,In_1759,In_465);
or U881 (N_881,In_93,In_1053);
nand U882 (N_882,In_1911,In_1675);
and U883 (N_883,In_2014,In_2184);
xor U884 (N_884,In_1741,In_239);
and U885 (N_885,In_1468,In_2295);
nor U886 (N_886,In_472,In_2372);
and U887 (N_887,In_1116,In_307);
or U888 (N_888,In_2764,In_2670);
xor U889 (N_889,In_809,In_2495);
or U890 (N_890,In_979,In_1454);
nand U891 (N_891,In_1790,In_240);
or U892 (N_892,In_1920,In_2973);
nor U893 (N_893,In_2130,In_2250);
nor U894 (N_894,In_2678,In_2509);
and U895 (N_895,In_2302,In_664);
nand U896 (N_896,In_2293,In_31);
xnor U897 (N_897,In_162,In_616);
nor U898 (N_898,In_1953,In_1342);
xnor U899 (N_899,In_2537,In_1638);
nand U900 (N_900,In_43,In_300);
and U901 (N_901,In_2425,In_1343);
nand U902 (N_902,In_950,In_1653);
or U903 (N_903,In_1775,In_2606);
xor U904 (N_904,In_2527,In_245);
xor U905 (N_905,In_2738,In_2204);
nand U906 (N_906,In_2925,In_223);
nand U907 (N_907,In_711,In_1540);
nand U908 (N_908,In_2357,In_2426);
nand U909 (N_909,In_1874,In_343);
or U910 (N_910,In_2617,In_926);
xnor U911 (N_911,In_1663,In_447);
nor U912 (N_912,In_1742,In_1028);
nand U913 (N_913,In_2977,In_227);
nor U914 (N_914,In_397,In_2092);
and U915 (N_915,In_1821,In_2989);
or U916 (N_916,In_1220,In_108);
or U917 (N_917,In_557,In_2198);
and U918 (N_918,In_2552,In_1671);
nor U919 (N_919,In_744,In_587);
xor U920 (N_920,In_2631,In_1841);
xor U921 (N_921,In_2345,In_166);
nor U922 (N_922,In_1489,In_1474);
or U923 (N_923,In_385,In_747);
and U924 (N_924,In_1752,In_2342);
or U925 (N_925,In_1242,In_2919);
and U926 (N_926,In_880,In_1763);
nand U927 (N_927,In_1162,In_1488);
xor U928 (N_928,In_1555,In_847);
nand U929 (N_929,In_2540,In_470);
or U930 (N_930,In_1238,In_1930);
xnor U931 (N_931,In_1459,In_2544);
or U932 (N_932,In_1627,In_934);
xor U933 (N_933,In_1719,In_387);
and U934 (N_934,In_2431,In_444);
and U935 (N_935,In_4,In_900);
or U936 (N_936,In_2773,In_2427);
or U937 (N_937,In_2969,In_2080);
and U938 (N_938,In_2725,In_1061);
nor U939 (N_939,In_2045,In_1216);
and U940 (N_940,In_2158,In_235);
nand U941 (N_941,In_1291,In_1361);
nand U942 (N_942,In_1580,In_2224);
nor U943 (N_943,In_187,In_1076);
nand U944 (N_944,In_210,In_1400);
or U945 (N_945,In_2605,In_1685);
xnor U946 (N_946,In_2731,In_1760);
nor U947 (N_947,In_1149,In_2714);
nor U948 (N_948,In_2752,In_1103);
nand U949 (N_949,In_179,In_665);
nor U950 (N_950,In_1029,In_2292);
and U951 (N_951,In_848,In_738);
nor U952 (N_952,In_990,In_1497);
nand U953 (N_953,In_2588,In_837);
nor U954 (N_954,In_1931,In_1592);
or U955 (N_955,In_1834,In_936);
or U956 (N_956,In_29,In_313);
nor U957 (N_957,In_736,In_1977);
or U958 (N_958,In_1967,In_825);
and U959 (N_959,In_1566,In_688);
and U960 (N_960,In_594,In_1204);
or U961 (N_961,In_2630,In_304);
nor U962 (N_962,In_1659,In_1025);
xnor U963 (N_963,In_1153,In_1891);
nand U964 (N_964,In_253,In_2041);
nand U965 (N_965,In_1768,In_781);
and U966 (N_966,In_419,In_1129);
and U967 (N_967,In_1046,In_2059);
nand U968 (N_968,In_2244,In_756);
nand U969 (N_969,In_818,In_2851);
nand U970 (N_970,In_1196,In_176);
nand U971 (N_971,In_538,In_1000);
nor U972 (N_972,In_2808,In_1045);
xor U973 (N_973,In_726,In_2207);
nand U974 (N_974,In_706,In_1368);
nor U975 (N_975,In_326,In_212);
xnor U976 (N_976,In_2802,In_1792);
nor U977 (N_977,In_1879,In_1379);
xnor U978 (N_978,In_2434,In_2033);
or U979 (N_979,In_2709,In_2771);
nor U980 (N_980,In_1762,In_359);
nor U981 (N_981,In_793,In_655);
nand U982 (N_982,In_2750,In_2700);
or U983 (N_983,In_580,In_614);
nor U984 (N_984,In_1626,In_2291);
or U985 (N_985,In_2398,In_1270);
or U986 (N_986,In_1808,In_1542);
nor U987 (N_987,In_2582,In_59);
nor U988 (N_988,In_2692,In_2278);
or U989 (N_989,In_2382,In_219);
xor U990 (N_990,In_1833,In_2782);
or U991 (N_991,In_1750,In_1791);
xor U992 (N_992,In_1516,In_33);
or U993 (N_993,In_1487,In_1482);
or U994 (N_994,In_964,In_1904);
nand U995 (N_995,In_1657,In_1544);
or U996 (N_996,In_400,In_224);
and U997 (N_997,In_320,In_2822);
or U998 (N_998,In_2911,In_1063);
or U999 (N_999,In_316,In_76);
or U1000 (N_1000,In_2415,In_2895);
and U1001 (N_1001,In_2696,In_2220);
nor U1002 (N_1002,In_2238,In_2559);
nor U1003 (N_1003,In_2416,In_252);
nor U1004 (N_1004,In_2116,In_390);
xnor U1005 (N_1005,In_1581,In_2488);
xnor U1006 (N_1006,In_2636,In_20);
nand U1007 (N_1007,In_2834,In_1423);
and U1008 (N_1008,In_772,In_1219);
xor U1009 (N_1009,In_2501,In_1951);
nand U1010 (N_1010,In_1585,In_2421);
nand U1011 (N_1011,In_388,In_653);
xor U1012 (N_1012,In_2095,In_2593);
or U1013 (N_1013,In_325,In_1100);
nor U1014 (N_1014,In_2104,In_2380);
and U1015 (N_1015,In_1157,In_340);
and U1016 (N_1016,In_2695,In_1513);
and U1017 (N_1017,In_128,In_2473);
and U1018 (N_1018,In_442,In_1431);
or U1019 (N_1019,In_2031,In_1027);
nor U1020 (N_1020,In_46,In_379);
xor U1021 (N_1021,In_1526,In_908);
and U1022 (N_1022,In_1803,In_1554);
xnor U1023 (N_1023,In_1138,In_2199);
nand U1024 (N_1024,In_2825,In_1373);
nor U1025 (N_1025,In_805,In_1255);
nand U1026 (N_1026,In_2005,In_1037);
nor U1027 (N_1027,In_884,In_2635);
or U1028 (N_1028,In_1734,In_2694);
nand U1029 (N_1029,In_1928,In_1083);
and U1030 (N_1030,In_79,In_2974);
xor U1031 (N_1031,In_2326,In_852);
nor U1032 (N_1032,In_2049,In_1559);
nand U1033 (N_1033,In_1799,In_2001);
and U1034 (N_1034,In_2983,In_1144);
or U1035 (N_1035,In_501,In_2337);
or U1036 (N_1036,In_1268,In_2534);
xnor U1037 (N_1037,In_335,In_2762);
xnor U1038 (N_1038,In_1856,In_1758);
nor U1039 (N_1039,In_822,In_232);
nand U1040 (N_1040,In_2682,In_530);
xnor U1041 (N_1041,In_1112,In_1633);
or U1042 (N_1042,In_2298,In_824);
and U1043 (N_1043,In_1855,In_696);
and U1044 (N_1044,In_118,In_45);
nand U1045 (N_1045,In_370,In_1150);
xor U1046 (N_1046,In_2076,In_431);
or U1047 (N_1047,In_2860,In_2564);
or U1048 (N_1048,In_510,In_509);
nand U1049 (N_1049,In_1944,In_1179);
nand U1050 (N_1050,In_945,In_428);
and U1051 (N_1051,In_113,In_184);
or U1052 (N_1052,In_1493,In_1367);
nor U1053 (N_1053,In_613,In_297);
nand U1054 (N_1054,In_543,In_1610);
xor U1055 (N_1055,In_1814,In_2838);
xnor U1056 (N_1056,In_2516,In_1429);
or U1057 (N_1057,In_2841,In_1822);
nand U1058 (N_1058,In_2909,In_2209);
or U1059 (N_1059,In_1124,In_860);
nor U1060 (N_1060,In_1068,In_1465);
xnor U1061 (N_1061,In_2444,In_1457);
nor U1062 (N_1062,In_1815,In_135);
xnor U1063 (N_1063,In_363,In_42);
and U1064 (N_1064,In_647,In_1304);
and U1065 (N_1065,In_1311,In_2324);
and U1066 (N_1066,In_351,In_369);
or U1067 (N_1067,In_2070,In_1805);
nor U1068 (N_1068,In_827,In_41);
nor U1069 (N_1069,In_2597,In_2460);
and U1070 (N_1070,In_373,In_1456);
nand U1071 (N_1071,In_5,In_534);
nand U1072 (N_1072,In_972,In_1201);
nor U1073 (N_1073,In_992,In_1887);
or U1074 (N_1074,In_2219,In_1158);
and U1075 (N_1075,In_2462,In_1549);
nand U1076 (N_1076,In_2975,In_1039);
and U1077 (N_1077,In_2575,In_576);
or U1078 (N_1078,In_2296,In_153);
or U1079 (N_1079,In_2200,In_2840);
and U1080 (N_1080,In_1440,In_2383);
or U1081 (N_1081,In_2098,In_612);
nand U1082 (N_1082,In_2465,In_2972);
nor U1083 (N_1083,In_2164,In_807);
or U1084 (N_1084,In_1503,In_2968);
xor U1085 (N_1085,In_2964,In_1923);
nor U1086 (N_1086,In_788,In_1001);
xnor U1087 (N_1087,In_1852,In_2335);
and U1088 (N_1088,In_2607,In_1517);
and U1089 (N_1089,In_2131,In_1699);
nor U1090 (N_1090,In_1945,In_646);
and U1091 (N_1091,In_515,In_1644);
nand U1092 (N_1092,In_1330,In_1993);
xnor U1093 (N_1093,In_1906,In_236);
xnor U1094 (N_1094,In_2982,In_2938);
nor U1095 (N_1095,In_2978,In_2574);
nor U1096 (N_1096,In_866,In_327);
and U1097 (N_1097,In_1226,In_2307);
nand U1098 (N_1098,In_1052,In_1131);
or U1099 (N_1099,In_2766,In_1597);
or U1100 (N_1100,In_1518,In_1892);
xnor U1101 (N_1101,In_52,In_2699);
and U1102 (N_1102,In_2942,In_2233);
and U1103 (N_1103,In_2146,In_724);
xnor U1104 (N_1104,In_720,In_1968);
or U1105 (N_1105,In_2197,In_2057);
and U1106 (N_1106,In_2149,In_1470);
nand U1107 (N_1107,In_2266,In_198);
and U1108 (N_1108,In_1140,In_500);
xor U1109 (N_1109,In_2402,In_1886);
and U1110 (N_1110,In_1356,In_620);
and U1111 (N_1111,In_2600,In_2019);
and U1112 (N_1112,In_1331,In_458);
and U1113 (N_1113,In_1506,In_2963);
nand U1114 (N_1114,In_312,In_578);
and U1115 (N_1115,In_418,In_1936);
and U1116 (N_1116,In_2652,In_2211);
and U1117 (N_1117,In_2737,In_682);
xnor U1118 (N_1118,In_2940,In_1491);
or U1119 (N_1119,In_103,In_1444);
xor U1120 (N_1120,In_1463,In_177);
or U1121 (N_1121,In_673,In_203);
and U1122 (N_1122,In_677,In_1434);
or U1123 (N_1123,In_2877,In_581);
or U1124 (N_1124,In_1441,In_427);
xor U1125 (N_1125,In_2697,In_577);
xor U1126 (N_1126,In_547,In_1709);
nand U1127 (N_1127,In_1492,In_488);
or U1128 (N_1128,In_586,In_2082);
nor U1129 (N_1129,In_466,In_2351);
nor U1130 (N_1130,In_13,In_592);
or U1131 (N_1131,In_294,In_814);
nor U1132 (N_1132,In_715,In_563);
nor U1133 (N_1133,In_450,In_641);
or U1134 (N_1134,In_2015,In_1346);
or U1135 (N_1135,In_1777,In_826);
nor U1136 (N_1136,In_2555,In_2050);
nor U1137 (N_1137,In_2658,In_739);
nor U1138 (N_1138,In_2780,In_2719);
or U1139 (N_1139,In_2910,In_1316);
or U1140 (N_1140,In_2018,In_2012);
xor U1141 (N_1141,In_1860,In_353);
and U1142 (N_1142,In_1435,In_2823);
xnor U1143 (N_1143,In_1288,In_1878);
nand U1144 (N_1144,In_2894,In_1514);
nor U1145 (N_1145,In_962,In_1510);
nand U1146 (N_1146,In_2455,In_405);
nor U1147 (N_1147,In_1461,In_2626);
nand U1148 (N_1148,In_1690,In_437);
or U1149 (N_1149,In_1641,In_2683);
or U1150 (N_1150,In_684,In_1900);
xor U1151 (N_1151,In_1916,In_911);
or U1152 (N_1152,In_2629,In_396);
or U1153 (N_1153,In_1225,In_732);
xor U1154 (N_1154,In_2043,In_2667);
nand U1155 (N_1155,In_1415,In_1617);
or U1156 (N_1156,In_2715,In_2627);
xor U1157 (N_1157,In_222,In_622);
xnor U1158 (N_1158,In_329,In_2687);
nor U1159 (N_1159,In_1976,In_1215);
xor U1160 (N_1160,In_134,In_891);
xor U1161 (N_1161,In_1293,In_1104);
xor U1162 (N_1162,In_2734,In_411);
or U1163 (N_1163,In_2848,In_579);
xor U1164 (N_1164,In_200,In_2000);
nand U1165 (N_1165,In_2301,In_946);
or U1166 (N_1166,In_1428,In_2138);
nor U1167 (N_1167,In_2048,In_2912);
or U1168 (N_1168,In_876,In_415);
or U1169 (N_1169,In_1591,In_1134);
nor U1170 (N_1170,In_1203,In_1003);
nand U1171 (N_1171,In_1152,In_1525);
or U1172 (N_1172,In_1306,In_154);
or U1173 (N_1173,In_1546,In_904);
or U1174 (N_1174,In_2451,In_498);
nand U1175 (N_1175,In_1347,In_1877);
nor U1176 (N_1176,In_1360,In_745);
xnor U1177 (N_1177,In_2646,In_1589);
nor U1178 (N_1178,In_2987,In_109);
nor U1179 (N_1179,In_1371,In_2741);
xor U1180 (N_1180,In_1128,In_737);
xnor U1181 (N_1181,In_753,In_467);
and U1182 (N_1182,In_2706,In_19);
xor U1183 (N_1183,In_2928,In_1198);
or U1184 (N_1184,In_2939,In_249);
xnor U1185 (N_1185,In_702,In_456);
and U1186 (N_1186,In_2665,In_1883);
xnor U1187 (N_1187,In_459,In_482);
nand U1188 (N_1188,In_640,In_261);
and U1189 (N_1189,In_1317,In_2159);
or U1190 (N_1190,In_833,In_1147);
and U1191 (N_1191,In_776,In_2028);
xnor U1192 (N_1192,In_2121,In_1101);
nor U1193 (N_1193,In_874,In_2847);
or U1194 (N_1194,In_2587,In_1590);
xor U1195 (N_1195,In_1893,In_39);
xnor U1196 (N_1196,In_2232,In_1846);
and U1197 (N_1197,In_1021,In_1091);
or U1198 (N_1198,In_768,In_318);
and U1199 (N_1199,In_923,In_636);
and U1200 (N_1200,In_1051,In_537);
nand U1201 (N_1201,In_2992,In_1529);
xor U1202 (N_1202,In_2642,In_2446);
nor U1203 (N_1203,In_1243,In_527);
xnor U1204 (N_1204,In_703,In_750);
and U1205 (N_1205,In_2639,In_541);
nand U1206 (N_1206,In_2420,In_2723);
nor U1207 (N_1207,In_591,In_1044);
nor U1208 (N_1208,In_102,In_1606);
xnor U1209 (N_1209,In_2867,In_804);
and U1210 (N_1210,In_658,In_2140);
nand U1211 (N_1211,In_286,In_839);
xor U1212 (N_1212,In_971,In_952);
xnor U1213 (N_1213,In_1180,In_595);
nand U1214 (N_1214,In_829,In_524);
or U1215 (N_1215,In_15,In_631);
and U1216 (N_1216,In_2870,In_1472);
xnor U1217 (N_1217,In_2660,In_1339);
nor U1218 (N_1218,In_1918,In_2309);
or U1219 (N_1219,In_1419,In_2815);
nand U1220 (N_1220,In_1385,In_2359);
xnor U1221 (N_1221,In_1726,In_1515);
and U1222 (N_1222,In_2729,In_1077);
and U1223 (N_1223,In_2674,In_1439);
and U1224 (N_1224,In_2874,In_305);
nor U1225 (N_1225,In_2558,In_1973);
or U1226 (N_1226,In_893,In_1778);
and U1227 (N_1227,In_315,In_2078);
nand U1228 (N_1228,In_265,In_906);
nor U1229 (N_1229,In_1557,In_342);
and U1230 (N_1230,In_2212,In_51);
nor U1231 (N_1231,In_2248,In_2311);
nand U1232 (N_1232,In_2718,In_690);
or U1233 (N_1233,In_1829,In_2565);
and U1234 (N_1234,In_2272,In_1981);
or U1235 (N_1235,In_1380,In_611);
xor U1236 (N_1236,In_114,In_399);
and U1237 (N_1237,In_1810,In_714);
xor U1238 (N_1238,In_1783,In_1334);
and U1239 (N_1239,In_2937,In_332);
xor U1240 (N_1240,In_2285,In_1223);
xnor U1241 (N_1241,In_867,In_269);
nand U1242 (N_1242,In_2518,In_468);
or U1243 (N_1243,In_2591,In_2644);
nand U1244 (N_1244,In_2021,In_1980);
and U1245 (N_1245,In_2467,In_2610);
nor U1246 (N_1246,In_2480,In_2286);
and U1247 (N_1247,In_169,In_1582);
or U1248 (N_1248,In_2899,In_186);
nand U1249 (N_1249,In_2852,In_965);
nor U1250 (N_1250,In_1688,In_2775);
nor U1251 (N_1251,In_1399,In_2061);
nand U1252 (N_1252,In_350,In_2103);
nand U1253 (N_1253,In_659,In_126);
or U1254 (N_1254,In_1214,In_1452);
nor U1255 (N_1255,In_1298,In_1745);
xor U1256 (N_1256,In_930,In_2855);
nand U1257 (N_1257,In_2727,In_2490);
and U1258 (N_1258,In_1240,In_80);
xor U1259 (N_1259,In_938,In_1827);
nand U1260 (N_1260,In_2206,In_632);
xor U1261 (N_1261,In_864,In_44);
or U1262 (N_1262,In_885,In_1889);
and U1263 (N_1263,In_931,In_1257);
or U1264 (N_1264,In_2795,In_1283);
nor U1265 (N_1265,In_1363,In_2811);
nor U1266 (N_1266,In_2781,In_999);
nand U1267 (N_1267,In_1065,In_9);
xnor U1268 (N_1268,In_1285,In_914);
or U1269 (N_1269,In_2541,In_2844);
or U1270 (N_1270,In_2265,In_1406);
xnor U1271 (N_1271,In_2638,In_2649);
and U1272 (N_1272,In_717,In_2476);
xnor U1273 (N_1273,In_1067,In_292);
nor U1274 (N_1274,In_2958,In_2182);
xnor U1275 (N_1275,In_2885,In_2733);
and U1276 (N_1276,In_2986,In_518);
or U1277 (N_1277,In_2890,In_2920);
and U1278 (N_1278,In_1442,In_691);
xnor U1279 (N_1279,In_2805,In_2872);
nor U1280 (N_1280,In_69,In_2016);
and U1281 (N_1281,In_544,In_1280);
nand U1282 (N_1282,In_905,In_484);
or U1283 (N_1283,In_2194,In_1321);
or U1284 (N_1284,In_1882,In_1173);
and U1285 (N_1285,In_1770,In_1340);
or U1286 (N_1286,In_943,In_1074);
xnor U1287 (N_1287,In_1940,In_96);
nor U1288 (N_1288,In_985,In_2067);
xor U1289 (N_1289,In_573,In_1609);
nor U1290 (N_1290,In_1058,In_951);
or U1291 (N_1291,In_901,In_932);
nand U1292 (N_1292,In_525,In_2757);
or U1293 (N_1293,In_2494,In_146);
and U1294 (N_1294,In_445,In_2505);
nor U1295 (N_1295,In_2573,In_1337);
or U1296 (N_1296,In_1410,In_1136);
nor U1297 (N_1297,In_18,In_841);
or U1298 (N_1298,In_54,In_1929);
or U1299 (N_1299,In_191,In_2581);
and U1300 (N_1300,In_1998,In_2903);
and U1301 (N_1301,In_994,In_705);
and U1302 (N_1302,In_1600,In_1631);
and U1303 (N_1303,In_758,In_77);
or U1304 (N_1304,In_894,In_1865);
nand U1305 (N_1305,In_770,In_448);
nand U1306 (N_1306,In_1781,In_2892);
xnor U1307 (N_1307,In_424,In_2249);
nand U1308 (N_1308,In_2688,In_2458);
nand U1309 (N_1309,In_1812,In_2956);
nand U1310 (N_1310,In_2837,In_735);
or U1311 (N_1311,In_1139,In_2743);
nor U1312 (N_1312,In_1070,In_2869);
nand U1313 (N_1313,In_2529,In_719);
and U1314 (N_1314,In_1187,In_1766);
nand U1315 (N_1315,In_2360,In_896);
xor U1316 (N_1316,In_2166,In_521);
or U1317 (N_1317,In_976,In_2701);
nor U1318 (N_1318,In_2921,In_1984);
or U1319 (N_1319,In_381,In_2772);
nor U1320 (N_1320,In_2418,In_2539);
nor U1321 (N_1321,In_997,In_220);
nor U1322 (N_1322,In_119,In_65);
or U1323 (N_1323,In_1048,In_1917);
xnor U1324 (N_1324,In_1744,In_1847);
nand U1325 (N_1325,In_2566,In_1550);
xnor U1326 (N_1326,In_1085,In_2819);
or U1327 (N_1327,In_1411,In_2117);
xnor U1328 (N_1328,In_1632,In_401);
nor U1329 (N_1329,In_572,In_1012);
and U1330 (N_1330,In_298,In_2276);
and U1331 (N_1331,In_2858,In_2297);
nor U1332 (N_1332,In_1274,In_2793);
nand U1333 (N_1333,In_1481,In_2254);
xnor U1334 (N_1334,In_559,In_731);
nand U1335 (N_1335,In_1107,In_495);
xor U1336 (N_1336,In_1082,In_1539);
nand U1337 (N_1337,In_476,In_2484);
nor U1338 (N_1338,In_2325,In_1473);
and U1339 (N_1339,In_2417,In_1056);
xor U1340 (N_1340,In_2512,In_2818);
nor U1341 (N_1341,In_2251,In_618);
xnor U1342 (N_1342,In_443,In_365);
or U1343 (N_1343,In_2252,In_752);
nand U1344 (N_1344,In_1924,In_963);
and U1345 (N_1345,In_2730,In_708);
xnor U1346 (N_1346,In_1935,In_2583);
nor U1347 (N_1347,In_2161,In_2330);
xor U1348 (N_1348,In_255,In_2483);
and U1349 (N_1349,In_267,In_1261);
nand U1350 (N_1350,In_663,In_2132);
nand U1351 (N_1351,In_1015,In_348);
nor U1352 (N_1352,In_78,In_2794);
and U1353 (N_1353,In_2468,In_336);
or U1354 (N_1354,In_1387,In_1445);
and U1355 (N_1355,In_2560,In_1211);
nor U1356 (N_1356,In_1996,In_372);
and U1357 (N_1357,In_213,In_2456);
nand U1358 (N_1358,In_2753,In_701);
nand U1359 (N_1359,In_1925,In_2530);
nor U1360 (N_1360,In_727,In_233);
nor U1361 (N_1361,In_850,In_2994);
xor U1362 (N_1362,In_1614,In_440);
nand U1363 (N_1363,In_540,In_276);
nand U1364 (N_1364,In_1681,In_2615);
or U1365 (N_1365,In_115,In_545);
nor U1366 (N_1366,In_1466,In_755);
or U1367 (N_1367,In_180,In_1159);
or U1368 (N_1368,In_1408,In_2528);
or U1369 (N_1369,In_2839,In_1414);
nor U1370 (N_1370,In_1575,In_1937);
nor U1371 (N_1371,In_1190,In_2689);
nor U1372 (N_1372,In_1884,In_463);
nand U1373 (N_1373,In_194,In_2178);
and U1374 (N_1374,In_637,In_197);
xor U1375 (N_1375,In_2133,In_1495);
or U1376 (N_1376,In_1616,In_2299);
nor U1377 (N_1377,In_1914,In_417);
or U1378 (N_1378,In_384,In_2308);
or U1379 (N_1379,In_2519,In_257);
nand U1380 (N_1380,In_492,In_1386);
or U1381 (N_1381,In_1601,In_927);
nand U1382 (N_1382,In_130,In_250);
and U1383 (N_1383,In_2230,In_1604);
nor U1384 (N_1384,In_2047,In_1963);
and U1385 (N_1385,In_2862,In_2933);
nor U1386 (N_1386,In_2260,In_2281);
nand U1387 (N_1387,In_1583,In_2929);
or U1388 (N_1388,In_2482,In_2270);
or U1389 (N_1389,In_2829,In_2006);
nand U1390 (N_1390,In_116,In_2361);
xnor U1391 (N_1391,In_1443,In_627);
or U1392 (N_1392,In_1333,In_284);
xor U1393 (N_1393,In_958,In_2262);
xnor U1394 (N_1394,In_2218,In_2596);
nor U1395 (N_1395,In_2025,In_2193);
nor U1396 (N_1396,In_1377,In_2896);
and U1397 (N_1397,In_477,In_1084);
nand U1398 (N_1398,In_689,In_1682);
nor U1399 (N_1399,In_494,In_2798);
xnor U1400 (N_1400,In_787,In_2826);
or U1401 (N_1401,In_989,In_924);
and U1402 (N_1402,In_303,In_2115);
or U1403 (N_1403,In_486,In_1476);
nor U1404 (N_1404,In_1862,In_1114);
or U1405 (N_1405,In_2569,In_62);
or U1406 (N_1406,In_383,In_910);
and U1407 (N_1407,In_2961,In_296);
xnor U1408 (N_1408,In_395,In_698);
nor U1409 (N_1409,In_2553,In_1177);
nand U1410 (N_1410,In_97,In_2225);
and U1411 (N_1411,In_1654,In_2747);
or U1412 (N_1412,In_1096,In_1660);
nor U1413 (N_1413,In_2409,In_2441);
nor U1414 (N_1414,In_2137,In_968);
or U1415 (N_1415,In_2390,In_2071);
and U1416 (N_1416,In_299,In_1072);
nand U1417 (N_1417,In_2181,In_1717);
and U1418 (N_1418,In_883,In_1636);
and U1419 (N_1419,In_933,In_27);
or U1420 (N_1420,In_2400,In_2685);
and U1421 (N_1421,In_1119,In_529);
nor U1422 (N_1422,In_1166,In_2332);
or U1423 (N_1423,In_1090,In_1375);
nor U1424 (N_1424,In_947,In_1120);
nand U1425 (N_1425,In_1868,In_2118);
and U1426 (N_1426,In_1013,In_1099);
xnor U1427 (N_1427,In_446,In_1329);
xor U1428 (N_1428,In_2440,In_1669);
nor U1429 (N_1429,In_2623,In_435);
xnor U1430 (N_1430,In_1871,In_2406);
or U1431 (N_1431,In_1761,In_1705);
nand U1432 (N_1432,In_531,In_823);
nor U1433 (N_1433,In_2960,In_1694);
xnor U1434 (N_1434,In_1797,In_716);
or U1435 (N_1435,In_2479,In_394);
or U1436 (N_1436,In_2832,In_2205);
nand U1437 (N_1437,In_293,In_160);
nor U1438 (N_1438,In_1230,In_430);
nor U1439 (N_1439,In_1776,In_389);
or U1440 (N_1440,In_289,In_1054);
nand U1441 (N_1441,In_1412,In_2576);
and U1442 (N_1442,In_2144,In_812);
xnor U1443 (N_1443,In_1109,In_334);
and U1444 (N_1444,In_713,In_2032);
xnor U1445 (N_1445,In_956,In_2404);
and U1446 (N_1446,In_796,In_1142);
nand U1447 (N_1447,In_532,In_1322);
nand U1448 (N_1448,In_2386,In_48);
and U1449 (N_1449,In_2997,In_1982);
xnor U1450 (N_1450,In_287,In_1824);
or U1451 (N_1451,In_625,In_535);
or U1452 (N_1452,In_100,In_863);
nand U1453 (N_1453,In_1715,In_260);
or U1454 (N_1454,In_1767,In_1896);
nor U1455 (N_1455,In_570,In_56);
or U1456 (N_1456,In_266,In_1055);
and U1457 (N_1457,In_406,In_707);
or U1458 (N_1458,In_462,In_1599);
and U1459 (N_1459,In_1047,In_785);
nor U1460 (N_1460,In_969,In_2162);
nor U1461 (N_1461,In_2310,In_131);
xor U1462 (N_1462,In_1958,In_1881);
and U1463 (N_1463,In_275,In_2268);
and U1464 (N_1464,In_2160,In_2672);
nor U1465 (N_1465,In_1328,In_2450);
nor U1466 (N_1466,In_2318,In_899);
and U1467 (N_1467,In_2363,In_2662);
and U1468 (N_1468,In_1712,In_403);
nor U1469 (N_1469,In_1205,In_2259);
or U1470 (N_1470,In_1999,In_2570);
nand U1471 (N_1471,In_555,In_1252);
and U1472 (N_1472,In_217,In_1080);
or U1473 (N_1473,In_375,In_845);
and U1474 (N_1474,In_722,In_810);
or U1475 (N_1475,In_1366,In_2195);
xnor U1476 (N_1476,In_1266,In_202);
or U1477 (N_1477,In_1448,In_2283);
and U1478 (N_1478,In_2504,In_2113);
nand U1479 (N_1479,In_1620,In_2423);
or U1480 (N_1480,In_2424,In_2275);
xnor U1481 (N_1481,In_1978,In_2090);
nor U1482 (N_1482,In_290,In_749);
and U1483 (N_1483,In_2550,In_551);
nor U1484 (N_1484,In_623,In_2273);
and U1485 (N_1485,In_314,In_633);
nor U1486 (N_1486,In_2744,In_2022);
xnor U1487 (N_1487,In_1965,In_2277);
and U1488 (N_1488,In_838,In_1772);
and U1489 (N_1489,In_2066,In_2323);
nand U1490 (N_1490,In_628,In_2329);
and U1491 (N_1491,In_474,In_432);
or U1492 (N_1492,In_1458,In_105);
and U1493 (N_1493,In_957,In_1290);
nand U1494 (N_1494,In_1396,In_1598);
and U1495 (N_1495,In_2981,In_1735);
xor U1496 (N_1496,In_2433,In_86);
and U1497 (N_1497,In_1248,In_1194);
or U1498 (N_1498,In_1727,In_2585);
nand U1499 (N_1499,In_769,In_526);
and U1500 (N_1500,In_867,In_144);
and U1501 (N_1501,In_2471,In_434);
nand U1502 (N_1502,In_2137,In_2891);
and U1503 (N_1503,In_794,In_800);
and U1504 (N_1504,In_2142,In_272);
and U1505 (N_1505,In_2234,In_952);
nand U1506 (N_1506,In_2815,In_2391);
or U1507 (N_1507,In_26,In_231);
or U1508 (N_1508,In_479,In_2163);
and U1509 (N_1509,In_1837,In_686);
and U1510 (N_1510,In_2026,In_771);
and U1511 (N_1511,In_2549,In_1106);
or U1512 (N_1512,In_403,In_729);
nand U1513 (N_1513,In_562,In_1391);
nand U1514 (N_1514,In_166,In_324);
or U1515 (N_1515,In_187,In_2813);
xnor U1516 (N_1516,In_1494,In_2830);
xnor U1517 (N_1517,In_1482,In_501);
nor U1518 (N_1518,In_1649,In_1822);
and U1519 (N_1519,In_515,In_590);
and U1520 (N_1520,In_2924,In_2335);
and U1521 (N_1521,In_565,In_1530);
or U1522 (N_1522,In_1837,In_855);
xor U1523 (N_1523,In_104,In_96);
and U1524 (N_1524,In_736,In_1348);
nand U1525 (N_1525,In_573,In_834);
nor U1526 (N_1526,In_1537,In_1809);
xor U1527 (N_1527,In_2213,In_1273);
nand U1528 (N_1528,In_621,In_2660);
nand U1529 (N_1529,In_58,In_2884);
nand U1530 (N_1530,In_2719,In_1269);
and U1531 (N_1531,In_471,In_2155);
nor U1532 (N_1532,In_1133,In_1260);
and U1533 (N_1533,In_2417,In_1100);
nand U1534 (N_1534,In_950,In_2485);
nor U1535 (N_1535,In_450,In_1611);
nor U1536 (N_1536,In_185,In_347);
xnor U1537 (N_1537,In_2075,In_407);
nand U1538 (N_1538,In_1348,In_1952);
nand U1539 (N_1539,In_85,In_1);
and U1540 (N_1540,In_674,In_600);
nor U1541 (N_1541,In_2302,In_2366);
nand U1542 (N_1542,In_2097,In_2853);
and U1543 (N_1543,In_1071,In_1903);
or U1544 (N_1544,In_1402,In_1934);
nand U1545 (N_1545,In_628,In_1234);
or U1546 (N_1546,In_1109,In_707);
xnor U1547 (N_1547,In_331,In_1172);
nand U1548 (N_1548,In_239,In_2476);
or U1549 (N_1549,In_969,In_2929);
nor U1550 (N_1550,In_138,In_2661);
and U1551 (N_1551,In_1204,In_873);
and U1552 (N_1552,In_2069,In_1359);
or U1553 (N_1553,In_1802,In_1586);
and U1554 (N_1554,In_2068,In_600);
xnor U1555 (N_1555,In_1083,In_128);
and U1556 (N_1556,In_2424,In_1618);
and U1557 (N_1557,In_2742,In_977);
nor U1558 (N_1558,In_1703,In_198);
xnor U1559 (N_1559,In_1686,In_2358);
and U1560 (N_1560,In_1701,In_346);
or U1561 (N_1561,In_2267,In_2123);
and U1562 (N_1562,In_1441,In_1412);
xnor U1563 (N_1563,In_2999,In_1697);
xnor U1564 (N_1564,In_1035,In_2081);
and U1565 (N_1565,In_1960,In_1833);
nand U1566 (N_1566,In_183,In_2597);
or U1567 (N_1567,In_1402,In_2438);
xor U1568 (N_1568,In_958,In_2832);
nand U1569 (N_1569,In_990,In_934);
xor U1570 (N_1570,In_2825,In_2217);
and U1571 (N_1571,In_1569,In_1272);
and U1572 (N_1572,In_2034,In_35);
or U1573 (N_1573,In_1941,In_308);
nand U1574 (N_1574,In_1095,In_2889);
nand U1575 (N_1575,In_2662,In_2546);
or U1576 (N_1576,In_910,In_2319);
nor U1577 (N_1577,In_2009,In_1562);
nand U1578 (N_1578,In_450,In_1295);
nor U1579 (N_1579,In_2653,In_2238);
nand U1580 (N_1580,In_1796,In_662);
nand U1581 (N_1581,In_2015,In_388);
nand U1582 (N_1582,In_2751,In_1585);
nand U1583 (N_1583,In_2643,In_424);
xnor U1584 (N_1584,In_916,In_472);
or U1585 (N_1585,In_222,In_2575);
or U1586 (N_1586,In_595,In_2928);
nand U1587 (N_1587,In_596,In_693);
and U1588 (N_1588,In_1206,In_2816);
and U1589 (N_1589,In_2314,In_567);
and U1590 (N_1590,In_1146,In_2838);
nor U1591 (N_1591,In_2459,In_834);
xor U1592 (N_1592,In_1450,In_2252);
nor U1593 (N_1593,In_1988,In_288);
nand U1594 (N_1594,In_484,In_1275);
or U1595 (N_1595,In_1767,In_1969);
and U1596 (N_1596,In_1530,In_2445);
nor U1597 (N_1597,In_2028,In_2585);
or U1598 (N_1598,In_2486,In_2494);
nand U1599 (N_1599,In_136,In_1657);
nand U1600 (N_1600,In_2967,In_115);
or U1601 (N_1601,In_323,In_1473);
or U1602 (N_1602,In_866,In_1712);
nor U1603 (N_1603,In_1689,In_554);
nand U1604 (N_1604,In_973,In_2966);
or U1605 (N_1605,In_894,In_2379);
and U1606 (N_1606,In_1291,In_1160);
and U1607 (N_1607,In_2544,In_1627);
xor U1608 (N_1608,In_2158,In_2989);
xor U1609 (N_1609,In_2296,In_1906);
and U1610 (N_1610,In_1688,In_1175);
xor U1611 (N_1611,In_2768,In_1885);
xnor U1612 (N_1612,In_2194,In_1749);
nor U1613 (N_1613,In_373,In_2301);
or U1614 (N_1614,In_1866,In_2919);
nand U1615 (N_1615,In_2825,In_2592);
nand U1616 (N_1616,In_1364,In_961);
and U1617 (N_1617,In_83,In_66);
and U1618 (N_1618,In_1235,In_2873);
nand U1619 (N_1619,In_2674,In_586);
nand U1620 (N_1620,In_1421,In_2414);
xor U1621 (N_1621,In_384,In_984);
xor U1622 (N_1622,In_2,In_2917);
nand U1623 (N_1623,In_2453,In_858);
nand U1624 (N_1624,In_2855,In_147);
xnor U1625 (N_1625,In_11,In_145);
nor U1626 (N_1626,In_1816,In_753);
nand U1627 (N_1627,In_1428,In_1884);
and U1628 (N_1628,In_788,In_1460);
nand U1629 (N_1629,In_113,In_2498);
and U1630 (N_1630,In_1149,In_588);
xnor U1631 (N_1631,In_1577,In_1102);
nand U1632 (N_1632,In_1715,In_1005);
nor U1633 (N_1633,In_2574,In_1535);
nor U1634 (N_1634,In_2800,In_1426);
nand U1635 (N_1635,In_877,In_386);
or U1636 (N_1636,In_2900,In_869);
or U1637 (N_1637,In_346,In_981);
nor U1638 (N_1638,In_1535,In_65);
and U1639 (N_1639,In_2101,In_1295);
or U1640 (N_1640,In_86,In_2368);
nor U1641 (N_1641,In_810,In_1937);
xor U1642 (N_1642,In_2025,In_2866);
nand U1643 (N_1643,In_903,In_2455);
xnor U1644 (N_1644,In_1841,In_1898);
nor U1645 (N_1645,In_950,In_2333);
and U1646 (N_1646,In_1616,In_2601);
xnor U1647 (N_1647,In_2397,In_236);
nand U1648 (N_1648,In_1630,In_1881);
and U1649 (N_1649,In_2997,In_2896);
nand U1650 (N_1650,In_869,In_116);
or U1651 (N_1651,In_1252,In_892);
and U1652 (N_1652,In_727,In_2819);
xnor U1653 (N_1653,In_2898,In_1567);
nand U1654 (N_1654,In_155,In_1880);
or U1655 (N_1655,In_2689,In_2345);
nor U1656 (N_1656,In_1280,In_2474);
or U1657 (N_1657,In_676,In_2618);
or U1658 (N_1658,In_1408,In_2412);
nand U1659 (N_1659,In_1231,In_2141);
and U1660 (N_1660,In_2394,In_2702);
xnor U1661 (N_1661,In_446,In_1747);
xnor U1662 (N_1662,In_2550,In_299);
or U1663 (N_1663,In_1331,In_1216);
xor U1664 (N_1664,In_836,In_2796);
nand U1665 (N_1665,In_1157,In_2568);
or U1666 (N_1666,In_2766,In_46);
and U1667 (N_1667,In_687,In_1555);
or U1668 (N_1668,In_1398,In_2524);
and U1669 (N_1669,In_1927,In_2356);
xor U1670 (N_1670,In_2554,In_892);
and U1671 (N_1671,In_2158,In_2122);
xnor U1672 (N_1672,In_277,In_1328);
xor U1673 (N_1673,In_2329,In_405);
nor U1674 (N_1674,In_574,In_2787);
nand U1675 (N_1675,In_553,In_1470);
xor U1676 (N_1676,In_2920,In_2409);
or U1677 (N_1677,In_1865,In_2140);
and U1678 (N_1678,In_1825,In_1559);
xnor U1679 (N_1679,In_28,In_344);
or U1680 (N_1680,In_2247,In_564);
and U1681 (N_1681,In_1414,In_2913);
nand U1682 (N_1682,In_878,In_2775);
and U1683 (N_1683,In_211,In_1481);
or U1684 (N_1684,In_578,In_1811);
or U1685 (N_1685,In_741,In_2687);
and U1686 (N_1686,In_2574,In_85);
xor U1687 (N_1687,In_1658,In_1908);
and U1688 (N_1688,In_554,In_1412);
or U1689 (N_1689,In_66,In_794);
nand U1690 (N_1690,In_112,In_1093);
nand U1691 (N_1691,In_2077,In_2382);
nor U1692 (N_1692,In_2582,In_795);
or U1693 (N_1693,In_1599,In_2748);
nand U1694 (N_1694,In_1088,In_560);
and U1695 (N_1695,In_1896,In_1305);
or U1696 (N_1696,In_1740,In_119);
or U1697 (N_1697,In_1705,In_2260);
xnor U1698 (N_1698,In_1379,In_111);
xor U1699 (N_1699,In_808,In_1222);
or U1700 (N_1700,In_2072,In_118);
nand U1701 (N_1701,In_405,In_2550);
or U1702 (N_1702,In_1661,In_793);
nand U1703 (N_1703,In_979,In_1435);
and U1704 (N_1704,In_1912,In_2445);
nor U1705 (N_1705,In_2762,In_1587);
and U1706 (N_1706,In_610,In_1849);
nor U1707 (N_1707,In_1569,In_1220);
xor U1708 (N_1708,In_2604,In_882);
and U1709 (N_1709,In_1368,In_77);
xnor U1710 (N_1710,In_2225,In_1300);
and U1711 (N_1711,In_1166,In_1020);
nand U1712 (N_1712,In_2189,In_1482);
and U1713 (N_1713,In_703,In_1594);
and U1714 (N_1714,In_1459,In_276);
nor U1715 (N_1715,In_249,In_2644);
nor U1716 (N_1716,In_710,In_337);
and U1717 (N_1717,In_511,In_2251);
nand U1718 (N_1718,In_1694,In_2436);
and U1719 (N_1719,In_1103,In_653);
or U1720 (N_1720,In_812,In_2475);
nor U1721 (N_1721,In_2387,In_1897);
and U1722 (N_1722,In_1112,In_2793);
and U1723 (N_1723,In_2786,In_542);
and U1724 (N_1724,In_571,In_1942);
or U1725 (N_1725,In_424,In_1568);
and U1726 (N_1726,In_957,In_2219);
or U1727 (N_1727,In_2324,In_2182);
xor U1728 (N_1728,In_1654,In_1139);
xnor U1729 (N_1729,In_898,In_1083);
nand U1730 (N_1730,In_537,In_2538);
nor U1731 (N_1731,In_926,In_114);
nor U1732 (N_1732,In_47,In_920);
nor U1733 (N_1733,In_834,In_1898);
and U1734 (N_1734,In_2387,In_299);
nor U1735 (N_1735,In_1116,In_473);
nor U1736 (N_1736,In_624,In_452);
nand U1737 (N_1737,In_1388,In_2759);
nand U1738 (N_1738,In_290,In_2457);
nor U1739 (N_1739,In_1243,In_349);
and U1740 (N_1740,In_179,In_2022);
and U1741 (N_1741,In_2356,In_2667);
and U1742 (N_1742,In_1895,In_1312);
nor U1743 (N_1743,In_1043,In_2363);
and U1744 (N_1744,In_1607,In_1496);
nor U1745 (N_1745,In_1237,In_1233);
or U1746 (N_1746,In_1964,In_2391);
or U1747 (N_1747,In_780,In_166);
and U1748 (N_1748,In_838,In_321);
xnor U1749 (N_1749,In_2046,In_2588);
and U1750 (N_1750,In_455,In_2634);
nor U1751 (N_1751,In_1872,In_2870);
nand U1752 (N_1752,In_228,In_1590);
xnor U1753 (N_1753,In_253,In_1348);
nand U1754 (N_1754,In_1229,In_1103);
xor U1755 (N_1755,In_625,In_1943);
or U1756 (N_1756,In_2305,In_1638);
and U1757 (N_1757,In_2787,In_242);
nor U1758 (N_1758,In_1405,In_294);
nand U1759 (N_1759,In_2511,In_1028);
nand U1760 (N_1760,In_2367,In_1433);
or U1761 (N_1761,In_1106,In_2232);
or U1762 (N_1762,In_742,In_301);
xnor U1763 (N_1763,In_2232,In_1226);
nand U1764 (N_1764,In_473,In_1727);
and U1765 (N_1765,In_149,In_786);
nand U1766 (N_1766,In_2445,In_2215);
xnor U1767 (N_1767,In_1799,In_278);
or U1768 (N_1768,In_1686,In_1453);
nor U1769 (N_1769,In_1569,In_324);
nand U1770 (N_1770,In_246,In_1972);
xnor U1771 (N_1771,In_1970,In_634);
xnor U1772 (N_1772,In_1631,In_2393);
xor U1773 (N_1773,In_1422,In_2484);
nand U1774 (N_1774,In_846,In_852);
nand U1775 (N_1775,In_2402,In_2141);
nor U1776 (N_1776,In_2863,In_1199);
xnor U1777 (N_1777,In_1467,In_807);
or U1778 (N_1778,In_463,In_1169);
or U1779 (N_1779,In_1923,In_2617);
xnor U1780 (N_1780,In_2850,In_1021);
or U1781 (N_1781,In_1125,In_1993);
and U1782 (N_1782,In_753,In_686);
and U1783 (N_1783,In_1738,In_1205);
or U1784 (N_1784,In_2018,In_2021);
and U1785 (N_1785,In_293,In_2318);
or U1786 (N_1786,In_207,In_406);
nor U1787 (N_1787,In_2949,In_1683);
xor U1788 (N_1788,In_2918,In_466);
or U1789 (N_1789,In_606,In_1929);
xor U1790 (N_1790,In_2602,In_1582);
and U1791 (N_1791,In_2252,In_1852);
or U1792 (N_1792,In_459,In_2574);
nor U1793 (N_1793,In_2040,In_875);
and U1794 (N_1794,In_1834,In_22);
xnor U1795 (N_1795,In_2440,In_2496);
and U1796 (N_1796,In_800,In_2122);
nand U1797 (N_1797,In_2095,In_1329);
nor U1798 (N_1798,In_2803,In_1380);
nor U1799 (N_1799,In_1935,In_24);
nand U1800 (N_1800,In_2923,In_1589);
nand U1801 (N_1801,In_2865,In_2032);
or U1802 (N_1802,In_185,In_2063);
nor U1803 (N_1803,In_2722,In_583);
and U1804 (N_1804,In_1868,In_337);
and U1805 (N_1805,In_234,In_1694);
or U1806 (N_1806,In_1832,In_2478);
xnor U1807 (N_1807,In_2354,In_1578);
xnor U1808 (N_1808,In_894,In_1341);
or U1809 (N_1809,In_1472,In_1615);
and U1810 (N_1810,In_399,In_827);
nor U1811 (N_1811,In_2506,In_484);
and U1812 (N_1812,In_2488,In_879);
and U1813 (N_1813,In_2833,In_503);
xnor U1814 (N_1814,In_68,In_2391);
nor U1815 (N_1815,In_957,In_1082);
and U1816 (N_1816,In_632,In_1490);
nor U1817 (N_1817,In_2445,In_1998);
or U1818 (N_1818,In_2459,In_723);
or U1819 (N_1819,In_2485,In_1141);
nand U1820 (N_1820,In_2049,In_1937);
and U1821 (N_1821,In_2399,In_667);
or U1822 (N_1822,In_2657,In_412);
or U1823 (N_1823,In_354,In_2065);
xnor U1824 (N_1824,In_2817,In_2894);
or U1825 (N_1825,In_2728,In_252);
nand U1826 (N_1826,In_1800,In_2070);
nor U1827 (N_1827,In_310,In_1962);
nor U1828 (N_1828,In_471,In_1793);
nand U1829 (N_1829,In_2833,In_128);
nand U1830 (N_1830,In_149,In_1889);
nand U1831 (N_1831,In_112,In_2765);
nand U1832 (N_1832,In_1735,In_2648);
or U1833 (N_1833,In_803,In_2784);
and U1834 (N_1834,In_1663,In_590);
xor U1835 (N_1835,In_238,In_1948);
or U1836 (N_1836,In_1816,In_2718);
or U1837 (N_1837,In_1982,In_923);
or U1838 (N_1838,In_681,In_2288);
or U1839 (N_1839,In_2784,In_1793);
or U1840 (N_1840,In_1336,In_1816);
and U1841 (N_1841,In_2658,In_143);
nand U1842 (N_1842,In_138,In_2638);
and U1843 (N_1843,In_2104,In_212);
xnor U1844 (N_1844,In_1267,In_2372);
nand U1845 (N_1845,In_1602,In_1757);
xor U1846 (N_1846,In_2427,In_1399);
nor U1847 (N_1847,In_2598,In_1528);
or U1848 (N_1848,In_129,In_1438);
nand U1849 (N_1849,In_1824,In_2218);
or U1850 (N_1850,In_1907,In_455);
nor U1851 (N_1851,In_309,In_1070);
xnor U1852 (N_1852,In_679,In_1001);
or U1853 (N_1853,In_490,In_478);
nor U1854 (N_1854,In_2754,In_2622);
or U1855 (N_1855,In_247,In_1064);
or U1856 (N_1856,In_2212,In_2033);
nand U1857 (N_1857,In_2659,In_153);
nor U1858 (N_1858,In_524,In_1365);
and U1859 (N_1859,In_232,In_2832);
nor U1860 (N_1860,In_1215,In_2402);
or U1861 (N_1861,In_494,In_1167);
nor U1862 (N_1862,In_647,In_2441);
nand U1863 (N_1863,In_2835,In_1464);
and U1864 (N_1864,In_729,In_1269);
nand U1865 (N_1865,In_1647,In_1728);
or U1866 (N_1866,In_2872,In_1336);
nand U1867 (N_1867,In_1549,In_338);
and U1868 (N_1868,In_2612,In_2751);
xnor U1869 (N_1869,In_1734,In_1377);
nor U1870 (N_1870,In_2276,In_1417);
nor U1871 (N_1871,In_1215,In_1502);
nand U1872 (N_1872,In_2591,In_14);
and U1873 (N_1873,In_2051,In_1082);
xnor U1874 (N_1874,In_2450,In_2814);
and U1875 (N_1875,In_1735,In_26);
xor U1876 (N_1876,In_1387,In_2321);
and U1877 (N_1877,In_560,In_2430);
or U1878 (N_1878,In_1189,In_624);
nand U1879 (N_1879,In_127,In_935);
xor U1880 (N_1880,In_682,In_94);
and U1881 (N_1881,In_2448,In_1805);
or U1882 (N_1882,In_1952,In_2073);
nand U1883 (N_1883,In_13,In_2217);
and U1884 (N_1884,In_2423,In_1894);
nand U1885 (N_1885,In_2789,In_29);
nor U1886 (N_1886,In_2048,In_2442);
nand U1887 (N_1887,In_905,In_2261);
nand U1888 (N_1888,In_482,In_1618);
xnor U1889 (N_1889,In_945,In_2957);
nand U1890 (N_1890,In_948,In_1901);
or U1891 (N_1891,In_398,In_2953);
nand U1892 (N_1892,In_1485,In_1985);
xor U1893 (N_1893,In_337,In_2099);
or U1894 (N_1894,In_898,In_251);
or U1895 (N_1895,In_2804,In_277);
nor U1896 (N_1896,In_406,In_1505);
and U1897 (N_1897,In_308,In_1715);
nor U1898 (N_1898,In_2669,In_1073);
xor U1899 (N_1899,In_2806,In_2703);
or U1900 (N_1900,In_474,In_2173);
or U1901 (N_1901,In_262,In_1402);
and U1902 (N_1902,In_1861,In_1724);
or U1903 (N_1903,In_528,In_1175);
or U1904 (N_1904,In_862,In_953);
xnor U1905 (N_1905,In_2270,In_397);
or U1906 (N_1906,In_1903,In_2787);
nor U1907 (N_1907,In_2116,In_2286);
or U1908 (N_1908,In_2890,In_365);
nor U1909 (N_1909,In_1458,In_1369);
nor U1910 (N_1910,In_2234,In_649);
nand U1911 (N_1911,In_1693,In_222);
xor U1912 (N_1912,In_862,In_900);
and U1913 (N_1913,In_1891,In_280);
nor U1914 (N_1914,In_2493,In_654);
or U1915 (N_1915,In_1155,In_143);
and U1916 (N_1916,In_1824,In_1369);
and U1917 (N_1917,In_1615,In_725);
nor U1918 (N_1918,In_1703,In_1640);
and U1919 (N_1919,In_2413,In_2744);
nor U1920 (N_1920,In_961,In_1933);
nand U1921 (N_1921,In_2701,In_945);
and U1922 (N_1922,In_1987,In_596);
nor U1923 (N_1923,In_547,In_1603);
xnor U1924 (N_1924,In_2624,In_686);
nor U1925 (N_1925,In_2754,In_1010);
or U1926 (N_1926,In_2326,In_2983);
and U1927 (N_1927,In_642,In_685);
or U1928 (N_1928,In_1223,In_817);
or U1929 (N_1929,In_1551,In_2676);
nand U1930 (N_1930,In_858,In_328);
and U1931 (N_1931,In_1022,In_2822);
nor U1932 (N_1932,In_429,In_1634);
nand U1933 (N_1933,In_2784,In_561);
nor U1934 (N_1934,In_694,In_846);
nand U1935 (N_1935,In_2172,In_1216);
xor U1936 (N_1936,In_253,In_2127);
or U1937 (N_1937,In_1474,In_1976);
or U1938 (N_1938,In_372,In_938);
and U1939 (N_1939,In_334,In_2151);
xnor U1940 (N_1940,In_743,In_648);
nand U1941 (N_1941,In_2505,In_21);
nor U1942 (N_1942,In_1342,In_2352);
nor U1943 (N_1943,In_1394,In_2627);
xor U1944 (N_1944,In_1155,In_664);
xnor U1945 (N_1945,In_2193,In_315);
nand U1946 (N_1946,In_59,In_1150);
nor U1947 (N_1947,In_2265,In_1155);
xnor U1948 (N_1948,In_261,In_2073);
or U1949 (N_1949,In_2957,In_42);
nand U1950 (N_1950,In_325,In_2514);
xor U1951 (N_1951,In_1859,In_2066);
or U1952 (N_1952,In_2189,In_1323);
and U1953 (N_1953,In_753,In_1023);
or U1954 (N_1954,In_825,In_2215);
xor U1955 (N_1955,In_1221,In_2601);
xnor U1956 (N_1956,In_1172,In_2086);
or U1957 (N_1957,In_2503,In_1817);
and U1958 (N_1958,In_774,In_2896);
nand U1959 (N_1959,In_1664,In_1733);
nand U1960 (N_1960,In_272,In_2633);
nand U1961 (N_1961,In_2526,In_917);
xor U1962 (N_1962,In_1390,In_2563);
nor U1963 (N_1963,In_2847,In_395);
xor U1964 (N_1964,In_1404,In_1750);
nor U1965 (N_1965,In_1187,In_2603);
xnor U1966 (N_1966,In_2512,In_994);
xnor U1967 (N_1967,In_606,In_1052);
and U1968 (N_1968,In_1039,In_592);
nor U1969 (N_1969,In_2869,In_420);
or U1970 (N_1970,In_948,In_1379);
nand U1971 (N_1971,In_2660,In_790);
and U1972 (N_1972,In_626,In_2653);
nand U1973 (N_1973,In_220,In_432);
or U1974 (N_1974,In_870,In_396);
nand U1975 (N_1975,In_2550,In_1056);
or U1976 (N_1976,In_2215,In_2907);
nor U1977 (N_1977,In_755,In_1085);
nor U1978 (N_1978,In_1494,In_2943);
and U1979 (N_1979,In_404,In_2886);
and U1980 (N_1980,In_304,In_2061);
nor U1981 (N_1981,In_1466,In_656);
or U1982 (N_1982,In_2132,In_2744);
xnor U1983 (N_1983,In_514,In_2306);
or U1984 (N_1984,In_455,In_2025);
nor U1985 (N_1985,In_105,In_1427);
and U1986 (N_1986,In_1777,In_2816);
nor U1987 (N_1987,In_2024,In_1038);
or U1988 (N_1988,In_1438,In_2348);
nand U1989 (N_1989,In_2763,In_1333);
nand U1990 (N_1990,In_1867,In_2674);
or U1991 (N_1991,In_1883,In_951);
nand U1992 (N_1992,In_1801,In_1956);
and U1993 (N_1993,In_1527,In_617);
xnor U1994 (N_1994,In_2103,In_2918);
nand U1995 (N_1995,In_1444,In_1484);
xnor U1996 (N_1996,In_220,In_2047);
nand U1997 (N_1997,In_2250,In_1371);
nor U1998 (N_1998,In_169,In_1199);
or U1999 (N_1999,In_2467,In_1940);
and U2000 (N_2000,In_1165,In_627);
or U2001 (N_2001,In_1388,In_982);
or U2002 (N_2002,In_607,In_246);
and U2003 (N_2003,In_1955,In_2486);
xnor U2004 (N_2004,In_1426,In_643);
nor U2005 (N_2005,In_2459,In_1772);
xor U2006 (N_2006,In_2340,In_2083);
nor U2007 (N_2007,In_1924,In_613);
nor U2008 (N_2008,In_2794,In_981);
nor U2009 (N_2009,In_43,In_2069);
nand U2010 (N_2010,In_2644,In_1643);
nor U2011 (N_2011,In_2155,In_1611);
xor U2012 (N_2012,In_135,In_1385);
nand U2013 (N_2013,In_1712,In_2965);
nand U2014 (N_2014,In_2335,In_2856);
or U2015 (N_2015,In_2534,In_2606);
nor U2016 (N_2016,In_2036,In_2583);
and U2017 (N_2017,In_1172,In_2100);
or U2018 (N_2018,In_2569,In_148);
xnor U2019 (N_2019,In_648,In_707);
nor U2020 (N_2020,In_833,In_2480);
xnor U2021 (N_2021,In_1973,In_1180);
and U2022 (N_2022,In_1880,In_2942);
xor U2023 (N_2023,In_302,In_1811);
nor U2024 (N_2024,In_1625,In_1820);
xnor U2025 (N_2025,In_1965,In_1051);
nor U2026 (N_2026,In_248,In_1437);
or U2027 (N_2027,In_84,In_1667);
and U2028 (N_2028,In_772,In_2501);
or U2029 (N_2029,In_2265,In_2558);
xor U2030 (N_2030,In_2163,In_2778);
and U2031 (N_2031,In_219,In_1983);
xor U2032 (N_2032,In_2564,In_13);
or U2033 (N_2033,In_1695,In_283);
nor U2034 (N_2034,In_2587,In_525);
xnor U2035 (N_2035,In_1194,In_905);
or U2036 (N_2036,In_1555,In_91);
or U2037 (N_2037,In_2253,In_1606);
nand U2038 (N_2038,In_1627,In_954);
nand U2039 (N_2039,In_1788,In_2245);
nor U2040 (N_2040,In_1372,In_1182);
or U2041 (N_2041,In_624,In_848);
and U2042 (N_2042,In_2896,In_1812);
or U2043 (N_2043,In_2877,In_1987);
and U2044 (N_2044,In_997,In_1040);
or U2045 (N_2045,In_45,In_1324);
or U2046 (N_2046,In_1963,In_2994);
or U2047 (N_2047,In_1916,In_2369);
or U2048 (N_2048,In_875,In_1276);
and U2049 (N_2049,In_1444,In_1726);
and U2050 (N_2050,In_1950,In_1168);
and U2051 (N_2051,In_2946,In_1373);
nand U2052 (N_2052,In_580,In_2889);
nand U2053 (N_2053,In_1000,In_2122);
nand U2054 (N_2054,In_1457,In_1117);
nor U2055 (N_2055,In_1559,In_328);
xnor U2056 (N_2056,In_43,In_1101);
nand U2057 (N_2057,In_971,In_1326);
nor U2058 (N_2058,In_2471,In_1077);
nand U2059 (N_2059,In_1089,In_1245);
nor U2060 (N_2060,In_2330,In_588);
and U2061 (N_2061,In_2671,In_2473);
nor U2062 (N_2062,In_1847,In_2761);
xnor U2063 (N_2063,In_2830,In_785);
xnor U2064 (N_2064,In_967,In_2100);
xnor U2065 (N_2065,In_475,In_2562);
xnor U2066 (N_2066,In_1041,In_2288);
xor U2067 (N_2067,In_1432,In_2482);
or U2068 (N_2068,In_933,In_84);
and U2069 (N_2069,In_1851,In_2103);
xnor U2070 (N_2070,In_2288,In_2828);
nand U2071 (N_2071,In_892,In_2057);
nand U2072 (N_2072,In_1978,In_2487);
xor U2073 (N_2073,In_87,In_1278);
nor U2074 (N_2074,In_1449,In_2133);
and U2075 (N_2075,In_2668,In_1968);
or U2076 (N_2076,In_60,In_1215);
and U2077 (N_2077,In_2761,In_1657);
nand U2078 (N_2078,In_2537,In_520);
xnor U2079 (N_2079,In_1023,In_2005);
nor U2080 (N_2080,In_2313,In_2926);
and U2081 (N_2081,In_1259,In_2221);
nand U2082 (N_2082,In_2680,In_1472);
nor U2083 (N_2083,In_558,In_1546);
nor U2084 (N_2084,In_2687,In_763);
xnor U2085 (N_2085,In_436,In_390);
nand U2086 (N_2086,In_1302,In_1037);
nor U2087 (N_2087,In_1757,In_2836);
xnor U2088 (N_2088,In_2536,In_1651);
and U2089 (N_2089,In_3,In_1093);
nor U2090 (N_2090,In_369,In_2693);
nand U2091 (N_2091,In_695,In_2349);
xor U2092 (N_2092,In_1634,In_2366);
nand U2093 (N_2093,In_952,In_1699);
xor U2094 (N_2094,In_2731,In_1579);
xor U2095 (N_2095,In_2530,In_1429);
nand U2096 (N_2096,In_2257,In_2379);
xor U2097 (N_2097,In_161,In_1688);
and U2098 (N_2098,In_97,In_909);
xnor U2099 (N_2099,In_2329,In_1590);
and U2100 (N_2100,In_2631,In_1431);
nor U2101 (N_2101,In_1646,In_2149);
nor U2102 (N_2102,In_137,In_2451);
xnor U2103 (N_2103,In_1118,In_896);
or U2104 (N_2104,In_214,In_2739);
nand U2105 (N_2105,In_2756,In_163);
nand U2106 (N_2106,In_2887,In_2768);
and U2107 (N_2107,In_1342,In_551);
xnor U2108 (N_2108,In_1716,In_2843);
and U2109 (N_2109,In_805,In_2807);
xor U2110 (N_2110,In_1491,In_1970);
nor U2111 (N_2111,In_1552,In_2780);
nor U2112 (N_2112,In_2028,In_2784);
nor U2113 (N_2113,In_2801,In_771);
nor U2114 (N_2114,In_593,In_1273);
nor U2115 (N_2115,In_547,In_1721);
or U2116 (N_2116,In_2765,In_1675);
or U2117 (N_2117,In_2007,In_2168);
or U2118 (N_2118,In_178,In_2501);
nor U2119 (N_2119,In_2760,In_1794);
nand U2120 (N_2120,In_2463,In_2717);
and U2121 (N_2121,In_1455,In_989);
or U2122 (N_2122,In_1680,In_93);
or U2123 (N_2123,In_27,In_910);
nor U2124 (N_2124,In_947,In_1361);
and U2125 (N_2125,In_1622,In_1627);
and U2126 (N_2126,In_180,In_438);
xnor U2127 (N_2127,In_102,In_2853);
and U2128 (N_2128,In_1035,In_969);
xnor U2129 (N_2129,In_460,In_1311);
nand U2130 (N_2130,In_168,In_626);
xor U2131 (N_2131,In_2734,In_1039);
or U2132 (N_2132,In_69,In_253);
nand U2133 (N_2133,In_165,In_1544);
nor U2134 (N_2134,In_1296,In_772);
xnor U2135 (N_2135,In_1747,In_2057);
or U2136 (N_2136,In_2623,In_2728);
nand U2137 (N_2137,In_1691,In_2699);
and U2138 (N_2138,In_934,In_6);
nand U2139 (N_2139,In_2283,In_585);
or U2140 (N_2140,In_2516,In_257);
or U2141 (N_2141,In_2165,In_1666);
and U2142 (N_2142,In_1939,In_933);
nand U2143 (N_2143,In_502,In_2617);
xor U2144 (N_2144,In_2687,In_587);
xor U2145 (N_2145,In_1637,In_48);
or U2146 (N_2146,In_2417,In_2151);
xor U2147 (N_2147,In_752,In_1115);
nand U2148 (N_2148,In_1620,In_2981);
or U2149 (N_2149,In_1262,In_303);
xnor U2150 (N_2150,In_793,In_817);
and U2151 (N_2151,In_833,In_366);
and U2152 (N_2152,In_1288,In_534);
and U2153 (N_2153,In_1862,In_1206);
and U2154 (N_2154,In_2503,In_1745);
or U2155 (N_2155,In_1902,In_2970);
or U2156 (N_2156,In_2792,In_1241);
nor U2157 (N_2157,In_1489,In_1415);
nor U2158 (N_2158,In_2013,In_420);
and U2159 (N_2159,In_2432,In_2209);
or U2160 (N_2160,In_859,In_181);
nor U2161 (N_2161,In_2446,In_1929);
nand U2162 (N_2162,In_136,In_1118);
xor U2163 (N_2163,In_1238,In_1380);
xor U2164 (N_2164,In_66,In_161);
nor U2165 (N_2165,In_775,In_662);
or U2166 (N_2166,In_611,In_1545);
nand U2167 (N_2167,In_2300,In_2172);
and U2168 (N_2168,In_1877,In_2304);
or U2169 (N_2169,In_2813,In_2629);
nand U2170 (N_2170,In_1468,In_1007);
nand U2171 (N_2171,In_232,In_2700);
and U2172 (N_2172,In_2410,In_2857);
and U2173 (N_2173,In_1439,In_2406);
and U2174 (N_2174,In_1054,In_2033);
nor U2175 (N_2175,In_1275,In_1343);
nand U2176 (N_2176,In_882,In_1268);
xnor U2177 (N_2177,In_887,In_2011);
and U2178 (N_2178,In_673,In_356);
nand U2179 (N_2179,In_416,In_2108);
xnor U2180 (N_2180,In_1804,In_252);
or U2181 (N_2181,In_1590,In_2051);
and U2182 (N_2182,In_2639,In_941);
nand U2183 (N_2183,In_2277,In_1066);
and U2184 (N_2184,In_261,In_2665);
nand U2185 (N_2185,In_2378,In_739);
or U2186 (N_2186,In_518,In_261);
or U2187 (N_2187,In_134,In_42);
nor U2188 (N_2188,In_2377,In_2758);
nand U2189 (N_2189,In_2849,In_129);
and U2190 (N_2190,In_1578,In_905);
or U2191 (N_2191,In_970,In_518);
nor U2192 (N_2192,In_2342,In_1966);
xnor U2193 (N_2193,In_2901,In_2280);
nand U2194 (N_2194,In_1811,In_411);
nor U2195 (N_2195,In_863,In_104);
nor U2196 (N_2196,In_1000,In_2670);
nand U2197 (N_2197,In_1280,In_2226);
xor U2198 (N_2198,In_419,In_723);
and U2199 (N_2199,In_216,In_845);
or U2200 (N_2200,In_2537,In_2342);
nand U2201 (N_2201,In_1432,In_2538);
nor U2202 (N_2202,In_1556,In_2802);
and U2203 (N_2203,In_1571,In_464);
and U2204 (N_2204,In_1335,In_311);
nand U2205 (N_2205,In_2850,In_2286);
xnor U2206 (N_2206,In_595,In_2523);
xnor U2207 (N_2207,In_1082,In_2703);
and U2208 (N_2208,In_1936,In_383);
and U2209 (N_2209,In_378,In_1831);
nand U2210 (N_2210,In_2530,In_1815);
nor U2211 (N_2211,In_1272,In_808);
and U2212 (N_2212,In_2331,In_474);
xnor U2213 (N_2213,In_2581,In_2535);
nor U2214 (N_2214,In_326,In_41);
nor U2215 (N_2215,In_774,In_2780);
nor U2216 (N_2216,In_517,In_972);
nand U2217 (N_2217,In_1482,In_123);
and U2218 (N_2218,In_2927,In_464);
or U2219 (N_2219,In_707,In_380);
nand U2220 (N_2220,In_1105,In_2377);
or U2221 (N_2221,In_1220,In_216);
and U2222 (N_2222,In_251,In_1367);
nand U2223 (N_2223,In_1044,In_1298);
xor U2224 (N_2224,In_383,In_1228);
xnor U2225 (N_2225,In_2485,In_1549);
or U2226 (N_2226,In_1476,In_1007);
or U2227 (N_2227,In_200,In_513);
or U2228 (N_2228,In_1017,In_2769);
xnor U2229 (N_2229,In_1226,In_796);
xnor U2230 (N_2230,In_2882,In_2070);
nor U2231 (N_2231,In_562,In_2229);
nand U2232 (N_2232,In_1602,In_919);
and U2233 (N_2233,In_2542,In_1018);
xor U2234 (N_2234,In_295,In_293);
xnor U2235 (N_2235,In_1591,In_408);
and U2236 (N_2236,In_253,In_1281);
nand U2237 (N_2237,In_871,In_462);
nor U2238 (N_2238,In_191,In_306);
xnor U2239 (N_2239,In_2467,In_1088);
or U2240 (N_2240,In_2877,In_2555);
and U2241 (N_2241,In_1375,In_1566);
or U2242 (N_2242,In_2174,In_115);
nor U2243 (N_2243,In_246,In_2586);
nand U2244 (N_2244,In_2906,In_1797);
and U2245 (N_2245,In_2563,In_2222);
nand U2246 (N_2246,In_1099,In_1059);
and U2247 (N_2247,In_716,In_53);
or U2248 (N_2248,In_2394,In_2021);
and U2249 (N_2249,In_2770,In_410);
nand U2250 (N_2250,In_2339,In_2371);
or U2251 (N_2251,In_2010,In_2134);
xnor U2252 (N_2252,In_1228,In_815);
xor U2253 (N_2253,In_305,In_2);
nand U2254 (N_2254,In_139,In_249);
or U2255 (N_2255,In_2197,In_2255);
and U2256 (N_2256,In_53,In_185);
or U2257 (N_2257,In_1371,In_2427);
xor U2258 (N_2258,In_1488,In_2706);
nand U2259 (N_2259,In_2714,In_456);
or U2260 (N_2260,In_2774,In_2372);
nand U2261 (N_2261,In_1124,In_1197);
nand U2262 (N_2262,In_472,In_1301);
nand U2263 (N_2263,In_1183,In_1557);
xnor U2264 (N_2264,In_2890,In_2112);
nand U2265 (N_2265,In_2797,In_2437);
nor U2266 (N_2266,In_882,In_2110);
or U2267 (N_2267,In_1815,In_2966);
xnor U2268 (N_2268,In_442,In_322);
or U2269 (N_2269,In_2667,In_1795);
xnor U2270 (N_2270,In_2687,In_2296);
or U2271 (N_2271,In_790,In_359);
nand U2272 (N_2272,In_870,In_625);
nand U2273 (N_2273,In_2743,In_2043);
nand U2274 (N_2274,In_535,In_1605);
nand U2275 (N_2275,In_1800,In_75);
xor U2276 (N_2276,In_1411,In_493);
nand U2277 (N_2277,In_1303,In_1274);
nor U2278 (N_2278,In_1583,In_2371);
and U2279 (N_2279,In_261,In_636);
xor U2280 (N_2280,In_2398,In_1876);
nand U2281 (N_2281,In_1481,In_1310);
nor U2282 (N_2282,In_2714,In_2275);
or U2283 (N_2283,In_5,In_2459);
nor U2284 (N_2284,In_718,In_2764);
nor U2285 (N_2285,In_2494,In_2691);
nand U2286 (N_2286,In_91,In_1507);
or U2287 (N_2287,In_541,In_2993);
or U2288 (N_2288,In_2178,In_1072);
nor U2289 (N_2289,In_1650,In_1898);
nor U2290 (N_2290,In_1169,In_2724);
xor U2291 (N_2291,In_761,In_1515);
nor U2292 (N_2292,In_1621,In_580);
nand U2293 (N_2293,In_1229,In_232);
and U2294 (N_2294,In_336,In_795);
xor U2295 (N_2295,In_2104,In_1531);
nand U2296 (N_2296,In_1277,In_1437);
or U2297 (N_2297,In_8,In_2220);
xnor U2298 (N_2298,In_674,In_1128);
nor U2299 (N_2299,In_2300,In_2771);
nor U2300 (N_2300,In_1366,In_1878);
nand U2301 (N_2301,In_834,In_1135);
nand U2302 (N_2302,In_2083,In_2842);
nand U2303 (N_2303,In_848,In_396);
xor U2304 (N_2304,In_2157,In_1232);
xor U2305 (N_2305,In_1832,In_1328);
and U2306 (N_2306,In_2992,In_415);
nor U2307 (N_2307,In_2965,In_2150);
nor U2308 (N_2308,In_2415,In_895);
and U2309 (N_2309,In_225,In_137);
and U2310 (N_2310,In_808,In_95);
nor U2311 (N_2311,In_1834,In_608);
nor U2312 (N_2312,In_251,In_1900);
xor U2313 (N_2313,In_240,In_565);
xnor U2314 (N_2314,In_416,In_807);
xnor U2315 (N_2315,In_395,In_1935);
and U2316 (N_2316,In_2111,In_265);
nor U2317 (N_2317,In_178,In_1606);
and U2318 (N_2318,In_1777,In_787);
xnor U2319 (N_2319,In_2881,In_675);
nand U2320 (N_2320,In_1085,In_1171);
nor U2321 (N_2321,In_71,In_144);
and U2322 (N_2322,In_680,In_1153);
nor U2323 (N_2323,In_2565,In_2212);
and U2324 (N_2324,In_1132,In_789);
xor U2325 (N_2325,In_641,In_694);
or U2326 (N_2326,In_1288,In_196);
nand U2327 (N_2327,In_2144,In_489);
nand U2328 (N_2328,In_1733,In_744);
or U2329 (N_2329,In_1217,In_799);
nor U2330 (N_2330,In_6,In_737);
xnor U2331 (N_2331,In_1381,In_1918);
and U2332 (N_2332,In_2431,In_1875);
xnor U2333 (N_2333,In_2451,In_2879);
or U2334 (N_2334,In_1708,In_1914);
xor U2335 (N_2335,In_1798,In_2596);
or U2336 (N_2336,In_2533,In_1063);
and U2337 (N_2337,In_547,In_376);
nor U2338 (N_2338,In_2451,In_774);
and U2339 (N_2339,In_824,In_392);
nor U2340 (N_2340,In_1456,In_2841);
xor U2341 (N_2341,In_1776,In_1415);
or U2342 (N_2342,In_513,In_2516);
nor U2343 (N_2343,In_424,In_2958);
xnor U2344 (N_2344,In_8,In_2255);
nand U2345 (N_2345,In_134,In_1911);
xor U2346 (N_2346,In_630,In_620);
xor U2347 (N_2347,In_910,In_582);
or U2348 (N_2348,In_2565,In_2638);
and U2349 (N_2349,In_2417,In_1214);
or U2350 (N_2350,In_2884,In_2045);
or U2351 (N_2351,In_977,In_193);
or U2352 (N_2352,In_119,In_543);
and U2353 (N_2353,In_2428,In_529);
nor U2354 (N_2354,In_963,In_1213);
nand U2355 (N_2355,In_2583,In_790);
or U2356 (N_2356,In_2634,In_1978);
nor U2357 (N_2357,In_2018,In_1224);
nor U2358 (N_2358,In_2172,In_1244);
or U2359 (N_2359,In_1036,In_2046);
nand U2360 (N_2360,In_2335,In_1699);
nor U2361 (N_2361,In_2037,In_2789);
or U2362 (N_2362,In_1603,In_2374);
or U2363 (N_2363,In_2067,In_2287);
or U2364 (N_2364,In_2943,In_1096);
or U2365 (N_2365,In_698,In_1263);
nor U2366 (N_2366,In_57,In_2707);
nor U2367 (N_2367,In_1366,In_1663);
and U2368 (N_2368,In_2926,In_882);
nor U2369 (N_2369,In_702,In_167);
nor U2370 (N_2370,In_2818,In_1157);
or U2371 (N_2371,In_869,In_1534);
nand U2372 (N_2372,In_711,In_1347);
nand U2373 (N_2373,In_531,In_1654);
nand U2374 (N_2374,In_1004,In_518);
and U2375 (N_2375,In_305,In_1662);
and U2376 (N_2376,In_1919,In_968);
and U2377 (N_2377,In_2140,In_722);
or U2378 (N_2378,In_2455,In_1445);
xor U2379 (N_2379,In_2413,In_2077);
and U2380 (N_2380,In_628,In_175);
nor U2381 (N_2381,In_2672,In_598);
xor U2382 (N_2382,In_458,In_1256);
or U2383 (N_2383,In_2874,In_2233);
xor U2384 (N_2384,In_1766,In_1439);
xnor U2385 (N_2385,In_568,In_300);
xnor U2386 (N_2386,In_2510,In_702);
nand U2387 (N_2387,In_1871,In_2523);
or U2388 (N_2388,In_2448,In_528);
nand U2389 (N_2389,In_1343,In_2737);
xor U2390 (N_2390,In_2821,In_1640);
nor U2391 (N_2391,In_1766,In_1577);
nand U2392 (N_2392,In_676,In_1554);
or U2393 (N_2393,In_118,In_1204);
xnor U2394 (N_2394,In_1116,In_2795);
nor U2395 (N_2395,In_1376,In_1057);
nand U2396 (N_2396,In_1717,In_437);
nor U2397 (N_2397,In_210,In_1806);
nor U2398 (N_2398,In_1541,In_1117);
nor U2399 (N_2399,In_1695,In_94);
nand U2400 (N_2400,In_1500,In_2412);
xnor U2401 (N_2401,In_2892,In_1672);
nor U2402 (N_2402,In_993,In_2627);
or U2403 (N_2403,In_1960,In_305);
or U2404 (N_2404,In_621,In_1058);
or U2405 (N_2405,In_1893,In_309);
nor U2406 (N_2406,In_983,In_1511);
and U2407 (N_2407,In_439,In_170);
xor U2408 (N_2408,In_940,In_2388);
xor U2409 (N_2409,In_1713,In_609);
and U2410 (N_2410,In_2986,In_1415);
nand U2411 (N_2411,In_1041,In_2037);
or U2412 (N_2412,In_269,In_185);
nor U2413 (N_2413,In_897,In_950);
nor U2414 (N_2414,In_1873,In_201);
or U2415 (N_2415,In_691,In_1138);
nor U2416 (N_2416,In_366,In_1748);
nand U2417 (N_2417,In_2319,In_2845);
xor U2418 (N_2418,In_1707,In_494);
nor U2419 (N_2419,In_2884,In_656);
xor U2420 (N_2420,In_2024,In_2564);
and U2421 (N_2421,In_1946,In_689);
nand U2422 (N_2422,In_1839,In_1922);
nor U2423 (N_2423,In_2519,In_410);
nand U2424 (N_2424,In_1414,In_904);
nor U2425 (N_2425,In_2234,In_177);
and U2426 (N_2426,In_1950,In_2656);
or U2427 (N_2427,In_876,In_955);
nor U2428 (N_2428,In_233,In_1421);
and U2429 (N_2429,In_1407,In_2522);
xnor U2430 (N_2430,In_1840,In_267);
nor U2431 (N_2431,In_363,In_2123);
xor U2432 (N_2432,In_1223,In_2910);
nor U2433 (N_2433,In_685,In_481);
xor U2434 (N_2434,In_2430,In_1046);
nand U2435 (N_2435,In_254,In_1440);
nor U2436 (N_2436,In_1658,In_315);
nand U2437 (N_2437,In_1964,In_2162);
nor U2438 (N_2438,In_854,In_2681);
or U2439 (N_2439,In_550,In_964);
or U2440 (N_2440,In_767,In_336);
nor U2441 (N_2441,In_535,In_826);
or U2442 (N_2442,In_2656,In_1602);
and U2443 (N_2443,In_896,In_1789);
xor U2444 (N_2444,In_2158,In_1634);
or U2445 (N_2445,In_326,In_2306);
and U2446 (N_2446,In_595,In_2400);
nand U2447 (N_2447,In_2432,In_2318);
xnor U2448 (N_2448,In_1021,In_1577);
and U2449 (N_2449,In_564,In_949);
and U2450 (N_2450,In_2624,In_1343);
nand U2451 (N_2451,In_2841,In_1057);
and U2452 (N_2452,In_1070,In_512);
or U2453 (N_2453,In_1257,In_460);
or U2454 (N_2454,In_621,In_2989);
xnor U2455 (N_2455,In_2047,In_797);
xor U2456 (N_2456,In_1531,In_2802);
nand U2457 (N_2457,In_2525,In_93);
nand U2458 (N_2458,In_196,In_1634);
nor U2459 (N_2459,In_1047,In_1387);
or U2460 (N_2460,In_829,In_2581);
nand U2461 (N_2461,In_2414,In_720);
nand U2462 (N_2462,In_1930,In_2982);
nand U2463 (N_2463,In_122,In_2169);
or U2464 (N_2464,In_712,In_555);
nor U2465 (N_2465,In_433,In_1178);
xor U2466 (N_2466,In_2673,In_2873);
xnor U2467 (N_2467,In_1603,In_2804);
xor U2468 (N_2468,In_2921,In_1694);
or U2469 (N_2469,In_599,In_2299);
nand U2470 (N_2470,In_1160,In_2060);
or U2471 (N_2471,In_1520,In_159);
or U2472 (N_2472,In_1904,In_1411);
and U2473 (N_2473,In_2593,In_2114);
and U2474 (N_2474,In_1939,In_2118);
xor U2475 (N_2475,In_2062,In_1990);
xor U2476 (N_2476,In_2811,In_1779);
or U2477 (N_2477,In_856,In_796);
nor U2478 (N_2478,In_2859,In_1955);
nand U2479 (N_2479,In_2189,In_903);
nand U2480 (N_2480,In_529,In_1813);
and U2481 (N_2481,In_2242,In_953);
nand U2482 (N_2482,In_1893,In_216);
xor U2483 (N_2483,In_1027,In_2009);
or U2484 (N_2484,In_1653,In_2307);
and U2485 (N_2485,In_208,In_145);
and U2486 (N_2486,In_1238,In_670);
or U2487 (N_2487,In_2981,In_981);
nand U2488 (N_2488,In_590,In_328);
nor U2489 (N_2489,In_367,In_1187);
nor U2490 (N_2490,In_778,In_2716);
nor U2491 (N_2491,In_1498,In_373);
and U2492 (N_2492,In_1329,In_1676);
and U2493 (N_2493,In_486,In_860);
nor U2494 (N_2494,In_1645,In_1359);
or U2495 (N_2495,In_2106,In_2305);
nand U2496 (N_2496,In_2360,In_2642);
or U2497 (N_2497,In_1222,In_1209);
and U2498 (N_2498,In_309,In_2364);
xor U2499 (N_2499,In_2404,In_66);
nand U2500 (N_2500,In_398,In_2340);
or U2501 (N_2501,In_2721,In_19);
or U2502 (N_2502,In_382,In_803);
nand U2503 (N_2503,In_1808,In_2585);
nor U2504 (N_2504,In_281,In_1795);
xnor U2505 (N_2505,In_446,In_1669);
and U2506 (N_2506,In_2864,In_1724);
nor U2507 (N_2507,In_2134,In_922);
or U2508 (N_2508,In_1916,In_563);
or U2509 (N_2509,In_2075,In_1216);
xor U2510 (N_2510,In_2127,In_1827);
nor U2511 (N_2511,In_1222,In_632);
or U2512 (N_2512,In_307,In_1531);
nand U2513 (N_2513,In_1991,In_2667);
xor U2514 (N_2514,In_1510,In_1177);
nand U2515 (N_2515,In_1785,In_2399);
nor U2516 (N_2516,In_395,In_1604);
xor U2517 (N_2517,In_1390,In_476);
nor U2518 (N_2518,In_888,In_1510);
or U2519 (N_2519,In_672,In_656);
xor U2520 (N_2520,In_631,In_214);
nor U2521 (N_2521,In_2223,In_393);
and U2522 (N_2522,In_1087,In_118);
or U2523 (N_2523,In_1017,In_294);
nor U2524 (N_2524,In_1879,In_2864);
nor U2525 (N_2525,In_1588,In_2968);
or U2526 (N_2526,In_622,In_2848);
nor U2527 (N_2527,In_972,In_2841);
nor U2528 (N_2528,In_2479,In_1481);
xnor U2529 (N_2529,In_475,In_2413);
or U2530 (N_2530,In_1733,In_1432);
nand U2531 (N_2531,In_965,In_2388);
or U2532 (N_2532,In_275,In_2241);
nand U2533 (N_2533,In_619,In_1641);
or U2534 (N_2534,In_2451,In_1497);
or U2535 (N_2535,In_418,In_632);
or U2536 (N_2536,In_680,In_2122);
and U2537 (N_2537,In_2291,In_2459);
xnor U2538 (N_2538,In_1301,In_443);
and U2539 (N_2539,In_292,In_2475);
and U2540 (N_2540,In_571,In_812);
nand U2541 (N_2541,In_1857,In_1942);
or U2542 (N_2542,In_10,In_358);
or U2543 (N_2543,In_2277,In_2095);
xnor U2544 (N_2544,In_2569,In_2673);
xnor U2545 (N_2545,In_2581,In_123);
nand U2546 (N_2546,In_192,In_1409);
nor U2547 (N_2547,In_1916,In_2449);
and U2548 (N_2548,In_2685,In_2589);
or U2549 (N_2549,In_480,In_1426);
nor U2550 (N_2550,In_1906,In_1983);
xnor U2551 (N_2551,In_1312,In_1572);
and U2552 (N_2552,In_1767,In_2645);
and U2553 (N_2553,In_1894,In_1164);
nor U2554 (N_2554,In_1584,In_1096);
and U2555 (N_2555,In_1252,In_179);
nor U2556 (N_2556,In_1706,In_1690);
nor U2557 (N_2557,In_1509,In_357);
nor U2558 (N_2558,In_1248,In_517);
or U2559 (N_2559,In_623,In_1146);
and U2560 (N_2560,In_2531,In_2299);
nor U2561 (N_2561,In_688,In_2390);
xnor U2562 (N_2562,In_2207,In_1716);
xnor U2563 (N_2563,In_2755,In_666);
xnor U2564 (N_2564,In_2117,In_2137);
nand U2565 (N_2565,In_2579,In_716);
nor U2566 (N_2566,In_2724,In_1731);
nor U2567 (N_2567,In_2352,In_2048);
or U2568 (N_2568,In_2,In_1822);
or U2569 (N_2569,In_1520,In_2886);
or U2570 (N_2570,In_1530,In_437);
xor U2571 (N_2571,In_2318,In_1068);
or U2572 (N_2572,In_307,In_2607);
or U2573 (N_2573,In_1228,In_2012);
nor U2574 (N_2574,In_2554,In_2440);
nand U2575 (N_2575,In_2225,In_919);
nor U2576 (N_2576,In_103,In_2117);
xor U2577 (N_2577,In_2321,In_1016);
and U2578 (N_2578,In_2972,In_1287);
xor U2579 (N_2579,In_1484,In_2328);
nor U2580 (N_2580,In_1398,In_768);
and U2581 (N_2581,In_1390,In_2682);
xor U2582 (N_2582,In_309,In_1452);
and U2583 (N_2583,In_2376,In_518);
xnor U2584 (N_2584,In_2650,In_2583);
nand U2585 (N_2585,In_2401,In_2044);
nand U2586 (N_2586,In_251,In_191);
and U2587 (N_2587,In_1685,In_828);
xnor U2588 (N_2588,In_1205,In_423);
and U2589 (N_2589,In_2417,In_1121);
and U2590 (N_2590,In_542,In_2163);
nand U2591 (N_2591,In_2565,In_1567);
or U2592 (N_2592,In_2903,In_2811);
or U2593 (N_2593,In_2816,In_421);
nor U2594 (N_2594,In_2287,In_1175);
and U2595 (N_2595,In_2147,In_2672);
or U2596 (N_2596,In_991,In_1001);
nor U2597 (N_2597,In_1537,In_262);
xor U2598 (N_2598,In_893,In_2900);
nor U2599 (N_2599,In_2601,In_1066);
and U2600 (N_2600,In_1361,In_1197);
and U2601 (N_2601,In_612,In_1977);
and U2602 (N_2602,In_593,In_1143);
and U2603 (N_2603,In_2318,In_298);
xnor U2604 (N_2604,In_556,In_2491);
xnor U2605 (N_2605,In_2611,In_1120);
nor U2606 (N_2606,In_723,In_91);
and U2607 (N_2607,In_294,In_1462);
or U2608 (N_2608,In_1861,In_36);
nor U2609 (N_2609,In_2027,In_1510);
or U2610 (N_2610,In_2120,In_2119);
and U2611 (N_2611,In_774,In_2053);
and U2612 (N_2612,In_2443,In_2849);
nand U2613 (N_2613,In_2368,In_1963);
xor U2614 (N_2614,In_593,In_821);
nor U2615 (N_2615,In_2920,In_20);
or U2616 (N_2616,In_1987,In_2357);
xor U2617 (N_2617,In_1462,In_2381);
or U2618 (N_2618,In_625,In_232);
xor U2619 (N_2619,In_2051,In_1142);
and U2620 (N_2620,In_1532,In_2938);
nand U2621 (N_2621,In_2690,In_2932);
or U2622 (N_2622,In_1150,In_79);
and U2623 (N_2623,In_966,In_1500);
nor U2624 (N_2624,In_1140,In_1943);
nor U2625 (N_2625,In_2340,In_2841);
xnor U2626 (N_2626,In_1300,In_348);
xor U2627 (N_2627,In_32,In_1602);
or U2628 (N_2628,In_2089,In_2908);
and U2629 (N_2629,In_1245,In_2295);
nand U2630 (N_2630,In_1038,In_1142);
nand U2631 (N_2631,In_1895,In_1888);
nor U2632 (N_2632,In_2,In_1845);
xnor U2633 (N_2633,In_2531,In_1416);
or U2634 (N_2634,In_37,In_2824);
and U2635 (N_2635,In_2823,In_115);
and U2636 (N_2636,In_187,In_2413);
xor U2637 (N_2637,In_2663,In_1024);
nor U2638 (N_2638,In_2934,In_1291);
nand U2639 (N_2639,In_1786,In_2585);
or U2640 (N_2640,In_1792,In_1784);
or U2641 (N_2641,In_1555,In_1270);
nand U2642 (N_2642,In_2084,In_1635);
xnor U2643 (N_2643,In_763,In_652);
or U2644 (N_2644,In_592,In_2091);
nand U2645 (N_2645,In_641,In_465);
and U2646 (N_2646,In_2822,In_1471);
or U2647 (N_2647,In_1745,In_2735);
nand U2648 (N_2648,In_1866,In_310);
and U2649 (N_2649,In_2858,In_1289);
xnor U2650 (N_2650,In_1290,In_2926);
nand U2651 (N_2651,In_1711,In_2451);
nand U2652 (N_2652,In_2414,In_2272);
nor U2653 (N_2653,In_1304,In_1184);
nor U2654 (N_2654,In_412,In_1457);
or U2655 (N_2655,In_1250,In_2682);
and U2656 (N_2656,In_1393,In_1635);
and U2657 (N_2657,In_579,In_2298);
nand U2658 (N_2658,In_2085,In_2248);
nor U2659 (N_2659,In_82,In_1284);
nor U2660 (N_2660,In_1817,In_1865);
nand U2661 (N_2661,In_976,In_651);
and U2662 (N_2662,In_2669,In_495);
and U2663 (N_2663,In_975,In_664);
nor U2664 (N_2664,In_657,In_1239);
and U2665 (N_2665,In_1509,In_1963);
xnor U2666 (N_2666,In_1034,In_1463);
nand U2667 (N_2667,In_293,In_51);
nand U2668 (N_2668,In_599,In_1179);
or U2669 (N_2669,In_545,In_255);
nor U2670 (N_2670,In_818,In_2323);
and U2671 (N_2671,In_1055,In_1761);
xnor U2672 (N_2672,In_794,In_2715);
xnor U2673 (N_2673,In_536,In_1055);
nand U2674 (N_2674,In_902,In_2694);
nor U2675 (N_2675,In_2519,In_603);
nand U2676 (N_2676,In_1810,In_1994);
xnor U2677 (N_2677,In_937,In_1815);
or U2678 (N_2678,In_1859,In_1394);
nor U2679 (N_2679,In_2156,In_982);
nor U2680 (N_2680,In_268,In_1779);
and U2681 (N_2681,In_2944,In_1514);
nand U2682 (N_2682,In_700,In_83);
xor U2683 (N_2683,In_1191,In_1354);
nand U2684 (N_2684,In_2260,In_783);
and U2685 (N_2685,In_2135,In_402);
nor U2686 (N_2686,In_1614,In_2324);
and U2687 (N_2687,In_821,In_1022);
xor U2688 (N_2688,In_289,In_1204);
nor U2689 (N_2689,In_2561,In_1403);
and U2690 (N_2690,In_1004,In_1395);
or U2691 (N_2691,In_1163,In_2993);
nor U2692 (N_2692,In_785,In_1978);
nor U2693 (N_2693,In_2872,In_223);
nor U2694 (N_2694,In_2070,In_40);
nand U2695 (N_2695,In_1024,In_190);
nor U2696 (N_2696,In_1825,In_863);
or U2697 (N_2697,In_1598,In_1885);
or U2698 (N_2698,In_1225,In_1955);
xnor U2699 (N_2699,In_2198,In_224);
xnor U2700 (N_2700,In_1261,In_358);
or U2701 (N_2701,In_1355,In_2924);
nor U2702 (N_2702,In_1512,In_1158);
or U2703 (N_2703,In_412,In_2547);
nand U2704 (N_2704,In_2848,In_2116);
or U2705 (N_2705,In_1923,In_2439);
xor U2706 (N_2706,In_2521,In_1101);
nand U2707 (N_2707,In_159,In_1845);
xor U2708 (N_2708,In_1396,In_2905);
xor U2709 (N_2709,In_187,In_2065);
or U2710 (N_2710,In_2925,In_2889);
and U2711 (N_2711,In_2287,In_1684);
xor U2712 (N_2712,In_1417,In_2805);
and U2713 (N_2713,In_814,In_2205);
and U2714 (N_2714,In_1594,In_744);
xor U2715 (N_2715,In_1056,In_933);
and U2716 (N_2716,In_1075,In_670);
xor U2717 (N_2717,In_1036,In_1300);
and U2718 (N_2718,In_1915,In_1748);
and U2719 (N_2719,In_1135,In_1377);
nor U2720 (N_2720,In_2835,In_1665);
or U2721 (N_2721,In_616,In_1944);
and U2722 (N_2722,In_889,In_1859);
xnor U2723 (N_2723,In_209,In_1580);
and U2724 (N_2724,In_1252,In_174);
nand U2725 (N_2725,In_2263,In_1256);
and U2726 (N_2726,In_1551,In_1919);
or U2727 (N_2727,In_2216,In_1072);
xor U2728 (N_2728,In_96,In_2929);
and U2729 (N_2729,In_2471,In_1555);
or U2730 (N_2730,In_2058,In_289);
nor U2731 (N_2731,In_721,In_1861);
or U2732 (N_2732,In_659,In_2838);
xnor U2733 (N_2733,In_2019,In_587);
or U2734 (N_2734,In_1648,In_2063);
nand U2735 (N_2735,In_2834,In_2868);
nor U2736 (N_2736,In_864,In_1444);
xnor U2737 (N_2737,In_461,In_781);
nand U2738 (N_2738,In_2384,In_1378);
nor U2739 (N_2739,In_2452,In_144);
or U2740 (N_2740,In_872,In_2849);
nand U2741 (N_2741,In_348,In_569);
or U2742 (N_2742,In_61,In_202);
xnor U2743 (N_2743,In_2346,In_493);
nor U2744 (N_2744,In_2756,In_2207);
nor U2745 (N_2745,In_2322,In_2214);
or U2746 (N_2746,In_1871,In_339);
nor U2747 (N_2747,In_624,In_760);
and U2748 (N_2748,In_1313,In_2614);
nand U2749 (N_2749,In_109,In_1279);
nand U2750 (N_2750,In_540,In_2981);
and U2751 (N_2751,In_2994,In_1808);
nor U2752 (N_2752,In_1622,In_2754);
and U2753 (N_2753,In_80,In_2596);
and U2754 (N_2754,In_1773,In_410);
nand U2755 (N_2755,In_1295,In_1797);
nand U2756 (N_2756,In_1232,In_585);
xnor U2757 (N_2757,In_1792,In_150);
xor U2758 (N_2758,In_2304,In_1319);
nand U2759 (N_2759,In_2413,In_1942);
nor U2760 (N_2760,In_7,In_230);
xor U2761 (N_2761,In_236,In_1014);
and U2762 (N_2762,In_1220,In_1662);
or U2763 (N_2763,In_1064,In_840);
nand U2764 (N_2764,In_1914,In_2661);
and U2765 (N_2765,In_1346,In_475);
nor U2766 (N_2766,In_1277,In_941);
or U2767 (N_2767,In_1583,In_456);
nand U2768 (N_2768,In_2717,In_727);
nor U2769 (N_2769,In_1592,In_1679);
nand U2770 (N_2770,In_2523,In_2775);
nor U2771 (N_2771,In_1992,In_9);
nor U2772 (N_2772,In_508,In_2535);
and U2773 (N_2773,In_1398,In_242);
or U2774 (N_2774,In_587,In_2498);
nor U2775 (N_2775,In_2284,In_1085);
nand U2776 (N_2776,In_897,In_177);
nand U2777 (N_2777,In_304,In_427);
nor U2778 (N_2778,In_1540,In_1856);
or U2779 (N_2779,In_1618,In_2345);
or U2780 (N_2780,In_1189,In_354);
xor U2781 (N_2781,In_954,In_1338);
nor U2782 (N_2782,In_1503,In_1453);
nor U2783 (N_2783,In_1999,In_2338);
and U2784 (N_2784,In_2259,In_769);
and U2785 (N_2785,In_62,In_1309);
nand U2786 (N_2786,In_1779,In_2519);
nand U2787 (N_2787,In_2634,In_1919);
nor U2788 (N_2788,In_2866,In_1755);
or U2789 (N_2789,In_610,In_570);
or U2790 (N_2790,In_2433,In_2881);
or U2791 (N_2791,In_16,In_431);
xor U2792 (N_2792,In_464,In_2379);
nor U2793 (N_2793,In_2691,In_2872);
nor U2794 (N_2794,In_779,In_405);
and U2795 (N_2795,In_2278,In_2899);
xor U2796 (N_2796,In_2406,In_2009);
xnor U2797 (N_2797,In_1581,In_330);
or U2798 (N_2798,In_1713,In_86);
or U2799 (N_2799,In_377,In_2216);
nand U2800 (N_2800,In_397,In_2759);
nand U2801 (N_2801,In_1397,In_265);
xnor U2802 (N_2802,In_1026,In_2558);
xor U2803 (N_2803,In_1238,In_850);
nor U2804 (N_2804,In_2049,In_594);
and U2805 (N_2805,In_1369,In_2549);
or U2806 (N_2806,In_2555,In_1487);
nand U2807 (N_2807,In_694,In_1080);
nand U2808 (N_2808,In_603,In_2506);
nand U2809 (N_2809,In_2324,In_1981);
nand U2810 (N_2810,In_1644,In_1568);
or U2811 (N_2811,In_2630,In_839);
nor U2812 (N_2812,In_492,In_2591);
and U2813 (N_2813,In_340,In_2778);
nand U2814 (N_2814,In_1179,In_1086);
xnor U2815 (N_2815,In_1067,In_2562);
xnor U2816 (N_2816,In_2131,In_2828);
or U2817 (N_2817,In_1388,In_5);
or U2818 (N_2818,In_2260,In_1506);
and U2819 (N_2819,In_2890,In_898);
xnor U2820 (N_2820,In_1725,In_2207);
xor U2821 (N_2821,In_2965,In_1127);
or U2822 (N_2822,In_2321,In_1069);
nor U2823 (N_2823,In_878,In_379);
and U2824 (N_2824,In_622,In_1416);
nor U2825 (N_2825,In_1059,In_1603);
or U2826 (N_2826,In_631,In_2050);
xor U2827 (N_2827,In_557,In_388);
or U2828 (N_2828,In_1704,In_2983);
nand U2829 (N_2829,In_2737,In_2247);
xor U2830 (N_2830,In_471,In_1320);
nand U2831 (N_2831,In_1830,In_767);
and U2832 (N_2832,In_1475,In_2128);
xnor U2833 (N_2833,In_190,In_2817);
or U2834 (N_2834,In_1791,In_669);
nand U2835 (N_2835,In_163,In_2409);
nand U2836 (N_2836,In_2061,In_1208);
nand U2837 (N_2837,In_276,In_1135);
nand U2838 (N_2838,In_2768,In_355);
and U2839 (N_2839,In_994,In_1271);
and U2840 (N_2840,In_1570,In_1069);
nor U2841 (N_2841,In_1990,In_2884);
and U2842 (N_2842,In_2571,In_2223);
nand U2843 (N_2843,In_642,In_2287);
xnor U2844 (N_2844,In_421,In_668);
nor U2845 (N_2845,In_2042,In_1135);
nand U2846 (N_2846,In_2631,In_843);
xor U2847 (N_2847,In_2251,In_2299);
or U2848 (N_2848,In_819,In_1744);
and U2849 (N_2849,In_706,In_2898);
nand U2850 (N_2850,In_2844,In_1009);
and U2851 (N_2851,In_41,In_1406);
xor U2852 (N_2852,In_2933,In_1575);
and U2853 (N_2853,In_2005,In_874);
and U2854 (N_2854,In_2617,In_684);
nand U2855 (N_2855,In_2858,In_1443);
nand U2856 (N_2856,In_2917,In_776);
xor U2857 (N_2857,In_222,In_2839);
nor U2858 (N_2858,In_2530,In_995);
nor U2859 (N_2859,In_1339,In_2706);
nor U2860 (N_2860,In_1262,In_485);
or U2861 (N_2861,In_1744,In_1331);
nor U2862 (N_2862,In_2626,In_2133);
nor U2863 (N_2863,In_79,In_2732);
nand U2864 (N_2864,In_522,In_538);
or U2865 (N_2865,In_2298,In_869);
or U2866 (N_2866,In_234,In_2127);
or U2867 (N_2867,In_2947,In_901);
and U2868 (N_2868,In_93,In_2686);
nand U2869 (N_2869,In_1063,In_1042);
and U2870 (N_2870,In_2730,In_2471);
and U2871 (N_2871,In_297,In_977);
xnor U2872 (N_2872,In_2206,In_900);
nor U2873 (N_2873,In_88,In_1005);
xnor U2874 (N_2874,In_2506,In_2044);
nor U2875 (N_2875,In_2097,In_657);
nor U2876 (N_2876,In_1305,In_1016);
nor U2877 (N_2877,In_2032,In_368);
xor U2878 (N_2878,In_2254,In_1124);
nand U2879 (N_2879,In_643,In_982);
nor U2880 (N_2880,In_2688,In_1562);
or U2881 (N_2881,In_1891,In_97);
nand U2882 (N_2882,In_55,In_1250);
xnor U2883 (N_2883,In_769,In_2361);
nand U2884 (N_2884,In_1853,In_1314);
or U2885 (N_2885,In_1538,In_1764);
xor U2886 (N_2886,In_1357,In_428);
nor U2887 (N_2887,In_2200,In_898);
xnor U2888 (N_2888,In_477,In_1281);
nor U2889 (N_2889,In_2828,In_1132);
xor U2890 (N_2890,In_552,In_833);
and U2891 (N_2891,In_379,In_834);
xnor U2892 (N_2892,In_2594,In_926);
nor U2893 (N_2893,In_2435,In_2237);
xor U2894 (N_2894,In_2777,In_2998);
xor U2895 (N_2895,In_473,In_1704);
or U2896 (N_2896,In_1360,In_1908);
xnor U2897 (N_2897,In_2784,In_1955);
nor U2898 (N_2898,In_430,In_2235);
xor U2899 (N_2899,In_1767,In_361);
or U2900 (N_2900,In_2299,In_426);
or U2901 (N_2901,In_81,In_697);
and U2902 (N_2902,In_297,In_2681);
and U2903 (N_2903,In_1265,In_2629);
nand U2904 (N_2904,In_1210,In_213);
and U2905 (N_2905,In_1872,In_2455);
and U2906 (N_2906,In_456,In_94);
or U2907 (N_2907,In_1436,In_2107);
xor U2908 (N_2908,In_660,In_366);
and U2909 (N_2909,In_878,In_1731);
nor U2910 (N_2910,In_2459,In_986);
and U2911 (N_2911,In_2283,In_849);
or U2912 (N_2912,In_631,In_338);
nand U2913 (N_2913,In_1177,In_565);
or U2914 (N_2914,In_102,In_788);
nor U2915 (N_2915,In_535,In_2284);
and U2916 (N_2916,In_2393,In_2301);
xnor U2917 (N_2917,In_1068,In_2497);
nand U2918 (N_2918,In_226,In_2462);
nor U2919 (N_2919,In_380,In_1440);
nand U2920 (N_2920,In_2141,In_1655);
nand U2921 (N_2921,In_2922,In_1530);
nand U2922 (N_2922,In_1227,In_650);
nor U2923 (N_2923,In_749,In_1162);
or U2924 (N_2924,In_2967,In_1995);
nand U2925 (N_2925,In_1367,In_2800);
nand U2926 (N_2926,In_485,In_1268);
or U2927 (N_2927,In_901,In_1480);
nand U2928 (N_2928,In_2259,In_1852);
xor U2929 (N_2929,In_517,In_2756);
and U2930 (N_2930,In_413,In_1355);
nand U2931 (N_2931,In_1468,In_949);
or U2932 (N_2932,In_1555,In_1790);
and U2933 (N_2933,In_2153,In_1973);
nor U2934 (N_2934,In_1943,In_1176);
nor U2935 (N_2935,In_346,In_2499);
xor U2936 (N_2936,In_2177,In_2775);
nor U2937 (N_2937,In_936,In_775);
xor U2938 (N_2938,In_1244,In_1178);
nand U2939 (N_2939,In_245,In_1472);
nand U2940 (N_2940,In_2207,In_1238);
and U2941 (N_2941,In_2218,In_415);
xnor U2942 (N_2942,In_1617,In_1184);
nand U2943 (N_2943,In_503,In_2682);
and U2944 (N_2944,In_2732,In_2655);
xor U2945 (N_2945,In_2071,In_2951);
and U2946 (N_2946,In_1482,In_1891);
and U2947 (N_2947,In_1319,In_676);
and U2948 (N_2948,In_2346,In_1412);
nand U2949 (N_2949,In_521,In_2358);
or U2950 (N_2950,In_583,In_374);
or U2951 (N_2951,In_1675,In_405);
nor U2952 (N_2952,In_2231,In_969);
nand U2953 (N_2953,In_2729,In_1401);
and U2954 (N_2954,In_1791,In_2735);
or U2955 (N_2955,In_340,In_2510);
nand U2956 (N_2956,In_701,In_2775);
xor U2957 (N_2957,In_1325,In_2873);
xnor U2958 (N_2958,In_769,In_1012);
nand U2959 (N_2959,In_155,In_423);
or U2960 (N_2960,In_2615,In_827);
nor U2961 (N_2961,In_1076,In_573);
xnor U2962 (N_2962,In_1560,In_2308);
nand U2963 (N_2963,In_733,In_2083);
nand U2964 (N_2964,In_747,In_688);
nor U2965 (N_2965,In_959,In_2300);
nand U2966 (N_2966,In_894,In_1705);
or U2967 (N_2967,In_255,In_2247);
nand U2968 (N_2968,In_189,In_2965);
nand U2969 (N_2969,In_1460,In_2047);
or U2970 (N_2970,In_1865,In_1694);
nor U2971 (N_2971,In_1946,In_1336);
or U2972 (N_2972,In_644,In_511);
or U2973 (N_2973,In_236,In_1129);
nand U2974 (N_2974,In_2292,In_1780);
xnor U2975 (N_2975,In_1789,In_1564);
nor U2976 (N_2976,In_1076,In_249);
nand U2977 (N_2977,In_2609,In_494);
and U2978 (N_2978,In_2655,In_771);
and U2979 (N_2979,In_1956,In_1196);
and U2980 (N_2980,In_1506,In_643);
nor U2981 (N_2981,In_123,In_217);
xnor U2982 (N_2982,In_2414,In_235);
and U2983 (N_2983,In_2227,In_653);
xor U2984 (N_2984,In_1386,In_167);
and U2985 (N_2985,In_2679,In_1578);
xnor U2986 (N_2986,In_611,In_2155);
and U2987 (N_2987,In_133,In_546);
nor U2988 (N_2988,In_2057,In_564);
nor U2989 (N_2989,In_1454,In_2071);
or U2990 (N_2990,In_754,In_2853);
nor U2991 (N_2991,In_33,In_1995);
and U2992 (N_2992,In_2973,In_1466);
nor U2993 (N_2993,In_592,In_274);
xnor U2994 (N_2994,In_2429,In_2188);
xnor U2995 (N_2995,In_294,In_854);
nand U2996 (N_2996,In_1562,In_2387);
nor U2997 (N_2997,In_922,In_392);
and U2998 (N_2998,In_2611,In_2849);
xor U2999 (N_2999,In_144,In_513);
nand U3000 (N_3000,N_1479,N_655);
or U3001 (N_3001,N_1645,N_638);
and U3002 (N_3002,N_2599,N_1572);
or U3003 (N_3003,N_150,N_1627);
xor U3004 (N_3004,N_304,N_1215);
and U3005 (N_3005,N_2681,N_1948);
xnor U3006 (N_3006,N_1502,N_2219);
xnor U3007 (N_3007,N_2875,N_2254);
xnor U3008 (N_3008,N_668,N_1469);
nand U3009 (N_3009,N_2364,N_2582);
xnor U3010 (N_3010,N_2863,N_2506);
nor U3011 (N_3011,N_1571,N_1087);
and U3012 (N_3012,N_1112,N_1935);
and U3013 (N_3013,N_2730,N_501);
xor U3014 (N_3014,N_2542,N_403);
or U3015 (N_3015,N_2787,N_2620);
xnor U3016 (N_3016,N_1093,N_742);
or U3017 (N_3017,N_473,N_2299);
nand U3018 (N_3018,N_2782,N_2492);
xor U3019 (N_3019,N_857,N_508);
and U3020 (N_3020,N_359,N_335);
and U3021 (N_3021,N_2615,N_2400);
xnor U3022 (N_3022,N_458,N_2797);
nor U3023 (N_3023,N_1091,N_1618);
xor U3024 (N_3024,N_842,N_2404);
xnor U3025 (N_3025,N_1314,N_551);
and U3026 (N_3026,N_214,N_2039);
nand U3027 (N_3027,N_783,N_456);
and U3028 (N_3028,N_858,N_2871);
nor U3029 (N_3029,N_754,N_2121);
or U3030 (N_3030,N_591,N_2712);
or U3031 (N_3031,N_432,N_1450);
xnor U3032 (N_3032,N_2849,N_980);
or U3033 (N_3033,N_2301,N_2557);
or U3034 (N_3034,N_496,N_429);
or U3035 (N_3035,N_695,N_1515);
or U3036 (N_3036,N_2067,N_27);
nor U3037 (N_3037,N_2230,N_1713);
nor U3038 (N_3038,N_992,N_1857);
and U3039 (N_3039,N_1794,N_6);
or U3040 (N_3040,N_131,N_60);
xnor U3041 (N_3041,N_2468,N_0);
nand U3042 (N_3042,N_128,N_2987);
xor U3043 (N_3043,N_2256,N_2840);
nand U3044 (N_3044,N_1675,N_1991);
nand U3045 (N_3045,N_1227,N_2489);
and U3046 (N_3046,N_1305,N_1108);
nor U3047 (N_3047,N_2537,N_2719);
and U3048 (N_3048,N_469,N_1357);
nor U3049 (N_3049,N_2372,N_2761);
or U3050 (N_3050,N_2523,N_190);
nor U3051 (N_3051,N_1149,N_1072);
nand U3052 (N_3052,N_868,N_662);
nand U3053 (N_3053,N_704,N_1252);
or U3054 (N_3054,N_1448,N_443);
and U3055 (N_3055,N_2798,N_1187);
xor U3056 (N_3056,N_2956,N_1975);
xnor U3057 (N_3057,N_2918,N_714);
nand U3058 (N_3058,N_622,N_149);
and U3059 (N_3059,N_1143,N_2041);
nand U3060 (N_3060,N_520,N_590);
and U3061 (N_3061,N_1811,N_899);
or U3062 (N_3062,N_570,N_2643);
nor U3063 (N_3063,N_360,N_1716);
nand U3064 (N_3064,N_1323,N_995);
nand U3065 (N_3065,N_2210,N_987);
nand U3066 (N_3066,N_1589,N_1233);
nor U3067 (N_3067,N_307,N_1429);
and U3068 (N_3068,N_2232,N_325);
and U3069 (N_3069,N_1275,N_2661);
or U3070 (N_3070,N_2988,N_2774);
or U3071 (N_3071,N_1582,N_2068);
nand U3072 (N_3072,N_1724,N_294);
or U3073 (N_3073,N_2870,N_1123);
nand U3074 (N_3074,N_2520,N_2541);
nand U3075 (N_3075,N_1082,N_2085);
nor U3076 (N_3076,N_1000,N_2486);
nand U3077 (N_3077,N_785,N_2517);
xnor U3078 (N_3078,N_510,N_2650);
or U3079 (N_3079,N_2487,N_1714);
nor U3080 (N_3080,N_2111,N_1613);
xnor U3081 (N_3081,N_635,N_971);
nor U3082 (N_3082,N_1525,N_2287);
nand U3083 (N_3083,N_465,N_1438);
and U3084 (N_3084,N_12,N_2737);
nor U3085 (N_3085,N_1051,N_828);
and U3086 (N_3086,N_804,N_2385);
nand U3087 (N_3087,N_2073,N_2954);
nand U3088 (N_3088,N_2663,N_641);
or U3089 (N_3089,N_1827,N_1818);
or U3090 (N_3090,N_2285,N_1245);
nand U3091 (N_3091,N_1770,N_1989);
nor U3092 (N_3092,N_1085,N_2509);
nand U3093 (N_3093,N_1126,N_1228);
nand U3094 (N_3094,N_880,N_422);
xnor U3095 (N_3095,N_2963,N_1522);
or U3096 (N_3096,N_2061,N_356);
and U3097 (N_3097,N_2654,N_724);
nor U3098 (N_3098,N_2595,N_1241);
nor U3099 (N_3099,N_2091,N_972);
and U3100 (N_3100,N_2181,N_395);
and U3101 (N_3101,N_2384,N_49);
xor U3102 (N_3102,N_1973,N_251);
nand U3103 (N_3103,N_546,N_556);
nor U3104 (N_3104,N_203,N_603);
nand U3105 (N_3105,N_2893,N_2311);
nor U3106 (N_3106,N_2501,N_2884);
xnor U3107 (N_3107,N_2156,N_2493);
and U3108 (N_3108,N_2469,N_763);
and U3109 (N_3109,N_1746,N_2142);
and U3110 (N_3110,N_1886,N_71);
and U3111 (N_3111,N_847,N_2152);
or U3112 (N_3112,N_1887,N_290);
xnor U3113 (N_3113,N_109,N_1505);
nand U3114 (N_3114,N_262,N_2332);
and U3115 (N_3115,N_2577,N_1136);
nor U3116 (N_3116,N_1045,N_74);
and U3117 (N_3117,N_1184,N_1974);
and U3118 (N_3118,N_770,N_2899);
or U3119 (N_3119,N_2170,N_2211);
nor U3120 (N_3120,N_2403,N_287);
or U3121 (N_3121,N_1608,N_2320);
and U3122 (N_3122,N_2164,N_1862);
nor U3123 (N_3123,N_1725,N_888);
and U3124 (N_3124,N_861,N_379);
or U3125 (N_3125,N_2873,N_891);
xnor U3126 (N_3126,N_2458,N_2155);
nor U3127 (N_3127,N_2692,N_1114);
nand U3128 (N_3128,N_2622,N_909);
nand U3129 (N_3129,N_253,N_2020);
nor U3130 (N_3130,N_1619,N_1993);
or U3131 (N_3131,N_2978,N_2017);
and U3132 (N_3132,N_2282,N_51);
xnor U3133 (N_3133,N_790,N_2079);
and U3134 (N_3134,N_1634,N_2904);
and U3135 (N_3135,N_924,N_560);
nand U3136 (N_3136,N_1248,N_1517);
nand U3137 (N_3137,N_536,N_2706);
xor U3138 (N_3138,N_2046,N_1674);
and U3139 (N_3139,N_1262,N_1617);
nand U3140 (N_3140,N_2652,N_2329);
nand U3141 (N_3141,N_478,N_1346);
or U3142 (N_3142,N_755,N_141);
xnor U3143 (N_3143,N_1990,N_1542);
nor U3144 (N_3144,N_2605,N_2066);
and U3145 (N_3145,N_1364,N_1162);
nor U3146 (N_3146,N_597,N_1445);
nand U3147 (N_3147,N_838,N_2209);
nor U3148 (N_3148,N_2445,N_1374);
nand U3149 (N_3149,N_1380,N_1351);
xnor U3150 (N_3150,N_1454,N_2003);
nor U3151 (N_3151,N_1947,N_910);
nand U3152 (N_3152,N_2388,N_1417);
nand U3153 (N_3153,N_563,N_1804);
nor U3154 (N_3154,N_2080,N_640);
nand U3155 (N_3155,N_2726,N_985);
xor U3156 (N_3156,N_2511,N_966);
and U3157 (N_3157,N_1319,N_1047);
or U3158 (N_3158,N_1740,N_2000);
nand U3159 (N_3159,N_548,N_174);
nor U3160 (N_3160,N_978,N_2810);
nand U3161 (N_3161,N_1992,N_1411);
or U3162 (N_3162,N_447,N_2392);
or U3163 (N_3163,N_1834,N_1906);
or U3164 (N_3164,N_2391,N_802);
xnor U3165 (N_3165,N_633,N_129);
xor U3166 (N_3166,N_1127,N_207);
or U3167 (N_3167,N_2901,N_140);
and U3168 (N_3168,N_20,N_352);
xnor U3169 (N_3169,N_2473,N_2122);
and U3170 (N_3170,N_1686,N_368);
and U3171 (N_3171,N_397,N_2860);
xor U3172 (N_3172,N_948,N_1977);
nand U3173 (N_3173,N_62,N_731);
or U3174 (N_3174,N_487,N_459);
xnor U3175 (N_3175,N_2109,N_2594);
nand U3176 (N_3176,N_1927,N_121);
nor U3177 (N_3177,N_2677,N_2762);
xor U3178 (N_3178,N_280,N_153);
and U3179 (N_3179,N_446,N_766);
xnor U3180 (N_3180,N_2365,N_1905);
and U3181 (N_3181,N_2946,N_2767);
and U3182 (N_3182,N_1587,N_2854);
and U3183 (N_3183,N_753,N_521);
nand U3184 (N_3184,N_2895,N_1223);
xnor U3185 (N_3185,N_35,N_2187);
nand U3186 (N_3186,N_1343,N_2488);
xnor U3187 (N_3187,N_1508,N_2283);
and U3188 (N_3188,N_1928,N_1509);
nand U3189 (N_3189,N_2932,N_1600);
and U3190 (N_3190,N_968,N_2031);
nor U3191 (N_3191,N_2081,N_1764);
or U3192 (N_3192,N_665,N_2915);
nand U3193 (N_3193,N_1148,N_86);
nand U3194 (N_3194,N_1877,N_120);
and U3195 (N_3195,N_954,N_2619);
and U3196 (N_3196,N_1579,N_1470);
and U3197 (N_3197,N_1658,N_215);
xor U3198 (N_3198,N_2834,N_1446);
and U3199 (N_3199,N_848,N_2830);
and U3200 (N_3200,N_40,N_1753);
or U3201 (N_3201,N_730,N_2218);
or U3202 (N_3202,N_2551,N_2885);
or U3203 (N_3203,N_2411,N_2442);
or U3204 (N_3204,N_498,N_644);
xor U3205 (N_3205,N_2981,N_338);
xnor U3206 (N_3206,N_415,N_1043);
and U3207 (N_3207,N_1427,N_2953);
or U3208 (N_3208,N_1595,N_751);
xnor U3209 (N_3209,N_2215,N_407);
xnor U3210 (N_3210,N_2564,N_2147);
or U3211 (N_3211,N_1354,N_2739);
nand U3212 (N_3212,N_442,N_1551);
and U3213 (N_3213,N_1489,N_1667);
or U3214 (N_3214,N_2010,N_2379);
xnor U3215 (N_3215,N_2515,N_1147);
and U3216 (N_3216,N_1003,N_2554);
or U3217 (N_3217,N_125,N_1745);
xnor U3218 (N_3218,N_1382,N_1699);
or U3219 (N_3219,N_1480,N_2641);
nor U3220 (N_3220,N_56,N_1702);
xnor U3221 (N_3221,N_339,N_1964);
nor U3222 (N_3222,N_834,N_2402);
nand U3223 (N_3223,N_2876,N_960);
or U3224 (N_3224,N_779,N_2927);
nor U3225 (N_3225,N_1520,N_2393);
or U3226 (N_3226,N_2573,N_305);
or U3227 (N_3227,N_2967,N_1695);
nor U3228 (N_3228,N_855,N_2322);
xor U3229 (N_3229,N_1757,N_2255);
nor U3230 (N_3230,N_669,N_1844);
xor U3231 (N_3231,N_613,N_630);
or U3232 (N_3232,N_1513,N_286);
nor U3233 (N_3233,N_38,N_1337);
or U3234 (N_3234,N_543,N_2984);
and U3235 (N_3235,N_470,N_2628);
and U3236 (N_3236,N_390,N_1036);
and U3237 (N_3237,N_2248,N_1883);
xnor U3238 (N_3238,N_2037,N_468);
and U3239 (N_3239,N_2169,N_2738);
nand U3240 (N_3240,N_1461,N_2314);
or U3241 (N_3241,N_1128,N_1316);
nand U3242 (N_3242,N_1939,N_2077);
nor U3243 (N_3243,N_358,N_2128);
or U3244 (N_3244,N_132,N_593);
nand U3245 (N_3245,N_2916,N_2349);
nand U3246 (N_3246,N_1097,N_2001);
and U3247 (N_3247,N_2366,N_1268);
nand U3248 (N_3248,N_488,N_371);
nand U3249 (N_3249,N_1599,N_612);
or U3250 (N_3250,N_1644,N_2114);
nand U3251 (N_3251,N_659,N_2363);
nand U3252 (N_3252,N_944,N_2262);
nor U3253 (N_3253,N_1192,N_1370);
and U3254 (N_3254,N_2693,N_2423);
and U3255 (N_3255,N_1201,N_1064);
xnor U3256 (N_3256,N_68,N_1604);
nor U3257 (N_3257,N_2380,N_1621);
nor U3258 (N_3258,N_990,N_1235);
xor U3259 (N_3259,N_1070,N_2013);
nand U3260 (N_3260,N_2191,N_2116);
xor U3261 (N_3261,N_2846,N_1829);
or U3262 (N_3262,N_2043,N_2653);
or U3263 (N_3263,N_2257,N_2752);
nand U3264 (N_3264,N_78,N_1996);
nor U3265 (N_3265,N_542,N_1612);
nand U3266 (N_3266,N_2133,N_418);
nor U3267 (N_3267,N_1751,N_673);
xnor U3268 (N_3268,N_565,N_2118);
xor U3269 (N_3269,N_1237,N_866);
and U3270 (N_3270,N_1843,N_816);
xor U3271 (N_3271,N_1656,N_2685);
and U3272 (N_3272,N_2408,N_1222);
nand U3273 (N_3273,N_2788,N_994);
xor U3274 (N_3274,N_524,N_1498);
nand U3275 (N_3275,N_2504,N_2836);
and U3276 (N_3276,N_2317,N_1298);
xor U3277 (N_3277,N_620,N_93);
nand U3278 (N_3278,N_2913,N_696);
nor U3279 (N_3279,N_1308,N_237);
and U3280 (N_3280,N_261,N_555);
or U3281 (N_3281,N_88,N_1435);
and U3282 (N_3282,N_2055,N_1849);
or U3283 (N_3283,N_2102,N_768);
nand U3284 (N_3284,N_2740,N_298);
xnor U3285 (N_3285,N_1913,N_2805);
nand U3286 (N_3286,N_2676,N_220);
xor U3287 (N_3287,N_119,N_1892);
nand U3288 (N_3288,N_1332,N_466);
and U3289 (N_3289,N_1179,N_2025);
nor U3290 (N_3290,N_2202,N_1917);
and U3291 (N_3291,N_2397,N_1637);
or U3292 (N_3292,N_1118,N_1543);
and U3293 (N_3293,N_1163,N_276);
or U3294 (N_3294,N_1688,N_2153);
or U3295 (N_3295,N_135,N_344);
nand U3296 (N_3296,N_1265,N_272);
nor U3297 (N_3297,N_1651,N_747);
and U3298 (N_3298,N_1146,N_1335);
or U3299 (N_3299,N_1856,N_181);
nor U3300 (N_3300,N_894,N_202);
xor U3301 (N_3301,N_2223,N_491);
and U3302 (N_3302,N_647,N_2290);
nand U3303 (N_3303,N_1558,N_719);
nand U3304 (N_3304,N_226,N_2867);
nand U3305 (N_3305,N_1959,N_1153);
xnor U3306 (N_3306,N_1793,N_1115);
nand U3307 (N_3307,N_2450,N_1698);
xor U3308 (N_3308,N_2375,N_873);
nand U3309 (N_3309,N_2950,N_2713);
and U3310 (N_3310,N_2640,N_284);
nand U3311 (N_3311,N_2896,N_1870);
xor U3312 (N_3312,N_2453,N_605);
nor U3313 (N_3313,N_330,N_1561);
xor U3314 (N_3314,N_1073,N_2226);
nor U3315 (N_3315,N_1904,N_2703);
nor U3316 (N_3316,N_239,N_917);
and U3317 (N_3317,N_2186,N_584);
nand U3318 (N_3318,N_1533,N_1309);
and U3319 (N_3319,N_331,N_1383);
nor U3320 (N_3320,N_2755,N_1413);
and U3321 (N_3321,N_2057,N_3);
and U3322 (N_3322,N_2278,N_378);
and U3323 (N_3323,N_2498,N_2044);
xor U3324 (N_3324,N_1664,N_2361);
xor U3325 (N_3325,N_1208,N_1061);
nor U3326 (N_3326,N_2416,N_186);
and U3327 (N_3327,N_2618,N_621);
nor U3328 (N_3328,N_1481,N_127);
and U3329 (N_3329,N_2502,N_2221);
or U3330 (N_3330,N_47,N_534);
xor U3331 (N_3331,N_1581,N_176);
xor U3332 (N_3332,N_955,N_831);
or U3333 (N_3333,N_2024,N_1806);
xor U3334 (N_3334,N_2945,N_1647);
nor U3335 (N_3335,N_2161,N_1919);
and U3336 (N_3336,N_625,N_1726);
and U3337 (N_3337,N_1689,N_2818);
or U3338 (N_3338,N_1573,N_1069);
and U3339 (N_3339,N_2724,N_1569);
nand U3340 (N_3340,N_1788,N_221);
or U3341 (N_3341,N_2892,N_2697);
and U3342 (N_3342,N_1577,N_16);
nand U3343 (N_3343,N_380,N_818);
and U3344 (N_3344,N_2548,N_1111);
nor U3345 (N_3345,N_2746,N_1117);
nor U3346 (N_3346,N_2700,N_2015);
nor U3347 (N_3347,N_2494,N_2496);
and U3348 (N_3348,N_2135,N_2766);
nand U3349 (N_3349,N_1137,N_1781);
xor U3350 (N_3350,N_1024,N_984);
and U3351 (N_3351,N_1727,N_919);
or U3352 (N_3352,N_1198,N_172);
nor U3353 (N_3353,N_2188,N_2644);
or U3354 (N_3354,N_2856,N_2800);
nand U3355 (N_3355,N_2233,N_2974);
xnor U3356 (N_3356,N_63,N_291);
and U3357 (N_3357,N_2410,N_913);
xor U3358 (N_3358,N_1735,N_1736);
nand U3359 (N_3359,N_2699,N_1020);
nor U3360 (N_3360,N_761,N_2524);
xnor U3361 (N_3361,N_902,N_1748);
nor U3362 (N_3362,N_688,N_2992);
nor U3363 (N_3363,N_860,N_2667);
nand U3364 (N_3364,N_1366,N_1185);
nor U3365 (N_3365,N_1283,N_1909);
and U3366 (N_3366,N_1865,N_2005);
xor U3367 (N_3367,N_2968,N_1120);
or U3368 (N_3368,N_1224,N_1326);
xor U3369 (N_3369,N_2247,N_871);
xnor U3370 (N_3370,N_1278,N_2086);
nor U3371 (N_3371,N_1221,N_775);
and U3372 (N_3372,N_1232,N_1226);
nand U3373 (N_3373,N_224,N_1015);
and U3374 (N_3374,N_1033,N_1320);
nand U3375 (N_3375,N_161,N_1315);
xor U3376 (N_3376,N_1367,N_1256);
and U3377 (N_3377,N_2606,N_606);
nor U3378 (N_3378,N_375,N_180);
xnor U3379 (N_3379,N_1575,N_2431);
nand U3380 (N_3380,N_205,N_1771);
nand U3381 (N_3381,N_716,N_2419);
nand U3382 (N_3382,N_930,N_2199);
nand U3383 (N_3383,N_2426,N_2467);
or U3384 (N_3384,N_303,N_2881);
or U3385 (N_3385,N_758,N_686);
and U3386 (N_3386,N_1902,N_2753);
xor U3387 (N_3387,N_2038,N_1463);
nand U3388 (N_3388,N_2725,N_7);
or U3389 (N_3389,N_2327,N_89);
xnor U3390 (N_3390,N_1155,N_2129);
and U3391 (N_3391,N_489,N_901);
xor U3392 (N_3392,N_1243,N_111);
and U3393 (N_3393,N_2065,N_2413);
and U3394 (N_3394,N_1144,N_53);
nand U3395 (N_3395,N_2894,N_2241);
or U3396 (N_3396,N_1334,N_778);
nand U3397 (N_3397,N_823,N_2679);
nor U3398 (N_3398,N_2747,N_2995);
xor U3399 (N_3399,N_2833,N_173);
xor U3400 (N_3400,N_1798,N_382);
nor U3401 (N_3401,N_2611,N_1641);
nor U3402 (N_3402,N_2801,N_249);
and U3403 (N_3403,N_2772,N_1017);
xnor U3404 (N_3404,N_2382,N_2824);
nand U3405 (N_3405,N_2985,N_1978);
nand U3406 (N_3406,N_1455,N_216);
or U3407 (N_3407,N_177,N_2796);
nor U3408 (N_3408,N_329,N_265);
nand U3409 (N_3409,N_2702,N_616);
or U3410 (N_3410,N_2602,N_1924);
nand U3411 (N_3411,N_1088,N_2645);
and U3412 (N_3412,N_676,N_729);
or U3413 (N_3413,N_1960,N_2414);
xor U3414 (N_3414,N_2386,N_315);
nor U3415 (N_3415,N_1559,N_482);
or U3416 (N_3416,N_1390,N_1290);
and U3417 (N_3417,N_1333,N_1066);
nand U3418 (N_3418,N_1690,N_2898);
or U3419 (N_3419,N_1526,N_2063);
and U3420 (N_3420,N_522,N_2276);
or U3421 (N_3421,N_1307,N_1471);
xor U3422 (N_3422,N_1918,N_467);
xnor U3423 (N_3423,N_1822,N_1396);
and U3424 (N_3424,N_2178,N_2369);
xor U3425 (N_3425,N_1188,N_1756);
and U3426 (N_3426,N_32,N_103);
and U3427 (N_3427,N_2456,N_2571);
xnor U3428 (N_3428,N_1760,N_614);
xor U3429 (N_3429,N_1946,N_2993);
xnor U3430 (N_3430,N_1339,N_2961);
or U3431 (N_3431,N_2714,N_2533);
xnor U3432 (N_3432,N_1601,N_610);
xor U3433 (N_3433,N_58,N_2351);
and U3434 (N_3434,N_2136,N_837);
nand U3435 (N_3435,N_2623,N_821);
nor U3436 (N_3436,N_2567,N_2246);
xnor U3437 (N_3437,N_327,N_2516);
nor U3438 (N_3438,N_2045,N_2269);
nor U3439 (N_3439,N_682,N_1912);
nor U3440 (N_3440,N_1504,N_2083);
or U3441 (N_3441,N_1018,N_1779);
nand U3442 (N_3442,N_784,N_2642);
nor U3443 (N_3443,N_225,N_1205);
nor U3444 (N_3444,N_1067,N_544);
and U3445 (N_3445,N_1773,N_208);
xnor U3446 (N_3446,N_1449,N_310);
or U3447 (N_3447,N_1156,N_989);
and U3448 (N_3448,N_2684,N_2708);
nand U3449 (N_3449,N_316,N_1331);
nor U3450 (N_3450,N_596,N_1405);
nor U3451 (N_3451,N_1789,N_2110);
nand U3452 (N_3452,N_2535,N_479);
or U3453 (N_3453,N_2733,N_1238);
nor U3454 (N_3454,N_907,N_2743);
and U3455 (N_3455,N_1660,N_194);
nand U3456 (N_3456,N_367,N_2326);
nor U3457 (N_3457,N_2244,N_2831);
nor U3458 (N_3458,N_1244,N_2949);
nand U3459 (N_3459,N_1467,N_817);
and U3460 (N_3460,N_1294,N_23);
xnor U3461 (N_3461,N_193,N_1197);
or U3462 (N_3462,N_1795,N_1052);
nand U3463 (N_3463,N_1538,N_1029);
and U3464 (N_3464,N_2197,N_525);
and U3465 (N_3465,N_295,N_2835);
or U3466 (N_3466,N_376,N_1322);
nand U3467 (N_3467,N_2261,N_2624);
or U3468 (N_3468,N_1869,N_2286);
nor U3469 (N_3469,N_997,N_139);
nor U3470 (N_3470,N_36,N_890);
nand U3471 (N_3471,N_2735,N_1068);
nor U3472 (N_3472,N_1058,N_266);
nor U3473 (N_3473,N_2828,N_490);
and U3474 (N_3474,N_1527,N_2050);
and U3475 (N_3475,N_1929,N_762);
nand U3476 (N_3476,N_571,N_2857);
xor U3477 (N_3477,N_2274,N_502);
xor U3478 (N_3478,N_1898,N_1620);
xnor U3479 (N_3479,N_64,N_2390);
or U3480 (N_3480,N_629,N_1583);
xor U3481 (N_3481,N_710,N_22);
nor U3482 (N_3482,N_1562,N_2549);
nor U3483 (N_3483,N_2373,N_2060);
and U3484 (N_3484,N_1442,N_797);
nand U3485 (N_3485,N_2959,N_1196);
xor U3486 (N_3486,N_2457,N_1828);
nand U3487 (N_3487,N_2666,N_879);
nand U3488 (N_3488,N_1739,N_2168);
xor U3489 (N_3489,N_2093,N_1327);
xor U3490 (N_3490,N_1096,N_183);
nand U3491 (N_3491,N_991,N_1436);
or U3492 (N_3492,N_2757,N_1026);
and U3493 (N_3493,N_387,N_532);
nor U3494 (N_3494,N_1565,N_815);
nand U3495 (N_3495,N_26,N_977);
or U3496 (N_3496,N_2742,N_1885);
nor U3497 (N_3497,N_1164,N_1590);
xor U3498 (N_3498,N_2358,N_122);
xnor U3499 (N_3499,N_28,N_362);
nor U3500 (N_3500,N_1672,N_155);
and U3501 (N_3501,N_2130,N_2497);
xnor U3502 (N_3502,N_830,N_1295);
xor U3503 (N_3503,N_2784,N_1836);
or U3504 (N_3504,N_1899,N_2662);
nand U3505 (N_3505,N_1682,N_1937);
nor U3506 (N_3506,N_2360,N_1488);
nor U3507 (N_3507,N_2310,N_2707);
or U3508 (N_3508,N_745,N_1010);
and U3509 (N_3509,N_2983,N_1805);
nand U3510 (N_3510,N_1650,N_529);
or U3511 (N_3511,N_2008,N_2238);
and U3512 (N_3512,N_1841,N_2789);
and U3513 (N_3513,N_451,N_1519);
nand U3514 (N_3514,N_2315,N_2097);
nor U3515 (N_3515,N_185,N_143);
nor U3516 (N_3516,N_1539,N_2033);
nor U3517 (N_3517,N_2051,N_2123);
or U3518 (N_3518,N_1810,N_2682);
and U3519 (N_3519,N_619,N_2688);
and U3520 (N_3520,N_2716,N_2750);
nand U3521 (N_3521,N_2664,N_1472);
and U3522 (N_3522,N_1847,N_1189);
nor U3523 (N_3523,N_1536,N_1271);
and U3524 (N_3524,N_1321,N_617);
nand U3525 (N_3525,N_2864,N_2580);
nor U3526 (N_3526,N_435,N_321);
or U3527 (N_3527,N_2629,N_1234);
nand U3528 (N_3528,N_1281,N_2087);
nor U3529 (N_3529,N_2819,N_2203);
nand U3530 (N_3530,N_1838,N_1433);
xor U3531 (N_3531,N_2204,N_744);
nand U3532 (N_3532,N_776,N_277);
and U3533 (N_3533,N_1421,N_1399);
nand U3534 (N_3534,N_1464,N_869);
nand U3535 (N_3535,N_1425,N_345);
nand U3536 (N_3536,N_1280,N_2141);
nand U3537 (N_3537,N_2334,N_840);
or U3538 (N_3538,N_1934,N_2575);
and U3539 (N_3539,N_297,N_1203);
and U3540 (N_3540,N_2715,N_2852);
or U3541 (N_3541,N_2082,N_437);
nor U3542 (N_3542,N_1749,N_936);
xnor U3543 (N_3543,N_685,N_2070);
nor U3544 (N_3544,N_2231,N_1388);
or U3545 (N_3545,N_795,N_2291);
nand U3546 (N_3546,N_1231,N_388);
nor U3547 (N_3547,N_1720,N_399);
xnor U3548 (N_3548,N_1514,N_1957);
or U3549 (N_3549,N_2975,N_782);
or U3550 (N_3550,N_1744,N_160);
nor U3551 (N_3551,N_2635,N_2691);
and U3552 (N_3552,N_2421,N_1451);
xnor U3553 (N_3553,N_933,N_599);
and U3554 (N_3554,N_2263,N_259);
nor U3555 (N_3555,N_771,N_1431);
and U3556 (N_3556,N_967,N_581);
nor U3557 (N_3557,N_323,N_1199);
xnor U3558 (N_3558,N_4,N_1385);
nor U3559 (N_3559,N_1785,N_1379);
nor U3560 (N_3560,N_1372,N_2521);
and U3561 (N_3561,N_248,N_1703);
xor U3562 (N_3562,N_1787,N_1282);
nand U3563 (N_3563,N_2304,N_854);
nand U3564 (N_3564,N_2160,N_25);
and U3565 (N_3565,N_1742,N_1610);
and U3566 (N_3566,N_895,N_749);
or U3567 (N_3567,N_1797,N_320);
nor U3568 (N_3568,N_2359,N_2185);
nor U3569 (N_3569,N_549,N_1585);
and U3570 (N_3570,N_1365,N_628);
xnor U3571 (N_3571,N_2721,N_1395);
nand U3572 (N_3572,N_1972,N_2324);
nand U3573 (N_3573,N_2944,N_1161);
xnor U3574 (N_3574,N_1330,N_1541);
nand U3575 (N_3575,N_1528,N_1440);
nor U3576 (N_3576,N_1219,N_2036);
and U3577 (N_3577,N_1673,N_707);
or U3578 (N_3578,N_2064,N_884);
or U3579 (N_3579,N_2925,N_2131);
or U3580 (N_3580,N_2455,N_2034);
xnor U3581 (N_3581,N_355,N_2921);
xor U3582 (N_3582,N_243,N_2855);
or U3583 (N_3583,N_1958,N_2446);
nand U3584 (N_3584,N_853,N_2822);
nor U3585 (N_3585,N_553,N_843);
xor U3586 (N_3586,N_2977,N_1850);
xnor U3587 (N_3587,N_667,N_2508);
and U3588 (N_3588,N_151,N_750);
nand U3589 (N_3589,N_219,N_723);
xnor U3590 (N_3590,N_580,N_2207);
or U3591 (N_3591,N_2701,N_2811);
and U3592 (N_3592,N_1871,N_2367);
nand U3593 (N_3593,N_2159,N_1594);
nand U3594 (N_3594,N_2874,N_1949);
nand U3595 (N_3595,N_2637,N_2378);
and U3596 (N_3596,N_974,N_1324);
nand U3597 (N_3597,N_1407,N_2720);
nor U3598 (N_3598,N_953,N_1681);
nor U3599 (N_3599,N_1549,N_975);
xor U3600 (N_3600,N_1933,N_312);
and U3601 (N_3601,N_2669,N_713);
xor U3602 (N_3602,N_1090,N_1150);
and U3603 (N_3603,N_1345,N_1537);
nor U3604 (N_3604,N_658,N_2220);
xor U3605 (N_3605,N_441,N_1596);
nor U3606 (N_3606,N_2173,N_634);
xnor U3607 (N_3607,N_650,N_2880);
nor U3608 (N_3608,N_903,N_361);
nand U3609 (N_3609,N_572,N_908);
xor U3610 (N_3610,N_671,N_2095);
or U3611 (N_3611,N_2108,N_2940);
nand U3612 (N_3612,N_2998,N_2795);
nor U3613 (N_3613,N_1982,N_1938);
xor U3614 (N_3614,N_2495,N_801);
and U3615 (N_3615,N_2357,N_1483);
xor U3616 (N_3616,N_2260,N_1037);
or U3617 (N_3617,N_1501,N_1263);
nor U3618 (N_3618,N_1888,N_1796);
and U3619 (N_3619,N_2049,N_1002);
xor U3620 (N_3620,N_1487,N_706);
and U3621 (N_3621,N_1955,N_718);
xnor U3622 (N_3622,N_2023,N_354);
xor U3623 (N_3623,N_1874,N_2399);
nand U3624 (N_3624,N_2558,N_809);
or U3625 (N_3625,N_1657,N_2323);
and U3626 (N_3626,N_698,N_2727);
or U3627 (N_3627,N_19,N_1598);
and U3628 (N_3628,N_2826,N_1923);
nand U3629 (N_3629,N_2972,N_829);
and U3630 (N_3630,N_1762,N_2418);
xor U3631 (N_3631,N_91,N_2483);
nor U3632 (N_3632,N_67,N_232);
nor U3633 (N_3633,N_2032,N_1158);
or U3634 (N_3634,N_1038,N_1820);
nor U3635 (N_3635,N_1772,N_951);
nor U3636 (N_3636,N_1900,N_527);
xnor U3637 (N_3637,N_2119,N_870);
and U3638 (N_3638,N_734,N_1139);
or U3639 (N_3639,N_1168,N_2302);
nand U3640 (N_3640,N_738,N_157);
xor U3641 (N_3641,N_701,N_1914);
xor U3642 (N_3642,N_1632,N_728);
xnor U3643 (N_3643,N_760,N_1790);
xnor U3644 (N_3644,N_611,N_507);
nand U3645 (N_3645,N_1220,N_2107);
nor U3646 (N_3646,N_1172,N_1415);
or U3647 (N_3647,N_741,N_169);
xnor U3648 (N_3648,N_631,N_1485);
nand U3649 (N_3649,N_1494,N_450);
or U3650 (N_3650,N_578,N_1605);
and U3651 (N_3651,N_2216,N_34);
or U3652 (N_3652,N_1813,N_1054);
xnor U3653 (N_3653,N_792,N_306);
xor U3654 (N_3654,N_1078,N_2534);
xor U3655 (N_3655,N_2149,N_1412);
nand U3656 (N_3656,N_2464,N_825);
or U3657 (N_3657,N_1206,N_341);
and U3658 (N_3658,N_166,N_2433);
and U3659 (N_3659,N_2773,N_264);
nand U3660 (N_3660,N_1500,N_1401);
xor U3661 (N_3661,N_493,N_844);
and U3662 (N_3662,N_1786,N_1560);
nand U3663 (N_3663,N_1132,N_545);
or U3664 (N_3664,N_244,N_2793);
xor U3665 (N_3665,N_113,N_1653);
nand U3666 (N_3666,N_2525,N_1174);
nor U3667 (N_3667,N_708,N_2965);
and U3668 (N_3668,N_872,N_44);
or U3669 (N_3669,N_705,N_2412);
xor U3670 (N_3670,N_732,N_1839);
nor U3671 (N_3671,N_1730,N_2354);
nor U3672 (N_3672,N_2933,N_1624);
nor U3673 (N_3673,N_279,N_31);
nand U3674 (N_3674,N_2882,N_1529);
nor U3675 (N_3675,N_30,N_2938);
nand U3676 (N_3676,N_1458,N_979);
and U3677 (N_3677,N_1999,N_2930);
or U3678 (N_3678,N_1563,N_2658);
or U3679 (N_3679,N_83,N_727);
and U3680 (N_3680,N_427,N_2790);
and U3681 (N_3681,N_2546,N_2125);
xnor U3682 (N_3682,N_1503,N_2853);
nor U3683 (N_3683,N_1842,N_1693);
or U3684 (N_3684,N_117,N_2775);
or U3685 (N_3685,N_293,N_2132);
and U3686 (N_3686,N_2689,N_1776);
and U3687 (N_3687,N_2579,N_2807);
xor U3688 (N_3688,N_102,N_1230);
xor U3689 (N_3689,N_836,N_1212);
or U3690 (N_3690,N_562,N_1022);
or U3691 (N_3691,N_75,N_1622);
or U3692 (N_3692,N_2303,N_938);
xnor U3693 (N_3693,N_1831,N_184);
nand U3694 (N_3694,N_1584,N_1936);
xnor U3695 (N_3695,N_1432,N_2195);
nand U3696 (N_3696,N_2448,N_2561);
xor U3697 (N_3697,N_552,N_1336);
or U3698 (N_3698,N_1103,N_2616);
or U3699 (N_3699,N_1260,N_2167);
nand U3700 (N_3700,N_9,N_1546);
or U3701 (N_3701,N_2019,N_1687);
or U3702 (N_3702,N_2345,N_2799);
nor U3703 (N_3703,N_425,N_959);
nand U3704 (N_3704,N_1406,N_1732);
nor U3705 (N_3705,N_112,N_2655);
nor U3706 (N_3706,N_1076,N_2103);
and U3707 (N_3707,N_1545,N_2480);
xnor U3708 (N_3708,N_2252,N_1341);
nor U3709 (N_3709,N_1109,N_2926);
or U3710 (N_3710,N_258,N_1893);
and U3711 (N_3711,N_1328,N_1141);
xor U3712 (N_3712,N_1576,N_2779);
nand U3713 (N_3713,N_70,N_1285);
nor U3714 (N_3714,N_1079,N_398);
and U3715 (N_3715,N_1950,N_846);
nor U3716 (N_3716,N_2671,N_567);
nand U3717 (N_3717,N_1094,N_2328);
and U3718 (N_3718,N_748,N_1356);
and U3719 (N_3719,N_2865,N_2672);
and U3720 (N_3720,N_1532,N_1);
xor U3721 (N_3721,N_1963,N_2071);
or U3722 (N_3722,N_2249,N_2004);
nand U3723 (N_3723,N_2398,N_574);
xor U3724 (N_3724,N_1961,N_1272);
and U3725 (N_3725,N_2396,N_2058);
and U3726 (N_3726,N_805,N_693);
nand U3727 (N_3727,N_764,N_689);
nand U3728 (N_3728,N_342,N_773);
or U3729 (N_3729,N_1879,N_2783);
or U3730 (N_3730,N_52,N_2765);
nand U3731 (N_3731,N_579,N_1631);
nand U3732 (N_3732,N_2928,N_1499);
nand U3733 (N_3733,N_95,N_1352);
nor U3734 (N_3734,N_1439,N_537);
or U3735 (N_3735,N_1550,N_1317);
nor U3736 (N_3736,N_643,N_947);
xnor U3737 (N_3737,N_179,N_1557);
nand U3738 (N_3738,N_1835,N_1291);
nand U3739 (N_3739,N_530,N_2578);
nand U3740 (N_3740,N_2817,N_218);
xor U3741 (N_3741,N_956,N_2964);
and U3742 (N_3742,N_878,N_392);
and U3743 (N_3743,N_2306,N_1077);
and U3744 (N_3744,N_2879,N_1211);
and U3745 (N_3745,N_2999,N_937);
or U3746 (N_3746,N_2934,N_993);
xnor U3747 (N_3747,N_1477,N_1765);
nor U3748 (N_3748,N_1381,N_2098);
nor U3749 (N_3749,N_2522,N_607);
nand U3750 (N_3750,N_281,N_142);
nand U3751 (N_3751,N_2866,N_2009);
or U3752 (N_3752,N_2659,N_108);
and U3753 (N_3753,N_2047,N_1895);
and U3754 (N_3754,N_2778,N_2556);
and U3755 (N_3755,N_2237,N_952);
nand U3756 (N_3756,N_865,N_900);
and U3757 (N_3757,N_1269,N_2991);
and U3758 (N_3758,N_2124,N_1606);
xor U3759 (N_3759,N_322,N_736);
and U3760 (N_3760,N_2929,N_2982);
xor U3761 (N_3761,N_72,N_1837);
and U3762 (N_3762,N_337,N_124);
and U3763 (N_3763,N_431,N_48);
and U3764 (N_3764,N_2514,N_484);
and U3765 (N_3765,N_1008,N_1394);
and U3766 (N_3766,N_309,N_2206);
nor U3767 (N_3767,N_2531,N_796);
xnor U3768 (N_3768,N_1507,N_1623);
xor U3769 (N_3769,N_1296,N_1484);
or U3770 (N_3770,N_1701,N_2791);
and U3771 (N_3771,N_2802,N_1521);
or U3772 (N_3772,N_2422,N_1251);
and U3773 (N_3773,N_1178,N_915);
nor U3774 (N_3774,N_1053,N_2844);
nor U3775 (N_3775,N_867,N_881);
nor U3776 (N_3776,N_2251,N_781);
nor U3777 (N_3777,N_1039,N_204);
nor U3778 (N_3778,N_2417,N_833);
nor U3779 (N_3779,N_2559,N_1261);
or U3780 (N_3780,N_1848,N_1236);
xnor U3781 (N_3781,N_2476,N_2510);
nand U3782 (N_3782,N_1534,N_2670);
and U3783 (N_3783,N_2309,N_499);
nor U3784 (N_3784,N_2429,N_2769);
nand U3785 (N_3785,N_1932,N_2395);
xnor U3786 (N_3786,N_96,N_434);
nor U3787 (N_3787,N_1277,N_2030);
and U3788 (N_3788,N_1253,N_2277);
and U3789 (N_3789,N_2213,N_1142);
xor U3790 (N_3790,N_2177,N_452);
xor U3791 (N_3791,N_1512,N_1134);
nor U3792 (N_3792,N_1016,N_2935);
xnor U3793 (N_3793,N_582,N_1025);
nand U3794 (N_3794,N_1635,N_2717);
or U3795 (N_3795,N_1200,N_2243);
xor U3796 (N_3796,N_550,N_637);
or U3797 (N_3797,N_752,N_2145);
nor U3798 (N_3798,N_1210,N_2673);
nand U3799 (N_3799,N_845,N_2563);
xnor U3800 (N_3800,N_1304,N_1830);
or U3801 (N_3801,N_656,N_1754);
xnor U3802 (N_3802,N_2014,N_2214);
or U3803 (N_3803,N_1833,N_85);
or U3804 (N_3804,N_2026,N_2002);
nor U3805 (N_3805,N_256,N_1074);
xor U3806 (N_3806,N_1802,N_2976);
nor U3807 (N_3807,N_492,N_197);
nor U3808 (N_3808,N_271,N_2909);
or U3809 (N_3809,N_1941,N_162);
and U3810 (N_3810,N_2021,N_137);
or U3811 (N_3811,N_2139,N_1552);
nand U3812 (N_3812,N_2201,N_2407);
or U3813 (N_3813,N_735,N_1671);
or U3814 (N_3814,N_700,N_1119);
xnor U3815 (N_3815,N_626,N_1750);
nor U3816 (N_3816,N_2869,N_1098);
or U3817 (N_3817,N_1191,N_1204);
and U3818 (N_3818,N_1654,N_1049);
or U3819 (N_3819,N_1611,N_2912);
and U3820 (N_3820,N_826,N_1410);
nand U3821 (N_3821,N_2271,N_2883);
and U3822 (N_3822,N_1292,N_2861);
and U3823 (N_3823,N_2171,N_1954);
nand U3824 (N_3824,N_167,N_107);
and U3825 (N_3825,N_1289,N_444);
and U3826 (N_3826,N_2052,N_1638);
xor U3827 (N_3827,N_1655,N_2858);
and U3828 (N_3828,N_2581,N_1403);
and U3829 (N_3829,N_1652,N_430);
nor U3830 (N_3830,N_1769,N_2194);
nand U3831 (N_3831,N_1987,N_402);
xor U3832 (N_3832,N_1057,N_1547);
nor U3833 (N_3833,N_969,N_357);
xor U3834 (N_3834,N_2265,N_2217);
nor U3835 (N_3835,N_191,N_2377);
nor U3836 (N_3836,N_332,N_42);
nor U3837 (N_3837,N_2292,N_1832);
xor U3838 (N_3838,N_2273,N_1264);
or U3839 (N_3839,N_506,N_601);
nand U3840 (N_3840,N_1023,N_2112);
or U3841 (N_3841,N_2910,N_2028);
xor U3842 (N_3842,N_2562,N_2751);
and U3843 (N_3843,N_1173,N_1930);
or U3844 (N_3844,N_1998,N_1766);
xnor U3845 (N_3845,N_2335,N_2227);
or U3846 (N_3846,N_2253,N_2729);
xnor U3847 (N_3847,N_2942,N_394);
xnor U3848 (N_3848,N_115,N_2074);
xor U3849 (N_3849,N_2971,N_462);
and U3850 (N_3850,N_2054,N_2512);
nand U3851 (N_3851,N_2040,N_328);
and U3852 (N_3852,N_916,N_1649);
and U3853 (N_3853,N_1213,N_759);
xor U3854 (N_3854,N_247,N_384);
or U3855 (N_3855,N_453,N_154);
nand U3856 (N_3856,N_2053,N_2889);
nand U3857 (N_3857,N_33,N_1759);
or U3858 (N_3858,N_41,N_210);
nand U3859 (N_3859,N_651,N_2505);
or U3860 (N_3860,N_1180,N_2694);
or U3861 (N_3861,N_2389,N_2042);
nor U3862 (N_3862,N_2472,N_1696);
or U3863 (N_3863,N_2657,N_2986);
xnor U3864 (N_3864,N_2348,N_1782);
nand U3865 (N_3865,N_201,N_2540);
and U3866 (N_3866,N_1071,N_2376);
nor U3867 (N_3867,N_564,N_391);
or U3868 (N_3868,N_2695,N_2827);
and U3869 (N_3869,N_1889,N_84);
xor U3870 (N_3870,N_1443,N_2610);
or U3871 (N_3871,N_666,N_1741);
or U3872 (N_3872,N_1680,N_983);
nand U3873 (N_3873,N_661,N_1777);
nor U3874 (N_3874,N_680,N_343);
or U3875 (N_3875,N_928,N_2532);
nand U3876 (N_3876,N_1864,N_2096);
nand U3877 (N_3877,N_1095,N_2843);
and U3878 (N_3878,N_50,N_1684);
xnor U3879 (N_3879,N_1591,N_2264);
and U3880 (N_3880,N_852,N_1266);
xnor U3881 (N_3881,N_2313,N_472);
nor U3882 (N_3882,N_875,N_409);
nor U3883 (N_3883,N_538,N_300);
and U3884 (N_3884,N_1145,N_254);
nor U3885 (N_3885,N_2786,N_2962);
nand U3886 (N_3886,N_1574,N_595);
or U3887 (N_3887,N_29,N_1801);
or U3888 (N_3888,N_1361,N_897);
nor U3889 (N_3889,N_2117,N_1970);
xnor U3890 (N_3890,N_1718,N_1997);
nand U3891 (N_3891,N_1780,N_963);
nand U3892 (N_3892,N_1824,N_2943);
nor U3893 (N_3893,N_182,N_2470);
nor U3894 (N_3894,N_2639,N_2528);
nor U3895 (N_3895,N_1677,N_2760);
nand U3896 (N_3896,N_962,N_2675);
or U3897 (N_3897,N_585,N_1665);
nand U3898 (N_3898,N_1194,N_2325);
or U3899 (N_3899,N_2381,N_217);
or U3900 (N_3900,N_2809,N_1217);
nand U3901 (N_3901,N_2270,N_2435);
and U3902 (N_3902,N_737,N_2897);
or U3903 (N_3903,N_1540,N_2405);
and U3904 (N_3904,N_460,N_554);
xnor U3905 (N_3905,N_267,N_586);
xor U3906 (N_3906,N_105,N_414);
or U3907 (N_3907,N_475,N_996);
and U3908 (N_3908,N_21,N_1708);
xor U3909 (N_3909,N_2434,N_1102);
xnor U3910 (N_3910,N_511,N_1712);
nor U3911 (N_3911,N_209,N_772);
and U3912 (N_3912,N_2776,N_898);
or U3913 (N_3913,N_1815,N_832);
and U3914 (N_3914,N_1592,N_664);
nor U3915 (N_3915,N_576,N_126);
nand U3916 (N_3916,N_45,N_1979);
xor U3917 (N_3917,N_1853,N_1778);
xor U3918 (N_3918,N_2718,N_1855);
and U3919 (N_3919,N_1694,N_2293);
nand U3920 (N_3920,N_152,N_539);
or U3921 (N_3921,N_146,N_278);
nor U3922 (N_3922,N_1434,N_559);
and U3923 (N_3923,N_2570,N_1216);
or U3924 (N_3924,N_2674,N_296);
nor U3925 (N_3925,N_740,N_236);
xnor U3926 (N_3926,N_1473,N_632);
and U3927 (N_3927,N_2951,N_609);
nand U3928 (N_3928,N_1190,N_1734);
nand U3929 (N_3929,N_820,N_351);
or U3930 (N_3930,N_859,N_156);
nand U3931 (N_3931,N_2461,N_800);
nor U3932 (N_3932,N_726,N_889);
nor U3933 (N_3933,N_850,N_1799);
and U3934 (N_3934,N_807,N_2955);
nor U3935 (N_3935,N_386,N_1884);
xor U3936 (N_3936,N_1868,N_2183);
xor U3937 (N_3937,N_340,N_212);
and U3938 (N_3938,N_623,N_2007);
xnor U3939 (N_3939,N_80,N_2792);
or U3940 (N_3940,N_657,N_2180);
and U3941 (N_3941,N_299,N_1625);
nor U3942 (N_3942,N_1101,N_1414);
and U3943 (N_3943,N_82,N_2686);
xor U3944 (N_3944,N_2312,N_98);
or U3945 (N_3945,N_1636,N_703);
or U3946 (N_3946,N_583,N_1728);
xnor U3947 (N_3947,N_906,N_2638);
xor U3948 (N_3948,N_263,N_2100);
and U3949 (N_3949,N_76,N_2960);
nor U3950 (N_3950,N_2948,N_2947);
nand U3951 (N_3951,N_926,N_1301);
nor U3952 (N_3952,N_2228,N_1218);
nand U3953 (N_3953,N_558,N_227);
nor U3954 (N_3954,N_1105,N_627);
or U3955 (N_3955,N_2475,N_1447);
or U3956 (N_3956,N_2279,N_1225);
xor U3957 (N_3957,N_2958,N_2979);
xor U3958 (N_3958,N_1683,N_2939);
nor U3959 (N_3959,N_1303,N_1107);
xor U3960 (N_3960,N_242,N_2126);
and U3961 (N_3961,N_1048,N_230);
or U3962 (N_3962,N_1983,N_373);
or U3963 (N_3963,N_283,N_934);
or U3964 (N_3964,N_946,N_2297);
and U3965 (N_3965,N_1858,N_1310);
nand U3966 (N_3966,N_717,N_1116);
or U3967 (N_3967,N_366,N_912);
nor U3968 (N_3968,N_2745,N_1851);
nand U3969 (N_3969,N_806,N_1423);
nor U3970 (N_3970,N_1242,N_1444);
nor U3971 (N_3971,N_2631,N_1710);
nor U3972 (N_3972,N_1896,N_1041);
or U3973 (N_3973,N_1497,N_1597);
xor U3974 (N_3974,N_165,N_369);
nand U3975 (N_3975,N_819,N_1492);
nand U3976 (N_3976,N_2970,N_2120);
or U3977 (N_3977,N_2343,N_2851);
or U3978 (N_3978,N_786,N_981);
and U3979 (N_3979,N_561,N_774);
or U3980 (N_3980,N_1988,N_1729);
nor U3981 (N_3981,N_2829,N_514);
nor U3982 (N_3982,N_2154,N_1792);
and U3983 (N_3983,N_2878,N_364);
xor U3984 (N_3984,N_17,N_2845);
nand U3985 (N_3985,N_931,N_876);
and U3986 (N_3986,N_813,N_233);
or U3987 (N_3987,N_2200,N_269);
xor U3988 (N_3988,N_1952,N_569);
nand U3989 (N_3989,N_2428,N_206);
or U3990 (N_3990,N_79,N_2439);
xnor U3991 (N_3991,N_835,N_757);
nand U3992 (N_3992,N_2891,N_2536);
nor U3993 (N_3993,N_257,N_2808);
xor U3994 (N_3994,N_1768,N_2665);
nand U3995 (N_3995,N_2432,N_240);
xor U3996 (N_3996,N_2603,N_533);
or U3997 (N_3997,N_2850,N_24);
or U3998 (N_3998,N_365,N_1872);
or U3999 (N_3999,N_1980,N_2319);
and U4000 (N_4000,N_2336,N_1389);
nand U4001 (N_4001,N_2454,N_1984);
nand U4002 (N_4002,N_1628,N_2996);
and U4003 (N_4003,N_504,N_1784);
nor U4004 (N_4004,N_2466,N_1816);
and U4005 (N_4005,N_1311,N_2415);
or U4006 (N_4006,N_739,N_1019);
xnor U4007 (N_4007,N_1138,N_1880);
or U4008 (N_4008,N_2056,N_1719);
or U4009 (N_4009,N_1926,N_421);
nor U4010 (N_4010,N_1666,N_811);
xnor U4011 (N_4011,N_2146,N_1005);
or U4012 (N_4012,N_715,N_652);
xor U4013 (N_4013,N_1195,N_2447);
and U4014 (N_4014,N_2756,N_228);
nand U4015 (N_4015,N_2174,N_1969);
nand U4016 (N_4016,N_2823,N_118);
or U4017 (N_4017,N_2587,N_998);
and U4018 (N_4018,N_1104,N_2424);
nand U4019 (N_4019,N_324,N_594);
nor U4020 (N_4020,N_463,N_2872);
xor U4021 (N_4021,N_2574,N_2048);
xor U4022 (N_4022,N_863,N_2816);
nor U4023 (N_4023,N_255,N_2566);
and U4024 (N_4024,N_2090,N_1925);
xnor U4025 (N_4025,N_178,N_2338);
nand U4026 (N_4026,N_2339,N_198);
and U4027 (N_4027,N_2471,N_2908);
and U4028 (N_4028,N_2409,N_2696);
xor U4029 (N_4029,N_927,N_448);
xnor U4030 (N_4030,N_2698,N_882);
nand U4031 (N_4031,N_1349,N_1812);
nor U4032 (N_4032,N_1129,N_2821);
nand U4033 (N_4033,N_1110,N_1376);
nor U4034 (N_4034,N_1821,N_2690);
nand U4035 (N_4035,N_2158,N_1465);
xnor U4036 (N_4036,N_957,N_1131);
or U4037 (N_4037,N_1475,N_59);
xnor U4038 (N_4038,N_2841,N_1258);
xor U4039 (N_4039,N_874,N_2519);
nor U4040 (N_4040,N_2307,N_2768);
nor U4041 (N_4041,N_566,N_2078);
and U4042 (N_4042,N_920,N_1466);
and U4043 (N_4043,N_711,N_660);
or U4044 (N_4044,N_1344,N_1081);
xor U4045 (N_4045,N_2632,N_2250);
nand U4046 (N_4046,N_1700,N_803);
nand U4047 (N_4047,N_2630,N_2842);
or U4048 (N_4048,N_654,N_2544);
nor U4049 (N_4049,N_2225,N_1353);
nand U4050 (N_4050,N_2887,N_1363);
nand U4051 (N_4051,N_2166,N_1706);
or U4052 (N_4052,N_648,N_1911);
xor U4053 (N_4053,N_1456,N_1176);
nand U4054 (N_4054,N_1030,N_531);
xor U4055 (N_4055,N_649,N_885);
or U4056 (N_4056,N_2815,N_918);
xnor U4057 (N_4057,N_1408,N_765);
or U4058 (N_4058,N_273,N_789);
or U4059 (N_4059,N_231,N_1386);
nor U4060 (N_4060,N_1287,N_1409);
and U4061 (N_4061,N_645,N_1416);
xnor U4062 (N_4062,N_1733,N_2905);
xor U4063 (N_4063,N_2094,N_2318);
nand U4064 (N_4064,N_241,N_2539);
nor U4065 (N_4065,N_483,N_573);
xnor U4066 (N_4066,N_1027,N_1373);
nor U4067 (N_4067,N_1011,N_8);
xnor U4068 (N_4068,N_353,N_1167);
or U4069 (N_4069,N_275,N_1080);
nor U4070 (N_4070,N_1616,N_699);
xnor U4071 (N_4071,N_2289,N_777);
nor U4072 (N_4072,N_2101,N_1523);
or U4073 (N_4073,N_393,N_400);
xor U4074 (N_4074,N_1945,N_568);
nand U4075 (N_4075,N_1878,N_1418);
or U4076 (N_4076,N_2212,N_2812);
xor U4077 (N_4077,N_1130,N_2838);
nand U4078 (N_4078,N_886,N_1704);
nand U4079 (N_4079,N_1084,N_2296);
xnor U4080 (N_4080,N_413,N_982);
and U4081 (N_4081,N_1299,N_1004);
nor U4082 (N_4082,N_1755,N_1685);
nor U4083 (N_4083,N_1495,N_2012);
xor U4084 (N_4084,N_2035,N_1288);
xor U4085 (N_4085,N_516,N_2138);
nand U4086 (N_4086,N_223,N_1239);
xnor U4087 (N_4087,N_433,N_2308);
nand U4088 (N_4088,N_1859,N_97);
nand U4089 (N_4089,N_2888,N_2436);
nor U4090 (N_4090,N_2804,N_416);
or U4091 (N_4091,N_2374,N_839);
and U4092 (N_4092,N_1021,N_1491);
or U4093 (N_4093,N_1861,N_133);
and U4094 (N_4094,N_2503,N_2182);
or U4095 (N_4095,N_2922,N_1707);
and U4096 (N_4096,N_1876,N_1055);
or U4097 (N_4097,N_14,N_347);
and U4098 (N_4098,N_1823,N_2479);
nor U4099 (N_4099,N_1274,N_528);
nand U4100 (N_4100,N_170,N_2825);
xor U4101 (N_4101,N_973,N_2208);
or U4102 (N_4102,N_2507,N_65);
xnor U4103 (N_4103,N_2018,N_1863);
nand U4104 (N_4104,N_624,N_318);
nand U4105 (N_4105,N_2383,N_1567);
xor U4106 (N_4106,N_1891,N_1170);
nor U4107 (N_4107,N_1391,N_2731);
and U4108 (N_4108,N_2890,N_1113);
xnor U4109 (N_4109,N_94,N_2877);
nand U4110 (N_4110,N_1511,N_1633);
or U4111 (N_4111,N_1273,N_288);
and U4112 (N_4112,N_1524,N_1133);
nand U4113 (N_4113,N_2941,N_246);
xor U4114 (N_4114,N_721,N_2491);
and U4115 (N_4115,N_746,N_1459);
nor U4116 (N_4116,N_2330,N_2420);
or U4117 (N_4117,N_381,N_106);
xnor U4118 (N_4118,N_2529,N_1800);
xor U4119 (N_4119,N_1486,N_1976);
xor U4120 (N_4120,N_958,N_2771);
or U4121 (N_4121,N_808,N_1518);
nor U4122 (N_4122,N_2242,N_2176);
nand U4123 (N_4123,N_1387,N_455);
or U4124 (N_4124,N_2683,N_1586);
nand U4125 (N_4125,N_672,N_37);
xor U4126 (N_4126,N_2687,N_2280);
or U4127 (N_4127,N_2759,N_2994);
nand U4128 (N_4128,N_313,N_2832);
nor U4129 (N_4129,N_2634,N_2137);
xor U4130 (N_4130,N_461,N_2914);
xor U4131 (N_4131,N_2481,N_2337);
nor U4132 (N_4132,N_1814,N_15);
nand U4133 (N_4133,N_2651,N_1430);
nor U4134 (N_4134,N_2584,N_720);
xor U4135 (N_4135,N_2462,N_168);
nor U4136 (N_4136,N_1437,N_2513);
xnor U4137 (N_4137,N_1229,N_2596);
xnor U4138 (N_4138,N_222,N_164);
and U4139 (N_4139,N_1915,N_1419);
nor U4140 (N_4140,N_1400,N_684);
nand U4141 (N_4141,N_423,N_1692);
xor U4142 (N_4142,N_1398,N_2900);
nand U4143 (N_4143,N_827,N_1663);
or U4144 (N_4144,N_940,N_961);
and U4145 (N_4145,N_100,N_2617);
nand U4146 (N_4146,N_694,N_2474);
nor U4147 (N_4147,N_302,N_1371);
nor U4148 (N_4148,N_454,N_77);
xor U4149 (N_4149,N_1506,N_2952);
xor U4150 (N_4150,N_1031,N_10);
or U4151 (N_4151,N_1378,N_1962);
and U4152 (N_4152,N_1154,N_1306);
and U4153 (N_4153,N_2585,N_743);
nand U4154 (N_4154,N_406,N_1840);
and U4155 (N_4155,N_712,N_1723);
or U4156 (N_4156,N_1639,N_457);
xnor U4157 (N_4157,N_1249,N_2552);
nor U4158 (N_4158,N_1564,N_314);
and U4159 (N_4159,N_57,N_2728);
nor U4160 (N_4160,N_2625,N_1968);
xnor U4161 (N_4161,N_1006,N_1721);
nand U4162 (N_4162,N_2920,N_642);
and U4163 (N_4163,N_2794,N_2140);
and U4164 (N_4164,N_822,N_1424);
nor U4165 (N_4165,N_2722,N_1014);
or U4166 (N_4166,N_2430,N_877);
and U4167 (N_4167,N_2780,N_1209);
xnor U4168 (N_4168,N_2538,N_2371);
or U4169 (N_4169,N_1809,N_588);
nor U4170 (N_4170,N_1342,N_1259);
nor U4171 (N_4171,N_1046,N_2347);
or U4172 (N_4172,N_2848,N_147);
and U4173 (N_4173,N_2613,N_66);
nand U4174 (N_4174,N_841,N_192);
nor U4175 (N_4175,N_199,N_2678);
xnor U4176 (N_4176,N_1580,N_600);
nor U4177 (N_4177,N_2011,N_2104);
or U4178 (N_4178,N_1916,N_663);
or U4179 (N_4179,N_541,N_480);
nand U4180 (N_4180,N_2478,N_2656);
xor U4181 (N_4181,N_1867,N_1157);
nor U4182 (N_4182,N_515,N_914);
nand U4183 (N_4183,N_921,N_2847);
nor U4184 (N_4184,N_904,N_1646);
nand U4185 (N_4185,N_2340,N_252);
xor U4186 (N_4186,N_1986,N_523);
and U4187 (N_4187,N_494,N_1075);
and U4188 (N_4188,N_988,N_722);
or U4189 (N_4189,N_2763,N_1044);
or U4190 (N_4190,N_976,N_2530);
nor U4191 (N_4191,N_814,N_474);
nand U4192 (N_4192,N_2192,N_495);
and U4193 (N_4193,N_55,N_935);
or U4194 (N_4194,N_2668,N_1312);
and U4195 (N_4195,N_950,N_1340);
nand U4196 (N_4196,N_1121,N_1808);
and U4197 (N_4197,N_2240,N_1426);
or U4198 (N_4198,N_2859,N_1348);
nor U4199 (N_4199,N_260,N_2163);
xnor U4200 (N_4200,N_2576,N_445);
nand U4201 (N_4201,N_509,N_2076);
or U4202 (N_4202,N_1355,N_350);
nand U4203 (N_4203,N_929,N_1151);
xor U4204 (N_4204,N_1940,N_171);
or U4205 (N_4205,N_46,N_1854);
and U4206 (N_4206,N_519,N_2526);
nand U4207 (N_4207,N_2597,N_2113);
or U4208 (N_4208,N_1122,N_363);
xor U4209 (N_4209,N_1626,N_2646);
nor U4210 (N_4210,N_2806,N_2368);
nand U4211 (N_4211,N_1152,N_2234);
and U4212 (N_4212,N_1042,N_1186);
xnor U4213 (N_4213,N_1775,N_2179);
or U4214 (N_4214,N_1099,N_334);
nor U4215 (N_4215,N_1207,N_1901);
or U4216 (N_4216,N_1944,N_697);
or U4217 (N_4217,N_1181,N_412);
and U4218 (N_4218,N_1882,N_464);
nor U4219 (N_4219,N_2741,N_1034);
nor U4220 (N_4220,N_1092,N_2553);
or U4221 (N_4221,N_2680,N_2268);
or U4222 (N_4222,N_2406,N_2649);
nor U4223 (N_4223,N_787,N_2906);
nor U4224 (N_4224,N_1516,N_1903);
xor U4225 (N_4225,N_1921,N_43);
or U4226 (N_4226,N_134,N_1284);
nor U4227 (N_4227,N_285,N_1165);
nand U4228 (N_4228,N_2189,N_864);
and U4229 (N_4229,N_608,N_2370);
or U4230 (N_4230,N_1056,N_1083);
nor U4231 (N_4231,N_196,N_477);
nor U4232 (N_4232,N_517,N_1193);
xnor U4233 (N_4233,N_158,N_1060);
or U4234 (N_4234,N_235,N_1166);
and U4235 (N_4235,N_1643,N_1731);
nand U4236 (N_4236,N_424,N_317);
nand U4237 (N_4237,N_145,N_893);
nor U4238 (N_4238,N_2449,N_1761);
and U4239 (N_4239,N_73,N_1566);
and U4240 (N_4240,N_942,N_1050);
nor U4241 (N_4241,N_1404,N_374);
nand U4242 (N_4242,N_1846,N_1035);
xnor U4243 (N_4243,N_1752,N_5);
xnor U4244 (N_4244,N_1825,N_2723);
xnor U4245 (N_4245,N_282,N_2957);
nor U4246 (N_4246,N_385,N_1255);
nand U4247 (N_4247,N_1670,N_2924);
xnor U4248 (N_4248,N_518,N_646);
xnor U4249 (N_4249,N_1493,N_702);
xnor U4250 (N_4250,N_2245,N_892);
or U4251 (N_4251,N_999,N_1602);
xor U4252 (N_4252,N_1819,N_2452);
nand U4253 (N_4253,N_1476,N_2997);
or U4254 (N_4254,N_2484,N_2485);
xor U4255 (N_4255,N_943,N_1826);
xor U4256 (N_4256,N_2,N_925);
nand U4257 (N_4257,N_2626,N_681);
xnor U4258 (N_4258,N_1803,N_1588);
xor U4259 (N_4259,N_2931,N_1758);
xor U4260 (N_4260,N_1845,N_90);
and U4261 (N_4261,N_200,N_1614);
or U4262 (N_4262,N_598,N_1737);
nor U4263 (N_4263,N_148,N_2814);
xor U4264 (N_4264,N_2499,N_1967);
nor U4265 (N_4265,N_234,N_1866);
nor U4266 (N_4266,N_2917,N_1368);
xor U4267 (N_4267,N_1607,N_2612);
nor U4268 (N_4268,N_2144,N_2593);
nor U4269 (N_4269,N_2711,N_2089);
and U4270 (N_4270,N_1293,N_211);
or U4271 (N_4271,N_2966,N_2239);
or U4272 (N_4272,N_856,N_2205);
nand U4273 (N_4273,N_639,N_2157);
nor U4274 (N_4274,N_798,N_396);
or U4275 (N_4275,N_2298,N_370);
nand U4276 (N_4276,N_725,N_92);
or U4277 (N_4277,N_2295,N_1890);
nand U4278 (N_4278,N_1065,N_1711);
and U4279 (N_4279,N_2106,N_1875);
or U4280 (N_4280,N_274,N_503);
xor U4281 (N_4281,N_1007,N_383);
and U4282 (N_4282,N_2660,N_2609);
xor U4283 (N_4283,N_1910,N_1994);
and U4284 (N_4284,N_1462,N_604);
or U4285 (N_4285,N_2591,N_1202);
and U4286 (N_4286,N_849,N_2919);
and U4287 (N_4287,N_1615,N_136);
and U4288 (N_4288,N_2709,N_1452);
nand U4289 (N_4289,N_2443,N_1358);
nor U4290 (N_4290,N_411,N_1807);
nor U4291 (N_4291,N_2222,N_2820);
or U4292 (N_4292,N_2165,N_39);
nor U4293 (N_4293,N_1086,N_2344);
and U4294 (N_4294,N_1659,N_2198);
xor U4295 (N_4295,N_1360,N_2175);
nor U4296 (N_4296,N_1490,N_2936);
nand U4297 (N_4297,N_1106,N_439);
and U4298 (N_4298,N_2777,N_2352);
xor U4299 (N_4299,N_862,N_1763);
nand U4300 (N_4300,N_2590,N_2172);
nand U4301 (N_4301,N_348,N_2572);
and U4302 (N_4302,N_1642,N_2980);
or U4303 (N_4303,N_1908,N_2288);
nor U4304 (N_4304,N_2550,N_1402);
or U4305 (N_4305,N_438,N_2275);
nand U4306 (N_4306,N_308,N_1679);
nor U4307 (N_4307,N_410,N_1279);
or U4308 (N_4308,N_485,N_1783);
nor U4309 (N_4309,N_2088,N_2321);
nand U4310 (N_4310,N_54,N_2438);
or U4311 (N_4311,N_116,N_1318);
and U4312 (N_4312,N_691,N_1593);
and U4313 (N_4313,N_336,N_2284);
or U4314 (N_4314,N_1548,N_2356);
nand U4315 (N_4315,N_449,N_389);
xor U4316 (N_4316,N_2150,N_1640);
xor U4317 (N_4317,N_577,N_2600);
and U4318 (N_4318,N_1482,N_2105);
xor U4319 (N_4319,N_405,N_1276);
xnor U4320 (N_4320,N_18,N_1369);
nand U4321 (N_4321,N_229,N_1059);
and U4322 (N_4322,N_1747,N_1531);
and U4323 (N_4323,N_2601,N_1743);
xor U4324 (N_4324,N_2029,N_87);
or U4325 (N_4325,N_592,N_1965);
xnor U4326 (N_4326,N_346,N_2196);
xor U4327 (N_4327,N_780,N_1297);
nand U4328 (N_4328,N_1556,N_2465);
nand U4329 (N_4329,N_144,N_2224);
and U4330 (N_4330,N_1338,N_1422);
and U4331 (N_4331,N_2608,N_2006);
nor U4332 (N_4332,N_1817,N_653);
xor U4333 (N_4333,N_851,N_677);
and U4334 (N_4334,N_2115,N_1032);
nor U4335 (N_4335,N_2749,N_13);
nand U4336 (N_4336,N_1894,N_2545);
nand U4337 (N_4337,N_2902,N_333);
nor U4338 (N_4338,N_2586,N_104);
nand U4339 (N_4339,N_2294,N_2316);
and U4340 (N_4340,N_1135,N_2923);
nor U4341 (N_4341,N_2764,N_319);
xnor U4342 (N_4342,N_1350,N_2440);
xor U4343 (N_4343,N_99,N_1971);
and U4344 (N_4344,N_709,N_675);
and U4345 (N_4345,N_2259,N_615);
and U4346 (N_4346,N_250,N_2084);
xnor U4347 (N_4347,N_2148,N_1603);
nand U4348 (N_4348,N_1668,N_2754);
nor U4349 (N_4349,N_2362,N_1240);
nand U4350 (N_4350,N_2394,N_793);
or U4351 (N_4351,N_2184,N_1555);
nand U4352 (N_4352,N_2614,N_1246);
and U4353 (N_4353,N_1347,N_1270);
nand U4354 (N_4354,N_408,N_2736);
and U4355 (N_4355,N_1384,N_2770);
nor U4356 (N_4356,N_500,N_1175);
nor U4357 (N_4357,N_1553,N_618);
nor U4358 (N_4358,N_965,N_2973);
and U4359 (N_4359,N_1774,N_1873);
and U4360 (N_4360,N_1767,N_2969);
xor U4361 (N_4361,N_540,N_213);
xor U4362 (N_4362,N_923,N_2463);
and U4363 (N_4363,N_2839,N_1791);
nand U4364 (N_4364,N_1907,N_932);
xnor U4365 (N_4365,N_767,N_1325);
and U4366 (N_4366,N_2589,N_794);
or U4367 (N_4367,N_2732,N_1881);
nor U4368 (N_4368,N_1942,N_2342);
nand U4369 (N_4369,N_2229,N_1100);
xor U4370 (N_4370,N_2633,N_1956);
nor U4371 (N_4371,N_2059,N_687);
nand U4372 (N_4372,N_426,N_292);
nor U4373 (N_4373,N_2636,N_1182);
nand U4374 (N_4374,N_2451,N_2813);
xor U4375 (N_4375,N_1302,N_1159);
and U4376 (N_4376,N_1609,N_1697);
nand U4377 (N_4377,N_1040,N_101);
or U4378 (N_4378,N_2190,N_2785);
and U4379 (N_4379,N_114,N_2990);
and U4380 (N_4380,N_130,N_1931);
nand U4381 (N_4381,N_481,N_535);
nor U4382 (N_4382,N_1177,N_2734);
or U4383 (N_4383,N_547,N_268);
or U4384 (N_4384,N_1669,N_2862);
or U4385 (N_4385,N_1089,N_1535);
nand U4386 (N_4386,N_289,N_2460);
and U4387 (N_4387,N_2092,N_1453);
xnor U4388 (N_4388,N_1920,N_1063);
nand U4389 (N_4389,N_2569,N_679);
xnor U4390 (N_4390,N_1169,N_1922);
and U4391 (N_4391,N_2236,N_513);
and U4392 (N_4392,N_2281,N_1257);
or U4393 (N_4393,N_2705,N_138);
and U4394 (N_4394,N_1286,N_2355);
and U4395 (N_4395,N_238,N_2134);
and U4396 (N_4396,N_692,N_1544);
nor U4397 (N_4397,N_2305,N_2401);
nand U4398 (N_4398,N_2027,N_2350);
nand U4399 (N_4399,N_2143,N_1062);
nand U4400 (N_4400,N_2346,N_2911);
nand U4401 (N_4401,N_911,N_1662);
and U4402 (N_4402,N_2837,N_2162);
nor U4403 (N_4403,N_1474,N_1985);
or U4404 (N_4404,N_1709,N_486);
and U4405 (N_4405,N_1377,N_788);
nand U4406 (N_4406,N_1359,N_159);
xor U4407 (N_4407,N_2333,N_1171);
or U4408 (N_4408,N_2272,N_428);
xnor U4409 (N_4409,N_1183,N_2543);
nor U4410 (N_4410,N_2258,N_2598);
xor U4411 (N_4411,N_2459,N_1943);
xor U4412 (N_4412,N_471,N_2235);
or U4413 (N_4413,N_1441,N_2069);
nand U4414 (N_4414,N_964,N_326);
xnor U4415 (N_4415,N_674,N_1691);
xnor U4416 (N_4416,N_2560,N_419);
nor U4417 (N_4417,N_1140,N_636);
or U4418 (N_4418,N_2437,N_2387);
nor U4419 (N_4419,N_670,N_1478);
xnor U4420 (N_4420,N_2565,N_1722);
nor U4421 (N_4421,N_2127,N_2062);
and U4422 (N_4422,N_1738,N_1375);
xor U4423 (N_4423,N_1125,N_1705);
xnor U4424 (N_4424,N_2648,N_922);
xnor U4425 (N_4425,N_2022,N_61);
nor U4426 (N_4426,N_1267,N_1570);
or U4427 (N_4427,N_939,N_2266);
and U4428 (N_4428,N_1630,N_81);
xor U4429 (N_4429,N_2353,N_557);
nor U4430 (N_4430,N_1860,N_1554);
and U4431 (N_4431,N_526,N_1578);
xor U4432 (N_4432,N_1568,N_1214);
nor U4433 (N_4433,N_1897,N_2588);
nor U4434 (N_4434,N_2710,N_372);
nand U4435 (N_4435,N_587,N_2647);
nand U4436 (N_4436,N_2758,N_824);
xnor U4437 (N_4437,N_683,N_311);
nand U4438 (N_4438,N_195,N_1393);
nor U4439 (N_4439,N_1676,N_123);
nor U4440 (N_4440,N_1510,N_1028);
and U4441 (N_4441,N_1124,N_2500);
and U4442 (N_4442,N_420,N_733);
xnor U4443 (N_4443,N_2621,N_678);
or U4444 (N_4444,N_1420,N_2341);
nor U4445 (N_4445,N_2803,N_2748);
xor U4446 (N_4446,N_941,N_2583);
nor U4447 (N_4447,N_589,N_505);
xnor U4448 (N_4448,N_11,N_1247);
and U4449 (N_4449,N_1254,N_949);
nor U4450 (N_4450,N_1951,N_377);
xnor U4451 (N_4451,N_1250,N_1460);
or U4452 (N_4452,N_2444,N_1717);
nor U4453 (N_4453,N_1160,N_2907);
and U4454 (N_4454,N_1392,N_2427);
xor U4455 (N_4455,N_2016,N_2555);
nand U4456 (N_4456,N_404,N_1953);
nor U4457 (N_4457,N_270,N_1678);
and U4458 (N_4458,N_2744,N_575);
xnor U4459 (N_4459,N_2490,N_1981);
nand U4460 (N_4460,N_436,N_2527);
xor U4461 (N_4461,N_175,N_1966);
and U4462 (N_4462,N_887,N_1428);
or U4463 (N_4463,N_2331,N_417);
nor U4464 (N_4464,N_440,N_2704);
or U4465 (N_4465,N_756,N_1715);
xnor U4466 (N_4466,N_1009,N_2627);
xnor U4467 (N_4467,N_2075,N_1300);
and U4468 (N_4468,N_476,N_1496);
nand U4469 (N_4469,N_2547,N_1329);
xnor U4470 (N_4470,N_188,N_812);
nand U4471 (N_4471,N_905,N_2441);
nand U4472 (N_4472,N_110,N_2604);
nor U4473 (N_4473,N_2886,N_1362);
nor U4474 (N_4474,N_2518,N_1852);
and U4475 (N_4475,N_1012,N_1313);
xnor U4476 (N_4476,N_2607,N_401);
or U4477 (N_4477,N_2267,N_602);
or U4478 (N_4478,N_970,N_2482);
or U4479 (N_4479,N_2477,N_1001);
and U4480 (N_4480,N_810,N_896);
nand U4481 (N_4481,N_2193,N_690);
or U4482 (N_4482,N_2300,N_883);
nand U4483 (N_4483,N_497,N_1397);
nor U4484 (N_4484,N_945,N_2072);
nand U4485 (N_4485,N_2989,N_2568);
xnor U4486 (N_4486,N_301,N_2151);
xor U4487 (N_4487,N_1530,N_2425);
nand U4488 (N_4488,N_799,N_2868);
nor U4489 (N_4489,N_2592,N_1648);
or U4490 (N_4490,N_2781,N_512);
nand U4491 (N_4491,N_187,N_1629);
nand U4492 (N_4492,N_189,N_1457);
nand U4493 (N_4493,N_1468,N_986);
and U4494 (N_4494,N_1661,N_2099);
nor U4495 (N_4495,N_2937,N_1995);
xor U4496 (N_4496,N_349,N_69);
and U4497 (N_4497,N_163,N_769);
nor U4498 (N_4498,N_1013,N_2903);
or U4499 (N_4499,N_245,N_791);
nand U4500 (N_4500,N_769,N_2299);
or U4501 (N_4501,N_2697,N_2925);
nor U4502 (N_4502,N_204,N_1623);
and U4503 (N_4503,N_1348,N_2592);
xnor U4504 (N_4504,N_1103,N_1326);
and U4505 (N_4505,N_93,N_1931);
nor U4506 (N_4506,N_2528,N_2542);
or U4507 (N_4507,N_885,N_250);
nor U4508 (N_4508,N_234,N_162);
or U4509 (N_4509,N_2862,N_1861);
xor U4510 (N_4510,N_1068,N_2402);
xor U4511 (N_4511,N_2581,N_334);
xor U4512 (N_4512,N_1044,N_2995);
xor U4513 (N_4513,N_2514,N_1670);
nand U4514 (N_4514,N_52,N_575);
xor U4515 (N_4515,N_1814,N_586);
or U4516 (N_4516,N_1958,N_2018);
or U4517 (N_4517,N_2783,N_2418);
xor U4518 (N_4518,N_1695,N_1091);
xnor U4519 (N_4519,N_943,N_2257);
xnor U4520 (N_4520,N_2858,N_2078);
or U4521 (N_4521,N_1921,N_1928);
or U4522 (N_4522,N_760,N_1687);
or U4523 (N_4523,N_1364,N_538);
xnor U4524 (N_4524,N_2417,N_669);
xnor U4525 (N_4525,N_440,N_1007);
or U4526 (N_4526,N_2628,N_1140);
and U4527 (N_4527,N_870,N_1675);
or U4528 (N_4528,N_2003,N_1136);
and U4529 (N_4529,N_686,N_2722);
and U4530 (N_4530,N_2607,N_1811);
nand U4531 (N_4531,N_1375,N_2113);
nor U4532 (N_4532,N_1016,N_597);
xor U4533 (N_4533,N_1436,N_1128);
nand U4534 (N_4534,N_69,N_1817);
or U4535 (N_4535,N_1397,N_2916);
and U4536 (N_4536,N_1053,N_167);
nor U4537 (N_4537,N_1430,N_1952);
xnor U4538 (N_4538,N_2686,N_1379);
and U4539 (N_4539,N_2066,N_2277);
and U4540 (N_4540,N_1134,N_2887);
nor U4541 (N_4541,N_2302,N_982);
and U4542 (N_4542,N_2416,N_1580);
nand U4543 (N_4543,N_375,N_1029);
nand U4544 (N_4544,N_34,N_2094);
xor U4545 (N_4545,N_2076,N_2262);
or U4546 (N_4546,N_1305,N_2985);
nor U4547 (N_4547,N_409,N_798);
nand U4548 (N_4548,N_2069,N_2036);
and U4549 (N_4549,N_773,N_2377);
xnor U4550 (N_4550,N_2203,N_2167);
and U4551 (N_4551,N_801,N_1094);
xnor U4552 (N_4552,N_1913,N_2947);
xor U4553 (N_4553,N_2371,N_2718);
and U4554 (N_4554,N_1614,N_83);
xor U4555 (N_4555,N_2734,N_2833);
and U4556 (N_4556,N_2633,N_486);
and U4557 (N_4557,N_1498,N_1500);
and U4558 (N_4558,N_1650,N_1323);
nor U4559 (N_4559,N_2333,N_1933);
nand U4560 (N_4560,N_2418,N_432);
nor U4561 (N_4561,N_590,N_1970);
and U4562 (N_4562,N_2277,N_508);
nand U4563 (N_4563,N_73,N_2563);
nor U4564 (N_4564,N_1748,N_163);
nor U4565 (N_4565,N_1550,N_80);
xnor U4566 (N_4566,N_2084,N_28);
and U4567 (N_4567,N_1673,N_1362);
nor U4568 (N_4568,N_1349,N_2702);
xnor U4569 (N_4569,N_2740,N_729);
xnor U4570 (N_4570,N_1400,N_2752);
and U4571 (N_4571,N_867,N_1955);
nand U4572 (N_4572,N_627,N_634);
xnor U4573 (N_4573,N_912,N_1835);
nand U4574 (N_4574,N_19,N_1896);
nor U4575 (N_4575,N_1117,N_1419);
and U4576 (N_4576,N_1033,N_2073);
xor U4577 (N_4577,N_1490,N_486);
nor U4578 (N_4578,N_918,N_2527);
xor U4579 (N_4579,N_262,N_242);
nand U4580 (N_4580,N_1692,N_287);
nand U4581 (N_4581,N_2323,N_232);
and U4582 (N_4582,N_1767,N_1354);
xor U4583 (N_4583,N_1291,N_1154);
nor U4584 (N_4584,N_96,N_561);
xor U4585 (N_4585,N_193,N_505);
nand U4586 (N_4586,N_1565,N_117);
nor U4587 (N_4587,N_286,N_625);
xnor U4588 (N_4588,N_2121,N_366);
and U4589 (N_4589,N_782,N_521);
nand U4590 (N_4590,N_2961,N_273);
nor U4591 (N_4591,N_1943,N_1281);
xnor U4592 (N_4592,N_480,N_1230);
xnor U4593 (N_4593,N_1911,N_257);
and U4594 (N_4594,N_1153,N_145);
nor U4595 (N_4595,N_2708,N_253);
or U4596 (N_4596,N_2158,N_2996);
or U4597 (N_4597,N_1868,N_2526);
or U4598 (N_4598,N_156,N_1810);
and U4599 (N_4599,N_1683,N_2776);
nor U4600 (N_4600,N_848,N_1160);
nor U4601 (N_4601,N_670,N_2159);
nor U4602 (N_4602,N_112,N_226);
xnor U4603 (N_4603,N_2967,N_350);
nor U4604 (N_4604,N_2117,N_1841);
xnor U4605 (N_4605,N_1744,N_1091);
or U4606 (N_4606,N_1841,N_2514);
or U4607 (N_4607,N_2,N_1128);
nand U4608 (N_4608,N_854,N_1880);
nand U4609 (N_4609,N_575,N_508);
or U4610 (N_4610,N_2747,N_1593);
nor U4611 (N_4611,N_595,N_1515);
or U4612 (N_4612,N_1,N_2159);
xnor U4613 (N_4613,N_1830,N_1882);
or U4614 (N_4614,N_1683,N_935);
xnor U4615 (N_4615,N_2391,N_2824);
or U4616 (N_4616,N_1622,N_117);
xor U4617 (N_4617,N_1483,N_270);
or U4618 (N_4618,N_2726,N_2596);
or U4619 (N_4619,N_2077,N_914);
nor U4620 (N_4620,N_2811,N_2169);
or U4621 (N_4621,N_2275,N_2986);
xnor U4622 (N_4622,N_2404,N_1382);
xor U4623 (N_4623,N_2011,N_2785);
xor U4624 (N_4624,N_1050,N_2322);
nor U4625 (N_4625,N_1177,N_2740);
and U4626 (N_4626,N_214,N_2310);
nor U4627 (N_4627,N_1399,N_1943);
or U4628 (N_4628,N_2966,N_1311);
nor U4629 (N_4629,N_166,N_2526);
and U4630 (N_4630,N_673,N_1317);
xor U4631 (N_4631,N_240,N_1232);
xor U4632 (N_4632,N_1974,N_589);
nand U4633 (N_4633,N_2519,N_1654);
nand U4634 (N_4634,N_778,N_653);
or U4635 (N_4635,N_1320,N_240);
and U4636 (N_4636,N_887,N_1536);
and U4637 (N_4637,N_1096,N_2125);
nand U4638 (N_4638,N_1261,N_1733);
or U4639 (N_4639,N_394,N_2929);
nand U4640 (N_4640,N_2872,N_1071);
and U4641 (N_4641,N_485,N_2972);
xor U4642 (N_4642,N_1325,N_2474);
and U4643 (N_4643,N_908,N_1489);
and U4644 (N_4644,N_1836,N_117);
xnor U4645 (N_4645,N_2252,N_2146);
nand U4646 (N_4646,N_1788,N_2336);
nand U4647 (N_4647,N_1349,N_318);
xnor U4648 (N_4648,N_1609,N_2583);
xnor U4649 (N_4649,N_791,N_2450);
and U4650 (N_4650,N_203,N_901);
nor U4651 (N_4651,N_2926,N_2529);
and U4652 (N_4652,N_382,N_1358);
nand U4653 (N_4653,N_1005,N_2066);
and U4654 (N_4654,N_1060,N_668);
xnor U4655 (N_4655,N_2698,N_2214);
or U4656 (N_4656,N_386,N_2174);
nor U4657 (N_4657,N_1685,N_2435);
nand U4658 (N_4658,N_584,N_2306);
xor U4659 (N_4659,N_828,N_1434);
xnor U4660 (N_4660,N_541,N_2787);
xor U4661 (N_4661,N_1239,N_1532);
xor U4662 (N_4662,N_837,N_1997);
and U4663 (N_4663,N_2651,N_1323);
nor U4664 (N_4664,N_409,N_743);
nand U4665 (N_4665,N_2787,N_1806);
and U4666 (N_4666,N_1390,N_2214);
nand U4667 (N_4667,N_1424,N_208);
or U4668 (N_4668,N_294,N_1713);
nand U4669 (N_4669,N_1273,N_1508);
nand U4670 (N_4670,N_625,N_1645);
nor U4671 (N_4671,N_1044,N_214);
nor U4672 (N_4672,N_750,N_2596);
nor U4673 (N_4673,N_289,N_1269);
xor U4674 (N_4674,N_2288,N_2974);
nor U4675 (N_4675,N_1159,N_2827);
and U4676 (N_4676,N_2170,N_1054);
or U4677 (N_4677,N_1676,N_2216);
xnor U4678 (N_4678,N_710,N_2034);
nand U4679 (N_4679,N_350,N_315);
or U4680 (N_4680,N_1417,N_1484);
nor U4681 (N_4681,N_1853,N_1912);
or U4682 (N_4682,N_2728,N_1677);
nand U4683 (N_4683,N_730,N_1295);
or U4684 (N_4684,N_899,N_164);
nor U4685 (N_4685,N_1977,N_644);
and U4686 (N_4686,N_2519,N_2755);
or U4687 (N_4687,N_1127,N_116);
xor U4688 (N_4688,N_2753,N_694);
xnor U4689 (N_4689,N_2343,N_369);
xor U4690 (N_4690,N_613,N_469);
nor U4691 (N_4691,N_1085,N_1690);
nand U4692 (N_4692,N_150,N_2105);
or U4693 (N_4693,N_1398,N_1285);
nor U4694 (N_4694,N_1087,N_1502);
nor U4695 (N_4695,N_2065,N_1895);
or U4696 (N_4696,N_2760,N_2707);
nand U4697 (N_4697,N_2551,N_2473);
or U4698 (N_4698,N_1260,N_2657);
and U4699 (N_4699,N_2708,N_1623);
or U4700 (N_4700,N_841,N_1795);
xnor U4701 (N_4701,N_2936,N_2643);
or U4702 (N_4702,N_1294,N_1069);
xnor U4703 (N_4703,N_2759,N_2069);
or U4704 (N_4704,N_653,N_1538);
or U4705 (N_4705,N_2316,N_1123);
xnor U4706 (N_4706,N_93,N_1626);
and U4707 (N_4707,N_125,N_46);
and U4708 (N_4708,N_1052,N_180);
xor U4709 (N_4709,N_2859,N_2926);
nand U4710 (N_4710,N_1924,N_1443);
nand U4711 (N_4711,N_2590,N_2405);
xor U4712 (N_4712,N_2778,N_2560);
nor U4713 (N_4713,N_2499,N_176);
nand U4714 (N_4714,N_2225,N_200);
nand U4715 (N_4715,N_2165,N_2925);
nor U4716 (N_4716,N_321,N_1106);
xor U4717 (N_4717,N_2211,N_698);
nand U4718 (N_4718,N_2756,N_2326);
or U4719 (N_4719,N_2702,N_2979);
nand U4720 (N_4720,N_2429,N_1296);
nor U4721 (N_4721,N_2871,N_1478);
nor U4722 (N_4722,N_305,N_2804);
nor U4723 (N_4723,N_1156,N_2927);
and U4724 (N_4724,N_30,N_2740);
nand U4725 (N_4725,N_1850,N_1514);
and U4726 (N_4726,N_1474,N_2872);
xor U4727 (N_4727,N_26,N_2001);
and U4728 (N_4728,N_2820,N_2053);
nand U4729 (N_4729,N_301,N_2089);
nor U4730 (N_4730,N_2385,N_2693);
xor U4731 (N_4731,N_1413,N_2925);
xnor U4732 (N_4732,N_1948,N_1081);
nor U4733 (N_4733,N_2878,N_1235);
xor U4734 (N_4734,N_1302,N_1200);
xor U4735 (N_4735,N_581,N_900);
xnor U4736 (N_4736,N_2952,N_105);
nand U4737 (N_4737,N_287,N_163);
xnor U4738 (N_4738,N_678,N_2473);
or U4739 (N_4739,N_914,N_2069);
or U4740 (N_4740,N_539,N_1796);
nand U4741 (N_4741,N_2205,N_2068);
or U4742 (N_4742,N_1877,N_485);
xor U4743 (N_4743,N_1103,N_2763);
xor U4744 (N_4744,N_1548,N_875);
and U4745 (N_4745,N_824,N_1499);
xnor U4746 (N_4746,N_864,N_978);
or U4747 (N_4747,N_1931,N_2709);
nor U4748 (N_4748,N_1536,N_1450);
nand U4749 (N_4749,N_1950,N_2993);
and U4750 (N_4750,N_2356,N_2481);
nand U4751 (N_4751,N_1362,N_2130);
xor U4752 (N_4752,N_111,N_1263);
and U4753 (N_4753,N_576,N_2911);
or U4754 (N_4754,N_1404,N_920);
and U4755 (N_4755,N_2190,N_840);
nor U4756 (N_4756,N_179,N_2083);
nor U4757 (N_4757,N_2377,N_1253);
xnor U4758 (N_4758,N_1513,N_1637);
nand U4759 (N_4759,N_1900,N_336);
and U4760 (N_4760,N_784,N_2679);
nand U4761 (N_4761,N_2110,N_1106);
and U4762 (N_4762,N_1425,N_732);
nand U4763 (N_4763,N_341,N_1559);
and U4764 (N_4764,N_1055,N_161);
nor U4765 (N_4765,N_2245,N_2060);
nand U4766 (N_4766,N_2897,N_1319);
and U4767 (N_4767,N_863,N_2584);
and U4768 (N_4768,N_605,N_506);
nand U4769 (N_4769,N_2592,N_1254);
or U4770 (N_4770,N_2866,N_369);
or U4771 (N_4771,N_2273,N_1844);
or U4772 (N_4772,N_638,N_2673);
xnor U4773 (N_4773,N_22,N_1724);
nand U4774 (N_4774,N_1018,N_2504);
and U4775 (N_4775,N_1582,N_628);
and U4776 (N_4776,N_141,N_2796);
nor U4777 (N_4777,N_1477,N_412);
nor U4778 (N_4778,N_1384,N_2638);
nor U4779 (N_4779,N_265,N_1931);
or U4780 (N_4780,N_450,N_2647);
xor U4781 (N_4781,N_2762,N_1141);
nor U4782 (N_4782,N_463,N_2221);
or U4783 (N_4783,N_2877,N_2077);
or U4784 (N_4784,N_1447,N_2064);
nor U4785 (N_4785,N_2280,N_2655);
nor U4786 (N_4786,N_1457,N_2051);
or U4787 (N_4787,N_2046,N_2061);
nand U4788 (N_4788,N_775,N_171);
nand U4789 (N_4789,N_1008,N_1943);
and U4790 (N_4790,N_1122,N_189);
nor U4791 (N_4791,N_1294,N_656);
or U4792 (N_4792,N_1141,N_2578);
xnor U4793 (N_4793,N_2579,N_2850);
and U4794 (N_4794,N_1763,N_1899);
xor U4795 (N_4795,N_2737,N_743);
or U4796 (N_4796,N_2555,N_1041);
and U4797 (N_4797,N_2563,N_2688);
nand U4798 (N_4798,N_2912,N_497);
nor U4799 (N_4799,N_1610,N_314);
xnor U4800 (N_4800,N_821,N_2896);
or U4801 (N_4801,N_1645,N_1621);
xnor U4802 (N_4802,N_2724,N_1966);
nand U4803 (N_4803,N_962,N_80);
nor U4804 (N_4804,N_1591,N_2081);
xor U4805 (N_4805,N_1243,N_1684);
nand U4806 (N_4806,N_900,N_2714);
and U4807 (N_4807,N_2332,N_2038);
nand U4808 (N_4808,N_550,N_564);
nand U4809 (N_4809,N_557,N_1325);
xnor U4810 (N_4810,N_2518,N_2196);
or U4811 (N_4811,N_2950,N_310);
nor U4812 (N_4812,N_2065,N_691);
nand U4813 (N_4813,N_136,N_873);
and U4814 (N_4814,N_1221,N_476);
and U4815 (N_4815,N_2557,N_2841);
xor U4816 (N_4816,N_106,N_1452);
nand U4817 (N_4817,N_13,N_1553);
and U4818 (N_4818,N_2865,N_1986);
xnor U4819 (N_4819,N_759,N_2181);
nor U4820 (N_4820,N_1091,N_636);
nor U4821 (N_4821,N_209,N_1756);
or U4822 (N_4822,N_145,N_593);
and U4823 (N_4823,N_1177,N_546);
nor U4824 (N_4824,N_1046,N_670);
nor U4825 (N_4825,N_2899,N_924);
nor U4826 (N_4826,N_999,N_2447);
or U4827 (N_4827,N_2539,N_1016);
xnor U4828 (N_4828,N_1160,N_2415);
nand U4829 (N_4829,N_295,N_1708);
nor U4830 (N_4830,N_1678,N_412);
nor U4831 (N_4831,N_2090,N_2129);
or U4832 (N_4832,N_69,N_2172);
nor U4833 (N_4833,N_1669,N_266);
nand U4834 (N_4834,N_2702,N_264);
or U4835 (N_4835,N_601,N_1166);
nand U4836 (N_4836,N_1544,N_367);
and U4837 (N_4837,N_1804,N_2762);
xnor U4838 (N_4838,N_2169,N_559);
and U4839 (N_4839,N_1995,N_1630);
nor U4840 (N_4840,N_319,N_2906);
nand U4841 (N_4841,N_1382,N_1021);
nand U4842 (N_4842,N_62,N_2580);
nand U4843 (N_4843,N_2781,N_2316);
xor U4844 (N_4844,N_1504,N_182);
nor U4845 (N_4845,N_1898,N_2047);
and U4846 (N_4846,N_246,N_1209);
or U4847 (N_4847,N_1619,N_1860);
nand U4848 (N_4848,N_2934,N_2602);
xor U4849 (N_4849,N_2299,N_2381);
nand U4850 (N_4850,N_2361,N_2260);
or U4851 (N_4851,N_1175,N_1);
nand U4852 (N_4852,N_2717,N_1160);
or U4853 (N_4853,N_1757,N_185);
nand U4854 (N_4854,N_1522,N_409);
xnor U4855 (N_4855,N_310,N_2794);
xor U4856 (N_4856,N_668,N_1455);
or U4857 (N_4857,N_2121,N_2113);
nor U4858 (N_4858,N_1270,N_815);
or U4859 (N_4859,N_1,N_2021);
nor U4860 (N_4860,N_168,N_2273);
and U4861 (N_4861,N_7,N_2894);
xor U4862 (N_4862,N_310,N_1193);
nor U4863 (N_4863,N_553,N_1658);
nand U4864 (N_4864,N_1798,N_144);
or U4865 (N_4865,N_2222,N_334);
nor U4866 (N_4866,N_884,N_929);
nand U4867 (N_4867,N_1192,N_1650);
xor U4868 (N_4868,N_2878,N_1636);
nand U4869 (N_4869,N_1815,N_2030);
or U4870 (N_4870,N_949,N_2067);
and U4871 (N_4871,N_407,N_1516);
and U4872 (N_4872,N_1951,N_2998);
nand U4873 (N_4873,N_87,N_1338);
nand U4874 (N_4874,N_2848,N_1088);
xnor U4875 (N_4875,N_130,N_1372);
and U4876 (N_4876,N_2128,N_383);
nand U4877 (N_4877,N_343,N_2748);
nor U4878 (N_4878,N_1350,N_2106);
nor U4879 (N_4879,N_1444,N_1351);
or U4880 (N_4880,N_2028,N_2715);
nor U4881 (N_4881,N_266,N_1542);
nand U4882 (N_4882,N_1320,N_473);
or U4883 (N_4883,N_1305,N_2618);
nor U4884 (N_4884,N_1733,N_673);
xnor U4885 (N_4885,N_1250,N_1388);
nor U4886 (N_4886,N_2169,N_1616);
xnor U4887 (N_4887,N_1086,N_196);
nor U4888 (N_4888,N_1386,N_1840);
nor U4889 (N_4889,N_2501,N_1028);
xnor U4890 (N_4890,N_2678,N_1621);
or U4891 (N_4891,N_2660,N_2093);
nor U4892 (N_4892,N_1694,N_2916);
and U4893 (N_4893,N_2103,N_1614);
and U4894 (N_4894,N_424,N_489);
xnor U4895 (N_4895,N_1546,N_1558);
xnor U4896 (N_4896,N_2754,N_2272);
or U4897 (N_4897,N_2004,N_585);
xor U4898 (N_4898,N_2090,N_1752);
xor U4899 (N_4899,N_246,N_2963);
xor U4900 (N_4900,N_814,N_191);
and U4901 (N_4901,N_1343,N_1251);
nand U4902 (N_4902,N_1673,N_1431);
or U4903 (N_4903,N_1400,N_2539);
or U4904 (N_4904,N_776,N_2328);
nand U4905 (N_4905,N_484,N_2302);
nand U4906 (N_4906,N_2817,N_587);
and U4907 (N_4907,N_2317,N_2177);
or U4908 (N_4908,N_2920,N_966);
and U4909 (N_4909,N_104,N_1290);
nand U4910 (N_4910,N_1353,N_777);
nor U4911 (N_4911,N_21,N_2455);
xor U4912 (N_4912,N_2822,N_2501);
and U4913 (N_4913,N_1686,N_2725);
xor U4914 (N_4914,N_1606,N_395);
or U4915 (N_4915,N_262,N_2520);
and U4916 (N_4916,N_2275,N_2930);
nor U4917 (N_4917,N_587,N_1002);
nor U4918 (N_4918,N_2125,N_1172);
nor U4919 (N_4919,N_1716,N_63);
or U4920 (N_4920,N_2998,N_720);
nor U4921 (N_4921,N_1285,N_2160);
nand U4922 (N_4922,N_670,N_761);
and U4923 (N_4923,N_1729,N_693);
nand U4924 (N_4924,N_1788,N_2576);
nor U4925 (N_4925,N_482,N_2418);
nand U4926 (N_4926,N_1659,N_2488);
nor U4927 (N_4927,N_2885,N_225);
xnor U4928 (N_4928,N_210,N_2575);
or U4929 (N_4929,N_667,N_1926);
xnor U4930 (N_4930,N_1617,N_2323);
xor U4931 (N_4931,N_823,N_2341);
and U4932 (N_4932,N_1092,N_1767);
nand U4933 (N_4933,N_751,N_2316);
xor U4934 (N_4934,N_795,N_1733);
and U4935 (N_4935,N_2796,N_2786);
or U4936 (N_4936,N_2424,N_1505);
xor U4937 (N_4937,N_1290,N_283);
and U4938 (N_4938,N_284,N_1195);
or U4939 (N_4939,N_2316,N_1646);
xor U4940 (N_4940,N_408,N_423);
xor U4941 (N_4941,N_1323,N_1468);
xnor U4942 (N_4942,N_686,N_1213);
nand U4943 (N_4943,N_1710,N_896);
or U4944 (N_4944,N_2256,N_326);
or U4945 (N_4945,N_975,N_1178);
xor U4946 (N_4946,N_2757,N_1823);
xnor U4947 (N_4947,N_1658,N_1199);
and U4948 (N_4948,N_1893,N_2361);
xnor U4949 (N_4949,N_206,N_731);
or U4950 (N_4950,N_1256,N_47);
and U4951 (N_4951,N_322,N_172);
or U4952 (N_4952,N_865,N_2435);
xnor U4953 (N_4953,N_261,N_2048);
or U4954 (N_4954,N_981,N_2284);
nand U4955 (N_4955,N_661,N_2692);
nor U4956 (N_4956,N_1235,N_493);
nand U4957 (N_4957,N_2478,N_1493);
xor U4958 (N_4958,N_1067,N_1142);
and U4959 (N_4959,N_1940,N_1024);
xnor U4960 (N_4960,N_2511,N_845);
xor U4961 (N_4961,N_767,N_2524);
and U4962 (N_4962,N_1889,N_2168);
or U4963 (N_4963,N_93,N_1024);
xor U4964 (N_4964,N_1702,N_2996);
xor U4965 (N_4965,N_1476,N_2954);
or U4966 (N_4966,N_1582,N_208);
nor U4967 (N_4967,N_744,N_1601);
xnor U4968 (N_4968,N_1560,N_1089);
xor U4969 (N_4969,N_1093,N_274);
or U4970 (N_4970,N_984,N_1011);
xnor U4971 (N_4971,N_65,N_220);
and U4972 (N_4972,N_109,N_2157);
nor U4973 (N_4973,N_332,N_2365);
and U4974 (N_4974,N_1511,N_96);
xor U4975 (N_4975,N_1128,N_695);
or U4976 (N_4976,N_1254,N_2482);
nand U4977 (N_4977,N_818,N_1824);
xnor U4978 (N_4978,N_2471,N_859);
or U4979 (N_4979,N_1925,N_2919);
nand U4980 (N_4980,N_655,N_1597);
nand U4981 (N_4981,N_2060,N_2131);
nand U4982 (N_4982,N_773,N_957);
nor U4983 (N_4983,N_1719,N_2832);
nand U4984 (N_4984,N_2303,N_251);
or U4985 (N_4985,N_1272,N_1215);
or U4986 (N_4986,N_2669,N_872);
and U4987 (N_4987,N_1197,N_2449);
and U4988 (N_4988,N_282,N_2942);
nand U4989 (N_4989,N_2653,N_351);
and U4990 (N_4990,N_2648,N_579);
or U4991 (N_4991,N_1816,N_1990);
xor U4992 (N_4992,N_858,N_951);
nor U4993 (N_4993,N_199,N_1650);
and U4994 (N_4994,N_1697,N_2289);
nand U4995 (N_4995,N_2609,N_2789);
nand U4996 (N_4996,N_322,N_1665);
or U4997 (N_4997,N_650,N_2984);
or U4998 (N_4998,N_1393,N_985);
xor U4999 (N_4999,N_711,N_2810);
nor U5000 (N_5000,N_1601,N_947);
nand U5001 (N_5001,N_2201,N_1949);
nand U5002 (N_5002,N_2319,N_16);
xnor U5003 (N_5003,N_1882,N_2941);
and U5004 (N_5004,N_337,N_1197);
and U5005 (N_5005,N_1959,N_628);
and U5006 (N_5006,N_646,N_101);
nand U5007 (N_5007,N_844,N_2533);
xor U5008 (N_5008,N_2810,N_2594);
and U5009 (N_5009,N_1634,N_2027);
and U5010 (N_5010,N_443,N_1946);
nor U5011 (N_5011,N_1726,N_2758);
xor U5012 (N_5012,N_2931,N_994);
nor U5013 (N_5013,N_1974,N_1572);
nor U5014 (N_5014,N_509,N_1530);
and U5015 (N_5015,N_2137,N_1188);
or U5016 (N_5016,N_1992,N_2600);
or U5017 (N_5017,N_837,N_2135);
or U5018 (N_5018,N_362,N_1026);
nand U5019 (N_5019,N_2803,N_730);
nor U5020 (N_5020,N_392,N_1750);
xnor U5021 (N_5021,N_29,N_2806);
and U5022 (N_5022,N_65,N_277);
or U5023 (N_5023,N_2504,N_2276);
and U5024 (N_5024,N_162,N_2238);
nand U5025 (N_5025,N_1545,N_2325);
or U5026 (N_5026,N_2370,N_1927);
nor U5027 (N_5027,N_1900,N_1127);
nor U5028 (N_5028,N_2645,N_1892);
and U5029 (N_5029,N_2583,N_875);
xor U5030 (N_5030,N_494,N_1533);
nand U5031 (N_5031,N_1541,N_2812);
or U5032 (N_5032,N_235,N_1779);
nor U5033 (N_5033,N_1268,N_2716);
xnor U5034 (N_5034,N_1680,N_1167);
xnor U5035 (N_5035,N_1710,N_1316);
nand U5036 (N_5036,N_1448,N_831);
and U5037 (N_5037,N_1549,N_1053);
and U5038 (N_5038,N_1627,N_2612);
xor U5039 (N_5039,N_2774,N_1104);
xor U5040 (N_5040,N_537,N_1538);
xnor U5041 (N_5041,N_2750,N_225);
nor U5042 (N_5042,N_1374,N_2390);
xor U5043 (N_5043,N_103,N_1510);
nand U5044 (N_5044,N_1400,N_2748);
or U5045 (N_5045,N_443,N_987);
nand U5046 (N_5046,N_2443,N_1035);
and U5047 (N_5047,N_114,N_2172);
and U5048 (N_5048,N_1801,N_1783);
nand U5049 (N_5049,N_2209,N_2212);
xor U5050 (N_5050,N_1031,N_1216);
nand U5051 (N_5051,N_1961,N_1118);
xnor U5052 (N_5052,N_1285,N_1424);
or U5053 (N_5053,N_1605,N_771);
and U5054 (N_5054,N_700,N_781);
or U5055 (N_5055,N_1200,N_2252);
nand U5056 (N_5056,N_1272,N_2171);
or U5057 (N_5057,N_1661,N_2730);
xor U5058 (N_5058,N_1058,N_2925);
and U5059 (N_5059,N_314,N_31);
nand U5060 (N_5060,N_2643,N_1822);
and U5061 (N_5061,N_1801,N_1232);
or U5062 (N_5062,N_2384,N_2192);
xnor U5063 (N_5063,N_2111,N_2554);
or U5064 (N_5064,N_210,N_2908);
nor U5065 (N_5065,N_598,N_26);
or U5066 (N_5066,N_2580,N_2665);
nor U5067 (N_5067,N_2962,N_1089);
or U5068 (N_5068,N_2266,N_36);
and U5069 (N_5069,N_257,N_583);
nor U5070 (N_5070,N_530,N_1149);
nand U5071 (N_5071,N_922,N_2509);
and U5072 (N_5072,N_339,N_1241);
and U5073 (N_5073,N_634,N_2391);
xnor U5074 (N_5074,N_695,N_335);
xor U5075 (N_5075,N_2375,N_455);
nand U5076 (N_5076,N_2326,N_685);
nand U5077 (N_5077,N_662,N_2904);
nor U5078 (N_5078,N_1718,N_1850);
and U5079 (N_5079,N_1675,N_11);
xor U5080 (N_5080,N_1752,N_1875);
xnor U5081 (N_5081,N_1809,N_252);
or U5082 (N_5082,N_2825,N_1387);
xnor U5083 (N_5083,N_1976,N_2726);
xnor U5084 (N_5084,N_2424,N_1572);
nand U5085 (N_5085,N_1790,N_1680);
nand U5086 (N_5086,N_794,N_373);
or U5087 (N_5087,N_276,N_936);
nor U5088 (N_5088,N_882,N_1547);
nor U5089 (N_5089,N_2083,N_2367);
nand U5090 (N_5090,N_2727,N_2572);
and U5091 (N_5091,N_1375,N_2724);
and U5092 (N_5092,N_293,N_1287);
xor U5093 (N_5093,N_230,N_2496);
nor U5094 (N_5094,N_1892,N_1481);
and U5095 (N_5095,N_554,N_325);
and U5096 (N_5096,N_1240,N_1366);
nor U5097 (N_5097,N_2081,N_2310);
xor U5098 (N_5098,N_841,N_433);
xor U5099 (N_5099,N_1150,N_2980);
or U5100 (N_5100,N_2010,N_467);
xor U5101 (N_5101,N_287,N_1329);
xnor U5102 (N_5102,N_1099,N_158);
nor U5103 (N_5103,N_1159,N_1408);
nor U5104 (N_5104,N_2774,N_1223);
or U5105 (N_5105,N_1047,N_56);
xnor U5106 (N_5106,N_2727,N_1604);
nor U5107 (N_5107,N_2108,N_2867);
nor U5108 (N_5108,N_69,N_1283);
xor U5109 (N_5109,N_1797,N_1628);
xnor U5110 (N_5110,N_485,N_1615);
nand U5111 (N_5111,N_495,N_972);
nand U5112 (N_5112,N_430,N_1750);
xor U5113 (N_5113,N_2245,N_2571);
or U5114 (N_5114,N_2673,N_2458);
and U5115 (N_5115,N_944,N_612);
nand U5116 (N_5116,N_1024,N_804);
or U5117 (N_5117,N_98,N_363);
xor U5118 (N_5118,N_1151,N_2633);
nor U5119 (N_5119,N_1599,N_1508);
or U5120 (N_5120,N_2434,N_1712);
xor U5121 (N_5121,N_94,N_4);
nor U5122 (N_5122,N_1414,N_1164);
xor U5123 (N_5123,N_1141,N_1175);
nand U5124 (N_5124,N_1775,N_234);
or U5125 (N_5125,N_693,N_41);
xor U5126 (N_5126,N_1437,N_1685);
xnor U5127 (N_5127,N_2747,N_1886);
or U5128 (N_5128,N_2350,N_100);
or U5129 (N_5129,N_2837,N_1400);
and U5130 (N_5130,N_1594,N_2821);
nand U5131 (N_5131,N_1548,N_266);
xnor U5132 (N_5132,N_561,N_2187);
or U5133 (N_5133,N_2149,N_2128);
nor U5134 (N_5134,N_2201,N_1647);
nor U5135 (N_5135,N_2053,N_1184);
nand U5136 (N_5136,N_587,N_1754);
xor U5137 (N_5137,N_190,N_2048);
nand U5138 (N_5138,N_84,N_1614);
or U5139 (N_5139,N_2411,N_546);
nand U5140 (N_5140,N_158,N_901);
xnor U5141 (N_5141,N_2397,N_610);
and U5142 (N_5142,N_529,N_914);
nand U5143 (N_5143,N_584,N_1433);
or U5144 (N_5144,N_1676,N_2645);
or U5145 (N_5145,N_1798,N_2246);
and U5146 (N_5146,N_170,N_1445);
or U5147 (N_5147,N_154,N_698);
xnor U5148 (N_5148,N_1272,N_1740);
xor U5149 (N_5149,N_2291,N_2565);
or U5150 (N_5150,N_1932,N_874);
nand U5151 (N_5151,N_2976,N_551);
xnor U5152 (N_5152,N_1423,N_1631);
and U5153 (N_5153,N_2339,N_2326);
or U5154 (N_5154,N_2375,N_2476);
xnor U5155 (N_5155,N_2875,N_851);
nor U5156 (N_5156,N_2614,N_2675);
or U5157 (N_5157,N_1997,N_1578);
xor U5158 (N_5158,N_2724,N_136);
nor U5159 (N_5159,N_1363,N_1726);
or U5160 (N_5160,N_1854,N_220);
and U5161 (N_5161,N_797,N_2478);
nor U5162 (N_5162,N_2044,N_463);
xnor U5163 (N_5163,N_1205,N_1869);
and U5164 (N_5164,N_802,N_1564);
or U5165 (N_5165,N_461,N_679);
or U5166 (N_5166,N_1239,N_1226);
and U5167 (N_5167,N_1753,N_1401);
xnor U5168 (N_5168,N_1251,N_1244);
nor U5169 (N_5169,N_2625,N_1485);
nand U5170 (N_5170,N_1539,N_620);
xnor U5171 (N_5171,N_348,N_1864);
nor U5172 (N_5172,N_573,N_1485);
nor U5173 (N_5173,N_666,N_2917);
or U5174 (N_5174,N_2054,N_647);
or U5175 (N_5175,N_1825,N_2911);
xnor U5176 (N_5176,N_2993,N_1357);
xor U5177 (N_5177,N_2505,N_1648);
nor U5178 (N_5178,N_2161,N_596);
and U5179 (N_5179,N_2061,N_807);
and U5180 (N_5180,N_1665,N_947);
and U5181 (N_5181,N_1701,N_2826);
nand U5182 (N_5182,N_2791,N_2388);
or U5183 (N_5183,N_1231,N_250);
or U5184 (N_5184,N_1704,N_2964);
or U5185 (N_5185,N_1620,N_2503);
nand U5186 (N_5186,N_2998,N_196);
nand U5187 (N_5187,N_2888,N_2209);
or U5188 (N_5188,N_364,N_2326);
nor U5189 (N_5189,N_1095,N_1322);
nand U5190 (N_5190,N_2443,N_208);
nand U5191 (N_5191,N_1403,N_343);
xnor U5192 (N_5192,N_521,N_2185);
nor U5193 (N_5193,N_1447,N_172);
nor U5194 (N_5194,N_2734,N_2945);
nand U5195 (N_5195,N_1811,N_1596);
nand U5196 (N_5196,N_2741,N_601);
xor U5197 (N_5197,N_307,N_32);
or U5198 (N_5198,N_2288,N_2350);
or U5199 (N_5199,N_1788,N_2442);
nand U5200 (N_5200,N_948,N_66);
and U5201 (N_5201,N_738,N_1695);
xor U5202 (N_5202,N_867,N_2872);
nand U5203 (N_5203,N_810,N_275);
xor U5204 (N_5204,N_1588,N_1926);
and U5205 (N_5205,N_651,N_2152);
or U5206 (N_5206,N_283,N_2262);
or U5207 (N_5207,N_2314,N_553);
or U5208 (N_5208,N_2898,N_102);
or U5209 (N_5209,N_1966,N_2756);
xor U5210 (N_5210,N_594,N_2338);
and U5211 (N_5211,N_361,N_2480);
xor U5212 (N_5212,N_1121,N_1159);
nor U5213 (N_5213,N_1987,N_804);
xnor U5214 (N_5214,N_573,N_2596);
nand U5215 (N_5215,N_2207,N_1923);
nand U5216 (N_5216,N_1494,N_676);
nand U5217 (N_5217,N_1128,N_71);
nor U5218 (N_5218,N_2987,N_511);
nor U5219 (N_5219,N_1936,N_1294);
nor U5220 (N_5220,N_276,N_2346);
and U5221 (N_5221,N_2876,N_2365);
xnor U5222 (N_5222,N_1322,N_1664);
and U5223 (N_5223,N_1852,N_1225);
or U5224 (N_5224,N_543,N_297);
and U5225 (N_5225,N_1559,N_267);
nor U5226 (N_5226,N_1078,N_121);
and U5227 (N_5227,N_2557,N_1621);
or U5228 (N_5228,N_87,N_2374);
xnor U5229 (N_5229,N_195,N_629);
and U5230 (N_5230,N_1847,N_738);
nor U5231 (N_5231,N_1793,N_2029);
nor U5232 (N_5232,N_2234,N_1351);
nor U5233 (N_5233,N_791,N_1784);
and U5234 (N_5234,N_248,N_2782);
xor U5235 (N_5235,N_2237,N_1693);
and U5236 (N_5236,N_2874,N_97);
or U5237 (N_5237,N_1160,N_517);
and U5238 (N_5238,N_58,N_2431);
nor U5239 (N_5239,N_209,N_1604);
or U5240 (N_5240,N_776,N_2289);
or U5241 (N_5241,N_170,N_2335);
nand U5242 (N_5242,N_1121,N_1506);
nor U5243 (N_5243,N_2938,N_158);
or U5244 (N_5244,N_2913,N_2942);
and U5245 (N_5245,N_2733,N_1739);
nand U5246 (N_5246,N_867,N_988);
and U5247 (N_5247,N_1746,N_2602);
xnor U5248 (N_5248,N_272,N_117);
nand U5249 (N_5249,N_768,N_560);
and U5250 (N_5250,N_601,N_2398);
nor U5251 (N_5251,N_1676,N_200);
and U5252 (N_5252,N_2230,N_309);
nand U5253 (N_5253,N_2319,N_250);
xnor U5254 (N_5254,N_585,N_2267);
nor U5255 (N_5255,N_436,N_138);
and U5256 (N_5256,N_1930,N_737);
xnor U5257 (N_5257,N_716,N_1496);
and U5258 (N_5258,N_1774,N_731);
nor U5259 (N_5259,N_1469,N_1939);
or U5260 (N_5260,N_279,N_496);
or U5261 (N_5261,N_2093,N_1806);
or U5262 (N_5262,N_721,N_1577);
nor U5263 (N_5263,N_768,N_2112);
nor U5264 (N_5264,N_817,N_1479);
xor U5265 (N_5265,N_524,N_243);
xor U5266 (N_5266,N_2518,N_597);
nand U5267 (N_5267,N_203,N_1486);
or U5268 (N_5268,N_228,N_775);
xor U5269 (N_5269,N_1889,N_1958);
and U5270 (N_5270,N_2155,N_607);
nand U5271 (N_5271,N_1415,N_1041);
and U5272 (N_5272,N_1682,N_1635);
and U5273 (N_5273,N_1078,N_1839);
nor U5274 (N_5274,N_211,N_2084);
xor U5275 (N_5275,N_2494,N_2399);
nor U5276 (N_5276,N_1031,N_826);
nand U5277 (N_5277,N_2482,N_2010);
nor U5278 (N_5278,N_2103,N_2322);
nor U5279 (N_5279,N_1376,N_338);
xnor U5280 (N_5280,N_1324,N_323);
nor U5281 (N_5281,N_1405,N_2381);
nand U5282 (N_5282,N_1998,N_1866);
and U5283 (N_5283,N_858,N_1757);
xnor U5284 (N_5284,N_1911,N_1077);
nand U5285 (N_5285,N_20,N_1724);
xnor U5286 (N_5286,N_1231,N_2683);
nor U5287 (N_5287,N_256,N_2343);
xor U5288 (N_5288,N_1192,N_1437);
nand U5289 (N_5289,N_784,N_2519);
nor U5290 (N_5290,N_1626,N_2559);
and U5291 (N_5291,N_1955,N_2343);
or U5292 (N_5292,N_1926,N_1974);
and U5293 (N_5293,N_26,N_2668);
and U5294 (N_5294,N_1937,N_1266);
nand U5295 (N_5295,N_84,N_2538);
nand U5296 (N_5296,N_2024,N_2936);
nor U5297 (N_5297,N_1152,N_968);
xor U5298 (N_5298,N_2419,N_2730);
nor U5299 (N_5299,N_1622,N_2100);
and U5300 (N_5300,N_626,N_2205);
xnor U5301 (N_5301,N_1060,N_2745);
or U5302 (N_5302,N_1605,N_534);
nor U5303 (N_5303,N_1215,N_2889);
nand U5304 (N_5304,N_2492,N_2648);
nor U5305 (N_5305,N_170,N_2105);
and U5306 (N_5306,N_522,N_2941);
xor U5307 (N_5307,N_1006,N_1588);
nor U5308 (N_5308,N_581,N_2748);
or U5309 (N_5309,N_219,N_1063);
nand U5310 (N_5310,N_2142,N_928);
nand U5311 (N_5311,N_620,N_1641);
nor U5312 (N_5312,N_196,N_2558);
nor U5313 (N_5313,N_2389,N_2256);
nand U5314 (N_5314,N_1677,N_701);
and U5315 (N_5315,N_1112,N_1235);
xnor U5316 (N_5316,N_1557,N_377);
and U5317 (N_5317,N_1170,N_25);
and U5318 (N_5318,N_218,N_2872);
nor U5319 (N_5319,N_228,N_204);
nor U5320 (N_5320,N_1727,N_2494);
xnor U5321 (N_5321,N_2360,N_247);
nand U5322 (N_5322,N_57,N_886);
xor U5323 (N_5323,N_2326,N_1801);
and U5324 (N_5324,N_2701,N_83);
xor U5325 (N_5325,N_2849,N_404);
nand U5326 (N_5326,N_700,N_611);
nand U5327 (N_5327,N_2603,N_654);
and U5328 (N_5328,N_1017,N_573);
nand U5329 (N_5329,N_1498,N_1280);
and U5330 (N_5330,N_1672,N_1995);
or U5331 (N_5331,N_2595,N_634);
or U5332 (N_5332,N_1905,N_851);
nand U5333 (N_5333,N_181,N_360);
xor U5334 (N_5334,N_1899,N_122);
and U5335 (N_5335,N_1894,N_781);
nand U5336 (N_5336,N_2141,N_747);
and U5337 (N_5337,N_1984,N_1282);
and U5338 (N_5338,N_1556,N_2641);
nand U5339 (N_5339,N_574,N_2484);
nand U5340 (N_5340,N_405,N_2442);
or U5341 (N_5341,N_2827,N_1145);
xor U5342 (N_5342,N_299,N_1347);
and U5343 (N_5343,N_2859,N_2447);
or U5344 (N_5344,N_2178,N_649);
or U5345 (N_5345,N_652,N_1042);
nor U5346 (N_5346,N_2040,N_1379);
or U5347 (N_5347,N_2635,N_1575);
nand U5348 (N_5348,N_2648,N_2903);
and U5349 (N_5349,N_1060,N_810);
xor U5350 (N_5350,N_606,N_1524);
or U5351 (N_5351,N_21,N_2856);
nor U5352 (N_5352,N_2614,N_2058);
xnor U5353 (N_5353,N_1085,N_113);
or U5354 (N_5354,N_1580,N_401);
nor U5355 (N_5355,N_2192,N_2059);
nand U5356 (N_5356,N_859,N_2080);
nor U5357 (N_5357,N_2224,N_722);
or U5358 (N_5358,N_1934,N_1226);
and U5359 (N_5359,N_57,N_1681);
xnor U5360 (N_5360,N_1557,N_335);
and U5361 (N_5361,N_131,N_1944);
nand U5362 (N_5362,N_1802,N_2193);
and U5363 (N_5363,N_2957,N_660);
nor U5364 (N_5364,N_1955,N_2510);
or U5365 (N_5365,N_1687,N_476);
or U5366 (N_5366,N_2236,N_2936);
and U5367 (N_5367,N_1236,N_1486);
or U5368 (N_5368,N_396,N_552);
and U5369 (N_5369,N_1479,N_1120);
and U5370 (N_5370,N_1168,N_2246);
and U5371 (N_5371,N_2533,N_67);
nor U5372 (N_5372,N_2114,N_2646);
nand U5373 (N_5373,N_107,N_1122);
nor U5374 (N_5374,N_1683,N_2859);
or U5375 (N_5375,N_2126,N_1258);
and U5376 (N_5376,N_116,N_2329);
or U5377 (N_5377,N_654,N_1002);
nor U5378 (N_5378,N_1900,N_2871);
or U5379 (N_5379,N_1657,N_789);
nand U5380 (N_5380,N_1514,N_2430);
nor U5381 (N_5381,N_1458,N_2734);
xor U5382 (N_5382,N_693,N_1759);
xnor U5383 (N_5383,N_686,N_153);
or U5384 (N_5384,N_1104,N_1650);
and U5385 (N_5385,N_1909,N_634);
nor U5386 (N_5386,N_2700,N_1053);
and U5387 (N_5387,N_2745,N_443);
xnor U5388 (N_5388,N_1259,N_2415);
xnor U5389 (N_5389,N_1702,N_2730);
and U5390 (N_5390,N_1144,N_2042);
or U5391 (N_5391,N_1775,N_1604);
or U5392 (N_5392,N_452,N_2273);
and U5393 (N_5393,N_2643,N_520);
and U5394 (N_5394,N_2167,N_239);
nand U5395 (N_5395,N_336,N_1216);
or U5396 (N_5396,N_1740,N_1176);
xnor U5397 (N_5397,N_43,N_1008);
and U5398 (N_5398,N_2570,N_2647);
or U5399 (N_5399,N_2350,N_1851);
nand U5400 (N_5400,N_1055,N_881);
and U5401 (N_5401,N_2331,N_1037);
nor U5402 (N_5402,N_2449,N_970);
nand U5403 (N_5403,N_1767,N_2667);
nor U5404 (N_5404,N_2059,N_226);
nor U5405 (N_5405,N_2460,N_1106);
nand U5406 (N_5406,N_1943,N_651);
nor U5407 (N_5407,N_1558,N_2403);
and U5408 (N_5408,N_1875,N_1627);
and U5409 (N_5409,N_115,N_2974);
or U5410 (N_5410,N_1396,N_309);
or U5411 (N_5411,N_526,N_1796);
xnor U5412 (N_5412,N_2290,N_97);
xor U5413 (N_5413,N_1690,N_2560);
nor U5414 (N_5414,N_429,N_2784);
nor U5415 (N_5415,N_1021,N_528);
xor U5416 (N_5416,N_2611,N_1951);
and U5417 (N_5417,N_2491,N_687);
and U5418 (N_5418,N_1381,N_286);
nand U5419 (N_5419,N_990,N_2293);
xnor U5420 (N_5420,N_1563,N_1003);
nand U5421 (N_5421,N_1863,N_510);
nor U5422 (N_5422,N_1614,N_1044);
nor U5423 (N_5423,N_1334,N_654);
nor U5424 (N_5424,N_279,N_293);
or U5425 (N_5425,N_1574,N_232);
xor U5426 (N_5426,N_2696,N_2986);
nor U5427 (N_5427,N_1138,N_625);
nor U5428 (N_5428,N_2636,N_942);
nand U5429 (N_5429,N_2140,N_2612);
xnor U5430 (N_5430,N_255,N_2758);
or U5431 (N_5431,N_826,N_440);
xor U5432 (N_5432,N_2968,N_405);
nand U5433 (N_5433,N_1031,N_2586);
xnor U5434 (N_5434,N_1769,N_428);
xor U5435 (N_5435,N_560,N_2301);
or U5436 (N_5436,N_1995,N_2613);
and U5437 (N_5437,N_2065,N_3);
nor U5438 (N_5438,N_1794,N_1297);
nor U5439 (N_5439,N_235,N_1157);
nand U5440 (N_5440,N_2232,N_669);
nand U5441 (N_5441,N_2763,N_2858);
nor U5442 (N_5442,N_2537,N_2643);
and U5443 (N_5443,N_97,N_1016);
or U5444 (N_5444,N_2276,N_689);
xnor U5445 (N_5445,N_1602,N_293);
or U5446 (N_5446,N_2338,N_1337);
nand U5447 (N_5447,N_2168,N_552);
and U5448 (N_5448,N_2022,N_2146);
and U5449 (N_5449,N_1964,N_1624);
and U5450 (N_5450,N_1907,N_118);
xor U5451 (N_5451,N_1786,N_618);
xnor U5452 (N_5452,N_2726,N_526);
nand U5453 (N_5453,N_23,N_2917);
xnor U5454 (N_5454,N_2037,N_1549);
or U5455 (N_5455,N_8,N_1811);
nand U5456 (N_5456,N_1066,N_855);
and U5457 (N_5457,N_2924,N_1319);
and U5458 (N_5458,N_1884,N_543);
or U5459 (N_5459,N_1517,N_2406);
or U5460 (N_5460,N_1928,N_1454);
nor U5461 (N_5461,N_2489,N_315);
nand U5462 (N_5462,N_261,N_205);
nand U5463 (N_5463,N_756,N_2387);
xnor U5464 (N_5464,N_2567,N_1216);
nand U5465 (N_5465,N_694,N_2511);
xnor U5466 (N_5466,N_266,N_2451);
and U5467 (N_5467,N_31,N_2113);
nand U5468 (N_5468,N_2305,N_1993);
or U5469 (N_5469,N_1187,N_689);
nor U5470 (N_5470,N_374,N_378);
and U5471 (N_5471,N_2829,N_1648);
nand U5472 (N_5472,N_1096,N_1523);
nand U5473 (N_5473,N_1005,N_516);
xor U5474 (N_5474,N_1079,N_1306);
nand U5475 (N_5475,N_2154,N_735);
and U5476 (N_5476,N_2519,N_2174);
or U5477 (N_5477,N_202,N_2628);
or U5478 (N_5478,N_547,N_796);
or U5479 (N_5479,N_1636,N_1171);
xor U5480 (N_5480,N_2735,N_824);
or U5481 (N_5481,N_1762,N_367);
nand U5482 (N_5482,N_1449,N_1858);
nor U5483 (N_5483,N_1285,N_1737);
nor U5484 (N_5484,N_2442,N_1295);
or U5485 (N_5485,N_2016,N_443);
or U5486 (N_5486,N_791,N_475);
and U5487 (N_5487,N_1933,N_2410);
nor U5488 (N_5488,N_1976,N_398);
and U5489 (N_5489,N_2130,N_1196);
xnor U5490 (N_5490,N_466,N_2288);
xnor U5491 (N_5491,N_2372,N_2258);
and U5492 (N_5492,N_616,N_1600);
xor U5493 (N_5493,N_2446,N_1583);
xor U5494 (N_5494,N_53,N_1397);
xnor U5495 (N_5495,N_2521,N_1233);
nor U5496 (N_5496,N_1749,N_2970);
nand U5497 (N_5497,N_1564,N_2430);
or U5498 (N_5498,N_2805,N_471);
nor U5499 (N_5499,N_142,N_1717);
xor U5500 (N_5500,N_932,N_1717);
nand U5501 (N_5501,N_2261,N_2808);
or U5502 (N_5502,N_623,N_2603);
and U5503 (N_5503,N_26,N_185);
and U5504 (N_5504,N_1003,N_1909);
nor U5505 (N_5505,N_1967,N_345);
nand U5506 (N_5506,N_787,N_387);
nand U5507 (N_5507,N_578,N_2268);
and U5508 (N_5508,N_567,N_874);
or U5509 (N_5509,N_2455,N_1125);
or U5510 (N_5510,N_1586,N_2413);
and U5511 (N_5511,N_154,N_895);
nor U5512 (N_5512,N_2555,N_289);
or U5513 (N_5513,N_504,N_1515);
or U5514 (N_5514,N_2663,N_2547);
and U5515 (N_5515,N_181,N_726);
xor U5516 (N_5516,N_1983,N_2402);
nor U5517 (N_5517,N_2069,N_1286);
and U5518 (N_5518,N_770,N_1855);
nand U5519 (N_5519,N_2531,N_2173);
nand U5520 (N_5520,N_1466,N_1285);
or U5521 (N_5521,N_1967,N_1035);
nor U5522 (N_5522,N_1173,N_1058);
xnor U5523 (N_5523,N_1082,N_357);
or U5524 (N_5524,N_1574,N_2161);
or U5525 (N_5525,N_590,N_794);
and U5526 (N_5526,N_1808,N_1447);
xor U5527 (N_5527,N_2281,N_2307);
and U5528 (N_5528,N_2077,N_2620);
xor U5529 (N_5529,N_1995,N_981);
and U5530 (N_5530,N_1761,N_235);
nand U5531 (N_5531,N_1848,N_1861);
nand U5532 (N_5532,N_1353,N_882);
and U5533 (N_5533,N_445,N_2295);
nand U5534 (N_5534,N_1781,N_987);
xnor U5535 (N_5535,N_707,N_1243);
and U5536 (N_5536,N_2309,N_2594);
nor U5537 (N_5537,N_1537,N_1917);
nand U5538 (N_5538,N_47,N_2388);
and U5539 (N_5539,N_2060,N_408);
or U5540 (N_5540,N_1525,N_545);
xnor U5541 (N_5541,N_420,N_120);
or U5542 (N_5542,N_2326,N_204);
nand U5543 (N_5543,N_1831,N_1389);
nor U5544 (N_5544,N_1349,N_210);
nor U5545 (N_5545,N_1503,N_1902);
nor U5546 (N_5546,N_941,N_1125);
nand U5547 (N_5547,N_1487,N_980);
xnor U5548 (N_5548,N_2117,N_2108);
nand U5549 (N_5549,N_2402,N_278);
nor U5550 (N_5550,N_1315,N_763);
xor U5551 (N_5551,N_1976,N_2922);
nand U5552 (N_5552,N_1040,N_191);
nor U5553 (N_5553,N_1268,N_2966);
nor U5554 (N_5554,N_890,N_810);
or U5555 (N_5555,N_2712,N_2740);
nor U5556 (N_5556,N_1000,N_2472);
or U5557 (N_5557,N_1712,N_2754);
nand U5558 (N_5558,N_2763,N_1980);
nor U5559 (N_5559,N_308,N_603);
or U5560 (N_5560,N_136,N_1649);
nor U5561 (N_5561,N_2928,N_1259);
and U5562 (N_5562,N_1425,N_2450);
xor U5563 (N_5563,N_922,N_1578);
and U5564 (N_5564,N_1884,N_2614);
and U5565 (N_5565,N_2788,N_1640);
or U5566 (N_5566,N_981,N_812);
xor U5567 (N_5567,N_478,N_2923);
or U5568 (N_5568,N_2049,N_1185);
nor U5569 (N_5569,N_2208,N_663);
and U5570 (N_5570,N_1498,N_2285);
nand U5571 (N_5571,N_1811,N_2779);
nor U5572 (N_5572,N_947,N_2634);
xnor U5573 (N_5573,N_1685,N_1502);
nor U5574 (N_5574,N_2606,N_1739);
nor U5575 (N_5575,N_1627,N_1749);
nor U5576 (N_5576,N_821,N_1426);
or U5577 (N_5577,N_2551,N_298);
xnor U5578 (N_5578,N_761,N_2376);
or U5579 (N_5579,N_1803,N_1462);
nor U5580 (N_5580,N_415,N_2654);
nor U5581 (N_5581,N_744,N_471);
nand U5582 (N_5582,N_1006,N_1482);
nand U5583 (N_5583,N_2192,N_1843);
or U5584 (N_5584,N_2287,N_758);
nand U5585 (N_5585,N_2506,N_2513);
nand U5586 (N_5586,N_2325,N_194);
and U5587 (N_5587,N_395,N_1882);
xor U5588 (N_5588,N_1026,N_2376);
nand U5589 (N_5589,N_2366,N_226);
nor U5590 (N_5590,N_295,N_1888);
and U5591 (N_5591,N_791,N_812);
nor U5592 (N_5592,N_1086,N_2418);
xnor U5593 (N_5593,N_2948,N_2199);
xor U5594 (N_5594,N_2061,N_1943);
or U5595 (N_5595,N_1080,N_695);
and U5596 (N_5596,N_2756,N_62);
or U5597 (N_5597,N_414,N_446);
nor U5598 (N_5598,N_2999,N_1126);
xnor U5599 (N_5599,N_2435,N_1307);
or U5600 (N_5600,N_2906,N_233);
nand U5601 (N_5601,N_81,N_2981);
nor U5602 (N_5602,N_1265,N_1624);
xnor U5603 (N_5603,N_218,N_1390);
nand U5604 (N_5604,N_742,N_453);
or U5605 (N_5605,N_1130,N_659);
nand U5606 (N_5606,N_2379,N_2167);
xnor U5607 (N_5607,N_763,N_1113);
nand U5608 (N_5608,N_2232,N_2342);
xor U5609 (N_5609,N_598,N_45);
and U5610 (N_5610,N_2061,N_1167);
nor U5611 (N_5611,N_120,N_2562);
and U5612 (N_5612,N_2907,N_2879);
or U5613 (N_5613,N_676,N_2968);
or U5614 (N_5614,N_999,N_2750);
and U5615 (N_5615,N_543,N_2808);
and U5616 (N_5616,N_301,N_2096);
and U5617 (N_5617,N_2784,N_373);
nand U5618 (N_5618,N_592,N_783);
nand U5619 (N_5619,N_484,N_2830);
and U5620 (N_5620,N_2164,N_578);
nor U5621 (N_5621,N_1408,N_2499);
nor U5622 (N_5622,N_785,N_2375);
and U5623 (N_5623,N_1556,N_636);
nand U5624 (N_5624,N_545,N_2475);
and U5625 (N_5625,N_1371,N_2065);
xor U5626 (N_5626,N_858,N_666);
xor U5627 (N_5627,N_1328,N_1232);
nand U5628 (N_5628,N_434,N_2547);
nor U5629 (N_5629,N_537,N_2693);
and U5630 (N_5630,N_2394,N_2912);
xor U5631 (N_5631,N_1433,N_1904);
xnor U5632 (N_5632,N_2481,N_176);
and U5633 (N_5633,N_1911,N_757);
nand U5634 (N_5634,N_2886,N_136);
nand U5635 (N_5635,N_2431,N_422);
and U5636 (N_5636,N_405,N_1774);
and U5637 (N_5637,N_1445,N_1059);
and U5638 (N_5638,N_685,N_1892);
nor U5639 (N_5639,N_2477,N_830);
nor U5640 (N_5640,N_2279,N_180);
nand U5641 (N_5641,N_968,N_2118);
nor U5642 (N_5642,N_2729,N_994);
nor U5643 (N_5643,N_1557,N_1194);
nor U5644 (N_5644,N_1400,N_159);
and U5645 (N_5645,N_1496,N_273);
xnor U5646 (N_5646,N_2470,N_1464);
nand U5647 (N_5647,N_145,N_1147);
and U5648 (N_5648,N_300,N_2786);
nand U5649 (N_5649,N_245,N_1749);
nand U5650 (N_5650,N_2622,N_1595);
nand U5651 (N_5651,N_45,N_827);
xor U5652 (N_5652,N_2275,N_2773);
nand U5653 (N_5653,N_2430,N_1225);
and U5654 (N_5654,N_786,N_2325);
and U5655 (N_5655,N_1358,N_683);
xor U5656 (N_5656,N_337,N_765);
and U5657 (N_5657,N_1336,N_1695);
or U5658 (N_5658,N_1828,N_105);
xor U5659 (N_5659,N_1209,N_2250);
or U5660 (N_5660,N_807,N_1379);
or U5661 (N_5661,N_2980,N_2648);
or U5662 (N_5662,N_2985,N_2489);
or U5663 (N_5663,N_947,N_1950);
xnor U5664 (N_5664,N_2026,N_2053);
or U5665 (N_5665,N_533,N_2877);
xor U5666 (N_5666,N_142,N_2006);
xor U5667 (N_5667,N_768,N_127);
xor U5668 (N_5668,N_2724,N_2139);
nand U5669 (N_5669,N_2107,N_1855);
or U5670 (N_5670,N_1183,N_977);
xor U5671 (N_5671,N_885,N_2222);
nor U5672 (N_5672,N_91,N_1912);
nor U5673 (N_5673,N_1916,N_1117);
nand U5674 (N_5674,N_414,N_1255);
nand U5675 (N_5675,N_2131,N_561);
nor U5676 (N_5676,N_2502,N_798);
or U5677 (N_5677,N_730,N_787);
or U5678 (N_5678,N_556,N_1815);
nand U5679 (N_5679,N_2573,N_2921);
nand U5680 (N_5680,N_728,N_905);
xnor U5681 (N_5681,N_2407,N_1980);
xor U5682 (N_5682,N_727,N_1614);
nand U5683 (N_5683,N_2503,N_695);
or U5684 (N_5684,N_297,N_1378);
xor U5685 (N_5685,N_2142,N_55);
and U5686 (N_5686,N_1433,N_2868);
nor U5687 (N_5687,N_990,N_1742);
or U5688 (N_5688,N_2563,N_2504);
xnor U5689 (N_5689,N_229,N_1310);
and U5690 (N_5690,N_1577,N_1980);
or U5691 (N_5691,N_2611,N_2980);
xnor U5692 (N_5692,N_2980,N_832);
xor U5693 (N_5693,N_2218,N_2241);
nor U5694 (N_5694,N_2836,N_67);
nand U5695 (N_5695,N_724,N_2568);
or U5696 (N_5696,N_1743,N_1914);
nor U5697 (N_5697,N_2759,N_1439);
xnor U5698 (N_5698,N_2875,N_2247);
and U5699 (N_5699,N_2689,N_1426);
nor U5700 (N_5700,N_250,N_128);
nand U5701 (N_5701,N_1552,N_476);
and U5702 (N_5702,N_2139,N_1093);
nand U5703 (N_5703,N_428,N_154);
or U5704 (N_5704,N_2688,N_1923);
nor U5705 (N_5705,N_1275,N_2161);
nand U5706 (N_5706,N_307,N_1089);
nor U5707 (N_5707,N_2821,N_209);
xnor U5708 (N_5708,N_2530,N_2093);
or U5709 (N_5709,N_2039,N_1536);
and U5710 (N_5710,N_610,N_1270);
and U5711 (N_5711,N_2642,N_2149);
nor U5712 (N_5712,N_728,N_2856);
nor U5713 (N_5713,N_1335,N_1706);
or U5714 (N_5714,N_152,N_217);
or U5715 (N_5715,N_1566,N_2190);
or U5716 (N_5716,N_1994,N_2489);
nand U5717 (N_5717,N_1246,N_2809);
xor U5718 (N_5718,N_2905,N_1558);
nor U5719 (N_5719,N_997,N_2428);
xor U5720 (N_5720,N_2485,N_745);
nor U5721 (N_5721,N_1047,N_514);
and U5722 (N_5722,N_2250,N_2457);
and U5723 (N_5723,N_2515,N_2834);
nor U5724 (N_5724,N_2003,N_1386);
nand U5725 (N_5725,N_1654,N_1082);
nand U5726 (N_5726,N_1862,N_2199);
and U5727 (N_5727,N_2051,N_1403);
nand U5728 (N_5728,N_2386,N_1926);
and U5729 (N_5729,N_1887,N_978);
nand U5730 (N_5730,N_2997,N_843);
or U5731 (N_5731,N_2761,N_2254);
nor U5732 (N_5732,N_1627,N_2376);
or U5733 (N_5733,N_2070,N_2144);
or U5734 (N_5734,N_43,N_647);
nand U5735 (N_5735,N_54,N_1334);
nand U5736 (N_5736,N_149,N_2705);
xnor U5737 (N_5737,N_1044,N_232);
nand U5738 (N_5738,N_2617,N_2726);
nand U5739 (N_5739,N_41,N_2026);
nand U5740 (N_5740,N_472,N_1412);
and U5741 (N_5741,N_931,N_2537);
nor U5742 (N_5742,N_947,N_1063);
nor U5743 (N_5743,N_2052,N_1783);
nand U5744 (N_5744,N_1171,N_2048);
xnor U5745 (N_5745,N_2986,N_919);
xnor U5746 (N_5746,N_1208,N_1870);
nand U5747 (N_5747,N_1927,N_2634);
nor U5748 (N_5748,N_258,N_1394);
or U5749 (N_5749,N_2839,N_990);
nor U5750 (N_5750,N_1504,N_1840);
and U5751 (N_5751,N_1044,N_189);
or U5752 (N_5752,N_400,N_1371);
nand U5753 (N_5753,N_2733,N_1413);
nor U5754 (N_5754,N_2469,N_2948);
xnor U5755 (N_5755,N_1013,N_454);
or U5756 (N_5756,N_2903,N_2138);
nand U5757 (N_5757,N_1823,N_611);
xor U5758 (N_5758,N_117,N_748);
and U5759 (N_5759,N_1964,N_1978);
nand U5760 (N_5760,N_1267,N_2769);
nor U5761 (N_5761,N_2783,N_199);
nand U5762 (N_5762,N_2535,N_2981);
nand U5763 (N_5763,N_1461,N_2453);
xnor U5764 (N_5764,N_2240,N_2739);
or U5765 (N_5765,N_872,N_1506);
nor U5766 (N_5766,N_1043,N_379);
or U5767 (N_5767,N_1446,N_1356);
or U5768 (N_5768,N_1363,N_968);
or U5769 (N_5769,N_880,N_594);
nor U5770 (N_5770,N_2434,N_1999);
xor U5771 (N_5771,N_173,N_1527);
xnor U5772 (N_5772,N_226,N_2613);
or U5773 (N_5773,N_2850,N_1322);
or U5774 (N_5774,N_700,N_1554);
or U5775 (N_5775,N_1999,N_641);
or U5776 (N_5776,N_1980,N_2463);
or U5777 (N_5777,N_831,N_2097);
xor U5778 (N_5778,N_735,N_1023);
and U5779 (N_5779,N_2902,N_811);
or U5780 (N_5780,N_2255,N_1840);
nand U5781 (N_5781,N_2905,N_2618);
nor U5782 (N_5782,N_2180,N_2801);
and U5783 (N_5783,N_456,N_945);
xor U5784 (N_5784,N_2486,N_2028);
nand U5785 (N_5785,N_2219,N_2637);
or U5786 (N_5786,N_1597,N_743);
or U5787 (N_5787,N_1928,N_2106);
nand U5788 (N_5788,N_522,N_2589);
or U5789 (N_5789,N_1913,N_1284);
xnor U5790 (N_5790,N_15,N_1623);
or U5791 (N_5791,N_2766,N_1863);
nor U5792 (N_5792,N_2655,N_2100);
nand U5793 (N_5793,N_1884,N_2167);
and U5794 (N_5794,N_2007,N_2080);
xnor U5795 (N_5795,N_2697,N_2278);
and U5796 (N_5796,N_263,N_269);
xor U5797 (N_5797,N_1851,N_350);
nor U5798 (N_5798,N_1670,N_2720);
xnor U5799 (N_5799,N_1159,N_297);
and U5800 (N_5800,N_1982,N_601);
xnor U5801 (N_5801,N_1945,N_1198);
nor U5802 (N_5802,N_669,N_2386);
xor U5803 (N_5803,N_2217,N_127);
nand U5804 (N_5804,N_1454,N_2254);
nand U5805 (N_5805,N_2570,N_1483);
nor U5806 (N_5806,N_988,N_2964);
and U5807 (N_5807,N_1309,N_2648);
xnor U5808 (N_5808,N_1168,N_2180);
nand U5809 (N_5809,N_101,N_709);
or U5810 (N_5810,N_1353,N_2335);
nand U5811 (N_5811,N_52,N_1054);
or U5812 (N_5812,N_2052,N_1265);
and U5813 (N_5813,N_1011,N_1444);
xor U5814 (N_5814,N_2644,N_1392);
and U5815 (N_5815,N_2106,N_722);
xor U5816 (N_5816,N_2240,N_2466);
and U5817 (N_5817,N_884,N_2569);
nand U5818 (N_5818,N_1743,N_1372);
or U5819 (N_5819,N_1718,N_2227);
xor U5820 (N_5820,N_64,N_1099);
nand U5821 (N_5821,N_2783,N_654);
xor U5822 (N_5822,N_592,N_602);
xnor U5823 (N_5823,N_215,N_2891);
xor U5824 (N_5824,N_2011,N_386);
xnor U5825 (N_5825,N_347,N_2811);
nor U5826 (N_5826,N_357,N_919);
xor U5827 (N_5827,N_2099,N_2170);
nor U5828 (N_5828,N_1851,N_2853);
or U5829 (N_5829,N_2215,N_1878);
xor U5830 (N_5830,N_1149,N_2492);
nand U5831 (N_5831,N_288,N_2784);
xor U5832 (N_5832,N_1135,N_2158);
nand U5833 (N_5833,N_2859,N_2388);
and U5834 (N_5834,N_192,N_203);
nand U5835 (N_5835,N_40,N_1429);
and U5836 (N_5836,N_28,N_364);
and U5837 (N_5837,N_87,N_2463);
xor U5838 (N_5838,N_1985,N_279);
and U5839 (N_5839,N_2843,N_2163);
nor U5840 (N_5840,N_1079,N_1315);
nand U5841 (N_5841,N_280,N_1195);
nand U5842 (N_5842,N_2733,N_918);
nor U5843 (N_5843,N_255,N_670);
nand U5844 (N_5844,N_903,N_575);
nand U5845 (N_5845,N_156,N_1373);
nor U5846 (N_5846,N_2890,N_1527);
and U5847 (N_5847,N_1367,N_1495);
or U5848 (N_5848,N_1402,N_2184);
and U5849 (N_5849,N_2132,N_294);
or U5850 (N_5850,N_2623,N_2790);
and U5851 (N_5851,N_2779,N_2800);
or U5852 (N_5852,N_2403,N_739);
or U5853 (N_5853,N_2932,N_942);
nor U5854 (N_5854,N_413,N_1383);
xnor U5855 (N_5855,N_1724,N_179);
xnor U5856 (N_5856,N_954,N_1665);
or U5857 (N_5857,N_502,N_1567);
nand U5858 (N_5858,N_2325,N_2228);
and U5859 (N_5859,N_71,N_2567);
xor U5860 (N_5860,N_1582,N_1491);
and U5861 (N_5861,N_129,N_859);
nor U5862 (N_5862,N_145,N_1862);
and U5863 (N_5863,N_1669,N_1201);
or U5864 (N_5864,N_414,N_1777);
nand U5865 (N_5865,N_2684,N_2449);
xor U5866 (N_5866,N_2158,N_513);
xnor U5867 (N_5867,N_1647,N_1810);
and U5868 (N_5868,N_2849,N_2295);
and U5869 (N_5869,N_104,N_1776);
nand U5870 (N_5870,N_1433,N_27);
nand U5871 (N_5871,N_734,N_2389);
xor U5872 (N_5872,N_1537,N_2184);
nor U5873 (N_5873,N_2391,N_1991);
nand U5874 (N_5874,N_1423,N_246);
nor U5875 (N_5875,N_2199,N_1974);
or U5876 (N_5876,N_1314,N_803);
or U5877 (N_5877,N_1397,N_2253);
and U5878 (N_5878,N_33,N_1743);
and U5879 (N_5879,N_1338,N_264);
xnor U5880 (N_5880,N_71,N_573);
or U5881 (N_5881,N_683,N_1816);
xor U5882 (N_5882,N_1583,N_2862);
nor U5883 (N_5883,N_17,N_1041);
or U5884 (N_5884,N_2107,N_2093);
xnor U5885 (N_5885,N_673,N_2470);
or U5886 (N_5886,N_2287,N_882);
or U5887 (N_5887,N_2180,N_130);
nand U5888 (N_5888,N_2512,N_1397);
or U5889 (N_5889,N_163,N_2064);
or U5890 (N_5890,N_234,N_1348);
nor U5891 (N_5891,N_2559,N_2520);
xor U5892 (N_5892,N_751,N_2691);
and U5893 (N_5893,N_1660,N_2680);
xnor U5894 (N_5894,N_1078,N_1296);
and U5895 (N_5895,N_1743,N_1463);
xnor U5896 (N_5896,N_1543,N_1403);
nand U5897 (N_5897,N_402,N_501);
nand U5898 (N_5898,N_727,N_2240);
and U5899 (N_5899,N_1879,N_1666);
and U5900 (N_5900,N_1352,N_2913);
or U5901 (N_5901,N_2819,N_1329);
xor U5902 (N_5902,N_2776,N_664);
nor U5903 (N_5903,N_393,N_238);
or U5904 (N_5904,N_1773,N_2375);
or U5905 (N_5905,N_2192,N_2136);
xnor U5906 (N_5906,N_1785,N_961);
and U5907 (N_5907,N_2248,N_910);
and U5908 (N_5908,N_2078,N_1179);
and U5909 (N_5909,N_716,N_1956);
nor U5910 (N_5910,N_1346,N_1329);
and U5911 (N_5911,N_910,N_2050);
nor U5912 (N_5912,N_2192,N_1510);
or U5913 (N_5913,N_2573,N_54);
or U5914 (N_5914,N_377,N_517);
and U5915 (N_5915,N_2599,N_1458);
and U5916 (N_5916,N_2776,N_985);
nand U5917 (N_5917,N_2738,N_2012);
or U5918 (N_5918,N_1686,N_2375);
nand U5919 (N_5919,N_651,N_448);
and U5920 (N_5920,N_967,N_2617);
and U5921 (N_5921,N_1541,N_2842);
or U5922 (N_5922,N_617,N_2348);
or U5923 (N_5923,N_314,N_2634);
and U5924 (N_5924,N_1789,N_460);
xor U5925 (N_5925,N_1873,N_830);
xor U5926 (N_5926,N_2039,N_522);
and U5927 (N_5927,N_2759,N_1956);
and U5928 (N_5928,N_887,N_1191);
xor U5929 (N_5929,N_2085,N_2057);
and U5930 (N_5930,N_138,N_2805);
and U5931 (N_5931,N_124,N_100);
and U5932 (N_5932,N_2457,N_1165);
nor U5933 (N_5933,N_205,N_1653);
or U5934 (N_5934,N_1581,N_1305);
xor U5935 (N_5935,N_1426,N_2630);
nand U5936 (N_5936,N_2459,N_2516);
nor U5937 (N_5937,N_2459,N_1898);
nor U5938 (N_5938,N_1013,N_1624);
nand U5939 (N_5939,N_2038,N_457);
xor U5940 (N_5940,N_1288,N_852);
and U5941 (N_5941,N_947,N_71);
xor U5942 (N_5942,N_214,N_2557);
nor U5943 (N_5943,N_883,N_2677);
xor U5944 (N_5944,N_1363,N_2761);
xnor U5945 (N_5945,N_683,N_1970);
nand U5946 (N_5946,N_307,N_333);
nor U5947 (N_5947,N_2835,N_460);
nand U5948 (N_5948,N_2027,N_2621);
xnor U5949 (N_5949,N_627,N_367);
nor U5950 (N_5950,N_1987,N_554);
and U5951 (N_5951,N_1913,N_2307);
xor U5952 (N_5952,N_728,N_1657);
and U5953 (N_5953,N_2024,N_158);
nor U5954 (N_5954,N_1055,N_1541);
xor U5955 (N_5955,N_2233,N_1632);
nand U5956 (N_5956,N_2466,N_2548);
and U5957 (N_5957,N_553,N_623);
xor U5958 (N_5958,N_591,N_1662);
or U5959 (N_5959,N_1521,N_1248);
and U5960 (N_5960,N_658,N_2680);
xnor U5961 (N_5961,N_2922,N_1649);
and U5962 (N_5962,N_1836,N_1333);
or U5963 (N_5963,N_1208,N_181);
and U5964 (N_5964,N_2078,N_2121);
or U5965 (N_5965,N_2711,N_571);
xnor U5966 (N_5966,N_2561,N_1291);
or U5967 (N_5967,N_1060,N_1947);
or U5968 (N_5968,N_2599,N_1870);
or U5969 (N_5969,N_368,N_1661);
nand U5970 (N_5970,N_2821,N_2384);
or U5971 (N_5971,N_227,N_2719);
nor U5972 (N_5972,N_2463,N_1830);
or U5973 (N_5973,N_2372,N_674);
nor U5974 (N_5974,N_1985,N_1835);
xor U5975 (N_5975,N_724,N_146);
xor U5976 (N_5976,N_2568,N_1122);
or U5977 (N_5977,N_1694,N_1086);
and U5978 (N_5978,N_2693,N_617);
and U5979 (N_5979,N_2170,N_1770);
xor U5980 (N_5980,N_997,N_474);
nand U5981 (N_5981,N_1978,N_231);
and U5982 (N_5982,N_2355,N_990);
or U5983 (N_5983,N_2435,N_785);
xor U5984 (N_5984,N_799,N_2739);
or U5985 (N_5985,N_2433,N_242);
nor U5986 (N_5986,N_2336,N_1270);
or U5987 (N_5987,N_45,N_189);
or U5988 (N_5988,N_2452,N_2314);
or U5989 (N_5989,N_1229,N_1567);
or U5990 (N_5990,N_718,N_1513);
xor U5991 (N_5991,N_2347,N_91);
nand U5992 (N_5992,N_117,N_806);
nand U5993 (N_5993,N_1498,N_2569);
nand U5994 (N_5994,N_811,N_1817);
and U5995 (N_5995,N_1909,N_1023);
xor U5996 (N_5996,N_1068,N_2404);
nand U5997 (N_5997,N_225,N_2463);
nor U5998 (N_5998,N_2347,N_1384);
nor U5999 (N_5999,N_156,N_30);
and U6000 (N_6000,N_3498,N_5353);
or U6001 (N_6001,N_3817,N_4773);
xor U6002 (N_6002,N_5108,N_4302);
nor U6003 (N_6003,N_5495,N_4751);
nor U6004 (N_6004,N_4019,N_4885);
nor U6005 (N_6005,N_3093,N_3082);
and U6006 (N_6006,N_4775,N_5464);
nor U6007 (N_6007,N_5135,N_5129);
nand U6008 (N_6008,N_5572,N_4383);
and U6009 (N_6009,N_5439,N_3346);
or U6010 (N_6010,N_3328,N_4635);
nand U6011 (N_6011,N_4009,N_4055);
xnor U6012 (N_6012,N_5753,N_4659);
xor U6013 (N_6013,N_5461,N_3601);
and U6014 (N_6014,N_3121,N_5574);
nand U6015 (N_6015,N_5845,N_4330);
and U6016 (N_6016,N_5412,N_4607);
nor U6017 (N_6017,N_3658,N_4040);
nand U6018 (N_6018,N_5898,N_5173);
nand U6019 (N_6019,N_4177,N_3831);
xor U6020 (N_6020,N_5023,N_4193);
nand U6021 (N_6021,N_3463,N_3253);
or U6022 (N_6022,N_3123,N_4792);
nor U6023 (N_6023,N_3245,N_4381);
or U6024 (N_6024,N_5921,N_3189);
nor U6025 (N_6025,N_3595,N_3260);
nand U6026 (N_6026,N_5150,N_5674);
nand U6027 (N_6027,N_3215,N_5823);
nand U6028 (N_6028,N_4220,N_4429);
nand U6029 (N_6029,N_4946,N_5838);
xor U6030 (N_6030,N_3235,N_5151);
or U6031 (N_6031,N_4991,N_3083);
nor U6032 (N_6032,N_3292,N_3434);
or U6033 (N_6033,N_4272,N_5097);
or U6034 (N_6034,N_4187,N_3876);
and U6035 (N_6035,N_4434,N_3839);
nor U6036 (N_6036,N_5250,N_4701);
and U6037 (N_6037,N_5923,N_5655);
and U6038 (N_6038,N_5643,N_4927);
nand U6039 (N_6039,N_4172,N_5628);
and U6040 (N_6040,N_4492,N_3792);
nand U6041 (N_6041,N_5208,N_4911);
nand U6042 (N_6042,N_5294,N_3154);
nand U6043 (N_6043,N_4063,N_5486);
nand U6044 (N_6044,N_5121,N_3425);
nand U6045 (N_6045,N_5858,N_3566);
and U6046 (N_6046,N_4795,N_5611);
xor U6047 (N_6047,N_3937,N_5962);
nor U6048 (N_6048,N_5679,N_4206);
xnor U6049 (N_6049,N_4839,N_4665);
nand U6050 (N_6050,N_3787,N_3870);
and U6051 (N_6051,N_3207,N_4028);
nor U6052 (N_6052,N_4630,N_4122);
xor U6053 (N_6053,N_4493,N_4866);
and U6054 (N_6054,N_5888,N_4616);
nor U6055 (N_6055,N_4244,N_5710);
nand U6056 (N_6056,N_4502,N_5180);
nand U6057 (N_6057,N_4550,N_3389);
xor U6058 (N_6058,N_5577,N_5992);
nand U6059 (N_6059,N_4241,N_5455);
or U6060 (N_6060,N_4279,N_4427);
nor U6061 (N_6061,N_3842,N_5816);
nand U6062 (N_6062,N_4274,N_5204);
or U6063 (N_6063,N_4849,N_3579);
or U6064 (N_6064,N_4370,N_3310);
nand U6065 (N_6065,N_4826,N_4237);
nand U6066 (N_6066,N_4819,N_4555);
nor U6067 (N_6067,N_3362,N_5546);
or U6068 (N_6068,N_3181,N_4915);
and U6069 (N_6069,N_3802,N_4075);
and U6070 (N_6070,N_3730,N_4534);
xnor U6071 (N_6071,N_5685,N_3963);
or U6072 (N_6072,N_3759,N_5201);
nor U6073 (N_6073,N_3195,N_5314);
xnor U6074 (N_6074,N_5553,N_3869);
nor U6075 (N_6075,N_5423,N_5926);
or U6076 (N_6076,N_4796,N_5080);
or U6077 (N_6077,N_4338,N_4877);
nand U6078 (N_6078,N_3496,N_3473);
nand U6079 (N_6079,N_4703,N_5531);
nand U6080 (N_6080,N_4571,N_4506);
and U6081 (N_6081,N_3893,N_4173);
xnor U6082 (N_6082,N_5182,N_5079);
and U6083 (N_6083,N_3594,N_5790);
and U6084 (N_6084,N_4987,N_4368);
nor U6085 (N_6085,N_3702,N_4322);
nor U6086 (N_6086,N_3138,N_5072);
nor U6087 (N_6087,N_5098,N_5882);
nand U6088 (N_6088,N_4830,N_5758);
and U6089 (N_6089,N_5467,N_5369);
and U6090 (N_6090,N_4566,N_3399);
nand U6091 (N_6091,N_4233,N_3677);
nor U6092 (N_6092,N_3353,N_4198);
xnor U6093 (N_6093,N_3222,N_3948);
nand U6094 (N_6094,N_5683,N_3731);
or U6095 (N_6095,N_4085,N_3533);
xor U6096 (N_6096,N_4988,N_4413);
xor U6097 (N_6097,N_3144,N_4867);
xor U6098 (N_6098,N_4903,N_5402);
or U6099 (N_6099,N_3768,N_3526);
and U6100 (N_6100,N_4336,N_3805);
or U6101 (N_6101,N_3846,N_3779);
and U6102 (N_6102,N_5945,N_5364);
nand U6103 (N_6103,N_3020,N_4704);
xnor U6104 (N_6104,N_4247,N_3429);
nor U6105 (N_6105,N_5367,N_3199);
xor U6106 (N_6106,N_3014,N_5307);
nand U6107 (N_6107,N_4437,N_3307);
nor U6108 (N_6108,N_5869,N_5030);
nor U6109 (N_6109,N_4045,N_5360);
nand U6110 (N_6110,N_4201,N_5184);
and U6111 (N_6111,N_3012,N_5510);
or U6112 (N_6112,N_4315,N_3524);
or U6113 (N_6113,N_5998,N_3085);
nor U6114 (N_6114,N_5465,N_5549);
nand U6115 (N_6115,N_3243,N_5269);
nor U6116 (N_6116,N_4746,N_4214);
or U6117 (N_6117,N_5871,N_3913);
nor U6118 (N_6118,N_3974,N_5948);
and U6119 (N_6119,N_3666,N_4949);
nor U6120 (N_6120,N_4408,N_3290);
nand U6121 (N_6121,N_3288,N_3391);
xnor U6122 (N_6122,N_3372,N_4916);
xnor U6123 (N_6123,N_5397,N_3572);
or U6124 (N_6124,N_4347,N_3849);
and U6125 (N_6125,N_5185,N_3190);
nor U6126 (N_6126,N_3981,N_4405);
or U6127 (N_6127,N_5094,N_3440);
and U6128 (N_6128,N_5985,N_4634);
and U6129 (N_6129,N_5291,N_4419);
or U6130 (N_6130,N_5015,N_4791);
nand U6131 (N_6131,N_5614,N_3487);
xnor U6132 (N_6132,N_3737,N_5386);
nor U6133 (N_6133,N_5444,N_3007);
or U6134 (N_6134,N_4475,N_5462);
and U6135 (N_6135,N_3646,N_4742);
nand U6136 (N_6136,N_4562,N_4275);
nor U6137 (N_6137,N_4878,N_4872);
xnor U6138 (N_6138,N_5558,N_4726);
or U6139 (N_6139,N_5138,N_3477);
nor U6140 (N_6140,N_5435,N_5761);
nor U6141 (N_6141,N_5528,N_3590);
xnor U6142 (N_6142,N_5914,N_3764);
nor U6143 (N_6143,N_3158,N_4887);
or U6144 (N_6144,N_3452,N_3823);
or U6145 (N_6145,N_5246,N_3006);
xnor U6146 (N_6146,N_4091,N_4990);
and U6147 (N_6147,N_4443,N_5885);
or U6148 (N_6148,N_5841,N_3616);
nand U6149 (N_6149,N_5339,N_5925);
and U6150 (N_6150,N_3311,N_4612);
or U6151 (N_6151,N_4137,N_3907);
or U6152 (N_6152,N_3920,N_3635);
nor U6153 (N_6153,N_4814,N_5934);
nor U6154 (N_6154,N_3044,N_5603);
and U6155 (N_6155,N_3280,N_4258);
xnor U6156 (N_6156,N_3567,N_4513);
and U6157 (N_6157,N_3274,N_3035);
nand U6158 (N_6158,N_3095,N_4891);
nand U6159 (N_6159,N_5209,N_4544);
xor U6160 (N_6160,N_3914,N_3697);
nand U6161 (N_6161,N_3358,N_4287);
nand U6162 (N_6162,N_5227,N_4467);
and U6163 (N_6163,N_3514,N_5740);
xor U6164 (N_6164,N_3556,N_4216);
nor U6165 (N_6165,N_3554,N_5379);
or U6166 (N_6166,N_5484,N_4813);
or U6167 (N_6167,N_4770,N_4442);
nor U6168 (N_6168,N_3850,N_3064);
and U6169 (N_6169,N_4962,N_5324);
and U6170 (N_6170,N_4453,N_5265);
nand U6171 (N_6171,N_5835,N_4471);
nand U6172 (N_6172,N_3972,N_5140);
or U6173 (N_6173,N_4108,N_5832);
or U6174 (N_6174,N_4376,N_5037);
nor U6175 (N_6175,N_3860,N_3909);
xnor U6176 (N_6176,N_5622,N_3987);
nand U6177 (N_6177,N_4595,N_3111);
nor U6178 (N_6178,N_4545,N_3874);
nand U6179 (N_6179,N_4426,N_5441);
or U6180 (N_6180,N_3977,N_5604);
nand U6181 (N_6181,N_4890,N_5113);
and U6182 (N_6182,N_4558,N_3157);
nand U6183 (N_6183,N_5124,N_5283);
nor U6184 (N_6184,N_5247,N_4357);
or U6185 (N_6185,N_4951,N_3406);
and U6186 (N_6186,N_5843,N_3669);
nand U6187 (N_6187,N_3332,N_4486);
nand U6188 (N_6188,N_3612,N_3667);
xnor U6189 (N_6189,N_4715,N_5300);
and U6190 (N_6190,N_4646,N_4133);
and U6191 (N_6191,N_3531,N_3967);
nor U6192 (N_6192,N_5449,N_5863);
and U6193 (N_6193,N_5220,N_3808);
and U6194 (N_6194,N_5489,N_4098);
or U6195 (N_6195,N_3439,N_3177);
or U6196 (N_6196,N_3132,N_3467);
xnor U6197 (N_6197,N_5183,N_4393);
and U6198 (N_6198,N_4359,N_4823);
xor U6199 (N_6199,N_5343,N_3286);
nor U6200 (N_6200,N_5957,N_4662);
xnor U6201 (N_6201,N_4447,N_3994);
xnor U6202 (N_6202,N_4304,N_3855);
and U6203 (N_6203,N_4253,N_3578);
nor U6204 (N_6204,N_5236,N_5366);
xor U6205 (N_6205,N_4208,N_3427);
nor U6206 (N_6206,N_4631,N_5984);
and U6207 (N_6207,N_5949,N_3386);
xnor U6208 (N_6208,N_3305,N_3945);
or U6209 (N_6209,N_5411,N_4879);
xor U6210 (N_6210,N_5468,N_3062);
and U6211 (N_6211,N_5652,N_5243);
and U6212 (N_6212,N_4568,N_5445);
xnor U6213 (N_6213,N_4228,N_5479);
xnor U6214 (N_6214,N_3300,N_4810);
nand U6215 (N_6215,N_3534,N_3668);
xor U6216 (N_6216,N_3219,N_3865);
or U6217 (N_6217,N_4356,N_5705);
nor U6218 (N_6218,N_5615,N_3150);
or U6219 (N_6219,N_4348,N_4976);
nand U6220 (N_6220,N_3344,N_3706);
and U6221 (N_6221,N_5211,N_3843);
or U6222 (N_6222,N_3308,N_3167);
nand U6223 (N_6223,N_3185,N_4025);
xnor U6224 (N_6224,N_5341,N_3387);
xnor U6225 (N_6225,N_3584,N_5975);
xor U6226 (N_6226,N_3693,N_4308);
nand U6227 (N_6227,N_5930,N_3117);
or U6228 (N_6228,N_4585,N_3170);
nor U6229 (N_6229,N_3866,N_5064);
nand U6230 (N_6230,N_3072,N_5126);
nand U6231 (N_6231,N_5706,N_5177);
and U6232 (N_6232,N_5387,N_3350);
nor U6233 (N_6233,N_4755,N_4231);
and U6234 (N_6234,N_4152,N_3797);
xor U6235 (N_6235,N_4886,N_4549);
nor U6236 (N_6236,N_4730,N_3890);
nand U6237 (N_6237,N_5487,N_3211);
or U6238 (N_6238,N_5480,N_3262);
nor U6239 (N_6239,N_3597,N_4160);
xor U6240 (N_6240,N_4226,N_3365);
or U6241 (N_6241,N_4473,N_4217);
nor U6242 (N_6242,N_3027,N_3106);
or U6243 (N_6243,N_5092,N_5349);
or U6244 (N_6244,N_3061,N_5867);
nor U6245 (N_6245,N_5280,N_4709);
and U6246 (N_6246,N_3281,N_3403);
and U6247 (N_6247,N_3562,N_5765);
or U6248 (N_6248,N_5844,N_3785);
xor U6249 (N_6249,N_3560,N_3873);
nand U6250 (N_6250,N_3796,N_5716);
nand U6251 (N_6251,N_5070,N_3337);
and U6252 (N_6252,N_5334,N_3136);
xnor U6253 (N_6253,N_3416,N_4954);
and U6254 (N_6254,N_5980,N_4981);
or U6255 (N_6255,N_5096,N_4968);
xor U6256 (N_6256,N_4093,N_3315);
nor U6257 (N_6257,N_5556,N_5703);
xnor U6258 (N_6258,N_4622,N_3047);
nand U6259 (N_6259,N_3564,N_4252);
or U6260 (N_6260,N_4711,N_3225);
and U6261 (N_6261,N_5218,N_4215);
xnor U6262 (N_6262,N_4477,N_5046);
and U6263 (N_6263,N_4515,N_4171);
or U6264 (N_6264,N_3793,N_3236);
or U6265 (N_6265,N_3322,N_5996);
and U6266 (N_6266,N_5315,N_5538);
xnor U6267 (N_6267,N_4606,N_3513);
nand U6268 (N_6268,N_5640,N_4260);
nor U6269 (N_6269,N_5336,N_5325);
nand U6270 (N_6270,N_4780,N_5348);
or U6271 (N_6271,N_5627,N_4331);
and U6272 (N_6272,N_4644,N_5646);
or U6273 (N_6273,N_5606,N_3885);
and U6274 (N_6274,N_5210,N_3806);
nor U6275 (N_6275,N_4116,N_4836);
nand U6276 (N_6276,N_3636,N_5191);
or U6277 (N_6277,N_4068,N_4015);
and U6278 (N_6278,N_3917,N_4176);
or U6279 (N_6279,N_4615,N_3816);
nand U6280 (N_6280,N_5401,N_3600);
xnor U6281 (N_6281,N_4871,N_4066);
nor U6282 (N_6282,N_3950,N_3747);
and U6283 (N_6283,N_5459,N_5517);
xnor U6284 (N_6284,N_4251,N_3475);
nor U6285 (N_6285,N_5273,N_5986);
nor U6286 (N_6286,N_3134,N_5632);
or U6287 (N_6287,N_3375,N_4863);
nor U6288 (N_6288,N_4065,N_4959);
nand U6289 (N_6289,N_5954,N_4933);
nor U6290 (N_6290,N_3443,N_3774);
and U6291 (N_6291,N_4067,N_4552);
nor U6292 (N_6292,N_3946,N_3544);
or U6293 (N_6293,N_5289,N_5678);
and U6294 (N_6294,N_3980,N_3645);
or U6295 (N_6295,N_4974,N_4759);
nor U6296 (N_6296,N_4969,N_3650);
or U6297 (N_6297,N_5785,N_5454);
or U6298 (N_6298,N_4194,N_5680);
and U6299 (N_6299,N_4827,N_5205);
or U6300 (N_6300,N_5071,N_5909);
or U6301 (N_6301,N_5125,N_4922);
or U6302 (N_6302,N_4488,N_3471);
or U6303 (N_6303,N_3238,N_4110);
xor U6304 (N_6304,N_3216,N_5817);
and U6305 (N_6305,N_4318,N_4594);
or U6306 (N_6306,N_4689,N_5372);
xor U6307 (N_6307,N_4124,N_3383);
and U6308 (N_6308,N_5702,N_4563);
xnor U6309 (N_6309,N_4501,N_3279);
or U6310 (N_6310,N_4569,N_4543);
or U6311 (N_6311,N_4710,N_5061);
nand U6312 (N_6312,N_5798,N_5158);
xnor U6313 (N_6313,N_3491,N_4485);
or U6314 (N_6314,N_5175,N_3825);
nor U6315 (N_6315,N_5049,N_4313);
nand U6316 (N_6316,N_3736,N_4151);
nor U6317 (N_6317,N_4103,N_5241);
xor U6318 (N_6318,N_5800,N_3413);
nor U6319 (N_6319,N_4465,N_4738);
xor U6320 (N_6320,N_3749,N_5176);
or U6321 (N_6321,N_5483,N_5115);
or U6322 (N_6322,N_5248,N_3244);
xor U6323 (N_6323,N_5769,N_4284);
nand U6324 (N_6324,N_5866,N_3700);
nand U6325 (N_6325,N_5697,N_4510);
nor U6326 (N_6326,N_3721,N_5195);
nor U6327 (N_6327,N_4170,N_4597);
nor U6328 (N_6328,N_3910,N_4530);
and U6329 (N_6329,N_3448,N_4668);
or U6330 (N_6330,N_3819,N_5249);
nor U6331 (N_6331,N_5935,N_5744);
and U6332 (N_6332,N_4736,N_3008);
nor U6333 (N_6333,N_4495,N_5997);
or U6334 (N_6334,N_5982,N_4483);
and U6335 (N_6335,N_5525,N_4538);
xor U6336 (N_6336,N_5752,N_5216);
or U6337 (N_6337,N_4683,N_5356);
nand U6338 (N_6338,N_5073,N_5965);
nor U6339 (N_6339,N_3940,N_3241);
or U6340 (N_6340,N_5764,N_3193);
nand U6341 (N_6341,N_3367,N_3795);
or U6342 (N_6342,N_5024,N_4306);
nand U6343 (N_6343,N_4999,N_5551);
xor U6344 (N_6344,N_3751,N_3101);
or U6345 (N_6345,N_5735,N_3735);
xor U6346 (N_6346,N_5013,N_3548);
nand U6347 (N_6347,N_3436,N_3428);
and U6348 (N_6348,N_5991,N_3951);
nor U6349 (N_6349,N_4006,N_5629);
nor U6350 (N_6350,N_4749,N_5178);
or U6351 (N_6351,N_5742,N_5554);
and U6352 (N_6352,N_5378,N_3761);
xnor U6353 (N_6353,N_5365,N_3649);
or U6354 (N_6354,N_4511,N_3485);
nand U6355 (N_6355,N_3714,N_3033);
or U6356 (N_6356,N_3188,N_5700);
or U6357 (N_6357,N_4280,N_3501);
or U6358 (N_6358,N_5292,N_4784);
nand U6359 (N_6359,N_5750,N_5899);
xor U6360 (N_6360,N_5575,N_3208);
xnor U6361 (N_6361,N_5598,N_3527);
nor U6362 (N_6362,N_4650,N_4654);
or U6363 (N_6363,N_3370,N_3187);
or U6364 (N_6364,N_3617,N_4599);
and U6365 (N_6365,N_5006,N_5815);
and U6366 (N_6366,N_4895,N_3986);
xor U6367 (N_6367,N_4817,N_5557);
nor U6368 (N_6368,N_5457,N_5805);
or U6369 (N_6369,N_4059,N_4084);
and U6370 (N_6370,N_4632,N_3517);
xor U6371 (N_6371,N_3511,N_4591);
and U6372 (N_6372,N_4460,N_4892);
and U6373 (N_6373,N_5145,N_5748);
nand U6374 (N_6374,N_4812,N_3343);
nor U6375 (N_6375,N_5880,N_5895);
nor U6376 (N_6376,N_4192,N_3979);
and U6377 (N_6377,N_5448,N_3329);
nor U6378 (N_6378,N_5268,N_3165);
nor U6379 (N_6379,N_5022,N_5533);
xnor U6380 (N_6380,N_5492,N_3031);
nand U6381 (N_6381,N_3934,N_3282);
or U6382 (N_6382,N_3586,N_4672);
nor U6383 (N_6383,N_5038,N_5395);
nand U6384 (N_6384,N_4620,N_3456);
nand U6385 (N_6385,N_3164,N_3541);
and U6386 (N_6386,N_3388,N_4870);
and U6387 (N_6387,N_3419,N_5482);
nand U6388 (N_6388,N_4123,N_3753);
nand U6389 (N_6389,N_3921,N_4404);
and U6390 (N_6390,N_4052,N_4760);
nand U6391 (N_6391,N_3720,N_5257);
xor U6392 (N_6392,N_5394,N_5668);
and U6393 (N_6393,N_5035,N_3906);
nand U6394 (N_6394,N_4708,N_3915);
or U6395 (N_6395,N_4986,N_3698);
nor U6396 (N_6396,N_3990,N_5213);
nor U6397 (N_6397,N_5593,N_4120);
or U6398 (N_6398,N_4663,N_4264);
nor U6399 (N_6399,N_5421,N_4167);
xnor U6400 (N_6400,N_3109,N_4929);
nor U6401 (N_6401,N_5864,N_5760);
xnor U6402 (N_6402,N_5424,N_5712);
and U6403 (N_6403,N_3856,N_5718);
and U6404 (N_6404,N_4833,N_5601);
and U6405 (N_6405,N_5146,N_3743);
nand U6406 (N_6406,N_3576,N_4029);
and U6407 (N_6407,N_4271,N_3287);
nor U6408 (N_6408,N_5561,N_5034);
xor U6409 (N_6409,N_5896,N_4535);
or U6410 (N_6410,N_3159,N_5266);
nor U6411 (N_6411,N_5131,N_3359);
nor U6412 (N_6412,N_5513,N_3005);
or U6413 (N_6413,N_3277,N_3203);
xor U6414 (N_6414,N_5407,N_3581);
and U6415 (N_6415,N_5578,N_4637);
nand U6416 (N_6416,N_3681,N_4536);
nand U6417 (N_6417,N_3297,N_4906);
and U6418 (N_6418,N_5739,N_3662);
or U6419 (N_6419,N_3458,N_3480);
nand U6420 (N_6420,N_3090,N_5103);
nor U6421 (N_6421,N_5335,N_4086);
nand U6422 (N_6422,N_3151,N_4223);
or U6423 (N_6423,N_3385,N_4853);
or U6424 (N_6424,N_4765,N_3896);
nor U6425 (N_6425,N_5074,N_5879);
nor U6426 (N_6426,N_5820,N_5347);
xnor U6427 (N_6427,N_5897,N_5605);
and U6428 (N_6428,N_5799,N_3392);
nand U6429 (N_6429,N_3537,N_5520);
nor U6430 (N_6430,N_4458,N_5919);
nor U6431 (N_6431,N_4802,N_4769);
nand U6432 (N_6432,N_5989,N_3004);
and U6433 (N_6433,N_3405,N_5729);
xnor U6434 (N_6434,N_4261,N_5978);
and U6435 (N_6435,N_3659,N_3997);
or U6436 (N_6436,N_5027,N_4582);
nor U6437 (N_6437,N_4380,N_5442);
nor U6438 (N_6438,N_5631,N_4387);
nor U6439 (N_6439,N_3989,N_4189);
or U6440 (N_6440,N_3587,N_3559);
xnor U6441 (N_6441,N_5833,N_3794);
nand U6442 (N_6442,N_4633,N_4466);
nand U6443 (N_6443,N_4428,N_3178);
nand U6444 (N_6444,N_5384,N_4130);
or U6445 (N_6445,N_4047,N_5304);
or U6446 (N_6446,N_5050,N_4245);
xnor U6447 (N_6447,N_4449,N_3663);
nor U6448 (N_6448,N_5009,N_5226);
and U6449 (N_6449,N_4482,N_5008);
nor U6450 (N_6450,N_5566,N_4923);
xnor U6451 (N_6451,N_3060,N_5245);
or U6452 (N_6452,N_3333,N_5704);
xor U6453 (N_6453,N_5390,N_4378);
nor U6454 (N_6454,N_4077,N_5824);
nor U6455 (N_6455,N_3326,N_4529);
and U6456 (N_6456,N_4840,N_3054);
nor U6457 (N_6457,N_4864,N_3438);
and U6458 (N_6458,N_5597,N_5618);
or U6459 (N_6459,N_5276,N_3933);
nand U6460 (N_6460,N_3727,N_4512);
xor U6461 (N_6461,N_5787,N_4145);
or U6462 (N_6462,N_5282,N_5796);
nand U6463 (N_6463,N_4003,N_5701);
nor U6464 (N_6464,N_3366,N_4756);
nand U6465 (N_6465,N_5795,N_5481);
xnor U6466 (N_6466,N_3461,N_4416);
or U6467 (N_6467,N_4459,N_3993);
xor U6468 (N_6468,N_4776,N_3045);
xor U6469 (N_6469,N_4869,N_3878);
nor U6470 (N_6470,N_3931,N_5144);
nand U6471 (N_6471,N_3112,N_3829);
nor U6472 (N_6472,N_4020,N_3113);
xnor U6473 (N_6473,N_3968,N_4551);
and U6474 (N_6474,N_5305,N_3409);
and U6475 (N_6475,N_3071,N_5583);
nand U6476 (N_6476,N_4143,N_5694);
xnor U6477 (N_6477,N_5950,N_5499);
or U6478 (N_6478,N_3686,N_4798);
and U6479 (N_6479,N_3445,N_3820);
xor U6480 (N_6480,N_5279,N_5648);
and U6481 (N_6481,N_3770,N_4178);
or U6482 (N_6482,N_5840,N_5532);
nor U6483 (N_6483,N_3074,N_4102);
nor U6484 (N_6484,N_3791,N_3381);
nand U6485 (N_6485,N_3745,N_3046);
and U6486 (N_6486,N_5418,N_4960);
nor U6487 (N_6487,N_5848,N_5901);
and U6488 (N_6488,N_5822,N_5792);
xor U6489 (N_6489,N_3361,N_5054);
nand U6490 (N_6490,N_4575,N_3153);
or U6491 (N_6491,N_4463,N_5156);
xnor U6492 (N_6492,N_3466,N_4517);
xnor U6493 (N_6493,N_5040,N_5726);
and U6494 (N_6494,N_5147,N_3271);
or U6495 (N_6495,N_5200,N_4600);
and U6496 (N_6496,N_5354,N_3563);
nand U6497 (N_6497,N_3276,N_3675);
xnor U6498 (N_6498,N_5987,N_4588);
xnor U6499 (N_6499,N_3536,N_5281);
and U6500 (N_6500,N_4246,N_5639);
nor U6501 (N_6501,N_4508,N_3710);
nor U6502 (N_6502,N_3168,N_5596);
nand U6503 (N_6503,N_5310,N_3613);
nor U6504 (N_6504,N_4844,N_5964);
and U6505 (N_6505,N_4311,N_5497);
and U6506 (N_6506,N_3695,N_5446);
nor U6507 (N_6507,N_3508,N_3573);
and U6508 (N_6508,N_5406,N_3380);
and U6509 (N_6509,N_3139,N_5306);
nor U6510 (N_6510,N_4398,N_5052);
or U6511 (N_6511,N_5186,N_4363);
nor U6512 (N_6512,N_4083,N_3146);
nor U6513 (N_6513,N_5337,N_3327);
xor U6514 (N_6514,N_5385,N_5666);
xnor U6515 (N_6515,N_4101,N_3063);
nor U6516 (N_6516,N_4257,N_3097);
nor U6517 (N_6517,N_5344,N_4125);
or U6518 (N_6518,N_4461,N_3431);
and U6519 (N_6519,N_3591,N_5906);
or U6520 (N_6520,N_4992,N_4388);
nor U6521 (N_6521,N_3551,N_3781);
nor U6522 (N_6522,N_3331,N_5883);
or U6523 (N_6523,N_5116,N_4937);
nor U6524 (N_6524,N_3773,N_3970);
xor U6525 (N_6525,N_5782,N_3098);
nand U6526 (N_6526,N_4438,N_3631);
xnor U6527 (N_6527,N_5212,N_4390);
nand U6528 (N_6528,N_4012,N_3529);
or U6529 (N_6529,N_3130,N_3261);
nand U6530 (N_6530,N_4050,N_4850);
and U6531 (N_6531,N_4344,N_4762);
and U6532 (N_6532,N_3499,N_3201);
or U6533 (N_6533,N_4785,N_5959);
and U6534 (N_6534,N_4115,N_4418);
and U6535 (N_6535,N_3246,N_3778);
xnor U6536 (N_6536,N_3127,N_3826);
xor U6537 (N_6537,N_3644,N_4195);
nand U6538 (N_6538,N_4129,N_3102);
xor U6539 (N_6539,N_5527,N_3003);
xnor U6540 (N_6540,N_4681,N_3204);
nor U6541 (N_6541,N_5788,N_5229);
nor U6542 (N_6542,N_4153,N_4693);
xnor U6543 (N_6543,N_3894,N_5550);
nor U6544 (N_6544,N_4462,N_4931);
and U6545 (N_6545,N_3887,N_3859);
nor U6546 (N_6546,N_5505,N_3393);
nand U6547 (N_6547,N_5960,N_5154);
nand U6548 (N_6548,N_3682,N_5828);
xnor U6549 (N_6549,N_4856,N_5107);
or U6550 (N_6550,N_3903,N_5889);
and U6551 (N_6551,N_5187,N_5399);
xnor U6552 (N_6552,N_5720,N_3918);
xor U6553 (N_6553,N_4300,N_4932);
and U6554 (N_6554,N_4384,N_3577);
and U6555 (N_6555,N_3451,N_4188);
or U6556 (N_6556,N_4598,N_4793);
xor U6557 (N_6557,N_5398,N_4329);
or U6558 (N_6558,N_5181,N_5298);
nor U6559 (N_6559,N_4786,N_4979);
and U6560 (N_6560,N_3379,N_3492);
nand U6561 (N_6561,N_3956,N_4452);
nor U6562 (N_6562,N_3857,N_5207);
xnor U6563 (N_6563,N_5228,N_4435);
and U6564 (N_6564,N_4702,N_4499);
xor U6565 (N_6565,N_5326,N_3639);
nand U6566 (N_6566,N_4079,N_5428);
and U6567 (N_6567,N_5734,N_4494);
nor U6568 (N_6568,N_3834,N_3943);
and U6569 (N_6569,N_3881,N_5222);
xor U6570 (N_6570,N_3032,N_5669);
xnor U6571 (N_6571,N_3641,N_5288);
and U6572 (N_6572,N_3512,N_5927);
nand U6573 (N_6573,N_5284,N_5903);
xor U6574 (N_6574,N_3205,N_5902);
and U6575 (N_6575,N_3395,N_4661);
nand U6576 (N_6576,N_3756,N_5252);
nor U6577 (N_6577,N_5916,N_4695);
or U6578 (N_6578,N_4829,N_5617);
and U6579 (N_6579,N_3852,N_4046);
xnor U6580 (N_6580,N_3627,N_5861);
or U6581 (N_6581,N_5893,N_4104);
and U6582 (N_6582,N_3437,N_4262);
xnor U6583 (N_6583,N_4044,N_5552);
nand U6584 (N_6584,N_3418,N_5779);
and U6585 (N_6585,N_3075,N_3051);
xnor U6586 (N_6586,N_5507,N_3019);
nor U6587 (N_6587,N_3861,N_4162);
xor U6588 (N_6588,N_3927,N_3103);
or U6589 (N_6589,N_3643,N_3209);
nor U6590 (N_6590,N_3854,N_3984);
or U6591 (N_6591,N_5842,N_5931);
nand U6592 (N_6592,N_4540,N_4034);
and U6593 (N_6593,N_4431,N_4945);
nand U6594 (N_6594,N_3814,N_5350);
nand U6595 (N_6595,N_4056,N_4614);
and U6596 (N_6596,N_4150,N_4647);
and U6597 (N_6597,N_5653,N_5104);
xnor U6598 (N_6598,N_5171,N_4561);
nand U6599 (N_6599,N_3010,N_5028);
and U6600 (N_6600,N_3574,N_4651);
nor U6601 (N_6601,N_5362,N_4277);
nor U6602 (N_6602,N_5469,N_5067);
xor U6603 (N_6603,N_5301,N_4327);
or U6604 (N_6604,N_4340,N_3615);
and U6605 (N_6605,N_3786,N_3804);
or U6606 (N_6606,N_3363,N_5657);
nand U6607 (N_6607,N_5846,N_4698);
nor U6608 (N_6608,N_4725,N_3030);
and U6609 (N_6609,N_5238,N_4432);
nand U6610 (N_6610,N_4234,N_4021);
xnor U6611 (N_6611,N_4367,N_3056);
nor U6612 (N_6612,N_3884,N_4298);
or U6613 (N_6613,N_4617,N_4670);
or U6614 (N_6614,N_3654,N_3299);
nand U6615 (N_6615,N_4847,N_4740);
nor U6616 (N_6616,N_4787,N_3259);
xor U6617 (N_6617,N_3478,N_3504);
and U6618 (N_6618,N_5755,N_4669);
xor U6619 (N_6619,N_3435,N_3449);
nor U6620 (N_6620,N_4956,N_5254);
or U6621 (N_6621,N_5834,N_5419);
or U6622 (N_6622,N_5771,N_3404);
nor U6623 (N_6623,N_3925,N_3765);
or U6624 (N_6624,N_4420,N_4901);
and U6625 (N_6625,N_3119,N_5784);
and U6626 (N_6626,N_4325,N_4169);
and U6627 (N_6627,N_4403,N_3828);
xor U6628 (N_6628,N_4675,N_4126);
or U6629 (N_6629,N_5660,N_4982);
and U6630 (N_6630,N_4642,N_3716);
or U6631 (N_6631,N_4842,N_4880);
nand U6632 (N_6632,N_4621,N_4970);
or U6633 (N_6633,N_4165,N_5966);
nor U6634 (N_6634,N_3585,N_3518);
nand U6635 (N_6635,N_3285,N_5837);
xor U6636 (N_6636,N_5952,N_3926);
nand U6637 (N_6637,N_4801,N_5117);
and U6638 (N_6638,N_5774,N_5477);
or U6639 (N_6639,N_3505,N_4586);
and U6640 (N_6640,N_5958,N_5509);
and U6641 (N_6641,N_4924,N_4832);
or U6642 (N_6642,N_5019,N_5410);
xnor U6643 (N_6643,N_3506,N_3995);
or U6644 (N_6644,N_5918,N_4790);
nand U6645 (N_6645,N_3000,N_5524);
nand U6646 (N_6646,N_5667,N_4478);
and U6647 (N_6647,N_5630,N_3464);
xor U6648 (N_6648,N_3470,N_3687);
and U6649 (N_6649,N_5634,N_5745);
nand U6650 (N_6650,N_5235,N_5961);
and U6651 (N_6651,N_4335,N_4392);
nand U6652 (N_6652,N_4476,N_5166);
nor U6653 (N_6653,N_4777,N_4334);
nand U6654 (N_6654,N_5346,N_5699);
nor U6655 (N_6655,N_3446,N_3827);
and U6656 (N_6656,N_3891,N_4565);
and U6657 (N_6657,N_3194,N_5970);
xor U6658 (N_6658,N_4035,N_3301);
xnor U6659 (N_6659,N_3542,N_4238);
or U6660 (N_6660,N_5773,N_3169);
xor U6661 (N_6661,N_3227,N_3034);
or U6662 (N_6662,N_4141,N_3957);
xor U6663 (N_6663,N_5005,N_5318);
and U6664 (N_6664,N_3621,N_3978);
xnor U6665 (N_6665,N_5388,N_4858);
or U6666 (N_6666,N_3502,N_5122);
or U6667 (N_6667,N_5374,N_3398);
or U6668 (N_6668,N_4389,N_4301);
nand U6669 (N_6669,N_5873,N_4324);
xnor U6670 (N_6670,N_4809,N_3415);
nor U6671 (N_6671,N_5036,N_5012);
xnor U6672 (N_6672,N_4016,N_4699);
or U6673 (N_6673,N_4008,N_5033);
xnor U6674 (N_6674,N_4884,N_4526);
and U6675 (N_6675,N_4352,N_4971);
xnor U6676 (N_6676,N_4855,N_4926);
nor U6677 (N_6677,N_5327,N_5619);
xnor U6678 (N_6678,N_3079,N_3886);
xnor U6679 (N_6679,N_5728,N_3630);
xnor U6680 (N_6680,N_3603,N_5594);
nand U6681 (N_6681,N_3976,N_3265);
and U6682 (N_6682,N_5002,N_5351);
nor U6683 (N_6683,N_3722,N_3629);
or U6684 (N_6684,N_4004,N_4846);
nor U6685 (N_6685,N_4935,N_4484);
or U6686 (N_6686,N_3543,N_4653);
or U6687 (N_6687,N_3408,N_4090);
nor U6688 (N_6688,N_4939,N_3073);
xor U6689 (N_6689,N_4677,N_5587);
nor U6690 (N_6690,N_3655,N_4716);
and U6691 (N_6691,N_3444,N_4094);
nand U6692 (N_6692,N_4142,N_5202);
or U6693 (N_6693,N_5414,N_4010);
xnor U6694 (N_6694,N_4754,N_5391);
and U6695 (N_6695,N_5751,N_3864);
or U6696 (N_6696,N_3783,N_3374);
nand U6697 (N_6697,N_3015,N_3678);
or U6698 (N_6698,N_3269,N_4557);
xnor U6699 (N_6699,N_5830,N_5658);
nor U6700 (N_6700,N_5541,N_5859);
or U6701 (N_6701,N_5225,N_3985);
nor U6702 (N_6702,N_3050,N_4722);
nor U6703 (N_6703,N_3877,N_3704);
and U6704 (N_6704,N_3345,N_3197);
nand U6705 (N_6705,N_4030,N_5540);
nand U6706 (N_6706,N_3705,N_5069);
nand U6707 (N_6707,N_4470,N_5812);
nand U6708 (N_6708,N_4207,N_5803);
or U6709 (N_6709,N_5416,N_3421);
and U6710 (N_6710,N_5854,N_5570);
nand U6711 (N_6711,N_4213,N_4026);
nor U6712 (N_6712,N_3742,N_4523);
or U6713 (N_6713,N_3067,N_3845);
nor U6714 (N_6714,N_3257,N_3672);
or U6715 (N_6715,N_4640,N_3422);
or U6716 (N_6716,N_3038,N_5039);
nand U6717 (N_6717,N_3247,N_4087);
nor U6718 (N_6718,N_3691,N_4673);
or U6719 (N_6719,N_4374,N_3029);
or U6720 (N_6720,N_5316,N_3609);
or U6721 (N_6721,N_3068,N_3206);
and U6722 (N_6722,N_4375,N_5526);
nor U6723 (N_6723,N_5319,N_3042);
and U6724 (N_6724,N_3200,N_3790);
xor U6725 (N_6725,N_4423,N_5234);
or U6726 (N_6726,N_4542,N_5971);
or U6727 (N_6727,N_5722,N_5295);
or U6728 (N_6728,N_4548,N_4527);
and U6729 (N_6729,N_5780,N_5322);
nand U6730 (N_6730,N_4309,N_4281);
or U6731 (N_6731,N_5673,N_3840);
nor U6732 (N_6732,N_4553,N_3988);
nand U6733 (N_6733,N_4161,N_4554);
or U6734 (N_6734,N_4514,N_3306);
and U6735 (N_6735,N_5886,N_5076);
and U6736 (N_6736,N_4039,N_5089);
or U6737 (N_6737,N_4800,N_5068);
or U6738 (N_6738,N_5299,N_4255);
and U6739 (N_6739,N_5692,N_3673);
and U6740 (N_6740,N_4692,N_3732);
nand U6741 (N_6741,N_5014,N_3728);
nor U6742 (N_6742,N_5681,N_4076);
and U6743 (N_6743,N_5650,N_5836);
xor U6744 (N_6744,N_4583,N_3510);
nand U6745 (N_6745,N_4996,N_3569);
and U6746 (N_6746,N_4626,N_4410);
xnor U6747 (N_6747,N_3191,N_3481);
or U6748 (N_6748,N_5189,N_3519);
and U6749 (N_6749,N_5713,N_5381);
xor U6750 (N_6750,N_5206,N_3213);
nor U6751 (N_6751,N_3614,N_4268);
and U6752 (N_6752,N_3348,N_4587);
nand U6753 (N_6753,N_3771,N_5642);
xnor U6754 (N_6754,N_3248,N_5677);
and U6755 (N_6755,N_3426,N_4944);
nor U6756 (N_6756,N_4119,N_4605);
xnor U6757 (N_6757,N_4851,N_5400);
nand U6758 (N_6758,N_4995,N_3642);
and U6759 (N_6759,N_5031,N_5732);
xor U6760 (N_6760,N_5777,N_3397);
or U6761 (N_6761,N_4731,N_5077);
xnor U6762 (N_6762,N_5093,N_4664);
nor U6763 (N_6763,N_3048,N_3904);
nor U6764 (N_6764,N_4350,N_3611);
nor U6765 (N_6765,N_4994,N_4180);
xnor U6766 (N_6766,N_4678,N_4837);
and U6767 (N_6767,N_5109,N_4031);
and U6768 (N_6768,N_3593,N_5881);
and U6769 (N_6769,N_4249,N_5904);
and U6770 (N_6770,N_4993,N_3637);
and U6771 (N_6771,N_5789,N_3037);
nand U6772 (N_6772,N_3760,N_5426);
xnor U6773 (N_6773,N_5911,N_5020);
nand U6774 (N_6774,N_4369,N_5682);
nand U6775 (N_6775,N_4627,N_4001);
xnor U6776 (N_6776,N_5083,N_4164);
nand U6777 (N_6777,N_3483,N_4341);
and U6778 (N_6778,N_5905,N_5219);
and U6779 (N_6779,N_4504,N_3958);
nor U6780 (N_6780,N_3851,N_4940);
and U6781 (N_6781,N_4386,N_5995);
nand U6782 (N_6782,N_5090,N_5261);
nor U6783 (N_6783,N_3135,N_3183);
and U6784 (N_6784,N_5270,N_4721);
and U6785 (N_6785,N_4883,N_4942);
and U6786 (N_6786,N_4748,N_5358);
nand U6787 (N_6787,N_3947,N_4436);
or U6788 (N_6788,N_4036,N_3484);
nand U6789 (N_6789,N_5264,N_3900);
xor U6790 (N_6790,N_4270,N_4815);
and U6791 (N_6791,N_4353,N_3407);
nand U6792 (N_6792,N_4295,N_4567);
xor U6793 (N_6793,N_3775,N_4794);
xnor U6794 (N_6794,N_5287,N_3717);
nor U6795 (N_6795,N_4316,N_5672);
or U6796 (N_6796,N_5707,N_5709);
or U6797 (N_6797,N_5297,N_5762);
and U6798 (N_6798,N_5624,N_5368);
nor U6799 (N_6799,N_5827,N_4589);
nand U6800 (N_6800,N_4317,N_4547);
or U6801 (N_6801,N_5352,N_4694);
xor U6802 (N_6802,N_4409,N_4894);
or U6803 (N_6803,N_3515,N_3298);
or U6804 (N_6804,N_4441,N_3973);
xnor U6805 (N_6805,N_4679,N_4337);
or U6806 (N_6806,N_3352,N_4804);
and U6807 (N_6807,N_4747,N_3497);
nor U6808 (N_6808,N_5065,N_3110);
or U6809 (N_6809,N_3684,N_3780);
xor U6810 (N_6810,N_5389,N_5613);
xor U6811 (N_6811,N_3897,N_3369);
or U6812 (N_6812,N_3822,N_3302);
nand U6813 (N_6813,N_4127,N_3351);
xor U6814 (N_6814,N_3129,N_4395);
and U6815 (N_6815,N_5043,N_5485);
nand U6816 (N_6816,N_4580,N_5503);
and U6817 (N_6817,N_4263,N_3763);
nor U6818 (N_6818,N_5727,N_5695);
or U6819 (N_6819,N_4190,N_4980);
and U6820 (N_6820,N_4875,N_3226);
nand U6821 (N_6821,N_3959,N_5277);
nor U6822 (N_6822,N_3088,N_5434);
xor U6823 (N_6823,N_5562,N_4181);
nor U6824 (N_6824,N_4022,N_4623);
or U6825 (N_6825,N_5818,N_4680);
xor U6826 (N_6826,N_5466,N_3671);
xor U6827 (N_6827,N_3690,N_4941);
xnor U6828 (N_6828,N_5519,N_3258);
and U6829 (N_6829,N_3545,N_5066);
nand U6830 (N_6830,N_3734,N_5118);
nand U6831 (N_6831,N_5874,N_4727);
nand U6832 (N_6832,N_5530,N_3122);
and U6833 (N_6833,N_3334,N_3100);
nand U6834 (N_6834,N_3394,N_5564);
and U6835 (N_6835,N_3803,N_4652);
or U6836 (N_6836,N_5662,N_3087);
nor U6837 (N_6837,N_4256,N_4292);
and U6838 (N_6838,N_5580,N_4024);
and U6839 (N_6839,N_4718,N_4307);
and U6840 (N_6840,N_5088,N_4789);
nand U6841 (N_6841,N_3357,N_3833);
nor U6842 (N_6842,N_4743,N_3490);
xor U6843 (N_6843,N_5167,N_5053);
and U6844 (N_6844,N_3086,N_3919);
nor U6845 (N_6845,N_3707,N_5801);
nand U6846 (N_6846,N_5953,N_3557);
xor U6847 (N_6847,N_4783,N_4095);
nor U6848 (N_6848,N_4479,N_4154);
nand U6849 (N_6849,N_5408,N_4379);
xnor U6850 (N_6850,N_3810,N_5003);
xor U6851 (N_6851,N_4532,N_3145);
xnor U6852 (N_6852,N_5821,N_5179);
nor U6853 (N_6853,N_3278,N_4186);
nor U6854 (N_6854,N_5738,N_3618);
nor U6855 (N_6855,N_3273,N_5849);
or U6856 (N_6856,N_3895,N_3800);
and U6857 (N_6857,N_5659,N_3830);
and U6858 (N_6858,N_5686,N_5396);
and U6859 (N_6859,N_4205,N_4266);
xnor U6860 (N_6860,N_5852,N_5579);
or U6861 (N_6861,N_3685,N_4963);
or U6862 (N_6862,N_4541,N_5591);
xor U6863 (N_6863,N_4613,N_5141);
or U6864 (N_6864,N_3952,N_4412);
xor U6865 (N_6865,N_3396,N_3217);
or U6866 (N_6866,N_4961,N_4224);
xor U6867 (N_6867,N_4291,N_5331);
xor U6868 (N_6868,N_3313,N_5670);
and U6869 (N_6869,N_3899,N_4572);
and U6870 (N_6870,N_5870,N_4717);
nand U6871 (N_6871,N_3916,N_5847);
and U6872 (N_6872,N_3442,N_4360);
nand U6873 (N_6873,N_5332,N_5160);
or U6874 (N_6874,N_4519,N_5025);
xnor U6875 (N_6875,N_5671,N_4820);
nor U6876 (N_6876,N_4321,N_3746);
and U6877 (N_6877,N_5983,N_4027);
nor U6878 (N_6878,N_3378,N_3224);
xnor U6879 (N_6879,N_4671,N_5475);
or U6880 (N_6880,N_4089,N_5420);
and U6881 (N_6881,N_5920,N_5851);
xor U6882 (N_6882,N_5649,N_5026);
nor U6883 (N_6883,N_4088,N_5193);
xor U6884 (N_6884,N_3949,N_5590);
xor U6885 (N_6885,N_4539,N_5689);
xor U6886 (N_6886,N_3142,N_5100);
xor U6887 (N_6887,N_3373,N_5447);
nor U6888 (N_6888,N_4868,N_5560);
xnor U6889 (N_6889,N_4364,N_4808);
and U6890 (N_6890,N_3186,N_5258);
nor U6891 (N_6891,N_5730,N_3718);
xnor U6892 (N_6892,N_5330,N_4406);
xnor U6893 (N_6893,N_3708,N_4714);
xor U6894 (N_6894,N_4105,N_4014);
and U6895 (N_6895,N_5778,N_5693);
and U6896 (N_6896,N_5568,N_5047);
xnor U6897 (N_6897,N_4339,N_5776);
nand U6898 (N_6898,N_5763,N_4952);
and U6899 (N_6899,N_4057,N_3143);
nor U6900 (N_6900,N_3929,N_4283);
or U6901 (N_6901,N_4112,N_4297);
or U6902 (N_6902,N_3212,N_5000);
nor U6903 (N_6903,N_4881,N_4767);
or U6904 (N_6904,N_5635,N_4211);
or U6905 (N_6905,N_3364,N_4147);
and U6906 (N_6906,N_5359,N_4054);
nand U6907 (N_6907,N_3229,N_4713);
or U6908 (N_6908,N_3782,N_5545);
nor U6909 (N_6909,N_4111,N_4928);
or U6910 (N_6910,N_4739,N_4362);
xnor U6911 (N_6911,N_3975,N_5132);
xnor U6912 (N_6912,N_3066,N_5783);
nor U6913 (N_6913,N_4707,N_4185);
and U6914 (N_6914,N_3726,N_5453);
and U6915 (N_6915,N_4584,N_3888);
nand U6916 (N_6916,N_3296,N_3107);
and U6917 (N_6917,N_5286,N_4265);
xnor U6918 (N_6918,N_4000,N_3960);
nand U6919 (N_6919,N_5119,N_5979);
nand U6920 (N_6920,N_3766,N_4958);
or U6921 (N_6921,N_4414,N_4314);
xnor U6922 (N_6922,N_4919,N_5675);
and U6923 (N_6923,N_4852,N_3176);
or U6924 (N_6924,N_4648,N_5955);
or U6925 (N_6925,N_4750,N_3930);
and U6926 (N_6926,N_4343,N_5810);
nor U6927 (N_6927,N_5190,N_3078);
and U6928 (N_6928,N_3625,N_4914);
nor U6929 (N_6929,N_5766,N_5794);
nand U6930 (N_6930,N_4472,N_5041);
or U6931 (N_6931,N_5255,N_3638);
nand U6932 (N_6932,N_4490,N_3998);
nor U6933 (N_6933,N_4666,N_5262);
and U6934 (N_6934,N_5915,N_3453);
xor U6935 (N_6935,N_4489,N_5749);
or U6936 (N_6936,N_5977,N_3433);
or U6937 (N_6937,N_5884,N_4874);
or U6938 (N_6938,N_3748,N_4069);
xor U6939 (N_6939,N_3547,N_3812);
nor U6940 (N_6940,N_3349,N_4966);
and U6941 (N_6941,N_3447,N_3376);
and U6942 (N_6942,N_5493,N_5263);
nand U6943 (N_6943,N_4696,N_5968);
nor U6944 (N_6944,N_3606,N_4732);
xnor U6945 (N_6945,N_4209,N_4570);
nor U6946 (N_6946,N_5451,N_5584);
and U6947 (N_6947,N_3482,N_5431);
or U6948 (N_6948,N_4761,N_4799);
or U6949 (N_6949,N_3689,N_3474);
nor U6950 (N_6950,N_3455,N_3026);
nor U6951 (N_6951,N_3493,N_5120);
nor U6952 (N_6952,N_3099,N_3237);
nand U6953 (N_6953,N_5941,N_4282);
or U6954 (N_6954,N_4766,N_3131);
nand U6955 (N_6955,N_4042,N_5515);
xor U6956 (N_6956,N_3233,N_4720);
xor U6957 (N_6957,N_4239,N_4682);
xnor U6958 (N_6958,N_5543,N_3772);
and U6959 (N_6959,N_3377,N_3124);
nand U6960 (N_6960,N_3390,N_5892);
and U6961 (N_6961,N_3715,N_4425);
nor U6962 (N_6962,N_3942,N_3479);
nor U6963 (N_6963,N_4107,N_3171);
nand U6964 (N_6964,N_4236,N_3648);
nand U6965 (N_6965,N_3001,N_5162);
and U6966 (N_6966,N_5430,N_4744);
nand U6967 (N_6967,N_4155,N_5203);
nand U6968 (N_6968,N_3239,N_4267);
and U6969 (N_6969,N_3116,N_5152);
xor U6970 (N_6970,N_4005,N_3314);
nor U6971 (N_6971,N_5062,N_3002);
nor U6972 (N_6972,N_4997,N_5224);
or U6973 (N_6973,N_5676,N_3049);
nand U6974 (N_6974,N_3991,N_5051);
xnor U6975 (N_6975,N_5111,N_3076);
xor U6976 (N_6976,N_5793,N_5490);
nand U6977 (N_6977,N_3411,N_5198);
or U6978 (N_6978,N_3105,N_5392);
nand U6979 (N_6979,N_5017,N_5626);
and U6980 (N_6980,N_3723,N_4402);
xnor U6981 (N_6981,N_4294,N_4071);
and U6982 (N_6982,N_4753,N_4782);
or U6983 (N_6983,N_5567,N_5427);
or U6984 (N_6984,N_5232,N_3516);
or U6985 (N_6985,N_3992,N_3509);
xnor U6986 (N_6986,N_5312,N_4609);
xnor U6987 (N_6987,N_3633,N_4168);
xor U6988 (N_6988,N_3198,N_3104);
or U6989 (N_6989,N_3555,N_3488);
nor U6990 (N_6990,N_4037,N_5375);
xor U6991 (N_6991,N_4326,N_4763);
and U6992 (N_6992,N_4422,N_4624);
nand U6993 (N_6993,N_4230,N_4109);
nor U6994 (N_6994,N_5944,N_3902);
nor U6995 (N_6995,N_5933,N_5684);
and U6996 (N_6996,N_4433,N_5361);
or U6997 (N_6997,N_5501,N_3676);
nor U6998 (N_6998,N_4053,N_3172);
or U6999 (N_6999,N_3935,N_4909);
nand U7000 (N_7000,N_4500,N_5589);
xor U7001 (N_7001,N_5539,N_4121);
nor U7002 (N_7002,N_5376,N_3798);
xnor U7003 (N_7003,N_5128,N_3148);
nor U7004 (N_7004,N_3620,N_3341);
nor U7005 (N_7005,N_3908,N_3228);
xnor U7006 (N_7006,N_3647,N_4841);
xor U7007 (N_7007,N_5114,N_5142);
or U7008 (N_7008,N_3546,N_3565);
or U7009 (N_7009,N_5809,N_4288);
and U7010 (N_7010,N_4876,N_3052);
xnor U7011 (N_7011,N_4454,N_5625);
or U7012 (N_7012,N_5586,N_5600);
nor U7013 (N_7013,N_4685,N_4774);
nor U7014 (N_7014,N_4645,N_4043);
and U7015 (N_7015,N_5172,N_3740);
and U7016 (N_7016,N_4222,N_5021);
xnor U7017 (N_7017,N_5075,N_5470);
nor U7018 (N_7018,N_3495,N_5059);
nand U7019 (N_7019,N_5518,N_4525);
and U7020 (N_7020,N_4888,N_3011);
or U7021 (N_7021,N_5664,N_4132);
xor U7022 (N_7022,N_5875,N_3220);
xor U7023 (N_7023,N_3848,N_4938);
nand U7024 (N_7024,N_5458,N_3494);
and U7025 (N_7025,N_4248,N_4182);
and U7026 (N_7026,N_3744,N_4312);
xor U7027 (N_7027,N_5791,N_3882);
nand U7028 (N_7028,N_4848,N_5045);
or U7029 (N_7029,N_3592,N_5278);
and U7030 (N_7030,N_3289,N_3267);
xnor U7031 (N_7031,N_4396,N_3599);
xnor U7032 (N_7032,N_4972,N_3454);
xor U7033 (N_7033,N_4146,N_4100);
and U7034 (N_7034,N_3080,N_4843);
nand U7035 (N_7035,N_5857,N_4349);
xnor U7036 (N_7036,N_4174,N_4602);
and U7037 (N_7037,N_3626,N_5967);
or U7038 (N_7038,N_5148,N_4700);
nand U7039 (N_7039,N_5993,N_3309);
and U7040 (N_7040,N_3462,N_5688);
nand U7041 (N_7041,N_3175,N_3863);
nor U7042 (N_7042,N_5826,N_5754);
nand U7043 (N_7043,N_3853,N_5938);
and U7044 (N_7044,N_4687,N_4657);
nand U7045 (N_7045,N_3041,N_4286);
and U7046 (N_7046,N_5409,N_4498);
nand U7047 (N_7047,N_5907,N_4975);
nor U7048 (N_7048,N_5928,N_3596);
nor U7049 (N_7049,N_4377,N_3476);
nand U7050 (N_7050,N_3254,N_5825);
and U7051 (N_7051,N_4503,N_3777);
and U7052 (N_7052,N_4191,N_5737);
xor U7053 (N_7053,N_4965,N_3841);
or U7054 (N_7054,N_4096,N_5990);
xor U7055 (N_7055,N_3040,N_4219);
nand U7056 (N_7056,N_5313,N_5240);
and U7057 (N_7057,N_5656,N_3173);
nand U7058 (N_7058,N_3712,N_4446);
nand U7059 (N_7059,N_5106,N_3750);
nor U7060 (N_7060,N_3837,N_4522);
nor U7061 (N_7061,N_5333,N_3303);
nor U7062 (N_7062,N_4254,N_4950);
nor U7063 (N_7063,N_3264,N_4577);
or U7064 (N_7064,N_5018,N_3114);
and U7065 (N_7065,N_4697,N_3465);
xor U7066 (N_7066,N_4342,N_3065);
nand U7067 (N_7067,N_3043,N_4537);
nor U7068 (N_7068,N_3457,N_4049);
or U7069 (N_7069,N_4451,N_5839);
and U7070 (N_7070,N_5086,N_5757);
nor U7071 (N_7071,N_5230,N_4781);
and U7072 (N_7072,N_5393,N_5081);
nor U7073 (N_7073,N_5855,N_5082);
xor U7074 (N_7074,N_4113,N_4546);
xnor U7075 (N_7075,N_5415,N_5731);
nand U7076 (N_7076,N_4608,N_5110);
nor U7077 (N_7077,N_5085,N_3016);
nor U7078 (N_7078,N_4803,N_3291);
and U7079 (N_7079,N_5221,N_4686);
and U7080 (N_7080,N_5452,N_3018);
and U7081 (N_7081,N_3954,N_5637);
nor U7082 (N_7082,N_4690,N_4183);
nand U7083 (N_7083,N_5929,N_3784);
nand U7084 (N_7084,N_4735,N_3953);
nand U7085 (N_7085,N_5161,N_3320);
xor U7086 (N_7086,N_4771,N_4033);
nand U7087 (N_7087,N_4741,N_5267);
nand U7088 (N_7088,N_5308,N_3836);
or U7089 (N_7089,N_5576,N_4705);
and U7090 (N_7090,N_4474,N_5342);
or U7091 (N_7091,N_4610,N_3084);
nand U7092 (N_7092,N_3182,N_5371);
nand U7093 (N_7093,N_3432,N_5621);
xor U7094 (N_7094,N_3709,N_3528);
nand U7095 (N_7095,N_5471,N_4656);
nand U7096 (N_7096,N_3719,N_5253);
nand U7097 (N_7097,N_3664,N_4072);
nand U7098 (N_7098,N_4074,N_4382);
and U7099 (N_7099,N_3738,N_3602);
xnor U7100 (N_7100,N_4507,N_5865);
nor U7101 (N_7101,N_5973,N_5196);
nand U7102 (N_7102,N_3340,N_3424);
or U7103 (N_7103,N_5894,N_3125);
nor U7104 (N_7104,N_4456,N_3623);
nor U7105 (N_7105,N_4407,N_4355);
nor U7106 (N_7106,N_5223,N_3402);
nor U7107 (N_7107,N_4900,N_3996);
and U7108 (N_7108,N_3232,N_4977);
xor U7109 (N_7109,N_3356,N_5813);
or U7110 (N_7110,N_5450,N_4857);
nor U7111 (N_7111,N_5476,N_5443);
xnor U7112 (N_7112,N_5942,N_4573);
or U7113 (N_7113,N_5756,N_4041);
nor U7114 (N_7114,N_4417,N_4590);
xnor U7115 (N_7115,N_3608,N_5506);
and U7116 (N_7116,N_3256,N_5174);
and U7117 (N_7117,N_3680,N_4032);
xnor U7118 (N_7118,N_4825,N_5862);
or U7119 (N_7119,N_4497,N_3939);
and U7120 (N_7120,N_3460,N_5623);
xnor U7121 (N_7121,N_5272,N_3525);
nor U7122 (N_7122,N_5581,N_4328);
nor U7123 (N_7123,N_4611,N_4601);
and U7124 (N_7124,N_4299,N_5797);
nor U7125 (N_7125,N_4345,N_5620);
xor U7126 (N_7126,N_4229,N_4131);
or U7127 (N_7127,N_3459,N_3414);
and U7128 (N_7128,N_3604,N_5829);
and U7129 (N_7129,N_5007,N_4983);
nor U7130 (N_7130,N_4835,N_5856);
nand U7131 (N_7131,N_3058,N_4333);
and U7132 (N_7132,N_4358,N_4706);
or U7133 (N_7133,N_5976,N_4989);
nor U7134 (N_7134,N_3640,N_4158);
nor U7135 (N_7135,N_5529,N_4688);
nand U7136 (N_7136,N_3218,N_5946);
nand U7137 (N_7137,N_3553,N_4221);
or U7138 (N_7138,N_3335,N_5403);
xor U7139 (N_7139,N_4480,N_3091);
nand U7140 (N_7140,N_3767,N_5696);
and U7141 (N_7141,N_3284,N_3520);
nor U7142 (N_7142,N_5029,N_4691);
and U7143 (N_7143,N_3653,N_4636);
xor U7144 (N_7144,N_4323,N_3371);
xnor U7145 (N_7145,N_3971,N_4468);
nand U7146 (N_7146,N_4156,N_5969);
nand U7147 (N_7147,N_5736,N_5743);
xnor U7148 (N_7148,N_4758,N_4455);
nor U7149 (N_7149,N_5143,N_5155);
nand U7150 (N_7150,N_5239,N_4896);
and U7151 (N_7151,N_3982,N_3752);
nor U7152 (N_7152,N_5474,N_3321);
and U7153 (N_7153,N_3550,N_5060);
xor U7154 (N_7154,N_3880,N_5436);
and U7155 (N_7155,N_3858,N_3558);
nor U7156 (N_7156,N_4772,N_5523);
and U7157 (N_7157,N_5544,N_4062);
nand U7158 (N_7158,N_5512,N_3912);
nor U7159 (N_7159,N_4373,N_3319);
and U7160 (N_7160,N_3283,N_5759);
xnor U7161 (N_7161,N_3688,N_3944);
xnor U7162 (N_7162,N_5947,N_3272);
nor U7163 (N_7163,N_3024,N_5807);
and U7164 (N_7164,N_3108,N_5105);
xnor U7165 (N_7165,N_4064,N_3255);
nand U7166 (N_7166,N_4889,N_5956);
or U7167 (N_7167,N_3251,N_3252);
and U7168 (N_7168,N_5504,N_5717);
xor U7169 (N_7169,N_4011,N_3149);
and U7170 (N_7170,N_4354,N_4925);
and U7171 (N_7171,N_4411,N_3500);
nand U7172 (N_7172,N_5569,N_4184);
or U7173 (N_7173,N_5853,N_3701);
and U7174 (N_7174,N_4985,N_5511);
xor U7175 (N_7175,N_5317,N_5432);
xnor U7176 (N_7176,N_5814,N_4964);
or U7177 (N_7177,N_4212,N_4509);
nor U7178 (N_7178,N_5663,N_4684);
xnor U7179 (N_7179,N_5460,N_3410);
and U7180 (N_7180,N_4197,N_4818);
nor U7181 (N_7181,N_5602,N_4893);
and U7182 (N_7182,N_4013,N_3342);
and U7183 (N_7183,N_4469,N_5887);
or U7184 (N_7184,N_4023,N_4415);
xor U7185 (N_7185,N_3055,N_4202);
nor U7186 (N_7186,N_3724,N_5733);
xor U7187 (N_7187,N_3683,N_4955);
xnor U7188 (N_7188,N_4674,N_4303);
and U7189 (N_7189,N_3703,N_3847);
nor U7190 (N_7190,N_5514,N_5296);
or U7191 (N_7191,N_5654,N_3570);
and U7192 (N_7192,N_3905,N_4556);
xnor U7193 (N_7193,N_4372,N_4521);
nor U7194 (N_7194,N_4276,N_5972);
nand U7195 (N_7195,N_4967,N_4907);
nor U7196 (N_7196,N_3420,N_3898);
and U7197 (N_7197,N_5498,N_5417);
xor U7198 (N_7198,N_3696,N_3711);
and U7199 (N_7199,N_4117,N_5687);
and U7200 (N_7200,N_3316,N_5917);
or U7201 (N_7201,N_4080,N_4505);
nand U7202 (N_7202,N_3401,N_3818);
and U7203 (N_7203,N_4604,N_3140);
nor U7204 (N_7204,N_5199,N_5786);
nand U7205 (N_7205,N_5329,N_5571);
and U7206 (N_7206,N_5363,N_3588);
or U7207 (N_7207,N_5011,N_5285);
nor U7208 (N_7208,N_5878,N_4081);
or U7209 (N_7209,N_3811,N_5163);
or U7210 (N_7210,N_5999,N_4520);
nor U7211 (N_7211,N_5644,N_4902);
xor U7212 (N_7212,N_5355,N_3266);
nor U7213 (N_7213,N_4018,N_3657);
xnor U7214 (N_7214,N_5215,N_4361);
nand U7215 (N_7215,N_4897,N_5715);
nor U7216 (N_7216,N_4051,N_4531);
and U7217 (N_7217,N_4399,N_4619);
and U7218 (N_7218,N_4934,N_5555);
or U7219 (N_7219,N_4366,N_3868);
or U7220 (N_7220,N_3589,N_4225);
nor U7221 (N_7221,N_4487,N_3472);
and U7222 (N_7222,N_4259,N_5382);
nor U7223 (N_7223,N_3115,N_3652);
xor U7224 (N_7224,N_3486,N_3163);
nor U7225 (N_7225,N_4319,N_4834);
nand U7226 (N_7226,N_3961,N_4278);
xnor U7227 (N_7227,N_5042,N_5645);
or U7228 (N_7228,N_5217,N_3053);
or U7229 (N_7229,N_5963,N_5500);
nand U7230 (N_7230,N_4737,N_4144);
or U7231 (N_7231,N_4854,N_5323);
and U7232 (N_7232,N_5413,N_5170);
xnor U7233 (N_7233,N_3094,N_5095);
xnor U7234 (N_7234,N_4097,N_5404);
nand U7235 (N_7235,N_5890,N_5698);
xnor U7236 (N_7236,N_4149,N_5599);
or U7237 (N_7237,N_5078,N_4421);
or U7238 (N_7238,N_3249,N_3240);
and U7239 (N_7239,N_4118,N_3441);
nand U7240 (N_7240,N_3867,N_4210);
or U7241 (N_7241,N_4899,N_3923);
xor U7242 (N_7242,N_5377,N_4385);
and U7243 (N_7243,N_3801,N_4947);
nand U7244 (N_7244,N_5536,N_4235);
nand U7245 (N_7245,N_3400,N_5711);
xor U7246 (N_7246,N_3725,N_5768);
or U7247 (N_7247,N_3758,N_3430);
nand U7248 (N_7248,N_4464,N_3417);
and U7249 (N_7249,N_3821,N_3202);
xnor U7250 (N_7250,N_4038,N_5321);
nor U7251 (N_7251,N_3523,N_5405);
and U7252 (N_7252,N_5437,N_4831);
and U7253 (N_7253,N_3275,N_5192);
or U7254 (N_7254,N_4724,N_4232);
nand U7255 (N_7255,N_4734,N_5781);
and U7256 (N_7256,N_5691,N_5099);
or U7257 (N_7257,N_4838,N_4641);
nand U7258 (N_7258,N_5302,N_5425);
xor U7259 (N_7259,N_3263,N_3538);
or U7260 (N_7260,N_4728,N_5438);
nor U7261 (N_7261,N_3166,N_4179);
xnor U7262 (N_7262,N_5032,N_5563);
and U7263 (N_7263,N_4073,N_5860);
and U7264 (N_7264,N_5237,N_3674);
and U7265 (N_7265,N_5522,N_3582);
and U7266 (N_7266,N_5357,N_5309);
or U7267 (N_7267,N_5665,N_3021);
nand U7268 (N_7268,N_3081,N_4140);
and U7269 (N_7269,N_4733,N_4060);
nor U7270 (N_7270,N_5502,N_4822);
and U7271 (N_7271,N_3789,N_3469);
or U7272 (N_7272,N_3872,N_4227);
nor U7273 (N_7273,N_5164,N_4629);
or U7274 (N_7274,N_4061,N_4581);
or U7275 (N_7275,N_5922,N_4163);
or U7276 (N_7276,N_3133,N_4953);
nand U7277 (N_7277,N_3180,N_5260);
xor U7278 (N_7278,N_4778,N_3384);
or U7279 (N_7279,N_3023,N_5194);
and U7280 (N_7280,N_3450,N_5271);
and U7281 (N_7281,N_4845,N_5440);
nand U7282 (N_7282,N_4524,N_5010);
or U7283 (N_7283,N_5850,N_3983);
or U7284 (N_7284,N_4918,N_4285);
xnor U7285 (N_7285,N_3741,N_3156);
or U7286 (N_7286,N_5133,N_5373);
nand U7287 (N_7287,N_5770,N_5542);
and U7288 (N_7288,N_4159,N_3552);
nor U7289 (N_7289,N_4092,N_4816);
nor U7290 (N_7290,N_4296,N_3338);
nand U7291 (N_7291,N_5811,N_5747);
nor U7292 (N_7292,N_4305,N_4625);
nand U7293 (N_7293,N_4289,N_3214);
nor U7294 (N_7294,N_4320,N_3670);
nor U7295 (N_7295,N_4806,N_5535);
or U7296 (N_7296,N_5725,N_3799);
nand U7297 (N_7297,N_3539,N_5016);
and U7298 (N_7298,N_3009,N_4365);
xnor U7299 (N_7299,N_3540,N_5932);
xnor U7300 (N_7300,N_4936,N_4618);
nor U7301 (N_7301,N_5951,N_3077);
and U7302 (N_7302,N_3561,N_4948);
or U7303 (N_7303,N_4048,N_3221);
or U7304 (N_7304,N_3330,N_3059);
nand U7305 (N_7305,N_5320,N_4579);
xor U7306 (N_7306,N_3813,N_3883);
or U7307 (N_7307,N_5912,N_4957);
nand U7308 (N_7308,N_4439,N_3788);
xor U7309 (N_7309,N_3210,N_4242);
nand U7310 (N_7310,N_3622,N_3507);
and U7311 (N_7311,N_3879,N_5472);
xnor U7312 (N_7312,N_5275,N_3607);
and U7313 (N_7313,N_4593,N_3969);
and U7314 (N_7314,N_3999,N_3580);
nor U7315 (N_7315,N_5429,N_3174);
nor U7316 (N_7316,N_3489,N_3234);
xor U7317 (N_7317,N_3535,N_5123);
and U7318 (N_7318,N_3755,N_4250);
nand U7319 (N_7319,N_5633,N_5806);
nor U7320 (N_7320,N_3769,N_5168);
or U7321 (N_7321,N_4904,N_3928);
nand U7322 (N_7322,N_4943,N_3871);
xnor U7323 (N_7323,N_3651,N_3656);
or U7324 (N_7324,N_4576,N_4596);
or U7325 (N_7325,N_5610,N_4218);
xnor U7326 (N_7326,N_5868,N_3118);
and U7327 (N_7327,N_4921,N_5708);
nand U7328 (N_7328,N_3325,N_4905);
nand U7329 (N_7329,N_5595,N_4444);
or U7330 (N_7330,N_3025,N_4138);
xnor U7331 (N_7331,N_3231,N_5831);
nor U7332 (N_7332,N_3809,N_4269);
nand U7333 (N_7333,N_5802,N_4430);
nor U7334 (N_7334,N_5651,N_5559);
or U7335 (N_7335,N_3815,N_5188);
nor U7336 (N_7336,N_3161,N_4824);
nand U7337 (N_7337,N_4082,N_3412);
nor U7338 (N_7338,N_4114,N_4978);
nor U7339 (N_7339,N_5746,N_3120);
xnor U7340 (N_7340,N_3838,N_5137);
nand U7341 (N_7341,N_3022,N_3962);
nand U7342 (N_7342,N_3571,N_4199);
nor U7343 (N_7343,N_5290,N_3354);
xor U7344 (N_7344,N_3368,N_3549);
xor U7345 (N_7345,N_4821,N_4106);
xor U7346 (N_7346,N_4058,N_3192);
xnor U7347 (N_7347,N_4779,N_4099);
or U7348 (N_7348,N_4882,N_4807);
xnor U7349 (N_7349,N_3339,N_4139);
and U7350 (N_7350,N_3665,N_3628);
nor U7351 (N_7351,N_5582,N_5876);
or U7352 (N_7352,N_5101,N_4860);
or U7353 (N_7353,N_3126,N_5690);
nor U7354 (N_7354,N_5274,N_3754);
or U7355 (N_7355,N_4371,N_5609);
nand U7356 (N_7356,N_3141,N_4293);
and U7357 (N_7357,N_5607,N_3832);
nor U7358 (N_7358,N_4070,N_4559);
nand U7359 (N_7359,N_5055,N_5139);
and U7360 (N_7360,N_4136,N_5548);
and U7361 (N_7361,N_5380,N_3605);
nor U7362 (N_7362,N_4729,N_5638);
or U7363 (N_7363,N_5877,N_3936);
or U7364 (N_7364,N_4017,N_4204);
or U7365 (N_7365,N_3147,N_4135);
nor U7366 (N_7366,N_4859,N_4638);
nand U7367 (N_7367,N_3355,N_3268);
nor U7368 (N_7368,N_3941,N_5157);
or U7369 (N_7369,N_4805,N_5345);
nor U7370 (N_7370,N_3938,N_3152);
or U7371 (N_7371,N_3757,N_3324);
or U7372 (N_7372,N_5872,N_4660);
or U7373 (N_7373,N_3568,N_5585);
nor U7374 (N_7374,N_5661,N_5775);
nor U7375 (N_7375,N_3317,N_4516);
or U7376 (N_7376,N_3250,N_3713);
nor U7377 (N_7377,N_3184,N_5153);
and U7378 (N_7378,N_5169,N_4481);
xnor U7379 (N_7379,N_5937,N_5647);
and U7380 (N_7380,N_5496,N_5473);
nor U7381 (N_7381,N_5244,N_4764);
nand U7382 (N_7382,N_4332,N_5936);
nand U7383 (N_7383,N_5370,N_4401);
nand U7384 (N_7384,N_4667,N_5608);
and U7385 (N_7385,N_4440,N_3729);
nand U7386 (N_7386,N_4450,N_5328);
or U7387 (N_7387,N_5136,N_3017);
or U7388 (N_7388,N_3911,N_5573);
nand U7389 (N_7389,N_3162,N_4200);
xnor U7390 (N_7390,N_5981,N_4148);
xnor U7391 (N_7391,N_4908,N_4861);
or U7392 (N_7392,N_5091,N_5338);
and U7393 (N_7393,N_4873,N_5165);
xnor U7394 (N_7394,N_3096,N_5001);
nor U7395 (N_7395,N_5340,N_5159);
and U7396 (N_7396,N_4811,N_5048);
xor U7397 (N_7397,N_3160,N_4448);
and U7398 (N_7398,N_5491,N_5943);
xor U7399 (N_7399,N_3699,N_5256);
nor U7400 (N_7400,N_3028,N_4788);
nor U7401 (N_7401,N_3965,N_4865);
and U7402 (N_7402,N_4723,N_3661);
or U7403 (N_7403,N_5494,N_4196);
and U7404 (N_7404,N_4346,N_3922);
nor U7405 (N_7405,N_5112,N_3522);
or U7406 (N_7406,N_4445,N_4757);
and U7407 (N_7407,N_3889,N_5641);
nor U7408 (N_7408,N_3230,N_4973);
or U7409 (N_7409,N_5516,N_3057);
or U7410 (N_7410,N_3196,N_3039);
or U7411 (N_7411,N_5988,N_5127);
or U7412 (N_7412,N_3835,N_4128);
nor U7413 (N_7413,N_5231,N_4920);
and U7414 (N_7414,N_4649,N_3155);
nand U7415 (N_7415,N_5383,N_5293);
nor U7416 (N_7416,N_4175,N_5463);
nand U7417 (N_7417,N_4310,N_5547);
nor U7418 (N_7418,N_5087,N_3955);
and U7419 (N_7419,N_4397,N_3521);
or U7420 (N_7420,N_3892,N_4533);
xnor U7421 (N_7421,N_3069,N_4712);
nor U7422 (N_7422,N_4828,N_4913);
and U7423 (N_7423,N_4643,N_3924);
xnor U7424 (N_7424,N_4002,N_5939);
or U7425 (N_7425,N_3619,N_5940);
nor U7426 (N_7426,N_3137,N_3128);
or U7427 (N_7427,N_3598,N_3293);
nor U7428 (N_7428,N_4240,N_5819);
or U7429 (N_7429,N_5772,N_5056);
nor U7430 (N_7430,N_3610,N_3070);
and U7431 (N_7431,N_3776,N_5303);
and U7432 (N_7432,N_5588,N_3964);
xor U7433 (N_7433,N_4628,N_5910);
and U7434 (N_7434,N_5004,N_5724);
and U7435 (N_7435,N_5456,N_5994);
or U7436 (N_7436,N_4157,N_5422);
and U7437 (N_7437,N_4491,N_3179);
and U7438 (N_7438,N_3318,N_4134);
nor U7439 (N_7439,N_3575,N_4007);
xnor U7440 (N_7440,N_4351,N_4290);
or U7441 (N_7441,N_5197,N_3089);
nand U7442 (N_7442,N_4998,N_5488);
xnor U7443 (N_7443,N_3304,N_5478);
nor U7444 (N_7444,N_5063,N_5908);
xor U7445 (N_7445,N_3807,N_4574);
nor U7446 (N_7446,N_5130,N_4603);
or U7447 (N_7447,N_5719,N_4898);
nor U7448 (N_7448,N_4203,N_5134);
and U7449 (N_7449,N_5900,N_3733);
or U7450 (N_7450,N_3336,N_5913);
xor U7451 (N_7451,N_3013,N_4528);
xor U7452 (N_7452,N_5714,N_5084);
xor U7453 (N_7453,N_5974,N_4243);
xnor U7454 (N_7454,N_5242,N_5058);
xnor U7455 (N_7455,N_4564,N_5565);
xor U7456 (N_7456,N_3824,N_3347);
and U7457 (N_7457,N_5534,N_4676);
or U7458 (N_7458,N_4984,N_4578);
nand U7459 (N_7459,N_3503,N_3862);
or U7460 (N_7460,N_4166,N_3468);
nor U7461 (N_7461,N_4745,N_5149);
or U7462 (N_7462,N_4394,N_5311);
and U7463 (N_7463,N_5233,N_3692);
nand U7464 (N_7464,N_4917,N_3360);
xor U7465 (N_7465,N_3966,N_3739);
nand U7466 (N_7466,N_5616,N_3632);
and U7467 (N_7467,N_4457,N_5259);
nor U7468 (N_7468,N_5537,N_3660);
nand U7469 (N_7469,N_3634,N_5767);
nor U7470 (N_7470,N_4078,N_5044);
nor U7471 (N_7471,N_3270,N_3092);
or U7472 (N_7472,N_4752,N_4496);
nor U7473 (N_7473,N_3242,N_3694);
nor U7474 (N_7474,N_3875,N_4400);
or U7475 (N_7475,N_4862,N_4424);
or U7476 (N_7476,N_5808,N_5804);
or U7477 (N_7477,N_3036,N_3312);
nor U7478 (N_7478,N_3844,N_3423);
xor U7479 (N_7479,N_3932,N_5891);
nand U7480 (N_7480,N_5057,N_3901);
nor U7481 (N_7481,N_4655,N_5433);
and U7482 (N_7482,N_5592,N_5636);
nand U7483 (N_7483,N_3294,N_4560);
nor U7484 (N_7484,N_3762,N_4518);
nand U7485 (N_7485,N_4273,N_5508);
nand U7486 (N_7486,N_4719,N_4797);
nand U7487 (N_7487,N_3532,N_4391);
or U7488 (N_7488,N_4930,N_4768);
or U7489 (N_7489,N_3382,N_5214);
or U7490 (N_7490,N_5721,N_3223);
or U7491 (N_7491,N_5102,N_5924);
and U7492 (N_7492,N_4639,N_5612);
and U7493 (N_7493,N_5251,N_3295);
or U7494 (N_7494,N_3583,N_4910);
and U7495 (N_7495,N_3624,N_3530);
nand U7496 (N_7496,N_5521,N_4592);
or U7497 (N_7497,N_3323,N_5741);
or U7498 (N_7498,N_5723,N_4912);
xor U7499 (N_7499,N_3679,N_4658);
nand U7500 (N_7500,N_4957,N_4357);
nand U7501 (N_7501,N_5450,N_4566);
nor U7502 (N_7502,N_4655,N_5099);
and U7503 (N_7503,N_4530,N_4782);
and U7504 (N_7504,N_5885,N_4254);
nand U7505 (N_7505,N_4696,N_4231);
nand U7506 (N_7506,N_5193,N_4207);
or U7507 (N_7507,N_4401,N_5880);
and U7508 (N_7508,N_3267,N_4994);
and U7509 (N_7509,N_5299,N_4087);
nor U7510 (N_7510,N_3425,N_4365);
and U7511 (N_7511,N_4201,N_5698);
xor U7512 (N_7512,N_4908,N_5705);
nor U7513 (N_7513,N_3781,N_3611);
nand U7514 (N_7514,N_5688,N_5852);
nand U7515 (N_7515,N_4018,N_5154);
and U7516 (N_7516,N_3653,N_5679);
nor U7517 (N_7517,N_3507,N_5030);
nand U7518 (N_7518,N_4394,N_4681);
and U7519 (N_7519,N_5454,N_4659);
nand U7520 (N_7520,N_4004,N_4439);
xor U7521 (N_7521,N_3789,N_3682);
xnor U7522 (N_7522,N_3348,N_5620);
nor U7523 (N_7523,N_5087,N_5658);
nor U7524 (N_7524,N_5790,N_5973);
or U7525 (N_7525,N_5195,N_5828);
xnor U7526 (N_7526,N_4415,N_5839);
xnor U7527 (N_7527,N_3608,N_5600);
or U7528 (N_7528,N_5200,N_5965);
or U7529 (N_7529,N_5930,N_3568);
nand U7530 (N_7530,N_4288,N_5176);
xor U7531 (N_7531,N_5074,N_3040);
and U7532 (N_7532,N_5227,N_5005);
nor U7533 (N_7533,N_4567,N_3760);
or U7534 (N_7534,N_3690,N_3183);
xor U7535 (N_7535,N_3688,N_4326);
or U7536 (N_7536,N_3584,N_4188);
xor U7537 (N_7537,N_5578,N_3956);
nor U7538 (N_7538,N_5132,N_4619);
nor U7539 (N_7539,N_3765,N_4202);
nand U7540 (N_7540,N_5149,N_4692);
or U7541 (N_7541,N_5936,N_4549);
nand U7542 (N_7542,N_5360,N_4864);
and U7543 (N_7543,N_3310,N_5598);
or U7544 (N_7544,N_4525,N_5243);
and U7545 (N_7545,N_3961,N_5640);
or U7546 (N_7546,N_5373,N_3872);
or U7547 (N_7547,N_4098,N_3366);
nand U7548 (N_7548,N_5508,N_4823);
nand U7549 (N_7549,N_4177,N_5935);
nor U7550 (N_7550,N_4920,N_4551);
and U7551 (N_7551,N_5060,N_3060);
or U7552 (N_7552,N_4086,N_4432);
nor U7553 (N_7553,N_4429,N_3758);
xor U7554 (N_7554,N_4147,N_4453);
or U7555 (N_7555,N_4264,N_5403);
or U7556 (N_7556,N_5264,N_3699);
xnor U7557 (N_7557,N_5258,N_5939);
nand U7558 (N_7558,N_3293,N_5651);
or U7559 (N_7559,N_4759,N_5266);
nand U7560 (N_7560,N_3641,N_3566);
nor U7561 (N_7561,N_5955,N_5699);
nand U7562 (N_7562,N_4590,N_5211);
nor U7563 (N_7563,N_4776,N_4662);
nor U7564 (N_7564,N_3235,N_3016);
nor U7565 (N_7565,N_3438,N_4461);
nand U7566 (N_7566,N_5189,N_5595);
or U7567 (N_7567,N_5680,N_3075);
nand U7568 (N_7568,N_3057,N_3020);
nand U7569 (N_7569,N_3848,N_4860);
xor U7570 (N_7570,N_4452,N_5991);
or U7571 (N_7571,N_3019,N_4823);
and U7572 (N_7572,N_5665,N_5448);
or U7573 (N_7573,N_5222,N_4473);
or U7574 (N_7574,N_4222,N_5527);
nor U7575 (N_7575,N_4206,N_5659);
xnor U7576 (N_7576,N_4552,N_3863);
nor U7577 (N_7577,N_5672,N_3214);
nand U7578 (N_7578,N_5639,N_3756);
nand U7579 (N_7579,N_4554,N_5195);
nand U7580 (N_7580,N_5142,N_4047);
nor U7581 (N_7581,N_3082,N_3415);
or U7582 (N_7582,N_5696,N_4032);
nand U7583 (N_7583,N_4948,N_4685);
nor U7584 (N_7584,N_4387,N_4903);
xnor U7585 (N_7585,N_4738,N_4202);
and U7586 (N_7586,N_4641,N_3342);
or U7587 (N_7587,N_5975,N_5910);
and U7588 (N_7588,N_4164,N_5180);
xnor U7589 (N_7589,N_4211,N_3655);
nand U7590 (N_7590,N_5013,N_5811);
xnor U7591 (N_7591,N_4973,N_3082);
and U7592 (N_7592,N_4774,N_3591);
or U7593 (N_7593,N_5319,N_4770);
xor U7594 (N_7594,N_4262,N_5356);
xor U7595 (N_7595,N_5916,N_4111);
and U7596 (N_7596,N_5836,N_3913);
and U7597 (N_7597,N_3619,N_5077);
xnor U7598 (N_7598,N_5597,N_5397);
or U7599 (N_7599,N_5412,N_5581);
xnor U7600 (N_7600,N_3301,N_3967);
xor U7601 (N_7601,N_3340,N_5251);
and U7602 (N_7602,N_3964,N_4338);
nor U7603 (N_7603,N_5138,N_4028);
nand U7604 (N_7604,N_3044,N_4645);
and U7605 (N_7605,N_4211,N_3749);
or U7606 (N_7606,N_5707,N_4129);
xor U7607 (N_7607,N_5026,N_3931);
nor U7608 (N_7608,N_4030,N_4677);
nor U7609 (N_7609,N_4675,N_5663);
and U7610 (N_7610,N_4316,N_5146);
nor U7611 (N_7611,N_4303,N_4143);
nand U7612 (N_7612,N_5100,N_4387);
and U7613 (N_7613,N_3624,N_4602);
xnor U7614 (N_7614,N_5462,N_5860);
or U7615 (N_7615,N_4020,N_5160);
nand U7616 (N_7616,N_5631,N_4617);
or U7617 (N_7617,N_3386,N_4346);
xnor U7618 (N_7618,N_3475,N_4122);
nor U7619 (N_7619,N_4685,N_3948);
and U7620 (N_7620,N_3467,N_4266);
or U7621 (N_7621,N_3300,N_4430);
nor U7622 (N_7622,N_4592,N_5062);
nor U7623 (N_7623,N_5873,N_5902);
xnor U7624 (N_7624,N_3154,N_3130);
or U7625 (N_7625,N_5280,N_3364);
and U7626 (N_7626,N_4585,N_3676);
nand U7627 (N_7627,N_4338,N_4866);
and U7628 (N_7628,N_3428,N_3140);
xnor U7629 (N_7629,N_3423,N_4821);
nor U7630 (N_7630,N_3097,N_3479);
nor U7631 (N_7631,N_3154,N_3714);
or U7632 (N_7632,N_5394,N_3337);
xnor U7633 (N_7633,N_3620,N_4692);
nand U7634 (N_7634,N_4990,N_4164);
nand U7635 (N_7635,N_3657,N_4225);
nor U7636 (N_7636,N_4709,N_3945);
and U7637 (N_7637,N_3022,N_5988);
and U7638 (N_7638,N_5581,N_5153);
xor U7639 (N_7639,N_5726,N_4304);
or U7640 (N_7640,N_5973,N_4727);
xnor U7641 (N_7641,N_3424,N_4562);
nand U7642 (N_7642,N_4035,N_3181);
xor U7643 (N_7643,N_3775,N_3846);
and U7644 (N_7644,N_5684,N_3074);
or U7645 (N_7645,N_4598,N_3728);
and U7646 (N_7646,N_5132,N_5635);
or U7647 (N_7647,N_5652,N_4963);
and U7648 (N_7648,N_3489,N_4961);
and U7649 (N_7649,N_5045,N_5784);
xnor U7650 (N_7650,N_4228,N_3384);
nor U7651 (N_7651,N_5912,N_4158);
nand U7652 (N_7652,N_3371,N_5162);
nand U7653 (N_7653,N_4082,N_5944);
or U7654 (N_7654,N_5238,N_5427);
nor U7655 (N_7655,N_4176,N_5548);
or U7656 (N_7656,N_5064,N_3481);
and U7657 (N_7657,N_5006,N_3662);
nand U7658 (N_7658,N_4687,N_3410);
nand U7659 (N_7659,N_4961,N_3701);
or U7660 (N_7660,N_4333,N_3598);
xor U7661 (N_7661,N_5599,N_5377);
xnor U7662 (N_7662,N_4902,N_3127);
and U7663 (N_7663,N_4077,N_4449);
or U7664 (N_7664,N_5385,N_3849);
xnor U7665 (N_7665,N_4891,N_4728);
xnor U7666 (N_7666,N_3835,N_5022);
nand U7667 (N_7667,N_4680,N_3916);
or U7668 (N_7668,N_3755,N_4089);
or U7669 (N_7669,N_3371,N_5315);
nand U7670 (N_7670,N_5854,N_4590);
xor U7671 (N_7671,N_4062,N_5676);
nand U7672 (N_7672,N_4149,N_5221);
or U7673 (N_7673,N_3154,N_5993);
nor U7674 (N_7674,N_4826,N_3186);
xnor U7675 (N_7675,N_4193,N_4801);
xnor U7676 (N_7676,N_5123,N_4112);
xnor U7677 (N_7677,N_4660,N_5685);
and U7678 (N_7678,N_4645,N_5920);
or U7679 (N_7679,N_4885,N_3675);
nor U7680 (N_7680,N_5668,N_3903);
nand U7681 (N_7681,N_4639,N_5322);
nand U7682 (N_7682,N_5954,N_3406);
and U7683 (N_7683,N_3541,N_3470);
and U7684 (N_7684,N_4795,N_3673);
or U7685 (N_7685,N_3637,N_5744);
xor U7686 (N_7686,N_4832,N_4766);
and U7687 (N_7687,N_5988,N_5501);
or U7688 (N_7688,N_5942,N_3744);
nor U7689 (N_7689,N_5491,N_4463);
and U7690 (N_7690,N_3069,N_3464);
nand U7691 (N_7691,N_5099,N_4568);
nand U7692 (N_7692,N_3098,N_4498);
nand U7693 (N_7693,N_5426,N_3956);
or U7694 (N_7694,N_4816,N_4494);
nand U7695 (N_7695,N_5876,N_4028);
and U7696 (N_7696,N_4336,N_4722);
nand U7697 (N_7697,N_4881,N_5462);
xnor U7698 (N_7698,N_5568,N_5970);
nor U7699 (N_7699,N_3578,N_3450);
and U7700 (N_7700,N_5858,N_3941);
or U7701 (N_7701,N_4472,N_5809);
and U7702 (N_7702,N_4030,N_5219);
and U7703 (N_7703,N_3032,N_4757);
nand U7704 (N_7704,N_3266,N_3753);
or U7705 (N_7705,N_3283,N_5449);
nor U7706 (N_7706,N_3846,N_3685);
xnor U7707 (N_7707,N_3393,N_3756);
and U7708 (N_7708,N_4198,N_4164);
or U7709 (N_7709,N_5309,N_3737);
nor U7710 (N_7710,N_3810,N_5102);
and U7711 (N_7711,N_3947,N_5295);
xor U7712 (N_7712,N_4297,N_5139);
and U7713 (N_7713,N_5636,N_4855);
or U7714 (N_7714,N_3037,N_3863);
or U7715 (N_7715,N_4021,N_3199);
and U7716 (N_7716,N_5370,N_5717);
nor U7717 (N_7717,N_3144,N_4421);
xor U7718 (N_7718,N_5810,N_3006);
nor U7719 (N_7719,N_4574,N_3015);
and U7720 (N_7720,N_5726,N_5706);
and U7721 (N_7721,N_5252,N_5607);
nand U7722 (N_7722,N_3240,N_5383);
or U7723 (N_7723,N_5528,N_4783);
and U7724 (N_7724,N_4907,N_3778);
nor U7725 (N_7725,N_4528,N_5564);
and U7726 (N_7726,N_5307,N_4149);
and U7727 (N_7727,N_4706,N_3752);
or U7728 (N_7728,N_3302,N_5693);
xnor U7729 (N_7729,N_5602,N_4122);
nor U7730 (N_7730,N_5717,N_3226);
nand U7731 (N_7731,N_4603,N_4534);
xnor U7732 (N_7732,N_5269,N_4952);
and U7733 (N_7733,N_5739,N_5777);
and U7734 (N_7734,N_5471,N_4143);
or U7735 (N_7735,N_5117,N_3874);
xnor U7736 (N_7736,N_4064,N_4812);
nor U7737 (N_7737,N_5504,N_5932);
and U7738 (N_7738,N_3031,N_4271);
and U7739 (N_7739,N_3118,N_3053);
xor U7740 (N_7740,N_5654,N_4956);
nor U7741 (N_7741,N_3079,N_4139);
xor U7742 (N_7742,N_4809,N_5867);
nor U7743 (N_7743,N_5113,N_5880);
or U7744 (N_7744,N_5025,N_3432);
xnor U7745 (N_7745,N_4137,N_3304);
xor U7746 (N_7746,N_5232,N_3896);
or U7747 (N_7747,N_5530,N_5420);
nand U7748 (N_7748,N_5132,N_4279);
xor U7749 (N_7749,N_4274,N_3837);
xor U7750 (N_7750,N_4197,N_3926);
and U7751 (N_7751,N_5926,N_5306);
nor U7752 (N_7752,N_4163,N_3804);
xor U7753 (N_7753,N_4033,N_3067);
nand U7754 (N_7754,N_3611,N_5760);
nand U7755 (N_7755,N_4785,N_5880);
nor U7756 (N_7756,N_4350,N_4253);
and U7757 (N_7757,N_4381,N_3633);
or U7758 (N_7758,N_5381,N_5093);
xor U7759 (N_7759,N_3130,N_3679);
and U7760 (N_7760,N_3960,N_4350);
xnor U7761 (N_7761,N_4633,N_3171);
xor U7762 (N_7762,N_4763,N_3788);
and U7763 (N_7763,N_5232,N_5349);
nand U7764 (N_7764,N_4034,N_5193);
or U7765 (N_7765,N_3006,N_3171);
nor U7766 (N_7766,N_4847,N_4225);
xor U7767 (N_7767,N_5087,N_3836);
or U7768 (N_7768,N_5357,N_5896);
nor U7769 (N_7769,N_3556,N_5574);
nor U7770 (N_7770,N_5641,N_4530);
or U7771 (N_7771,N_4182,N_5585);
nand U7772 (N_7772,N_3131,N_3711);
and U7773 (N_7773,N_3344,N_4178);
nor U7774 (N_7774,N_5048,N_4578);
nand U7775 (N_7775,N_5844,N_4150);
nand U7776 (N_7776,N_5769,N_5010);
nor U7777 (N_7777,N_5652,N_4355);
and U7778 (N_7778,N_3912,N_4269);
nand U7779 (N_7779,N_3739,N_4241);
nor U7780 (N_7780,N_3024,N_3816);
nand U7781 (N_7781,N_3653,N_5491);
or U7782 (N_7782,N_3112,N_5886);
xor U7783 (N_7783,N_5019,N_5293);
or U7784 (N_7784,N_3176,N_3817);
and U7785 (N_7785,N_4556,N_5940);
and U7786 (N_7786,N_5681,N_4490);
xnor U7787 (N_7787,N_4160,N_3301);
xnor U7788 (N_7788,N_4782,N_4323);
nor U7789 (N_7789,N_4376,N_4800);
or U7790 (N_7790,N_5582,N_4017);
nand U7791 (N_7791,N_3401,N_4353);
or U7792 (N_7792,N_3043,N_3270);
nor U7793 (N_7793,N_3181,N_5221);
nor U7794 (N_7794,N_4111,N_4166);
nor U7795 (N_7795,N_3960,N_5572);
nor U7796 (N_7796,N_5159,N_4166);
and U7797 (N_7797,N_3774,N_5131);
nand U7798 (N_7798,N_3863,N_4904);
nor U7799 (N_7799,N_4196,N_5094);
xor U7800 (N_7800,N_5902,N_4477);
nand U7801 (N_7801,N_5137,N_3395);
nor U7802 (N_7802,N_4728,N_3151);
xnor U7803 (N_7803,N_3932,N_5125);
nor U7804 (N_7804,N_4213,N_5053);
nor U7805 (N_7805,N_3714,N_4217);
nand U7806 (N_7806,N_4062,N_4757);
nand U7807 (N_7807,N_5269,N_5749);
or U7808 (N_7808,N_5725,N_4327);
or U7809 (N_7809,N_4173,N_4236);
nor U7810 (N_7810,N_3997,N_3670);
xnor U7811 (N_7811,N_4719,N_5989);
xor U7812 (N_7812,N_4017,N_5629);
xnor U7813 (N_7813,N_5450,N_5911);
and U7814 (N_7814,N_4947,N_3306);
and U7815 (N_7815,N_3378,N_5446);
or U7816 (N_7816,N_5453,N_4287);
nand U7817 (N_7817,N_4616,N_5805);
xnor U7818 (N_7818,N_3175,N_3561);
nand U7819 (N_7819,N_4575,N_3408);
or U7820 (N_7820,N_5045,N_4584);
and U7821 (N_7821,N_5344,N_5235);
xor U7822 (N_7822,N_4404,N_3869);
or U7823 (N_7823,N_3878,N_3309);
nand U7824 (N_7824,N_3285,N_4175);
nand U7825 (N_7825,N_5415,N_5335);
xor U7826 (N_7826,N_4119,N_4948);
and U7827 (N_7827,N_5397,N_4970);
nor U7828 (N_7828,N_5800,N_3854);
and U7829 (N_7829,N_3579,N_3849);
nor U7830 (N_7830,N_4311,N_5829);
nor U7831 (N_7831,N_5770,N_5854);
and U7832 (N_7832,N_5172,N_3332);
xnor U7833 (N_7833,N_3279,N_4264);
xor U7834 (N_7834,N_5444,N_3352);
xnor U7835 (N_7835,N_5069,N_5381);
nand U7836 (N_7836,N_4531,N_5928);
or U7837 (N_7837,N_4370,N_3864);
nand U7838 (N_7838,N_3740,N_4780);
nor U7839 (N_7839,N_3567,N_5871);
nand U7840 (N_7840,N_3958,N_4131);
nor U7841 (N_7841,N_4745,N_3585);
nand U7842 (N_7842,N_4442,N_3405);
nand U7843 (N_7843,N_3976,N_4816);
xnor U7844 (N_7844,N_5914,N_3640);
nor U7845 (N_7845,N_5647,N_3936);
xnor U7846 (N_7846,N_4601,N_5785);
xor U7847 (N_7847,N_3435,N_3347);
and U7848 (N_7848,N_3534,N_4764);
nand U7849 (N_7849,N_3595,N_5656);
nor U7850 (N_7850,N_4625,N_5557);
or U7851 (N_7851,N_4255,N_5387);
xnor U7852 (N_7852,N_4817,N_5247);
nor U7853 (N_7853,N_4396,N_3166);
nor U7854 (N_7854,N_4193,N_5167);
nand U7855 (N_7855,N_3714,N_3716);
xor U7856 (N_7856,N_3591,N_3887);
nor U7857 (N_7857,N_3593,N_3423);
and U7858 (N_7858,N_3706,N_3518);
nor U7859 (N_7859,N_3916,N_5494);
and U7860 (N_7860,N_5069,N_4538);
or U7861 (N_7861,N_4683,N_3849);
or U7862 (N_7862,N_4694,N_3838);
or U7863 (N_7863,N_5414,N_4845);
nor U7864 (N_7864,N_5568,N_4933);
nand U7865 (N_7865,N_5534,N_3161);
or U7866 (N_7866,N_4458,N_3285);
xor U7867 (N_7867,N_5921,N_5767);
and U7868 (N_7868,N_3133,N_3231);
and U7869 (N_7869,N_3948,N_5832);
or U7870 (N_7870,N_3211,N_4809);
nand U7871 (N_7871,N_4295,N_4509);
nor U7872 (N_7872,N_4602,N_4665);
nand U7873 (N_7873,N_5727,N_3297);
xor U7874 (N_7874,N_5061,N_5362);
xnor U7875 (N_7875,N_4724,N_5714);
nand U7876 (N_7876,N_5299,N_4770);
nor U7877 (N_7877,N_4906,N_4433);
xnor U7878 (N_7878,N_4437,N_3821);
nand U7879 (N_7879,N_4328,N_3955);
xnor U7880 (N_7880,N_4179,N_3439);
and U7881 (N_7881,N_3509,N_4899);
nand U7882 (N_7882,N_4617,N_5546);
nor U7883 (N_7883,N_5191,N_5636);
nor U7884 (N_7884,N_3830,N_3552);
xor U7885 (N_7885,N_4636,N_5724);
or U7886 (N_7886,N_5428,N_5209);
nand U7887 (N_7887,N_4554,N_3255);
xor U7888 (N_7888,N_4297,N_5776);
and U7889 (N_7889,N_5098,N_4309);
nor U7890 (N_7890,N_4121,N_5504);
nand U7891 (N_7891,N_3740,N_4412);
nand U7892 (N_7892,N_3234,N_5525);
nor U7893 (N_7893,N_4371,N_5369);
and U7894 (N_7894,N_5275,N_4423);
and U7895 (N_7895,N_4130,N_5357);
nand U7896 (N_7896,N_5019,N_4572);
xor U7897 (N_7897,N_3136,N_4315);
and U7898 (N_7898,N_5297,N_3529);
nand U7899 (N_7899,N_4864,N_5554);
and U7900 (N_7900,N_3833,N_5999);
or U7901 (N_7901,N_5667,N_5660);
nor U7902 (N_7902,N_4236,N_4794);
nor U7903 (N_7903,N_5395,N_5548);
or U7904 (N_7904,N_3871,N_4139);
and U7905 (N_7905,N_4160,N_4994);
or U7906 (N_7906,N_5410,N_5147);
nand U7907 (N_7907,N_5998,N_5405);
nor U7908 (N_7908,N_3252,N_4764);
or U7909 (N_7909,N_5388,N_5304);
xor U7910 (N_7910,N_5149,N_3720);
xor U7911 (N_7911,N_4183,N_3724);
nor U7912 (N_7912,N_3903,N_3706);
nor U7913 (N_7913,N_5899,N_3158);
nor U7914 (N_7914,N_3912,N_4440);
and U7915 (N_7915,N_3305,N_5909);
or U7916 (N_7916,N_5680,N_3420);
nand U7917 (N_7917,N_5968,N_3950);
or U7918 (N_7918,N_3198,N_3390);
and U7919 (N_7919,N_4192,N_5417);
nand U7920 (N_7920,N_4716,N_4595);
or U7921 (N_7921,N_3216,N_3591);
nand U7922 (N_7922,N_3393,N_5029);
nand U7923 (N_7923,N_5516,N_5577);
nor U7924 (N_7924,N_5874,N_3907);
nor U7925 (N_7925,N_5010,N_4748);
nand U7926 (N_7926,N_4928,N_3169);
or U7927 (N_7927,N_4956,N_5768);
nor U7928 (N_7928,N_5505,N_5222);
nor U7929 (N_7929,N_5017,N_3182);
or U7930 (N_7930,N_3774,N_4206);
and U7931 (N_7931,N_4251,N_4619);
nor U7932 (N_7932,N_5666,N_5814);
nor U7933 (N_7933,N_4448,N_3457);
and U7934 (N_7934,N_5790,N_3635);
nand U7935 (N_7935,N_5945,N_4143);
and U7936 (N_7936,N_3091,N_5965);
nor U7937 (N_7937,N_4204,N_5459);
and U7938 (N_7938,N_5239,N_4413);
and U7939 (N_7939,N_3971,N_4201);
or U7940 (N_7940,N_5814,N_5538);
and U7941 (N_7941,N_3639,N_3679);
nand U7942 (N_7942,N_3606,N_4664);
and U7943 (N_7943,N_4862,N_4373);
nand U7944 (N_7944,N_5208,N_4217);
xor U7945 (N_7945,N_3744,N_3821);
or U7946 (N_7946,N_5831,N_3611);
or U7947 (N_7947,N_3748,N_3830);
and U7948 (N_7948,N_4799,N_5650);
nand U7949 (N_7949,N_5622,N_3115);
and U7950 (N_7950,N_3109,N_4292);
nor U7951 (N_7951,N_3305,N_5102);
and U7952 (N_7952,N_4400,N_5576);
nand U7953 (N_7953,N_4099,N_3342);
and U7954 (N_7954,N_4741,N_3873);
or U7955 (N_7955,N_4803,N_3796);
or U7956 (N_7956,N_4847,N_3100);
nor U7957 (N_7957,N_4353,N_5385);
nand U7958 (N_7958,N_3109,N_3539);
nand U7959 (N_7959,N_3366,N_5102);
xnor U7960 (N_7960,N_4413,N_4579);
nor U7961 (N_7961,N_4244,N_4907);
nor U7962 (N_7962,N_5667,N_3686);
xor U7963 (N_7963,N_5082,N_5935);
or U7964 (N_7964,N_3330,N_3402);
or U7965 (N_7965,N_4979,N_5132);
nor U7966 (N_7966,N_5266,N_3686);
or U7967 (N_7967,N_3867,N_5942);
or U7968 (N_7968,N_3439,N_3323);
and U7969 (N_7969,N_3214,N_5058);
nor U7970 (N_7970,N_3245,N_5817);
nand U7971 (N_7971,N_3199,N_4104);
and U7972 (N_7972,N_5236,N_4126);
nand U7973 (N_7973,N_4218,N_5629);
nor U7974 (N_7974,N_5315,N_5990);
and U7975 (N_7975,N_5846,N_5635);
nor U7976 (N_7976,N_5494,N_4699);
nand U7977 (N_7977,N_3881,N_3196);
and U7978 (N_7978,N_3710,N_3401);
nand U7979 (N_7979,N_4096,N_4568);
nand U7980 (N_7980,N_3000,N_4970);
xor U7981 (N_7981,N_3979,N_5569);
or U7982 (N_7982,N_4926,N_3984);
and U7983 (N_7983,N_4201,N_4499);
or U7984 (N_7984,N_3332,N_5188);
nand U7985 (N_7985,N_4409,N_4813);
and U7986 (N_7986,N_4165,N_5509);
nand U7987 (N_7987,N_5120,N_5242);
or U7988 (N_7988,N_4521,N_4627);
xnor U7989 (N_7989,N_3861,N_5642);
or U7990 (N_7990,N_5135,N_3521);
and U7991 (N_7991,N_3130,N_5387);
nand U7992 (N_7992,N_4898,N_4516);
xor U7993 (N_7993,N_3126,N_3979);
or U7994 (N_7994,N_4355,N_3258);
and U7995 (N_7995,N_4289,N_4801);
or U7996 (N_7996,N_3274,N_3595);
nand U7997 (N_7997,N_3323,N_5610);
xnor U7998 (N_7998,N_3401,N_3258);
xor U7999 (N_7999,N_3625,N_4479);
xnor U8000 (N_8000,N_4522,N_4219);
and U8001 (N_8001,N_4173,N_5370);
and U8002 (N_8002,N_4767,N_3343);
nor U8003 (N_8003,N_4972,N_4765);
nand U8004 (N_8004,N_4585,N_3289);
and U8005 (N_8005,N_4813,N_4898);
xor U8006 (N_8006,N_4401,N_4311);
nand U8007 (N_8007,N_4893,N_4580);
and U8008 (N_8008,N_4795,N_4457);
xor U8009 (N_8009,N_3189,N_3761);
nor U8010 (N_8010,N_3171,N_4971);
xnor U8011 (N_8011,N_5040,N_3369);
or U8012 (N_8012,N_4740,N_3060);
and U8013 (N_8013,N_5654,N_3525);
nand U8014 (N_8014,N_5680,N_5040);
nor U8015 (N_8015,N_3089,N_5591);
and U8016 (N_8016,N_3913,N_3520);
nand U8017 (N_8017,N_3701,N_4523);
nor U8018 (N_8018,N_5398,N_5774);
nor U8019 (N_8019,N_5654,N_3374);
nand U8020 (N_8020,N_4520,N_4456);
nand U8021 (N_8021,N_5198,N_5975);
xor U8022 (N_8022,N_3770,N_4368);
nor U8023 (N_8023,N_4127,N_5060);
xor U8024 (N_8024,N_4519,N_3868);
nor U8025 (N_8025,N_4433,N_3709);
nand U8026 (N_8026,N_4883,N_3225);
xor U8027 (N_8027,N_3771,N_3769);
nor U8028 (N_8028,N_5195,N_4820);
nand U8029 (N_8029,N_5733,N_3686);
and U8030 (N_8030,N_4810,N_4054);
xnor U8031 (N_8031,N_5635,N_3753);
or U8032 (N_8032,N_5322,N_4170);
nand U8033 (N_8033,N_3902,N_4455);
or U8034 (N_8034,N_3141,N_3064);
nand U8035 (N_8035,N_5066,N_4356);
or U8036 (N_8036,N_3783,N_4188);
or U8037 (N_8037,N_5484,N_5696);
or U8038 (N_8038,N_5942,N_4704);
nand U8039 (N_8039,N_4703,N_3697);
xnor U8040 (N_8040,N_3526,N_4595);
nand U8041 (N_8041,N_5619,N_3178);
and U8042 (N_8042,N_3706,N_5403);
nand U8043 (N_8043,N_3583,N_3723);
and U8044 (N_8044,N_4681,N_4824);
nor U8045 (N_8045,N_3908,N_5800);
nor U8046 (N_8046,N_5933,N_3814);
or U8047 (N_8047,N_3207,N_4032);
xnor U8048 (N_8048,N_3737,N_5911);
or U8049 (N_8049,N_5704,N_4458);
nand U8050 (N_8050,N_3131,N_4002);
nand U8051 (N_8051,N_4453,N_5476);
or U8052 (N_8052,N_5733,N_4226);
xor U8053 (N_8053,N_4221,N_5546);
and U8054 (N_8054,N_3645,N_4427);
and U8055 (N_8055,N_3492,N_3215);
xor U8056 (N_8056,N_5018,N_3283);
and U8057 (N_8057,N_3775,N_4785);
and U8058 (N_8058,N_3374,N_5389);
nand U8059 (N_8059,N_4470,N_4497);
or U8060 (N_8060,N_5280,N_3511);
or U8061 (N_8061,N_3117,N_4025);
xnor U8062 (N_8062,N_4619,N_3830);
nor U8063 (N_8063,N_3564,N_5894);
nand U8064 (N_8064,N_5189,N_3948);
nand U8065 (N_8065,N_4461,N_5995);
xor U8066 (N_8066,N_3268,N_4709);
or U8067 (N_8067,N_5376,N_4891);
or U8068 (N_8068,N_5146,N_3529);
and U8069 (N_8069,N_3776,N_4138);
nand U8070 (N_8070,N_5884,N_5372);
or U8071 (N_8071,N_4717,N_5479);
or U8072 (N_8072,N_3384,N_4087);
nand U8073 (N_8073,N_3540,N_3665);
nand U8074 (N_8074,N_3098,N_4993);
nand U8075 (N_8075,N_4790,N_3288);
xor U8076 (N_8076,N_3906,N_4829);
nor U8077 (N_8077,N_5042,N_3179);
nand U8078 (N_8078,N_5923,N_5535);
or U8079 (N_8079,N_3433,N_4124);
nand U8080 (N_8080,N_4836,N_5903);
xor U8081 (N_8081,N_5446,N_4331);
and U8082 (N_8082,N_4432,N_4002);
and U8083 (N_8083,N_4568,N_4169);
nor U8084 (N_8084,N_3190,N_3067);
xnor U8085 (N_8085,N_3865,N_3217);
and U8086 (N_8086,N_5554,N_3367);
xor U8087 (N_8087,N_3979,N_4752);
nor U8088 (N_8088,N_5264,N_4315);
nand U8089 (N_8089,N_3688,N_5679);
or U8090 (N_8090,N_3381,N_3617);
nand U8091 (N_8091,N_5202,N_3727);
xnor U8092 (N_8092,N_5670,N_4466);
and U8093 (N_8093,N_5503,N_3530);
and U8094 (N_8094,N_4743,N_5149);
and U8095 (N_8095,N_3865,N_3195);
xor U8096 (N_8096,N_5292,N_4148);
xor U8097 (N_8097,N_5979,N_3028);
xnor U8098 (N_8098,N_4586,N_4875);
nand U8099 (N_8099,N_5700,N_4141);
xor U8100 (N_8100,N_5739,N_4472);
nor U8101 (N_8101,N_3474,N_5255);
xnor U8102 (N_8102,N_3721,N_5121);
and U8103 (N_8103,N_5288,N_5364);
nor U8104 (N_8104,N_5739,N_3293);
nor U8105 (N_8105,N_5648,N_4983);
nand U8106 (N_8106,N_4098,N_4730);
xor U8107 (N_8107,N_3700,N_4695);
nor U8108 (N_8108,N_5307,N_5702);
and U8109 (N_8109,N_4246,N_4576);
nor U8110 (N_8110,N_3646,N_3644);
or U8111 (N_8111,N_4225,N_3714);
or U8112 (N_8112,N_4849,N_4653);
xor U8113 (N_8113,N_3099,N_5471);
xnor U8114 (N_8114,N_5313,N_5056);
or U8115 (N_8115,N_3627,N_4169);
nand U8116 (N_8116,N_5899,N_4924);
and U8117 (N_8117,N_3518,N_5349);
xnor U8118 (N_8118,N_5183,N_4997);
nor U8119 (N_8119,N_3469,N_4441);
nand U8120 (N_8120,N_4448,N_5213);
and U8121 (N_8121,N_4864,N_5519);
nand U8122 (N_8122,N_3010,N_3083);
nand U8123 (N_8123,N_5810,N_4477);
nor U8124 (N_8124,N_4637,N_5971);
nor U8125 (N_8125,N_5340,N_5766);
and U8126 (N_8126,N_3158,N_3073);
and U8127 (N_8127,N_4029,N_4800);
and U8128 (N_8128,N_3085,N_5683);
nor U8129 (N_8129,N_4662,N_4359);
or U8130 (N_8130,N_3600,N_4547);
nor U8131 (N_8131,N_4248,N_5045);
or U8132 (N_8132,N_4305,N_3059);
nor U8133 (N_8133,N_3552,N_5024);
nand U8134 (N_8134,N_5055,N_3823);
and U8135 (N_8135,N_4540,N_3422);
and U8136 (N_8136,N_3226,N_4582);
xor U8137 (N_8137,N_4333,N_4652);
xor U8138 (N_8138,N_5456,N_3951);
xnor U8139 (N_8139,N_5646,N_4134);
and U8140 (N_8140,N_5779,N_3497);
or U8141 (N_8141,N_4848,N_5411);
xor U8142 (N_8142,N_5192,N_3410);
and U8143 (N_8143,N_4792,N_4743);
or U8144 (N_8144,N_4849,N_5028);
xor U8145 (N_8145,N_4421,N_4979);
nand U8146 (N_8146,N_5379,N_3814);
nor U8147 (N_8147,N_3104,N_3588);
nand U8148 (N_8148,N_4795,N_5133);
and U8149 (N_8149,N_4613,N_4636);
nand U8150 (N_8150,N_5056,N_4810);
and U8151 (N_8151,N_4284,N_3793);
xnor U8152 (N_8152,N_3565,N_4497);
or U8153 (N_8153,N_4723,N_5359);
and U8154 (N_8154,N_5789,N_3893);
xor U8155 (N_8155,N_3375,N_4066);
or U8156 (N_8156,N_4902,N_3337);
nor U8157 (N_8157,N_3713,N_4073);
nand U8158 (N_8158,N_3373,N_5523);
nand U8159 (N_8159,N_5648,N_4564);
nor U8160 (N_8160,N_5059,N_4266);
xor U8161 (N_8161,N_4065,N_5337);
nand U8162 (N_8162,N_4790,N_4133);
nor U8163 (N_8163,N_5636,N_3719);
xor U8164 (N_8164,N_4860,N_3740);
xor U8165 (N_8165,N_3289,N_3769);
xor U8166 (N_8166,N_3321,N_3963);
or U8167 (N_8167,N_4229,N_4081);
and U8168 (N_8168,N_5365,N_4862);
nand U8169 (N_8169,N_4187,N_3200);
nor U8170 (N_8170,N_3537,N_3964);
and U8171 (N_8171,N_3714,N_4092);
nand U8172 (N_8172,N_3625,N_5946);
nand U8173 (N_8173,N_5483,N_3570);
xnor U8174 (N_8174,N_4175,N_5156);
and U8175 (N_8175,N_5645,N_5665);
nor U8176 (N_8176,N_5480,N_5256);
xnor U8177 (N_8177,N_5892,N_5195);
nor U8178 (N_8178,N_4507,N_3206);
or U8179 (N_8179,N_3497,N_4069);
or U8180 (N_8180,N_5297,N_4633);
nor U8181 (N_8181,N_5432,N_3875);
nor U8182 (N_8182,N_3240,N_3241);
xnor U8183 (N_8183,N_4369,N_5626);
nand U8184 (N_8184,N_5942,N_4765);
nand U8185 (N_8185,N_4302,N_3707);
nor U8186 (N_8186,N_4276,N_5927);
nand U8187 (N_8187,N_3294,N_3724);
nand U8188 (N_8188,N_5051,N_4732);
xor U8189 (N_8189,N_5312,N_3317);
nand U8190 (N_8190,N_3353,N_3298);
nand U8191 (N_8191,N_5213,N_4396);
or U8192 (N_8192,N_3506,N_4330);
nand U8193 (N_8193,N_3319,N_4070);
or U8194 (N_8194,N_5360,N_4899);
and U8195 (N_8195,N_4040,N_5768);
nand U8196 (N_8196,N_3672,N_3011);
and U8197 (N_8197,N_3281,N_3327);
or U8198 (N_8198,N_4755,N_3348);
nor U8199 (N_8199,N_3246,N_4325);
xnor U8200 (N_8200,N_4174,N_5979);
xor U8201 (N_8201,N_5129,N_4914);
xor U8202 (N_8202,N_3538,N_5588);
xnor U8203 (N_8203,N_5175,N_4175);
nor U8204 (N_8204,N_3970,N_4541);
nor U8205 (N_8205,N_3104,N_5090);
nor U8206 (N_8206,N_4149,N_5691);
nand U8207 (N_8207,N_5946,N_3164);
and U8208 (N_8208,N_4335,N_3427);
nor U8209 (N_8209,N_4563,N_3447);
nor U8210 (N_8210,N_5911,N_4354);
xnor U8211 (N_8211,N_4651,N_5050);
or U8212 (N_8212,N_4236,N_4701);
xor U8213 (N_8213,N_3436,N_3361);
nand U8214 (N_8214,N_5401,N_3729);
nand U8215 (N_8215,N_5621,N_4782);
xor U8216 (N_8216,N_3196,N_3900);
nand U8217 (N_8217,N_3524,N_5796);
xor U8218 (N_8218,N_3256,N_4871);
and U8219 (N_8219,N_4670,N_4132);
xnor U8220 (N_8220,N_4763,N_4297);
or U8221 (N_8221,N_3650,N_5049);
nand U8222 (N_8222,N_4204,N_4255);
or U8223 (N_8223,N_3472,N_5234);
nand U8224 (N_8224,N_3565,N_3204);
xnor U8225 (N_8225,N_4018,N_3135);
nor U8226 (N_8226,N_3052,N_4374);
and U8227 (N_8227,N_5318,N_3200);
and U8228 (N_8228,N_4255,N_4500);
or U8229 (N_8229,N_5112,N_5533);
xor U8230 (N_8230,N_5646,N_5054);
and U8231 (N_8231,N_5573,N_3009);
xnor U8232 (N_8232,N_4834,N_3256);
nand U8233 (N_8233,N_4913,N_5705);
nor U8234 (N_8234,N_5476,N_3103);
and U8235 (N_8235,N_4375,N_3464);
and U8236 (N_8236,N_5497,N_4875);
or U8237 (N_8237,N_5565,N_4172);
or U8238 (N_8238,N_3253,N_3349);
xor U8239 (N_8239,N_3347,N_4612);
nor U8240 (N_8240,N_4828,N_3032);
nor U8241 (N_8241,N_3101,N_3666);
nor U8242 (N_8242,N_3855,N_5094);
or U8243 (N_8243,N_5996,N_3254);
and U8244 (N_8244,N_5294,N_3398);
and U8245 (N_8245,N_4809,N_5434);
and U8246 (N_8246,N_4666,N_4345);
and U8247 (N_8247,N_4615,N_3013);
xor U8248 (N_8248,N_4814,N_3612);
nand U8249 (N_8249,N_5725,N_5435);
or U8250 (N_8250,N_3220,N_5149);
and U8251 (N_8251,N_3980,N_4714);
nor U8252 (N_8252,N_4020,N_4713);
nor U8253 (N_8253,N_3239,N_4097);
and U8254 (N_8254,N_5204,N_5851);
xor U8255 (N_8255,N_4817,N_3021);
or U8256 (N_8256,N_5687,N_3060);
and U8257 (N_8257,N_4830,N_5619);
nor U8258 (N_8258,N_4472,N_3609);
and U8259 (N_8259,N_3136,N_3424);
and U8260 (N_8260,N_4155,N_5798);
or U8261 (N_8261,N_5548,N_3391);
or U8262 (N_8262,N_5363,N_5152);
xor U8263 (N_8263,N_5544,N_3656);
xor U8264 (N_8264,N_5150,N_5034);
and U8265 (N_8265,N_4466,N_5876);
xor U8266 (N_8266,N_4962,N_3134);
xnor U8267 (N_8267,N_5052,N_4029);
nand U8268 (N_8268,N_4543,N_4050);
and U8269 (N_8269,N_3013,N_3920);
and U8270 (N_8270,N_5749,N_5904);
xor U8271 (N_8271,N_5998,N_5205);
xor U8272 (N_8272,N_4937,N_5353);
and U8273 (N_8273,N_5060,N_4997);
xor U8274 (N_8274,N_4823,N_3738);
or U8275 (N_8275,N_5068,N_4510);
nor U8276 (N_8276,N_5808,N_4783);
nor U8277 (N_8277,N_4605,N_5727);
xnor U8278 (N_8278,N_5725,N_5690);
and U8279 (N_8279,N_3844,N_4711);
or U8280 (N_8280,N_4184,N_3907);
or U8281 (N_8281,N_4781,N_4153);
and U8282 (N_8282,N_4027,N_5836);
nor U8283 (N_8283,N_5726,N_3342);
and U8284 (N_8284,N_5910,N_4208);
or U8285 (N_8285,N_3508,N_5159);
or U8286 (N_8286,N_4723,N_4351);
xor U8287 (N_8287,N_3283,N_3083);
xnor U8288 (N_8288,N_3699,N_5132);
nand U8289 (N_8289,N_5315,N_3847);
and U8290 (N_8290,N_3611,N_4869);
or U8291 (N_8291,N_4466,N_5930);
xor U8292 (N_8292,N_4005,N_3147);
or U8293 (N_8293,N_5206,N_5462);
and U8294 (N_8294,N_5773,N_3876);
xnor U8295 (N_8295,N_5755,N_5101);
nor U8296 (N_8296,N_3638,N_5004);
or U8297 (N_8297,N_4399,N_4837);
or U8298 (N_8298,N_5969,N_5941);
nor U8299 (N_8299,N_5546,N_5760);
nand U8300 (N_8300,N_4442,N_4231);
nand U8301 (N_8301,N_5172,N_3135);
or U8302 (N_8302,N_4401,N_4594);
nand U8303 (N_8303,N_5939,N_3930);
xnor U8304 (N_8304,N_5429,N_4767);
nor U8305 (N_8305,N_5941,N_3957);
and U8306 (N_8306,N_4012,N_4028);
or U8307 (N_8307,N_3733,N_4485);
or U8308 (N_8308,N_3292,N_5811);
nand U8309 (N_8309,N_3077,N_5559);
xnor U8310 (N_8310,N_3950,N_5746);
nand U8311 (N_8311,N_4156,N_5311);
or U8312 (N_8312,N_4274,N_4198);
or U8313 (N_8313,N_4797,N_3558);
xor U8314 (N_8314,N_5237,N_3493);
or U8315 (N_8315,N_3351,N_5884);
and U8316 (N_8316,N_3818,N_4242);
xor U8317 (N_8317,N_3135,N_4561);
xor U8318 (N_8318,N_3706,N_5606);
or U8319 (N_8319,N_4700,N_5376);
or U8320 (N_8320,N_4184,N_3398);
xnor U8321 (N_8321,N_3827,N_4635);
or U8322 (N_8322,N_5589,N_4340);
and U8323 (N_8323,N_3687,N_5523);
nor U8324 (N_8324,N_4023,N_5997);
xor U8325 (N_8325,N_5909,N_3733);
xnor U8326 (N_8326,N_4610,N_5609);
xor U8327 (N_8327,N_3315,N_4892);
xnor U8328 (N_8328,N_4813,N_4926);
xnor U8329 (N_8329,N_3679,N_5429);
and U8330 (N_8330,N_3063,N_4289);
or U8331 (N_8331,N_5669,N_5446);
xnor U8332 (N_8332,N_3777,N_4251);
and U8333 (N_8333,N_5058,N_5770);
or U8334 (N_8334,N_5212,N_3874);
or U8335 (N_8335,N_5163,N_3436);
or U8336 (N_8336,N_3376,N_3927);
nor U8337 (N_8337,N_3093,N_4519);
nor U8338 (N_8338,N_3015,N_5688);
or U8339 (N_8339,N_4011,N_5589);
and U8340 (N_8340,N_4403,N_5951);
xnor U8341 (N_8341,N_4714,N_3187);
or U8342 (N_8342,N_5308,N_5369);
and U8343 (N_8343,N_4044,N_4697);
nor U8344 (N_8344,N_3485,N_5487);
and U8345 (N_8345,N_4662,N_3991);
and U8346 (N_8346,N_5286,N_4059);
nand U8347 (N_8347,N_3346,N_3567);
or U8348 (N_8348,N_4921,N_3487);
nand U8349 (N_8349,N_4395,N_3965);
and U8350 (N_8350,N_4339,N_3744);
or U8351 (N_8351,N_5514,N_5289);
or U8352 (N_8352,N_3229,N_3732);
or U8353 (N_8353,N_3388,N_3897);
and U8354 (N_8354,N_3515,N_3193);
or U8355 (N_8355,N_3631,N_4617);
and U8356 (N_8356,N_3036,N_3709);
nor U8357 (N_8357,N_3856,N_4593);
or U8358 (N_8358,N_4143,N_5620);
xor U8359 (N_8359,N_5213,N_4197);
xnor U8360 (N_8360,N_4707,N_5357);
xor U8361 (N_8361,N_3550,N_5417);
xnor U8362 (N_8362,N_4636,N_4842);
xnor U8363 (N_8363,N_3394,N_5916);
nand U8364 (N_8364,N_3752,N_4345);
nor U8365 (N_8365,N_4622,N_4855);
or U8366 (N_8366,N_5427,N_4904);
xnor U8367 (N_8367,N_5939,N_3988);
nand U8368 (N_8368,N_4176,N_4516);
nand U8369 (N_8369,N_5994,N_4982);
xnor U8370 (N_8370,N_4334,N_4490);
nor U8371 (N_8371,N_4028,N_4989);
nand U8372 (N_8372,N_3530,N_4388);
xor U8373 (N_8373,N_4505,N_4088);
and U8374 (N_8374,N_5831,N_3044);
or U8375 (N_8375,N_4859,N_3455);
and U8376 (N_8376,N_4096,N_3389);
and U8377 (N_8377,N_4259,N_5449);
and U8378 (N_8378,N_3284,N_3879);
or U8379 (N_8379,N_5203,N_5751);
or U8380 (N_8380,N_4078,N_5716);
or U8381 (N_8381,N_3500,N_4995);
and U8382 (N_8382,N_3288,N_3907);
nor U8383 (N_8383,N_4351,N_4076);
and U8384 (N_8384,N_3041,N_4242);
nor U8385 (N_8385,N_4272,N_4192);
or U8386 (N_8386,N_3759,N_3555);
xnor U8387 (N_8387,N_4648,N_5714);
nand U8388 (N_8388,N_5555,N_3354);
xor U8389 (N_8389,N_5445,N_3577);
xor U8390 (N_8390,N_4642,N_4169);
xor U8391 (N_8391,N_5019,N_5823);
and U8392 (N_8392,N_5455,N_4334);
or U8393 (N_8393,N_5728,N_5784);
xor U8394 (N_8394,N_5871,N_5732);
and U8395 (N_8395,N_4809,N_4069);
xor U8396 (N_8396,N_5212,N_3513);
or U8397 (N_8397,N_5681,N_3361);
xor U8398 (N_8398,N_4657,N_4655);
xnor U8399 (N_8399,N_3975,N_5446);
nor U8400 (N_8400,N_5303,N_4056);
or U8401 (N_8401,N_3370,N_4183);
nand U8402 (N_8402,N_4260,N_5405);
or U8403 (N_8403,N_4489,N_3593);
or U8404 (N_8404,N_5714,N_3041);
nor U8405 (N_8405,N_3331,N_5096);
xnor U8406 (N_8406,N_4379,N_3327);
nand U8407 (N_8407,N_3182,N_5756);
or U8408 (N_8408,N_3336,N_4429);
and U8409 (N_8409,N_4516,N_4957);
or U8410 (N_8410,N_4314,N_5181);
or U8411 (N_8411,N_4057,N_5327);
or U8412 (N_8412,N_3174,N_3332);
and U8413 (N_8413,N_5577,N_3798);
nor U8414 (N_8414,N_5451,N_5948);
xor U8415 (N_8415,N_5157,N_5318);
nand U8416 (N_8416,N_4734,N_4867);
nand U8417 (N_8417,N_3997,N_4988);
nor U8418 (N_8418,N_5172,N_5490);
nand U8419 (N_8419,N_3540,N_3128);
xor U8420 (N_8420,N_5511,N_4958);
nand U8421 (N_8421,N_3814,N_3433);
nor U8422 (N_8422,N_5574,N_5056);
xnor U8423 (N_8423,N_5696,N_4172);
xnor U8424 (N_8424,N_5980,N_4361);
nor U8425 (N_8425,N_4186,N_3128);
or U8426 (N_8426,N_4362,N_5057);
and U8427 (N_8427,N_5451,N_4665);
nor U8428 (N_8428,N_4751,N_3556);
or U8429 (N_8429,N_3283,N_5380);
nand U8430 (N_8430,N_4184,N_3262);
and U8431 (N_8431,N_5184,N_3863);
xnor U8432 (N_8432,N_5983,N_4980);
xnor U8433 (N_8433,N_3964,N_3803);
or U8434 (N_8434,N_4233,N_3434);
or U8435 (N_8435,N_5328,N_5888);
or U8436 (N_8436,N_3946,N_4837);
nand U8437 (N_8437,N_4308,N_5484);
nor U8438 (N_8438,N_3210,N_3991);
and U8439 (N_8439,N_3809,N_4606);
nor U8440 (N_8440,N_4579,N_3441);
and U8441 (N_8441,N_5362,N_3597);
xnor U8442 (N_8442,N_5657,N_3173);
or U8443 (N_8443,N_4638,N_4518);
and U8444 (N_8444,N_3136,N_5356);
or U8445 (N_8445,N_5125,N_4396);
nand U8446 (N_8446,N_3398,N_3577);
xor U8447 (N_8447,N_5288,N_4689);
and U8448 (N_8448,N_5320,N_4044);
nor U8449 (N_8449,N_3369,N_3004);
xnor U8450 (N_8450,N_3627,N_5192);
and U8451 (N_8451,N_4911,N_4926);
xnor U8452 (N_8452,N_4638,N_5092);
nand U8453 (N_8453,N_5448,N_3228);
nand U8454 (N_8454,N_4601,N_5475);
xor U8455 (N_8455,N_4219,N_3699);
nand U8456 (N_8456,N_3107,N_5591);
or U8457 (N_8457,N_3619,N_5373);
or U8458 (N_8458,N_5995,N_3648);
nor U8459 (N_8459,N_3388,N_4213);
xnor U8460 (N_8460,N_4637,N_4452);
and U8461 (N_8461,N_4238,N_4936);
or U8462 (N_8462,N_5557,N_5925);
and U8463 (N_8463,N_5515,N_5282);
nand U8464 (N_8464,N_5258,N_5390);
nand U8465 (N_8465,N_5805,N_3063);
or U8466 (N_8466,N_4711,N_3938);
xor U8467 (N_8467,N_4507,N_5128);
or U8468 (N_8468,N_3552,N_3204);
xor U8469 (N_8469,N_5515,N_4487);
nor U8470 (N_8470,N_3960,N_5351);
nand U8471 (N_8471,N_4557,N_5205);
nand U8472 (N_8472,N_3183,N_5948);
xor U8473 (N_8473,N_3090,N_5009);
and U8474 (N_8474,N_3862,N_4071);
and U8475 (N_8475,N_3347,N_3520);
or U8476 (N_8476,N_3928,N_5081);
nor U8477 (N_8477,N_4835,N_3882);
nor U8478 (N_8478,N_4596,N_5887);
or U8479 (N_8479,N_4620,N_3233);
nand U8480 (N_8480,N_4553,N_4934);
nor U8481 (N_8481,N_3888,N_4008);
nor U8482 (N_8482,N_4972,N_3450);
or U8483 (N_8483,N_5681,N_4504);
or U8484 (N_8484,N_3101,N_5617);
nand U8485 (N_8485,N_4871,N_4722);
nand U8486 (N_8486,N_5763,N_4049);
or U8487 (N_8487,N_4591,N_4788);
xor U8488 (N_8488,N_3332,N_3239);
xnor U8489 (N_8489,N_4446,N_4245);
xor U8490 (N_8490,N_5150,N_4142);
nand U8491 (N_8491,N_3549,N_5063);
nor U8492 (N_8492,N_5685,N_3861);
nand U8493 (N_8493,N_3016,N_5794);
nand U8494 (N_8494,N_5559,N_4566);
xnor U8495 (N_8495,N_5444,N_5662);
nor U8496 (N_8496,N_4715,N_3774);
nor U8497 (N_8497,N_5968,N_3539);
nand U8498 (N_8498,N_5475,N_5547);
nand U8499 (N_8499,N_3766,N_3687);
xnor U8500 (N_8500,N_3465,N_4662);
or U8501 (N_8501,N_4521,N_4454);
nand U8502 (N_8502,N_3321,N_5576);
or U8503 (N_8503,N_3953,N_5309);
nand U8504 (N_8504,N_5078,N_3863);
nand U8505 (N_8505,N_5149,N_3863);
nand U8506 (N_8506,N_5637,N_3130);
or U8507 (N_8507,N_5780,N_4113);
nor U8508 (N_8508,N_4500,N_4873);
nand U8509 (N_8509,N_4758,N_5213);
xor U8510 (N_8510,N_4390,N_4538);
or U8511 (N_8511,N_3735,N_3318);
or U8512 (N_8512,N_4942,N_4484);
and U8513 (N_8513,N_5947,N_4611);
xnor U8514 (N_8514,N_3665,N_4004);
or U8515 (N_8515,N_4008,N_4878);
or U8516 (N_8516,N_5126,N_4071);
xor U8517 (N_8517,N_4481,N_3118);
nor U8518 (N_8518,N_5532,N_5161);
and U8519 (N_8519,N_4970,N_5056);
and U8520 (N_8520,N_3004,N_4719);
or U8521 (N_8521,N_5151,N_4032);
xor U8522 (N_8522,N_4338,N_3917);
and U8523 (N_8523,N_5497,N_5463);
and U8524 (N_8524,N_3492,N_4568);
nor U8525 (N_8525,N_3672,N_3611);
and U8526 (N_8526,N_5787,N_4853);
or U8527 (N_8527,N_4901,N_4246);
nor U8528 (N_8528,N_4601,N_3009);
xnor U8529 (N_8529,N_3821,N_5477);
xor U8530 (N_8530,N_5345,N_4592);
and U8531 (N_8531,N_4517,N_5481);
or U8532 (N_8532,N_4822,N_4044);
nand U8533 (N_8533,N_5659,N_3587);
nand U8534 (N_8534,N_5249,N_4717);
nor U8535 (N_8535,N_5853,N_5534);
nor U8536 (N_8536,N_5006,N_4170);
and U8537 (N_8537,N_4820,N_5192);
or U8538 (N_8538,N_5665,N_3861);
xnor U8539 (N_8539,N_3770,N_5426);
or U8540 (N_8540,N_5477,N_5580);
nand U8541 (N_8541,N_4422,N_4314);
and U8542 (N_8542,N_4169,N_3596);
nand U8543 (N_8543,N_3456,N_4862);
xnor U8544 (N_8544,N_5814,N_4640);
nor U8545 (N_8545,N_5271,N_4439);
xnor U8546 (N_8546,N_5028,N_3222);
nand U8547 (N_8547,N_4005,N_3182);
and U8548 (N_8548,N_3965,N_3422);
or U8549 (N_8549,N_5178,N_4223);
nand U8550 (N_8550,N_3843,N_3106);
or U8551 (N_8551,N_3948,N_5089);
nor U8552 (N_8552,N_4810,N_3753);
or U8553 (N_8553,N_4431,N_3147);
nand U8554 (N_8554,N_5752,N_4797);
or U8555 (N_8555,N_4603,N_5322);
and U8556 (N_8556,N_3106,N_3874);
nand U8557 (N_8557,N_3297,N_3674);
xor U8558 (N_8558,N_4467,N_5886);
nand U8559 (N_8559,N_4709,N_5580);
nand U8560 (N_8560,N_4750,N_4625);
nand U8561 (N_8561,N_5139,N_5717);
xnor U8562 (N_8562,N_4527,N_5179);
xnor U8563 (N_8563,N_5142,N_4013);
nand U8564 (N_8564,N_5766,N_4295);
and U8565 (N_8565,N_3217,N_5193);
xor U8566 (N_8566,N_3505,N_4715);
nor U8567 (N_8567,N_4690,N_3967);
nor U8568 (N_8568,N_3949,N_3531);
nand U8569 (N_8569,N_5427,N_4674);
xnor U8570 (N_8570,N_3160,N_4290);
or U8571 (N_8571,N_3970,N_5862);
nand U8572 (N_8572,N_5877,N_5161);
and U8573 (N_8573,N_3950,N_5645);
xnor U8574 (N_8574,N_4537,N_5107);
nand U8575 (N_8575,N_3270,N_4382);
xor U8576 (N_8576,N_4282,N_4341);
and U8577 (N_8577,N_3427,N_4454);
and U8578 (N_8578,N_4962,N_4204);
xnor U8579 (N_8579,N_4582,N_4020);
nor U8580 (N_8580,N_5823,N_5337);
xnor U8581 (N_8581,N_5017,N_5981);
nor U8582 (N_8582,N_3416,N_4701);
or U8583 (N_8583,N_3341,N_5174);
nor U8584 (N_8584,N_5029,N_4426);
nand U8585 (N_8585,N_4572,N_4862);
nand U8586 (N_8586,N_4016,N_5162);
xnor U8587 (N_8587,N_3444,N_5854);
or U8588 (N_8588,N_3643,N_5025);
or U8589 (N_8589,N_3498,N_5990);
nor U8590 (N_8590,N_4280,N_5942);
nand U8591 (N_8591,N_3783,N_4240);
nor U8592 (N_8592,N_5864,N_5809);
nor U8593 (N_8593,N_4086,N_3714);
xnor U8594 (N_8594,N_3833,N_5815);
xor U8595 (N_8595,N_4469,N_4570);
or U8596 (N_8596,N_4198,N_3950);
nand U8597 (N_8597,N_4837,N_3215);
nor U8598 (N_8598,N_3894,N_5795);
xnor U8599 (N_8599,N_4058,N_5770);
nand U8600 (N_8600,N_3214,N_5668);
nor U8601 (N_8601,N_3509,N_4018);
nor U8602 (N_8602,N_3559,N_5790);
and U8603 (N_8603,N_5867,N_3235);
and U8604 (N_8604,N_5068,N_4721);
and U8605 (N_8605,N_4334,N_5039);
xor U8606 (N_8606,N_4173,N_5453);
or U8607 (N_8607,N_5763,N_3792);
or U8608 (N_8608,N_5073,N_4193);
and U8609 (N_8609,N_3527,N_5818);
nor U8610 (N_8610,N_4076,N_4696);
and U8611 (N_8611,N_5808,N_4053);
xnor U8612 (N_8612,N_5167,N_4256);
and U8613 (N_8613,N_5653,N_4446);
and U8614 (N_8614,N_3789,N_4665);
and U8615 (N_8615,N_5723,N_3584);
nor U8616 (N_8616,N_3487,N_3617);
nand U8617 (N_8617,N_5663,N_3797);
or U8618 (N_8618,N_4188,N_5342);
and U8619 (N_8619,N_4420,N_3870);
nor U8620 (N_8620,N_3264,N_3633);
nor U8621 (N_8621,N_5397,N_5948);
nand U8622 (N_8622,N_5296,N_5190);
and U8623 (N_8623,N_5141,N_4615);
xnor U8624 (N_8624,N_4001,N_5358);
nand U8625 (N_8625,N_3623,N_5248);
xnor U8626 (N_8626,N_3531,N_3707);
and U8627 (N_8627,N_3865,N_3590);
xor U8628 (N_8628,N_4188,N_3042);
and U8629 (N_8629,N_3592,N_5205);
or U8630 (N_8630,N_5888,N_3653);
nor U8631 (N_8631,N_5740,N_5380);
and U8632 (N_8632,N_4608,N_4457);
nor U8633 (N_8633,N_4058,N_3427);
nor U8634 (N_8634,N_4873,N_3273);
nand U8635 (N_8635,N_4692,N_3404);
or U8636 (N_8636,N_4324,N_4835);
or U8637 (N_8637,N_4587,N_4382);
xor U8638 (N_8638,N_5028,N_5155);
nand U8639 (N_8639,N_3244,N_5051);
or U8640 (N_8640,N_4989,N_4716);
xor U8641 (N_8641,N_4605,N_5891);
xor U8642 (N_8642,N_3272,N_4927);
xnor U8643 (N_8643,N_5021,N_4426);
nand U8644 (N_8644,N_4186,N_3608);
nor U8645 (N_8645,N_3930,N_3231);
or U8646 (N_8646,N_3536,N_5262);
nor U8647 (N_8647,N_5790,N_4429);
nor U8648 (N_8648,N_4130,N_4453);
or U8649 (N_8649,N_5141,N_4816);
or U8650 (N_8650,N_3990,N_5500);
and U8651 (N_8651,N_4366,N_4986);
xor U8652 (N_8652,N_5887,N_5639);
xor U8653 (N_8653,N_4511,N_3483);
nor U8654 (N_8654,N_5400,N_4042);
xnor U8655 (N_8655,N_3240,N_4660);
or U8656 (N_8656,N_5605,N_4552);
nor U8657 (N_8657,N_4498,N_4797);
xor U8658 (N_8658,N_4972,N_5068);
or U8659 (N_8659,N_5264,N_4635);
nand U8660 (N_8660,N_4325,N_3147);
nor U8661 (N_8661,N_3159,N_3330);
xnor U8662 (N_8662,N_3214,N_3415);
xnor U8663 (N_8663,N_4203,N_4118);
or U8664 (N_8664,N_4406,N_5676);
nor U8665 (N_8665,N_5567,N_5588);
nand U8666 (N_8666,N_5961,N_5462);
or U8667 (N_8667,N_5331,N_4042);
nor U8668 (N_8668,N_3267,N_5885);
or U8669 (N_8669,N_5128,N_4770);
nand U8670 (N_8670,N_3615,N_4816);
xor U8671 (N_8671,N_5881,N_4590);
nand U8672 (N_8672,N_4514,N_5038);
or U8673 (N_8673,N_3621,N_3912);
or U8674 (N_8674,N_3635,N_5450);
xnor U8675 (N_8675,N_5375,N_3145);
nand U8676 (N_8676,N_5724,N_3983);
nand U8677 (N_8677,N_5378,N_4014);
xor U8678 (N_8678,N_4733,N_4811);
and U8679 (N_8679,N_4701,N_4644);
nor U8680 (N_8680,N_3017,N_4183);
or U8681 (N_8681,N_5122,N_4767);
or U8682 (N_8682,N_4355,N_5822);
and U8683 (N_8683,N_3309,N_4648);
nor U8684 (N_8684,N_3627,N_5265);
nand U8685 (N_8685,N_4294,N_3114);
and U8686 (N_8686,N_4158,N_4807);
nor U8687 (N_8687,N_3309,N_4060);
or U8688 (N_8688,N_3411,N_5694);
xor U8689 (N_8689,N_5028,N_4608);
nand U8690 (N_8690,N_3034,N_4428);
and U8691 (N_8691,N_5261,N_4504);
and U8692 (N_8692,N_3815,N_5622);
and U8693 (N_8693,N_3202,N_4653);
xnor U8694 (N_8694,N_4193,N_3434);
nor U8695 (N_8695,N_5795,N_3881);
or U8696 (N_8696,N_3568,N_4444);
and U8697 (N_8697,N_3936,N_3351);
nand U8698 (N_8698,N_4502,N_5386);
or U8699 (N_8699,N_5419,N_5451);
nor U8700 (N_8700,N_4072,N_3916);
xnor U8701 (N_8701,N_5703,N_3163);
or U8702 (N_8702,N_3979,N_3245);
or U8703 (N_8703,N_3536,N_5027);
and U8704 (N_8704,N_3513,N_5287);
or U8705 (N_8705,N_3979,N_3300);
and U8706 (N_8706,N_3876,N_3865);
nor U8707 (N_8707,N_5306,N_4129);
nand U8708 (N_8708,N_4986,N_5770);
or U8709 (N_8709,N_3572,N_5111);
nand U8710 (N_8710,N_4370,N_5670);
xor U8711 (N_8711,N_3374,N_4872);
nor U8712 (N_8712,N_3676,N_4541);
and U8713 (N_8713,N_3557,N_3639);
or U8714 (N_8714,N_5429,N_4322);
nor U8715 (N_8715,N_5004,N_5160);
nand U8716 (N_8716,N_5344,N_5719);
nand U8717 (N_8717,N_3690,N_5948);
and U8718 (N_8718,N_5527,N_5032);
nor U8719 (N_8719,N_3828,N_4312);
xnor U8720 (N_8720,N_3894,N_4793);
nor U8721 (N_8721,N_4424,N_5517);
xnor U8722 (N_8722,N_3818,N_5023);
or U8723 (N_8723,N_3892,N_3477);
nor U8724 (N_8724,N_3971,N_5926);
or U8725 (N_8725,N_5026,N_3190);
xnor U8726 (N_8726,N_3142,N_5260);
nor U8727 (N_8727,N_4179,N_4730);
and U8728 (N_8728,N_5066,N_3508);
nor U8729 (N_8729,N_3266,N_3102);
and U8730 (N_8730,N_4556,N_3997);
xor U8731 (N_8731,N_5807,N_5438);
or U8732 (N_8732,N_5553,N_5304);
nor U8733 (N_8733,N_5216,N_3237);
nand U8734 (N_8734,N_5330,N_4570);
nor U8735 (N_8735,N_5548,N_3215);
and U8736 (N_8736,N_3492,N_4738);
and U8737 (N_8737,N_5268,N_3951);
or U8738 (N_8738,N_4969,N_3966);
and U8739 (N_8739,N_3512,N_5439);
nand U8740 (N_8740,N_3357,N_5548);
or U8741 (N_8741,N_5126,N_5897);
nand U8742 (N_8742,N_5704,N_3267);
or U8743 (N_8743,N_5590,N_3019);
nand U8744 (N_8744,N_3288,N_5232);
nor U8745 (N_8745,N_3942,N_5574);
nor U8746 (N_8746,N_5682,N_3677);
nor U8747 (N_8747,N_3984,N_5793);
or U8748 (N_8748,N_4492,N_3050);
or U8749 (N_8749,N_3730,N_4623);
or U8750 (N_8750,N_3479,N_3901);
nor U8751 (N_8751,N_4757,N_3521);
or U8752 (N_8752,N_4552,N_5661);
xor U8753 (N_8753,N_3909,N_5834);
xor U8754 (N_8754,N_5069,N_3420);
and U8755 (N_8755,N_3335,N_5325);
xnor U8756 (N_8756,N_3180,N_4477);
or U8757 (N_8757,N_3211,N_3311);
nor U8758 (N_8758,N_5756,N_4818);
xnor U8759 (N_8759,N_3211,N_4376);
or U8760 (N_8760,N_3241,N_4009);
or U8761 (N_8761,N_4904,N_4102);
xnor U8762 (N_8762,N_5672,N_3633);
nand U8763 (N_8763,N_3478,N_3367);
xnor U8764 (N_8764,N_3813,N_4629);
and U8765 (N_8765,N_5764,N_4855);
xor U8766 (N_8766,N_4907,N_4356);
xnor U8767 (N_8767,N_5426,N_5556);
nor U8768 (N_8768,N_3352,N_4031);
nand U8769 (N_8769,N_5796,N_5678);
and U8770 (N_8770,N_5208,N_4487);
nor U8771 (N_8771,N_5501,N_3479);
xor U8772 (N_8772,N_4985,N_4774);
nor U8773 (N_8773,N_3378,N_5328);
and U8774 (N_8774,N_3752,N_5159);
nor U8775 (N_8775,N_3789,N_3956);
xnor U8776 (N_8776,N_4147,N_4188);
or U8777 (N_8777,N_3352,N_5736);
and U8778 (N_8778,N_5553,N_4204);
nor U8779 (N_8779,N_3381,N_5989);
and U8780 (N_8780,N_3209,N_4166);
xor U8781 (N_8781,N_4127,N_3480);
nor U8782 (N_8782,N_3926,N_4684);
nor U8783 (N_8783,N_5334,N_3571);
xnor U8784 (N_8784,N_3682,N_4965);
nor U8785 (N_8785,N_3411,N_5447);
nand U8786 (N_8786,N_5641,N_3368);
or U8787 (N_8787,N_5638,N_5284);
xor U8788 (N_8788,N_4344,N_5018);
xnor U8789 (N_8789,N_3020,N_4504);
and U8790 (N_8790,N_3901,N_3809);
or U8791 (N_8791,N_5633,N_4321);
or U8792 (N_8792,N_5669,N_3354);
nor U8793 (N_8793,N_4612,N_3839);
and U8794 (N_8794,N_5608,N_3190);
nand U8795 (N_8795,N_4370,N_5888);
nor U8796 (N_8796,N_3771,N_5950);
xnor U8797 (N_8797,N_5522,N_5243);
xor U8798 (N_8798,N_4098,N_5878);
xor U8799 (N_8799,N_5050,N_3389);
xnor U8800 (N_8800,N_4044,N_4919);
nor U8801 (N_8801,N_5189,N_3453);
and U8802 (N_8802,N_3570,N_4108);
nor U8803 (N_8803,N_3708,N_5903);
nand U8804 (N_8804,N_5986,N_3816);
or U8805 (N_8805,N_3054,N_5612);
and U8806 (N_8806,N_3363,N_3375);
nand U8807 (N_8807,N_5465,N_4983);
or U8808 (N_8808,N_3764,N_4117);
xnor U8809 (N_8809,N_3686,N_3547);
or U8810 (N_8810,N_5079,N_4485);
or U8811 (N_8811,N_3600,N_4682);
nand U8812 (N_8812,N_5358,N_5682);
nand U8813 (N_8813,N_3017,N_3347);
nand U8814 (N_8814,N_5584,N_5404);
and U8815 (N_8815,N_5710,N_4560);
xnor U8816 (N_8816,N_4473,N_3742);
and U8817 (N_8817,N_5363,N_3534);
or U8818 (N_8818,N_5347,N_5583);
nor U8819 (N_8819,N_5695,N_4808);
nor U8820 (N_8820,N_4648,N_3713);
or U8821 (N_8821,N_4838,N_3787);
xor U8822 (N_8822,N_3960,N_4664);
xnor U8823 (N_8823,N_3164,N_3615);
and U8824 (N_8824,N_3754,N_5128);
and U8825 (N_8825,N_5494,N_4216);
or U8826 (N_8826,N_4712,N_4208);
or U8827 (N_8827,N_4553,N_3956);
xor U8828 (N_8828,N_5545,N_3666);
or U8829 (N_8829,N_3733,N_4789);
xnor U8830 (N_8830,N_3121,N_5746);
or U8831 (N_8831,N_4502,N_4354);
and U8832 (N_8832,N_4629,N_3331);
or U8833 (N_8833,N_5172,N_5253);
xor U8834 (N_8834,N_5116,N_5168);
or U8835 (N_8835,N_4200,N_4949);
and U8836 (N_8836,N_5814,N_5588);
xnor U8837 (N_8837,N_5799,N_5937);
or U8838 (N_8838,N_3419,N_3757);
xnor U8839 (N_8839,N_3646,N_3488);
xor U8840 (N_8840,N_4619,N_4316);
nand U8841 (N_8841,N_4824,N_5690);
or U8842 (N_8842,N_5589,N_5897);
and U8843 (N_8843,N_4254,N_3409);
or U8844 (N_8844,N_5485,N_3520);
and U8845 (N_8845,N_4663,N_5182);
and U8846 (N_8846,N_3910,N_3619);
xor U8847 (N_8847,N_4622,N_5942);
nand U8848 (N_8848,N_3292,N_5575);
and U8849 (N_8849,N_4922,N_3993);
and U8850 (N_8850,N_4406,N_4601);
or U8851 (N_8851,N_3434,N_5166);
nand U8852 (N_8852,N_4152,N_3257);
xnor U8853 (N_8853,N_4680,N_5748);
xor U8854 (N_8854,N_5398,N_5898);
xor U8855 (N_8855,N_3917,N_5214);
and U8856 (N_8856,N_4608,N_4739);
nor U8857 (N_8857,N_5383,N_3565);
and U8858 (N_8858,N_4675,N_3385);
xnor U8859 (N_8859,N_5160,N_5210);
nand U8860 (N_8860,N_4758,N_3540);
or U8861 (N_8861,N_3897,N_3709);
nor U8862 (N_8862,N_5582,N_4030);
and U8863 (N_8863,N_4575,N_5572);
or U8864 (N_8864,N_3662,N_4657);
nand U8865 (N_8865,N_3367,N_4216);
xnor U8866 (N_8866,N_3285,N_5323);
nand U8867 (N_8867,N_4099,N_5883);
nor U8868 (N_8868,N_3454,N_4698);
nand U8869 (N_8869,N_3327,N_4176);
xnor U8870 (N_8870,N_5459,N_5335);
nand U8871 (N_8871,N_4725,N_5546);
nand U8872 (N_8872,N_4475,N_3902);
nor U8873 (N_8873,N_5558,N_4940);
and U8874 (N_8874,N_5600,N_4517);
xor U8875 (N_8875,N_4947,N_5850);
or U8876 (N_8876,N_5303,N_5806);
or U8877 (N_8877,N_3452,N_5547);
nand U8878 (N_8878,N_3582,N_5869);
nor U8879 (N_8879,N_3415,N_3467);
or U8880 (N_8880,N_4358,N_5057);
or U8881 (N_8881,N_4619,N_3723);
and U8882 (N_8882,N_5750,N_5291);
or U8883 (N_8883,N_5455,N_4959);
and U8884 (N_8884,N_5829,N_4183);
xor U8885 (N_8885,N_4731,N_5443);
and U8886 (N_8886,N_3722,N_4217);
or U8887 (N_8887,N_3316,N_3025);
or U8888 (N_8888,N_3548,N_4127);
and U8889 (N_8889,N_5748,N_3556);
nand U8890 (N_8890,N_3128,N_4893);
or U8891 (N_8891,N_3951,N_3062);
xor U8892 (N_8892,N_4807,N_5657);
and U8893 (N_8893,N_3671,N_4228);
or U8894 (N_8894,N_5836,N_4279);
and U8895 (N_8895,N_4085,N_3651);
nor U8896 (N_8896,N_3696,N_5854);
nand U8897 (N_8897,N_4204,N_4539);
and U8898 (N_8898,N_3245,N_3605);
and U8899 (N_8899,N_5452,N_3485);
or U8900 (N_8900,N_3268,N_4172);
or U8901 (N_8901,N_5824,N_4944);
xnor U8902 (N_8902,N_3366,N_5610);
xor U8903 (N_8903,N_4405,N_5542);
and U8904 (N_8904,N_3897,N_5579);
nor U8905 (N_8905,N_4844,N_3983);
nor U8906 (N_8906,N_3809,N_3658);
xor U8907 (N_8907,N_3514,N_4264);
or U8908 (N_8908,N_5567,N_5123);
or U8909 (N_8909,N_4021,N_3120);
nor U8910 (N_8910,N_5031,N_4278);
or U8911 (N_8911,N_3020,N_3730);
xnor U8912 (N_8912,N_3862,N_5183);
nand U8913 (N_8913,N_3145,N_3682);
nand U8914 (N_8914,N_5319,N_3253);
nor U8915 (N_8915,N_4837,N_3104);
nand U8916 (N_8916,N_3305,N_5601);
nor U8917 (N_8917,N_3324,N_3036);
and U8918 (N_8918,N_4764,N_4099);
nand U8919 (N_8919,N_4122,N_3566);
xor U8920 (N_8920,N_5274,N_4935);
and U8921 (N_8921,N_3204,N_3631);
or U8922 (N_8922,N_5630,N_4671);
xnor U8923 (N_8923,N_4640,N_5116);
nand U8924 (N_8924,N_5964,N_3050);
or U8925 (N_8925,N_4033,N_5512);
nand U8926 (N_8926,N_5484,N_5840);
and U8927 (N_8927,N_3498,N_3906);
and U8928 (N_8928,N_5787,N_5755);
or U8929 (N_8929,N_4881,N_3824);
or U8930 (N_8930,N_4938,N_4191);
or U8931 (N_8931,N_3029,N_5081);
and U8932 (N_8932,N_3604,N_4149);
or U8933 (N_8933,N_4162,N_5406);
nand U8934 (N_8934,N_3187,N_3054);
or U8935 (N_8935,N_3531,N_3988);
nor U8936 (N_8936,N_3969,N_4281);
xnor U8937 (N_8937,N_3474,N_5071);
or U8938 (N_8938,N_4445,N_3633);
nor U8939 (N_8939,N_3925,N_5347);
nor U8940 (N_8940,N_4794,N_5614);
nand U8941 (N_8941,N_5679,N_3274);
or U8942 (N_8942,N_4532,N_5597);
nand U8943 (N_8943,N_5883,N_4635);
and U8944 (N_8944,N_4421,N_3062);
nor U8945 (N_8945,N_3422,N_3338);
or U8946 (N_8946,N_4613,N_5000);
or U8947 (N_8947,N_5353,N_3724);
and U8948 (N_8948,N_3788,N_3607);
nand U8949 (N_8949,N_4343,N_3100);
nand U8950 (N_8950,N_4807,N_4860);
nand U8951 (N_8951,N_3331,N_4245);
nor U8952 (N_8952,N_3578,N_5699);
or U8953 (N_8953,N_3542,N_4785);
and U8954 (N_8954,N_4911,N_3152);
or U8955 (N_8955,N_3553,N_5899);
or U8956 (N_8956,N_5007,N_5225);
and U8957 (N_8957,N_3087,N_5147);
nor U8958 (N_8958,N_3916,N_3389);
nor U8959 (N_8959,N_3030,N_3561);
and U8960 (N_8960,N_4996,N_4821);
nand U8961 (N_8961,N_4428,N_4890);
xor U8962 (N_8962,N_3099,N_3995);
nor U8963 (N_8963,N_4008,N_4392);
and U8964 (N_8964,N_5395,N_5728);
or U8965 (N_8965,N_5772,N_5113);
or U8966 (N_8966,N_5509,N_3155);
xnor U8967 (N_8967,N_4837,N_3917);
xor U8968 (N_8968,N_3756,N_4893);
nand U8969 (N_8969,N_5567,N_5094);
or U8970 (N_8970,N_5191,N_3394);
nand U8971 (N_8971,N_3649,N_3565);
xor U8972 (N_8972,N_3208,N_4571);
xor U8973 (N_8973,N_5158,N_5174);
nand U8974 (N_8974,N_3496,N_4530);
nor U8975 (N_8975,N_5939,N_4738);
nand U8976 (N_8976,N_4084,N_4585);
or U8977 (N_8977,N_5175,N_3321);
or U8978 (N_8978,N_4323,N_3308);
or U8979 (N_8979,N_5204,N_4491);
nor U8980 (N_8980,N_4544,N_4427);
nor U8981 (N_8981,N_4216,N_4566);
and U8982 (N_8982,N_4814,N_4735);
xor U8983 (N_8983,N_3376,N_4414);
nor U8984 (N_8984,N_5624,N_4206);
xor U8985 (N_8985,N_4912,N_3536);
nor U8986 (N_8986,N_3465,N_3262);
nand U8987 (N_8987,N_3594,N_3835);
nand U8988 (N_8988,N_4047,N_3631);
or U8989 (N_8989,N_3122,N_5572);
and U8990 (N_8990,N_5243,N_4416);
xor U8991 (N_8991,N_5403,N_3102);
or U8992 (N_8992,N_3162,N_4852);
and U8993 (N_8993,N_3524,N_4894);
and U8994 (N_8994,N_4000,N_3898);
nand U8995 (N_8995,N_4384,N_3545);
xnor U8996 (N_8996,N_5711,N_4773);
nor U8997 (N_8997,N_5002,N_4540);
and U8998 (N_8998,N_5053,N_3264);
nor U8999 (N_8999,N_3290,N_5265);
and U9000 (N_9000,N_6511,N_7977);
and U9001 (N_9001,N_8818,N_7059);
xnor U9002 (N_9002,N_8213,N_6958);
and U9003 (N_9003,N_6514,N_8290);
xnor U9004 (N_9004,N_7934,N_7857);
nor U9005 (N_9005,N_6712,N_6944);
nor U9006 (N_9006,N_8266,N_8583);
nand U9007 (N_9007,N_7657,N_7118);
and U9008 (N_9008,N_7963,N_6593);
nand U9009 (N_9009,N_7204,N_6885);
xor U9010 (N_9010,N_8298,N_6891);
nand U9011 (N_9011,N_6683,N_8069);
and U9012 (N_9012,N_6191,N_6022);
xor U9013 (N_9013,N_6829,N_7948);
xor U9014 (N_9014,N_7903,N_6259);
or U9015 (N_9015,N_8557,N_8270);
or U9016 (N_9016,N_7980,N_7699);
nor U9017 (N_9017,N_8684,N_6541);
xnor U9018 (N_9018,N_6933,N_6008);
nor U9019 (N_9019,N_8620,N_7420);
and U9020 (N_9020,N_7325,N_6006);
nand U9021 (N_9021,N_6711,N_7203);
or U9022 (N_9022,N_8842,N_6677);
or U9023 (N_9023,N_8797,N_7408);
nand U9024 (N_9024,N_8956,N_8005);
or U9025 (N_9025,N_6974,N_8918);
nor U9026 (N_9026,N_8475,N_8963);
or U9027 (N_9027,N_8057,N_6169);
or U9028 (N_9028,N_7061,N_7532);
xnor U9029 (N_9029,N_7080,N_8606);
and U9030 (N_9030,N_7888,N_8470);
and U9031 (N_9031,N_7595,N_6109);
xor U9032 (N_9032,N_7205,N_7904);
and U9033 (N_9033,N_6399,N_6066);
and U9034 (N_9034,N_7232,N_8959);
xor U9035 (N_9035,N_6766,N_6285);
xor U9036 (N_9036,N_8838,N_8616);
or U9037 (N_9037,N_7721,N_8677);
or U9038 (N_9038,N_8917,N_6681);
xor U9039 (N_9039,N_7461,N_8232);
nand U9040 (N_9040,N_6192,N_8610);
and U9041 (N_9041,N_7466,N_6032);
nor U9042 (N_9042,N_7833,N_7747);
nand U9043 (N_9043,N_7083,N_8191);
and U9044 (N_9044,N_8722,N_6397);
nor U9045 (N_9045,N_8010,N_6557);
or U9046 (N_9046,N_6193,N_6709);
nand U9047 (N_9047,N_8467,N_6838);
xor U9048 (N_9048,N_6143,N_8612);
nor U9049 (N_9049,N_8679,N_6645);
nor U9050 (N_9050,N_8229,N_8405);
nor U9051 (N_9051,N_6433,N_7592);
and U9052 (N_9052,N_6135,N_6226);
or U9053 (N_9053,N_6505,N_6095);
and U9054 (N_9054,N_7445,N_8389);
or U9055 (N_9055,N_6884,N_6435);
or U9056 (N_9056,N_7809,N_6993);
nand U9057 (N_9057,N_6189,N_6003);
xor U9058 (N_9058,N_6756,N_8782);
or U9059 (N_9059,N_8170,N_8989);
nor U9060 (N_9060,N_6897,N_6662);
and U9061 (N_9061,N_6949,N_7503);
nor U9062 (N_9062,N_8273,N_8481);
nand U9063 (N_9063,N_6940,N_8625);
xor U9064 (N_9064,N_6020,N_7051);
xnor U9065 (N_9065,N_7633,N_8385);
or U9066 (N_9066,N_6001,N_7071);
and U9067 (N_9067,N_8310,N_8231);
nand U9068 (N_9068,N_6607,N_7358);
nand U9069 (N_9069,N_6333,N_6782);
and U9070 (N_9070,N_8940,N_8076);
xor U9071 (N_9071,N_7309,N_8638);
and U9072 (N_9072,N_7910,N_7546);
nand U9073 (N_9073,N_6195,N_7797);
nor U9074 (N_9074,N_7545,N_7818);
xnor U9075 (N_9075,N_7561,N_7007);
nand U9076 (N_9076,N_8947,N_8858);
xor U9077 (N_9077,N_8082,N_8168);
xnor U9078 (N_9078,N_7851,N_8631);
xor U9079 (N_9079,N_7054,N_6786);
nor U9080 (N_9080,N_6703,N_6754);
or U9081 (N_9081,N_8259,N_8516);
and U9082 (N_9082,N_8787,N_6350);
or U9083 (N_9083,N_8707,N_8255);
nor U9084 (N_9084,N_8223,N_7202);
and U9085 (N_9085,N_8379,N_8401);
or U9086 (N_9086,N_8330,N_8466);
or U9087 (N_9087,N_6159,N_8031);
nor U9088 (N_9088,N_8474,N_8404);
or U9089 (N_9089,N_8868,N_6826);
or U9090 (N_9090,N_7612,N_8418);
nor U9091 (N_9091,N_6905,N_7622);
nor U9092 (N_9092,N_6516,N_8196);
xor U9093 (N_9093,N_6706,N_6243);
and U9094 (N_9094,N_6956,N_7498);
xnor U9095 (N_9095,N_6018,N_8634);
or U9096 (N_9096,N_8975,N_7748);
nor U9097 (N_9097,N_7336,N_8629);
nand U9098 (N_9098,N_7429,N_6911);
nor U9099 (N_9099,N_8655,N_7608);
xnor U9100 (N_9100,N_6459,N_8119);
nand U9101 (N_9101,N_6443,N_6051);
nor U9102 (N_9102,N_6871,N_6305);
and U9103 (N_9103,N_7401,N_7655);
xnor U9104 (N_9104,N_7572,N_7342);
or U9105 (N_9105,N_6724,N_7823);
xor U9106 (N_9106,N_8957,N_8443);
nor U9107 (N_9107,N_6306,N_6280);
nand U9108 (N_9108,N_7653,N_7192);
and U9109 (N_9109,N_6233,N_6722);
nand U9110 (N_9110,N_7994,N_7368);
or U9111 (N_9111,N_6588,N_8400);
and U9112 (N_9112,N_7863,N_6733);
nand U9113 (N_9113,N_7951,N_8598);
or U9114 (N_9114,N_6598,N_6361);
nand U9115 (N_9115,N_6522,N_8575);
and U9116 (N_9116,N_6980,N_6811);
xnor U9117 (N_9117,N_7236,N_8427);
nor U9118 (N_9118,N_6047,N_8271);
nand U9119 (N_9119,N_8128,N_8942);
nand U9120 (N_9120,N_8499,N_6672);
and U9121 (N_9121,N_8827,N_7104);
and U9122 (N_9122,N_8225,N_7941);
xnor U9123 (N_9123,N_8632,N_7933);
or U9124 (N_9124,N_8037,N_7929);
nand U9125 (N_9125,N_7257,N_7046);
nand U9126 (N_9126,N_7898,N_8094);
or U9127 (N_9127,N_6465,N_8413);
nand U9128 (N_9128,N_8072,N_8214);
nand U9129 (N_9129,N_6988,N_7850);
and U9130 (N_9130,N_7506,N_8239);
or U9131 (N_9131,N_7728,N_7154);
and U9132 (N_9132,N_8760,N_8093);
nor U9133 (N_9133,N_7892,N_7844);
or U9134 (N_9134,N_8162,N_7637);
xnor U9135 (N_9135,N_8314,N_6021);
xor U9136 (N_9136,N_7835,N_6416);
nor U9137 (N_9137,N_8185,N_7399);
xnor U9138 (N_9138,N_6521,N_6320);
nand U9139 (N_9139,N_7463,N_7746);
and U9140 (N_9140,N_7878,N_7226);
nand U9141 (N_9141,N_7068,N_6610);
nand U9142 (N_9142,N_8830,N_8937);
nor U9143 (N_9143,N_8016,N_8786);
xnor U9144 (N_9144,N_6764,N_6542);
xor U9145 (N_9145,N_6673,N_8546);
nand U9146 (N_9146,N_7028,N_7263);
nand U9147 (N_9147,N_7596,N_7352);
or U9148 (N_9148,N_7162,N_6346);
xnor U9149 (N_9149,N_7604,N_7533);
nor U9150 (N_9150,N_6262,N_6242);
and U9151 (N_9151,N_7914,N_6369);
and U9152 (N_9152,N_8837,N_7122);
nor U9153 (N_9153,N_6410,N_6312);
nand U9154 (N_9154,N_8052,N_6422);
nand U9155 (N_9155,N_7393,N_8608);
or U9156 (N_9156,N_8884,N_7534);
xnor U9157 (N_9157,N_8784,N_7755);
nand U9158 (N_9158,N_7765,N_7098);
and U9159 (N_9159,N_7187,N_8995);
nand U9160 (N_9160,N_8179,N_6310);
nand U9161 (N_9161,N_8319,N_6668);
and U9162 (N_9162,N_6821,N_7185);
or U9163 (N_9163,N_8504,N_6245);
xnor U9164 (N_9164,N_8484,N_8030);
and U9165 (N_9165,N_6094,N_8049);
and U9166 (N_9166,N_7978,N_8727);
xnor U9167 (N_9167,N_8805,N_6752);
xor U9168 (N_9168,N_7489,N_6629);
and U9169 (N_9169,N_7846,N_8336);
xnor U9170 (N_9170,N_6458,N_7327);
nor U9171 (N_9171,N_7491,N_8067);
and U9172 (N_9172,N_6042,N_6418);
nand U9173 (N_9173,N_6656,N_7740);
nor U9174 (N_9174,N_6163,N_6792);
or U9175 (N_9175,N_7119,N_7509);
and U9176 (N_9176,N_6105,N_6406);
nor U9177 (N_9177,N_8735,N_7411);
nand U9178 (N_9178,N_6166,N_6248);
nand U9179 (N_9179,N_8023,N_7126);
and U9180 (N_9180,N_7344,N_8145);
and U9181 (N_9181,N_8397,N_8253);
or U9182 (N_9182,N_6460,N_6010);
nor U9183 (N_9183,N_8437,N_7547);
and U9184 (N_9184,N_8833,N_7855);
nand U9185 (N_9185,N_6247,N_7840);
or U9186 (N_9186,N_8494,N_6295);
and U9187 (N_9187,N_8251,N_8566);
and U9188 (N_9188,N_8083,N_8247);
xor U9189 (N_9189,N_8487,N_6383);
nor U9190 (N_9190,N_7548,N_8012);
nand U9191 (N_9191,N_6049,N_6358);
nand U9192 (N_9192,N_6064,N_8281);
and U9193 (N_9193,N_7177,N_6203);
nand U9194 (N_9194,N_7998,N_8647);
or U9195 (N_9195,N_8525,N_6217);
and U9196 (N_9196,N_7551,N_8421);
nor U9197 (N_9197,N_8038,N_6874);
and U9198 (N_9198,N_6876,N_6145);
xnor U9199 (N_9199,N_6196,N_8372);
and U9200 (N_9200,N_6405,N_6033);
and U9201 (N_9201,N_7381,N_8131);
and U9202 (N_9202,N_8801,N_6715);
or U9203 (N_9203,N_8406,N_8249);
xnor U9204 (N_9204,N_7219,N_6046);
and U9205 (N_9205,N_6809,N_6293);
xnor U9206 (N_9206,N_8855,N_6455);
xor U9207 (N_9207,N_7813,N_8994);
or U9208 (N_9208,N_7335,N_8976);
nand U9209 (N_9209,N_7673,N_8667);
nand U9210 (N_9210,N_8682,N_7820);
and U9211 (N_9211,N_7964,N_8831);
and U9212 (N_9212,N_7238,N_7026);
xor U9213 (N_9213,N_7583,N_8199);
nand U9214 (N_9214,N_8071,N_6990);
xnor U9215 (N_9215,N_6206,N_7827);
xor U9216 (N_9216,N_7448,N_6190);
nor U9217 (N_9217,N_7379,N_6849);
and U9218 (N_9218,N_8675,N_6776);
nor U9219 (N_9219,N_6844,N_7953);
nand U9220 (N_9220,N_8844,N_6583);
and U9221 (N_9221,N_6537,N_7896);
xor U9222 (N_9222,N_8154,N_8045);
nand U9223 (N_9223,N_8283,N_6146);
nand U9224 (N_9224,N_6496,N_7101);
and U9225 (N_9225,N_7213,N_6710);
or U9226 (N_9226,N_8498,N_8116);
and U9227 (N_9227,N_7067,N_8680);
xnor U9228 (N_9228,N_7306,N_6225);
and U9229 (N_9229,N_6340,N_7178);
xnor U9230 (N_9230,N_6650,N_7716);
nand U9231 (N_9231,N_8936,N_8316);
xnor U9232 (N_9232,N_6533,N_7175);
xor U9233 (N_9233,N_7714,N_6393);
or U9234 (N_9234,N_7758,N_6401);
xor U9235 (N_9235,N_8099,N_6915);
and U9236 (N_9236,N_8890,N_6117);
and U9237 (N_9237,N_8803,N_8408);
nand U9238 (N_9238,N_8384,N_8268);
or U9239 (N_9239,N_8350,N_8896);
nand U9240 (N_9240,N_8780,N_8866);
nor U9241 (N_9241,N_6917,N_8469);
and U9242 (N_9242,N_7666,N_6270);
nor U9243 (N_9243,N_7042,N_6743);
or U9244 (N_9244,N_7974,N_6556);
nor U9245 (N_9245,N_6512,N_7412);
xor U9246 (N_9246,N_8690,N_8501);
and U9247 (N_9247,N_7522,N_8258);
and U9248 (N_9248,N_8059,N_8870);
nand U9249 (N_9249,N_6799,N_7705);
nand U9250 (N_9250,N_7012,N_6255);
nand U9251 (N_9251,N_8476,N_8195);
and U9252 (N_9252,N_7826,N_8013);
or U9253 (N_9253,N_7004,N_8799);
xor U9254 (N_9254,N_7879,N_7337);
nor U9255 (N_9255,N_8233,N_7750);
or U9256 (N_9256,N_6419,N_6395);
xor U9257 (N_9257,N_8718,N_8303);
or U9258 (N_9258,N_8627,N_8519);
xnor U9259 (N_9259,N_8553,N_8449);
nand U9260 (N_9260,N_8361,N_8728);
xor U9261 (N_9261,N_8674,N_6814);
and U9262 (N_9262,N_6839,N_7708);
nand U9263 (N_9263,N_6336,N_8441);
and U9264 (N_9264,N_8576,N_8460);
xnor U9265 (N_9265,N_7715,N_8860);
nand U9266 (N_9266,N_8969,N_6274);
xor U9267 (N_9267,N_7233,N_8246);
and U9268 (N_9268,N_7663,N_6284);
or U9269 (N_9269,N_7667,N_8104);
nand U9270 (N_9270,N_8160,N_6646);
or U9271 (N_9271,N_7229,N_6755);
or U9272 (N_9272,N_6389,N_7761);
or U9273 (N_9273,N_7348,N_6605);
xor U9274 (N_9274,N_6567,N_6791);
or U9275 (N_9275,N_6981,N_7529);
xor U9276 (N_9276,N_6689,N_7447);
xnor U9277 (N_9277,N_7284,N_8327);
nand U9278 (N_9278,N_7117,N_7693);
or U9279 (N_9279,N_6342,N_8176);
xnor U9280 (N_9280,N_7085,N_8528);
xnor U9281 (N_9281,N_8286,N_8425);
and U9282 (N_9282,N_7505,N_6609);
xor U9283 (N_9283,N_7395,N_6819);
and U9284 (N_9284,N_8177,N_8025);
nand U9285 (N_9285,N_8077,N_8053);
and U9286 (N_9286,N_7485,N_7365);
nand U9287 (N_9287,N_7985,N_7299);
or U9288 (N_9288,N_6173,N_7282);
or U9289 (N_9289,N_8265,N_8946);
nand U9290 (N_9290,N_6843,N_7504);
nand U9291 (N_9291,N_8256,N_6479);
xor U9292 (N_9292,N_7726,N_8112);
nand U9293 (N_9293,N_6977,N_6158);
xor U9294 (N_9294,N_8714,N_7567);
nor U9295 (N_9295,N_6497,N_7323);
nand U9296 (N_9296,N_6337,N_6882);
xor U9297 (N_9297,N_7651,N_8056);
xnor U9298 (N_9298,N_7132,N_7610);
and U9299 (N_9299,N_8597,N_8423);
xnor U9300 (N_9300,N_7450,N_7152);
or U9301 (N_9301,N_6367,N_6235);
xor U9302 (N_9302,N_6761,N_7795);
nand U9303 (N_9303,N_7856,N_8335);
or U9304 (N_9304,N_8088,N_7201);
and U9305 (N_9305,N_6445,N_8141);
nor U9306 (N_9306,N_8894,N_7524);
xnor U9307 (N_9307,N_8121,N_7021);
or U9308 (N_9308,N_6138,N_8245);
or U9309 (N_9309,N_8706,N_8514);
or U9310 (N_9310,N_7273,N_6576);
or U9311 (N_9311,N_8288,N_7707);
and U9312 (N_9312,N_6725,N_8070);
nand U9313 (N_9313,N_7664,N_6936);
or U9314 (N_9314,N_6488,N_6734);
nand U9315 (N_9315,N_6555,N_8346);
nor U9316 (N_9316,N_6691,N_7157);
and U9317 (N_9317,N_7246,N_6631);
xor U9318 (N_9318,N_6589,N_6075);
or U9319 (N_9319,N_8819,N_6078);
nor U9320 (N_9320,N_7292,N_6390);
xnor U9321 (N_9321,N_6851,N_7523);
nor U9322 (N_9322,N_7945,N_6457);
nor U9323 (N_9323,N_7770,N_7718);
nand U9324 (N_9324,N_7940,N_6315);
or U9325 (N_9325,N_7932,N_7156);
nand U9326 (N_9326,N_8793,N_7121);
xor U9327 (N_9327,N_8587,N_6486);
or U9328 (N_9328,N_8923,N_6165);
or U9329 (N_9329,N_6536,N_7609);
and U9330 (N_9330,N_7084,N_6368);
nand U9331 (N_9331,N_6469,N_8186);
nand U9332 (N_9332,N_7731,N_8517);
nand U9333 (N_9333,N_8991,N_7074);
and U9334 (N_9334,N_7375,N_7640);
nor U9335 (N_9335,N_6198,N_8280);
nor U9336 (N_9336,N_7389,N_8895);
nand U9337 (N_9337,N_6881,N_6321);
or U9338 (N_9338,N_6987,N_7993);
xnor U9339 (N_9339,N_6437,N_7573);
xnor U9340 (N_9340,N_8681,N_7488);
nand U9341 (N_9341,N_7115,N_7422);
xnor U9342 (N_9342,N_6113,N_8847);
xor U9343 (N_9343,N_6059,N_8115);
xor U9344 (N_9344,N_8132,N_7931);
nor U9345 (N_9345,N_6836,N_6760);
xor U9346 (N_9346,N_6380,N_6388);
xnor U9347 (N_9347,N_7347,N_8747);
and U9348 (N_9348,N_8986,N_6563);
nor U9349 (N_9349,N_7737,N_7180);
and U9350 (N_9350,N_6124,N_7254);
xnor U9351 (N_9351,N_6114,N_7446);
or U9352 (N_9352,N_7513,N_8163);
nor U9353 (N_9353,N_6942,N_8188);
or U9354 (N_9354,N_6793,N_8834);
and U9355 (N_9355,N_7227,N_6492);
xor U9356 (N_9356,N_7922,N_6526);
nand U9357 (N_9357,N_7882,N_7947);
xor U9358 (N_9358,N_8407,N_8078);
nor U9359 (N_9359,N_7796,N_7486);
nand U9360 (N_9360,N_8430,N_7587);
and U9361 (N_9361,N_8635,N_6702);
nand U9362 (N_9362,N_6149,N_7153);
xnor U9363 (N_9363,N_7698,N_6540);
nand U9364 (N_9364,N_8551,N_7955);
nand U9365 (N_9365,N_8201,N_6498);
xor U9366 (N_9366,N_8712,N_8263);
or U9367 (N_9367,N_8084,N_8355);
nand U9368 (N_9368,N_7217,N_7995);
and U9369 (N_9369,N_8042,N_8457);
nor U9370 (N_9370,N_7671,N_7430);
xnor U9371 (N_9371,N_8447,N_8305);
or U9372 (N_9372,N_6737,N_8720);
nor U9373 (N_9373,N_6220,N_8933);
nand U9374 (N_9374,N_6955,N_6996);
nand U9375 (N_9375,N_7475,N_7790);
and U9376 (N_9376,N_7553,N_7908);
nor U9377 (N_9377,N_8694,N_8017);
and U9378 (N_9378,N_8851,N_7419);
and U9379 (N_9379,N_7366,N_8530);
nor U9380 (N_9380,N_6447,N_7457);
xor U9381 (N_9381,N_6865,N_8966);
and U9382 (N_9382,N_8291,N_8426);
nand U9383 (N_9383,N_6083,N_6510);
and U9384 (N_9384,N_6466,N_8046);
xor U9385 (N_9385,N_7810,N_6575);
nor U9386 (N_9386,N_8843,N_7346);
nand U9387 (N_9387,N_7030,N_8126);
and U9388 (N_9388,N_7597,N_7027);
nor U9389 (N_9389,N_8428,N_7170);
or U9390 (N_9390,N_7570,N_7560);
and U9391 (N_9391,N_6774,N_6900);
and U9392 (N_9392,N_8020,N_8795);
xor U9393 (N_9393,N_6903,N_6532);
or U9394 (N_9394,N_6396,N_8061);
nor U9395 (N_9395,N_8511,N_7946);
or U9396 (N_9396,N_7997,N_8865);
or U9397 (N_9397,N_6129,N_6950);
and U9398 (N_9398,N_6494,N_7741);
xor U9399 (N_9399,N_7191,N_7235);
or U9400 (N_9400,N_8357,N_7063);
nand U9401 (N_9401,N_8565,N_8624);
and U9402 (N_9402,N_7502,N_7989);
xnor U9403 (N_9403,N_8877,N_7973);
or U9404 (N_9404,N_6637,N_6840);
xor U9405 (N_9405,N_6892,N_8526);
nor U9406 (N_9406,N_6595,N_8611);
nand U9407 (N_9407,N_8006,N_7681);
xnor U9408 (N_9408,N_6027,N_8533);
nor U9409 (N_9409,N_8887,N_7869);
or U9410 (N_9410,N_8885,N_8791);
or U9411 (N_9411,N_7926,N_7318);
xnor U9412 (N_9412,N_7853,N_6757);
xor U9413 (N_9413,N_6928,N_6023);
and U9414 (N_9414,N_8338,N_8605);
nor U9415 (N_9415,N_7465,N_7166);
xor U9416 (N_9416,N_7979,N_6824);
nand U9417 (N_9417,N_6197,N_7047);
or U9418 (N_9418,N_7692,N_7555);
or U9419 (N_9419,N_7427,N_8816);
or U9420 (N_9420,N_6954,N_7982);
and U9421 (N_9421,N_7659,N_8452);
xor U9422 (N_9422,N_6810,N_8113);
nand U9423 (N_9423,N_6354,N_8641);
nor U9424 (N_9424,N_7376,N_8987);
nand U9425 (N_9425,N_7064,N_8143);
nor U9426 (N_9426,N_6931,N_7672);
nand U9427 (N_9427,N_8236,N_6922);
xor U9428 (N_9428,N_6670,N_8951);
xnor U9429 (N_9429,N_7537,N_7865);
nand U9430 (N_9430,N_8507,N_6188);
nor U9431 (N_9431,N_6887,N_7848);
nor U9432 (N_9432,N_8783,N_6058);
and U9433 (N_9433,N_6212,N_7276);
nand U9434 (N_9434,N_6326,N_7437);
or U9435 (N_9435,N_8888,N_7009);
or U9436 (N_9436,N_7173,N_6328);
and U9437 (N_9437,N_6485,N_7942);
and U9438 (N_9438,N_6181,N_8593);
nand U9439 (N_9439,N_8703,N_8189);
nor U9440 (N_9440,N_6490,N_6088);
and U9441 (N_9441,N_8345,N_6071);
nor U9442 (N_9442,N_6153,N_8802);
xor U9443 (N_9443,N_7444,N_6057);
and U9444 (N_9444,N_7367,N_7384);
nand U9445 (N_9445,N_8881,N_7680);
nand U9446 (N_9446,N_8648,N_6500);
nor U9447 (N_9447,N_6294,N_8035);
and U9448 (N_9448,N_6417,N_6907);
or U9449 (N_9449,N_6880,N_7244);
and U9450 (N_9450,N_8014,N_8980);
or U9451 (N_9451,N_8171,N_8394);
nand U9452 (N_9452,N_6654,N_7843);
and U9453 (N_9453,N_8118,N_8395);
nand U9454 (N_9454,N_8552,N_7378);
nand U9455 (N_9455,N_7052,N_7106);
xnor U9456 (N_9456,N_6831,N_6921);
and U9457 (N_9457,N_8390,N_6504);
nand U9458 (N_9458,N_7158,N_7829);
or U9459 (N_9459,N_7214,N_7895);
nor U9460 (N_9460,N_8510,N_8901);
nor U9461 (N_9461,N_8633,N_8961);
nand U9462 (N_9462,N_8022,N_8767);
or U9463 (N_9463,N_8536,N_6176);
nand U9464 (N_9464,N_6144,N_6365);
nand U9465 (N_9465,N_6731,N_8719);
and U9466 (N_9466,N_7635,N_7764);
and U9467 (N_9467,N_6258,N_7308);
and U9468 (N_9468,N_8815,N_7812);
nor U9469 (N_9469,N_6787,N_8490);
xor U9470 (N_9470,N_7243,N_8874);
xnor U9471 (N_9471,N_8175,N_6484);
and U9472 (N_9472,N_7792,N_6596);
or U9473 (N_9473,N_6223,N_6888);
or U9474 (N_9474,N_8410,N_6775);
nand U9475 (N_9475,N_7441,N_6122);
and U9476 (N_9476,N_6442,N_6969);
nor U9477 (N_9477,N_6713,N_8660);
nand U9478 (N_9478,N_6693,N_8602);
and U9479 (N_9479,N_8841,N_6916);
nand U9480 (N_9480,N_7999,N_7760);
nand U9481 (N_9481,N_8324,N_8872);
nand U9482 (N_9482,N_8532,N_7738);
and U9483 (N_9483,N_8211,N_8431);
xor U9484 (N_9484,N_8238,N_7508);
and U9485 (N_9485,N_7195,N_6561);
nor U9486 (N_9486,N_6552,N_8348);
xnor U9487 (N_9487,N_6652,N_6207);
nand U9488 (N_9488,N_6864,N_6584);
or U9489 (N_9489,N_7255,N_6666);
nand U9490 (N_9490,N_6883,N_6818);
or U9491 (N_9491,N_6592,N_6932);
nor U9492 (N_9492,N_8965,N_6948);
xnor U9493 (N_9493,N_6093,N_8461);
or U9494 (N_9494,N_7440,N_8770);
nor U9495 (N_9495,N_6440,N_6454);
and U9496 (N_9496,N_8311,N_8852);
nor U9497 (N_9497,N_6366,N_7674);
nand U9498 (N_9498,N_6606,N_7902);
nand U9499 (N_9499,N_6965,N_8763);
nor U9500 (N_9500,N_7332,N_6464);
nand U9501 (N_9501,N_8731,N_6694);
nand U9502 (N_9502,N_7811,N_8262);
or U9503 (N_9503,N_8315,N_8623);
nor U9504 (N_9504,N_7403,N_8008);
nor U9505 (N_9505,N_6718,N_8645);
nand U9506 (N_9506,N_6009,N_7527);
nand U9507 (N_9507,N_6089,N_8585);
or U9508 (N_9508,N_6096,N_7300);
or U9509 (N_9509,N_7702,N_8275);
and U9510 (N_9510,N_7864,N_8244);
or U9511 (N_9511,N_6133,N_8708);
or U9512 (N_9512,N_6651,N_7141);
nand U9513 (N_9513,N_6983,N_7464);
nand U9514 (N_9514,N_8559,N_8619);
nor U9515 (N_9515,N_6381,N_8317);
nand U9516 (N_9516,N_6509,N_8689);
and U9517 (N_9517,N_6420,N_6957);
nor U9518 (N_9518,N_7688,N_8215);
or U9519 (N_9519,N_7291,N_8287);
and U9520 (N_9520,N_6069,N_7986);
nand U9521 (N_9521,N_6000,N_8592);
xnor U9522 (N_9522,N_8221,N_6276);
xor U9523 (N_9523,N_8666,N_8978);
and U9524 (N_9524,N_6551,N_7209);
nor U9525 (N_9525,N_7632,N_6998);
nor U9526 (N_9526,N_6081,N_8451);
xor U9527 (N_9527,N_7163,N_8644);
or U9528 (N_9528,N_8109,N_7036);
or U9529 (N_9529,N_7469,N_6183);
and U9530 (N_9530,N_8352,N_6720);
nand U9531 (N_9531,N_8846,N_8144);
or U9532 (N_9532,N_8698,N_7821);
xnor U9533 (N_9533,N_8864,N_7656);
and U9534 (N_9534,N_7689,N_8326);
and U9535 (N_9535,N_8668,N_6172);
nand U9536 (N_9536,N_7517,N_6044);
and U9537 (N_9537,N_7142,N_7041);
xnor U9538 (N_9538,N_8962,N_6301);
and U9539 (N_9539,N_7563,N_6319);
nor U9540 (N_9540,N_7139,N_7507);
xor U9541 (N_9541,N_7787,N_6527);
xnor U9542 (N_9542,N_6216,N_8065);
nand U9543 (N_9543,N_7093,N_8309);
nand U9544 (N_9544,N_7271,N_6349);
xnor U9545 (N_9545,N_8347,N_8920);
nor U9546 (N_9546,N_6665,N_8134);
nor U9547 (N_9547,N_8809,N_8321);
nor U9548 (N_9548,N_6986,N_7521);
xnor U9549 (N_9549,N_7087,N_8166);
nor U9550 (N_9550,N_8222,N_7630);
nor U9551 (N_9551,N_7601,N_7500);
xnor U9552 (N_9552,N_6277,N_6570);
xnor U9553 (N_9553,N_8489,N_8759);
nand U9554 (N_9554,N_7515,N_8092);
nor U9555 (N_9555,N_6717,N_6130);
and U9556 (N_9556,N_6394,N_7458);
and U9557 (N_9557,N_8482,N_6160);
nor U9558 (N_9558,N_8756,N_8640);
or U9559 (N_9559,N_7939,N_8172);
nand U9560 (N_9560,N_7002,N_7134);
nand U9561 (N_9561,N_8560,N_7594);
xnor U9562 (N_9562,N_8823,N_8228);
xnor U9563 (N_9563,N_6275,N_8002);
xor U9564 (N_9564,N_6562,N_6444);
or U9565 (N_9565,N_7405,N_8044);
and U9566 (N_9566,N_7103,N_6641);
and U9567 (N_9567,N_6061,N_8601);
xor U9568 (N_9568,N_8968,N_8102);
or U9569 (N_9569,N_8733,N_8549);
or U9570 (N_9570,N_8739,N_8029);
nand U9571 (N_9571,N_7380,N_6853);
nand U9572 (N_9572,N_6909,N_6269);
or U9573 (N_9573,N_6244,N_6152);
xnor U9574 (N_9574,N_8916,N_8669);
and U9575 (N_9575,N_8219,N_8279);
xor U9576 (N_9576,N_7396,N_6221);
nor U9577 (N_9577,N_6035,N_6491);
nand U9578 (N_9578,N_8110,N_8241);
xnor U9579 (N_9579,N_7712,N_8435);
and U9580 (N_9580,N_7220,N_8654);
and U9581 (N_9581,N_7875,N_6817);
or U9582 (N_9582,N_6241,N_7566);
nand U9583 (N_9583,N_7834,N_6507);
and U9584 (N_9584,N_7438,N_8579);
nand U9585 (N_9585,N_7578,N_6402);
and U9586 (N_9586,N_7894,N_8203);
or U9587 (N_9587,N_7481,N_6926);
nor U9588 (N_9588,N_6157,N_8325);
nor U9589 (N_9589,N_8261,N_7436);
nor U9590 (N_9590,N_8626,N_8911);
nand U9591 (N_9591,N_8495,N_8604);
nor U9592 (N_9592,N_7022,N_8151);
xor U9593 (N_9593,N_7208,N_6803);
xnor U9594 (N_9594,N_8125,N_6898);
nor U9595 (N_9595,N_6999,N_7415);
xor U9596 (N_9596,N_8304,N_6282);
or U9597 (N_9597,N_8313,N_8448);
nor U9598 (N_9598,N_7782,N_8891);
nand U9599 (N_9599,N_6430,N_6966);
nand U9600 (N_9600,N_6586,N_8857);
or U9601 (N_9601,N_6287,N_8967);
nor U9602 (N_9602,N_7176,N_8282);
nand U9603 (N_9603,N_6456,N_7144);
nand U9604 (N_9604,N_7312,N_8984);
xor U9605 (N_9605,N_8301,N_8970);
and U9606 (N_9606,N_8135,N_8485);
or U9607 (N_9607,N_6102,N_7355);
nand U9608 (N_9608,N_7248,N_6228);
and U9609 (N_9609,N_7013,N_7452);
nand U9610 (N_9610,N_8652,N_8302);
or U9611 (N_9611,N_7143,N_7240);
or U9612 (N_9612,N_6816,N_6742);
or U9613 (N_9613,N_6832,N_8398);
nand U9614 (N_9614,N_7091,N_7096);
and U9615 (N_9615,N_7800,N_8055);
and U9616 (N_9616,N_7972,N_8964);
and U9617 (N_9617,N_7643,N_6753);
xor U9618 (N_9618,N_6126,N_7779);
and U9619 (N_9619,N_6648,N_6483);
xor U9620 (N_9620,N_6450,N_7329);
and U9621 (N_9621,N_8934,N_7772);
xnor U9622 (N_9622,N_8187,N_8075);
xnor U9623 (N_9623,N_7650,N_7073);
nor U9624 (N_9624,N_7988,N_6327);
nand U9625 (N_9625,N_7302,N_7120);
xnor U9626 (N_9626,N_8875,N_8101);
xor U9627 (N_9627,N_8277,N_6746);
or U9628 (N_9628,N_7351,N_6125);
or U9629 (N_9629,N_6168,N_6623);
and U9630 (N_9630,N_8785,N_8993);
and U9631 (N_9631,N_6739,N_7362);
or U9632 (N_9632,N_6309,N_8673);
nand U9633 (N_9633,N_7793,N_6852);
or U9634 (N_9634,N_8839,N_7127);
and U9635 (N_9635,N_8915,N_6875);
or U9636 (N_9636,N_8123,N_7294);
nor U9637 (N_9637,N_7230,N_8550);
or U9638 (N_9638,N_6421,N_7370);
xor U9639 (N_9639,N_7222,N_7849);
nor U9640 (N_9640,N_7418,N_6002);
nor U9641 (N_9641,N_6600,N_7281);
or U9642 (N_9642,N_6446,N_8367);
and U9643 (N_9643,N_6378,N_6886);
nand U9644 (N_9644,N_6184,N_7876);
or U9645 (N_9645,N_8019,N_7038);
or U9646 (N_9646,N_8621,N_7645);
nor U9647 (N_9647,N_8555,N_8840);
nor U9648 (N_9648,N_6789,N_7343);
xor U9649 (N_9649,N_8505,N_7077);
and U9650 (N_9650,N_7320,N_8477);
or U9651 (N_9651,N_8403,N_7615);
nor U9652 (N_9652,N_6846,N_8826);
nand U9653 (N_9653,N_6566,N_7421);
nand U9654 (N_9654,N_8562,N_7258);
or U9655 (N_9655,N_6796,N_8440);
or U9656 (N_9656,N_8863,N_8699);
or U9657 (N_9657,N_7328,N_6612);
xnor U9658 (N_9658,N_8582,N_7526);
nor U9659 (N_9659,N_7828,N_6695);
nor U9660 (N_9660,N_8971,N_8804);
nor U9661 (N_9661,N_8369,N_8436);
and U9662 (N_9662,N_6302,N_7701);
nand U9663 (N_9663,N_8331,N_8243);
xor U9664 (N_9664,N_7497,N_8411);
xor U9665 (N_9665,N_6531,N_7668);
nand U9666 (N_9666,N_8429,N_7357);
nor U9667 (N_9667,N_8568,N_7261);
xnor U9668 (N_9668,N_6530,N_7373);
xor U9669 (N_9669,N_8488,N_7025);
and U9670 (N_9670,N_8200,N_7614);
xor U9671 (N_9671,N_6544,N_7413);
nor U9672 (N_9672,N_6861,N_6107);
nand U9673 (N_9673,N_7684,N_6704);
and U9674 (N_9674,N_8778,N_7268);
nand U9675 (N_9675,N_6628,N_8704);
xnor U9676 (N_9676,N_6857,N_8434);
nand U9677 (N_9677,N_6210,N_6213);
nand U9678 (N_9678,N_6741,N_8506);
nor U9679 (N_9679,N_8148,N_6847);
or U9680 (N_9680,N_6240,N_7626);
nand U9681 (N_9681,N_8992,N_7685);
nand U9682 (N_9682,N_8473,N_8524);
or U9683 (N_9683,N_8912,N_6053);
nand U9684 (N_9684,N_7613,N_8353);
nor U9685 (N_9685,N_8146,N_8307);
or U9686 (N_9686,N_6565,N_8328);
xnor U9687 (N_9687,N_6748,N_7815);
nand U9688 (N_9688,N_8764,N_6608);
xor U9689 (N_9689,N_7303,N_6997);
nor U9690 (N_9690,N_7231,N_6268);
xor U9691 (N_9691,N_7428,N_7100);
or U9692 (N_9692,N_6918,N_7055);
or U9693 (N_9693,N_8064,N_6873);
nand U9694 (N_9694,N_7033,N_7713);
nand U9695 (N_9695,N_7092,N_6781);
xnor U9696 (N_9696,N_8859,N_6963);
and U9697 (N_9697,N_7053,N_6613);
or U9698 (N_9698,N_8205,N_6322);
xor U9699 (N_9699,N_8609,N_6664);
nor U9700 (N_9700,N_8122,N_7155);
or U9701 (N_9701,N_7550,N_7791);
nor U9702 (N_9702,N_6679,N_8825);
nand U9703 (N_9703,N_7962,N_6959);
nor U9704 (N_9704,N_8480,N_6599);
and U9705 (N_9705,N_6175,N_6823);
nor U9706 (N_9706,N_7516,N_8085);
and U9707 (N_9707,N_7298,N_7181);
and U9708 (N_9708,N_6611,N_7260);
or U9709 (N_9709,N_6701,N_8670);
xnor U9710 (N_9710,N_7472,N_6360);
or U9711 (N_9711,N_8672,N_6026);
or U9712 (N_9712,N_6250,N_8563);
and U9713 (N_9713,N_7221,N_7710);
or U9714 (N_9714,N_8950,N_7388);
or U9715 (N_9715,N_8285,N_7531);
nand U9716 (N_9716,N_8212,N_7188);
and U9717 (N_9717,N_7024,N_6041);
nand U9718 (N_9718,N_8716,N_7784);
xnor U9719 (N_9719,N_8771,N_7575);
xnor U9720 (N_9720,N_6855,N_8746);
xor U9721 (N_9721,N_8364,N_7679);
and U9722 (N_9722,N_8363,N_8695);
or U9723 (N_9723,N_8033,N_8845);
and U9724 (N_9724,N_7709,N_8960);
and U9725 (N_9725,N_8152,N_8018);
or U9726 (N_9726,N_6127,N_7768);
or U9727 (N_9727,N_6513,N_8812);
nor U9728 (N_9728,N_8958,N_8973);
nor U9729 (N_9729,N_6630,N_8757);
xnor U9730 (N_9730,N_8547,N_8433);
nand U9731 (N_9731,N_7097,N_7961);
nand U9732 (N_9732,N_7259,N_6194);
nor U9733 (N_9733,N_7353,N_7167);
or U9734 (N_9734,N_7907,N_8124);
xor U9735 (N_9735,N_7321,N_7799);
and U9736 (N_9736,N_8943,N_6749);
or U9737 (N_9737,N_8167,N_6528);
or U9738 (N_9738,N_8832,N_6506);
or U9739 (N_9739,N_8529,N_8414);
nor U9740 (N_9740,N_8486,N_8133);
nand U9741 (N_9741,N_6700,N_6943);
xor U9742 (N_9742,N_6048,N_7858);
nor U9743 (N_9743,N_7145,N_7473);
nor U9744 (N_9744,N_6970,N_7562);
nand U9745 (N_9745,N_6906,N_8700);
and U9746 (N_9746,N_7133,N_7211);
nor U9747 (N_9747,N_7404,N_6868);
xor U9748 (N_9748,N_8897,N_6979);
nor U9749 (N_9749,N_7275,N_8817);
nand U9750 (N_9750,N_6441,N_8341);
xnor U9751 (N_9751,N_8798,N_6571);
nand U9752 (N_9752,N_7172,N_6050);
xor U9753 (N_9753,N_7687,N_8811);
xor U9754 (N_9754,N_8807,N_8174);
and U9755 (N_9755,N_8938,N_8366);
xnor U9756 (N_9756,N_7242,N_6845);
nand U9757 (N_9757,N_8471,N_8028);
and U9758 (N_9758,N_6964,N_7194);
nand U9759 (N_9759,N_8329,N_8009);
and U9760 (N_9760,N_7218,N_8103);
xnor U9761 (N_9761,N_7417,N_7490);
nor U9762 (N_9762,N_6636,N_7317);
and U9763 (N_9763,N_7045,N_7582);
nor U9764 (N_9764,N_7842,N_7987);
nor U9765 (N_9765,N_7773,N_6896);
and U9766 (N_9766,N_6414,N_7719);
nor U9767 (N_9767,N_6156,N_6187);
or U9768 (N_9768,N_7788,N_7996);
and U9769 (N_9769,N_7542,N_7510);
or U9770 (N_9770,N_7732,N_6525);
nand U9771 (N_9771,N_7207,N_8908);
or U9772 (N_9772,N_6150,N_6111);
or U9773 (N_9773,N_6827,N_8508);
xnor U9774 (N_9774,N_7225,N_6054);
nand U9775 (N_9775,N_8906,N_8068);
xor U9776 (N_9776,N_7745,N_7090);
and U9777 (N_9777,N_7493,N_8438);
xnor U9778 (N_9778,N_7965,N_7756);
or U9779 (N_9779,N_8821,N_7044);
or U9780 (N_9780,N_7111,N_6549);
or U9781 (N_9781,N_7862,N_8442);
nor U9782 (N_9782,N_7338,N_8358);
xnor U9783 (N_9783,N_8416,N_8646);
and U9784 (N_9784,N_8381,N_6092);
nand U9785 (N_9785,N_6474,N_8242);
xnor U9786 (N_9786,N_8781,N_8534);
and U9787 (N_9787,N_6034,N_8545);
nor U9788 (N_9788,N_8306,N_7138);
or U9789 (N_9789,N_7636,N_8907);
xor U9790 (N_9790,N_8713,N_6182);
xor U9791 (N_9791,N_6290,N_6449);
and U9792 (N_9792,N_7881,N_8573);
nand U9793 (N_9793,N_7586,N_8063);
nor U9794 (N_9794,N_7019,N_8034);
nor U9795 (N_9795,N_6934,N_7836);
xor U9796 (N_9796,N_6324,N_8493);
and U9797 (N_9797,N_7330,N_7623);
and U9798 (N_9798,N_7079,N_8157);
xnor U9799 (N_9799,N_6655,N_7223);
or U9800 (N_9800,N_7016,N_8412);
or U9801 (N_9801,N_8456,N_7182);
and U9802 (N_9802,N_7029,N_8693);
and U9803 (N_9803,N_7599,N_8492);
nor U9804 (N_9804,N_7442,N_8382);
nor U9805 (N_9805,N_6097,N_7584);
nor U9806 (N_9806,N_8661,N_7288);
or U9807 (N_9807,N_8376,N_8349);
nor U9808 (N_9808,N_6499,N_7264);
or U9809 (N_9809,N_6870,N_8297);
nand U9810 (N_9810,N_7638,N_6927);
and U9811 (N_9811,N_7265,N_8790);
nand U9812 (N_9812,N_7927,N_8949);
or U9813 (N_9813,N_6351,N_8761);
and U9814 (N_9814,N_6475,N_6205);
and U9815 (N_9815,N_6332,N_8914);
or U9816 (N_9816,N_8387,N_6476);
nor U9817 (N_9817,N_6669,N_6850);
nor U9818 (N_9818,N_6426,N_6660);
nand U9819 (N_9819,N_6356,N_8880);
xor U9820 (N_9820,N_6015,N_7371);
and U9821 (N_9821,N_7588,N_6162);
or U9822 (N_9822,N_8930,N_8032);
nor U9823 (N_9823,N_6331,N_6436);
or U9824 (N_9824,N_6558,N_6696);
or U9825 (N_9825,N_8883,N_7354);
xnor U9826 (N_9826,N_8856,N_7769);
or U9827 (N_9827,N_8450,N_7917);
or U9828 (N_9828,N_6292,N_8948);
and U9829 (N_9829,N_6224,N_6547);
xor U9830 (N_9830,N_6283,N_7744);
or U9831 (N_9831,N_7459,N_8089);
xor U9832 (N_9832,N_6139,N_8079);
nand U9833 (N_9833,N_6572,N_7558);
nand U9834 (N_9834,N_6030,N_6769);
and U9835 (N_9835,N_8999,N_8047);
xnor U9836 (N_9836,N_7060,N_7035);
nor U9837 (N_9837,N_6894,N_7911);
or U9838 (N_9838,N_8753,N_6338);
nand U9839 (N_9839,N_7621,N_6108);
nand U9840 (N_9840,N_6914,N_8614);
and U9841 (N_9841,N_7589,N_7174);
or U9842 (N_9842,N_8540,N_8744);
xor U9843 (N_9843,N_7564,N_8388);
nor U9844 (N_9844,N_7971,N_7579);
nand U9845 (N_9845,N_6313,N_8849);
and U9846 (N_9846,N_6101,N_6200);
nor U9847 (N_9847,N_7754,N_7619);
nand U9848 (N_9848,N_6487,N_7478);
or U9849 (N_9849,N_6232,N_8502);
xnor U9850 (N_9850,N_8040,N_6594);
or U9851 (N_9851,N_8792,N_8909);
nor U9852 (N_9852,N_7877,N_8600);
and U9853 (N_9853,N_7923,N_7819);
nand U9854 (N_9854,N_6772,N_7976);
or U9855 (N_9855,N_8337,N_8308);
and U9856 (N_9856,N_6618,N_6807);
and U9857 (N_9857,N_6415,N_7198);
xor U9858 (N_9858,N_8683,N_6967);
or U9859 (N_9859,N_8472,N_6622);
nand U9860 (N_9860,N_7683,N_8226);
or U9861 (N_9861,N_7250,N_7094);
and U9862 (N_9862,N_7169,N_6869);
nand U9863 (N_9863,N_7131,N_6234);
nand U9864 (N_9864,N_8541,N_7734);
nor U9865 (N_9865,N_8007,N_7723);
nand U9866 (N_9866,N_6685,N_7539);
or U9867 (N_9867,N_8207,N_6837);
nand U9868 (N_9868,N_7631,N_6123);
and U9869 (N_9869,N_8653,N_7968);
nor U9870 (N_9870,N_7752,N_6289);
and U9871 (N_9871,N_8178,N_8622);
nand U9872 (N_9872,N_7786,N_7660);
nor U9873 (N_9873,N_7816,N_6913);
nor U9874 (N_9874,N_8137,N_8048);
nand U9875 (N_9875,N_6068,N_7400);
nand U9876 (N_9876,N_6055,N_8813);
xnor U9877 (N_9877,N_7267,N_8824);
and U9878 (N_9878,N_6830,N_8129);
or U9879 (N_9879,N_8479,N_7757);
nand U9880 (N_9880,N_7642,N_7184);
nand U9881 (N_9881,N_7499,N_8111);
and U9882 (N_9882,N_8312,N_8463);
and U9883 (N_9883,N_7950,N_8402);
or U9884 (N_9884,N_6266,N_8155);
and U9885 (N_9885,N_6564,N_6073);
nor U9886 (N_9886,N_8156,N_8276);
nand U9887 (N_9887,N_6227,N_8227);
xor U9888 (N_9888,N_7585,N_8500);
xnor U9889 (N_9889,N_6935,N_7720);
nand U9890 (N_9890,N_6398,N_8491);
xor U9891 (N_9891,N_7706,N_8898);
or U9892 (N_9892,N_8181,N_6121);
xnor U9893 (N_9893,N_7686,N_7893);
nor U9894 (N_9894,N_8990,N_7385);
nor U9895 (N_9895,N_8869,N_7252);
xnor U9896 (N_9896,N_6863,N_7000);
xor U9897 (N_9897,N_6919,N_6052);
nor U9898 (N_9898,N_8997,N_8977);
or U9899 (N_9899,N_7043,N_6825);
nor U9900 (N_9900,N_7387,N_6249);
and U9901 (N_9901,N_6011,N_7196);
and U9902 (N_9902,N_7899,N_7477);
xor U9903 (N_9903,N_8000,N_7749);
nand U9904 (N_9904,N_8905,N_6750);
nand U9905 (N_9905,N_7629,N_7808);
nand U9906 (N_9906,N_6477,N_6573);
nand U9907 (N_9907,N_6901,N_7915);
xnor U9908 (N_9908,N_6344,N_8886);
and U9909 (N_9909,N_7966,N_6263);
and U9910 (N_9910,N_8100,N_7423);
xnor U9911 (N_9911,N_6834,N_7032);
nor U9912 (N_9912,N_6686,N_6732);
nor U9913 (N_9913,N_6676,N_6503);
nand U9914 (N_9914,N_6297,N_8789);
nor U9915 (N_9915,N_7479,N_6649);
xnor U9916 (N_9916,N_8998,N_7050);
nand U9917 (N_9917,N_7967,N_7627);
or U9918 (N_9918,N_6005,N_7669);
nor U9919 (N_9919,N_6120,N_8512);
nand U9920 (N_9920,N_8574,N_6545);
or U9921 (N_9921,N_8774,N_7057);
or U9922 (N_9922,N_7886,N_7854);
nor U9923 (N_9923,N_7543,N_6619);
nor U9924 (N_9924,N_8015,N_6132);
or U9925 (N_9925,N_6403,N_8260);
and U9926 (N_9926,N_8097,N_8446);
or U9927 (N_9927,N_6842,N_7700);
xor U9928 (N_9928,N_7775,N_7724);
nor U9929 (N_9929,N_6771,N_7206);
xor U9930 (N_9930,N_8095,N_6076);
nor U9931 (N_9931,N_8284,N_7277);
xor U9932 (N_9932,N_7771,N_8081);
and U9933 (N_9933,N_7556,N_6273);
or U9934 (N_9934,N_6627,N_6341);
xnor U9935 (N_9935,N_6738,N_8054);
or U9936 (N_9936,N_8724,N_6208);
nand U9937 (N_9937,N_7164,N_8444);
xor U9938 (N_9938,N_7109,N_8254);
xor U9939 (N_9939,N_7861,N_7783);
and U9940 (N_9940,N_8235,N_6682);
nor U9941 (N_9941,N_8983,N_7780);
or U9942 (N_9942,N_7890,N_8854);
nor U9943 (N_9943,N_6451,N_8836);
and U9944 (N_9944,N_8658,N_6778);
nand U9945 (N_9945,N_7216,N_6579);
xnor U9946 (N_9946,N_7224,N_7831);
nand U9947 (N_9947,N_8419,N_8899);
and U9948 (N_9948,N_7339,N_6763);
nand U9949 (N_9949,N_8544,N_7644);
nand U9950 (N_9950,N_6508,N_6675);
and U9951 (N_9951,N_7072,N_6899);
nand U9952 (N_9952,N_7901,N_6281);
nor U9953 (N_9953,N_6687,N_7424);
nor U9954 (N_9954,N_7189,N_6889);
and U9955 (N_9955,N_8705,N_6084);
nor U9956 (N_9956,N_7058,N_8105);
or U9957 (N_9957,N_6674,N_7739);
and U9958 (N_9958,N_8206,N_8808);
nor U9959 (N_9959,N_8586,N_7557);
xor U9960 (N_9960,N_6128,N_8656);
or U9961 (N_9961,N_7039,N_8120);
nor U9962 (N_9962,N_6495,N_6178);
xnor U9963 (N_9963,N_6317,N_8458);
nor U9964 (N_9964,N_7495,N_6642);
and U9965 (N_9965,N_8928,N_6582);
xor U9966 (N_9966,N_7646,N_8086);
or U9967 (N_9967,N_7676,N_6246);
and U9968 (N_9968,N_8107,N_8272);
nand U9969 (N_9969,N_8922,N_6267);
and U9970 (N_9970,N_6377,N_7397);
or U9971 (N_9971,N_6604,N_6924);
xor U9972 (N_9972,N_6251,N_8026);
xnor U9973 (N_9973,N_6214,N_8043);
nand U9974 (N_9974,N_8383,N_6995);
and U9975 (N_9975,N_6820,N_7340);
nand U9976 (N_9976,N_8996,N_7838);
or U9977 (N_9977,N_6780,N_7634);
nor U9978 (N_9978,N_7565,N_6632);
or U9979 (N_9979,N_6264,N_6735);
and U9980 (N_9980,N_7935,N_6063);
xnor U9981 (N_9981,N_6574,N_7070);
or U9982 (N_9982,N_8932,N_6439);
or U9983 (N_9983,N_7290,N_8333);
or U9984 (N_9984,N_6569,N_7762);
nand U9985 (N_9985,N_7616,N_7247);
or U9986 (N_9986,N_6708,N_8210);
nand U9987 (N_9987,N_6953,N_6971);
xnor U9988 (N_9988,N_7374,N_6759);
and U9989 (N_9989,N_7487,N_6237);
nor U9990 (N_9990,N_7984,N_6329);
nor U9991 (N_9991,N_6288,N_8396);
or U9992 (N_9992,N_7372,N_7249);
or U9993 (N_9993,N_7228,N_7576);
nand U9994 (N_9994,N_6520,N_7241);
nand U9995 (N_9995,N_7909,N_6370);
nor U9996 (N_9996,N_7006,N_6534);
or U9997 (N_9997,N_7781,N_8871);
nand U9998 (N_9998,N_8299,N_7912);
nand U9999 (N_9999,N_6991,N_8386);
nand U10000 (N_10000,N_6867,N_8230);
nor U10001 (N_10001,N_8036,N_7920);
nand U10002 (N_10002,N_8717,N_7874);
nor U10003 (N_10003,N_6946,N_6031);
and U10004 (N_10004,N_7349,N_7536);
nor U10005 (N_10005,N_7313,N_7677);
or U10006 (N_10006,N_8264,N_7324);
nand U10007 (N_10007,N_8945,N_7525);
xnor U10008 (N_10008,N_8011,N_7467);
or U10009 (N_10009,N_7197,N_7652);
xnor U10010 (N_10010,N_8636,N_8090);
nor U10011 (N_10011,N_8750,N_7274);
nor U10012 (N_10012,N_7839,N_6895);
nor U10013 (N_10013,N_7552,N_7280);
and U10014 (N_10014,N_7005,N_6099);
nand U10015 (N_10015,N_6653,N_8749);
nor U10016 (N_10016,N_8665,N_7146);
nand U10017 (N_10017,N_8359,N_7970);
xnor U10018 (N_10018,N_7076,N_7123);
nand U10019 (N_10019,N_6471,N_8850);
and U10020 (N_10020,N_8953,N_7954);
and U10021 (N_10021,N_7540,N_7369);
and U10022 (N_10022,N_8929,N_8740);
and U10023 (N_10023,N_6678,N_6872);
nor U10024 (N_10024,N_7830,N_8548);
and U10025 (N_10025,N_8127,N_6204);
and U10026 (N_10026,N_6056,N_8796);
nor U10027 (N_10027,N_7014,N_8972);
or U10028 (N_10028,N_6100,N_7010);
and U10029 (N_10029,N_8879,N_8257);
xnor U10030 (N_10030,N_6489,N_6524);
and U10031 (N_10031,N_6758,N_8926);
nor U10032 (N_10032,N_8224,N_6468);
or U10033 (N_10033,N_7620,N_6878);
nor U10034 (N_10034,N_7345,N_8725);
or U10035 (N_10035,N_7245,N_6429);
nor U10036 (N_10036,N_7137,N_8692);
and U10037 (N_10037,N_8736,N_7480);
and U10038 (N_10038,N_6098,N_8531);
or U10039 (N_10039,N_8685,N_8422);
and U10040 (N_10040,N_6773,N_6452);
xnor U10041 (N_10041,N_8459,N_6923);
nor U10042 (N_10042,N_8117,N_8439);
or U10043 (N_10043,N_6517,N_6386);
xor U10044 (N_10044,N_6091,N_7866);
nor U10045 (N_10045,N_6539,N_8050);
xnor U10046 (N_10046,N_7190,N_8375);
nand U10047 (N_10047,N_6384,N_7433);
nor U10048 (N_10048,N_6272,N_6412);
or U10049 (N_10049,N_6515,N_8062);
xnor U10050 (N_10050,N_6659,N_7670);
and U10051 (N_10051,N_8096,N_6300);
and U10052 (N_10052,N_6848,N_7150);
xnor U10053 (N_10053,N_6007,N_7804);
or U10054 (N_10054,N_6529,N_7814);
xor U10055 (N_10055,N_7889,N_7179);
and U10056 (N_10056,N_7462,N_6721);
nand U10057 (N_10057,N_7598,N_8853);
or U10058 (N_10058,N_7600,N_8639);
or U10059 (N_10059,N_6973,N_6587);
and U10060 (N_10060,N_7736,N_7735);
nor U10061 (N_10061,N_8882,N_6585);
or U10062 (N_10062,N_6453,N_8613);
or U10063 (N_10063,N_8618,N_8216);
xor U10064 (N_10064,N_6409,N_8775);
nor U10065 (N_10065,N_8149,N_6077);
nand U10066 (N_10066,N_7402,N_8074);
xnor U10067 (N_10067,N_6790,N_8686);
xor U10068 (N_10068,N_8368,N_8320);
and U10069 (N_10069,N_8721,N_6580);
nor U10070 (N_10070,N_6858,N_6621);
nand U10071 (N_10071,N_7870,N_7959);
nand U10072 (N_10072,N_7099,N_6373);
xnor U10073 (N_10073,N_7322,N_8710);
nor U10074 (N_10074,N_8737,N_7767);
and U10075 (N_10075,N_7711,N_8342);
and U10076 (N_10076,N_6318,N_8392);
nor U10077 (N_10077,N_7654,N_6364);
xor U10078 (N_10078,N_7140,N_7278);
nor U10079 (N_10079,N_6253,N_6601);
xor U10080 (N_10080,N_7416,N_6470);
nand U10081 (N_10081,N_8829,N_7037);
and U10082 (N_10082,N_7766,N_7580);
or U10083 (N_10083,N_6148,N_8954);
xor U10084 (N_10084,N_6822,N_8391);
or U10085 (N_10085,N_8365,N_8659);
and U10086 (N_10086,N_8590,N_7069);
or U10087 (N_10087,N_8711,N_6201);
and U10088 (N_10088,N_7606,N_7386);
nand U10089 (N_10089,N_7704,N_7618);
nor U10090 (N_10090,N_8603,N_8190);
and U10091 (N_10091,N_7647,N_6879);
or U10092 (N_10092,N_7969,N_8726);
and U10093 (N_10093,N_8889,N_7617);
nor U10094 (N_10094,N_6908,N_7802);
and U10095 (N_10095,N_8913,N_6085);
and U10096 (N_10096,N_7975,N_8591);
xor U10097 (N_10097,N_6798,N_8738);
nand U10098 (N_10098,N_7990,N_6952);
nor U10099 (N_10099,N_6866,N_6472);
nand U10100 (N_10100,N_6663,N_8322);
nor U10101 (N_10101,N_6634,N_7649);
and U10102 (N_10102,N_6112,N_6994);
or U10103 (N_10103,N_6805,N_8183);
nand U10104 (N_10104,N_7148,N_8921);
nand U10105 (N_10105,N_6371,N_7682);
xnor U10106 (N_10106,N_7880,N_6218);
or U10107 (N_10107,N_8130,N_6777);
nor U10108 (N_10108,N_7730,N_8981);
and U10109 (N_10109,N_7625,N_8250);
nand U10110 (N_10110,N_6154,N_6037);
nor U10111 (N_10111,N_7301,N_7496);
and U10112 (N_10112,N_6813,N_7286);
and U10113 (N_10113,N_6640,N_6559);
or U10114 (N_10114,N_8772,N_7295);
and U10115 (N_10115,N_7648,N_7581);
xor U10116 (N_10116,N_7777,N_6087);
or U10117 (N_10117,N_8001,N_8745);
nand U10118 (N_10118,N_8919,N_7307);
and U10119 (N_10119,N_7774,N_7763);
nand U10120 (N_10120,N_8204,N_6142);
and U10121 (N_10121,N_6347,N_6359);
nor U10122 (N_10122,N_7798,N_6762);
nand U10123 (N_10123,N_6065,N_6025);
nor U10124 (N_10124,N_6385,N_6177);
xnor U10125 (N_10125,N_6751,N_7559);
nand U10126 (N_10126,N_8318,N_6765);
xor U10127 (N_10127,N_6438,N_8935);
nor U10128 (N_10128,N_7341,N_7590);
nand U10129 (N_10129,N_6794,N_7930);
xor U10130 (N_10130,N_8202,N_7717);
xor U10131 (N_10131,N_8087,N_6745);
and U10132 (N_10132,N_6345,N_6978);
xor U10133 (N_10133,N_8098,N_8378);
xor U10134 (N_10134,N_8776,N_7088);
or U10135 (N_10135,N_6119,N_7825);
nand U10136 (N_10136,N_8542,N_6684);
nand U10137 (N_10137,N_8571,N_6134);
and U10138 (N_10138,N_8924,N_7722);
nor U10139 (N_10139,N_8554,N_8873);
nor U10140 (N_10140,N_8734,N_7453);
or U10141 (N_10141,N_8373,N_6939);
nor U10142 (N_10142,N_8194,N_7919);
or U10143 (N_10143,N_6335,N_6638);
nand U10144 (N_10144,N_6236,N_8344);
nor U10145 (N_10145,N_8664,N_6411);
xor U10146 (N_10146,N_6815,N_6975);
xor U10147 (N_10147,N_7943,N_8377);
and U10148 (N_10148,N_8217,N_8748);
or U10149 (N_10149,N_8513,N_6968);
nand U10150 (N_10150,N_7319,N_8432);
and U10151 (N_10151,N_7293,N_6382);
xnor U10152 (N_10152,N_8024,N_7001);
and U10153 (N_10153,N_8393,N_8709);
nor U10154 (N_10154,N_6304,N_6785);
or U10155 (N_10155,N_8165,N_7776);
nor U10156 (N_10156,N_8580,N_7200);
nor U10157 (N_10157,N_8354,N_6808);
nand U10158 (N_10158,N_8773,N_8269);
or U10159 (N_10159,N_8715,N_8876);
nor U10160 (N_10160,N_8220,N_8409);
or U10161 (N_10161,N_7285,N_8732);
nor U10162 (N_10162,N_6938,N_7483);
nand U10163 (N_10163,N_6467,N_8300);
or U10164 (N_10164,N_8939,N_6960);
or U10165 (N_10165,N_7159,N_6362);
xnor U10166 (N_10166,N_8688,N_8292);
or U10167 (N_10167,N_7287,N_6167);
nand U10168 (N_10168,N_6992,N_7409);
xor U10169 (N_10169,N_6783,N_8820);
and U10170 (N_10170,N_7883,N_6116);
xnor U10171 (N_10171,N_7432,N_7751);
or U10172 (N_10172,N_6620,N_8687);
nand U10173 (N_10173,N_6797,N_8543);
nand U10174 (N_10174,N_8931,N_8399);
and U10175 (N_10175,N_7398,N_6311);
and U10176 (N_10176,N_8523,N_6256);
nor U10177 (N_10177,N_6904,N_7186);
xnor U10178 (N_10178,N_7040,N_6800);
and U10179 (N_10179,N_7136,N_7326);
and U10180 (N_10180,N_6854,N_7316);
xnor U10181 (N_10181,N_7639,N_7049);
or U10182 (N_10182,N_6578,N_6768);
nor U10183 (N_10183,N_6493,N_8417);
nand U10184 (N_10184,N_7520,N_8595);
nor U10185 (N_10185,N_8567,N_6590);
and U10186 (N_10186,N_6339,N_6812);
or U10187 (N_10187,N_8106,N_7460);
and U10188 (N_10188,N_7859,N_8777);
xnor U10189 (N_10189,N_8955,N_6140);
nand U10190 (N_10190,N_6286,N_6079);
xnor U10191 (N_10191,N_6180,N_7803);
xor U10192 (N_10192,N_7128,N_6633);
and U10193 (N_10193,N_6667,N_7885);
xor U10194 (N_10194,N_8140,N_6719);
and U10195 (N_10195,N_7314,N_7334);
nor U10196 (N_10196,N_6523,N_6951);
or U10197 (N_10197,N_7017,N_8743);
and U10198 (N_10198,N_6298,N_7957);
xnor U10199 (N_10199,N_7981,N_6501);
xor U10200 (N_10200,N_6067,N_6828);
and U10201 (N_10201,N_8810,N_6391);
nand U10202 (N_10202,N_6518,N_6835);
nand U10203 (N_10203,N_6643,N_7066);
nor U10204 (N_10204,N_7210,N_6728);
or U10205 (N_10205,N_6890,N_6577);
xor U10206 (N_10206,N_8108,N_7873);
or U10207 (N_10207,N_8334,N_7107);
and U10208 (N_10208,N_6186,N_6136);
and U10209 (N_10209,N_7918,N_6461);
nor U10210 (N_10210,N_6252,N_8584);
and U10211 (N_10211,N_8518,N_8637);
xor U10212 (N_10212,N_7822,N_6546);
xnor U10213 (N_10213,N_7251,N_7394);
nand U10214 (N_10214,N_7778,N_7333);
nor U10215 (N_10215,N_8558,N_8158);
xor U10216 (N_10216,N_6375,N_7082);
nor U10217 (N_10217,N_8910,N_8356);
and U10218 (N_10218,N_8768,N_6372);
or U10219 (N_10219,N_7125,N_7130);
nand U10220 (N_10220,N_8515,N_8903);
nor U10221 (N_10221,N_7124,N_7482);
xnor U10222 (N_10222,N_8615,N_6802);
nand U10223 (N_10223,N_8765,N_7283);
nor U10224 (N_10224,N_7310,N_6278);
or U10225 (N_10225,N_7160,N_7845);
nor U10226 (N_10226,N_8293,N_7256);
and U10227 (N_10227,N_7568,N_8769);
and U10228 (N_10228,N_8788,N_8578);
nand U10229 (N_10229,N_6860,N_6647);
xnor U10230 (N_10230,N_7315,N_6554);
xor U10231 (N_10231,N_8594,N_7852);
and U10232 (N_10232,N_7867,N_7925);
nor U10233 (N_10233,N_8702,N_8161);
and U10234 (N_10234,N_8208,N_6548);
or U10235 (N_10235,N_8114,N_8497);
or U10236 (N_10236,N_6972,N_6736);
xor U10237 (N_10237,N_8169,N_8900);
and U10238 (N_10238,N_8371,N_6379);
nand U10239 (N_10239,N_7129,N_8332);
nand U10240 (N_10240,N_7476,N_6308);
nor U10241 (N_10241,N_7470,N_7456);
and U10242 (N_10242,N_7535,N_6019);
nand U10243 (N_10243,N_7414,N_8073);
nand U10244 (N_10244,N_7171,N_8453);
nor U10245 (N_10245,N_6788,N_8729);
nand U10246 (N_10246,N_7135,N_7960);
nand U10247 (N_10247,N_7662,N_7086);
nand U10248 (N_10248,N_6202,N_6045);
xnor U10249 (N_10249,N_8751,N_8153);
nor U10250 (N_10250,N_7116,N_6219);
xnor U10251 (N_10251,N_8521,N_6314);
nor U10252 (N_10252,N_6291,N_6716);
nor U10253 (N_10253,N_8800,N_7603);
and U10254 (N_10254,N_7311,N_7847);
nor U10255 (N_10255,N_7383,N_7665);
xor U10256 (N_10256,N_6744,N_8561);
nor U10257 (N_10257,N_7519,N_7364);
and U10258 (N_10258,N_7952,N_6699);
xor U10259 (N_10259,N_6303,N_8066);
nor U10260 (N_10260,N_7439,N_8267);
or U10261 (N_10261,N_6481,N_6603);
nor U10262 (N_10262,N_6238,N_6104);
and U10263 (N_10263,N_6910,N_7554);
nor U10264 (N_10264,N_6480,N_8522);
and U10265 (N_10265,N_6040,N_8520);
nand U10266 (N_10266,N_6231,N_7270);
xnor U10267 (N_10267,N_7501,N_6945);
and U10268 (N_10268,N_7492,N_7089);
or U10269 (N_10269,N_6423,N_6036);
xor U10270 (N_10270,N_6432,N_6462);
nor U10271 (N_10271,N_7983,N_8691);
xnor U10272 (N_10272,N_6062,N_8589);
nand U10273 (N_10273,N_8340,N_6538);
nor U10274 (N_10274,N_7785,N_7742);
xnor U10275 (N_10275,N_7916,N_7837);
nor U10276 (N_10276,N_6363,N_7753);
or U10277 (N_10277,N_6543,N_7571);
xor U10278 (N_10278,N_7361,N_7020);
xor U10279 (N_10279,N_7936,N_6161);
or U10280 (N_10280,N_6038,N_7110);
nand U10281 (N_10281,N_7102,N_6833);
nand U10282 (N_10282,N_6141,N_8462);
or U10283 (N_10283,N_7183,N_7872);
nand U10284 (N_10284,N_7449,N_7794);
xor U10285 (N_10285,N_8136,N_8142);
nand U10286 (N_10286,N_6617,N_8138);
and U10287 (N_10287,N_7887,N_6427);
or U10288 (N_10288,N_8150,N_6714);
or U10289 (N_10289,N_8588,N_7081);
and U10290 (N_10290,N_8193,N_7474);
and U10291 (N_10291,N_6070,N_8758);
nand U10292 (N_10292,N_7897,N_6185);
and U10293 (N_10293,N_6553,N_8878);
or U10294 (N_10294,N_6074,N_6080);
nand U10295 (N_10295,N_8904,N_8607);
xor U10296 (N_10296,N_8483,N_8237);
and U10297 (N_10297,N_6325,N_6086);
nand U10298 (N_10298,N_8198,N_6591);
and U10299 (N_10299,N_6260,N_6697);
nor U10300 (N_10300,N_8445,N_8952);
nand U10301 (N_10301,N_8828,N_8577);
and U10302 (N_10302,N_6387,N_7253);
xor U10303 (N_10303,N_8581,N_6323);
and U10304 (N_10304,N_8657,N_7434);
or U10305 (N_10305,N_8173,N_8509);
xor U10306 (N_10306,N_6170,N_7691);
or U10307 (N_10307,N_6060,N_8164);
and U10308 (N_10308,N_6985,N_6103);
nor U10309 (N_10309,N_7924,N_8234);
nor U10310 (N_10310,N_6639,N_7003);
nor U10311 (N_10311,N_8537,N_7471);
and U10312 (N_10312,N_7360,N_7297);
xor U10313 (N_10313,N_6602,N_8766);
and U10314 (N_10314,N_7451,N_7193);
nand U10315 (N_10315,N_7921,N_7518);
or U10316 (N_10316,N_8599,N_6043);
or U10317 (N_10317,N_7678,N_6355);
nand U10318 (N_10318,N_6925,N_6615);
nor U10319 (N_10319,N_6353,N_6425);
or U10320 (N_10320,N_8343,N_6376);
xnor U10321 (N_10321,N_7591,N_7725);
xor U10322 (N_10322,N_6017,N_6012);
or U10323 (N_10323,N_6343,N_6016);
nand U10324 (N_10324,N_8218,N_8630);
and U10325 (N_10325,N_7569,N_7611);
or U10326 (N_10326,N_6478,N_8822);
or U10327 (N_10327,N_8192,N_8572);
or U10328 (N_10328,N_7435,N_6624);
nand U10329 (N_10329,N_7807,N_6698);
and U10330 (N_10330,N_6279,N_8454);
nand U10331 (N_10331,N_7008,N_6296);
or U10332 (N_10332,N_6726,N_6434);
xnor U10333 (N_10333,N_8650,N_6729);
nor U10334 (N_10334,N_6334,N_6209);
nor U10335 (N_10335,N_6131,N_7860);
nor U10336 (N_10336,N_6730,N_6014);
xnor U10337 (N_10337,N_6947,N_7593);
and U10338 (N_10338,N_7906,N_8380);
or U10339 (N_10339,N_6413,N_7410);
nor U10340 (N_10340,N_6357,N_6155);
xor U10341 (N_10341,N_6961,N_7884);
nor U10342 (N_10342,N_8139,N_8643);
nor U10343 (N_10343,N_8159,N_6560);
and U10344 (N_10344,N_8892,N_6841);
nand U10345 (N_10345,N_8424,N_7661);
and U10346 (N_10346,N_8941,N_7891);
and U10347 (N_10347,N_7305,N_6473);
or U10348 (N_10348,N_7832,N_7905);
or U10349 (N_10349,N_7949,N_7212);
nor U10350 (N_10350,N_8374,N_7296);
xnor U10351 (N_10351,N_6707,N_7390);
nor U10352 (N_10352,N_6271,N_7658);
or U10353 (N_10353,N_6502,N_6374);
or U10354 (N_10354,N_8478,N_7356);
and U10355 (N_10355,N_7377,N_7031);
nor U10356 (N_10356,N_7801,N_7468);
nand U10357 (N_10357,N_6982,N_7607);
nand U10358 (N_10358,N_6407,N_7938);
and U10359 (N_10359,N_7105,N_8080);
and U10360 (N_10360,N_6039,N_6705);
nand U10361 (N_10361,N_8678,N_8041);
nand U10362 (N_10362,N_7868,N_6348);
and U10363 (N_10363,N_7697,N_7112);
xnor U10364 (N_10364,N_7075,N_7062);
and U10365 (N_10365,N_7018,N_7605);
or U10366 (N_10366,N_7494,N_8617);
and U10367 (N_10367,N_7729,N_8147);
xor U10368 (N_10368,N_7382,N_8893);
nor U10369 (N_10369,N_8295,N_8806);
xor U10370 (N_10370,N_6199,N_6090);
and U10371 (N_10371,N_7541,N_8252);
or U10372 (N_10372,N_6976,N_7363);
nor U10373 (N_10373,N_7426,N_6299);
nand U10374 (N_10374,N_8539,N_6174);
and U10375 (N_10375,N_8730,N_8339);
or U10376 (N_10376,N_7455,N_7165);
nand U10377 (N_10377,N_7628,N_7331);
and U10378 (N_10378,N_6147,N_8925);
nor U10379 (N_10379,N_7065,N_6801);
xor U10380 (N_10380,N_8862,N_8779);
nor U10381 (N_10381,N_8197,N_7048);
and U10382 (N_10382,N_6519,N_6404);
nor U10383 (N_10383,N_7900,N_6671);
nor U10384 (N_10384,N_7690,N_7431);
or U10385 (N_10385,N_7406,N_8814);
nor U10386 (N_10386,N_8927,N_6625);
nor U10387 (N_10387,N_6930,N_6767);
or U10388 (N_10388,N_6661,N_7023);
nor U10389 (N_10389,N_7817,N_8742);
xnor U10390 (N_10390,N_6115,N_7443);
or U10391 (N_10391,N_8628,N_8794);
and U10392 (N_10392,N_6550,N_6795);
and U10393 (N_10393,N_8370,N_6937);
xor U10394 (N_10394,N_7528,N_6431);
nor U10395 (N_10395,N_8004,N_8671);
and U10396 (N_10396,N_8496,N_8362);
xor U10397 (N_10397,N_6230,N_6463);
nand U10398 (N_10398,N_6024,N_7544);
or U10399 (N_10399,N_7727,N_8415);
nor U10400 (N_10400,N_6261,N_8835);
and U10401 (N_10401,N_7011,N_6179);
and U10402 (N_10402,N_8696,N_6215);
nand U10403 (N_10403,N_8564,N_7937);
or U10404 (N_10404,N_6941,N_8182);
and U10405 (N_10405,N_7991,N_8723);
nor U10406 (N_10406,N_8360,N_8323);
nand U10407 (N_10407,N_8701,N_7237);
nor U10408 (N_10408,N_6597,N_7928);
nor U10409 (N_10409,N_6164,N_8985);
xor U10410 (N_10410,N_6657,N_7454);
or U10411 (N_10411,N_7733,N_7199);
xor U10412 (N_10412,N_8278,N_6644);
nor U10413 (N_10413,N_8974,N_7806);
xor U10414 (N_10414,N_8503,N_6229);
nand U10415 (N_10415,N_7696,N_6806);
and U10416 (N_10416,N_8058,N_7641);
and U10417 (N_10417,N_7113,N_6110);
and U10418 (N_10418,N_7759,N_6912);
or U10419 (N_10419,N_6727,N_8755);
xnor U10420 (N_10420,N_6424,N_8596);
nor U10421 (N_10421,N_6330,N_7272);
nand U10422 (N_10422,N_6254,N_7530);
nand U10423 (N_10423,N_6028,N_7694);
nand U10424 (N_10424,N_8676,N_7168);
or U10425 (N_10425,N_6307,N_7624);
and U10426 (N_10426,N_7574,N_7512);
nand U10427 (N_10427,N_8651,N_8697);
or U10428 (N_10428,N_7407,N_7992);
xnor U10429 (N_10429,N_7359,N_6171);
nand U10430 (N_10430,N_7034,N_7675);
nor U10431 (N_10431,N_8741,N_7304);
and U10432 (N_10432,N_8468,N_6029);
nand U10433 (N_10433,N_6893,N_7149);
nor U10434 (N_10434,N_7944,N_6392);
or U10435 (N_10435,N_6877,N_7215);
nor U10436 (N_10436,N_8538,N_7239);
xor U10437 (N_10437,N_8003,N_8570);
nor U10438 (N_10438,N_8902,N_8535);
nand U10439 (N_10439,N_8180,N_6118);
xnor U10440 (N_10440,N_7602,N_8021);
nor U10441 (N_10441,N_7538,N_7425);
or U10442 (N_10442,N_8663,N_6626);
nand U10443 (N_10443,N_6984,N_6856);
xor U10444 (N_10444,N_6137,N_7266);
or U10445 (N_10445,N_7279,N_6151);
nor U10446 (N_10446,N_6680,N_7514);
or U10447 (N_10447,N_8091,N_8240);
nor U10448 (N_10448,N_8569,N_6779);
nand U10449 (N_10449,N_7056,N_6859);
xnor U10450 (N_10450,N_6072,N_8027);
and U10451 (N_10451,N_6688,N_8455);
xnor U10452 (N_10452,N_6920,N_6784);
or U10453 (N_10453,N_6408,N_8296);
nand U10454 (N_10454,N_6352,N_6400);
xor U10455 (N_10455,N_6614,N_7147);
or U10456 (N_10456,N_8944,N_8351);
and U10457 (N_10457,N_8754,N_8420);
or U10458 (N_10458,N_8662,N_6723);
xor U10459 (N_10459,N_6013,N_7695);
xnor U10460 (N_10460,N_7078,N_8465);
and U10461 (N_10461,N_8988,N_8248);
xnor U10462 (N_10462,N_6902,N_8039);
or U10463 (N_10463,N_7956,N_6989);
and U10464 (N_10464,N_6747,N_6635);
and U10465 (N_10465,N_7484,N_6581);
nand U10466 (N_10466,N_8848,N_6316);
nand U10467 (N_10467,N_7703,N_8649);
and U10468 (N_10468,N_8294,N_7015);
nor U10469 (N_10469,N_7350,N_6690);
nor U10470 (N_10470,N_7095,N_8060);
nor U10471 (N_10471,N_8051,N_6692);
and U10472 (N_10472,N_6004,N_7511);
xor U10473 (N_10473,N_6616,N_8867);
nand U10474 (N_10474,N_8752,N_7391);
nor U10475 (N_10475,N_6211,N_6082);
nor U10476 (N_10476,N_7958,N_8982);
nand U10477 (N_10477,N_7871,N_8184);
or U10478 (N_10478,N_7577,N_6804);
xor U10479 (N_10479,N_7234,N_7289);
or U10480 (N_10480,N_7392,N_8762);
and U10481 (N_10481,N_6448,N_6740);
and U10482 (N_10482,N_8289,N_6106);
xor U10483 (N_10483,N_7913,N_7262);
nor U10484 (N_10484,N_6239,N_7108);
nor U10485 (N_10485,N_6482,N_6257);
nor U10486 (N_10486,N_6962,N_6770);
or U10487 (N_10487,N_7805,N_8979);
or U10488 (N_10488,N_6929,N_8274);
and U10489 (N_10489,N_6222,N_7151);
xnor U10490 (N_10490,N_7549,N_7789);
xnor U10491 (N_10491,N_8464,N_6265);
and U10492 (N_10492,N_6862,N_7743);
xor U10493 (N_10493,N_6535,N_8527);
and U10494 (N_10494,N_6568,N_8556);
nand U10495 (N_10495,N_8861,N_8209);
nand U10496 (N_10496,N_7269,N_6658);
or U10497 (N_10497,N_8642,N_7841);
or U10498 (N_10498,N_6428,N_7161);
or U10499 (N_10499,N_7824,N_7114);
or U10500 (N_10500,N_8033,N_7838);
nand U10501 (N_10501,N_7634,N_8107);
nand U10502 (N_10502,N_6002,N_6734);
xnor U10503 (N_10503,N_6146,N_8763);
nand U10504 (N_10504,N_6920,N_8016);
nor U10505 (N_10505,N_8774,N_6833);
nand U10506 (N_10506,N_8231,N_8577);
or U10507 (N_10507,N_7284,N_8844);
or U10508 (N_10508,N_8947,N_7606);
or U10509 (N_10509,N_7605,N_8428);
nand U10510 (N_10510,N_7527,N_6467);
nor U10511 (N_10511,N_6238,N_7431);
and U10512 (N_10512,N_8621,N_8576);
xor U10513 (N_10513,N_7221,N_7331);
nand U10514 (N_10514,N_6412,N_7066);
and U10515 (N_10515,N_7482,N_6878);
nor U10516 (N_10516,N_6084,N_8997);
xor U10517 (N_10517,N_8632,N_8841);
and U10518 (N_10518,N_7889,N_7671);
and U10519 (N_10519,N_7457,N_6819);
nor U10520 (N_10520,N_8541,N_6430);
or U10521 (N_10521,N_6649,N_6392);
nand U10522 (N_10522,N_8311,N_7217);
xor U10523 (N_10523,N_6139,N_8517);
or U10524 (N_10524,N_7510,N_6399);
nand U10525 (N_10525,N_6504,N_8046);
and U10526 (N_10526,N_7614,N_6237);
nor U10527 (N_10527,N_8028,N_7172);
and U10528 (N_10528,N_8789,N_6728);
xor U10529 (N_10529,N_6351,N_7477);
nand U10530 (N_10530,N_7442,N_7868);
nand U10531 (N_10531,N_8321,N_6052);
and U10532 (N_10532,N_8932,N_8291);
nor U10533 (N_10533,N_7778,N_6281);
nor U10534 (N_10534,N_6716,N_6760);
nor U10535 (N_10535,N_8263,N_8649);
nand U10536 (N_10536,N_6502,N_6129);
nand U10537 (N_10537,N_7555,N_6848);
xnor U10538 (N_10538,N_7632,N_6810);
nand U10539 (N_10539,N_7845,N_6536);
and U10540 (N_10540,N_8809,N_7605);
and U10541 (N_10541,N_7685,N_7585);
or U10542 (N_10542,N_8650,N_8952);
nand U10543 (N_10543,N_8463,N_7125);
nor U10544 (N_10544,N_7977,N_6438);
or U10545 (N_10545,N_6983,N_6389);
or U10546 (N_10546,N_7176,N_7375);
and U10547 (N_10547,N_8732,N_7115);
nor U10548 (N_10548,N_7162,N_8595);
nor U10549 (N_10549,N_6448,N_7871);
nand U10550 (N_10550,N_8650,N_8033);
or U10551 (N_10551,N_7249,N_8622);
xnor U10552 (N_10552,N_6443,N_6465);
and U10553 (N_10553,N_7772,N_8195);
nand U10554 (N_10554,N_7514,N_7935);
nand U10555 (N_10555,N_7315,N_8683);
xnor U10556 (N_10556,N_6193,N_8421);
xor U10557 (N_10557,N_7105,N_8232);
nor U10558 (N_10558,N_7936,N_6556);
and U10559 (N_10559,N_7583,N_6339);
or U10560 (N_10560,N_8787,N_7200);
nand U10561 (N_10561,N_6213,N_7005);
xor U10562 (N_10562,N_8807,N_8172);
or U10563 (N_10563,N_8921,N_7394);
and U10564 (N_10564,N_7339,N_7830);
nor U10565 (N_10565,N_8553,N_7002);
xor U10566 (N_10566,N_6851,N_7773);
and U10567 (N_10567,N_7287,N_6191);
or U10568 (N_10568,N_8860,N_6396);
nand U10569 (N_10569,N_6155,N_8041);
nor U10570 (N_10570,N_6121,N_7581);
and U10571 (N_10571,N_8995,N_8808);
nor U10572 (N_10572,N_7458,N_8486);
xnor U10573 (N_10573,N_8492,N_7660);
and U10574 (N_10574,N_7418,N_8543);
nand U10575 (N_10575,N_8664,N_6700);
nand U10576 (N_10576,N_8134,N_7320);
xor U10577 (N_10577,N_6720,N_6382);
nand U10578 (N_10578,N_7071,N_8161);
xnor U10579 (N_10579,N_8358,N_7058);
nand U10580 (N_10580,N_6425,N_7431);
xnor U10581 (N_10581,N_7000,N_7323);
xnor U10582 (N_10582,N_8047,N_6803);
xnor U10583 (N_10583,N_7008,N_6587);
or U10584 (N_10584,N_7238,N_8674);
or U10585 (N_10585,N_6959,N_7342);
or U10586 (N_10586,N_8760,N_6564);
and U10587 (N_10587,N_8284,N_8299);
or U10588 (N_10588,N_7128,N_6933);
or U10589 (N_10589,N_8561,N_7823);
nand U10590 (N_10590,N_6357,N_7547);
or U10591 (N_10591,N_6924,N_7389);
nor U10592 (N_10592,N_7605,N_8646);
or U10593 (N_10593,N_6424,N_6933);
nand U10594 (N_10594,N_8920,N_8017);
xnor U10595 (N_10595,N_8105,N_6236);
or U10596 (N_10596,N_6350,N_7728);
nand U10597 (N_10597,N_6087,N_8280);
or U10598 (N_10598,N_8776,N_6487);
and U10599 (N_10599,N_6037,N_8645);
or U10600 (N_10600,N_6015,N_7785);
and U10601 (N_10601,N_7978,N_7937);
or U10602 (N_10602,N_8107,N_7998);
nand U10603 (N_10603,N_6445,N_8192);
xnor U10604 (N_10604,N_8822,N_7852);
and U10605 (N_10605,N_6099,N_8246);
nand U10606 (N_10606,N_8986,N_6294);
and U10607 (N_10607,N_6138,N_6211);
and U10608 (N_10608,N_6638,N_6625);
nor U10609 (N_10609,N_8562,N_7453);
xnor U10610 (N_10610,N_7002,N_8632);
xnor U10611 (N_10611,N_6603,N_6019);
nor U10612 (N_10612,N_8891,N_6864);
nor U10613 (N_10613,N_6133,N_7012);
nand U10614 (N_10614,N_8746,N_8489);
nand U10615 (N_10615,N_7463,N_8069);
or U10616 (N_10616,N_8001,N_7494);
and U10617 (N_10617,N_8737,N_6641);
nand U10618 (N_10618,N_6088,N_8470);
nand U10619 (N_10619,N_7979,N_7751);
nand U10620 (N_10620,N_7541,N_6939);
and U10621 (N_10621,N_8970,N_6489);
and U10622 (N_10622,N_6442,N_7559);
nand U10623 (N_10623,N_8867,N_6836);
xnor U10624 (N_10624,N_7606,N_8333);
nor U10625 (N_10625,N_8085,N_7265);
nand U10626 (N_10626,N_7773,N_6938);
or U10627 (N_10627,N_7687,N_6840);
or U10628 (N_10628,N_8243,N_7033);
or U10629 (N_10629,N_6359,N_7011);
or U10630 (N_10630,N_7910,N_7732);
xnor U10631 (N_10631,N_6991,N_8156);
nand U10632 (N_10632,N_8596,N_6050);
nand U10633 (N_10633,N_6974,N_7501);
nor U10634 (N_10634,N_8480,N_6398);
or U10635 (N_10635,N_7630,N_8984);
xor U10636 (N_10636,N_6234,N_7668);
nand U10637 (N_10637,N_8524,N_6071);
nand U10638 (N_10638,N_6556,N_8813);
nor U10639 (N_10639,N_8611,N_6617);
or U10640 (N_10640,N_6681,N_7761);
nand U10641 (N_10641,N_8333,N_8547);
xor U10642 (N_10642,N_8765,N_7879);
or U10643 (N_10643,N_6942,N_8156);
nor U10644 (N_10644,N_8254,N_8649);
or U10645 (N_10645,N_7966,N_8153);
and U10646 (N_10646,N_6748,N_8504);
and U10647 (N_10647,N_7270,N_6365);
or U10648 (N_10648,N_6986,N_6446);
or U10649 (N_10649,N_6416,N_6643);
nand U10650 (N_10650,N_6402,N_8591);
nand U10651 (N_10651,N_7718,N_7007);
xnor U10652 (N_10652,N_8939,N_7867);
nand U10653 (N_10653,N_8894,N_7613);
or U10654 (N_10654,N_6474,N_6312);
and U10655 (N_10655,N_8428,N_8940);
xor U10656 (N_10656,N_7220,N_8417);
and U10657 (N_10657,N_7294,N_8822);
and U10658 (N_10658,N_6545,N_8116);
xnor U10659 (N_10659,N_7191,N_7925);
xor U10660 (N_10660,N_8479,N_6164);
nor U10661 (N_10661,N_8507,N_7416);
nor U10662 (N_10662,N_8004,N_8067);
nor U10663 (N_10663,N_8424,N_8658);
or U10664 (N_10664,N_7286,N_8306);
nor U10665 (N_10665,N_7070,N_7052);
or U10666 (N_10666,N_8095,N_7810);
xor U10667 (N_10667,N_8503,N_7825);
and U10668 (N_10668,N_8684,N_8687);
or U10669 (N_10669,N_6039,N_6207);
or U10670 (N_10670,N_7584,N_8363);
and U10671 (N_10671,N_7962,N_8163);
nand U10672 (N_10672,N_7104,N_8744);
nand U10673 (N_10673,N_8001,N_8760);
or U10674 (N_10674,N_8483,N_7491);
nor U10675 (N_10675,N_6721,N_7481);
or U10676 (N_10676,N_8522,N_7900);
nand U10677 (N_10677,N_6618,N_6206);
or U10678 (N_10678,N_8916,N_7906);
nor U10679 (N_10679,N_8217,N_7771);
or U10680 (N_10680,N_8145,N_8546);
xor U10681 (N_10681,N_7598,N_7279);
and U10682 (N_10682,N_6960,N_7247);
and U10683 (N_10683,N_7373,N_8815);
nor U10684 (N_10684,N_6100,N_7829);
and U10685 (N_10685,N_6771,N_7227);
nor U10686 (N_10686,N_7015,N_7168);
nand U10687 (N_10687,N_7144,N_8647);
or U10688 (N_10688,N_7685,N_6922);
or U10689 (N_10689,N_7319,N_7686);
nor U10690 (N_10690,N_7179,N_8514);
nor U10691 (N_10691,N_8595,N_8576);
xor U10692 (N_10692,N_6304,N_7373);
xnor U10693 (N_10693,N_7744,N_7147);
nand U10694 (N_10694,N_6661,N_7442);
xnor U10695 (N_10695,N_6675,N_7592);
nor U10696 (N_10696,N_7512,N_6711);
nand U10697 (N_10697,N_7348,N_7219);
and U10698 (N_10698,N_7657,N_7949);
or U10699 (N_10699,N_6172,N_8346);
xnor U10700 (N_10700,N_6617,N_6991);
and U10701 (N_10701,N_7718,N_7735);
nor U10702 (N_10702,N_6600,N_8223);
and U10703 (N_10703,N_6563,N_6717);
nand U10704 (N_10704,N_7764,N_6795);
nand U10705 (N_10705,N_6508,N_6350);
nor U10706 (N_10706,N_7047,N_7544);
nand U10707 (N_10707,N_8804,N_6542);
nand U10708 (N_10708,N_8914,N_6154);
nor U10709 (N_10709,N_8674,N_8316);
nand U10710 (N_10710,N_7518,N_7615);
nand U10711 (N_10711,N_8282,N_7078);
nor U10712 (N_10712,N_8377,N_6223);
nor U10713 (N_10713,N_6629,N_7394);
nor U10714 (N_10714,N_8221,N_6856);
and U10715 (N_10715,N_7248,N_6448);
nor U10716 (N_10716,N_6278,N_8344);
xor U10717 (N_10717,N_6040,N_7583);
xnor U10718 (N_10718,N_6887,N_8134);
and U10719 (N_10719,N_6988,N_8217);
nand U10720 (N_10720,N_8250,N_6450);
and U10721 (N_10721,N_8477,N_6867);
or U10722 (N_10722,N_7266,N_7487);
and U10723 (N_10723,N_7507,N_6261);
or U10724 (N_10724,N_8232,N_6073);
or U10725 (N_10725,N_7493,N_7926);
nor U10726 (N_10726,N_6289,N_8329);
or U10727 (N_10727,N_8631,N_8602);
nand U10728 (N_10728,N_6709,N_6988);
xor U10729 (N_10729,N_7223,N_8680);
xnor U10730 (N_10730,N_8405,N_6724);
xnor U10731 (N_10731,N_8648,N_7985);
or U10732 (N_10732,N_7849,N_8163);
or U10733 (N_10733,N_7464,N_7248);
xnor U10734 (N_10734,N_6188,N_6661);
xor U10735 (N_10735,N_8701,N_6437);
nand U10736 (N_10736,N_7122,N_6586);
and U10737 (N_10737,N_8648,N_6358);
or U10738 (N_10738,N_8277,N_8415);
nor U10739 (N_10739,N_6884,N_6650);
xor U10740 (N_10740,N_8939,N_8556);
or U10741 (N_10741,N_8431,N_7033);
nor U10742 (N_10742,N_6885,N_8041);
xor U10743 (N_10743,N_7488,N_7238);
and U10744 (N_10744,N_8656,N_7017);
nand U10745 (N_10745,N_6570,N_7951);
nor U10746 (N_10746,N_7791,N_7815);
nor U10747 (N_10747,N_7703,N_7066);
xor U10748 (N_10748,N_7606,N_7773);
and U10749 (N_10749,N_7753,N_8494);
or U10750 (N_10750,N_8137,N_6868);
or U10751 (N_10751,N_7449,N_8101);
xnor U10752 (N_10752,N_7892,N_7519);
or U10753 (N_10753,N_8895,N_8410);
or U10754 (N_10754,N_8801,N_6087);
nand U10755 (N_10755,N_7989,N_8194);
nor U10756 (N_10756,N_7334,N_7575);
xnor U10757 (N_10757,N_7103,N_6961);
nand U10758 (N_10758,N_8789,N_7723);
nand U10759 (N_10759,N_8337,N_7779);
xor U10760 (N_10760,N_6348,N_8519);
or U10761 (N_10761,N_8118,N_6119);
or U10762 (N_10762,N_6807,N_6504);
or U10763 (N_10763,N_8153,N_8229);
nand U10764 (N_10764,N_7443,N_7134);
nand U10765 (N_10765,N_6149,N_7528);
nand U10766 (N_10766,N_6211,N_6634);
xor U10767 (N_10767,N_6980,N_6983);
xor U10768 (N_10768,N_7583,N_8612);
or U10769 (N_10769,N_7236,N_6180);
xor U10770 (N_10770,N_6770,N_6185);
xnor U10771 (N_10771,N_6923,N_8584);
nand U10772 (N_10772,N_6452,N_8481);
nand U10773 (N_10773,N_6359,N_6030);
nand U10774 (N_10774,N_7945,N_6418);
or U10775 (N_10775,N_8985,N_7267);
nand U10776 (N_10776,N_6778,N_7464);
nand U10777 (N_10777,N_7623,N_7449);
nor U10778 (N_10778,N_7136,N_7386);
nand U10779 (N_10779,N_7370,N_7432);
or U10780 (N_10780,N_8792,N_7692);
nand U10781 (N_10781,N_7286,N_7164);
nand U10782 (N_10782,N_7853,N_7431);
and U10783 (N_10783,N_8141,N_8728);
and U10784 (N_10784,N_8469,N_8361);
xnor U10785 (N_10785,N_7991,N_7368);
nand U10786 (N_10786,N_6406,N_7115);
or U10787 (N_10787,N_6638,N_7327);
xnor U10788 (N_10788,N_7715,N_6562);
and U10789 (N_10789,N_6121,N_8488);
and U10790 (N_10790,N_7462,N_8862);
and U10791 (N_10791,N_8670,N_6773);
or U10792 (N_10792,N_7048,N_7430);
nor U10793 (N_10793,N_7243,N_6466);
nand U10794 (N_10794,N_6956,N_6196);
xor U10795 (N_10795,N_8397,N_6930);
nand U10796 (N_10796,N_6955,N_8078);
nor U10797 (N_10797,N_6430,N_7509);
xnor U10798 (N_10798,N_7277,N_7298);
and U10799 (N_10799,N_7393,N_6624);
or U10800 (N_10800,N_6943,N_7404);
nor U10801 (N_10801,N_7871,N_8700);
and U10802 (N_10802,N_7838,N_8908);
xnor U10803 (N_10803,N_6170,N_6245);
xnor U10804 (N_10804,N_7407,N_7222);
or U10805 (N_10805,N_7424,N_8333);
nand U10806 (N_10806,N_8674,N_8628);
nor U10807 (N_10807,N_6494,N_6931);
nand U10808 (N_10808,N_8825,N_8481);
nand U10809 (N_10809,N_6332,N_8181);
nor U10810 (N_10810,N_6475,N_8095);
nand U10811 (N_10811,N_8679,N_6024);
and U10812 (N_10812,N_6538,N_6185);
nand U10813 (N_10813,N_6493,N_6720);
and U10814 (N_10814,N_8839,N_8358);
nand U10815 (N_10815,N_7768,N_7109);
or U10816 (N_10816,N_7057,N_6915);
nand U10817 (N_10817,N_7128,N_8036);
nand U10818 (N_10818,N_6582,N_8855);
and U10819 (N_10819,N_7945,N_6308);
xor U10820 (N_10820,N_7369,N_8460);
nor U10821 (N_10821,N_6874,N_8996);
and U10822 (N_10822,N_6844,N_8678);
xor U10823 (N_10823,N_7604,N_7061);
xnor U10824 (N_10824,N_8509,N_6443);
nand U10825 (N_10825,N_7005,N_7025);
nor U10826 (N_10826,N_7475,N_7354);
nor U10827 (N_10827,N_6674,N_8405);
nor U10828 (N_10828,N_7530,N_8936);
and U10829 (N_10829,N_7498,N_8169);
nand U10830 (N_10830,N_8000,N_8682);
nor U10831 (N_10831,N_7574,N_8950);
nor U10832 (N_10832,N_6925,N_8257);
xor U10833 (N_10833,N_6554,N_6112);
and U10834 (N_10834,N_6228,N_8666);
nor U10835 (N_10835,N_6324,N_8756);
or U10836 (N_10836,N_7878,N_8997);
and U10837 (N_10837,N_6386,N_6091);
nand U10838 (N_10838,N_7230,N_8876);
nand U10839 (N_10839,N_8547,N_7811);
xnor U10840 (N_10840,N_7205,N_7195);
and U10841 (N_10841,N_6771,N_6057);
xor U10842 (N_10842,N_7443,N_6656);
and U10843 (N_10843,N_6998,N_6088);
xor U10844 (N_10844,N_8632,N_8839);
or U10845 (N_10845,N_8326,N_6843);
and U10846 (N_10846,N_8997,N_6195);
or U10847 (N_10847,N_8216,N_8848);
and U10848 (N_10848,N_8461,N_7641);
nor U10849 (N_10849,N_6221,N_8852);
and U10850 (N_10850,N_7455,N_7652);
xnor U10851 (N_10851,N_8467,N_7549);
xnor U10852 (N_10852,N_6241,N_8773);
nand U10853 (N_10853,N_7709,N_6088);
and U10854 (N_10854,N_7448,N_8598);
xnor U10855 (N_10855,N_7800,N_7657);
xor U10856 (N_10856,N_7773,N_6706);
xnor U10857 (N_10857,N_6391,N_8890);
nor U10858 (N_10858,N_6386,N_6565);
or U10859 (N_10859,N_7946,N_8918);
or U10860 (N_10860,N_8504,N_8341);
nand U10861 (N_10861,N_8059,N_7226);
and U10862 (N_10862,N_6022,N_8476);
nand U10863 (N_10863,N_8463,N_8934);
nand U10864 (N_10864,N_6055,N_6095);
or U10865 (N_10865,N_8591,N_7918);
and U10866 (N_10866,N_6289,N_6130);
or U10867 (N_10867,N_8513,N_7685);
nand U10868 (N_10868,N_6712,N_7440);
nor U10869 (N_10869,N_6358,N_7705);
nand U10870 (N_10870,N_6722,N_7154);
xnor U10871 (N_10871,N_6754,N_6103);
nor U10872 (N_10872,N_8896,N_8547);
or U10873 (N_10873,N_8247,N_7764);
xor U10874 (N_10874,N_7282,N_6923);
nand U10875 (N_10875,N_7020,N_7707);
or U10876 (N_10876,N_8357,N_6973);
nor U10877 (N_10877,N_6454,N_7977);
nor U10878 (N_10878,N_6865,N_8626);
or U10879 (N_10879,N_8160,N_7812);
nand U10880 (N_10880,N_7299,N_8074);
nand U10881 (N_10881,N_8051,N_8430);
nor U10882 (N_10882,N_8448,N_7023);
and U10883 (N_10883,N_7182,N_7091);
xnor U10884 (N_10884,N_8332,N_7759);
nand U10885 (N_10885,N_6453,N_6859);
or U10886 (N_10886,N_8390,N_6140);
nand U10887 (N_10887,N_8220,N_6004);
nor U10888 (N_10888,N_8742,N_6898);
or U10889 (N_10889,N_8291,N_7167);
nand U10890 (N_10890,N_7419,N_8825);
and U10891 (N_10891,N_7984,N_7341);
nand U10892 (N_10892,N_8421,N_6166);
or U10893 (N_10893,N_6843,N_7881);
nand U10894 (N_10894,N_6073,N_7927);
nand U10895 (N_10895,N_7682,N_8545);
nand U10896 (N_10896,N_6866,N_6541);
xor U10897 (N_10897,N_8361,N_8441);
or U10898 (N_10898,N_8778,N_7065);
nand U10899 (N_10899,N_8102,N_8565);
nor U10900 (N_10900,N_8624,N_6887);
nor U10901 (N_10901,N_7175,N_8774);
xor U10902 (N_10902,N_6218,N_7714);
and U10903 (N_10903,N_7073,N_7761);
or U10904 (N_10904,N_6491,N_8811);
nand U10905 (N_10905,N_6544,N_8940);
xor U10906 (N_10906,N_8249,N_8065);
nor U10907 (N_10907,N_6751,N_7670);
xor U10908 (N_10908,N_8494,N_6887);
and U10909 (N_10909,N_7844,N_8829);
nor U10910 (N_10910,N_7177,N_8437);
xor U10911 (N_10911,N_6630,N_8379);
and U10912 (N_10912,N_8039,N_7733);
nor U10913 (N_10913,N_6768,N_8832);
xor U10914 (N_10914,N_7412,N_7697);
nand U10915 (N_10915,N_7826,N_8929);
xnor U10916 (N_10916,N_6490,N_8922);
and U10917 (N_10917,N_8857,N_8286);
and U10918 (N_10918,N_6498,N_8473);
nor U10919 (N_10919,N_7382,N_6024);
nor U10920 (N_10920,N_8116,N_8570);
xor U10921 (N_10921,N_8924,N_6178);
xnor U10922 (N_10922,N_7205,N_7655);
nand U10923 (N_10923,N_6337,N_8706);
nand U10924 (N_10924,N_7447,N_8921);
or U10925 (N_10925,N_7180,N_8739);
xnor U10926 (N_10926,N_8439,N_7845);
and U10927 (N_10927,N_8853,N_6584);
nand U10928 (N_10928,N_8720,N_6043);
or U10929 (N_10929,N_8008,N_8273);
nand U10930 (N_10930,N_6673,N_8899);
nor U10931 (N_10931,N_8262,N_7892);
or U10932 (N_10932,N_8096,N_7451);
and U10933 (N_10933,N_8220,N_7108);
xnor U10934 (N_10934,N_7565,N_7297);
or U10935 (N_10935,N_7129,N_8329);
nand U10936 (N_10936,N_8766,N_6714);
and U10937 (N_10937,N_7139,N_7353);
and U10938 (N_10938,N_7333,N_6303);
xnor U10939 (N_10939,N_7414,N_8311);
or U10940 (N_10940,N_6931,N_6723);
nor U10941 (N_10941,N_7881,N_7130);
or U10942 (N_10942,N_6054,N_6956);
or U10943 (N_10943,N_8961,N_6707);
nor U10944 (N_10944,N_7460,N_6407);
xor U10945 (N_10945,N_8863,N_8293);
nand U10946 (N_10946,N_6691,N_8705);
nor U10947 (N_10947,N_8196,N_7269);
nor U10948 (N_10948,N_6861,N_7660);
xnor U10949 (N_10949,N_7289,N_8620);
xor U10950 (N_10950,N_8445,N_7439);
and U10951 (N_10951,N_6277,N_8270);
or U10952 (N_10952,N_6469,N_7870);
and U10953 (N_10953,N_8521,N_6719);
or U10954 (N_10954,N_6987,N_8559);
nor U10955 (N_10955,N_8463,N_7673);
nor U10956 (N_10956,N_6571,N_6430);
or U10957 (N_10957,N_6866,N_6479);
nor U10958 (N_10958,N_8661,N_8993);
and U10959 (N_10959,N_6262,N_7479);
nor U10960 (N_10960,N_7070,N_8147);
nor U10961 (N_10961,N_6313,N_6861);
xnor U10962 (N_10962,N_8286,N_7719);
or U10963 (N_10963,N_6706,N_8110);
or U10964 (N_10964,N_8926,N_6416);
nor U10965 (N_10965,N_7468,N_8237);
and U10966 (N_10966,N_8538,N_8554);
xor U10967 (N_10967,N_7478,N_6709);
or U10968 (N_10968,N_8149,N_6144);
or U10969 (N_10969,N_6453,N_6966);
or U10970 (N_10970,N_7868,N_7314);
xnor U10971 (N_10971,N_6601,N_8449);
or U10972 (N_10972,N_8957,N_8813);
and U10973 (N_10973,N_7827,N_6846);
or U10974 (N_10974,N_8868,N_8634);
xor U10975 (N_10975,N_6430,N_7197);
and U10976 (N_10976,N_8768,N_8429);
nand U10977 (N_10977,N_7389,N_7607);
nand U10978 (N_10978,N_6488,N_7091);
nand U10979 (N_10979,N_8138,N_6051);
and U10980 (N_10980,N_6266,N_8605);
xor U10981 (N_10981,N_8604,N_8396);
nand U10982 (N_10982,N_7797,N_6653);
and U10983 (N_10983,N_8759,N_6727);
or U10984 (N_10984,N_7691,N_8457);
or U10985 (N_10985,N_7700,N_8628);
and U10986 (N_10986,N_8120,N_6227);
nand U10987 (N_10987,N_6057,N_6142);
nor U10988 (N_10988,N_7325,N_6350);
nand U10989 (N_10989,N_7831,N_8306);
or U10990 (N_10990,N_8196,N_7787);
and U10991 (N_10991,N_6895,N_6263);
xnor U10992 (N_10992,N_8664,N_8031);
nor U10993 (N_10993,N_8063,N_7490);
xnor U10994 (N_10994,N_8279,N_7310);
xor U10995 (N_10995,N_7528,N_8918);
nor U10996 (N_10996,N_7661,N_7697);
and U10997 (N_10997,N_8594,N_8496);
nor U10998 (N_10998,N_6182,N_6390);
xor U10999 (N_10999,N_7518,N_8703);
and U11000 (N_11000,N_8162,N_7569);
nand U11001 (N_11001,N_8124,N_6118);
nor U11002 (N_11002,N_6802,N_6735);
xor U11003 (N_11003,N_7841,N_8340);
or U11004 (N_11004,N_7191,N_6855);
nand U11005 (N_11005,N_7910,N_8849);
and U11006 (N_11006,N_7767,N_6534);
or U11007 (N_11007,N_8446,N_6817);
nand U11008 (N_11008,N_7281,N_6221);
nand U11009 (N_11009,N_6688,N_7617);
and U11010 (N_11010,N_6063,N_7792);
or U11011 (N_11011,N_7178,N_6458);
or U11012 (N_11012,N_7729,N_7876);
and U11013 (N_11013,N_6135,N_6697);
or U11014 (N_11014,N_7050,N_7618);
and U11015 (N_11015,N_7355,N_8610);
and U11016 (N_11016,N_8973,N_8155);
or U11017 (N_11017,N_7737,N_6163);
xor U11018 (N_11018,N_6294,N_6833);
nor U11019 (N_11019,N_8016,N_7282);
nor U11020 (N_11020,N_7167,N_6738);
nor U11021 (N_11021,N_6842,N_6139);
nand U11022 (N_11022,N_7124,N_7277);
nor U11023 (N_11023,N_7837,N_8922);
nor U11024 (N_11024,N_8596,N_6749);
nor U11025 (N_11025,N_8483,N_6576);
or U11026 (N_11026,N_8379,N_8797);
nand U11027 (N_11027,N_6267,N_7565);
and U11028 (N_11028,N_8104,N_6734);
nand U11029 (N_11029,N_8724,N_7076);
nand U11030 (N_11030,N_8301,N_7216);
nand U11031 (N_11031,N_7979,N_8898);
or U11032 (N_11032,N_7110,N_7467);
nand U11033 (N_11033,N_8760,N_7451);
nand U11034 (N_11034,N_7304,N_7745);
nor U11035 (N_11035,N_8415,N_6254);
nor U11036 (N_11036,N_6036,N_8290);
and U11037 (N_11037,N_6320,N_6930);
or U11038 (N_11038,N_8969,N_8935);
nand U11039 (N_11039,N_8360,N_8279);
or U11040 (N_11040,N_7600,N_8809);
nand U11041 (N_11041,N_8695,N_8715);
or U11042 (N_11042,N_8155,N_6339);
and U11043 (N_11043,N_8410,N_7132);
nor U11044 (N_11044,N_6848,N_8799);
nor U11045 (N_11045,N_6899,N_7306);
xnor U11046 (N_11046,N_7579,N_6138);
nor U11047 (N_11047,N_7783,N_6401);
nand U11048 (N_11048,N_7684,N_7107);
xnor U11049 (N_11049,N_8065,N_6083);
or U11050 (N_11050,N_6502,N_6182);
nor U11051 (N_11051,N_8816,N_7328);
nand U11052 (N_11052,N_6007,N_6639);
or U11053 (N_11053,N_6481,N_8389);
nor U11054 (N_11054,N_8094,N_6575);
xor U11055 (N_11055,N_6071,N_8647);
nand U11056 (N_11056,N_7496,N_6981);
nor U11057 (N_11057,N_6809,N_8582);
and U11058 (N_11058,N_6030,N_8840);
and U11059 (N_11059,N_6462,N_8845);
and U11060 (N_11060,N_6332,N_7722);
and U11061 (N_11061,N_7243,N_7633);
or U11062 (N_11062,N_8296,N_6410);
xnor U11063 (N_11063,N_6223,N_6453);
and U11064 (N_11064,N_6748,N_8534);
nor U11065 (N_11065,N_8271,N_7607);
or U11066 (N_11066,N_8463,N_6901);
xnor U11067 (N_11067,N_6702,N_7336);
xor U11068 (N_11068,N_7013,N_7868);
xor U11069 (N_11069,N_7046,N_8565);
nor U11070 (N_11070,N_6443,N_7136);
nor U11071 (N_11071,N_7890,N_7719);
nor U11072 (N_11072,N_8748,N_6178);
nand U11073 (N_11073,N_7958,N_7866);
nor U11074 (N_11074,N_7440,N_8997);
xnor U11075 (N_11075,N_6149,N_8750);
xor U11076 (N_11076,N_7818,N_6938);
nand U11077 (N_11077,N_8802,N_8211);
nand U11078 (N_11078,N_6492,N_6121);
xnor U11079 (N_11079,N_8335,N_8950);
xnor U11080 (N_11080,N_7132,N_6780);
and U11081 (N_11081,N_8552,N_7646);
or U11082 (N_11082,N_8930,N_8475);
and U11083 (N_11083,N_6218,N_7376);
nand U11084 (N_11084,N_6682,N_6924);
or U11085 (N_11085,N_7308,N_7350);
nor U11086 (N_11086,N_6697,N_7326);
or U11087 (N_11087,N_8671,N_7933);
nor U11088 (N_11088,N_8303,N_6765);
nand U11089 (N_11089,N_6983,N_6439);
nor U11090 (N_11090,N_7586,N_6101);
nor U11091 (N_11091,N_7585,N_6798);
xnor U11092 (N_11092,N_8407,N_8820);
and U11093 (N_11093,N_7308,N_7656);
nand U11094 (N_11094,N_8241,N_7513);
nor U11095 (N_11095,N_7342,N_8004);
nor U11096 (N_11096,N_7949,N_7781);
or U11097 (N_11097,N_7166,N_6291);
or U11098 (N_11098,N_6439,N_8570);
and U11099 (N_11099,N_6991,N_7591);
nand U11100 (N_11100,N_6956,N_6832);
xnor U11101 (N_11101,N_6972,N_6580);
nor U11102 (N_11102,N_7142,N_6045);
nand U11103 (N_11103,N_7831,N_7023);
or U11104 (N_11104,N_7348,N_6617);
or U11105 (N_11105,N_6342,N_8157);
or U11106 (N_11106,N_8987,N_8927);
or U11107 (N_11107,N_8578,N_6530);
or U11108 (N_11108,N_8101,N_8034);
or U11109 (N_11109,N_7021,N_8843);
or U11110 (N_11110,N_8379,N_8296);
or U11111 (N_11111,N_8742,N_8619);
nand U11112 (N_11112,N_6328,N_7962);
and U11113 (N_11113,N_6331,N_7565);
or U11114 (N_11114,N_6913,N_6952);
nor U11115 (N_11115,N_6035,N_6834);
xor U11116 (N_11116,N_6426,N_8893);
xor U11117 (N_11117,N_8808,N_8420);
nor U11118 (N_11118,N_6101,N_7524);
nand U11119 (N_11119,N_8687,N_8233);
nor U11120 (N_11120,N_6301,N_6629);
nand U11121 (N_11121,N_7852,N_6771);
nand U11122 (N_11122,N_7725,N_7634);
and U11123 (N_11123,N_7410,N_8608);
and U11124 (N_11124,N_6927,N_7276);
nor U11125 (N_11125,N_7439,N_6301);
nor U11126 (N_11126,N_7308,N_6857);
nor U11127 (N_11127,N_6423,N_8471);
and U11128 (N_11128,N_8751,N_7725);
or U11129 (N_11129,N_8498,N_8782);
nor U11130 (N_11130,N_6999,N_8790);
xnor U11131 (N_11131,N_8548,N_6608);
and U11132 (N_11132,N_6536,N_7426);
xor U11133 (N_11133,N_6534,N_7044);
xnor U11134 (N_11134,N_7728,N_8376);
nor U11135 (N_11135,N_8373,N_6103);
or U11136 (N_11136,N_8203,N_7466);
and U11137 (N_11137,N_6291,N_6030);
and U11138 (N_11138,N_7053,N_6161);
or U11139 (N_11139,N_8124,N_7623);
and U11140 (N_11140,N_8420,N_7098);
and U11141 (N_11141,N_6186,N_7981);
and U11142 (N_11142,N_6301,N_7591);
nor U11143 (N_11143,N_8550,N_7907);
and U11144 (N_11144,N_7202,N_7451);
and U11145 (N_11145,N_8362,N_7724);
xor U11146 (N_11146,N_7428,N_8205);
nand U11147 (N_11147,N_8033,N_8694);
or U11148 (N_11148,N_7234,N_8801);
nand U11149 (N_11149,N_6308,N_7754);
or U11150 (N_11150,N_8254,N_8459);
nand U11151 (N_11151,N_6944,N_8558);
xor U11152 (N_11152,N_7384,N_7648);
nor U11153 (N_11153,N_8834,N_8552);
and U11154 (N_11154,N_6575,N_8263);
nor U11155 (N_11155,N_7341,N_8901);
nor U11156 (N_11156,N_6551,N_7985);
and U11157 (N_11157,N_6855,N_7986);
or U11158 (N_11158,N_7606,N_7492);
nand U11159 (N_11159,N_7386,N_6139);
nor U11160 (N_11160,N_7326,N_7173);
nor U11161 (N_11161,N_6548,N_7435);
nor U11162 (N_11162,N_6472,N_8836);
nor U11163 (N_11163,N_6255,N_8966);
nor U11164 (N_11164,N_7931,N_6247);
xor U11165 (N_11165,N_7355,N_6380);
and U11166 (N_11166,N_7507,N_6246);
and U11167 (N_11167,N_6878,N_7081);
or U11168 (N_11168,N_7314,N_8599);
xnor U11169 (N_11169,N_7645,N_6977);
or U11170 (N_11170,N_7054,N_8936);
xnor U11171 (N_11171,N_8453,N_6502);
xnor U11172 (N_11172,N_6151,N_8528);
and U11173 (N_11173,N_7603,N_6600);
nand U11174 (N_11174,N_8616,N_6677);
nand U11175 (N_11175,N_7317,N_7502);
or U11176 (N_11176,N_7021,N_6213);
xor U11177 (N_11177,N_7254,N_7718);
xnor U11178 (N_11178,N_7565,N_7127);
nor U11179 (N_11179,N_6219,N_7129);
and U11180 (N_11180,N_8375,N_8511);
nand U11181 (N_11181,N_7319,N_7720);
xor U11182 (N_11182,N_8421,N_8553);
nor U11183 (N_11183,N_8372,N_7554);
nor U11184 (N_11184,N_6452,N_6951);
nand U11185 (N_11185,N_6965,N_7368);
nand U11186 (N_11186,N_6362,N_8965);
and U11187 (N_11187,N_8534,N_7383);
xnor U11188 (N_11188,N_6590,N_6528);
and U11189 (N_11189,N_8544,N_6151);
nor U11190 (N_11190,N_8910,N_8476);
nor U11191 (N_11191,N_8833,N_6715);
or U11192 (N_11192,N_7666,N_7828);
or U11193 (N_11193,N_8955,N_7118);
nand U11194 (N_11194,N_7560,N_7833);
nand U11195 (N_11195,N_8585,N_8751);
nand U11196 (N_11196,N_6356,N_8076);
and U11197 (N_11197,N_7422,N_7621);
nor U11198 (N_11198,N_7873,N_6712);
nand U11199 (N_11199,N_7439,N_7316);
nand U11200 (N_11200,N_7691,N_8881);
and U11201 (N_11201,N_7680,N_6599);
or U11202 (N_11202,N_8686,N_7244);
xor U11203 (N_11203,N_6034,N_6811);
and U11204 (N_11204,N_7025,N_6165);
nand U11205 (N_11205,N_8517,N_6087);
nor U11206 (N_11206,N_8107,N_7937);
xor U11207 (N_11207,N_7625,N_8216);
nor U11208 (N_11208,N_8816,N_7174);
xor U11209 (N_11209,N_6353,N_7149);
xnor U11210 (N_11210,N_8576,N_7236);
xor U11211 (N_11211,N_7388,N_8492);
xnor U11212 (N_11212,N_6157,N_6483);
nand U11213 (N_11213,N_7508,N_6651);
nor U11214 (N_11214,N_7730,N_8203);
xor U11215 (N_11215,N_6269,N_8793);
xnor U11216 (N_11216,N_7361,N_6213);
or U11217 (N_11217,N_6416,N_6665);
xor U11218 (N_11218,N_7274,N_8788);
nor U11219 (N_11219,N_6315,N_6435);
nand U11220 (N_11220,N_7322,N_6709);
and U11221 (N_11221,N_7048,N_8173);
nand U11222 (N_11222,N_8012,N_6895);
xnor U11223 (N_11223,N_8294,N_7262);
nor U11224 (N_11224,N_7069,N_8677);
nor U11225 (N_11225,N_6211,N_8332);
and U11226 (N_11226,N_7010,N_8051);
nand U11227 (N_11227,N_6020,N_8773);
and U11228 (N_11228,N_6857,N_6686);
xnor U11229 (N_11229,N_8982,N_6489);
nand U11230 (N_11230,N_6447,N_8758);
or U11231 (N_11231,N_7232,N_7999);
xor U11232 (N_11232,N_8689,N_8822);
nor U11233 (N_11233,N_7426,N_7946);
nand U11234 (N_11234,N_6221,N_7052);
xnor U11235 (N_11235,N_6592,N_8790);
nand U11236 (N_11236,N_6908,N_8135);
nor U11237 (N_11237,N_7722,N_8363);
or U11238 (N_11238,N_7937,N_7636);
xnor U11239 (N_11239,N_6882,N_6744);
and U11240 (N_11240,N_6943,N_8540);
or U11241 (N_11241,N_8240,N_7544);
nor U11242 (N_11242,N_7435,N_6366);
nor U11243 (N_11243,N_7279,N_8202);
nand U11244 (N_11244,N_7683,N_7620);
and U11245 (N_11245,N_6711,N_7579);
or U11246 (N_11246,N_6990,N_8345);
nor U11247 (N_11247,N_6583,N_6408);
nor U11248 (N_11248,N_6686,N_6099);
or U11249 (N_11249,N_8225,N_7654);
or U11250 (N_11250,N_6095,N_8066);
xor U11251 (N_11251,N_6712,N_8491);
and U11252 (N_11252,N_6131,N_6996);
or U11253 (N_11253,N_7177,N_8331);
nand U11254 (N_11254,N_7573,N_7220);
and U11255 (N_11255,N_8091,N_7380);
nand U11256 (N_11256,N_6325,N_6695);
nor U11257 (N_11257,N_6426,N_6830);
nand U11258 (N_11258,N_8615,N_6437);
or U11259 (N_11259,N_7295,N_7178);
nand U11260 (N_11260,N_6429,N_7704);
and U11261 (N_11261,N_8068,N_8060);
xnor U11262 (N_11262,N_6978,N_8723);
xnor U11263 (N_11263,N_7097,N_7343);
and U11264 (N_11264,N_8266,N_6146);
or U11265 (N_11265,N_8234,N_7309);
nand U11266 (N_11266,N_7466,N_8748);
xnor U11267 (N_11267,N_8916,N_7530);
and U11268 (N_11268,N_6894,N_6352);
nand U11269 (N_11269,N_7503,N_7107);
xor U11270 (N_11270,N_6772,N_8134);
nor U11271 (N_11271,N_8754,N_7489);
xor U11272 (N_11272,N_7427,N_8694);
nor U11273 (N_11273,N_6682,N_7608);
or U11274 (N_11274,N_6759,N_8644);
xor U11275 (N_11275,N_8426,N_6048);
nor U11276 (N_11276,N_7230,N_7577);
nand U11277 (N_11277,N_8189,N_6358);
nand U11278 (N_11278,N_8778,N_7139);
nand U11279 (N_11279,N_7539,N_6834);
or U11280 (N_11280,N_8710,N_8820);
nand U11281 (N_11281,N_8907,N_7952);
xnor U11282 (N_11282,N_8433,N_7968);
nor U11283 (N_11283,N_7351,N_7777);
or U11284 (N_11284,N_6760,N_7491);
nand U11285 (N_11285,N_7976,N_8726);
or U11286 (N_11286,N_6016,N_6843);
xor U11287 (N_11287,N_7581,N_7820);
xor U11288 (N_11288,N_8165,N_8764);
nor U11289 (N_11289,N_7954,N_6579);
nor U11290 (N_11290,N_8157,N_7885);
nor U11291 (N_11291,N_7786,N_8978);
nor U11292 (N_11292,N_6869,N_8395);
nand U11293 (N_11293,N_6388,N_6213);
nor U11294 (N_11294,N_6900,N_8359);
or U11295 (N_11295,N_8560,N_6346);
nor U11296 (N_11296,N_6276,N_6222);
or U11297 (N_11297,N_6281,N_6775);
xnor U11298 (N_11298,N_7101,N_7393);
and U11299 (N_11299,N_8810,N_7616);
nor U11300 (N_11300,N_8356,N_6939);
xnor U11301 (N_11301,N_7057,N_7314);
nand U11302 (N_11302,N_8471,N_7083);
and U11303 (N_11303,N_7254,N_8248);
and U11304 (N_11304,N_7950,N_7952);
nand U11305 (N_11305,N_8160,N_6390);
nor U11306 (N_11306,N_7116,N_7726);
nor U11307 (N_11307,N_6895,N_6506);
and U11308 (N_11308,N_8854,N_6749);
and U11309 (N_11309,N_7267,N_6036);
nand U11310 (N_11310,N_8555,N_7538);
nor U11311 (N_11311,N_8316,N_8202);
and U11312 (N_11312,N_7318,N_6936);
xor U11313 (N_11313,N_8030,N_8631);
nor U11314 (N_11314,N_8295,N_7217);
xor U11315 (N_11315,N_7909,N_6235);
nor U11316 (N_11316,N_6981,N_6984);
and U11317 (N_11317,N_7663,N_8824);
or U11318 (N_11318,N_7537,N_7194);
nand U11319 (N_11319,N_8667,N_8495);
nor U11320 (N_11320,N_8741,N_6530);
or U11321 (N_11321,N_8378,N_6225);
and U11322 (N_11322,N_8202,N_7369);
xnor U11323 (N_11323,N_8745,N_7328);
nor U11324 (N_11324,N_6867,N_8446);
xnor U11325 (N_11325,N_7380,N_6191);
xnor U11326 (N_11326,N_6208,N_6653);
nor U11327 (N_11327,N_6572,N_6429);
or U11328 (N_11328,N_6726,N_7291);
nor U11329 (N_11329,N_8622,N_7344);
nand U11330 (N_11330,N_8371,N_8760);
nand U11331 (N_11331,N_7030,N_7034);
nand U11332 (N_11332,N_6243,N_6410);
and U11333 (N_11333,N_6698,N_8426);
nand U11334 (N_11334,N_8426,N_8332);
nor U11335 (N_11335,N_8630,N_8615);
and U11336 (N_11336,N_6453,N_8937);
nand U11337 (N_11337,N_8175,N_7370);
nand U11338 (N_11338,N_8428,N_6002);
nand U11339 (N_11339,N_7259,N_7977);
or U11340 (N_11340,N_7071,N_8890);
nand U11341 (N_11341,N_8313,N_8055);
xnor U11342 (N_11342,N_6885,N_7079);
xor U11343 (N_11343,N_8201,N_7842);
nand U11344 (N_11344,N_6040,N_6075);
or U11345 (N_11345,N_7710,N_6125);
xor U11346 (N_11346,N_7824,N_6400);
xnor U11347 (N_11347,N_7066,N_8062);
xnor U11348 (N_11348,N_8464,N_7012);
and U11349 (N_11349,N_7189,N_8850);
or U11350 (N_11350,N_6140,N_8326);
and U11351 (N_11351,N_7549,N_8681);
xnor U11352 (N_11352,N_6391,N_8166);
nor U11353 (N_11353,N_8075,N_8077);
nor U11354 (N_11354,N_6358,N_7989);
nand U11355 (N_11355,N_6975,N_6048);
nand U11356 (N_11356,N_6657,N_8904);
and U11357 (N_11357,N_8995,N_7617);
nor U11358 (N_11358,N_6939,N_6127);
or U11359 (N_11359,N_8116,N_6733);
or U11360 (N_11360,N_8570,N_7524);
or U11361 (N_11361,N_6563,N_6927);
or U11362 (N_11362,N_8706,N_8688);
nand U11363 (N_11363,N_8085,N_8641);
or U11364 (N_11364,N_8345,N_7107);
nand U11365 (N_11365,N_8033,N_7526);
nor U11366 (N_11366,N_6981,N_6666);
nor U11367 (N_11367,N_8353,N_8685);
or U11368 (N_11368,N_6851,N_8203);
and U11369 (N_11369,N_7583,N_6745);
nor U11370 (N_11370,N_8831,N_8949);
nor U11371 (N_11371,N_7040,N_7294);
nand U11372 (N_11372,N_6832,N_6582);
and U11373 (N_11373,N_6816,N_6024);
nand U11374 (N_11374,N_7470,N_7407);
and U11375 (N_11375,N_8672,N_6405);
nand U11376 (N_11376,N_7652,N_8314);
or U11377 (N_11377,N_7578,N_8034);
nand U11378 (N_11378,N_8052,N_8371);
xnor U11379 (N_11379,N_7466,N_6491);
and U11380 (N_11380,N_8153,N_6569);
or U11381 (N_11381,N_8027,N_8325);
and U11382 (N_11382,N_8390,N_6940);
nand U11383 (N_11383,N_8130,N_8900);
nand U11384 (N_11384,N_7365,N_8006);
and U11385 (N_11385,N_6211,N_6228);
or U11386 (N_11386,N_8320,N_8660);
nor U11387 (N_11387,N_7813,N_7409);
nor U11388 (N_11388,N_6066,N_7393);
nand U11389 (N_11389,N_8664,N_8136);
nor U11390 (N_11390,N_7275,N_8556);
xor U11391 (N_11391,N_7826,N_8515);
nor U11392 (N_11392,N_6818,N_8483);
nand U11393 (N_11393,N_6629,N_6278);
xor U11394 (N_11394,N_6667,N_6565);
xor U11395 (N_11395,N_7684,N_7077);
xor U11396 (N_11396,N_8954,N_6404);
nand U11397 (N_11397,N_7218,N_8433);
nand U11398 (N_11398,N_7250,N_6142);
nand U11399 (N_11399,N_6533,N_7593);
xnor U11400 (N_11400,N_6869,N_8978);
nand U11401 (N_11401,N_7552,N_7205);
and U11402 (N_11402,N_8915,N_8462);
xnor U11403 (N_11403,N_6801,N_8710);
or U11404 (N_11404,N_8861,N_8446);
nor U11405 (N_11405,N_6403,N_7371);
or U11406 (N_11406,N_6201,N_7639);
or U11407 (N_11407,N_7509,N_8727);
or U11408 (N_11408,N_7414,N_6430);
nand U11409 (N_11409,N_7605,N_8326);
and U11410 (N_11410,N_6347,N_8106);
or U11411 (N_11411,N_6581,N_8303);
or U11412 (N_11412,N_8607,N_7312);
nand U11413 (N_11413,N_7356,N_8944);
nand U11414 (N_11414,N_8449,N_7889);
nand U11415 (N_11415,N_6656,N_8944);
and U11416 (N_11416,N_7892,N_7992);
xor U11417 (N_11417,N_7875,N_6330);
xor U11418 (N_11418,N_6291,N_6299);
or U11419 (N_11419,N_6456,N_7246);
nand U11420 (N_11420,N_6705,N_7783);
or U11421 (N_11421,N_7365,N_8080);
nor U11422 (N_11422,N_8750,N_7302);
and U11423 (N_11423,N_6177,N_7904);
or U11424 (N_11424,N_6515,N_8628);
nand U11425 (N_11425,N_6683,N_7582);
nand U11426 (N_11426,N_7513,N_7681);
and U11427 (N_11427,N_8481,N_7049);
and U11428 (N_11428,N_8172,N_6244);
and U11429 (N_11429,N_6304,N_6850);
and U11430 (N_11430,N_8467,N_7712);
nor U11431 (N_11431,N_7191,N_8414);
and U11432 (N_11432,N_8682,N_8826);
nor U11433 (N_11433,N_7503,N_8266);
or U11434 (N_11434,N_8925,N_7880);
nor U11435 (N_11435,N_6372,N_7822);
or U11436 (N_11436,N_7465,N_7232);
and U11437 (N_11437,N_6101,N_6078);
xnor U11438 (N_11438,N_8480,N_6811);
and U11439 (N_11439,N_6534,N_6825);
or U11440 (N_11440,N_7581,N_8380);
and U11441 (N_11441,N_6699,N_6500);
and U11442 (N_11442,N_6415,N_8159);
nor U11443 (N_11443,N_8175,N_6865);
and U11444 (N_11444,N_6395,N_8003);
nor U11445 (N_11445,N_6256,N_8727);
nand U11446 (N_11446,N_6891,N_7109);
nor U11447 (N_11447,N_7437,N_7949);
xor U11448 (N_11448,N_8521,N_8542);
xor U11449 (N_11449,N_6262,N_8136);
and U11450 (N_11450,N_8025,N_8694);
nand U11451 (N_11451,N_8872,N_8119);
and U11452 (N_11452,N_7114,N_6471);
or U11453 (N_11453,N_7890,N_6798);
nor U11454 (N_11454,N_7990,N_6139);
and U11455 (N_11455,N_8713,N_7981);
and U11456 (N_11456,N_7671,N_8667);
or U11457 (N_11457,N_6500,N_6379);
nand U11458 (N_11458,N_8390,N_7862);
nor U11459 (N_11459,N_6894,N_8684);
nor U11460 (N_11460,N_7126,N_8585);
and U11461 (N_11461,N_6947,N_6837);
nand U11462 (N_11462,N_7698,N_8774);
nand U11463 (N_11463,N_7462,N_6235);
nor U11464 (N_11464,N_6600,N_8161);
and U11465 (N_11465,N_7196,N_6845);
nor U11466 (N_11466,N_8442,N_6400);
nand U11467 (N_11467,N_6934,N_8374);
nand U11468 (N_11468,N_7501,N_8178);
nand U11469 (N_11469,N_6869,N_8663);
and U11470 (N_11470,N_8523,N_6632);
nor U11471 (N_11471,N_8359,N_7358);
and U11472 (N_11472,N_6005,N_8135);
and U11473 (N_11473,N_8199,N_7358);
or U11474 (N_11474,N_7233,N_7882);
nor U11475 (N_11475,N_8388,N_8692);
xnor U11476 (N_11476,N_8038,N_6478);
nor U11477 (N_11477,N_7574,N_8174);
and U11478 (N_11478,N_7169,N_6654);
nor U11479 (N_11479,N_6005,N_7901);
xnor U11480 (N_11480,N_6946,N_7894);
nor U11481 (N_11481,N_8870,N_6083);
or U11482 (N_11482,N_7971,N_7120);
nor U11483 (N_11483,N_8987,N_7375);
nand U11484 (N_11484,N_6454,N_6326);
nor U11485 (N_11485,N_6305,N_7775);
or U11486 (N_11486,N_7271,N_7811);
and U11487 (N_11487,N_6583,N_7876);
and U11488 (N_11488,N_6576,N_6636);
nor U11489 (N_11489,N_6064,N_6396);
nor U11490 (N_11490,N_6065,N_6798);
nor U11491 (N_11491,N_7740,N_6462);
nand U11492 (N_11492,N_6963,N_7367);
xnor U11493 (N_11493,N_8941,N_7501);
nand U11494 (N_11494,N_8454,N_7736);
xor U11495 (N_11495,N_7286,N_6933);
or U11496 (N_11496,N_8268,N_6481);
nor U11497 (N_11497,N_6094,N_6058);
or U11498 (N_11498,N_6749,N_6518);
and U11499 (N_11499,N_7884,N_7379);
xor U11500 (N_11500,N_6440,N_7819);
nand U11501 (N_11501,N_6517,N_7158);
and U11502 (N_11502,N_8113,N_7258);
xnor U11503 (N_11503,N_7284,N_8425);
nand U11504 (N_11504,N_8949,N_7538);
xor U11505 (N_11505,N_7452,N_6883);
xor U11506 (N_11506,N_8981,N_7196);
xor U11507 (N_11507,N_7408,N_6415);
and U11508 (N_11508,N_7784,N_7333);
nand U11509 (N_11509,N_7768,N_6235);
nor U11510 (N_11510,N_7464,N_7711);
or U11511 (N_11511,N_7657,N_8754);
and U11512 (N_11512,N_7534,N_8921);
xor U11513 (N_11513,N_8296,N_7570);
nor U11514 (N_11514,N_6164,N_7307);
nor U11515 (N_11515,N_6384,N_7308);
xnor U11516 (N_11516,N_8081,N_7316);
nand U11517 (N_11517,N_8542,N_6579);
nand U11518 (N_11518,N_8702,N_8256);
or U11519 (N_11519,N_7715,N_7441);
xnor U11520 (N_11520,N_7730,N_8079);
nor U11521 (N_11521,N_8000,N_7981);
xor U11522 (N_11522,N_8824,N_6651);
and U11523 (N_11523,N_7355,N_6191);
or U11524 (N_11524,N_6420,N_8992);
nand U11525 (N_11525,N_6793,N_7071);
nor U11526 (N_11526,N_7391,N_8405);
nor U11527 (N_11527,N_7814,N_8112);
nand U11528 (N_11528,N_6029,N_6523);
nor U11529 (N_11529,N_6779,N_8490);
nand U11530 (N_11530,N_7145,N_8862);
and U11531 (N_11531,N_6844,N_8037);
nand U11532 (N_11532,N_6462,N_8218);
or U11533 (N_11533,N_7349,N_8196);
and U11534 (N_11534,N_6246,N_7510);
or U11535 (N_11535,N_7839,N_7317);
or U11536 (N_11536,N_7690,N_6720);
xnor U11537 (N_11537,N_7712,N_7164);
xnor U11538 (N_11538,N_7376,N_6830);
or U11539 (N_11539,N_7836,N_8681);
nor U11540 (N_11540,N_6277,N_7029);
or U11541 (N_11541,N_8171,N_6047);
xnor U11542 (N_11542,N_6871,N_7357);
and U11543 (N_11543,N_6484,N_8486);
nand U11544 (N_11544,N_8345,N_7172);
and U11545 (N_11545,N_8289,N_8491);
and U11546 (N_11546,N_8944,N_8455);
nor U11547 (N_11547,N_8447,N_7806);
nor U11548 (N_11548,N_7001,N_6623);
or U11549 (N_11549,N_6575,N_6017);
and U11550 (N_11550,N_6460,N_8985);
or U11551 (N_11551,N_6229,N_6909);
nor U11552 (N_11552,N_7585,N_8228);
xnor U11553 (N_11553,N_8949,N_8263);
or U11554 (N_11554,N_8831,N_7636);
nand U11555 (N_11555,N_8165,N_7725);
xnor U11556 (N_11556,N_6940,N_6934);
and U11557 (N_11557,N_8729,N_7021);
and U11558 (N_11558,N_8249,N_6748);
and U11559 (N_11559,N_8535,N_6719);
and U11560 (N_11560,N_7613,N_6553);
nand U11561 (N_11561,N_6383,N_8104);
xnor U11562 (N_11562,N_6660,N_8343);
and U11563 (N_11563,N_7335,N_7324);
and U11564 (N_11564,N_6769,N_8920);
nand U11565 (N_11565,N_6756,N_8287);
nor U11566 (N_11566,N_8449,N_6478);
nor U11567 (N_11567,N_7344,N_8070);
xnor U11568 (N_11568,N_7024,N_7552);
nand U11569 (N_11569,N_6359,N_8464);
nor U11570 (N_11570,N_8773,N_6136);
xnor U11571 (N_11571,N_8125,N_8403);
and U11572 (N_11572,N_7858,N_8199);
nand U11573 (N_11573,N_7590,N_8403);
nor U11574 (N_11574,N_8905,N_8393);
or U11575 (N_11575,N_6996,N_8142);
nand U11576 (N_11576,N_7218,N_7895);
and U11577 (N_11577,N_7282,N_8518);
nor U11578 (N_11578,N_6388,N_7715);
nor U11579 (N_11579,N_6883,N_6067);
nand U11580 (N_11580,N_7987,N_7103);
or U11581 (N_11581,N_6160,N_6035);
nor U11582 (N_11582,N_7681,N_8717);
nand U11583 (N_11583,N_7057,N_7562);
nor U11584 (N_11584,N_8645,N_6927);
nor U11585 (N_11585,N_7622,N_7027);
nand U11586 (N_11586,N_8123,N_7281);
and U11587 (N_11587,N_8977,N_7685);
nand U11588 (N_11588,N_7296,N_7320);
nor U11589 (N_11589,N_8726,N_8630);
and U11590 (N_11590,N_7130,N_7399);
and U11591 (N_11591,N_7589,N_6655);
nand U11592 (N_11592,N_6030,N_7445);
xnor U11593 (N_11593,N_7899,N_6511);
xor U11594 (N_11594,N_7424,N_6617);
and U11595 (N_11595,N_8359,N_6362);
and U11596 (N_11596,N_8700,N_6356);
nor U11597 (N_11597,N_8980,N_6041);
and U11598 (N_11598,N_8566,N_7612);
nor U11599 (N_11599,N_6257,N_7244);
and U11600 (N_11600,N_7925,N_7585);
nor U11601 (N_11601,N_8038,N_8245);
xor U11602 (N_11602,N_8716,N_6415);
and U11603 (N_11603,N_7011,N_6640);
xor U11604 (N_11604,N_8667,N_6459);
or U11605 (N_11605,N_8058,N_7025);
nor U11606 (N_11606,N_8817,N_8758);
nor U11607 (N_11607,N_7490,N_7065);
or U11608 (N_11608,N_6771,N_8404);
xor U11609 (N_11609,N_8134,N_6473);
and U11610 (N_11610,N_8327,N_8463);
xor U11611 (N_11611,N_7804,N_6199);
nand U11612 (N_11612,N_7970,N_7161);
nor U11613 (N_11613,N_8378,N_6279);
nand U11614 (N_11614,N_7263,N_7859);
or U11615 (N_11615,N_8493,N_6477);
nor U11616 (N_11616,N_8404,N_8595);
nor U11617 (N_11617,N_6892,N_6432);
nor U11618 (N_11618,N_7248,N_7150);
or U11619 (N_11619,N_6934,N_7998);
and U11620 (N_11620,N_6532,N_6105);
or U11621 (N_11621,N_8283,N_8057);
or U11622 (N_11622,N_7948,N_8779);
or U11623 (N_11623,N_7660,N_7647);
nor U11624 (N_11624,N_7388,N_8094);
xor U11625 (N_11625,N_8061,N_6349);
nor U11626 (N_11626,N_8127,N_7608);
xor U11627 (N_11627,N_7331,N_6772);
nor U11628 (N_11628,N_6523,N_8975);
nor U11629 (N_11629,N_7882,N_8811);
and U11630 (N_11630,N_8144,N_6790);
and U11631 (N_11631,N_8214,N_7620);
nand U11632 (N_11632,N_8617,N_8651);
nand U11633 (N_11633,N_6984,N_6415);
nor U11634 (N_11634,N_6538,N_6079);
nand U11635 (N_11635,N_8771,N_8268);
nor U11636 (N_11636,N_6722,N_8831);
or U11637 (N_11637,N_8239,N_7144);
and U11638 (N_11638,N_7004,N_8493);
nor U11639 (N_11639,N_7879,N_7479);
or U11640 (N_11640,N_8604,N_7868);
and U11641 (N_11641,N_6074,N_7287);
or U11642 (N_11642,N_6372,N_6948);
xor U11643 (N_11643,N_6357,N_7595);
or U11644 (N_11644,N_6874,N_7256);
nor U11645 (N_11645,N_6127,N_7957);
and U11646 (N_11646,N_8951,N_7606);
xnor U11647 (N_11647,N_8024,N_7165);
or U11648 (N_11648,N_6964,N_8195);
or U11649 (N_11649,N_6290,N_6145);
or U11650 (N_11650,N_8343,N_8732);
or U11651 (N_11651,N_8139,N_8182);
nor U11652 (N_11652,N_6536,N_6785);
nand U11653 (N_11653,N_7442,N_6727);
nor U11654 (N_11654,N_7873,N_8473);
or U11655 (N_11655,N_8032,N_6524);
xor U11656 (N_11656,N_6985,N_6171);
xor U11657 (N_11657,N_8801,N_7475);
and U11658 (N_11658,N_8500,N_8266);
nand U11659 (N_11659,N_6400,N_8141);
nand U11660 (N_11660,N_6078,N_8683);
or U11661 (N_11661,N_7498,N_7226);
or U11662 (N_11662,N_6218,N_6899);
or U11663 (N_11663,N_6869,N_8717);
or U11664 (N_11664,N_7346,N_7590);
or U11665 (N_11665,N_8168,N_7676);
or U11666 (N_11666,N_8425,N_7677);
nor U11667 (N_11667,N_6773,N_6861);
nand U11668 (N_11668,N_8995,N_6075);
and U11669 (N_11669,N_7002,N_7261);
nor U11670 (N_11670,N_6940,N_8576);
nand U11671 (N_11671,N_6206,N_6144);
nor U11672 (N_11672,N_7116,N_8215);
nor U11673 (N_11673,N_6242,N_8073);
nand U11674 (N_11674,N_8798,N_7198);
nor U11675 (N_11675,N_8101,N_6055);
or U11676 (N_11676,N_8832,N_6140);
nand U11677 (N_11677,N_7718,N_6482);
and U11678 (N_11678,N_7803,N_8944);
nor U11679 (N_11679,N_6107,N_7587);
nand U11680 (N_11680,N_8858,N_6290);
xnor U11681 (N_11681,N_8750,N_6437);
xor U11682 (N_11682,N_7061,N_6960);
xor U11683 (N_11683,N_6696,N_8428);
xnor U11684 (N_11684,N_8890,N_6691);
and U11685 (N_11685,N_8426,N_6665);
and U11686 (N_11686,N_6827,N_7468);
or U11687 (N_11687,N_8583,N_7586);
or U11688 (N_11688,N_7916,N_8040);
nand U11689 (N_11689,N_7323,N_6364);
xnor U11690 (N_11690,N_7652,N_7760);
nor U11691 (N_11691,N_6165,N_6652);
nand U11692 (N_11692,N_7673,N_6065);
nor U11693 (N_11693,N_8847,N_7817);
xor U11694 (N_11694,N_6944,N_7424);
nand U11695 (N_11695,N_6777,N_6950);
and U11696 (N_11696,N_7362,N_7356);
or U11697 (N_11697,N_8011,N_7864);
nand U11698 (N_11698,N_7120,N_7368);
nor U11699 (N_11699,N_8080,N_7197);
nor U11700 (N_11700,N_7749,N_6926);
nand U11701 (N_11701,N_7954,N_6193);
xor U11702 (N_11702,N_7561,N_7777);
nand U11703 (N_11703,N_7729,N_7668);
xnor U11704 (N_11704,N_8631,N_8809);
or U11705 (N_11705,N_6916,N_6008);
and U11706 (N_11706,N_7690,N_6942);
and U11707 (N_11707,N_8131,N_7432);
or U11708 (N_11708,N_6674,N_6114);
or U11709 (N_11709,N_8298,N_8496);
nor U11710 (N_11710,N_6834,N_8419);
xnor U11711 (N_11711,N_8034,N_6376);
nor U11712 (N_11712,N_6438,N_8878);
nand U11713 (N_11713,N_7292,N_8300);
and U11714 (N_11714,N_8478,N_8301);
and U11715 (N_11715,N_7764,N_6638);
nand U11716 (N_11716,N_8844,N_6912);
and U11717 (N_11717,N_7862,N_6450);
nor U11718 (N_11718,N_8053,N_7187);
and U11719 (N_11719,N_6990,N_7084);
and U11720 (N_11720,N_7121,N_8488);
xor U11721 (N_11721,N_7301,N_6331);
nor U11722 (N_11722,N_8289,N_8793);
and U11723 (N_11723,N_6947,N_8357);
nand U11724 (N_11724,N_7442,N_7053);
or U11725 (N_11725,N_6787,N_6621);
and U11726 (N_11726,N_6039,N_8414);
xor U11727 (N_11727,N_8380,N_7887);
and U11728 (N_11728,N_7785,N_6758);
xnor U11729 (N_11729,N_7044,N_8964);
or U11730 (N_11730,N_6022,N_7942);
and U11731 (N_11731,N_8043,N_8888);
and U11732 (N_11732,N_6060,N_6690);
nor U11733 (N_11733,N_8522,N_7879);
or U11734 (N_11734,N_8924,N_8446);
and U11735 (N_11735,N_8089,N_8739);
or U11736 (N_11736,N_8417,N_8620);
nor U11737 (N_11737,N_6004,N_6971);
or U11738 (N_11738,N_6919,N_8956);
and U11739 (N_11739,N_8671,N_7469);
nand U11740 (N_11740,N_8700,N_6673);
xor U11741 (N_11741,N_8510,N_6920);
nor U11742 (N_11742,N_6681,N_8706);
and U11743 (N_11743,N_6934,N_8898);
or U11744 (N_11744,N_7588,N_6851);
xor U11745 (N_11745,N_6370,N_8997);
and U11746 (N_11746,N_8121,N_8861);
nor U11747 (N_11747,N_6290,N_8045);
nand U11748 (N_11748,N_6893,N_6871);
nand U11749 (N_11749,N_7196,N_7344);
or U11750 (N_11750,N_8887,N_6823);
nor U11751 (N_11751,N_8520,N_8429);
nor U11752 (N_11752,N_6953,N_8531);
and U11753 (N_11753,N_8952,N_6004);
xor U11754 (N_11754,N_7847,N_6967);
nor U11755 (N_11755,N_8618,N_7981);
xnor U11756 (N_11756,N_7716,N_7958);
and U11757 (N_11757,N_7267,N_6898);
and U11758 (N_11758,N_8310,N_7553);
nand U11759 (N_11759,N_7155,N_8081);
xor U11760 (N_11760,N_7481,N_8406);
or U11761 (N_11761,N_7314,N_7010);
nor U11762 (N_11762,N_8872,N_8636);
or U11763 (N_11763,N_7058,N_6755);
nand U11764 (N_11764,N_8938,N_7659);
nor U11765 (N_11765,N_7797,N_7714);
and U11766 (N_11766,N_8884,N_8912);
nand U11767 (N_11767,N_8366,N_7811);
and U11768 (N_11768,N_8827,N_6526);
and U11769 (N_11769,N_8597,N_6344);
and U11770 (N_11770,N_7101,N_6579);
or U11771 (N_11771,N_6245,N_8571);
and U11772 (N_11772,N_8253,N_7601);
xor U11773 (N_11773,N_8479,N_7334);
nand U11774 (N_11774,N_6615,N_7118);
xor U11775 (N_11775,N_8449,N_6970);
nor U11776 (N_11776,N_6520,N_7204);
and U11777 (N_11777,N_7054,N_7081);
or U11778 (N_11778,N_8491,N_6978);
nand U11779 (N_11779,N_7989,N_7619);
xor U11780 (N_11780,N_6727,N_6444);
xnor U11781 (N_11781,N_7748,N_8608);
nand U11782 (N_11782,N_6231,N_6976);
nand U11783 (N_11783,N_6868,N_6020);
nand U11784 (N_11784,N_8324,N_7147);
nor U11785 (N_11785,N_7894,N_8934);
nor U11786 (N_11786,N_6743,N_6605);
nand U11787 (N_11787,N_8329,N_8356);
and U11788 (N_11788,N_6997,N_8184);
nand U11789 (N_11789,N_8828,N_6587);
and U11790 (N_11790,N_8768,N_6827);
and U11791 (N_11791,N_7634,N_6966);
or U11792 (N_11792,N_6936,N_6637);
and U11793 (N_11793,N_6743,N_6552);
nor U11794 (N_11794,N_7385,N_6600);
nor U11795 (N_11795,N_7303,N_6854);
xnor U11796 (N_11796,N_8322,N_8645);
or U11797 (N_11797,N_8257,N_7024);
or U11798 (N_11798,N_7842,N_8922);
xnor U11799 (N_11799,N_8101,N_6725);
nor U11800 (N_11800,N_6649,N_8617);
and U11801 (N_11801,N_7332,N_6124);
nand U11802 (N_11802,N_7323,N_6177);
or U11803 (N_11803,N_6544,N_8609);
and U11804 (N_11804,N_6920,N_8450);
nand U11805 (N_11805,N_8582,N_7757);
and U11806 (N_11806,N_7984,N_6323);
and U11807 (N_11807,N_8678,N_7673);
nand U11808 (N_11808,N_7583,N_6774);
and U11809 (N_11809,N_8122,N_8612);
nand U11810 (N_11810,N_6490,N_6842);
and U11811 (N_11811,N_6185,N_7545);
nand U11812 (N_11812,N_8051,N_7751);
xor U11813 (N_11813,N_6095,N_6805);
nand U11814 (N_11814,N_8702,N_7691);
and U11815 (N_11815,N_8320,N_8435);
nand U11816 (N_11816,N_7511,N_8086);
xnor U11817 (N_11817,N_6821,N_8287);
or U11818 (N_11818,N_6369,N_7687);
xor U11819 (N_11819,N_7951,N_8139);
nor U11820 (N_11820,N_8637,N_6342);
nand U11821 (N_11821,N_6900,N_7777);
nor U11822 (N_11822,N_8022,N_6740);
or U11823 (N_11823,N_7109,N_6480);
nor U11824 (N_11824,N_8982,N_6511);
and U11825 (N_11825,N_7713,N_6387);
or U11826 (N_11826,N_7706,N_7430);
nor U11827 (N_11827,N_7883,N_7460);
nand U11828 (N_11828,N_6713,N_8121);
xor U11829 (N_11829,N_6825,N_8873);
nor U11830 (N_11830,N_7588,N_6149);
or U11831 (N_11831,N_8453,N_7389);
nand U11832 (N_11832,N_8204,N_6983);
nor U11833 (N_11833,N_6768,N_7158);
nand U11834 (N_11834,N_7466,N_6119);
nor U11835 (N_11835,N_6523,N_8788);
or U11836 (N_11836,N_6335,N_6056);
or U11837 (N_11837,N_6590,N_8805);
xor U11838 (N_11838,N_7833,N_8241);
and U11839 (N_11839,N_6012,N_7557);
or U11840 (N_11840,N_7583,N_8062);
nor U11841 (N_11841,N_6377,N_6085);
and U11842 (N_11842,N_6802,N_6104);
xor U11843 (N_11843,N_6150,N_7846);
nand U11844 (N_11844,N_7762,N_6513);
and U11845 (N_11845,N_7718,N_8602);
nor U11846 (N_11846,N_6164,N_7608);
nand U11847 (N_11847,N_6108,N_6480);
nand U11848 (N_11848,N_8334,N_7082);
nor U11849 (N_11849,N_8858,N_6633);
nor U11850 (N_11850,N_8639,N_7184);
or U11851 (N_11851,N_7917,N_8139);
or U11852 (N_11852,N_8811,N_7029);
xor U11853 (N_11853,N_6970,N_7661);
nor U11854 (N_11854,N_7244,N_8736);
xnor U11855 (N_11855,N_8483,N_7480);
xnor U11856 (N_11856,N_8073,N_7688);
and U11857 (N_11857,N_8407,N_8892);
and U11858 (N_11858,N_7617,N_7189);
xor U11859 (N_11859,N_7787,N_6861);
and U11860 (N_11860,N_6389,N_8221);
or U11861 (N_11861,N_7959,N_8741);
and U11862 (N_11862,N_7393,N_8248);
nand U11863 (N_11863,N_7645,N_7853);
nor U11864 (N_11864,N_6706,N_8980);
nand U11865 (N_11865,N_6638,N_7299);
xnor U11866 (N_11866,N_7581,N_6934);
xnor U11867 (N_11867,N_8629,N_7754);
nor U11868 (N_11868,N_8398,N_7143);
nand U11869 (N_11869,N_8138,N_8939);
or U11870 (N_11870,N_8440,N_7184);
or U11871 (N_11871,N_8911,N_7643);
nand U11872 (N_11872,N_6733,N_7169);
or U11873 (N_11873,N_8695,N_7504);
or U11874 (N_11874,N_8366,N_8495);
xor U11875 (N_11875,N_6770,N_8277);
nand U11876 (N_11876,N_8347,N_8209);
and U11877 (N_11877,N_8277,N_6705);
nand U11878 (N_11878,N_8510,N_7845);
and U11879 (N_11879,N_8315,N_6643);
nor U11880 (N_11880,N_6032,N_6176);
nand U11881 (N_11881,N_7408,N_8894);
xnor U11882 (N_11882,N_6787,N_7371);
or U11883 (N_11883,N_7771,N_7381);
xnor U11884 (N_11884,N_7724,N_8730);
or U11885 (N_11885,N_8446,N_8733);
nand U11886 (N_11886,N_6039,N_7319);
xnor U11887 (N_11887,N_6574,N_7398);
nand U11888 (N_11888,N_8900,N_7826);
or U11889 (N_11889,N_6435,N_8190);
or U11890 (N_11890,N_7014,N_7043);
and U11891 (N_11891,N_6738,N_7902);
or U11892 (N_11892,N_7058,N_8023);
nand U11893 (N_11893,N_7339,N_6440);
nor U11894 (N_11894,N_6127,N_7628);
xor U11895 (N_11895,N_6187,N_8570);
nor U11896 (N_11896,N_8023,N_7164);
or U11897 (N_11897,N_6087,N_6565);
and U11898 (N_11898,N_8402,N_8981);
or U11899 (N_11899,N_8121,N_6761);
nor U11900 (N_11900,N_6336,N_6595);
xnor U11901 (N_11901,N_7110,N_8659);
or U11902 (N_11902,N_6220,N_6920);
and U11903 (N_11903,N_6232,N_6206);
nand U11904 (N_11904,N_8798,N_7663);
nand U11905 (N_11905,N_8499,N_7002);
nor U11906 (N_11906,N_8671,N_8419);
nand U11907 (N_11907,N_6010,N_6497);
xnor U11908 (N_11908,N_7730,N_7180);
and U11909 (N_11909,N_7497,N_7986);
xor U11910 (N_11910,N_6681,N_7005);
xnor U11911 (N_11911,N_8128,N_8139);
and U11912 (N_11912,N_6321,N_8018);
nor U11913 (N_11913,N_7976,N_8359);
and U11914 (N_11914,N_8826,N_7684);
and U11915 (N_11915,N_7610,N_6181);
xor U11916 (N_11916,N_8679,N_7892);
nor U11917 (N_11917,N_6075,N_8770);
and U11918 (N_11918,N_7978,N_7251);
and U11919 (N_11919,N_6938,N_7950);
and U11920 (N_11920,N_8333,N_7706);
nor U11921 (N_11921,N_7234,N_6397);
or U11922 (N_11922,N_6718,N_8508);
nor U11923 (N_11923,N_7920,N_7593);
and U11924 (N_11924,N_8337,N_6047);
nand U11925 (N_11925,N_6801,N_6390);
nor U11926 (N_11926,N_6930,N_7364);
or U11927 (N_11927,N_8919,N_7188);
xnor U11928 (N_11928,N_6302,N_6445);
nand U11929 (N_11929,N_8796,N_6795);
xnor U11930 (N_11930,N_7109,N_6884);
and U11931 (N_11931,N_6959,N_6649);
xor U11932 (N_11932,N_8647,N_6291);
xnor U11933 (N_11933,N_7515,N_6022);
or U11934 (N_11934,N_8764,N_7144);
nand U11935 (N_11935,N_8396,N_8470);
or U11936 (N_11936,N_8744,N_7184);
nor U11937 (N_11937,N_6649,N_8651);
xnor U11938 (N_11938,N_8785,N_8246);
nand U11939 (N_11939,N_7942,N_6738);
nand U11940 (N_11940,N_6312,N_8337);
nor U11941 (N_11941,N_6709,N_8967);
and U11942 (N_11942,N_8943,N_6103);
and U11943 (N_11943,N_7906,N_6990);
xor U11944 (N_11944,N_8961,N_7871);
or U11945 (N_11945,N_7200,N_7140);
or U11946 (N_11946,N_8087,N_6813);
nand U11947 (N_11947,N_7356,N_6678);
nand U11948 (N_11948,N_6235,N_7492);
nor U11949 (N_11949,N_6933,N_7014);
xor U11950 (N_11950,N_7153,N_8153);
xnor U11951 (N_11951,N_8163,N_7219);
nor U11952 (N_11952,N_8982,N_7631);
xnor U11953 (N_11953,N_7438,N_8406);
xor U11954 (N_11954,N_6147,N_7261);
and U11955 (N_11955,N_6825,N_6064);
and U11956 (N_11956,N_8971,N_7466);
or U11957 (N_11957,N_6481,N_7515);
nor U11958 (N_11958,N_7787,N_7520);
xnor U11959 (N_11959,N_6077,N_6069);
or U11960 (N_11960,N_8647,N_6999);
or U11961 (N_11961,N_8096,N_8613);
or U11962 (N_11962,N_7722,N_6757);
xor U11963 (N_11963,N_7999,N_7522);
nor U11964 (N_11964,N_8169,N_7638);
and U11965 (N_11965,N_7007,N_8892);
and U11966 (N_11966,N_6480,N_6832);
xor U11967 (N_11967,N_8742,N_8959);
xnor U11968 (N_11968,N_6348,N_7539);
nand U11969 (N_11969,N_6770,N_7937);
and U11970 (N_11970,N_7496,N_7036);
nand U11971 (N_11971,N_8190,N_6254);
nor U11972 (N_11972,N_8376,N_8618);
and U11973 (N_11973,N_7216,N_7019);
and U11974 (N_11974,N_8669,N_8354);
xor U11975 (N_11975,N_6629,N_6385);
and U11976 (N_11976,N_8299,N_8705);
xnor U11977 (N_11977,N_7406,N_6507);
nand U11978 (N_11978,N_6118,N_7227);
xor U11979 (N_11979,N_6445,N_7788);
nand U11980 (N_11980,N_6662,N_6621);
nand U11981 (N_11981,N_8004,N_8558);
nor U11982 (N_11982,N_6867,N_7873);
nor U11983 (N_11983,N_7548,N_7472);
and U11984 (N_11984,N_8382,N_6933);
nand U11985 (N_11985,N_8869,N_6191);
xor U11986 (N_11986,N_8559,N_7282);
and U11987 (N_11987,N_8989,N_6361);
xor U11988 (N_11988,N_6036,N_6397);
nor U11989 (N_11989,N_7205,N_8889);
and U11990 (N_11990,N_8970,N_6594);
or U11991 (N_11991,N_8517,N_6451);
xor U11992 (N_11992,N_8190,N_7418);
and U11993 (N_11993,N_7271,N_6750);
nand U11994 (N_11994,N_6436,N_8023);
and U11995 (N_11995,N_6232,N_7845);
and U11996 (N_11996,N_8141,N_7503);
and U11997 (N_11997,N_7900,N_8933);
nand U11998 (N_11998,N_7825,N_6020);
nor U11999 (N_11999,N_8854,N_6356);
or U12000 (N_12000,N_10145,N_10625);
xor U12001 (N_12001,N_10451,N_10214);
nor U12002 (N_12002,N_11177,N_10830);
nand U12003 (N_12003,N_10762,N_9344);
nor U12004 (N_12004,N_9092,N_9737);
or U12005 (N_12005,N_10493,N_10473);
xnor U12006 (N_12006,N_9840,N_11578);
nand U12007 (N_12007,N_9098,N_9922);
and U12008 (N_12008,N_11333,N_11310);
nand U12009 (N_12009,N_10382,N_9968);
nor U12010 (N_12010,N_9567,N_10458);
nand U12011 (N_12011,N_11789,N_10018);
nor U12012 (N_12012,N_10648,N_11465);
and U12013 (N_12013,N_11258,N_10710);
or U12014 (N_12014,N_11893,N_10770);
nand U12015 (N_12015,N_10836,N_11372);
nor U12016 (N_12016,N_9990,N_9045);
nor U12017 (N_12017,N_9039,N_11937);
xnor U12018 (N_12018,N_11238,N_9655);
nor U12019 (N_12019,N_11999,N_9096);
xnor U12020 (N_12020,N_9759,N_9299);
xor U12021 (N_12021,N_10713,N_11751);
xor U12022 (N_12022,N_11025,N_11883);
nor U12023 (N_12023,N_9306,N_11252);
or U12024 (N_12024,N_9860,N_10035);
nand U12025 (N_12025,N_9276,N_11041);
nand U12026 (N_12026,N_10300,N_9554);
nor U12027 (N_12027,N_11168,N_9172);
and U12028 (N_12028,N_11331,N_9322);
or U12029 (N_12029,N_11544,N_10691);
and U12030 (N_12030,N_10076,N_11290);
nor U12031 (N_12031,N_10450,N_11430);
nand U12032 (N_12032,N_10129,N_10862);
xor U12033 (N_12033,N_9855,N_9366);
nand U12034 (N_12034,N_11795,N_10902);
nor U12035 (N_12035,N_9961,N_10607);
xor U12036 (N_12036,N_10913,N_9674);
nand U12037 (N_12037,N_11039,N_10667);
nor U12038 (N_12038,N_10573,N_11462);
nand U12039 (N_12039,N_9296,N_11126);
xnor U12040 (N_12040,N_9404,N_11065);
nor U12041 (N_12041,N_9771,N_11428);
or U12042 (N_12042,N_11558,N_10707);
xor U12043 (N_12043,N_10668,N_9820);
nor U12044 (N_12044,N_11075,N_11621);
and U12045 (N_12045,N_11996,N_11400);
nor U12046 (N_12046,N_11997,N_10047);
or U12047 (N_12047,N_11125,N_9339);
or U12048 (N_12048,N_10455,N_10860);
nand U12049 (N_12049,N_10333,N_10079);
nand U12050 (N_12050,N_11680,N_9001);
nand U12051 (N_12051,N_9287,N_10271);
nand U12052 (N_12052,N_10213,N_9883);
nand U12053 (N_12053,N_9474,N_9364);
nand U12054 (N_12054,N_10995,N_11181);
nor U12055 (N_12055,N_10327,N_9686);
nand U12056 (N_12056,N_11485,N_10528);
xnor U12057 (N_12057,N_10312,N_11182);
xnor U12058 (N_12058,N_11388,N_10972);
nor U12059 (N_12059,N_9529,N_10436);
or U12060 (N_12060,N_9200,N_10060);
nor U12061 (N_12061,N_10576,N_10928);
and U12062 (N_12062,N_11443,N_10805);
xor U12063 (N_12063,N_10407,N_9218);
nand U12064 (N_12064,N_10099,N_10177);
or U12065 (N_12065,N_9424,N_10751);
nand U12066 (N_12066,N_11165,N_9748);
nor U12067 (N_12067,N_11634,N_10046);
and U12068 (N_12068,N_10235,N_9891);
nor U12069 (N_12069,N_9470,N_9488);
nor U12070 (N_12070,N_11747,N_10133);
or U12071 (N_12071,N_11092,N_9621);
and U12072 (N_12072,N_11198,N_10577);
or U12073 (N_12073,N_10408,N_10949);
or U12074 (N_12074,N_9120,N_9518);
and U12075 (N_12075,N_11414,N_10636);
nor U12076 (N_12076,N_11959,N_11395);
xnor U12077 (N_12077,N_10364,N_11268);
nor U12078 (N_12078,N_11037,N_11345);
nand U12079 (N_12079,N_11088,N_9266);
and U12080 (N_12080,N_9446,N_10238);
and U12081 (N_12081,N_11242,N_10866);
nand U12082 (N_12082,N_11944,N_11974);
nand U12083 (N_12083,N_9485,N_11691);
xnor U12084 (N_12084,N_9274,N_10037);
and U12085 (N_12085,N_10260,N_9901);
and U12086 (N_12086,N_9176,N_9282);
nand U12087 (N_12087,N_10325,N_9784);
or U12088 (N_12088,N_10804,N_9613);
and U12089 (N_12089,N_11033,N_11952);
or U12090 (N_12090,N_11067,N_9556);
nand U12091 (N_12091,N_11197,N_9965);
xor U12092 (N_12092,N_10582,N_10870);
xor U12093 (N_12093,N_11029,N_11890);
or U12094 (N_12094,N_10175,N_10077);
xor U12095 (N_12095,N_10523,N_11149);
nand U12096 (N_12096,N_11275,N_11616);
nand U12097 (N_12097,N_9414,N_10721);
and U12098 (N_12098,N_10356,N_9689);
or U12099 (N_12099,N_9225,N_10033);
xor U12100 (N_12100,N_11353,N_11250);
nand U12101 (N_12101,N_10156,N_11803);
nand U12102 (N_12102,N_11729,N_11061);
and U12103 (N_12103,N_9046,N_9808);
nor U12104 (N_12104,N_9230,N_9641);
nor U12105 (N_12105,N_10499,N_11627);
or U12106 (N_12106,N_10571,N_9328);
nor U12107 (N_12107,N_10551,N_11721);
nand U12108 (N_12108,N_9050,N_11245);
nand U12109 (N_12109,N_9033,N_11507);
or U12110 (N_12110,N_9833,N_11363);
nand U12111 (N_12111,N_11594,N_10242);
nand U12112 (N_12112,N_11506,N_10354);
or U12113 (N_12113,N_11230,N_11051);
xor U12114 (N_12114,N_9249,N_9354);
nand U12115 (N_12115,N_10525,N_10485);
nand U12116 (N_12116,N_10967,N_9233);
and U12117 (N_12117,N_11956,N_11362);
and U12118 (N_12118,N_11313,N_11184);
and U12119 (N_12119,N_10218,N_11934);
and U12120 (N_12120,N_9437,N_9450);
nor U12121 (N_12121,N_9247,N_10651);
and U12122 (N_12122,N_10178,N_11385);
xor U12123 (N_12123,N_10943,N_9338);
xnor U12124 (N_12124,N_11450,N_10696);
and U12125 (N_12125,N_9234,N_11718);
nand U12126 (N_12126,N_9924,N_10012);
or U12127 (N_12127,N_11024,N_10687);
or U12128 (N_12128,N_10587,N_10802);
nand U12129 (N_12129,N_11137,N_11292);
nor U12130 (N_12130,N_11672,N_10011);
nor U12131 (N_12131,N_11328,N_11530);
nand U12132 (N_12132,N_10392,N_9459);
or U12133 (N_12133,N_9169,N_11114);
and U12134 (N_12134,N_10555,N_10813);
nand U12135 (N_12135,N_11917,N_10518);
nand U12136 (N_12136,N_11214,N_11264);
xnor U12137 (N_12137,N_9892,N_11563);
and U12138 (N_12138,N_10224,N_10909);
and U12139 (N_12139,N_10069,N_9810);
xnor U12140 (N_12140,N_11471,N_10665);
nand U12141 (N_12141,N_10210,N_9976);
nor U12142 (N_12142,N_9167,N_9850);
xor U12143 (N_12143,N_10960,N_9876);
nand U12144 (N_12144,N_11112,N_10282);
nand U12145 (N_12145,N_11743,N_9563);
or U12146 (N_12146,N_11581,N_10944);
nor U12147 (N_12147,N_11677,N_10064);
or U12148 (N_12148,N_11063,N_11723);
and U12149 (N_12149,N_11246,N_9580);
and U12150 (N_12150,N_11322,N_11459);
nor U12151 (N_12151,N_10811,N_10381);
and U12152 (N_12152,N_9941,N_9240);
xor U12153 (N_12153,N_10106,N_9762);
nand U12154 (N_12154,N_10112,N_9914);
and U12155 (N_12155,N_9515,N_9889);
nor U12156 (N_12156,N_10876,N_10581);
and U12157 (N_12157,N_11495,N_10301);
nand U12158 (N_12158,N_10789,N_10510);
and U12159 (N_12159,N_10367,N_10918);
and U12160 (N_12160,N_9995,N_11938);
nor U12161 (N_12161,N_9503,N_10790);
and U12162 (N_12162,N_11018,N_10633);
or U12163 (N_12163,N_9704,N_11622);
xnor U12164 (N_12164,N_10136,N_9314);
nor U12165 (N_12165,N_9479,N_11083);
and U12166 (N_12166,N_10647,N_11570);
xnor U12167 (N_12167,N_9177,N_11875);
and U12168 (N_12168,N_11637,N_9464);
and U12169 (N_12169,N_10150,N_11183);
or U12170 (N_12170,N_10245,N_10671);
nand U12171 (N_12171,N_9357,N_11923);
and U12172 (N_12172,N_10754,N_9619);
or U12173 (N_12173,N_11518,N_10706);
nor U12174 (N_12174,N_9003,N_11925);
xor U12175 (N_12175,N_11800,N_10722);
nor U12176 (N_12176,N_9264,N_11087);
xnor U12177 (N_12177,N_9009,N_9930);
and U12178 (N_12178,N_9998,N_11244);
and U12179 (N_12179,N_11864,N_10292);
xnor U12180 (N_12180,N_11775,N_9008);
or U12181 (N_12181,N_11638,N_11505);
or U12182 (N_12182,N_10073,N_10094);
nor U12183 (N_12183,N_9504,N_10021);
nor U12184 (N_12184,N_10773,N_9368);
nand U12185 (N_12185,N_10534,N_9259);
xor U12186 (N_12186,N_10769,N_9236);
nor U12187 (N_12187,N_11633,N_9956);
and U12188 (N_12188,N_10997,N_9679);
and U12189 (N_12189,N_10546,N_10098);
nor U12190 (N_12190,N_10236,N_9035);
xor U12191 (N_12191,N_11030,N_11548);
nand U12192 (N_12192,N_10640,N_11300);
and U12193 (N_12193,N_11138,N_9809);
xnor U12194 (N_12194,N_11208,N_9477);
xnor U12195 (N_12195,N_11907,N_9644);
xor U12196 (N_12196,N_11872,N_9603);
nor U12197 (N_12197,N_11437,N_11920);
nor U12198 (N_12198,N_9238,N_11675);
and U12199 (N_12199,N_9125,N_9138);
or U12200 (N_12200,N_10663,N_11220);
or U12201 (N_12201,N_10514,N_9020);
nor U12202 (N_12202,N_9760,N_11496);
nor U12203 (N_12203,N_9973,N_11109);
nand U12204 (N_12204,N_11528,N_10978);
xor U12205 (N_12205,N_11717,N_9918);
nand U12206 (N_12206,N_11737,N_11591);
or U12207 (N_12207,N_9847,N_11164);
nor U12208 (N_12208,N_11210,N_10222);
nor U12209 (N_12209,N_9559,N_10783);
xor U12210 (N_12210,N_11825,N_11968);
and U12211 (N_12211,N_10730,N_9885);
nor U12212 (N_12212,N_9447,N_11306);
nand U12213 (N_12213,N_11909,N_10677);
nor U12214 (N_12214,N_10384,N_9921);
or U12215 (N_12215,N_9653,N_9182);
nor U12216 (N_12216,N_10290,N_10863);
nand U12217 (N_12217,N_11019,N_11498);
xnor U12218 (N_12218,N_9946,N_11269);
or U12219 (N_12219,N_9409,N_9297);
nor U12220 (N_12220,N_11945,N_9991);
or U12221 (N_12221,N_11641,N_10462);
xor U12222 (N_12222,N_9533,N_11131);
xor U12223 (N_12223,N_10597,N_11396);
and U12224 (N_12224,N_11086,N_11988);
or U12225 (N_12225,N_11546,N_10467);
or U12226 (N_12226,N_9852,N_9508);
xnor U12227 (N_12227,N_11779,N_10448);
and U12228 (N_12228,N_9435,N_9960);
and U12229 (N_12229,N_10919,N_9104);
and U12230 (N_12230,N_11969,N_11735);
nand U12231 (N_12231,N_9849,N_10516);
nor U12232 (N_12232,N_10419,N_9173);
xnor U12233 (N_12233,N_9154,N_11191);
or U12234 (N_12234,N_9523,N_10760);
or U12235 (N_12235,N_9895,N_11812);
nand U12236 (N_12236,N_10296,N_10153);
nand U12237 (N_12237,N_9461,N_10227);
nor U12238 (N_12238,N_10686,N_11798);
and U12239 (N_12239,N_10422,N_9419);
and U12240 (N_12240,N_11059,N_11008);
or U12241 (N_12241,N_9609,N_11116);
nand U12242 (N_12242,N_11480,N_11871);
nand U12243 (N_12243,N_9528,N_11253);
xnor U12244 (N_12244,N_9939,N_9698);
and U12245 (N_12245,N_10501,N_10644);
xor U12246 (N_12246,N_11084,N_9693);
nand U12247 (N_12247,N_9077,N_11984);
nand U12248 (N_12248,N_10067,N_11753);
and U12249 (N_12249,N_10446,N_11719);
xor U12250 (N_12250,N_9324,N_11688);
xnor U12251 (N_12251,N_9040,N_9288);
xnor U12252 (N_12252,N_9627,N_11508);
nor U12253 (N_12253,N_10456,N_11816);
and U12254 (N_12254,N_10299,N_11102);
and U12255 (N_12255,N_9959,N_9842);
nor U12256 (N_12256,N_10093,N_10371);
xnor U12257 (N_12257,N_9822,N_11284);
or U12258 (N_12258,N_9909,N_9325);
or U12259 (N_12259,N_11314,N_10015);
xnor U12260 (N_12260,N_9618,N_10414);
xnor U12261 (N_12261,N_9473,N_11874);
or U12262 (N_12262,N_11017,N_11919);
nand U12263 (N_12263,N_11010,N_10946);
and U12264 (N_12264,N_9545,N_11143);
xnor U12265 (N_12265,N_10947,N_11100);
nor U12266 (N_12266,N_11992,N_10942);
or U12267 (N_12267,N_11884,N_10846);
or U12268 (N_12268,N_10558,N_11689);
xor U12269 (N_12269,N_11998,N_11754);
nand U12270 (N_12270,N_11186,N_9439);
and U12271 (N_12271,N_11993,N_9220);
xor U12272 (N_12272,N_10090,N_11365);
or U12273 (N_12273,N_11673,N_9055);
or U12274 (N_12274,N_10631,N_10981);
or U12275 (N_12275,N_9433,N_10532);
nand U12276 (N_12276,N_9215,N_10190);
or U12277 (N_12277,N_11656,N_10858);
xnor U12278 (N_12278,N_9090,N_10932);
nand U12279 (N_12279,N_9513,N_9100);
and U12280 (N_12280,N_9872,N_11877);
nor U12281 (N_12281,N_9486,N_9662);
nor U12282 (N_12282,N_11575,N_11135);
nand U12283 (N_12283,N_11712,N_10759);
nand U12284 (N_12284,N_9780,N_10645);
xor U12285 (N_12285,N_9517,N_10600);
or U12286 (N_12286,N_11731,N_10729);
xnor U12287 (N_12287,N_11840,N_10383);
nand U12288 (N_12288,N_10971,N_9925);
or U12289 (N_12289,N_10225,N_9659);
xnor U12290 (N_12290,N_11730,N_9813);
and U12291 (N_12291,N_10678,N_10562);
nor U12292 (N_12292,N_11889,N_10491);
or U12293 (N_12293,N_9937,N_11287);
or U12294 (N_12294,N_11739,N_9676);
and U12295 (N_12295,N_10431,N_11440);
nand U12296 (N_12296,N_11232,N_9766);
or U12297 (N_12297,N_11200,N_10684);
xnor U12298 (N_12298,N_10814,N_10063);
and U12299 (N_12299,N_9664,N_10809);
xnor U12300 (N_12300,N_11107,N_9048);
nor U12301 (N_12301,N_11778,N_10536);
nor U12302 (N_12302,N_11733,N_11270);
nand U12303 (N_12303,N_10374,N_11478);
and U12304 (N_12304,N_9629,N_10617);
or U12305 (N_12305,N_9119,N_10748);
and U12306 (N_12306,N_11377,N_10922);
or U12307 (N_12307,N_9067,N_9049);
xnor U12308 (N_12308,N_9058,N_9928);
nand U12309 (N_12309,N_11048,N_9761);
nor U12310 (N_12310,N_11077,N_9560);
and U12311 (N_12311,N_10520,N_11315);
and U12312 (N_12312,N_9795,N_10579);
and U12313 (N_12313,N_11601,N_9178);
nor U12314 (N_12314,N_10480,N_9981);
nand U12315 (N_12315,N_10416,N_10857);
nand U12316 (N_12316,N_10052,N_11750);
xor U12317 (N_12317,N_9188,N_10262);
xnor U12318 (N_12318,N_11399,N_9511);
or U12319 (N_12319,N_11144,N_11845);
or U12320 (N_12320,N_11141,N_9611);
nand U12321 (N_12321,N_10270,N_9384);
nand U12322 (N_12322,N_11127,N_10138);
nor U12323 (N_12323,N_11625,N_10165);
nand U12324 (N_12324,N_11604,N_10482);
and U12325 (N_12325,N_10572,N_10346);
nand U12326 (N_12326,N_10362,N_9544);
and U12327 (N_12327,N_11341,N_10940);
or U12328 (N_12328,N_9815,N_9696);
xor U12329 (N_12329,N_10883,N_9951);
nor U12330 (N_12330,N_10817,N_11914);
nor U12331 (N_12331,N_11068,N_9083);
nand U12332 (N_12332,N_10659,N_11096);
xor U12333 (N_12333,N_10295,N_10660);
xor U12334 (N_12334,N_9974,N_10786);
and U12335 (N_12335,N_11301,N_9642);
nor U12336 (N_12336,N_9223,N_10761);
xnor U12337 (N_12337,N_11967,N_10247);
nor U12338 (N_12338,N_9275,N_11364);
xnor U12339 (N_12339,N_10702,N_11291);
nand U12340 (N_12340,N_9987,N_10741);
and U12341 (N_12341,N_10237,N_11658);
nor U12342 (N_12342,N_10358,N_9212);
nor U12343 (N_12343,N_10329,N_9073);
or U12344 (N_12344,N_10310,N_10560);
and U12345 (N_12345,N_9345,N_10610);
or U12346 (N_12346,N_10767,N_10303);
or U12347 (N_12347,N_9183,N_10612);
nand U12348 (N_12348,N_10894,N_10147);
nand U12349 (N_12349,N_11663,N_9301);
nand U12350 (N_12350,N_9490,N_10843);
nand U12351 (N_12351,N_10143,N_10319);
nor U12352 (N_12352,N_10641,N_9286);
xnor U12353 (N_12353,N_10954,N_11928);
nor U12354 (N_12354,N_11547,N_10544);
nor U12355 (N_12355,N_9400,N_9165);
nor U12356 (N_12356,N_11681,N_11326);
nor U12357 (N_12357,N_9405,N_9564);
nand U12358 (N_12358,N_10887,N_9415);
nand U12359 (N_12359,N_9330,N_10091);
and U12360 (N_12360,N_11987,N_9227);
and U12361 (N_12361,N_11206,N_11768);
and U12362 (N_12362,N_9245,N_10221);
or U12363 (N_12363,N_9174,N_11281);
xor U12364 (N_12364,N_11774,N_9625);
xor U12365 (N_12365,N_10062,N_10251);
xor U12366 (N_12366,N_9062,N_10987);
nand U12367 (N_12367,N_10807,N_10839);
or U12368 (N_12368,N_10342,N_11078);
and U12369 (N_12369,N_11796,N_10249);
and U12370 (N_12370,N_11456,N_9129);
and U12371 (N_12371,N_9697,N_10965);
nand U12372 (N_12372,N_9536,N_11776);
nor U12373 (N_12373,N_11136,N_11091);
nor U12374 (N_12374,N_9992,N_9196);
nor U12375 (N_12375,N_9570,N_9670);
nor U12376 (N_12376,N_10925,N_9658);
and U12377 (N_12377,N_11943,N_10736);
nor U12378 (N_12378,N_11703,N_9380);
nand U12379 (N_12379,N_10041,N_9031);
xnor U12380 (N_12380,N_10731,N_10912);
and U12381 (N_12381,N_10475,N_11389);
xor U12382 (N_12382,N_11057,N_11271);
xor U12383 (N_12383,N_11603,N_9351);
or U12384 (N_12384,N_11299,N_9327);
and U12385 (N_12385,N_10939,N_11529);
nor U12386 (N_12386,N_10726,N_11043);
nand U12387 (N_12387,N_9298,N_11757);
and U12388 (N_12388,N_9730,N_9478);
or U12389 (N_12389,N_10599,N_10901);
and U12390 (N_12390,N_9255,N_10897);
and U12391 (N_12391,N_9391,N_11808);
and U12392 (N_12392,N_9445,N_9476);
xor U12393 (N_12393,N_10353,N_11879);
nand U12394 (N_12394,N_10435,N_11935);
nor U12395 (N_12395,N_9512,N_9436);
or U12396 (N_12396,N_10421,N_9416);
and U12397 (N_12397,N_9920,N_9871);
nand U12398 (N_12398,N_10543,N_10845);
nor U12399 (N_12399,N_10410,N_10026);
or U12400 (N_12400,N_10822,N_9421);
nand U12401 (N_12401,N_9688,N_11404);
xnor U12402 (N_12402,N_9019,N_9814);
xor U12403 (N_12403,N_11302,N_10935);
nor U12404 (N_12404,N_10183,N_9350);
or U12405 (N_12405,N_11015,N_9029);
or U12406 (N_12406,N_9806,N_9955);
nor U12407 (N_12407,N_10994,N_10465);
xor U12408 (N_12408,N_10698,N_9668);
nor U12409 (N_12409,N_10970,N_10505);
xnor U12410 (N_12410,N_10714,N_9673);
nor U12411 (N_12411,N_10893,N_9043);
or U12412 (N_12412,N_9831,N_11780);
nand U12413 (N_12413,N_10293,N_11076);
nand U12414 (N_12414,N_9783,N_10399);
nor U12415 (N_12415,N_10083,N_10350);
xor U12416 (N_12416,N_10287,N_10500);
or U12417 (N_12417,N_9546,N_9557);
xor U12418 (N_12418,N_11817,N_10793);
xnor U12419 (N_12419,N_9336,N_9816);
or U12420 (N_12420,N_9317,N_9495);
xor U12421 (N_12421,N_10208,N_9086);
nor U12422 (N_12422,N_9005,N_9051);
xnor U12423 (N_12423,N_10137,N_11202);
or U12424 (N_12424,N_11454,N_9422);
and U12425 (N_12425,N_9132,N_9037);
and U12426 (N_12426,N_10019,N_11892);
and U12427 (N_12427,N_10277,N_11585);
nand U12428 (N_12428,N_9811,N_9054);
and U12429 (N_12429,N_10892,N_10487);
xnor U12430 (N_12430,N_9047,N_10205);
xnor U12431 (N_12431,N_11110,N_9499);
xor U12432 (N_12432,N_9028,N_10345);
and U12433 (N_12433,N_10844,N_11806);
nor U12434 (N_12434,N_9701,N_9595);
nand U12435 (N_12435,N_9209,N_11439);
or U12436 (N_12436,N_9988,N_10801);
and U12437 (N_12437,N_9458,N_10693);
nor U12438 (N_12438,N_11312,N_10497);
or U12439 (N_12439,N_11720,N_10728);
or U12440 (N_12440,N_10005,N_11249);
nand U12441 (N_12441,N_11390,N_11766);
xor U12442 (N_12442,N_10771,N_10373);
xor U12443 (N_12443,N_11490,N_10996);
nor U12444 (N_12444,N_10874,N_10439);
xnor U12445 (N_12445,N_11488,N_10618);
nor U12446 (N_12446,N_11932,N_10232);
xor U12447 (N_12447,N_11105,N_10873);
or U12448 (N_12448,N_11229,N_11560);
or U12449 (N_12449,N_9402,N_10733);
xnor U12450 (N_12450,N_11148,N_10658);
or U12451 (N_12451,N_10288,N_11374);
or U12452 (N_12452,N_11976,N_9709);
or U12453 (N_12453,N_11749,N_9251);
nor U12454 (N_12454,N_11626,N_11429);
xor U12455 (N_12455,N_9752,N_10766);
xor U12456 (N_12456,N_11701,N_11784);
nor U12457 (N_12457,N_11908,N_10828);
and U12458 (N_12458,N_11128,N_9870);
or U12459 (N_12459,N_11402,N_11397);
and U12460 (N_12460,N_10621,N_10529);
or U12461 (N_12461,N_11477,N_11553);
or U12462 (N_12462,N_10923,N_9703);
nor U12463 (N_12463,N_11413,N_10402);
and U12464 (N_12464,N_11464,N_11123);
and U12465 (N_12465,N_10425,N_10256);
nand U12466 (N_12466,N_10952,N_9411);
or U12467 (N_12467,N_11042,N_10724);
and U12468 (N_12468,N_9294,N_11394);
or U12469 (N_12469,N_9004,N_10782);
xnor U12470 (N_12470,N_10157,N_11145);
or U12471 (N_12471,N_11915,N_10070);
and U12472 (N_12472,N_10979,N_9650);
or U12473 (N_12473,N_10168,N_10378);
xor U12474 (N_12474,N_10144,N_10865);
nor U12475 (N_12475,N_10081,N_10494);
nor U12476 (N_12476,N_9293,N_11347);
or U12477 (N_12477,N_10246,N_10102);
or U12478 (N_12478,N_10778,N_9950);
nor U12479 (N_12479,N_10438,N_11865);
xor U12480 (N_12480,N_11133,N_11205);
xnor U12481 (N_12481,N_9952,N_9520);
nand U12482 (N_12482,N_10200,N_11103);
nand U12483 (N_12483,N_10385,N_10524);
nor U12484 (N_12484,N_10082,N_11522);
nand U12485 (N_12485,N_11949,N_11421);
nand U12486 (N_12486,N_11631,N_10459);
and U12487 (N_12487,N_10001,N_11767);
xnor U12488 (N_12488,N_11847,N_10348);
nor U12489 (N_12489,N_9143,N_10634);
nor U12490 (N_12490,N_11339,N_9094);
nor U12491 (N_12491,N_11973,N_10962);
nor U12492 (N_12492,N_9455,N_9827);
xnor U12493 (N_12493,N_9615,N_9015);
nand U12494 (N_12494,N_10132,N_11455);
nand U12495 (N_12495,N_9329,N_10565);
xor U12496 (N_12496,N_11012,N_9856);
nand U12497 (N_12497,N_10492,N_10444);
and U12498 (N_12498,N_10688,N_9623);
and U12499 (N_12499,N_10241,N_9318);
and U12500 (N_12500,N_9597,N_11317);
xor U12501 (N_12501,N_10167,N_10498);
and U12502 (N_12502,N_10248,N_9708);
and U12503 (N_12503,N_10915,N_10420);
and U12504 (N_12504,N_11885,N_11446);
and U12505 (N_12505,N_9152,N_9389);
nand U12506 (N_12506,N_11159,N_9792);
nor U12507 (N_12507,N_10993,N_9149);
and U12508 (N_12508,N_9449,N_9017);
or U12509 (N_12509,N_9887,N_9427);
or U12510 (N_12510,N_11419,N_10298);
nand U12511 (N_12511,N_9309,N_10888);
nor U12512 (N_12512,N_10533,N_11081);
and U12513 (N_12513,N_9337,N_10240);
nand U12514 (N_12514,N_11922,N_11927);
nand U12515 (N_12515,N_9428,N_10715);
xor U12516 (N_12516,N_9630,N_11584);
nor U12517 (N_12517,N_9878,N_10530);
and U12518 (N_12518,N_10437,N_11398);
nor U12519 (N_12519,N_11280,N_9541);
and U12520 (N_12520,N_11572,N_9505);
xor U12521 (N_12521,N_10413,N_9304);
nand U12522 (N_12522,N_9095,N_11423);
and U12523 (N_12523,N_11157,N_11288);
nand U12524 (N_12524,N_11004,N_11234);
xnor U12525 (N_12525,N_10948,N_9977);
and U12526 (N_12526,N_11671,N_11866);
nand U12527 (N_12527,N_9694,N_10105);
nor U12528 (N_12528,N_9064,N_11684);
and U12529 (N_12529,N_11022,N_9857);
or U12530 (N_12530,N_9131,N_10119);
nand U12531 (N_12531,N_10095,N_10531);
nor U12532 (N_12532,N_11263,N_9371);
nor U12533 (N_12533,N_11327,N_10481);
xnor U12534 (N_12534,N_10363,N_9489);
nand U12535 (N_12535,N_11282,N_11755);
or U12536 (N_12536,N_9647,N_10116);
nand U12537 (N_12537,N_11378,N_10139);
nand U12538 (N_12538,N_10743,N_9678);
nand U12539 (N_12539,N_9616,N_10825);
nor U12540 (N_12540,N_11602,N_11140);
nor U12541 (N_12541,N_9861,N_11254);
and U12542 (N_12542,N_9553,N_11223);
and U12543 (N_12543,N_11824,N_9726);
nand U12544 (N_12544,N_9160,N_10429);
nor U12545 (N_12545,N_10567,N_10685);
nand U12546 (N_12546,N_9369,N_11352);
and U12547 (N_12547,N_11501,N_10896);
xor U12548 (N_12548,N_9824,N_9797);
and U12549 (N_12549,N_11196,N_9599);
nand U12550 (N_12550,N_9863,N_11849);
xnor U12551 (N_12551,N_11513,N_9184);
or U12552 (N_12552,N_9738,N_11823);
and U12553 (N_12553,N_9242,N_10750);
nand U12554 (N_12554,N_11316,N_9168);
and U12555 (N_12555,N_11119,N_11700);
and U12556 (N_12556,N_9983,N_10154);
nand U12557 (N_12557,N_9442,N_10191);
or U12558 (N_12558,N_11903,N_11697);
xnor U12559 (N_12559,N_11930,N_10197);
nor U12560 (N_12560,N_9507,N_10694);
xor U12561 (N_12561,N_10050,N_10903);
nand U12562 (N_12562,N_9851,N_10611);
or U12563 (N_12563,N_11525,N_9044);
xnor U12564 (N_12564,N_10072,N_10406);
or U12565 (N_12565,N_11303,N_11947);
or U12566 (N_12566,N_9101,N_10320);
and U12567 (N_12567,N_11901,N_11690);
nand U12568 (N_12568,N_9501,N_11325);
nand U12569 (N_12569,N_10936,N_11511);
and U12570 (N_12570,N_10110,N_10933);
nand U12571 (N_12571,N_11055,N_11367);
xnor U12572 (N_12572,N_11369,N_10606);
or U12573 (N_12573,N_9363,N_11714);
and U12574 (N_12574,N_11964,N_10910);
and U12575 (N_12575,N_11405,N_10590);
and U12576 (N_12576,N_10871,N_10788);
nor U12577 (N_12577,N_9190,N_10326);
and U12578 (N_12578,N_10261,N_9530);
xor U12579 (N_12579,N_11438,N_10220);
nor U12580 (N_12580,N_10624,N_10742);
nand U12581 (N_12581,N_11512,N_11646);
nand U12582 (N_12582,N_9395,N_10423);
nand U12583 (N_12583,N_11759,N_9605);
and U12584 (N_12584,N_11668,N_10244);
nand U12585 (N_12585,N_11989,N_9890);
xor U12586 (N_12586,N_10953,N_9097);
and U12587 (N_12587,N_9375,N_10286);
or U12588 (N_12588,N_10723,N_11071);
nor U12589 (N_12589,N_11896,N_10768);
nor U12590 (N_12590,N_9724,N_10718);
xnor U12591 (N_12591,N_9940,N_9588);
xor U12592 (N_12592,N_11176,N_9802);
nor U12593 (N_12593,N_10921,N_10331);
nor U12594 (N_12594,N_9569,N_11227);
xor U12595 (N_12595,N_9999,N_9151);
nor U12596 (N_12596,N_11278,N_11657);
nand U12597 (N_12597,N_9295,N_11873);
xnor U12598 (N_12598,N_11929,N_11910);
and U12599 (N_12599,N_11261,N_9202);
and U12600 (N_12600,N_10151,N_9253);
nor U12601 (N_12601,N_9313,N_9583);
or U12602 (N_12602,N_11203,N_10652);
nor U12603 (N_12603,N_9542,N_9030);
xnor U12604 (N_12604,N_11382,N_11773);
nand U12605 (N_12605,N_10539,N_10080);
or U12606 (N_12606,N_9122,N_9224);
xor U12607 (N_12607,N_10661,N_10330);
or U12608 (N_12608,N_11106,N_9341);
nand U12609 (N_12609,N_11062,N_11375);
and U12610 (N_12610,N_11842,N_10442);
or U12611 (N_12611,N_11047,N_9463);
or U12612 (N_12612,N_9656,N_9099);
nand U12613 (N_12613,N_10441,N_11225);
or U12614 (N_12614,N_10716,N_11589);
nand U12615 (N_12615,N_10864,N_11134);
xor U12616 (N_12616,N_11682,N_10537);
nand U12617 (N_12617,N_10049,N_10460);
xor U12618 (N_12618,N_11870,N_9355);
or U12619 (N_12619,N_9964,N_10302);
nor U12620 (N_12620,N_9263,N_10074);
xnor U12621 (N_12621,N_9980,N_10488);
or U12622 (N_12622,N_10044,N_11318);
nand U12623 (N_12623,N_11053,N_10810);
nand U12624 (N_12624,N_10700,N_9285);
or U12625 (N_12625,N_10628,N_11624);
or U12626 (N_12626,N_10917,N_10973);
and U12627 (N_12627,N_9448,N_11003);
nor U12628 (N_12628,N_11034,N_9651);
xnor U12629 (N_12629,N_9118,N_9397);
xnor U12630 (N_12630,N_9805,N_9607);
or U12631 (N_12631,N_9828,N_11777);
nor U12632 (N_12632,N_11822,N_11858);
and U12633 (N_12633,N_11412,N_10229);
nand U12634 (N_12634,N_11607,N_10194);
or U12635 (N_12635,N_9899,N_9141);
xnor U12636 (N_12636,N_11441,N_9103);
and U12637 (N_12637,N_9213,N_9565);
nand U12638 (N_12638,N_11898,N_9586);
or U12639 (N_12639,N_9754,N_10443);
and U12640 (N_12640,N_10690,N_11586);
xor U12641 (N_12641,N_10614,N_9365);
nand U12642 (N_12642,N_9024,N_9181);
and U12643 (N_12643,N_11595,N_11173);
or U12644 (N_12644,N_10604,N_9158);
xor U12645 (N_12645,N_10483,N_9953);
and U12646 (N_12646,N_11212,N_9578);
nor U12647 (N_12647,N_10040,N_10914);
or U12648 (N_12648,N_10017,N_11211);
and U12649 (N_12649,N_10638,N_10071);
nand U12650 (N_12650,N_10440,N_10841);
nor U12651 (N_12651,N_11069,N_9057);
xnor U12652 (N_12652,N_11573,N_9500);
nor U12653 (N_12653,N_11435,N_11502);
nor U12654 (N_12654,N_10349,N_9739);
xor U12655 (N_12655,N_9127,N_9270);
nor U12656 (N_12656,N_9390,N_10267);
and U12657 (N_12657,N_9066,N_9429);
and U12658 (N_12658,N_9034,N_11746);
and U12659 (N_12659,N_10605,N_9845);
nor U12660 (N_12660,N_9023,N_9430);
xor U12661 (N_12661,N_10526,N_10215);
and U12662 (N_12662,N_11539,N_11826);
or U12663 (N_12663,N_9787,N_9880);
nor U12664 (N_12664,N_11676,N_10596);
xor U12665 (N_12665,N_10365,N_11130);
or U12666 (N_12666,N_10471,N_9088);
xor U12667 (N_12667,N_11918,N_11576);
and U12668 (N_12668,N_10502,N_11537);
nor U12669 (N_12669,N_11770,N_10198);
nand U12670 (N_12670,N_11476,N_10827);
xnor U12671 (N_12671,N_9021,N_11645);
nor U12672 (N_12672,N_9133,N_9769);
or U12673 (N_12673,N_11966,N_10679);
and U12674 (N_12674,N_10785,N_10317);
or U12675 (N_12675,N_10400,N_9041);
nor U12676 (N_12676,N_10124,N_11336);
or U12677 (N_12677,N_9764,N_9982);
and U12678 (N_12678,N_10162,N_11283);
xnor U12679 (N_12679,N_9214,N_10449);
and U12680 (N_12680,N_11702,N_11970);
nor U12681 (N_12681,N_10574,N_9614);
and U12682 (N_12682,N_10022,N_9244);
and U12683 (N_12683,N_10988,N_9626);
and U12684 (N_12684,N_9823,N_10812);
and U12685 (N_12685,N_10798,N_11451);
nand U12686 (N_12686,N_11216,N_9381);
or U12687 (N_12687,N_11171,N_10032);
nand U12688 (N_12688,N_9487,N_10906);
or U12689 (N_12689,N_11349,N_10586);
and U12690 (N_12690,N_11834,N_11707);
nand U12691 (N_12691,N_9969,N_10272);
and U12692 (N_12692,N_9271,N_9592);
nor U12693 (N_12693,N_10507,N_10603);
or U12694 (N_12694,N_9012,N_9821);
nand U12695 (N_12695,N_9519,N_10609);
or U12696 (N_12696,N_11981,N_9643);
and U12697 (N_12697,N_9532,N_11361);
xor U12698 (N_12698,N_10039,N_10930);
and U12699 (N_12699,N_9466,N_10057);
or U12700 (N_12700,N_10990,N_11384);
nand U12701 (N_12701,N_11695,N_10547);
or U12702 (N_12702,N_9514,N_10155);
or U12703 (N_12703,N_11309,N_10055);
nand U12704 (N_12704,N_10484,N_10254);
or U12705 (N_12705,N_9175,N_10486);
nor U12706 (N_12706,N_9742,N_11577);
xnor U12707 (N_12707,N_9291,N_10206);
nand U12708 (N_12708,N_9864,N_11050);
and U12709 (N_12709,N_10130,N_9936);
xor U12710 (N_12710,N_9640,N_9745);
nor U12711 (N_12711,N_11659,N_10720);
nor U12712 (N_12712,N_11948,N_10622);
xor U12713 (N_12713,N_10253,N_10334);
nor U12714 (N_12714,N_9734,N_11342);
nor U12715 (N_12715,N_10010,N_11965);
or U12716 (N_12716,N_10956,N_10166);
nand U12717 (N_12717,N_10613,N_10852);
and U12718 (N_12718,N_10905,N_10008);
or U12719 (N_12719,N_11763,N_9123);
and U12720 (N_12720,N_11289,N_9835);
nor U12721 (N_12721,N_11426,N_9721);
or U12722 (N_12722,N_9460,N_9231);
xnor U12723 (N_12723,N_11785,N_9370);
and U12724 (N_12724,N_9632,N_11162);
and U12725 (N_12725,N_11393,N_11726);
and U12726 (N_12726,N_10837,N_11129);
nand U12727 (N_12727,N_9273,N_9228);
xor U12728 (N_12728,N_10212,N_9915);
nand U12729 (N_12729,N_9690,N_11355);
or U12730 (N_12730,N_11744,N_11598);
nand U12731 (N_12731,N_9916,N_9957);
or U12732 (N_12732,N_9204,N_11474);
xor U12733 (N_12733,N_11222,N_11980);
or U12734 (N_12734,N_10890,N_11085);
or U12735 (N_12735,N_11497,N_11597);
xnor U12736 (N_12736,N_11237,N_10279);
and U12737 (N_12737,N_11523,N_10740);
and U12738 (N_12738,N_9434,N_9566);
or U12739 (N_12739,N_11359,N_11756);
nor U12740 (N_12740,N_11562,N_11297);
xor U12741 (N_12741,N_9777,N_9074);
nor U12742 (N_12742,N_11178,N_10265);
xnor U12743 (N_12743,N_10563,N_9812);
or U12744 (N_12744,N_11556,N_10580);
nor U12745 (N_12745,N_9741,N_10369);
xnor U12746 (N_12746,N_11859,N_11960);
and U12747 (N_12747,N_11962,N_9216);
and U12748 (N_12748,N_9598,N_11118);
or U12749 (N_12749,N_10375,N_11642);
xor U12750 (N_12750,N_11273,N_9226);
or U12751 (N_12751,N_10038,N_11418);
and U12752 (N_12752,N_11855,N_10998);
and U12753 (N_12753,N_9912,N_10469);
xor U12754 (N_12754,N_11978,N_9758);
nand U12755 (N_12755,N_11592,N_11054);
and U12756 (N_12756,N_10043,N_10466);
or U12757 (N_12757,N_10774,N_9727);
nand U12758 (N_12758,N_10239,N_10682);
and U12759 (N_12759,N_10308,N_9666);
nand U12760 (N_12760,N_11666,N_10615);
nor U12761 (N_12761,N_11307,N_11623);
or U12762 (N_12762,N_10226,N_10370);
nor U12763 (N_12763,N_10669,N_9604);
xor U12764 (N_12764,N_9444,N_11117);
nor U12765 (N_12765,N_11590,N_10900);
or U12766 (N_12766,N_11783,N_11991);
xnor U12767 (N_12767,N_10086,N_11963);
nand U12768 (N_12768,N_9082,N_10635);
nor U12769 (N_12769,N_10732,N_10907);
or U12770 (N_12770,N_10643,N_9198);
and U12771 (N_12771,N_11955,N_9134);
or U12772 (N_12772,N_9874,N_9423);
nand U12773 (N_12773,N_9388,N_9743);
nand U12774 (N_12774,N_11332,N_9187);
xor U12775 (N_12775,N_11566,N_11152);
nand U12776 (N_12776,N_10511,N_9506);
nand U12777 (N_12777,N_10983,N_10794);
nor U12778 (N_12778,N_10695,N_10311);
nand U12779 (N_12779,N_10127,N_10192);
or U12780 (N_12780,N_10068,N_11120);
or U12781 (N_12781,N_9826,N_11259);
nand U12782 (N_12782,N_10395,N_11836);
nor U12783 (N_12783,N_10339,N_11357);
or U12784 (N_12784,N_11811,N_11829);
or U12785 (N_12785,N_10024,N_9775);
nor U12786 (N_12786,N_9022,N_9610);
and U12787 (N_12787,N_10445,N_11320);
xnor U12788 (N_12788,N_11156,N_10332);
or U12789 (N_12789,N_10966,N_10566);
xnor U12790 (N_12790,N_10172,N_11401);
nand U12791 (N_12791,N_10020,N_11606);
and U12792 (N_12792,N_11533,N_11155);
nor U12793 (N_12793,N_9989,N_9465);
and U12794 (N_12794,N_10705,N_9654);
xor U12795 (N_12795,N_9944,N_9740);
nor U12796 (N_12796,N_10717,N_10269);
nand U12797 (N_12797,N_10065,N_10428);
nand U12798 (N_12798,N_11588,N_11056);
xor U12799 (N_12799,N_10053,N_11819);
nor U12800 (N_12800,N_11706,N_11122);
or U12801 (N_12801,N_10351,N_9219);
and U12802 (N_12802,N_10535,N_9114);
and U12803 (N_12803,N_11936,N_10087);
nand U12804 (N_12804,N_11236,N_9081);
xor U12805 (N_12805,N_10538,N_9080);
and U12806 (N_12806,N_11392,N_9746);
xnor U12807 (N_12807,N_9631,N_9897);
nand U12808 (N_12808,N_10075,N_9392);
and U12809 (N_12809,N_11950,N_10297);
nor U12810 (N_12810,N_10642,N_9014);
nand U12811 (N_12811,N_11612,N_11406);
and U12812 (N_12812,N_9652,N_11442);
or U12813 (N_12813,N_11639,N_10664);
nor U12814 (N_12814,N_9113,N_10961);
and U12815 (N_12815,N_9549,N_11209);
or U12816 (N_12816,N_10003,N_11805);
xnor U12817 (N_12817,N_11740,N_11295);
nand U12818 (N_12818,N_10409,N_11804);
or U12819 (N_12819,N_9281,N_10704);
or U12820 (N_12820,N_11447,N_10430);
nor U12821 (N_12821,N_9779,N_11820);
nor U12822 (N_12822,N_11079,N_10818);
nand U12823 (N_12823,N_11685,N_11160);
nor U12824 (N_12824,N_11481,N_11146);
or U12825 (N_12825,N_9839,N_9000);
nor U12826 (N_12826,N_11408,N_11736);
nor U12827 (N_12827,N_10826,N_10389);
or U12828 (N_12828,N_11058,N_10992);
nand U12829 (N_12829,N_9819,N_9408);
nor U12830 (N_12830,N_9157,N_9834);
nand U12831 (N_12831,N_10234,N_10676);
and U12832 (N_12832,N_11233,N_10433);
and U12833 (N_12833,N_9581,N_11432);
xnor U12834 (N_12834,N_9888,N_11380);
nor U12835 (N_12835,N_10808,N_9483);
nor U12836 (N_12836,N_10747,N_9323);
xnor U12837 (N_12837,N_9170,N_9648);
xnor U12838 (N_12838,N_10030,N_11189);
or U12839 (N_12839,N_10404,N_9879);
and U12840 (N_12840,N_11436,N_11240);
or U12841 (N_12841,N_11605,N_11887);
nand U12842 (N_12842,N_11013,N_9711);
xnor U12843 (N_12843,N_10233,N_9772);
nand U12844 (N_12844,N_9996,N_10159);
nor U12845 (N_12845,N_10689,N_10107);
xor U12846 (N_12846,N_9691,N_11049);
nor U12847 (N_12847,N_10655,N_11792);
nor U12848 (N_12848,N_10877,N_10196);
xnor U12849 (N_12849,N_11911,N_11007);
xnor U12850 (N_12850,N_11569,N_11142);
nand U12851 (N_12851,N_11848,N_9671);
xnor U12852 (N_12852,N_10508,N_11520);
and U12853 (N_12853,N_10379,N_9521);
xor U12854 (N_12854,N_11073,N_11921);
nor U12855 (N_12855,N_10777,N_9908);
nand U12856 (N_12856,N_11001,N_10911);
and U12857 (N_12857,N_11801,N_11231);
and U12858 (N_12858,N_11734,N_11699);
xnor U12859 (N_12859,N_10174,N_11235);
or U12860 (N_12860,N_9417,N_10666);
or U12861 (N_12861,N_10223,N_9252);
or U12862 (N_12862,N_11678,N_9975);
or U12863 (N_12863,N_10393,N_9716);
or U12864 (N_12864,N_11256,N_10727);
or U12865 (N_12865,N_9262,N_9862);
and U12866 (N_12866,N_9348,N_10309);
or U12867 (N_12867,N_10784,N_10541);
xnor U12868 (N_12868,N_10889,N_9602);
nor U12869 (N_12869,N_11837,N_9237);
xnor U12870 (N_12870,N_10202,N_10059);
and U12871 (N_12871,N_11686,N_11667);
or U12872 (N_12872,N_10034,N_9106);
xor U12873 (N_12873,N_10869,N_11431);
nor U12874 (N_12874,N_9770,N_9087);
xor U12875 (N_12875,N_10029,N_9089);
nor U12876 (N_12876,N_11204,N_11491);
and U12877 (N_12877,N_10368,N_10595);
xnor U12878 (N_12878,N_11113,N_9582);
nor U12879 (N_12879,N_9837,N_10591);
or U12880 (N_12880,N_11669,N_9622);
nor U12881 (N_12881,N_11147,N_11188);
nor U12882 (N_12882,N_10274,N_9222);
nand U12883 (N_12883,N_11985,N_11217);
and U12884 (N_12884,N_10602,N_9594);
nor U12885 (N_12885,N_9302,N_11221);
nand U12886 (N_12886,N_11387,N_9239);
nand U12887 (N_12887,N_9025,N_11070);
or U12888 (N_12888,N_9166,N_10120);
or U12889 (N_12889,N_11904,N_9881);
and U12890 (N_12890,N_11489,N_9886);
nor U12891 (N_12891,N_10337,N_10758);
nand U12892 (N_12892,N_9868,N_10719);
nor U12893 (N_12893,N_10149,N_9705);
or U12894 (N_12894,N_9931,N_9283);
and U12895 (N_12895,N_11354,N_9744);
or U12896 (N_12896,N_9036,N_10745);
xnor U12897 (N_12897,N_9902,N_10977);
xor U12898 (N_12898,N_10824,N_9866);
and U12899 (N_12899,N_9665,N_9778);
nand U12900 (N_12900,N_11745,N_9986);
or U12901 (N_12901,N_10683,N_9207);
nand U12902 (N_12902,N_11555,N_10850);
nand U12903 (N_12903,N_9260,N_10128);
xnor U12904 (N_12904,N_10169,N_11926);
nor U12905 (N_12905,N_11036,N_9774);
nand U12906 (N_12906,N_9153,N_10426);
or U12907 (N_12907,N_11665,N_9180);
nand U12908 (N_12908,N_9913,N_11711);
nor U12909 (N_12909,N_9700,N_10879);
nor U12910 (N_12910,N_9750,N_9942);
nor U12911 (N_12911,N_9710,N_11201);
xor U12912 (N_12912,N_10273,N_9531);
nand U12913 (N_12913,N_10820,N_11381);
nand U12914 (N_12914,N_10737,N_11340);
nor U12915 (N_12915,N_10649,N_10851);
nor U12916 (N_12916,N_11167,N_11986);
nand U12917 (N_12917,N_10097,N_10757);
nor U12918 (N_12918,N_11619,N_10424);
and U12919 (N_12919,N_11571,N_10630);
nand U12920 (N_12920,N_11611,N_9186);
or U12921 (N_12921,N_11664,N_9675);
nor U12922 (N_12922,N_10211,N_11483);
xnor U12923 (N_12923,N_10938,N_11199);
nand U12924 (N_12924,N_10927,N_11653);
xnor U12925 (N_12925,N_9818,N_11521);
nand U12926 (N_12926,N_10048,N_11696);
and U12927 (N_12927,N_11554,N_11536);
nand U12928 (N_12928,N_10318,N_9137);
nor U12929 (N_12929,N_10780,N_11247);
nor U12930 (N_12930,N_9326,N_11031);
nor U12931 (N_12931,N_11457,N_9398);
xnor U12932 (N_12932,N_11635,N_11644);
xnor U12933 (N_12933,N_9333,N_11139);
xor U12934 (N_12934,N_10123,N_10829);
nand U12935 (N_12935,N_9418,N_10673);
nand U12936 (N_12936,N_9116,N_11542);
nand U12937 (N_12937,N_11881,N_9707);
nor U12938 (N_12938,N_10115,N_10945);
xnor U12939 (N_12939,N_11906,N_10209);
or U12940 (N_12940,N_10289,N_10899);
nor U12941 (N_12941,N_10461,N_10898);
xor U12942 (N_12942,N_10575,N_11272);
or U12943 (N_12943,N_10588,N_9789);
nor U12944 (N_12944,N_9002,N_9756);
and U12945 (N_12945,N_11821,N_9527);
or U12946 (N_12946,N_9203,N_10255);
nand U12947 (N_12947,N_11500,N_9246);
and U12948 (N_12948,N_10182,N_11466);
and U12949 (N_12949,N_9663,N_11613);
nand U12950 (N_12950,N_9112,N_11933);
and U12951 (N_12951,N_11503,N_11009);
and U12952 (N_12952,N_9929,N_10797);
nor U12953 (N_12953,N_9300,N_9334);
nor U12954 (N_12954,N_9765,N_9751);
nor U12955 (N_12955,N_11738,N_10545);
or U12956 (N_12956,N_9199,N_11579);
xor U12957 (N_12957,N_11308,N_10054);
and U12958 (N_12958,N_9933,N_10281);
nand U12959 (N_12959,N_9853,N_9492);
nor U12960 (N_12960,N_10916,N_10185);
nor U12961 (N_12961,N_10594,N_11329);
or U12962 (N_12962,N_9452,N_11175);
nand U12963 (N_12963,N_9934,N_9349);
xor U12964 (N_12964,N_9052,N_10527);
nand U12965 (N_12965,N_10042,N_10114);
and U12966 (N_12966,N_10268,N_9185);
nor U12967 (N_12967,N_9372,N_10266);
nand U12968 (N_12968,N_11032,N_10620);
and U12969 (N_12969,N_11169,N_11293);
nand U12970 (N_12970,N_9893,N_11951);
nor U12971 (N_12971,N_10315,N_11487);
or U12972 (N_12972,N_9164,N_10335);
and U12973 (N_12973,N_11888,N_9194);
xor U12974 (N_12974,N_10557,N_10418);
or U12975 (N_12975,N_11407,N_11344);
nand U12976 (N_12976,N_9359,N_10964);
and U12977 (N_12977,N_11524,N_11020);
or U12978 (N_12978,N_9016,N_9406);
or U12979 (N_12979,N_10772,N_11698);
xor U12980 (N_12980,N_11274,N_11163);
xor U12981 (N_12981,N_10427,N_9798);
nand U12982 (N_12982,N_10709,N_11311);
xor U12983 (N_12983,N_11337,N_11080);
xor U12984 (N_12984,N_11338,N_11193);
xor U12985 (N_12985,N_10521,N_10085);
nand U12986 (N_12986,N_9192,N_9393);
or U12987 (N_12987,N_11267,N_10522);
nor U12988 (N_12988,N_11535,N_9451);
xnor U12989 (N_12989,N_10556,N_11704);
nand U12990 (N_12990,N_9491,N_11104);
or U12991 (N_12991,N_10103,N_10061);
or U12992 (N_12992,N_10324,N_9718);
or U12993 (N_12993,N_10146,N_11350);
or U12994 (N_12994,N_9938,N_10951);
nor U12995 (N_12995,N_10204,N_10569);
nand U12996 (N_12996,N_9026,N_10725);
nor U12997 (N_12997,N_10025,N_11538);
nand U12998 (N_12998,N_11224,N_11549);
nand U12999 (N_12999,N_9243,N_9269);
or U13000 (N_13000,N_10398,N_9431);
or U13001 (N_13001,N_9907,N_9032);
nor U13002 (N_13002,N_9712,N_11095);
xnor U13003 (N_13003,N_10160,N_9107);
and U13004 (N_13004,N_11279,N_9494);
nand U13005 (N_13005,N_10764,N_11111);
nor U13006 (N_13006,N_9193,N_9068);
nand U13007 (N_13007,N_11294,N_10680);
or U13008 (N_13008,N_9612,N_10104);
nand U13009 (N_13009,N_9053,N_9747);
or U13010 (N_13010,N_11827,N_10164);
or U13011 (N_13011,N_11445,N_9425);
nor U13012 (N_13012,N_9018,N_11265);
nand U13013 (N_13013,N_9682,N_9949);
and U13014 (N_13014,N_9799,N_9606);
xnor U13015 (N_13015,N_11540,N_9684);
nor U13016 (N_13016,N_10623,N_9076);
and U13017 (N_13017,N_11433,N_10821);
and U13018 (N_13018,N_9256,N_9573);
xnor U13019 (N_13019,N_10882,N_9475);
xor U13020 (N_13020,N_9681,N_10561);
and U13021 (N_13021,N_10559,N_10738);
and U13022 (N_13022,N_10867,N_9561);
xnor U13023 (N_13023,N_9267,N_9620);
and U13024 (N_13024,N_10472,N_11862);
or U13025 (N_13025,N_10999,N_10639);
nand U13026 (N_13026,N_10650,N_11021);
nand U13027 (N_13027,N_11983,N_9894);
nor U13028 (N_13028,N_11617,N_11851);
nand U13029 (N_13029,N_9793,N_10734);
xor U13030 (N_13030,N_9343,N_10832);
xnor U13031 (N_13031,N_11545,N_10181);
and U13032 (N_13032,N_11764,N_9562);
nor U13033 (N_13033,N_9715,N_10975);
nand U13034 (N_13034,N_9589,N_11850);
or U13035 (N_13035,N_9373,N_10654);
or U13036 (N_13036,N_9210,N_10470);
or U13037 (N_13037,N_10158,N_11853);
nand U13038 (N_13038,N_11788,N_9069);
and U13039 (N_13039,N_10023,N_10478);
or U13040 (N_13040,N_11660,N_11532);
nor U13041 (N_13041,N_11504,N_10853);
xor U13042 (N_13042,N_11153,N_11161);
nor U13043 (N_13043,N_11942,N_9702);
or U13044 (N_13044,N_11124,N_9865);
and U13045 (N_13045,N_9584,N_9781);
xor U13046 (N_13046,N_9680,N_11090);
xnor U13047 (N_13047,N_9687,N_10263);
and U13048 (N_13048,N_10316,N_11321);
and U13049 (N_13049,N_11762,N_10849);
nand U13050 (N_13050,N_9006,N_11228);
nand U13051 (N_13051,N_9163,N_11239);
nor U13052 (N_13052,N_9854,N_9538);
and U13053 (N_13053,N_9978,N_11376);
nor U13054 (N_13054,N_9150,N_11422);
nor U13055 (N_13055,N_10904,N_11979);
and U13056 (N_13056,N_10840,N_11424);
or U13057 (N_13057,N_9763,N_11975);
nor U13058 (N_13058,N_9972,N_10161);
or U13059 (N_13059,N_10796,N_10217);
nand U13060 (N_13060,N_10066,N_10681);
nor U13061 (N_13061,N_9496,N_11728);
nand U13062 (N_13062,N_9467,N_9394);
and U13063 (N_13063,N_10028,N_9832);
xor U13064 (N_13064,N_11499,N_10031);
or U13065 (N_13065,N_9593,N_11482);
nand U13066 (N_13066,N_10434,N_9007);
and U13067 (N_13067,N_10264,N_10230);
nor U13068 (N_13068,N_10347,N_9966);
nor U13069 (N_13069,N_10564,N_9723);
and U13070 (N_13070,N_10637,N_9841);
and U13071 (N_13071,N_9065,N_10078);
xnor U13072 (N_13072,N_11716,N_9800);
nor U13073 (N_13073,N_10924,N_11151);
and U13074 (N_13074,N_11649,N_11793);
or U13075 (N_13075,N_11958,N_11260);
or U13076 (N_13076,N_11732,N_9970);
nor U13077 (N_13077,N_10007,N_9732);
or U13078 (N_13078,N_10294,N_10341);
nor U13079 (N_13079,N_9156,N_9526);
nand U13080 (N_13080,N_11218,N_10454);
nand U13081 (N_13081,N_9159,N_9321);
nand U13082 (N_13082,N_9672,N_9539);
nand U13083 (N_13083,N_11818,N_9587);
nor U13084 (N_13084,N_9367,N_9830);
or U13085 (N_13085,N_9695,N_10135);
nor U13086 (N_13086,N_10795,N_9522);
and U13087 (N_13087,N_11895,N_10489);
nand U13088 (N_13088,N_9699,N_9525);
nand U13089 (N_13089,N_11832,N_9201);
xor U13090 (N_13090,N_11972,N_11797);
nand U13091 (N_13091,N_10672,N_10819);
xor U13092 (N_13092,N_11648,N_9420);
or U13093 (N_13093,N_11409,N_11860);
nand U13094 (N_13094,N_10359,N_10142);
nand U13095 (N_13095,N_10711,N_10476);
nand U13096 (N_13096,N_9608,N_9075);
nor U13097 (N_13097,N_9510,N_10861);
xor U13098 (N_13098,N_11194,N_11610);
xnor U13099 (N_13099,N_10657,N_11831);
nor U13100 (N_13100,N_9265,N_11190);
xnor U13101 (N_13101,N_9801,N_9963);
xor U13102 (N_13102,N_10985,N_9807);
nor U13103 (N_13103,N_9910,N_9534);
and U13104 (N_13104,N_11346,N_10626);
xor U13105 (N_13105,N_9195,N_10816);
nor U13106 (N_13106,N_10092,N_10377);
or U13107 (N_13107,N_9407,N_9482);
nor U13108 (N_13108,N_10504,N_10386);
or U13109 (N_13109,N_10134,N_10343);
or U13110 (N_13110,N_11940,N_11946);
xor U13111 (N_13111,N_10199,N_9755);
nor U13112 (N_13112,N_11006,N_11121);
nand U13113 (N_13113,N_9502,N_10969);
nand U13114 (N_13114,N_10366,N_11296);
xnor U13115 (N_13115,N_11005,N_10173);
nand U13116 (N_13116,N_11931,N_9646);
xnor U13117 (N_13117,N_11469,N_11662);
nand U13118 (N_13118,N_11559,N_10401);
and U13119 (N_13119,N_9898,N_11629);
nor U13120 (N_13120,N_11670,N_11694);
or U13121 (N_13121,N_9692,N_11630);
nor U13122 (N_13122,N_11550,N_11215);
and U13123 (N_13123,N_9063,N_11052);
nor U13124 (N_13124,N_11982,N_11596);
and U13125 (N_13125,N_10352,N_10131);
or U13126 (N_13126,N_9926,N_11580);
nor U13127 (N_13127,N_9757,N_9413);
nand U13128 (N_13128,N_11961,N_11802);
or U13129 (N_13129,N_9804,N_10187);
or U13130 (N_13130,N_9601,N_10823);
or U13131 (N_13131,N_10895,N_10847);
and U13132 (N_13132,N_9590,N_9385);
and U13133 (N_13133,N_10468,N_9817);
or U13134 (N_13134,N_11154,N_10304);
nor U13135 (N_13135,N_9356,N_9335);
nand U13136 (N_13136,N_10632,N_11787);
xor U13137 (N_13137,N_9958,N_11852);
or U13138 (N_13138,N_10959,N_11386);
and U13139 (N_13139,N_11448,N_9753);
nand U13140 (N_13140,N_11683,N_9072);
xnor U13141 (N_13141,N_10036,N_11844);
nor U13142 (N_13142,N_10503,N_10259);
nor U13143 (N_13143,N_9683,N_11108);
xor U13144 (N_13144,N_10372,N_9140);
or U13145 (N_13145,N_9241,N_9382);
or U13146 (N_13146,N_9657,N_9059);
nand U13147 (N_13147,N_9310,N_11356);
xnor U13148 (N_13148,N_9248,N_9277);
nand U13149 (N_13149,N_10592,N_9873);
nor U13150 (N_13150,N_10872,N_9027);
or U13151 (N_13151,N_10674,N_11574);
nand U13152 (N_13152,N_9585,N_9791);
nand U13153 (N_13153,N_9967,N_11781);
or U13154 (N_13154,N_11724,N_9617);
xnor U13155 (N_13155,N_11534,N_9305);
and U13156 (N_13156,N_9145,N_9634);
or U13157 (N_13157,N_10307,N_11861);
and U13158 (N_13158,N_9462,N_11902);
xor U13159 (N_13159,N_11527,N_9208);
xor U13160 (N_13160,N_9121,N_9497);
and U13161 (N_13161,N_11814,N_11568);
or U13162 (N_13162,N_9628,N_11101);
or U13163 (N_13163,N_10457,N_10675);
and U13164 (N_13164,N_9136,N_9189);
and U13165 (N_13165,N_9162,N_10170);
and U13166 (N_13166,N_9624,N_10006);
nor U13167 (N_13167,N_9882,N_9579);
and U13168 (N_13168,N_9139,N_10275);
nand U13169 (N_13169,N_9410,N_10117);
nand U13170 (N_13170,N_9205,N_11000);
or U13171 (N_13171,N_10515,N_11510);
nor U13172 (N_13172,N_11044,N_10880);
xor U13173 (N_13173,N_10540,N_9441);
nand U13174 (N_13174,N_11046,N_11379);
and U13175 (N_13175,N_11710,N_10776);
or U13176 (N_13176,N_11241,N_11913);
nor U13177 (N_13177,N_9979,N_10744);
and U13178 (N_13178,N_10148,N_10171);
nand U13179 (N_13179,N_10886,N_9279);
xnor U13180 (N_13180,N_9102,N_11132);
or U13181 (N_13181,N_10495,N_9179);
xnor U13182 (N_13182,N_11150,N_10756);
xnor U13183 (N_13183,N_11064,N_9749);
nor U13184 (N_13184,N_11593,N_9639);
nand U13185 (N_13185,N_10568,N_9638);
nor U13186 (N_13186,N_11174,N_9191);
or U13187 (N_13187,N_10390,N_11484);
xor U13188 (N_13188,N_9146,N_11463);
nor U13189 (N_13189,N_10291,N_9555);
nor U13190 (N_13190,N_10258,N_9353);
xor U13191 (N_13191,N_9307,N_11709);
or U13192 (N_13192,N_11257,N_10765);
xor U13193 (N_13193,N_11643,N_11179);
or U13194 (N_13194,N_11587,N_10088);
or U13195 (N_13195,N_10490,N_9984);
or U13196 (N_13196,N_11411,N_10257);
nor U13197 (N_13197,N_11066,N_9877);
nor U13198 (N_13198,N_10108,N_11531);
or U13199 (N_13199,N_11172,N_9110);
nor U13200 (N_13200,N_10815,N_9374);
xor U13201 (N_13201,N_11358,N_10188);
xor U13202 (N_13202,N_11567,N_11452);
or U13203 (N_13203,N_10084,N_9829);
nand U13204 (N_13204,N_9061,N_10752);
xor U13205 (N_13205,N_11782,N_9316);
or U13206 (N_13206,N_11226,N_9843);
nor U13207 (N_13207,N_11994,N_10336);
or U13208 (N_13208,N_10884,N_10201);
nand U13209 (N_13209,N_9685,N_9105);
or U13210 (N_13210,N_11614,N_10712);
and U13211 (N_13211,N_9403,N_9426);
or U13212 (N_13212,N_9558,N_9254);
nand U13213 (N_13213,N_9869,N_11323);
nand U13214 (N_13214,N_9660,N_9312);
or U13215 (N_13215,N_9457,N_9126);
xor U13216 (N_13216,N_10321,N_10121);
nor U13217 (N_13217,N_10984,N_11561);
nand U13218 (N_13218,N_10125,N_10937);
xor U13219 (N_13219,N_11843,N_10989);
nand U13220 (N_13220,N_9577,N_11708);
and U13221 (N_13221,N_9733,N_9456);
nand U13222 (N_13222,N_10692,N_11760);
xnor U13223 (N_13223,N_11552,N_9284);
xnor U13224 (N_13224,N_10934,N_10552);
nor U13225 (N_13225,N_10627,N_11158);
and U13226 (N_13226,N_10252,N_11516);
nor U13227 (N_13227,N_10662,N_10403);
xnor U13228 (N_13228,N_10834,N_11028);
xor U13229 (N_13229,N_11403,N_10670);
nor U13230 (N_13230,N_9171,N_9844);
xor U13231 (N_13231,N_9905,N_9115);
nor U13232 (N_13232,N_9985,N_9884);
or U13233 (N_13233,N_11741,N_9635);
nand U13234 (N_13234,N_10891,N_10955);
nand U13235 (N_13235,N_9790,N_11868);
or U13236 (N_13236,N_11897,N_11765);
xor U13237 (N_13237,N_10180,N_9144);
xnor U13238 (N_13238,N_9268,N_10856);
xnor U13239 (N_13239,N_11416,N_10122);
nand U13240 (N_13240,N_10875,N_10931);
nand U13241 (N_13241,N_11458,N_11099);
nor U13242 (N_13242,N_11854,N_10957);
nor U13243 (N_13243,N_11040,N_11027);
nor U13244 (N_13244,N_9221,N_10340);
and U13245 (N_13245,N_10968,N_11026);
xor U13246 (N_13246,N_9292,N_11742);
and U13247 (N_13247,N_10656,N_11509);
and U13248 (N_13248,N_10735,N_11425);
nor U13249 (N_13249,N_10111,N_9725);
or U13250 (N_13250,N_11519,N_10002);
xnor U13251 (N_13251,N_10513,N_11251);
nand U13252 (N_13252,N_11195,N_10929);
nand U13253 (N_13253,N_10859,N_11319);
nand U13254 (N_13254,N_11654,N_11334);
nor U13255 (N_13255,N_9399,N_9788);
or U13256 (N_13256,N_9480,N_11551);
xor U13257 (N_13257,N_9669,N_9278);
or U13258 (N_13258,N_9875,N_10746);
or U13259 (N_13259,N_9923,N_11899);
nor U13260 (N_13260,N_9155,N_11492);
nor U13261 (N_13261,N_10186,N_10100);
xnor U13262 (N_13262,N_9838,N_10708);
xnor U13263 (N_13263,N_10549,N_10550);
and U13264 (N_13264,N_9111,N_9386);
and U13265 (N_13265,N_11841,N_10616);
xnor U13266 (N_13266,N_11651,N_9471);
xnor U13267 (N_13267,N_9331,N_10854);
nor U13268 (N_13268,N_10548,N_9997);
xnor U13269 (N_13269,N_10554,N_9383);
nor U13270 (N_13270,N_9235,N_9148);
and U13271 (N_13271,N_11900,N_11366);
nand U13272 (N_13272,N_9935,N_9340);
nor U13273 (N_13273,N_11679,N_9468);
or U13274 (N_13274,N_10193,N_9661);
nor U13275 (N_13275,N_11285,N_10243);
and U13276 (N_13276,N_9311,N_9342);
or U13277 (N_13277,N_10000,N_9859);
or U13278 (N_13278,N_9911,N_11060);
and U13279 (N_13279,N_10397,N_11444);
and U13280 (N_13280,N_10593,N_10509);
xor U13281 (N_13281,N_10051,N_9729);
or U13282 (N_13282,N_10976,N_11045);
xor U13283 (N_13283,N_10388,N_10878);
and U13284 (N_13284,N_11494,N_10344);
and U13285 (N_13285,N_10219,N_10464);
nor U13286 (N_13286,N_11486,N_11219);
nand U13287 (N_13287,N_11599,N_11886);
or U13288 (N_13288,N_11772,N_11725);
and U13289 (N_13289,N_10963,N_11192);
and U13290 (N_13290,N_10991,N_10141);
or U13291 (N_13291,N_10881,N_9011);
nand U13292 (N_13292,N_11835,N_11304);
or U13293 (N_13293,N_10447,N_9289);
nand U13294 (N_13294,N_9332,N_9315);
xor U13295 (N_13295,N_10739,N_11828);
nand U13296 (N_13296,N_11207,N_9927);
xnor U13297 (N_13297,N_9261,N_10838);
or U13298 (N_13298,N_9493,N_10361);
nand U13299 (N_13299,N_10176,N_10405);
and U13300 (N_13300,N_11248,N_10519);
nor U13301 (N_13301,N_11514,N_9432);
nand U13302 (N_13302,N_11809,N_9013);
nand U13303 (N_13303,N_11761,N_9078);
or U13304 (N_13304,N_9917,N_11472);
nand U13305 (N_13305,N_11391,N_11351);
or U13306 (N_13306,N_9649,N_11493);
xnor U13307 (N_13307,N_11035,N_11335);
nor U13308 (N_13308,N_10216,N_10842);
xnor U13309 (N_13309,N_9358,N_9290);
and U13310 (N_13310,N_10179,N_11846);
xor U13311 (N_13311,N_9962,N_10753);
nor U13312 (N_13312,N_10152,N_9948);
or U13313 (N_13313,N_10014,N_9667);
or U13314 (N_13314,N_9387,N_9645);
nand U13315 (N_13315,N_9258,N_9600);
nor U13316 (N_13316,N_11373,N_9147);
or U13317 (N_13317,N_11014,N_10394);
and U13318 (N_13318,N_11170,N_11891);
nor U13319 (N_13319,N_10646,N_10697);
xnor U13320 (N_13320,N_10619,N_9401);
and U13321 (N_13321,N_9361,N_10791);
and U13322 (N_13322,N_11632,N_9848);
or U13323 (N_13323,N_9109,N_9135);
and U13324 (N_13324,N_9229,N_10506);
nand U13325 (N_13325,N_11343,N_11794);
xnor U13326 (N_13326,N_11790,N_9537);
or U13327 (N_13327,N_11954,N_9091);
xnor U13328 (N_13328,N_10140,N_10027);
or U13329 (N_13329,N_9550,N_10920);
nand U13330 (N_13330,N_10387,N_9714);
nand U13331 (N_13331,N_9782,N_10417);
nor U13332 (N_13332,N_11468,N_10184);
nor U13333 (N_13333,N_11867,N_9776);
and U13334 (N_13334,N_11434,N_10376);
and U13335 (N_13335,N_11415,N_11276);
and U13336 (N_13336,N_10338,N_11786);
nand U13337 (N_13337,N_11583,N_10412);
and U13338 (N_13338,N_9232,N_10908);
xor U13339 (N_13339,N_9346,N_10781);
nor U13340 (N_13340,N_10452,N_10800);
and U13341 (N_13341,N_9376,N_11360);
or U13342 (N_13342,N_11543,N_9575);
and U13343 (N_13343,N_9728,N_10755);
and U13344 (N_13344,N_10328,N_11185);
and U13345 (N_13345,N_11687,N_11460);
xor U13346 (N_13346,N_10013,N_10453);
and U13347 (N_13347,N_9794,N_11905);
nor U13348 (N_13348,N_9117,N_11417);
and U13349 (N_13349,N_9906,N_9568);
nand U13350 (N_13350,N_9919,N_11941);
xor U13351 (N_13351,N_11758,N_10806);
nand U13352 (N_13352,N_9540,N_10835);
nor U13353 (N_13353,N_9308,N_9010);
nor U13354 (N_13354,N_10779,N_11957);
or U13355 (N_13355,N_10278,N_9085);
and U13356 (N_13356,N_11093,N_9551);
or U13357 (N_13357,N_11791,N_10250);
nor U13358 (N_13358,N_10799,N_11713);
and U13359 (N_13359,N_10982,N_9509);
nand U13360 (N_13360,N_10792,N_10855);
and U13361 (N_13361,N_10699,N_9722);
nand U13362 (N_13362,N_11410,N_11180);
nor U13363 (N_13363,N_10056,N_9903);
or U13364 (N_13364,N_9596,N_9280);
nand U13365 (N_13365,N_11876,N_11262);
nor U13366 (N_13366,N_9250,N_11912);
xnor U13367 (N_13367,N_9320,N_11869);
and U13368 (N_13368,N_9217,N_10512);
xor U13369 (N_13369,N_9272,N_10980);
or U13370 (N_13370,N_11693,N_10045);
nor U13371 (N_13371,N_9706,N_11748);
and U13372 (N_13372,N_11011,N_11628);
nor U13373 (N_13373,N_10589,N_10284);
xor U13374 (N_13374,N_9038,N_11072);
or U13375 (N_13375,N_11769,N_9637);
xnor U13376 (N_13376,N_11449,N_11371);
nor U13377 (N_13377,N_10950,N_10189);
nand U13378 (N_13378,N_9932,N_10285);
or U13379 (N_13379,N_10986,N_10885);
xor U13380 (N_13380,N_9206,N_9731);
or U13381 (N_13381,N_10322,N_10868);
and U13382 (N_13382,N_11038,N_11023);
nand U13383 (N_13383,N_9142,N_9543);
and U13384 (N_13384,N_9571,N_10276);
or U13385 (N_13385,N_11565,N_11383);
nor U13386 (N_13386,N_9803,N_11266);
and U13387 (N_13387,N_9524,N_11074);
and U13388 (N_13388,N_11810,N_11977);
nor U13389 (N_13389,N_10496,N_10411);
xnor U13390 (N_13390,N_10803,N_10306);
or U13391 (N_13391,N_10517,N_10089);
and U13392 (N_13392,N_9786,N_11600);
and U13393 (N_13393,N_11752,N_11097);
nand U13394 (N_13394,N_9719,N_11799);
nand U13395 (N_13395,N_9971,N_10775);
xor U13396 (N_13396,N_11833,N_9767);
nor U13397 (N_13397,N_9498,N_9443);
nand U13398 (N_13398,N_9896,N_9257);
and U13399 (N_13399,N_10280,N_10203);
or U13400 (N_13400,N_11615,N_11692);
nor U13401 (N_13401,N_10323,N_10113);
nand U13402 (N_13402,N_11016,N_11995);
or U13403 (N_13403,N_10283,N_11324);
nand U13404 (N_13404,N_9858,N_11815);
nand U13405 (N_13405,N_11370,N_9056);
nor U13406 (N_13406,N_11348,N_9128);
nand U13407 (N_13407,N_11557,N_11971);
nand U13408 (N_13408,N_9825,N_9124);
or U13409 (N_13409,N_10477,N_11661);
or U13410 (N_13410,N_10109,N_11939);
nor U13411 (N_13411,N_9060,N_9846);
nor U13412 (N_13412,N_9484,N_11475);
nor U13413 (N_13413,N_9472,N_9836);
and U13414 (N_13414,N_9360,N_10974);
xor U13415 (N_13415,N_10305,N_10474);
xnor U13416 (N_13416,N_10629,N_9591);
nor U13417 (N_13417,N_9161,N_10228);
or U13418 (N_13418,N_10926,N_10096);
xor U13419 (N_13419,N_9440,N_10357);
and U13420 (N_13420,N_9943,N_10958);
nor U13421 (N_13421,N_10701,N_10598);
nor U13422 (N_13422,N_10578,N_9993);
or U13423 (N_13423,N_11807,N_9469);
or U13424 (N_13424,N_9454,N_10585);
xnor U13425 (N_13425,N_9633,N_11298);
nand U13426 (N_13426,N_9945,N_9535);
and U13427 (N_13427,N_9773,N_10195);
nand U13428 (N_13428,N_9378,N_11609);
xnor U13429 (N_13429,N_10570,N_10703);
and U13430 (N_13430,N_11098,N_11727);
or U13431 (N_13431,N_11166,N_11115);
nor U13432 (N_13432,N_10608,N_9548);
xor U13433 (N_13433,N_10163,N_10380);
nor U13434 (N_13434,N_10207,N_11420);
nand U13435 (N_13435,N_9717,N_11771);
nand U13436 (N_13436,N_10763,N_11277);
xnor U13437 (N_13437,N_11479,N_9516);
or U13438 (N_13438,N_10396,N_11243);
nor U13439 (N_13439,N_10355,N_10653);
and U13440 (N_13440,N_10360,N_9319);
xor U13441 (N_13441,N_11856,N_9396);
and U13442 (N_13442,N_10542,N_11655);
and U13443 (N_13443,N_11368,N_11082);
nand U13444 (N_13444,N_10415,N_10584);
xnor U13445 (N_13445,N_10118,N_10787);
or U13446 (N_13446,N_11894,N_11564);
or U13447 (N_13447,N_9900,N_9736);
xor U13448 (N_13448,N_10583,N_9947);
nor U13449 (N_13449,N_10553,N_11916);
or U13450 (N_13450,N_9079,N_10848);
nor U13451 (N_13451,N_10831,N_9362);
or U13452 (N_13452,N_10009,N_11526);
xor U13453 (N_13453,N_9108,N_11620);
nor U13454 (N_13454,N_11652,N_11990);
or U13455 (N_13455,N_9677,N_9412);
and U13456 (N_13456,N_11213,N_11882);
and U13457 (N_13457,N_10313,N_9197);
or U13458 (N_13458,N_11636,N_11722);
and U13459 (N_13459,N_10941,N_9574);
nand U13460 (N_13460,N_9453,N_11461);
nand U13461 (N_13461,N_11541,N_11880);
nand U13462 (N_13462,N_9130,N_10101);
and U13463 (N_13463,N_11857,N_9572);
nand U13464 (N_13464,N_11515,N_11582);
nor U13465 (N_13465,N_11089,N_11255);
or U13466 (N_13466,N_11187,N_9785);
and U13467 (N_13467,N_11839,N_10833);
xnor U13468 (N_13468,N_10391,N_9636);
nand U13469 (N_13469,N_11715,N_11863);
nor U13470 (N_13470,N_11470,N_11608);
nand U13471 (N_13471,N_11473,N_11618);
or U13472 (N_13472,N_11674,N_11640);
xor U13473 (N_13473,N_11878,N_9735);
or U13474 (N_13474,N_11813,N_11453);
nand U13475 (N_13475,N_11467,N_11305);
nand U13476 (N_13476,N_11838,N_11647);
or U13477 (N_13477,N_9552,N_9347);
xnor U13478 (N_13478,N_11705,N_10601);
xor U13479 (N_13479,N_9352,N_9994);
nand U13480 (N_13480,N_9438,N_11650);
xnor U13481 (N_13481,N_11330,N_9042);
or U13482 (N_13482,N_11924,N_10479);
nor U13483 (N_13483,N_9954,N_11094);
xnor U13484 (N_13484,N_9481,N_9070);
or U13485 (N_13485,N_9303,N_9379);
nor U13486 (N_13486,N_10463,N_9867);
and U13487 (N_13487,N_9071,N_11830);
and U13488 (N_13488,N_9796,N_9576);
nand U13489 (N_13489,N_11427,N_9904);
or U13490 (N_13490,N_10016,N_10004);
xor U13491 (N_13491,N_11953,N_9377);
xor U13492 (N_13492,N_10231,N_10126);
nor U13493 (N_13493,N_9547,N_11517);
xor U13494 (N_13494,N_9084,N_10432);
or U13495 (N_13495,N_9768,N_10058);
or U13496 (N_13496,N_9713,N_10314);
and U13497 (N_13497,N_11002,N_9720);
nand U13498 (N_13498,N_9093,N_9211);
nor U13499 (N_13499,N_11286,N_10749);
or U13500 (N_13500,N_11910,N_10865);
xnor U13501 (N_13501,N_11174,N_10704);
or U13502 (N_13502,N_11378,N_9595);
xor U13503 (N_13503,N_9152,N_11585);
nand U13504 (N_13504,N_10355,N_11269);
nor U13505 (N_13505,N_9395,N_9935);
or U13506 (N_13506,N_10229,N_11496);
xor U13507 (N_13507,N_11542,N_10805);
or U13508 (N_13508,N_10347,N_11746);
or U13509 (N_13509,N_11415,N_9289);
or U13510 (N_13510,N_9765,N_10643);
nand U13511 (N_13511,N_11678,N_10839);
or U13512 (N_13512,N_9191,N_9038);
nand U13513 (N_13513,N_9980,N_11563);
or U13514 (N_13514,N_10126,N_11373);
or U13515 (N_13515,N_10450,N_11609);
nor U13516 (N_13516,N_11392,N_10557);
and U13517 (N_13517,N_9133,N_10552);
nor U13518 (N_13518,N_9988,N_10435);
nor U13519 (N_13519,N_9026,N_10944);
and U13520 (N_13520,N_11080,N_10707);
xnor U13521 (N_13521,N_10125,N_11883);
nand U13522 (N_13522,N_9655,N_11113);
or U13523 (N_13523,N_10428,N_11142);
xnor U13524 (N_13524,N_11254,N_11056);
nor U13525 (N_13525,N_11703,N_11651);
nand U13526 (N_13526,N_9920,N_9307);
nand U13527 (N_13527,N_9921,N_11763);
nor U13528 (N_13528,N_10167,N_10772);
xor U13529 (N_13529,N_9405,N_10301);
and U13530 (N_13530,N_9851,N_11936);
xor U13531 (N_13531,N_9785,N_11974);
or U13532 (N_13532,N_9483,N_9488);
and U13533 (N_13533,N_9182,N_10990);
nand U13534 (N_13534,N_9497,N_9722);
xnor U13535 (N_13535,N_10104,N_10614);
nand U13536 (N_13536,N_10598,N_9251);
and U13537 (N_13537,N_11208,N_9522);
and U13538 (N_13538,N_9582,N_9014);
and U13539 (N_13539,N_11105,N_9498);
nand U13540 (N_13540,N_11353,N_10294);
or U13541 (N_13541,N_9701,N_11565);
or U13542 (N_13542,N_9471,N_11153);
xnor U13543 (N_13543,N_10751,N_9590);
or U13544 (N_13544,N_11477,N_11039);
or U13545 (N_13545,N_10236,N_11567);
and U13546 (N_13546,N_10487,N_11459);
or U13547 (N_13547,N_10296,N_11304);
nand U13548 (N_13548,N_9086,N_9031);
nand U13549 (N_13549,N_10863,N_11526);
or U13550 (N_13550,N_9989,N_9466);
or U13551 (N_13551,N_9026,N_9485);
and U13552 (N_13552,N_9405,N_10151);
nand U13553 (N_13553,N_9224,N_10503);
and U13554 (N_13554,N_10679,N_9595);
nor U13555 (N_13555,N_10456,N_9843);
or U13556 (N_13556,N_10818,N_9265);
xnor U13557 (N_13557,N_10907,N_10778);
nor U13558 (N_13558,N_11953,N_11102);
and U13559 (N_13559,N_11734,N_10818);
and U13560 (N_13560,N_9550,N_11299);
and U13561 (N_13561,N_9471,N_9311);
nand U13562 (N_13562,N_11373,N_10657);
and U13563 (N_13563,N_10384,N_11085);
or U13564 (N_13564,N_9026,N_10680);
xnor U13565 (N_13565,N_9062,N_10669);
or U13566 (N_13566,N_9499,N_9053);
nand U13567 (N_13567,N_11654,N_9321);
nor U13568 (N_13568,N_10747,N_10804);
nor U13569 (N_13569,N_9043,N_9233);
and U13570 (N_13570,N_10297,N_10079);
nand U13571 (N_13571,N_10879,N_11983);
and U13572 (N_13572,N_11098,N_9757);
xor U13573 (N_13573,N_11549,N_9399);
or U13574 (N_13574,N_9219,N_9335);
nand U13575 (N_13575,N_11372,N_10789);
nand U13576 (N_13576,N_11135,N_10838);
and U13577 (N_13577,N_10127,N_11022);
xnor U13578 (N_13578,N_11834,N_10380);
xor U13579 (N_13579,N_10977,N_10256);
nand U13580 (N_13580,N_9668,N_11099);
xor U13581 (N_13581,N_9898,N_10034);
and U13582 (N_13582,N_10142,N_9297);
nor U13583 (N_13583,N_10064,N_9616);
and U13584 (N_13584,N_9357,N_10384);
nor U13585 (N_13585,N_10296,N_10631);
or U13586 (N_13586,N_9294,N_10072);
or U13587 (N_13587,N_11744,N_11875);
nor U13588 (N_13588,N_10523,N_11330);
or U13589 (N_13589,N_9333,N_10037);
xnor U13590 (N_13590,N_10510,N_9886);
or U13591 (N_13591,N_11262,N_11376);
and U13592 (N_13592,N_10776,N_9080);
or U13593 (N_13593,N_9238,N_10825);
nor U13594 (N_13594,N_9216,N_11292);
nor U13595 (N_13595,N_11576,N_11967);
xnor U13596 (N_13596,N_9703,N_9592);
and U13597 (N_13597,N_10848,N_11916);
and U13598 (N_13598,N_9803,N_11690);
xor U13599 (N_13599,N_10218,N_9462);
xor U13600 (N_13600,N_11206,N_9222);
xor U13601 (N_13601,N_11565,N_11567);
and U13602 (N_13602,N_9877,N_11852);
or U13603 (N_13603,N_9958,N_11648);
xor U13604 (N_13604,N_11959,N_10428);
and U13605 (N_13605,N_11980,N_9722);
and U13606 (N_13606,N_11639,N_9118);
and U13607 (N_13607,N_10320,N_9009);
nand U13608 (N_13608,N_11953,N_9361);
nor U13609 (N_13609,N_11011,N_11576);
nand U13610 (N_13610,N_10365,N_10078);
or U13611 (N_13611,N_9116,N_9694);
nor U13612 (N_13612,N_10061,N_9978);
xor U13613 (N_13613,N_11430,N_11260);
nand U13614 (N_13614,N_11894,N_11532);
or U13615 (N_13615,N_9554,N_11640);
and U13616 (N_13616,N_9191,N_10508);
xor U13617 (N_13617,N_10299,N_11319);
or U13618 (N_13618,N_10396,N_9896);
nor U13619 (N_13619,N_9177,N_11643);
xor U13620 (N_13620,N_10735,N_9663);
or U13621 (N_13621,N_10083,N_10958);
nor U13622 (N_13622,N_9516,N_11342);
xor U13623 (N_13623,N_10616,N_10673);
or U13624 (N_13624,N_9974,N_11527);
and U13625 (N_13625,N_11550,N_11369);
nor U13626 (N_13626,N_9845,N_10273);
and U13627 (N_13627,N_10171,N_11102);
and U13628 (N_13628,N_11671,N_11733);
nor U13629 (N_13629,N_11856,N_10495);
or U13630 (N_13630,N_10854,N_11721);
nand U13631 (N_13631,N_10212,N_11694);
nor U13632 (N_13632,N_9790,N_11156);
nor U13633 (N_13633,N_9552,N_9531);
nor U13634 (N_13634,N_11929,N_9336);
nand U13635 (N_13635,N_9385,N_11383);
nand U13636 (N_13636,N_11508,N_11736);
nor U13637 (N_13637,N_11792,N_9862);
nand U13638 (N_13638,N_10099,N_11525);
or U13639 (N_13639,N_11250,N_9061);
xnor U13640 (N_13640,N_10668,N_9630);
nor U13641 (N_13641,N_11935,N_10968);
or U13642 (N_13642,N_11439,N_9133);
or U13643 (N_13643,N_11073,N_11315);
xor U13644 (N_13644,N_9288,N_9540);
xnor U13645 (N_13645,N_11384,N_11194);
nand U13646 (N_13646,N_10249,N_11616);
nor U13647 (N_13647,N_10020,N_11731);
xnor U13648 (N_13648,N_10958,N_11787);
xor U13649 (N_13649,N_9495,N_9051);
or U13650 (N_13650,N_10640,N_9792);
or U13651 (N_13651,N_9796,N_11714);
and U13652 (N_13652,N_11668,N_10578);
and U13653 (N_13653,N_11766,N_10314);
xnor U13654 (N_13654,N_9089,N_10633);
nor U13655 (N_13655,N_10288,N_10694);
or U13656 (N_13656,N_9617,N_11156);
nand U13657 (N_13657,N_10343,N_10950);
nand U13658 (N_13658,N_11721,N_11570);
nor U13659 (N_13659,N_9298,N_11591);
and U13660 (N_13660,N_11685,N_11202);
xor U13661 (N_13661,N_9322,N_11551);
or U13662 (N_13662,N_11372,N_11095);
nor U13663 (N_13663,N_11226,N_10485);
and U13664 (N_13664,N_10712,N_10413);
or U13665 (N_13665,N_10557,N_9168);
xor U13666 (N_13666,N_11043,N_10739);
nand U13667 (N_13667,N_11301,N_11059);
nand U13668 (N_13668,N_10748,N_11839);
nand U13669 (N_13669,N_11291,N_11101);
and U13670 (N_13670,N_11135,N_9736);
nor U13671 (N_13671,N_11739,N_11487);
xor U13672 (N_13672,N_11273,N_9063);
nor U13673 (N_13673,N_11582,N_10564);
xor U13674 (N_13674,N_10648,N_11997);
nand U13675 (N_13675,N_11275,N_10830);
xor U13676 (N_13676,N_9628,N_11671);
nor U13677 (N_13677,N_9944,N_9362);
and U13678 (N_13678,N_11199,N_11227);
nor U13679 (N_13679,N_11224,N_11873);
nand U13680 (N_13680,N_9936,N_11492);
and U13681 (N_13681,N_9317,N_9225);
nand U13682 (N_13682,N_10726,N_10391);
or U13683 (N_13683,N_11088,N_9866);
nand U13684 (N_13684,N_11440,N_10114);
and U13685 (N_13685,N_10660,N_11287);
xor U13686 (N_13686,N_9254,N_10007);
nand U13687 (N_13687,N_9352,N_10784);
or U13688 (N_13688,N_11178,N_10730);
nor U13689 (N_13689,N_10668,N_9951);
and U13690 (N_13690,N_10067,N_9093);
or U13691 (N_13691,N_11679,N_11445);
or U13692 (N_13692,N_9873,N_11590);
nor U13693 (N_13693,N_9865,N_10881);
or U13694 (N_13694,N_9788,N_10218);
nand U13695 (N_13695,N_11392,N_10703);
and U13696 (N_13696,N_10344,N_10957);
xor U13697 (N_13697,N_10898,N_9048);
nor U13698 (N_13698,N_11685,N_9195);
xor U13699 (N_13699,N_9632,N_10614);
or U13700 (N_13700,N_11340,N_10683);
nor U13701 (N_13701,N_9342,N_11836);
nor U13702 (N_13702,N_10471,N_10396);
nand U13703 (N_13703,N_9579,N_10692);
xnor U13704 (N_13704,N_9529,N_11381);
xnor U13705 (N_13705,N_10553,N_9655);
nand U13706 (N_13706,N_9161,N_9570);
and U13707 (N_13707,N_9240,N_10829);
nor U13708 (N_13708,N_9356,N_10505);
nor U13709 (N_13709,N_11494,N_10084);
and U13710 (N_13710,N_11070,N_10503);
nor U13711 (N_13711,N_9022,N_11272);
or U13712 (N_13712,N_11610,N_9668);
nand U13713 (N_13713,N_10276,N_11466);
xnor U13714 (N_13714,N_11849,N_10537);
xnor U13715 (N_13715,N_9183,N_10875);
xnor U13716 (N_13716,N_9776,N_11738);
nand U13717 (N_13717,N_9712,N_9436);
nand U13718 (N_13718,N_9997,N_9016);
nand U13719 (N_13719,N_11673,N_10181);
nand U13720 (N_13720,N_9135,N_11372);
and U13721 (N_13721,N_9642,N_10546);
or U13722 (N_13722,N_9291,N_11258);
nor U13723 (N_13723,N_10743,N_10130);
and U13724 (N_13724,N_10794,N_11360);
nor U13725 (N_13725,N_10999,N_11306);
nor U13726 (N_13726,N_10188,N_11141);
nor U13727 (N_13727,N_9033,N_10314);
xnor U13728 (N_13728,N_10651,N_9681);
nand U13729 (N_13729,N_10024,N_9145);
and U13730 (N_13730,N_9608,N_10141);
xnor U13731 (N_13731,N_11015,N_11787);
nand U13732 (N_13732,N_11058,N_10631);
and U13733 (N_13733,N_11867,N_11548);
nor U13734 (N_13734,N_11153,N_10390);
xor U13735 (N_13735,N_9673,N_10964);
nand U13736 (N_13736,N_11748,N_9379);
nand U13737 (N_13737,N_10772,N_11616);
or U13738 (N_13738,N_11174,N_11050);
nand U13739 (N_13739,N_9866,N_11047);
and U13740 (N_13740,N_10270,N_11791);
xnor U13741 (N_13741,N_9635,N_11315);
or U13742 (N_13742,N_11996,N_11286);
nand U13743 (N_13743,N_11140,N_9816);
xnor U13744 (N_13744,N_10229,N_11713);
xor U13745 (N_13745,N_9779,N_11003);
xor U13746 (N_13746,N_11850,N_11115);
xor U13747 (N_13747,N_10668,N_11359);
nand U13748 (N_13748,N_11850,N_9195);
or U13749 (N_13749,N_9316,N_11822);
or U13750 (N_13750,N_11282,N_11371);
and U13751 (N_13751,N_9866,N_10994);
xnor U13752 (N_13752,N_9580,N_11417);
xor U13753 (N_13753,N_11249,N_10898);
and U13754 (N_13754,N_9298,N_9307);
nor U13755 (N_13755,N_9209,N_10134);
nand U13756 (N_13756,N_9006,N_10750);
and U13757 (N_13757,N_9497,N_11243);
and U13758 (N_13758,N_10987,N_10964);
nor U13759 (N_13759,N_11958,N_9559);
and U13760 (N_13760,N_9863,N_10622);
nand U13761 (N_13761,N_10093,N_10659);
xor U13762 (N_13762,N_11801,N_11208);
and U13763 (N_13763,N_10746,N_9465);
xnor U13764 (N_13764,N_9969,N_9124);
xnor U13765 (N_13765,N_9998,N_11709);
or U13766 (N_13766,N_11192,N_11264);
xnor U13767 (N_13767,N_10559,N_10655);
xor U13768 (N_13768,N_11498,N_10205);
and U13769 (N_13769,N_11524,N_11426);
xnor U13770 (N_13770,N_9634,N_9933);
and U13771 (N_13771,N_10095,N_11025);
xnor U13772 (N_13772,N_10717,N_11117);
nor U13773 (N_13773,N_9331,N_10221);
xor U13774 (N_13774,N_11614,N_10042);
or U13775 (N_13775,N_10751,N_9592);
xnor U13776 (N_13776,N_10672,N_9265);
or U13777 (N_13777,N_10417,N_11547);
xnor U13778 (N_13778,N_11816,N_10948);
or U13779 (N_13779,N_11375,N_9884);
nor U13780 (N_13780,N_11286,N_11603);
nor U13781 (N_13781,N_11818,N_10530);
or U13782 (N_13782,N_11158,N_11782);
xnor U13783 (N_13783,N_11741,N_11233);
and U13784 (N_13784,N_11559,N_9226);
and U13785 (N_13785,N_9082,N_10930);
nor U13786 (N_13786,N_9778,N_9507);
xor U13787 (N_13787,N_9160,N_9545);
or U13788 (N_13788,N_10602,N_11545);
nor U13789 (N_13789,N_9187,N_10115);
nand U13790 (N_13790,N_10281,N_11623);
or U13791 (N_13791,N_9682,N_10096);
and U13792 (N_13792,N_10856,N_10658);
or U13793 (N_13793,N_11127,N_9904);
and U13794 (N_13794,N_9647,N_10477);
and U13795 (N_13795,N_9044,N_9258);
nor U13796 (N_13796,N_11469,N_9688);
or U13797 (N_13797,N_10270,N_11038);
and U13798 (N_13798,N_9884,N_11972);
nor U13799 (N_13799,N_10618,N_11867);
xor U13800 (N_13800,N_9295,N_11009);
or U13801 (N_13801,N_9487,N_11396);
nor U13802 (N_13802,N_9463,N_9622);
nor U13803 (N_13803,N_11172,N_10469);
nor U13804 (N_13804,N_11884,N_9920);
nand U13805 (N_13805,N_10695,N_11882);
nor U13806 (N_13806,N_9762,N_11824);
and U13807 (N_13807,N_10176,N_10673);
and U13808 (N_13808,N_11920,N_10478);
and U13809 (N_13809,N_11362,N_11204);
xnor U13810 (N_13810,N_10682,N_11013);
xnor U13811 (N_13811,N_10663,N_9459);
nand U13812 (N_13812,N_11750,N_9602);
nor U13813 (N_13813,N_11786,N_10310);
nand U13814 (N_13814,N_10719,N_9718);
and U13815 (N_13815,N_10229,N_10252);
or U13816 (N_13816,N_9937,N_10565);
or U13817 (N_13817,N_10359,N_11606);
xor U13818 (N_13818,N_10524,N_11680);
nand U13819 (N_13819,N_10146,N_11521);
nand U13820 (N_13820,N_9323,N_11239);
and U13821 (N_13821,N_10568,N_11475);
nand U13822 (N_13822,N_10958,N_9516);
and U13823 (N_13823,N_10784,N_11164);
or U13824 (N_13824,N_9031,N_11205);
or U13825 (N_13825,N_11130,N_10233);
nor U13826 (N_13826,N_9666,N_11258);
and U13827 (N_13827,N_9445,N_9274);
xnor U13828 (N_13828,N_9782,N_9229);
or U13829 (N_13829,N_11651,N_10443);
nor U13830 (N_13830,N_11369,N_10969);
xor U13831 (N_13831,N_11832,N_9108);
nor U13832 (N_13832,N_10153,N_10110);
and U13833 (N_13833,N_10100,N_9533);
nand U13834 (N_13834,N_11644,N_10898);
nand U13835 (N_13835,N_9174,N_9889);
xor U13836 (N_13836,N_10147,N_9310);
or U13837 (N_13837,N_11506,N_10306);
xor U13838 (N_13838,N_10300,N_10442);
xor U13839 (N_13839,N_9431,N_10978);
and U13840 (N_13840,N_10179,N_11894);
nor U13841 (N_13841,N_10627,N_9117);
or U13842 (N_13842,N_9933,N_11221);
and U13843 (N_13843,N_9667,N_10703);
nor U13844 (N_13844,N_10226,N_10237);
nor U13845 (N_13845,N_9010,N_9935);
xor U13846 (N_13846,N_11623,N_9743);
xor U13847 (N_13847,N_11942,N_11125);
and U13848 (N_13848,N_11913,N_9820);
or U13849 (N_13849,N_11960,N_9396);
xnor U13850 (N_13850,N_9380,N_11991);
nand U13851 (N_13851,N_10293,N_9942);
or U13852 (N_13852,N_9716,N_10161);
nand U13853 (N_13853,N_10224,N_10552);
nor U13854 (N_13854,N_9524,N_10537);
nand U13855 (N_13855,N_11374,N_10973);
nor U13856 (N_13856,N_11830,N_9330);
xor U13857 (N_13857,N_10825,N_11377);
or U13858 (N_13858,N_10634,N_11166);
nor U13859 (N_13859,N_10707,N_11854);
and U13860 (N_13860,N_10094,N_11268);
nor U13861 (N_13861,N_9592,N_10922);
nand U13862 (N_13862,N_10295,N_11876);
xor U13863 (N_13863,N_11938,N_9343);
nor U13864 (N_13864,N_11193,N_9078);
nor U13865 (N_13865,N_11627,N_9001);
xnor U13866 (N_13866,N_10743,N_10452);
or U13867 (N_13867,N_10845,N_9589);
nor U13868 (N_13868,N_9122,N_10846);
and U13869 (N_13869,N_11723,N_10707);
xor U13870 (N_13870,N_11497,N_11354);
and U13871 (N_13871,N_9852,N_9764);
and U13872 (N_13872,N_10635,N_11134);
nor U13873 (N_13873,N_11629,N_9959);
nand U13874 (N_13874,N_11788,N_10001);
and U13875 (N_13875,N_10810,N_10914);
nand U13876 (N_13876,N_10370,N_10681);
xor U13877 (N_13877,N_10556,N_10870);
xor U13878 (N_13878,N_11957,N_9626);
or U13879 (N_13879,N_9676,N_11232);
and U13880 (N_13880,N_9089,N_10274);
nand U13881 (N_13881,N_10099,N_10365);
xor U13882 (N_13882,N_11805,N_11430);
and U13883 (N_13883,N_9827,N_11497);
nor U13884 (N_13884,N_10674,N_11750);
nand U13885 (N_13885,N_9741,N_10342);
and U13886 (N_13886,N_11475,N_10779);
and U13887 (N_13887,N_11526,N_10056);
and U13888 (N_13888,N_10960,N_10025);
or U13889 (N_13889,N_9520,N_9820);
nand U13890 (N_13890,N_9876,N_11312);
and U13891 (N_13891,N_9189,N_9203);
xnor U13892 (N_13892,N_11330,N_9207);
nor U13893 (N_13893,N_10675,N_10091);
xor U13894 (N_13894,N_11892,N_11026);
nor U13895 (N_13895,N_10981,N_11293);
or U13896 (N_13896,N_9205,N_11111);
nor U13897 (N_13897,N_11055,N_10340);
or U13898 (N_13898,N_10819,N_11851);
nor U13899 (N_13899,N_10061,N_10663);
nand U13900 (N_13900,N_10449,N_9797);
xor U13901 (N_13901,N_11942,N_11352);
and U13902 (N_13902,N_11384,N_10175);
nand U13903 (N_13903,N_11926,N_10518);
nor U13904 (N_13904,N_9447,N_10796);
xnor U13905 (N_13905,N_10519,N_9218);
and U13906 (N_13906,N_9604,N_9939);
xnor U13907 (N_13907,N_11455,N_11175);
xnor U13908 (N_13908,N_11511,N_11635);
nor U13909 (N_13909,N_9742,N_11336);
or U13910 (N_13910,N_11163,N_11125);
nand U13911 (N_13911,N_10935,N_11706);
xnor U13912 (N_13912,N_10654,N_10091);
xor U13913 (N_13913,N_10164,N_9732);
and U13914 (N_13914,N_10727,N_11802);
xnor U13915 (N_13915,N_11379,N_10576);
nand U13916 (N_13916,N_9686,N_10625);
or U13917 (N_13917,N_11448,N_11001);
xor U13918 (N_13918,N_9421,N_10696);
xnor U13919 (N_13919,N_9547,N_9414);
and U13920 (N_13920,N_9323,N_10889);
xnor U13921 (N_13921,N_9371,N_9856);
nor U13922 (N_13922,N_10041,N_10956);
nor U13923 (N_13923,N_11673,N_9114);
or U13924 (N_13924,N_10805,N_9803);
and U13925 (N_13925,N_11964,N_9145);
or U13926 (N_13926,N_10100,N_10163);
nor U13927 (N_13927,N_9622,N_9451);
xor U13928 (N_13928,N_9074,N_10164);
or U13929 (N_13929,N_9286,N_9942);
and U13930 (N_13930,N_10079,N_10967);
xnor U13931 (N_13931,N_9331,N_10392);
xor U13932 (N_13932,N_10636,N_10667);
xor U13933 (N_13933,N_9895,N_10007);
nand U13934 (N_13934,N_9176,N_10768);
xor U13935 (N_13935,N_10239,N_9978);
and U13936 (N_13936,N_10206,N_11328);
xnor U13937 (N_13937,N_9228,N_9279);
nand U13938 (N_13938,N_11181,N_9252);
or U13939 (N_13939,N_9134,N_11123);
xnor U13940 (N_13940,N_9154,N_11608);
xor U13941 (N_13941,N_10719,N_11741);
or U13942 (N_13942,N_11596,N_9695);
nor U13943 (N_13943,N_11979,N_9918);
and U13944 (N_13944,N_10026,N_9403);
nor U13945 (N_13945,N_9179,N_10410);
and U13946 (N_13946,N_11687,N_10209);
nand U13947 (N_13947,N_9307,N_9812);
nand U13948 (N_13948,N_10329,N_9328);
nor U13949 (N_13949,N_9691,N_11442);
xnor U13950 (N_13950,N_11874,N_9464);
or U13951 (N_13951,N_11929,N_11939);
or U13952 (N_13952,N_11332,N_11139);
or U13953 (N_13953,N_11357,N_9444);
xnor U13954 (N_13954,N_10092,N_11181);
or U13955 (N_13955,N_10737,N_9522);
nand U13956 (N_13956,N_9029,N_11198);
nand U13957 (N_13957,N_10108,N_9854);
and U13958 (N_13958,N_11669,N_9463);
or U13959 (N_13959,N_9697,N_10193);
nand U13960 (N_13960,N_11072,N_10943);
and U13961 (N_13961,N_9586,N_10077);
xor U13962 (N_13962,N_10218,N_10571);
and U13963 (N_13963,N_11627,N_11321);
nor U13964 (N_13964,N_10435,N_10030);
nand U13965 (N_13965,N_9122,N_10207);
and U13966 (N_13966,N_11470,N_10106);
or U13967 (N_13967,N_11831,N_9972);
nand U13968 (N_13968,N_11671,N_9546);
nand U13969 (N_13969,N_10712,N_10321);
nor U13970 (N_13970,N_9036,N_11928);
xnor U13971 (N_13971,N_9191,N_9238);
nor U13972 (N_13972,N_9174,N_11346);
nand U13973 (N_13973,N_9730,N_11345);
nor U13974 (N_13974,N_11034,N_9724);
nand U13975 (N_13975,N_11579,N_10527);
nor U13976 (N_13976,N_11043,N_10400);
xnor U13977 (N_13977,N_10242,N_11407);
xor U13978 (N_13978,N_10217,N_11996);
xnor U13979 (N_13979,N_10928,N_9047);
and U13980 (N_13980,N_11250,N_10213);
nor U13981 (N_13981,N_10943,N_10567);
nand U13982 (N_13982,N_9749,N_9518);
and U13983 (N_13983,N_9708,N_11437);
nor U13984 (N_13984,N_10011,N_9514);
or U13985 (N_13985,N_10086,N_9705);
and U13986 (N_13986,N_9763,N_10187);
nor U13987 (N_13987,N_10656,N_9194);
nand U13988 (N_13988,N_9920,N_11531);
nor U13989 (N_13989,N_9271,N_10050);
nand U13990 (N_13990,N_10033,N_10811);
xor U13991 (N_13991,N_9367,N_9713);
and U13992 (N_13992,N_10534,N_10162);
or U13993 (N_13993,N_10673,N_10004);
and U13994 (N_13994,N_9868,N_11596);
or U13995 (N_13995,N_11581,N_9825);
and U13996 (N_13996,N_10619,N_10218);
or U13997 (N_13997,N_9809,N_9993);
or U13998 (N_13998,N_9161,N_11776);
nand U13999 (N_13999,N_10472,N_9247);
and U14000 (N_14000,N_10099,N_10169);
xnor U14001 (N_14001,N_11280,N_9262);
nor U14002 (N_14002,N_10522,N_11483);
and U14003 (N_14003,N_10647,N_11747);
xor U14004 (N_14004,N_10514,N_11022);
or U14005 (N_14005,N_10350,N_9139);
xnor U14006 (N_14006,N_9280,N_10516);
and U14007 (N_14007,N_9110,N_10685);
nor U14008 (N_14008,N_11404,N_11345);
xor U14009 (N_14009,N_11731,N_11565);
or U14010 (N_14010,N_11290,N_10078);
nor U14011 (N_14011,N_11968,N_10197);
nor U14012 (N_14012,N_10134,N_10877);
or U14013 (N_14013,N_9235,N_11804);
nand U14014 (N_14014,N_9923,N_10401);
and U14015 (N_14015,N_10254,N_9587);
and U14016 (N_14016,N_10107,N_11218);
nand U14017 (N_14017,N_10559,N_9391);
nand U14018 (N_14018,N_9944,N_9366);
xor U14019 (N_14019,N_10361,N_9690);
or U14020 (N_14020,N_10991,N_11606);
nor U14021 (N_14021,N_9245,N_9298);
nor U14022 (N_14022,N_10441,N_9157);
nand U14023 (N_14023,N_10179,N_10882);
nor U14024 (N_14024,N_9222,N_10923);
or U14025 (N_14025,N_10141,N_11655);
or U14026 (N_14026,N_11260,N_11091);
nor U14027 (N_14027,N_9152,N_11009);
and U14028 (N_14028,N_9587,N_9619);
and U14029 (N_14029,N_10036,N_11703);
and U14030 (N_14030,N_11413,N_11987);
xor U14031 (N_14031,N_9847,N_11472);
nor U14032 (N_14032,N_10653,N_10799);
xor U14033 (N_14033,N_9225,N_9382);
or U14034 (N_14034,N_9008,N_9207);
and U14035 (N_14035,N_10446,N_9390);
nor U14036 (N_14036,N_10396,N_9287);
and U14037 (N_14037,N_9725,N_11409);
nand U14038 (N_14038,N_11573,N_10703);
nand U14039 (N_14039,N_9829,N_9246);
xor U14040 (N_14040,N_10153,N_9752);
xnor U14041 (N_14041,N_11685,N_11893);
xor U14042 (N_14042,N_9996,N_9655);
or U14043 (N_14043,N_11753,N_11559);
xnor U14044 (N_14044,N_11581,N_10936);
or U14045 (N_14045,N_9487,N_11632);
nor U14046 (N_14046,N_10096,N_10892);
nor U14047 (N_14047,N_10318,N_9450);
and U14048 (N_14048,N_9222,N_10587);
and U14049 (N_14049,N_9707,N_10262);
xor U14050 (N_14050,N_10575,N_10174);
nand U14051 (N_14051,N_11221,N_10194);
or U14052 (N_14052,N_9440,N_11466);
nand U14053 (N_14053,N_10293,N_9389);
nor U14054 (N_14054,N_9208,N_11771);
nor U14055 (N_14055,N_11041,N_9078);
nand U14056 (N_14056,N_9102,N_9661);
and U14057 (N_14057,N_9242,N_9218);
or U14058 (N_14058,N_9388,N_10175);
or U14059 (N_14059,N_9603,N_9690);
nand U14060 (N_14060,N_11270,N_9245);
nor U14061 (N_14061,N_10854,N_10660);
nand U14062 (N_14062,N_10101,N_11621);
nand U14063 (N_14063,N_10272,N_9575);
and U14064 (N_14064,N_10127,N_11002);
or U14065 (N_14065,N_10243,N_9102);
and U14066 (N_14066,N_11918,N_9496);
nor U14067 (N_14067,N_10595,N_10444);
nor U14068 (N_14068,N_11023,N_11479);
nor U14069 (N_14069,N_10860,N_10644);
nor U14070 (N_14070,N_9610,N_10137);
xnor U14071 (N_14071,N_9372,N_9192);
and U14072 (N_14072,N_10904,N_9141);
xor U14073 (N_14073,N_11508,N_9922);
nor U14074 (N_14074,N_11204,N_11215);
xnor U14075 (N_14075,N_9026,N_9337);
nand U14076 (N_14076,N_10373,N_10581);
or U14077 (N_14077,N_9113,N_10658);
and U14078 (N_14078,N_11279,N_9043);
nand U14079 (N_14079,N_11333,N_11911);
and U14080 (N_14080,N_11512,N_11003);
nor U14081 (N_14081,N_10910,N_10454);
and U14082 (N_14082,N_10667,N_11484);
nor U14083 (N_14083,N_11140,N_11053);
nand U14084 (N_14084,N_11520,N_11844);
nand U14085 (N_14085,N_10231,N_10603);
nand U14086 (N_14086,N_10120,N_9018);
and U14087 (N_14087,N_9747,N_10256);
nand U14088 (N_14088,N_9542,N_9831);
nor U14089 (N_14089,N_9267,N_11477);
or U14090 (N_14090,N_10379,N_9694);
or U14091 (N_14091,N_9499,N_11691);
and U14092 (N_14092,N_11953,N_10332);
and U14093 (N_14093,N_11205,N_10900);
nand U14094 (N_14094,N_9146,N_10706);
nand U14095 (N_14095,N_10501,N_11085);
and U14096 (N_14096,N_9979,N_11904);
nand U14097 (N_14097,N_9110,N_11585);
and U14098 (N_14098,N_9890,N_11652);
xnor U14099 (N_14099,N_9855,N_10217);
or U14100 (N_14100,N_11843,N_10307);
xnor U14101 (N_14101,N_11042,N_9744);
nor U14102 (N_14102,N_10809,N_11229);
or U14103 (N_14103,N_9844,N_11406);
xnor U14104 (N_14104,N_9736,N_9723);
and U14105 (N_14105,N_11890,N_11038);
or U14106 (N_14106,N_11653,N_10855);
and U14107 (N_14107,N_11973,N_11407);
and U14108 (N_14108,N_9380,N_11436);
and U14109 (N_14109,N_9205,N_9786);
nand U14110 (N_14110,N_9202,N_11485);
or U14111 (N_14111,N_9764,N_11240);
or U14112 (N_14112,N_11830,N_9104);
or U14113 (N_14113,N_10586,N_9897);
or U14114 (N_14114,N_11403,N_9928);
nand U14115 (N_14115,N_11251,N_9145);
or U14116 (N_14116,N_9608,N_11961);
nor U14117 (N_14117,N_11610,N_10859);
nor U14118 (N_14118,N_10363,N_10493);
and U14119 (N_14119,N_10496,N_9105);
nor U14120 (N_14120,N_10658,N_10632);
or U14121 (N_14121,N_11138,N_11770);
or U14122 (N_14122,N_9563,N_10708);
or U14123 (N_14123,N_10934,N_9289);
xor U14124 (N_14124,N_9122,N_11038);
nand U14125 (N_14125,N_11921,N_10733);
nand U14126 (N_14126,N_11984,N_11108);
and U14127 (N_14127,N_11526,N_11621);
or U14128 (N_14128,N_11673,N_11899);
and U14129 (N_14129,N_11891,N_11629);
and U14130 (N_14130,N_11245,N_11444);
or U14131 (N_14131,N_9574,N_10519);
xor U14132 (N_14132,N_11898,N_9068);
nor U14133 (N_14133,N_9660,N_9327);
xor U14134 (N_14134,N_11669,N_11048);
or U14135 (N_14135,N_10925,N_10122);
and U14136 (N_14136,N_10885,N_9378);
and U14137 (N_14137,N_10671,N_9982);
xor U14138 (N_14138,N_11088,N_9394);
and U14139 (N_14139,N_9023,N_10075);
nand U14140 (N_14140,N_11001,N_10346);
xor U14141 (N_14141,N_9546,N_9731);
or U14142 (N_14142,N_10949,N_11970);
and U14143 (N_14143,N_11794,N_11711);
xnor U14144 (N_14144,N_10813,N_9135);
nand U14145 (N_14145,N_11592,N_11693);
xnor U14146 (N_14146,N_9574,N_11678);
nand U14147 (N_14147,N_10538,N_10123);
xor U14148 (N_14148,N_9241,N_10116);
nand U14149 (N_14149,N_10524,N_11476);
nand U14150 (N_14150,N_11834,N_11447);
xnor U14151 (N_14151,N_10292,N_11492);
nand U14152 (N_14152,N_11110,N_10421);
nor U14153 (N_14153,N_10542,N_11255);
xor U14154 (N_14154,N_9629,N_9236);
or U14155 (N_14155,N_9571,N_11727);
or U14156 (N_14156,N_11577,N_10439);
and U14157 (N_14157,N_11873,N_10039);
xor U14158 (N_14158,N_10563,N_11440);
and U14159 (N_14159,N_10850,N_9739);
or U14160 (N_14160,N_10640,N_11175);
and U14161 (N_14161,N_11062,N_10863);
or U14162 (N_14162,N_9553,N_9925);
nor U14163 (N_14163,N_11895,N_9912);
nor U14164 (N_14164,N_10722,N_9952);
nand U14165 (N_14165,N_10891,N_11207);
or U14166 (N_14166,N_11833,N_9811);
or U14167 (N_14167,N_10923,N_9449);
nor U14168 (N_14168,N_11242,N_11324);
nand U14169 (N_14169,N_9406,N_9667);
nand U14170 (N_14170,N_11803,N_11808);
or U14171 (N_14171,N_9628,N_10415);
xnor U14172 (N_14172,N_11216,N_9853);
or U14173 (N_14173,N_9476,N_9999);
nand U14174 (N_14174,N_10029,N_10644);
or U14175 (N_14175,N_9855,N_10658);
or U14176 (N_14176,N_11868,N_10634);
nor U14177 (N_14177,N_11008,N_11800);
and U14178 (N_14178,N_9158,N_10553);
nand U14179 (N_14179,N_11717,N_11187);
or U14180 (N_14180,N_10190,N_9807);
or U14181 (N_14181,N_11272,N_9447);
and U14182 (N_14182,N_9021,N_11878);
nor U14183 (N_14183,N_11774,N_11816);
xor U14184 (N_14184,N_9621,N_9651);
or U14185 (N_14185,N_11197,N_9222);
nor U14186 (N_14186,N_9016,N_9173);
nand U14187 (N_14187,N_10104,N_11425);
and U14188 (N_14188,N_11963,N_9001);
or U14189 (N_14189,N_9613,N_11943);
nand U14190 (N_14190,N_10273,N_10081);
and U14191 (N_14191,N_11114,N_10666);
nand U14192 (N_14192,N_11353,N_11521);
nand U14193 (N_14193,N_11660,N_11590);
or U14194 (N_14194,N_9156,N_11523);
xnor U14195 (N_14195,N_9994,N_11748);
nor U14196 (N_14196,N_10185,N_9037);
and U14197 (N_14197,N_11049,N_10120);
nand U14198 (N_14198,N_11315,N_10960);
and U14199 (N_14199,N_9311,N_9154);
nand U14200 (N_14200,N_11105,N_10970);
nand U14201 (N_14201,N_9131,N_9059);
nand U14202 (N_14202,N_10271,N_10916);
nand U14203 (N_14203,N_11539,N_10944);
or U14204 (N_14204,N_9068,N_11331);
and U14205 (N_14205,N_10585,N_10104);
nand U14206 (N_14206,N_11273,N_11291);
nor U14207 (N_14207,N_11065,N_10417);
and U14208 (N_14208,N_10396,N_10764);
nor U14209 (N_14209,N_9994,N_9849);
xnor U14210 (N_14210,N_11803,N_10092);
nor U14211 (N_14211,N_11637,N_10360);
and U14212 (N_14212,N_11218,N_9529);
nand U14213 (N_14213,N_10003,N_10114);
and U14214 (N_14214,N_9362,N_9033);
and U14215 (N_14215,N_11599,N_11798);
nand U14216 (N_14216,N_10728,N_10376);
nor U14217 (N_14217,N_10519,N_11224);
and U14218 (N_14218,N_10677,N_9749);
and U14219 (N_14219,N_10938,N_9097);
or U14220 (N_14220,N_9753,N_9961);
nor U14221 (N_14221,N_11257,N_9376);
or U14222 (N_14222,N_11466,N_9094);
xor U14223 (N_14223,N_10310,N_11644);
and U14224 (N_14224,N_10267,N_10260);
xor U14225 (N_14225,N_11257,N_10845);
nand U14226 (N_14226,N_9857,N_9102);
nor U14227 (N_14227,N_9357,N_9295);
nor U14228 (N_14228,N_10744,N_10878);
nand U14229 (N_14229,N_9647,N_9681);
nand U14230 (N_14230,N_9835,N_11303);
or U14231 (N_14231,N_10913,N_11523);
xnor U14232 (N_14232,N_11314,N_9139);
or U14233 (N_14233,N_9156,N_11687);
or U14234 (N_14234,N_10448,N_9289);
and U14235 (N_14235,N_11565,N_11309);
and U14236 (N_14236,N_9388,N_10821);
nor U14237 (N_14237,N_11539,N_11313);
nor U14238 (N_14238,N_10241,N_9553);
nor U14239 (N_14239,N_10613,N_11377);
nand U14240 (N_14240,N_11877,N_9505);
and U14241 (N_14241,N_9499,N_11010);
nand U14242 (N_14242,N_11844,N_9168);
or U14243 (N_14243,N_9566,N_9193);
nand U14244 (N_14244,N_9046,N_9330);
nand U14245 (N_14245,N_9047,N_10640);
xnor U14246 (N_14246,N_10835,N_11224);
nor U14247 (N_14247,N_11144,N_10076);
and U14248 (N_14248,N_11741,N_11518);
xnor U14249 (N_14249,N_10094,N_9192);
or U14250 (N_14250,N_9382,N_10145);
nor U14251 (N_14251,N_10545,N_9028);
and U14252 (N_14252,N_9373,N_10147);
and U14253 (N_14253,N_11296,N_10513);
nand U14254 (N_14254,N_10860,N_9063);
nor U14255 (N_14255,N_11843,N_11593);
nor U14256 (N_14256,N_11548,N_10468);
and U14257 (N_14257,N_11449,N_11078);
or U14258 (N_14258,N_9827,N_10269);
xor U14259 (N_14259,N_11833,N_9707);
and U14260 (N_14260,N_10876,N_10818);
nor U14261 (N_14261,N_10663,N_10969);
nand U14262 (N_14262,N_10005,N_9707);
xnor U14263 (N_14263,N_9420,N_9141);
xor U14264 (N_14264,N_10848,N_9473);
or U14265 (N_14265,N_9803,N_9559);
xor U14266 (N_14266,N_9116,N_9416);
nand U14267 (N_14267,N_10828,N_10335);
xnor U14268 (N_14268,N_10141,N_10967);
nor U14269 (N_14269,N_9273,N_9366);
or U14270 (N_14270,N_11700,N_11031);
nand U14271 (N_14271,N_10216,N_11223);
or U14272 (N_14272,N_11129,N_11388);
nor U14273 (N_14273,N_11537,N_10257);
nor U14274 (N_14274,N_10233,N_11591);
nor U14275 (N_14275,N_10418,N_11500);
or U14276 (N_14276,N_9465,N_9979);
nor U14277 (N_14277,N_11637,N_10291);
nand U14278 (N_14278,N_10783,N_10193);
nor U14279 (N_14279,N_11466,N_11558);
or U14280 (N_14280,N_11647,N_11227);
and U14281 (N_14281,N_10643,N_10106);
nor U14282 (N_14282,N_11514,N_9639);
nand U14283 (N_14283,N_9147,N_9971);
or U14284 (N_14284,N_11144,N_10760);
and U14285 (N_14285,N_11993,N_9455);
and U14286 (N_14286,N_10423,N_9932);
and U14287 (N_14287,N_10665,N_11875);
or U14288 (N_14288,N_9634,N_9513);
or U14289 (N_14289,N_10287,N_11645);
nor U14290 (N_14290,N_9693,N_11477);
and U14291 (N_14291,N_11346,N_11189);
or U14292 (N_14292,N_10505,N_9414);
xor U14293 (N_14293,N_10913,N_10330);
or U14294 (N_14294,N_9209,N_9093);
nand U14295 (N_14295,N_11069,N_9638);
nand U14296 (N_14296,N_10158,N_10898);
xor U14297 (N_14297,N_9426,N_9612);
nand U14298 (N_14298,N_11716,N_9559);
nand U14299 (N_14299,N_11360,N_10160);
xnor U14300 (N_14300,N_10021,N_11013);
nor U14301 (N_14301,N_11509,N_11627);
nand U14302 (N_14302,N_10556,N_10135);
and U14303 (N_14303,N_9468,N_9917);
nand U14304 (N_14304,N_10289,N_11139);
nand U14305 (N_14305,N_11253,N_11678);
and U14306 (N_14306,N_11271,N_11842);
nand U14307 (N_14307,N_9837,N_10929);
and U14308 (N_14308,N_11934,N_9895);
or U14309 (N_14309,N_10084,N_11492);
nor U14310 (N_14310,N_10386,N_10943);
and U14311 (N_14311,N_10815,N_10026);
nand U14312 (N_14312,N_9468,N_10383);
nand U14313 (N_14313,N_11756,N_9894);
nand U14314 (N_14314,N_11581,N_9465);
nand U14315 (N_14315,N_9052,N_10565);
xor U14316 (N_14316,N_9890,N_11321);
xnor U14317 (N_14317,N_10599,N_11960);
nand U14318 (N_14318,N_11572,N_9456);
nand U14319 (N_14319,N_11922,N_10599);
nand U14320 (N_14320,N_9927,N_11839);
nand U14321 (N_14321,N_10971,N_9734);
or U14322 (N_14322,N_10030,N_10369);
nand U14323 (N_14323,N_10328,N_11804);
or U14324 (N_14324,N_9950,N_11410);
or U14325 (N_14325,N_9134,N_10260);
or U14326 (N_14326,N_9189,N_9226);
nand U14327 (N_14327,N_11049,N_9428);
nor U14328 (N_14328,N_9105,N_9472);
or U14329 (N_14329,N_11969,N_10347);
xnor U14330 (N_14330,N_9820,N_11227);
nand U14331 (N_14331,N_11890,N_10588);
and U14332 (N_14332,N_9638,N_10084);
nand U14333 (N_14333,N_9375,N_11441);
nand U14334 (N_14334,N_11996,N_10078);
and U14335 (N_14335,N_9056,N_10813);
and U14336 (N_14336,N_9692,N_10097);
and U14337 (N_14337,N_9322,N_10904);
xnor U14338 (N_14338,N_9165,N_11714);
nor U14339 (N_14339,N_10633,N_9469);
and U14340 (N_14340,N_11524,N_10970);
xnor U14341 (N_14341,N_9039,N_9424);
nor U14342 (N_14342,N_10287,N_11508);
nand U14343 (N_14343,N_9933,N_10923);
nand U14344 (N_14344,N_9828,N_10682);
and U14345 (N_14345,N_11040,N_10518);
and U14346 (N_14346,N_9793,N_9245);
nor U14347 (N_14347,N_10864,N_10593);
nand U14348 (N_14348,N_11274,N_10498);
and U14349 (N_14349,N_9836,N_11804);
or U14350 (N_14350,N_11232,N_10138);
nand U14351 (N_14351,N_9365,N_9389);
and U14352 (N_14352,N_9000,N_9520);
and U14353 (N_14353,N_9733,N_10996);
and U14354 (N_14354,N_11497,N_11536);
nand U14355 (N_14355,N_11029,N_9650);
or U14356 (N_14356,N_9288,N_11232);
nand U14357 (N_14357,N_9719,N_11434);
and U14358 (N_14358,N_11017,N_10271);
xor U14359 (N_14359,N_9414,N_10741);
nor U14360 (N_14360,N_11887,N_9487);
xnor U14361 (N_14361,N_11049,N_11806);
or U14362 (N_14362,N_11754,N_10940);
or U14363 (N_14363,N_9919,N_11177);
nand U14364 (N_14364,N_11482,N_11371);
xnor U14365 (N_14365,N_10296,N_9006);
nor U14366 (N_14366,N_10634,N_10732);
nor U14367 (N_14367,N_9844,N_9158);
nand U14368 (N_14368,N_11950,N_10634);
xnor U14369 (N_14369,N_9854,N_9639);
nor U14370 (N_14370,N_11503,N_9886);
nor U14371 (N_14371,N_10786,N_10938);
xor U14372 (N_14372,N_11409,N_10963);
and U14373 (N_14373,N_10151,N_10550);
nor U14374 (N_14374,N_11917,N_10113);
nand U14375 (N_14375,N_11175,N_10540);
and U14376 (N_14376,N_11082,N_9487);
nor U14377 (N_14377,N_10828,N_11566);
nor U14378 (N_14378,N_9968,N_11780);
and U14379 (N_14379,N_10866,N_11673);
and U14380 (N_14380,N_9479,N_10782);
xnor U14381 (N_14381,N_11099,N_9629);
nor U14382 (N_14382,N_9946,N_9471);
nand U14383 (N_14383,N_10896,N_11742);
and U14384 (N_14384,N_11297,N_10170);
or U14385 (N_14385,N_11020,N_10891);
nand U14386 (N_14386,N_11654,N_10832);
and U14387 (N_14387,N_11869,N_11876);
and U14388 (N_14388,N_11181,N_11291);
or U14389 (N_14389,N_10111,N_9985);
xor U14390 (N_14390,N_9853,N_9533);
nand U14391 (N_14391,N_9654,N_10817);
nor U14392 (N_14392,N_9270,N_10858);
nor U14393 (N_14393,N_9472,N_11291);
nand U14394 (N_14394,N_11313,N_11560);
or U14395 (N_14395,N_9794,N_9007);
or U14396 (N_14396,N_11920,N_9030);
xnor U14397 (N_14397,N_10519,N_10091);
and U14398 (N_14398,N_10602,N_11195);
and U14399 (N_14399,N_10938,N_9859);
nand U14400 (N_14400,N_11875,N_10657);
or U14401 (N_14401,N_11100,N_9816);
and U14402 (N_14402,N_11947,N_10938);
and U14403 (N_14403,N_9846,N_9345);
nand U14404 (N_14404,N_11560,N_10384);
or U14405 (N_14405,N_9517,N_11798);
xor U14406 (N_14406,N_10735,N_10864);
xor U14407 (N_14407,N_10728,N_9356);
or U14408 (N_14408,N_11524,N_10126);
and U14409 (N_14409,N_9977,N_9479);
nor U14410 (N_14410,N_11534,N_9397);
and U14411 (N_14411,N_10394,N_9929);
and U14412 (N_14412,N_10304,N_11235);
xnor U14413 (N_14413,N_11510,N_11293);
xnor U14414 (N_14414,N_9240,N_11528);
or U14415 (N_14415,N_10893,N_9580);
and U14416 (N_14416,N_9921,N_10002);
nand U14417 (N_14417,N_10343,N_11706);
xor U14418 (N_14418,N_11128,N_9443);
nand U14419 (N_14419,N_10003,N_11450);
nor U14420 (N_14420,N_10525,N_9645);
or U14421 (N_14421,N_9776,N_9291);
or U14422 (N_14422,N_10023,N_10273);
and U14423 (N_14423,N_9996,N_11860);
nand U14424 (N_14424,N_9219,N_9580);
nor U14425 (N_14425,N_9069,N_9780);
nand U14426 (N_14426,N_10651,N_9007);
or U14427 (N_14427,N_11770,N_10086);
xnor U14428 (N_14428,N_9886,N_10990);
xnor U14429 (N_14429,N_9781,N_9798);
nand U14430 (N_14430,N_9751,N_11808);
and U14431 (N_14431,N_10232,N_9297);
nor U14432 (N_14432,N_10622,N_10923);
or U14433 (N_14433,N_10813,N_10895);
nor U14434 (N_14434,N_10351,N_10982);
nor U14435 (N_14435,N_11649,N_10944);
nand U14436 (N_14436,N_10815,N_11236);
and U14437 (N_14437,N_10485,N_9207);
and U14438 (N_14438,N_9350,N_9922);
nand U14439 (N_14439,N_10216,N_9234);
or U14440 (N_14440,N_10027,N_11422);
or U14441 (N_14441,N_10045,N_11483);
or U14442 (N_14442,N_11502,N_11558);
and U14443 (N_14443,N_10058,N_10130);
nor U14444 (N_14444,N_10952,N_10019);
and U14445 (N_14445,N_11129,N_10572);
xnor U14446 (N_14446,N_9825,N_11859);
xnor U14447 (N_14447,N_11855,N_10143);
xor U14448 (N_14448,N_10191,N_9043);
xor U14449 (N_14449,N_11738,N_11874);
xor U14450 (N_14450,N_9936,N_9008);
nor U14451 (N_14451,N_9743,N_11345);
nor U14452 (N_14452,N_11065,N_11465);
nor U14453 (N_14453,N_10752,N_9179);
nand U14454 (N_14454,N_11623,N_11349);
or U14455 (N_14455,N_10109,N_10011);
and U14456 (N_14456,N_10535,N_9080);
nor U14457 (N_14457,N_9399,N_11775);
nor U14458 (N_14458,N_10409,N_11099);
or U14459 (N_14459,N_10857,N_9036);
and U14460 (N_14460,N_10203,N_9463);
xnor U14461 (N_14461,N_10665,N_11296);
xor U14462 (N_14462,N_10135,N_10090);
or U14463 (N_14463,N_9889,N_9302);
nand U14464 (N_14464,N_10857,N_10634);
xor U14465 (N_14465,N_10329,N_9401);
nand U14466 (N_14466,N_10348,N_10908);
and U14467 (N_14467,N_9096,N_9997);
nor U14468 (N_14468,N_9004,N_9425);
or U14469 (N_14469,N_9511,N_10597);
and U14470 (N_14470,N_11207,N_11730);
or U14471 (N_14471,N_10811,N_11451);
or U14472 (N_14472,N_9486,N_10941);
nand U14473 (N_14473,N_9866,N_10119);
xnor U14474 (N_14474,N_9394,N_10148);
nand U14475 (N_14475,N_10451,N_10426);
and U14476 (N_14476,N_9486,N_11587);
nand U14477 (N_14477,N_11453,N_11648);
xnor U14478 (N_14478,N_9951,N_11131);
nor U14479 (N_14479,N_11135,N_10757);
nand U14480 (N_14480,N_10305,N_11806);
nor U14481 (N_14481,N_11525,N_11825);
nor U14482 (N_14482,N_9100,N_10178);
nor U14483 (N_14483,N_11889,N_11868);
or U14484 (N_14484,N_9577,N_9542);
nand U14485 (N_14485,N_9922,N_11638);
xor U14486 (N_14486,N_11861,N_11853);
nand U14487 (N_14487,N_9816,N_11738);
and U14488 (N_14488,N_10147,N_9740);
nor U14489 (N_14489,N_10483,N_11679);
and U14490 (N_14490,N_9163,N_9021);
and U14491 (N_14491,N_10694,N_9077);
nor U14492 (N_14492,N_9026,N_10196);
nor U14493 (N_14493,N_9103,N_9014);
and U14494 (N_14494,N_9268,N_9295);
and U14495 (N_14495,N_9564,N_11987);
nor U14496 (N_14496,N_9971,N_9614);
or U14497 (N_14497,N_10324,N_10051);
xnor U14498 (N_14498,N_10401,N_11558);
nand U14499 (N_14499,N_9949,N_9759);
or U14500 (N_14500,N_11693,N_10442);
nor U14501 (N_14501,N_9513,N_11589);
xnor U14502 (N_14502,N_9656,N_10787);
nor U14503 (N_14503,N_11913,N_10438);
or U14504 (N_14504,N_9442,N_11187);
xnor U14505 (N_14505,N_10996,N_9576);
xor U14506 (N_14506,N_11844,N_9784);
and U14507 (N_14507,N_11247,N_11004);
or U14508 (N_14508,N_9151,N_11013);
xor U14509 (N_14509,N_10439,N_10782);
nor U14510 (N_14510,N_9746,N_10876);
xnor U14511 (N_14511,N_9376,N_10789);
and U14512 (N_14512,N_11978,N_9731);
nand U14513 (N_14513,N_9332,N_11644);
and U14514 (N_14514,N_10457,N_9218);
or U14515 (N_14515,N_10100,N_11745);
or U14516 (N_14516,N_10912,N_10097);
nand U14517 (N_14517,N_9895,N_9699);
nand U14518 (N_14518,N_9232,N_9731);
and U14519 (N_14519,N_10427,N_11647);
nand U14520 (N_14520,N_11025,N_9553);
nand U14521 (N_14521,N_11989,N_11966);
or U14522 (N_14522,N_9516,N_11536);
nor U14523 (N_14523,N_11084,N_10508);
xor U14524 (N_14524,N_9845,N_11572);
xnor U14525 (N_14525,N_11803,N_11218);
nand U14526 (N_14526,N_11129,N_9188);
or U14527 (N_14527,N_11409,N_11263);
nand U14528 (N_14528,N_11341,N_9752);
nand U14529 (N_14529,N_9532,N_10468);
nand U14530 (N_14530,N_10761,N_9557);
or U14531 (N_14531,N_11422,N_11338);
or U14532 (N_14532,N_10604,N_9246);
or U14533 (N_14533,N_9877,N_11353);
xnor U14534 (N_14534,N_10598,N_11073);
and U14535 (N_14535,N_10719,N_10569);
or U14536 (N_14536,N_9016,N_9323);
or U14537 (N_14537,N_10047,N_11790);
nand U14538 (N_14538,N_10628,N_9706);
xnor U14539 (N_14539,N_10648,N_11461);
nor U14540 (N_14540,N_11123,N_11399);
and U14541 (N_14541,N_11066,N_9540);
or U14542 (N_14542,N_9301,N_9703);
nand U14543 (N_14543,N_11104,N_9167);
nor U14544 (N_14544,N_9935,N_10649);
xor U14545 (N_14545,N_9866,N_10586);
nand U14546 (N_14546,N_11121,N_10525);
nor U14547 (N_14547,N_11593,N_11006);
nand U14548 (N_14548,N_10086,N_9270);
or U14549 (N_14549,N_10265,N_11150);
nor U14550 (N_14550,N_11286,N_9078);
and U14551 (N_14551,N_9905,N_11692);
and U14552 (N_14552,N_10605,N_9703);
nor U14553 (N_14553,N_10496,N_10515);
nor U14554 (N_14554,N_10611,N_11577);
nand U14555 (N_14555,N_11355,N_10849);
or U14556 (N_14556,N_10952,N_10188);
nand U14557 (N_14557,N_9588,N_11594);
or U14558 (N_14558,N_11012,N_10906);
nand U14559 (N_14559,N_9343,N_9572);
or U14560 (N_14560,N_10412,N_10171);
and U14561 (N_14561,N_10431,N_9725);
and U14562 (N_14562,N_9747,N_11944);
xnor U14563 (N_14563,N_11779,N_10594);
nor U14564 (N_14564,N_9518,N_11520);
nor U14565 (N_14565,N_11420,N_9425);
or U14566 (N_14566,N_9004,N_11924);
xnor U14567 (N_14567,N_9459,N_11317);
and U14568 (N_14568,N_11930,N_10934);
and U14569 (N_14569,N_10934,N_9660);
xor U14570 (N_14570,N_11510,N_11801);
and U14571 (N_14571,N_10626,N_10085);
nand U14572 (N_14572,N_11396,N_10035);
xor U14573 (N_14573,N_10599,N_10190);
or U14574 (N_14574,N_11242,N_11374);
and U14575 (N_14575,N_10796,N_11221);
and U14576 (N_14576,N_9315,N_10158);
or U14577 (N_14577,N_11593,N_11324);
nor U14578 (N_14578,N_11503,N_11200);
nand U14579 (N_14579,N_11324,N_9813);
nand U14580 (N_14580,N_11645,N_10473);
and U14581 (N_14581,N_11902,N_11913);
nand U14582 (N_14582,N_9207,N_9246);
xnor U14583 (N_14583,N_9755,N_11436);
nand U14584 (N_14584,N_11627,N_10675);
nand U14585 (N_14585,N_10514,N_9700);
and U14586 (N_14586,N_9086,N_11419);
and U14587 (N_14587,N_10301,N_11402);
and U14588 (N_14588,N_9751,N_9152);
or U14589 (N_14589,N_9252,N_10155);
and U14590 (N_14590,N_11244,N_10115);
nand U14591 (N_14591,N_10197,N_9468);
and U14592 (N_14592,N_11975,N_9594);
and U14593 (N_14593,N_11915,N_9568);
nand U14594 (N_14594,N_9143,N_11151);
and U14595 (N_14595,N_11925,N_9576);
or U14596 (N_14596,N_9420,N_9736);
xnor U14597 (N_14597,N_11592,N_11957);
xnor U14598 (N_14598,N_10702,N_10845);
nand U14599 (N_14599,N_10503,N_10866);
or U14600 (N_14600,N_9533,N_9903);
nand U14601 (N_14601,N_9705,N_10659);
or U14602 (N_14602,N_9716,N_11363);
xnor U14603 (N_14603,N_10888,N_9332);
nor U14604 (N_14604,N_9307,N_10618);
and U14605 (N_14605,N_9128,N_10943);
xor U14606 (N_14606,N_9148,N_9728);
and U14607 (N_14607,N_10117,N_11852);
nor U14608 (N_14608,N_11806,N_11292);
xor U14609 (N_14609,N_11596,N_11975);
nor U14610 (N_14610,N_11931,N_10482);
nor U14611 (N_14611,N_9852,N_9465);
or U14612 (N_14612,N_10115,N_11976);
nand U14613 (N_14613,N_10001,N_9626);
and U14614 (N_14614,N_11885,N_11888);
xnor U14615 (N_14615,N_9481,N_10780);
and U14616 (N_14616,N_11125,N_10998);
xor U14617 (N_14617,N_10452,N_9818);
and U14618 (N_14618,N_11360,N_9352);
nand U14619 (N_14619,N_11175,N_9140);
nor U14620 (N_14620,N_11514,N_11035);
and U14621 (N_14621,N_10705,N_10816);
and U14622 (N_14622,N_11537,N_10026);
and U14623 (N_14623,N_11661,N_11885);
nor U14624 (N_14624,N_9166,N_10283);
nor U14625 (N_14625,N_11318,N_10939);
or U14626 (N_14626,N_10209,N_10473);
nor U14627 (N_14627,N_10897,N_11340);
xnor U14628 (N_14628,N_10910,N_9711);
xnor U14629 (N_14629,N_11737,N_10449);
nor U14630 (N_14630,N_11112,N_10550);
nand U14631 (N_14631,N_10681,N_11277);
nand U14632 (N_14632,N_9180,N_11209);
nand U14633 (N_14633,N_11661,N_9436);
nor U14634 (N_14634,N_10999,N_10789);
and U14635 (N_14635,N_10808,N_10755);
or U14636 (N_14636,N_11998,N_10127);
and U14637 (N_14637,N_11438,N_9198);
xor U14638 (N_14638,N_10350,N_11136);
or U14639 (N_14639,N_9967,N_11224);
or U14640 (N_14640,N_11209,N_10931);
nor U14641 (N_14641,N_10072,N_10214);
nand U14642 (N_14642,N_9877,N_11502);
nor U14643 (N_14643,N_10094,N_10696);
nor U14644 (N_14644,N_10763,N_11564);
nand U14645 (N_14645,N_11968,N_9529);
nand U14646 (N_14646,N_9209,N_11287);
xnor U14647 (N_14647,N_11611,N_10711);
nand U14648 (N_14648,N_10382,N_10242);
and U14649 (N_14649,N_11849,N_10899);
xnor U14650 (N_14650,N_10338,N_11266);
and U14651 (N_14651,N_11904,N_10936);
nand U14652 (N_14652,N_10552,N_10236);
nor U14653 (N_14653,N_9551,N_11734);
nor U14654 (N_14654,N_11820,N_9315);
and U14655 (N_14655,N_9665,N_10659);
nor U14656 (N_14656,N_9795,N_11749);
and U14657 (N_14657,N_9756,N_10109);
xnor U14658 (N_14658,N_11718,N_11460);
nand U14659 (N_14659,N_10094,N_11581);
nor U14660 (N_14660,N_10387,N_11208);
xnor U14661 (N_14661,N_9542,N_10893);
nor U14662 (N_14662,N_10715,N_9959);
nor U14663 (N_14663,N_9273,N_9483);
xnor U14664 (N_14664,N_11412,N_10107);
or U14665 (N_14665,N_10578,N_9579);
xor U14666 (N_14666,N_9666,N_10149);
and U14667 (N_14667,N_9611,N_9419);
nor U14668 (N_14668,N_10207,N_10062);
and U14669 (N_14669,N_9514,N_11959);
or U14670 (N_14670,N_10994,N_11544);
xor U14671 (N_14671,N_9020,N_10077);
nand U14672 (N_14672,N_10082,N_9239);
xnor U14673 (N_14673,N_11989,N_9155);
or U14674 (N_14674,N_9318,N_11560);
xnor U14675 (N_14675,N_9923,N_11607);
nor U14676 (N_14676,N_10047,N_10346);
nand U14677 (N_14677,N_9247,N_9563);
or U14678 (N_14678,N_11379,N_9501);
nand U14679 (N_14679,N_11947,N_11107);
or U14680 (N_14680,N_9757,N_11315);
nor U14681 (N_14681,N_10566,N_10643);
and U14682 (N_14682,N_10851,N_9815);
nor U14683 (N_14683,N_11026,N_10793);
xnor U14684 (N_14684,N_9101,N_11263);
nand U14685 (N_14685,N_9258,N_9359);
xor U14686 (N_14686,N_10396,N_11291);
or U14687 (N_14687,N_11689,N_9935);
or U14688 (N_14688,N_9919,N_11164);
nand U14689 (N_14689,N_10759,N_11866);
nand U14690 (N_14690,N_9358,N_10305);
xnor U14691 (N_14691,N_9376,N_9545);
and U14692 (N_14692,N_9887,N_10871);
nor U14693 (N_14693,N_10810,N_9829);
xor U14694 (N_14694,N_11040,N_10567);
and U14695 (N_14695,N_10264,N_10850);
nor U14696 (N_14696,N_11551,N_10820);
xnor U14697 (N_14697,N_11886,N_9003);
nand U14698 (N_14698,N_10144,N_10738);
and U14699 (N_14699,N_11656,N_11727);
nand U14700 (N_14700,N_10193,N_11253);
or U14701 (N_14701,N_9963,N_11478);
nand U14702 (N_14702,N_11536,N_11555);
xor U14703 (N_14703,N_10989,N_9295);
nand U14704 (N_14704,N_11833,N_9214);
or U14705 (N_14705,N_11966,N_9645);
or U14706 (N_14706,N_11652,N_10751);
xor U14707 (N_14707,N_11786,N_10089);
nor U14708 (N_14708,N_11314,N_11577);
nor U14709 (N_14709,N_10202,N_9917);
or U14710 (N_14710,N_10289,N_10405);
xnor U14711 (N_14711,N_10486,N_11729);
xor U14712 (N_14712,N_11268,N_9768);
nand U14713 (N_14713,N_11071,N_9121);
nor U14714 (N_14714,N_10186,N_9020);
and U14715 (N_14715,N_10833,N_10725);
xnor U14716 (N_14716,N_10607,N_10976);
xnor U14717 (N_14717,N_10709,N_9957);
or U14718 (N_14718,N_9957,N_9128);
xor U14719 (N_14719,N_10796,N_11010);
and U14720 (N_14720,N_10488,N_10192);
or U14721 (N_14721,N_10351,N_11965);
and U14722 (N_14722,N_11014,N_10530);
xor U14723 (N_14723,N_9281,N_11393);
nand U14724 (N_14724,N_10245,N_10896);
nor U14725 (N_14725,N_11506,N_9832);
and U14726 (N_14726,N_11992,N_9680);
and U14727 (N_14727,N_10501,N_11761);
and U14728 (N_14728,N_10853,N_11875);
nand U14729 (N_14729,N_10262,N_11820);
or U14730 (N_14730,N_10340,N_9956);
and U14731 (N_14731,N_10438,N_10014);
nand U14732 (N_14732,N_10389,N_9133);
nor U14733 (N_14733,N_9313,N_10210);
nor U14734 (N_14734,N_11759,N_9419);
nor U14735 (N_14735,N_10392,N_11961);
and U14736 (N_14736,N_10172,N_11582);
or U14737 (N_14737,N_10160,N_10862);
nor U14738 (N_14738,N_9525,N_11085);
xor U14739 (N_14739,N_9414,N_9677);
nand U14740 (N_14740,N_9447,N_9469);
or U14741 (N_14741,N_11346,N_9919);
nand U14742 (N_14742,N_10498,N_10000);
nand U14743 (N_14743,N_11983,N_10592);
nand U14744 (N_14744,N_9647,N_10852);
xnor U14745 (N_14745,N_10387,N_9211);
or U14746 (N_14746,N_11422,N_10179);
nor U14747 (N_14747,N_10085,N_9181);
and U14748 (N_14748,N_9495,N_9221);
nor U14749 (N_14749,N_9775,N_11857);
and U14750 (N_14750,N_10533,N_10679);
xor U14751 (N_14751,N_10213,N_11241);
xnor U14752 (N_14752,N_10828,N_11919);
and U14753 (N_14753,N_11623,N_9354);
and U14754 (N_14754,N_11629,N_9557);
or U14755 (N_14755,N_9471,N_11711);
xnor U14756 (N_14756,N_10484,N_9303);
nand U14757 (N_14757,N_11439,N_10339);
nand U14758 (N_14758,N_11882,N_10701);
or U14759 (N_14759,N_11934,N_11019);
nor U14760 (N_14760,N_11391,N_9241);
xor U14761 (N_14761,N_10081,N_9659);
nor U14762 (N_14762,N_9470,N_9138);
nor U14763 (N_14763,N_9562,N_11669);
nand U14764 (N_14764,N_10641,N_10744);
or U14765 (N_14765,N_10064,N_10650);
nand U14766 (N_14766,N_11158,N_11319);
nand U14767 (N_14767,N_9894,N_9958);
and U14768 (N_14768,N_11674,N_10059);
nor U14769 (N_14769,N_10954,N_11423);
xnor U14770 (N_14770,N_11363,N_10024);
nor U14771 (N_14771,N_10352,N_10975);
nor U14772 (N_14772,N_9212,N_9618);
nor U14773 (N_14773,N_11329,N_9697);
nand U14774 (N_14774,N_11155,N_10127);
and U14775 (N_14775,N_10004,N_11548);
nor U14776 (N_14776,N_10175,N_9609);
nand U14777 (N_14777,N_9320,N_9180);
nand U14778 (N_14778,N_11342,N_11924);
and U14779 (N_14779,N_10158,N_9981);
nor U14780 (N_14780,N_11215,N_11873);
or U14781 (N_14781,N_9141,N_10884);
nand U14782 (N_14782,N_9372,N_10003);
nand U14783 (N_14783,N_9719,N_11813);
and U14784 (N_14784,N_10089,N_11822);
and U14785 (N_14785,N_9236,N_10619);
nor U14786 (N_14786,N_11558,N_11290);
and U14787 (N_14787,N_10214,N_10480);
or U14788 (N_14788,N_9623,N_9392);
nor U14789 (N_14789,N_10110,N_11874);
or U14790 (N_14790,N_9942,N_9832);
or U14791 (N_14791,N_10647,N_9856);
xor U14792 (N_14792,N_9955,N_10832);
or U14793 (N_14793,N_11872,N_11469);
nand U14794 (N_14794,N_10257,N_10148);
or U14795 (N_14795,N_11980,N_9852);
or U14796 (N_14796,N_10990,N_9254);
xor U14797 (N_14797,N_9532,N_9987);
and U14798 (N_14798,N_10435,N_10975);
nand U14799 (N_14799,N_10804,N_11838);
and U14800 (N_14800,N_9170,N_11137);
xor U14801 (N_14801,N_9944,N_9619);
and U14802 (N_14802,N_11351,N_10720);
and U14803 (N_14803,N_9514,N_11904);
xor U14804 (N_14804,N_9569,N_10464);
nor U14805 (N_14805,N_9115,N_10072);
xnor U14806 (N_14806,N_11318,N_11480);
and U14807 (N_14807,N_10145,N_10922);
nand U14808 (N_14808,N_9955,N_9922);
nand U14809 (N_14809,N_11619,N_11254);
nor U14810 (N_14810,N_11425,N_10893);
and U14811 (N_14811,N_11161,N_10089);
or U14812 (N_14812,N_11429,N_10208);
nand U14813 (N_14813,N_11336,N_10499);
xor U14814 (N_14814,N_11915,N_10318);
nand U14815 (N_14815,N_10821,N_9660);
or U14816 (N_14816,N_9541,N_10480);
and U14817 (N_14817,N_11952,N_10037);
nand U14818 (N_14818,N_10128,N_9382);
and U14819 (N_14819,N_10303,N_9814);
nand U14820 (N_14820,N_11551,N_10529);
nor U14821 (N_14821,N_11014,N_11873);
xor U14822 (N_14822,N_11198,N_9786);
nor U14823 (N_14823,N_10171,N_10184);
xnor U14824 (N_14824,N_9043,N_10509);
and U14825 (N_14825,N_11203,N_9622);
and U14826 (N_14826,N_9182,N_10827);
xor U14827 (N_14827,N_11289,N_9766);
and U14828 (N_14828,N_10309,N_9637);
xor U14829 (N_14829,N_11832,N_11705);
or U14830 (N_14830,N_11731,N_10464);
xor U14831 (N_14831,N_10919,N_11833);
nor U14832 (N_14832,N_11901,N_10935);
and U14833 (N_14833,N_11014,N_11916);
nand U14834 (N_14834,N_11411,N_10339);
and U14835 (N_14835,N_9738,N_11566);
nand U14836 (N_14836,N_11144,N_11486);
nor U14837 (N_14837,N_10869,N_11826);
nor U14838 (N_14838,N_11358,N_10597);
xor U14839 (N_14839,N_9269,N_9209);
and U14840 (N_14840,N_9764,N_11544);
xor U14841 (N_14841,N_11690,N_11153);
and U14842 (N_14842,N_11254,N_9791);
nor U14843 (N_14843,N_9117,N_10015);
nor U14844 (N_14844,N_9519,N_9035);
nand U14845 (N_14845,N_10499,N_10290);
or U14846 (N_14846,N_9261,N_10240);
and U14847 (N_14847,N_11674,N_9422);
nor U14848 (N_14848,N_10336,N_11774);
xnor U14849 (N_14849,N_11054,N_11192);
and U14850 (N_14850,N_10408,N_9270);
xnor U14851 (N_14851,N_9745,N_11706);
and U14852 (N_14852,N_9591,N_11766);
xor U14853 (N_14853,N_11729,N_10061);
nand U14854 (N_14854,N_11215,N_11635);
xnor U14855 (N_14855,N_11212,N_9494);
xor U14856 (N_14856,N_10657,N_9296);
xor U14857 (N_14857,N_9751,N_10918);
or U14858 (N_14858,N_9864,N_11734);
xor U14859 (N_14859,N_11314,N_10758);
nand U14860 (N_14860,N_9190,N_11887);
and U14861 (N_14861,N_10862,N_10694);
and U14862 (N_14862,N_11196,N_9751);
nor U14863 (N_14863,N_11870,N_10728);
xnor U14864 (N_14864,N_9159,N_9599);
nand U14865 (N_14865,N_9696,N_10799);
or U14866 (N_14866,N_10256,N_11035);
nor U14867 (N_14867,N_10393,N_10852);
nor U14868 (N_14868,N_11958,N_9273);
nor U14869 (N_14869,N_9424,N_9692);
nor U14870 (N_14870,N_9045,N_11731);
nand U14871 (N_14871,N_11994,N_11691);
xor U14872 (N_14872,N_9952,N_9444);
and U14873 (N_14873,N_10436,N_9346);
and U14874 (N_14874,N_11279,N_9808);
or U14875 (N_14875,N_11438,N_9405);
nand U14876 (N_14876,N_10277,N_11389);
and U14877 (N_14877,N_11305,N_11065);
xnor U14878 (N_14878,N_9748,N_11219);
and U14879 (N_14879,N_10737,N_9278);
or U14880 (N_14880,N_9829,N_9843);
or U14881 (N_14881,N_11417,N_9309);
nand U14882 (N_14882,N_10867,N_10064);
xnor U14883 (N_14883,N_9164,N_10269);
nor U14884 (N_14884,N_9671,N_9815);
and U14885 (N_14885,N_9146,N_9989);
xnor U14886 (N_14886,N_11792,N_9487);
nor U14887 (N_14887,N_11884,N_9126);
or U14888 (N_14888,N_11317,N_11324);
or U14889 (N_14889,N_11157,N_9225);
nand U14890 (N_14890,N_10109,N_9172);
or U14891 (N_14891,N_9652,N_11063);
xnor U14892 (N_14892,N_11444,N_11908);
xor U14893 (N_14893,N_11376,N_11311);
xor U14894 (N_14894,N_10396,N_9737);
xnor U14895 (N_14895,N_11338,N_10683);
nand U14896 (N_14896,N_11984,N_10915);
nor U14897 (N_14897,N_9461,N_9148);
nor U14898 (N_14898,N_10761,N_10055);
and U14899 (N_14899,N_10352,N_11160);
nand U14900 (N_14900,N_9735,N_11578);
nand U14901 (N_14901,N_9075,N_10824);
nand U14902 (N_14902,N_11446,N_10894);
nand U14903 (N_14903,N_9219,N_9661);
xnor U14904 (N_14904,N_11657,N_9769);
nor U14905 (N_14905,N_11504,N_9679);
or U14906 (N_14906,N_9312,N_11336);
xor U14907 (N_14907,N_11861,N_11433);
or U14908 (N_14908,N_10044,N_9908);
and U14909 (N_14909,N_9519,N_10224);
and U14910 (N_14910,N_10962,N_11150);
xor U14911 (N_14911,N_10104,N_10723);
and U14912 (N_14912,N_11301,N_9281);
xnor U14913 (N_14913,N_11902,N_10604);
xnor U14914 (N_14914,N_9775,N_10254);
xnor U14915 (N_14915,N_11998,N_9074);
xor U14916 (N_14916,N_10300,N_11497);
or U14917 (N_14917,N_10898,N_10169);
or U14918 (N_14918,N_11843,N_11785);
nand U14919 (N_14919,N_10294,N_11343);
nand U14920 (N_14920,N_11359,N_10670);
nor U14921 (N_14921,N_10729,N_9811);
and U14922 (N_14922,N_10149,N_11094);
nor U14923 (N_14923,N_10527,N_9999);
xor U14924 (N_14924,N_9267,N_11322);
and U14925 (N_14925,N_9239,N_11825);
nand U14926 (N_14926,N_9699,N_10505);
nor U14927 (N_14927,N_10368,N_10480);
nand U14928 (N_14928,N_9573,N_9726);
xor U14929 (N_14929,N_11594,N_11388);
and U14930 (N_14930,N_9009,N_11574);
or U14931 (N_14931,N_9941,N_11219);
nand U14932 (N_14932,N_10306,N_9789);
xnor U14933 (N_14933,N_9700,N_11721);
nand U14934 (N_14934,N_11710,N_11403);
and U14935 (N_14935,N_11413,N_11844);
or U14936 (N_14936,N_9534,N_10669);
nor U14937 (N_14937,N_11489,N_10847);
or U14938 (N_14938,N_11715,N_9216);
nor U14939 (N_14939,N_10498,N_11720);
nor U14940 (N_14940,N_10218,N_11412);
or U14941 (N_14941,N_11143,N_11346);
or U14942 (N_14942,N_10397,N_9293);
and U14943 (N_14943,N_11954,N_10268);
and U14944 (N_14944,N_11658,N_10902);
and U14945 (N_14945,N_9871,N_9701);
nor U14946 (N_14946,N_11638,N_9452);
or U14947 (N_14947,N_9347,N_10727);
and U14948 (N_14948,N_11215,N_9445);
nor U14949 (N_14949,N_9916,N_9872);
or U14950 (N_14950,N_10104,N_11397);
xnor U14951 (N_14951,N_9054,N_10722);
nor U14952 (N_14952,N_11917,N_9850);
and U14953 (N_14953,N_9905,N_9423);
or U14954 (N_14954,N_9312,N_11076);
or U14955 (N_14955,N_10897,N_11253);
nor U14956 (N_14956,N_10631,N_9104);
nand U14957 (N_14957,N_10282,N_9425);
xor U14958 (N_14958,N_10013,N_10162);
and U14959 (N_14959,N_11093,N_10123);
nand U14960 (N_14960,N_9413,N_9990);
nand U14961 (N_14961,N_9781,N_9932);
or U14962 (N_14962,N_11875,N_11466);
or U14963 (N_14963,N_11885,N_11656);
or U14964 (N_14964,N_9658,N_10519);
nor U14965 (N_14965,N_11154,N_11384);
xor U14966 (N_14966,N_10357,N_11585);
xnor U14967 (N_14967,N_9396,N_11399);
nor U14968 (N_14968,N_11582,N_11632);
nand U14969 (N_14969,N_10400,N_9096);
nor U14970 (N_14970,N_10923,N_10423);
nor U14971 (N_14971,N_10850,N_9183);
nand U14972 (N_14972,N_11225,N_10933);
xor U14973 (N_14973,N_10835,N_11818);
xnor U14974 (N_14974,N_10520,N_11253);
and U14975 (N_14975,N_11517,N_10886);
or U14976 (N_14976,N_11105,N_11623);
nand U14977 (N_14977,N_9449,N_11955);
nor U14978 (N_14978,N_11357,N_9730);
or U14979 (N_14979,N_11215,N_9208);
nor U14980 (N_14980,N_10685,N_11881);
nor U14981 (N_14981,N_9293,N_11433);
or U14982 (N_14982,N_11629,N_10273);
xor U14983 (N_14983,N_10787,N_9448);
nand U14984 (N_14984,N_10591,N_9125);
xor U14985 (N_14985,N_10730,N_10537);
nor U14986 (N_14986,N_11289,N_9954);
or U14987 (N_14987,N_10896,N_9615);
xnor U14988 (N_14988,N_11086,N_11844);
nand U14989 (N_14989,N_9364,N_11753);
nor U14990 (N_14990,N_10590,N_10675);
xnor U14991 (N_14991,N_9371,N_9857);
xor U14992 (N_14992,N_10060,N_9626);
xor U14993 (N_14993,N_10961,N_9301);
nor U14994 (N_14994,N_9426,N_9384);
xor U14995 (N_14995,N_10468,N_9782);
nand U14996 (N_14996,N_10154,N_11629);
or U14997 (N_14997,N_11061,N_10127);
nor U14998 (N_14998,N_10677,N_9136);
nand U14999 (N_14999,N_9573,N_10462);
nand U15000 (N_15000,N_14771,N_12296);
nand U15001 (N_15001,N_12292,N_12764);
xor U15002 (N_15002,N_14471,N_12055);
and U15003 (N_15003,N_13649,N_14162);
nand U15004 (N_15004,N_13604,N_12576);
nand U15005 (N_15005,N_14353,N_13836);
and U15006 (N_15006,N_14462,N_12769);
nand U15007 (N_15007,N_13833,N_13442);
xor U15008 (N_15008,N_14830,N_12114);
nand U15009 (N_15009,N_12862,N_14036);
and U15010 (N_15010,N_14695,N_12210);
nand U15011 (N_15011,N_13124,N_12207);
nor U15012 (N_15012,N_14596,N_13876);
or U15013 (N_15013,N_12911,N_14292);
xor U15014 (N_15014,N_12627,N_14950);
and U15015 (N_15015,N_14870,N_12496);
xor U15016 (N_15016,N_14285,N_14959);
or U15017 (N_15017,N_13643,N_14061);
or U15018 (N_15018,N_14661,N_14675);
nor U15019 (N_15019,N_12806,N_12886);
or U15020 (N_15020,N_12070,N_14835);
xor U15021 (N_15021,N_12714,N_14760);
or U15022 (N_15022,N_13663,N_12614);
or U15023 (N_15023,N_14704,N_13157);
xor U15024 (N_15024,N_14603,N_12030);
xor U15025 (N_15025,N_13476,N_14310);
and U15026 (N_15026,N_12646,N_14159);
nor U15027 (N_15027,N_13976,N_12303);
nand U15028 (N_15028,N_13421,N_13725);
nand U15029 (N_15029,N_13408,N_13794);
or U15030 (N_15030,N_13808,N_13204);
xnor U15031 (N_15031,N_14026,N_14534);
and U15032 (N_15032,N_14081,N_13728);
nand U15033 (N_15033,N_13016,N_14803);
nor U15034 (N_15034,N_14203,N_12887);
and U15035 (N_15035,N_14982,N_12565);
and U15036 (N_15036,N_13630,N_14670);
nand U15037 (N_15037,N_12486,N_12703);
and U15038 (N_15038,N_14338,N_13650);
or U15039 (N_15039,N_13196,N_14384);
or U15040 (N_15040,N_14883,N_12403);
xnor U15041 (N_15041,N_12766,N_12038);
nor U15042 (N_15042,N_14598,N_14891);
nand U15043 (N_15043,N_14755,N_12608);
nor U15044 (N_15044,N_14696,N_14811);
and U15045 (N_15045,N_13647,N_12276);
nor U15046 (N_15046,N_13482,N_13293);
nand U15047 (N_15047,N_14067,N_13822);
nand U15048 (N_15048,N_13548,N_14770);
xor U15049 (N_15049,N_14634,N_12432);
nor U15050 (N_15050,N_12449,N_13942);
or U15051 (N_15051,N_14132,N_13273);
nand U15052 (N_15052,N_12297,N_13325);
xor U15053 (N_15053,N_14482,N_13475);
xnor U15054 (N_15054,N_12270,N_14594);
or U15055 (N_15055,N_13358,N_12939);
or U15056 (N_15056,N_12651,N_13573);
nor U15057 (N_15057,N_12082,N_14712);
or U15058 (N_15058,N_12568,N_12801);
nor U15059 (N_15059,N_12416,N_13661);
nand U15060 (N_15060,N_12983,N_12340);
xnor U15061 (N_15061,N_13884,N_14046);
xor U15062 (N_15062,N_12294,N_13451);
xor U15063 (N_15063,N_13623,N_12360);
xor U15064 (N_15064,N_13017,N_12421);
xor U15065 (N_15065,N_13207,N_14645);
xnor U15066 (N_15066,N_12420,N_14711);
or U15067 (N_15067,N_12366,N_13802);
or U15068 (N_15068,N_12238,N_14642);
and U15069 (N_15069,N_14457,N_14300);
xnor U15070 (N_15070,N_13436,N_14391);
nand U15071 (N_15071,N_12049,N_12811);
nor U15072 (N_15072,N_13188,N_13312);
or U15073 (N_15073,N_14239,N_12822);
nand U15074 (N_15074,N_14312,N_13973);
xnor U15075 (N_15075,N_13185,N_14946);
nand U15076 (N_15076,N_13299,N_12864);
and U15077 (N_15077,N_14004,N_13128);
and U15078 (N_15078,N_12230,N_12320);
nor U15079 (N_15079,N_14996,N_13422);
and U15080 (N_15080,N_14914,N_14437);
xor U15081 (N_15081,N_13275,N_14703);
or U15082 (N_15082,N_12059,N_13353);
nor U15083 (N_15083,N_12935,N_14054);
nor U15084 (N_15084,N_12922,N_14990);
and U15085 (N_15085,N_12448,N_14541);
nand U15086 (N_15086,N_13637,N_12702);
or U15087 (N_15087,N_14301,N_14268);
and U15088 (N_15088,N_12890,N_12657);
xnor U15089 (N_15089,N_13787,N_13918);
nand U15090 (N_15090,N_12955,N_12741);
xor U15091 (N_15091,N_13211,N_12832);
or U15092 (N_15092,N_13321,N_12918);
or U15093 (N_15093,N_14658,N_14813);
xor U15094 (N_15094,N_13988,N_13804);
or U15095 (N_15095,N_13463,N_13512);
nor U15096 (N_15096,N_14082,N_14442);
nand U15097 (N_15097,N_13372,N_13403);
or U15098 (N_15098,N_13898,N_14084);
nor U15099 (N_15099,N_14524,N_14466);
or U15100 (N_15100,N_14971,N_12845);
xnor U15101 (N_15101,N_14791,N_14907);
nand U15102 (N_15102,N_14753,N_12986);
nor U15103 (N_15103,N_14308,N_13670);
xor U15104 (N_15104,N_14339,N_12966);
nand U15105 (N_15105,N_12690,N_12122);
xor U15106 (N_15106,N_14343,N_14931);
and U15107 (N_15107,N_14359,N_13152);
nand U15108 (N_15108,N_13444,N_14049);
and U15109 (N_15109,N_12633,N_12944);
nand U15110 (N_15110,N_13595,N_14341);
or U15111 (N_15111,N_12869,N_14627);
and U15112 (N_15112,N_13935,N_13539);
and U15113 (N_15113,N_12119,N_14792);
nor U15114 (N_15114,N_14629,N_12020);
nand U15115 (N_15115,N_12200,N_14826);
and U15116 (N_15116,N_13731,N_13316);
nand U15117 (N_15117,N_14477,N_12708);
and U15118 (N_15118,N_12293,N_13845);
xor U15119 (N_15119,N_14796,N_12325);
nand U15120 (N_15120,N_14323,N_13335);
nor U15121 (N_15121,N_12251,N_14702);
xnor U15122 (N_15122,N_13525,N_12662);
or U15123 (N_15123,N_12156,N_14861);
and U15124 (N_15124,N_13025,N_14684);
nand U15125 (N_15125,N_14587,N_14106);
nor U15126 (N_15126,N_13428,N_12816);
and U15127 (N_15127,N_12733,N_12850);
nor U15128 (N_15128,N_13151,N_14983);
or U15129 (N_15129,N_12613,N_12726);
nor U15130 (N_15130,N_14230,N_12826);
and U15131 (N_15131,N_13399,N_14052);
or U15132 (N_15132,N_14839,N_13896);
nand U15133 (N_15133,N_12794,N_12670);
xor U15134 (N_15134,N_12438,N_14757);
nand U15135 (N_15135,N_14352,N_14032);
nor U15136 (N_15136,N_14577,N_13668);
xor U15137 (N_15137,N_14389,N_12335);
and U15138 (N_15138,N_14947,N_13089);
xor U15139 (N_15139,N_12245,N_12218);
or U15140 (N_15140,N_13302,N_13447);
and U15141 (N_15141,N_12900,N_13400);
nor U15142 (N_15142,N_12434,N_12511);
nand U15143 (N_15143,N_14250,N_14936);
nor U15144 (N_15144,N_13813,N_13270);
and U15145 (N_15145,N_13798,N_12593);
or U15146 (N_15146,N_12023,N_14179);
nor U15147 (N_15147,N_13900,N_14655);
nor U15148 (N_15148,N_13734,N_14868);
nor U15149 (N_15149,N_13491,N_12555);
nor U15150 (N_15150,N_14922,N_13772);
nor U15151 (N_15151,N_13298,N_14354);
xnor U15152 (N_15152,N_13111,N_13245);
nand U15153 (N_15153,N_13379,N_14356);
and U15154 (N_15154,N_13799,N_14360);
nand U15155 (N_15155,N_13954,N_13891);
nor U15156 (N_15156,N_14657,N_12202);
nor U15157 (N_15157,N_14433,N_14881);
nor U15158 (N_15158,N_14663,N_12760);
xnor U15159 (N_15159,N_14255,N_13021);
or U15160 (N_15160,N_14664,N_14681);
nor U15161 (N_15161,N_14593,N_12800);
nor U15162 (N_15162,N_13061,N_13176);
nor U15163 (N_15163,N_13425,N_14365);
nand U15164 (N_15164,N_14824,N_12780);
or U15165 (N_15165,N_14428,N_13240);
xor U15166 (N_15166,N_13177,N_14966);
xnor U15167 (N_15167,N_12962,N_14610);
nor U15168 (N_15168,N_14137,N_13378);
nand U15169 (N_15169,N_13878,N_13116);
xor U15170 (N_15170,N_12285,N_13112);
nand U15171 (N_15171,N_13354,N_12765);
or U15172 (N_15172,N_12088,N_12799);
and U15173 (N_15173,N_13989,N_12013);
or U15174 (N_15174,N_13059,N_13076);
or U15175 (N_15175,N_12923,N_13655);
nand U15176 (N_15176,N_13713,N_12880);
and U15177 (N_15177,N_13214,N_12570);
or U15178 (N_15178,N_13841,N_14709);
nor U15179 (N_15179,N_12594,N_14731);
nand U15180 (N_15180,N_13824,N_13559);
xnor U15181 (N_15181,N_14238,N_12635);
nand U15182 (N_15182,N_12424,N_13707);
or U15183 (N_15183,N_13938,N_13764);
nand U15184 (N_15184,N_12569,N_12129);
and U15185 (N_15185,N_13856,N_12740);
nor U15186 (N_15186,N_14463,N_13598);
and U15187 (N_15187,N_13727,N_13518);
and U15188 (N_15188,N_13170,N_13955);
xnor U15189 (N_15189,N_12179,N_13979);
xor U15190 (N_15190,N_14960,N_13102);
xor U15191 (N_15191,N_13513,N_13641);
xnor U15192 (N_15192,N_14993,N_13117);
xor U15193 (N_15193,N_12560,N_13404);
or U15194 (N_15194,N_14799,N_13737);
nand U15195 (N_15195,N_14409,N_13004);
or U15196 (N_15196,N_13178,N_12804);
nand U15197 (N_15197,N_14837,N_12561);
or U15198 (N_15198,N_12056,N_12895);
nand U15199 (N_15199,N_13012,N_13949);
nor U15200 (N_15200,N_13168,N_13415);
xor U15201 (N_15201,N_12399,N_12228);
xor U15202 (N_15202,N_14079,N_12326);
xnor U15203 (N_15203,N_12332,N_14977);
nand U15204 (N_15204,N_14388,N_12357);
xnor U15205 (N_15205,N_12379,N_12289);
xnor U15206 (N_15206,N_13295,N_14019);
and U15207 (N_15207,N_12819,N_14633);
xor U15208 (N_15208,N_14175,N_12339);
and U15209 (N_15209,N_13816,N_13420);
nor U15210 (N_15210,N_13768,N_12308);
nor U15211 (N_15211,N_12351,N_13143);
nor U15212 (N_15212,N_13801,N_12108);
nor U15213 (N_15213,N_14143,N_12543);
xnor U15214 (N_15214,N_12290,N_13703);
nor U15215 (N_15215,N_14855,N_13550);
and U15216 (N_15216,N_13137,N_14348);
nor U15217 (N_15217,N_13592,N_12976);
or U15218 (N_15218,N_13278,N_14333);
xnor U15219 (N_15219,N_14403,N_13626);
nor U15220 (N_15220,N_12281,N_14125);
nor U15221 (N_15221,N_13908,N_14274);
and U15222 (N_15222,N_13258,N_14958);
and U15223 (N_15223,N_14859,N_14314);
xnor U15224 (N_15224,N_14267,N_12791);
xnor U15225 (N_15225,N_14850,N_12134);
nand U15226 (N_15226,N_13115,N_13098);
or U15227 (N_15227,N_13138,N_12444);
nor U15228 (N_15228,N_14509,N_12749);
and U15229 (N_15229,N_13907,N_14406);
nor U15230 (N_15230,N_13602,N_12622);
nor U15231 (N_15231,N_14010,N_12380);
nand U15232 (N_15232,N_13712,N_13291);
nor U15233 (N_15233,N_14030,N_12321);
nand U15234 (N_15234,N_12871,N_13029);
xnor U15235 (N_15235,N_14932,N_13120);
nand U15236 (N_15236,N_14926,N_13110);
and U15237 (N_15237,N_12792,N_12658);
xor U15238 (N_15238,N_13458,N_13292);
and U15239 (N_15239,N_12313,N_14035);
nor U15240 (N_15240,N_13580,N_14317);
nand U15241 (N_15241,N_14176,N_14022);
nor U15242 (N_15242,N_12010,N_12393);
or U15243 (N_15243,N_13984,N_14337);
nor U15244 (N_15244,N_12268,N_14748);
nand U15245 (N_15245,N_14808,N_12096);
xor U15246 (N_15246,N_12323,N_14319);
nand U15247 (N_15247,N_14804,N_13683);
xnor U15248 (N_15248,N_14849,N_13346);
nand U15249 (N_15249,N_14491,N_13577);
nand U15250 (N_15250,N_13790,N_12884);
xnor U15251 (N_15251,N_12773,N_12542);
xor U15252 (N_15252,N_14361,N_14078);
or U15253 (N_15253,N_14586,N_14258);
and U15254 (N_15254,N_12720,N_13108);
nor U15255 (N_15255,N_12778,N_13666);
and U15256 (N_15256,N_14862,N_13121);
xnor U15257 (N_15257,N_12781,N_14847);
nand U15258 (N_15258,N_14766,N_14579);
nor U15259 (N_15259,N_12162,N_13125);
nor U15260 (N_15260,N_13838,N_13597);
nor U15261 (N_15261,N_14028,N_13113);
nand U15262 (N_15262,N_12751,N_14631);
nand U15263 (N_15263,N_14426,N_13035);
nor U15264 (N_15264,N_13462,N_13269);
xnor U15265 (N_15265,N_12194,N_14979);
and U15266 (N_15266,N_12539,N_12697);
nand U15267 (N_15267,N_13285,N_13235);
xor U15268 (N_15268,N_14559,N_12676);
nand U15269 (N_15269,N_12534,N_12305);
and U15270 (N_15270,N_14318,N_12430);
or U15271 (N_15271,N_14015,N_13583);
xnor U15272 (N_15272,N_13259,N_13165);
and U15273 (N_15273,N_13495,N_13546);
nand U15274 (N_15274,N_13504,N_12798);
nand U15275 (N_15275,N_14505,N_13407);
nor U15276 (N_15276,N_12971,N_13893);
nand U15277 (N_15277,N_12965,N_14309);
nor U15278 (N_15278,N_12437,N_14941);
or U15279 (N_15279,N_13771,N_12926);
nor U15280 (N_15280,N_14867,N_13960);
nor U15281 (N_15281,N_12034,N_13239);
nand U15282 (N_15282,N_13470,N_12219);
xor U15283 (N_15283,N_13237,N_14145);
xor U15284 (N_15284,N_12288,N_14845);
and U15285 (N_15285,N_13926,N_14368);
nand U15286 (N_15286,N_12615,N_12402);
or U15287 (N_15287,N_12789,N_13007);
or U15288 (N_15288,N_14825,N_14674);
or U15289 (N_15289,N_14628,N_14988);
and U15290 (N_15290,N_13310,N_12835);
and U15291 (N_15291,N_14648,N_12875);
nand U15292 (N_15292,N_12311,N_13700);
nor U15293 (N_15293,N_12171,N_14069);
and U15294 (N_15294,N_14820,N_14168);
xor U15295 (N_15295,N_14893,N_12151);
and U15296 (N_15296,N_13208,N_14727);
or U15297 (N_15297,N_12390,N_13465);
and U15298 (N_15298,N_14265,N_13001);
nand U15299 (N_15299,N_12282,N_12808);
xnor U15300 (N_15300,N_13279,N_14497);
nor U15301 (N_15301,N_13754,N_13077);
nand U15302 (N_15302,N_14163,N_12404);
and U15303 (N_15303,N_13367,N_12943);
or U15304 (N_15304,N_12295,N_12361);
or U15305 (N_15305,N_14817,N_14844);
nand U15306 (N_15306,N_14795,N_12685);
and U15307 (N_15307,N_12704,N_12021);
or U15308 (N_15308,N_14000,N_12626);
or U15309 (N_15309,N_13429,N_12092);
nor U15310 (N_15310,N_13141,N_14422);
xor U15311 (N_15311,N_13714,N_13968);
or U15312 (N_15312,N_14955,N_13622);
or U15313 (N_15313,N_14398,N_14528);
or U15314 (N_15314,N_13921,N_13311);
and U15315 (N_15315,N_12725,N_14646);
xor U15316 (N_15316,N_13167,N_14330);
xnor U15317 (N_15317,N_13656,N_13693);
xor U15318 (N_15318,N_12941,N_12896);
nand U15319 (N_15319,N_14560,N_12371);
or U15320 (N_15320,N_14735,N_12718);
nand U15321 (N_15321,N_13639,N_13369);
or U15322 (N_15322,N_12968,N_13906);
and U15323 (N_15323,N_14011,N_12497);
or U15324 (N_15324,N_13756,N_13455);
xor U15325 (N_15325,N_14189,N_12573);
xnor U15326 (N_15326,N_12465,N_12375);
nand U15327 (N_15327,N_14713,N_12852);
and U15328 (N_15328,N_12990,N_13410);
and U15329 (N_15329,N_14277,N_14751);
nand U15330 (N_15330,N_13540,N_14362);
and U15331 (N_15331,N_13277,N_14730);
or U15332 (N_15332,N_13452,N_12748);
xnor U15333 (N_15333,N_12788,N_14066);
and U15334 (N_15334,N_13232,N_14978);
xnor U15335 (N_15335,N_13651,N_14242);
and U15336 (N_15336,N_13571,N_12909);
nor U15337 (N_15337,N_14710,N_13952);
and U15338 (N_15338,N_13609,N_12536);
xor U15339 (N_15339,N_12652,N_14903);
and U15340 (N_15340,N_14266,N_12048);
nand U15341 (N_15341,N_14515,N_12090);
nand U15342 (N_15342,N_14974,N_13032);
and U15343 (N_15343,N_14493,N_14172);
and U15344 (N_15344,N_13294,N_14894);
or U15345 (N_15345,N_13381,N_14815);
and U15346 (N_15346,N_12903,N_13052);
xnor U15347 (N_15347,N_14374,N_14720);
nor U15348 (N_15348,N_13881,N_12991);
and U15349 (N_15349,N_13361,N_12478);
nand U15350 (N_15350,N_13423,N_12002);
nor U15351 (N_15351,N_12498,N_13266);
nand U15352 (N_15352,N_13081,N_14937);
xnor U15353 (N_15353,N_14269,N_14083);
and U15354 (N_15354,N_12262,N_13855);
and U15355 (N_15355,N_12975,N_13691);
and U15356 (N_15356,N_14334,N_12553);
and U15357 (N_15357,N_13153,N_14716);
nor U15358 (N_15358,N_14480,N_12127);
nand U15359 (N_15359,N_12182,N_13966);
xor U15360 (N_15360,N_13281,N_12216);
nor U15361 (N_15361,N_12540,N_12865);
nor U15362 (N_15362,N_13184,N_14547);
or U15363 (N_15363,N_12563,N_12669);
or U15364 (N_15364,N_13603,N_14569);
nand U15365 (N_15365,N_14597,N_14536);
nor U15366 (N_15366,N_12805,N_13566);
and U15367 (N_15367,N_13645,N_14486);
nor U15368 (N_15368,N_14369,N_13697);
nor U15369 (N_15369,N_12828,N_12074);
or U15370 (N_15370,N_14110,N_12771);
xnor U15371 (N_15371,N_12458,N_14326);
nand U15372 (N_15372,N_12972,N_14245);
nor U15373 (N_15373,N_13049,N_12885);
xnor U15374 (N_15374,N_13871,N_12045);
xnor U15375 (N_15375,N_13044,N_14008);
or U15376 (N_15376,N_14842,N_14871);
nand U15377 (N_15377,N_14717,N_12167);
or U15378 (N_15378,N_12970,N_12770);
nor U15379 (N_15379,N_13522,N_14227);
xnor U15380 (N_15380,N_14719,N_13387);
nor U15381 (N_15381,N_12364,N_14431);
or U15382 (N_15382,N_14037,N_12642);
xnor U15383 (N_15383,N_14953,N_13368);
xnor U15384 (N_15384,N_12024,N_14568);
or U15385 (N_15385,N_13657,N_14131);
xnor U15386 (N_15386,N_14376,N_13746);
nand U15387 (N_15387,N_13520,N_13026);
and U15388 (N_15388,N_13435,N_12664);
nand U15389 (N_15389,N_12619,N_13570);
xnor U15390 (N_15390,N_14371,N_12104);
nor U15391 (N_15391,N_13675,N_12521);
xor U15392 (N_15392,N_14439,N_14373);
or U15393 (N_15393,N_13313,N_14784);
nor U15394 (N_15394,N_12649,N_14165);
nand U15395 (N_15395,N_14616,N_14345);
nor U15396 (N_15396,N_13156,N_13565);
nand U15397 (N_15397,N_14991,N_13624);
or U15398 (N_15398,N_12206,N_14563);
nand U15399 (N_15399,N_12397,N_12041);
xor U15400 (N_15400,N_14892,N_12863);
xor U15401 (N_15401,N_12929,N_13528);
and U15402 (N_15402,N_14943,N_12981);
nor U15403 (N_15403,N_12445,N_14782);
and U15404 (N_15404,N_12732,N_13412);
xnor U15405 (N_15405,N_12324,N_14758);
xor U15406 (N_15406,N_14889,N_13449);
nor U15407 (N_15407,N_13956,N_12666);
nand U15408 (N_15408,N_13382,N_14228);
nand U15409 (N_15409,N_13223,N_12101);
nor U15410 (N_15410,N_12000,N_13684);
and U15411 (N_15411,N_12846,N_12736);
or U15412 (N_15412,N_13010,N_12455);
xor U15413 (N_15413,N_12695,N_13811);
xnor U15414 (N_15414,N_12261,N_12988);
or U15415 (N_15415,N_13123,N_12915);
and U15416 (N_15416,N_12541,N_12747);
nand U15417 (N_15417,N_14538,N_14408);
or U15418 (N_15418,N_13183,N_12879);
and U15419 (N_15419,N_13586,N_12567);
or U15420 (N_15420,N_12532,N_13832);
or U15421 (N_15421,N_12843,N_14694);
or U15422 (N_15422,N_14906,N_14447);
or U15423 (N_15423,N_12388,N_14556);
nand U15424 (N_15424,N_13501,N_13051);
and U15425 (N_15425,N_12349,N_12821);
nor U15426 (N_15426,N_12693,N_13883);
and U15427 (N_15427,N_13995,N_14697);
or U15428 (N_15428,N_13024,N_13191);
and U15429 (N_15429,N_14043,N_13231);
or U15430 (N_15430,N_14257,N_14031);
nand U15431 (N_15431,N_12522,N_12777);
and U15432 (N_15432,N_13796,N_12558);
xor U15433 (N_15433,N_14086,N_13594);
and U15434 (N_15434,N_12980,N_12338);
and U15435 (N_15435,N_13692,N_14542);
nor U15436 (N_15436,N_12064,N_13497);
nand U15437 (N_15437,N_13541,N_14800);
or U15438 (N_15438,N_14156,N_12706);
nor U15439 (N_15439,N_14303,N_14209);
or U15440 (N_15440,N_13241,N_13660);
xnor U15441 (N_15441,N_13911,N_12817);
or U15442 (N_15442,N_13558,N_13662);
or U15443 (N_15443,N_14136,N_13752);
or U15444 (N_15444,N_13890,N_13735);
or U15445 (N_15445,N_13377,N_14745);
and U15446 (N_15446,N_13352,N_14549);
nor U15447 (N_15447,N_13305,N_14945);
or U15448 (N_15448,N_12271,N_13561);
nor U15449 (N_15449,N_14632,N_13336);
nand U15450 (N_15450,N_14246,N_12954);
nor U15451 (N_15451,N_14511,N_14260);
nand U15452 (N_15452,N_13870,N_14688);
nor U15453 (N_15453,N_13895,N_12359);
and U15454 (N_15454,N_13129,N_13395);
xor U15455 (N_15455,N_13057,N_13503);
nand U15456 (N_15456,N_13033,N_14525);
nand U15457 (N_15457,N_12136,N_12181);
and U15458 (N_15458,N_13236,N_13744);
xor U15459 (N_15459,N_12431,N_13992);
nand U15460 (N_15460,N_14498,N_14933);
or U15461 (N_15461,N_14148,N_14884);
nor U15462 (N_15462,N_12223,N_14653);
or U15463 (N_15463,N_12501,N_14450);
xor U15464 (N_15464,N_13766,N_14150);
nor U15465 (N_15465,N_14866,N_13197);
and U15466 (N_15466,N_12389,N_12727);
nand U15467 (N_15467,N_14591,N_13357);
xnor U15468 (N_15468,N_13082,N_14876);
and U15469 (N_15469,N_14965,N_12920);
nor U15470 (N_15470,N_13434,N_12411);
nand U15471 (N_15471,N_14805,N_14857);
xnor U15472 (N_15472,N_13364,N_14638);
nor U15473 (N_15473,N_12902,N_12668);
nor U15474 (N_15474,N_12786,N_12930);
or U15475 (N_15475,N_14909,N_12675);
or U15476 (N_15476,N_14916,N_12963);
nor U15477 (N_15477,N_14927,N_13005);
and U15478 (N_15478,N_14581,N_14370);
or U15479 (N_15479,N_14313,N_12274);
or U15480 (N_15480,N_14548,N_13509);
and U15481 (N_15481,N_13679,N_12456);
and U15482 (N_15482,N_12934,N_14651);
nor U15483 (N_15483,N_12953,N_13226);
nor U15484 (N_15484,N_13070,N_12208);
or U15485 (N_15485,N_12439,N_14677);
nand U15486 (N_15486,N_14212,N_14829);
nand U15487 (N_15487,N_12286,N_14773);
xnor U15488 (N_15488,N_12423,N_13371);
nand U15489 (N_15489,N_13489,N_12509);
xor U15490 (N_15490,N_13251,N_13591);
nor U15491 (N_15491,N_13182,N_13783);
nor U15492 (N_15492,N_12503,N_13545);
nand U15493 (N_15493,N_12109,N_13248);
and U15494 (N_15494,N_12121,N_12547);
nor U15495 (N_15495,N_13773,N_12995);
nor U15496 (N_15496,N_12905,N_12050);
nor U15497 (N_15497,N_12204,N_12065);
or U15498 (N_15498,N_14554,N_13175);
xor U15499 (N_15499,N_13103,N_14572);
nor U15500 (N_15500,N_12061,N_13616);
nor U15501 (N_15501,N_13481,N_12327);
and U15502 (N_15502,N_13826,N_14405);
or U15503 (N_15503,N_13390,N_12999);
xnor U15504 (N_15504,N_14899,N_13478);
nor U15505 (N_15505,N_13324,N_13542);
nor U15506 (N_15506,N_13393,N_12605);
or U15507 (N_15507,N_14366,N_12422);
or U15508 (N_15508,N_12660,N_12154);
and U15509 (N_15509,N_14951,N_13724);
xnor U15510 (N_15510,N_12142,N_14520);
and U15511 (N_15511,N_13987,N_13015);
nor U15512 (N_15512,N_12284,N_13466);
and U15513 (N_15513,N_12415,N_14939);
or U15514 (N_15514,N_13902,N_13306);
xnor U15515 (N_15515,N_12461,N_14689);
nand U15516 (N_15516,N_14321,N_12086);
and U15517 (N_15517,N_12709,N_13187);
or U15518 (N_15518,N_13406,N_12705);
nor U15519 (N_15519,N_14149,N_13142);
xor U15520 (N_15520,N_13963,N_13039);
nand U15521 (N_15521,N_12037,N_12960);
nand U15522 (N_15522,N_14420,N_13722);
and U15523 (N_15523,N_12011,N_14691);
xnor U15524 (N_15524,N_14286,N_12647);
and U15525 (N_15525,N_13326,N_12504);
xor U15526 (N_15526,N_12807,N_14506);
and U15527 (N_15527,N_14397,N_14501);
xor U15528 (N_15528,N_13747,N_14169);
nor U15529 (N_15529,N_13341,N_12837);
and U15530 (N_15530,N_13671,N_13830);
nand U15531 (N_15531,N_12514,N_12535);
and U15532 (N_15532,N_14734,N_13654);
xnor U15533 (N_15533,N_13262,N_12039);
nor U15534 (N_15534,N_12743,N_14544);
and U15535 (N_15535,N_14700,N_14822);
and U15536 (N_15536,N_14231,N_13741);
and U15537 (N_15537,N_14438,N_14832);
and U15538 (N_15538,N_13613,N_14381);
xor U15539 (N_15539,N_14552,N_14574);
or U15540 (N_15540,N_12112,N_13200);
nand U15541 (N_15541,N_13217,N_13507);
nand U15542 (N_15542,N_12744,N_12169);
nand U15543 (N_15543,N_12442,N_14229);
nor U15544 (N_15544,N_12318,N_13426);
and U15545 (N_15545,N_12484,N_14473);
nand U15546 (N_15546,N_12607,N_12027);
or U15547 (N_15547,N_14060,N_14736);
nor U15548 (N_15548,N_12130,N_12198);
nand U15549 (N_15549,N_13118,N_13710);
xor U15550 (N_15550,N_13862,N_12047);
and U15551 (N_15551,N_13831,N_12759);
xnor U15552 (N_15552,N_14109,N_13517);
and U15553 (N_15553,N_13394,N_14608);
and U15554 (N_15554,N_14461,N_13563);
and U15555 (N_15555,N_12952,N_13342);
nand U15556 (N_15556,N_13843,N_14396);
nor U15557 (N_15557,N_13718,N_13795);
nor U15558 (N_15558,N_14686,N_12518);
or U15559 (N_15559,N_14492,N_14929);
and U15560 (N_15560,N_14901,N_12060);
nor U15561 (N_15561,N_14489,N_13864);
or U15562 (N_15562,N_13446,N_13221);
or U15563 (N_15563,N_13549,N_13409);
xor U15564 (N_15564,N_13601,N_13272);
and U15565 (N_15565,N_13402,N_12146);
nor U15566 (N_15566,N_14173,N_13047);
nor U15567 (N_15567,N_14532,N_14017);
and U15568 (N_15568,N_14503,N_13366);
nand U15569 (N_15569,N_13776,N_12739);
or U15570 (N_15570,N_13874,N_14928);
and U15571 (N_15571,N_13983,N_12054);
or U15572 (N_15572,N_13308,N_13450);
nand U15573 (N_15573,N_14539,N_12761);
and U15574 (N_15574,N_14404,N_13944);
nor U15575 (N_15575,N_12029,N_14630);
nor U15576 (N_15576,N_12620,N_12077);
nor U15577 (N_15577,N_12958,N_13686);
nand U15578 (N_15578,N_13105,N_13538);
xor U15579 (N_15579,N_13014,N_14660);
xnor U15580 (N_15580,N_13351,N_13585);
nand U15581 (N_15581,N_12758,N_12717);
nor U15582 (N_15582,N_14726,N_14202);
and U15583 (N_15583,N_14890,N_13498);
or U15584 (N_15584,N_13687,N_14589);
xnor U15585 (N_15585,N_13205,N_13823);
nor U15586 (N_15586,N_12710,N_14819);
or U15587 (N_15587,N_12488,N_14877);
xor U15588 (N_15588,N_12435,N_13946);
nor U15589 (N_15589,N_14275,N_14789);
xor U15590 (N_15590,N_13508,N_14806);
nand U15591 (N_15591,N_13694,N_14526);
or U15592 (N_15592,N_14073,N_12590);
and U15593 (N_15593,N_14276,N_14272);
or U15594 (N_15594,N_13084,N_12650);
xor U15595 (N_15595,N_14797,N_13080);
nor U15596 (N_15596,N_13287,N_13701);
or U15597 (N_15597,N_14023,N_14522);
nand U15598 (N_15598,N_14747,N_12183);
xor U15599 (N_15599,N_14259,N_14108);
nand U15600 (N_15600,N_12687,N_13031);
nor U15601 (N_15601,N_14123,N_12969);
and U15602 (N_15602,N_14659,N_13981);
nand U15603 (N_15603,N_12653,N_13531);
or U15604 (N_15604,N_12495,N_12317);
nand U15605 (N_15605,N_12623,N_12278);
xnor U15606 (N_15606,N_14235,N_14625);
xnor U15607 (N_15607,N_14705,N_12394);
and U15608 (N_15608,N_12260,N_13380);
nor U15609 (N_15609,N_13362,N_14298);
nand U15610 (N_15610,N_14793,N_13356);
nor U15611 (N_15611,N_14938,N_13877);
and U15612 (N_15612,N_12125,N_14247);
nand U15613 (N_15613,N_12937,N_13774);
or U15614 (N_15614,N_13792,N_12414);
nor U15615 (N_15615,N_13999,N_13730);
or U15616 (N_15616,N_14540,N_13271);
or U15617 (N_15617,N_14025,N_12384);
or U15618 (N_15618,N_12728,N_12838);
or U15619 (N_15619,N_13685,N_14551);
nor U15620 (N_15620,N_12492,N_12724);
xnor U15621 (N_15621,N_13145,N_12110);
nand U15622 (N_15622,N_13284,N_14455);
nand U15623 (N_15623,N_14407,N_13327);
nand U15624 (N_15624,N_13468,N_14042);
and U15625 (N_15625,N_13642,N_14412);
nand U15626 (N_15626,N_13629,N_14508);
xor U15627 (N_15627,N_12409,N_13042);
nand U15628 (N_15628,N_13536,N_13488);
nor U15629 (N_15629,N_12924,N_12528);
or U15630 (N_15630,N_14529,N_13347);
nor U15631 (N_15631,N_14446,N_12046);
nor U15632 (N_15632,N_13767,N_12689);
and U15633 (N_15633,N_12433,N_12485);
nor U15634 (N_15634,N_13073,N_14585);
or U15635 (N_15635,N_14872,N_14200);
nand U15636 (N_15636,N_14833,N_12836);
and U15637 (N_15637,N_14831,N_14207);
xor U15638 (N_15638,N_14912,N_12464);
and U15639 (N_15639,N_14399,N_12036);
nand U15640 (N_15640,N_13094,N_13300);
or U15641 (N_15641,N_14853,N_12117);
nor U15642 (N_15642,N_12564,N_14913);
nor U15643 (N_15643,N_13194,N_13030);
xor U15644 (N_15644,N_12967,N_14690);
nor U15645 (N_15645,N_12247,N_12333);
nor U15646 (N_15646,N_14270,N_13959);
nand U15647 (N_15647,N_13726,N_12466);
and U15648 (N_15648,N_14129,N_13268);
nor U15649 (N_15649,N_13682,N_12446);
or U15650 (N_15650,N_14485,N_14652);
xor U15651 (N_15651,N_13345,N_13800);
nor U15652 (N_15652,N_12042,N_13290);
and U15653 (N_15653,N_13456,N_14530);
and U15654 (N_15654,N_14972,N_12562);
nand U15655 (N_15655,N_12193,N_14701);
and U15656 (N_15656,N_12354,N_12595);
nor U15657 (N_15657,N_14192,N_12191);
xor U15658 (N_15658,N_14087,N_12382);
and U15659 (N_15659,N_12159,N_13514);
nor U15660 (N_15660,N_13579,N_12150);
xnor U15661 (N_15661,N_13582,N_12225);
nand U15662 (N_15662,N_13350,N_12602);
nand U15663 (N_15663,N_14013,N_14698);
xnor U15664 (N_15664,N_13846,N_13667);
xnor U15665 (N_15665,N_14271,N_14127);
nor U15666 (N_15666,N_13496,N_13427);
and U15667 (N_15667,N_14107,N_12457);
and U15668 (N_15668,N_14496,N_13535);
or U15669 (N_15669,N_13909,N_12933);
nor U15670 (N_15670,N_13062,N_14863);
nand U15671 (N_15671,N_12878,N_13631);
or U15672 (N_15672,N_14284,N_12221);
xor U15673 (N_15673,N_13490,N_12447);
nor U15674 (N_15674,N_12355,N_14478);
xnor U15675 (N_15675,N_13873,N_14614);
xnor U15676 (N_15676,N_14287,N_13471);
nand U15677 (N_15677,N_13201,N_14056);
or U15678 (N_15678,N_12347,N_12330);
nand U15679 (N_15679,N_14448,N_12189);
and U15680 (N_15680,N_13365,N_14320);
nand U15681 (N_15681,N_12005,N_14311);
nor U15682 (N_15682,N_13699,N_12322);
or U15683 (N_15683,N_13562,N_14807);
nor U15684 (N_15684,N_13392,N_12517);
nor U15685 (N_15685,N_12145,N_13706);
nand U15686 (N_15686,N_14742,N_13872);
and U15687 (N_15687,N_12358,N_13419);
xnor U15688 (N_15688,N_13765,N_13155);
nand U15689 (N_15689,N_13689,N_13100);
xnor U15690 (N_15690,N_12166,N_13897);
or U15691 (N_15691,N_12094,N_13958);
or U15692 (N_15692,N_13927,N_14908);
and U15693 (N_15693,N_14858,N_14555);
nand U15694 (N_15694,N_13524,N_12287);
nand U15695 (N_15695,N_13303,N_13499);
or U15696 (N_15696,N_12063,N_14562);
nor U15697 (N_15697,N_13933,N_12494);
and U15698 (N_15698,N_12184,N_12874);
xor U15699 (N_15699,N_12467,N_14981);
nand U15700 (N_15700,N_12849,N_14316);
xor U15701 (N_15701,N_12078,N_13739);
or U15702 (N_15702,N_14640,N_12899);
nor U15703 (N_15703,N_14919,N_14372);
nand U15704 (N_15704,N_12148,N_14053);
nand U15705 (N_15705,N_12405,N_13213);
nor U15706 (N_15706,N_12796,N_12606);
and U15707 (N_15707,N_13793,N_14208);
or U15708 (N_15708,N_13457,N_14774);
xnor U15709 (N_15709,N_13560,N_14293);
nand U15710 (N_15710,N_14612,N_12812);
xnor U15711 (N_15711,N_14788,N_12707);
nand U15712 (N_15712,N_13615,N_12003);
xor U15713 (N_15713,N_12919,N_13617);
nor U15714 (N_15714,N_12453,N_12892);
or U15715 (N_15715,N_13915,N_13180);
xor U15716 (N_15716,N_14783,N_13106);
and U15717 (N_15717,N_14851,N_14886);
xnor U15718 (N_15718,N_13569,N_12132);
and U15719 (N_15719,N_14865,N_14418);
xor U15720 (N_15720,N_13132,N_12641);
nand U15721 (N_15721,N_13721,N_14954);
nand U15722 (N_15722,N_12100,N_14142);
xnor U15723 (N_15723,N_13122,N_13977);
nand U15724 (N_15724,N_14236,N_12701);
or U15725 (N_15725,N_13162,N_13009);
or U15726 (N_15726,N_12723,N_12499);
nor U15727 (N_15727,N_12214,N_12586);
nor U15728 (N_15728,N_14211,N_14786);
or U15729 (N_15729,N_14364,N_13091);
and U15730 (N_15730,N_13166,N_14048);
or U15731 (N_15731,N_14051,N_12681);
or U15732 (N_15732,N_14523,N_12715);
and U15733 (N_15733,N_13931,N_13551);
xnor U15734 (N_15734,N_12451,N_12731);
and U15735 (N_15735,N_13140,N_14521);
nand U15736 (N_15736,N_12115,N_14402);
or U15737 (N_15737,N_14869,N_14400);
nor U15738 (N_15738,N_13653,N_14882);
or U15739 (N_15739,N_13186,N_14852);
nor U15740 (N_15740,N_14779,N_14722);
xnor U15741 (N_15741,N_14178,N_13243);
xor U15742 (N_15742,N_14527,N_13620);
and U15743 (N_15743,N_14248,N_12538);
or U15744 (N_15744,N_12734,N_14636);
nand U15745 (N_15745,N_12914,N_12277);
nor U15746 (N_15746,N_13136,N_13097);
nor U15747 (N_15747,N_12913,N_14262);
xnor U15748 (N_15748,N_13729,N_14380);
nor U15749 (N_15749,N_14183,N_12672);
or U15750 (N_15750,N_14294,N_14186);
nor U15751 (N_15751,N_13533,N_13376);
xor U15752 (N_15752,N_12350,N_12557);
and U15753 (N_15753,N_13119,N_13477);
xor U15754 (N_15754,N_14454,N_12336);
or U15755 (N_15755,N_14117,N_14992);
and U15756 (N_15756,N_13006,N_12477);
or U15757 (N_15757,N_14692,N_13819);
xnor U15758 (N_15758,N_13738,N_14395);
nand U15759 (N_15759,N_13230,N_12479);
xor U15760 (N_15760,N_12574,N_13716);
or U15761 (N_15761,N_13511,N_13370);
nand U15762 (N_15762,N_12242,N_14089);
or U15763 (N_15763,N_13812,N_14456);
nand U15764 (N_15764,N_14504,N_12505);
and U15765 (N_15765,N_13993,N_13034);
and U15766 (N_15766,N_13510,N_13092);
and U15767 (N_15767,N_12009,N_14327);
nor U15768 (N_15768,N_14464,N_14963);
xor U15769 (N_15769,N_13593,N_14930);
nor U15770 (N_15770,N_12755,N_13543);
and U15771 (N_15771,N_14024,N_14746);
or U15772 (N_15772,N_13078,N_12601);
nand U15773 (N_15773,N_12927,N_14944);
xor U15774 (N_15774,N_14607,N_13333);
and U15775 (N_15775,N_12643,N_12168);
or U15776 (N_15776,N_12436,N_13676);
xnor U15777 (N_15777,N_14096,N_13702);
xnor U15778 (N_15778,N_12158,N_14133);
nand U15779 (N_15779,N_12269,N_13806);
and U15780 (N_15780,N_14743,N_12571);
and U15781 (N_15781,N_12018,N_12314);
and U15782 (N_15782,N_14198,N_13552);
or U15783 (N_15783,N_14613,N_14623);
or U15784 (N_15784,N_12636,N_12377);
nand U15785 (N_15785,N_12679,N_14072);
nand U15786 (N_15786,N_12001,N_13673);
nor U15787 (N_15787,N_12712,N_14092);
or U15788 (N_15788,N_14305,N_12300);
xor U15789 (N_15789,N_14481,N_14592);
xor U15790 (N_15790,N_13578,N_12655);
nor U15791 (N_15791,N_14902,N_12596);
xor U15792 (N_15792,N_12123,N_14888);
and U15793 (N_15793,N_12263,N_14961);
nand U15794 (N_15794,N_13868,N_13206);
xnor U15795 (N_15795,N_13863,N_13202);
nor U15796 (N_15796,N_12917,N_12797);
nand U15797 (N_15797,N_12684,N_13777);
nor U15798 (N_15798,N_14683,N_12212);
and U15799 (N_15799,N_13093,N_12428);
nand U15800 (N_15800,N_13920,N_14533);
xnor U15801 (N_15801,N_13901,N_14475);
and U15802 (N_15802,N_12856,N_12683);
xor U15803 (N_15803,N_13331,N_14322);
xor U15804 (N_15804,N_14969,N_13065);
nand U15805 (N_15805,N_13815,N_12400);
nor U15806 (N_15806,N_14411,N_13947);
and U15807 (N_15807,N_12017,N_13315);
nor U15808 (N_15808,N_14976,N_13564);
nand U15809 (N_15809,N_13632,N_14077);
and U15810 (N_15810,N_14104,N_14502);
nor U15811 (N_15811,N_12631,N_13418);
nand U15812 (N_15812,N_12031,N_12334);
nor U15813 (N_15813,N_12901,N_12639);
and U15814 (N_15814,N_13072,N_12839);
xor U15815 (N_15815,N_13865,N_12938);
nand U15816 (N_15816,N_13708,N_13437);
nor U15817 (N_15817,N_12459,N_12719);
or U15818 (N_15818,N_14114,N_14995);
xnor U15819 (N_15819,N_12775,N_13441);
nor U15820 (N_15820,N_12722,N_14134);
or U15821 (N_15821,N_14546,N_12113);
nor U15822 (N_15822,N_12418,N_13041);
nand U15823 (N_15823,N_12237,N_14476);
and U15824 (N_15824,N_13788,N_12147);
nand U15825 (N_15825,N_13951,N_12363);
nor U15826 (N_15826,N_13195,N_12443);
or U15827 (N_15827,N_13492,N_14254);
nor U15828 (N_15828,N_14041,N_12376);
or U15829 (N_15829,N_12490,N_14561);
nor U15830 (N_15830,N_12946,N_13181);
or U15831 (N_15831,N_12531,N_13709);
and U15832 (N_15832,N_13486,N_12138);
nand U15833 (N_15833,N_14470,N_12353);
and U15834 (N_15834,N_13717,N_12910);
nand U15835 (N_15835,N_13763,N_13556);
or U15836 (N_15836,N_13431,N_12475);
xnor U15837 (N_15837,N_14199,N_12813);
nand U15838 (N_15838,N_12673,N_13505);
and U15839 (N_15839,N_14975,N_13939);
and U15840 (N_15840,N_14900,N_13319);
nor U15841 (N_15841,N_14641,N_13869);
and U15842 (N_15842,N_13674,N_13320);
nand U15843 (N_15843,N_12205,N_12429);
xnor U15844 (N_15844,N_14768,N_12985);
xor U15845 (N_15845,N_12152,N_12283);
nand U15846 (N_15846,N_13844,N_13375);
and U15847 (N_15847,N_12131,N_14014);
nand U15848 (N_15848,N_14606,N_12057);
nand U15849 (N_15849,N_12266,N_13957);
xnor U15850 (N_15850,N_13479,N_14355);
nand U15851 (N_15851,N_12463,N_12599);
and U15852 (N_15852,N_14967,N_13723);
xor U15853 (N_15853,N_13567,N_14879);
xor U15854 (N_15854,N_14545,N_14898);
nand U15855 (N_15855,N_12040,N_14102);
or U15856 (N_15856,N_14467,N_12959);
nand U15857 (N_15857,N_13019,N_13769);
or U15858 (N_15858,N_12255,N_14576);
nor U15859 (N_15859,N_13104,N_14425);
nand U15860 (N_15860,N_12381,N_12095);
and U15861 (N_15861,N_12921,N_12211);
or U15862 (N_15862,N_14225,N_13923);
or U15863 (N_15863,N_14621,N_14295);
or U15864 (N_15864,N_12936,N_13523);
xor U15865 (N_15865,N_12091,N_12783);
or U15866 (N_15866,N_12637,N_12254);
nor U15867 (N_15867,N_12951,N_13814);
or U15868 (N_15868,N_12291,N_13304);
and U15869 (N_15869,N_14672,N_13473);
nand U15870 (N_15870,N_13834,N_12141);
and U15871 (N_15871,N_12473,N_14531);
nor U15872 (N_15872,N_12298,N_12025);
or U15873 (N_15873,N_13555,N_12076);
xor U15874 (N_15874,N_13967,N_12827);
nand U15875 (N_15875,N_14195,N_14667);
nor U15876 (N_15876,N_12250,N_13929);
and U15877 (N_15877,N_12016,N_14413);
or U15878 (N_15878,N_12694,N_12549);
or U15879 (N_15879,N_12940,N_13107);
nand U15880 (N_15880,N_12868,N_12634);
nand U15881 (N_15881,N_13860,N_14739);
nand U15882 (N_15882,N_14058,N_12105);
and U15883 (N_15883,N_13753,N_14517);
and U15884 (N_15884,N_12861,N_13633);
xor U15885 (N_15885,N_13330,N_12089);
xnor U15886 (N_15886,N_13391,N_13867);
nor U15887 (N_15887,N_14139,N_12588);
nor U15888 (N_15888,N_14999,N_13460);
nor U15889 (N_15889,N_12227,N_13998);
nor U15890 (N_15890,N_14693,N_12889);
or U15891 (N_15891,N_12795,N_13500);
nor U15892 (N_15892,N_13600,N_14662);
xnor U15893 (N_15893,N_14801,N_13257);
and U15894 (N_15894,N_13440,N_14622);
nor U15895 (N_15895,N_14363,N_12654);
or U15896 (N_15896,N_13994,N_12007);
or U15897 (N_15897,N_14307,N_12222);
xnor U15898 (N_15898,N_13373,N_12257);
nand U15899 (N_15899,N_14282,N_14429);
and U15900 (N_15900,N_12545,N_12548);
nand U15901 (N_15901,N_14873,N_14340);
or U15902 (N_15902,N_14973,N_13775);
and U15903 (N_15903,N_13835,N_12667);
xor U15904 (N_15904,N_13256,N_14904);
nand U15905 (N_15905,N_14427,N_13854);
xnor U15906 (N_15906,N_13133,N_13348);
nor U15907 (N_15907,N_14479,N_14767);
and U15908 (N_15908,N_13698,N_13413);
nand U15909 (N_15909,N_12203,N_13945);
xnor U15910 (N_15910,N_14816,N_14382);
or U15911 (N_15911,N_12591,N_12855);
xor U15912 (N_15912,N_13340,N_13572);
xor U15913 (N_15913,N_12472,N_13172);
xnor U15914 (N_15914,N_14840,N_12346);
xnor U15915 (N_15915,N_14994,N_12107);
nor U15916 (N_15916,N_13058,N_13619);
nor U15917 (N_15917,N_14215,N_13307);
and U15918 (N_15918,N_13762,N_13997);
or U15919 (N_15919,N_13758,N_14392);
xor U15920 (N_15920,N_13914,N_14626);
nor U15921 (N_15921,N_13250,N_12302);
nor U15922 (N_15922,N_13842,N_12957);
or U15923 (N_15923,N_14205,N_13264);
xor U15924 (N_15924,N_14005,N_13848);
nor U15925 (N_15925,N_13283,N_12120);
nand U15926 (N_15926,N_12677,N_12006);
nand U15927 (N_15927,N_13075,N_12128);
nand U15928 (N_15928,N_12721,N_12192);
xnor U15929 (N_15929,N_13253,N_13557);
xnor U15930 (N_15930,N_14201,N_12582);
nor U15931 (N_15931,N_13487,N_14306);
nor U15932 (N_15932,N_13389,N_12392);
and U15933 (N_15933,N_12616,N_12502);
xnor U15934 (N_15934,N_13018,N_12928);
nor U15935 (N_15935,N_13480,N_13695);
and U15936 (N_15936,N_13821,N_13904);
nor U15937 (N_15937,N_14685,N_13553);
xor U15938 (N_15938,N_12556,N_14158);
nand U15939 (N_15939,N_12093,N_12177);
nand U15940 (N_15940,N_13894,N_12226);
nor U15941 (N_15941,N_12580,N_13453);
nand U15942 (N_15942,N_14949,N_14682);
xnor U15943 (N_15943,N_14222,N_12356);
and U15944 (N_15944,N_13233,N_14027);
and U15945 (N_15945,N_14070,N_14090);
xor U15946 (N_15946,N_14378,N_14206);
xnor U15947 (N_15947,N_14458,N_14401);
nor U15948 (N_15948,N_13975,N_12632);
or U15949 (N_15949,N_12408,N_12698);
xor U15950 (N_15950,N_14920,N_13755);
xnor U15951 (N_15951,N_13411,N_14980);
nand U15952 (N_15952,N_14098,N_14002);
xnor U15953 (N_15953,N_13199,N_12947);
xor U15954 (N_15954,N_14105,N_13610);
and U15955 (N_15955,N_14219,N_14776);
or U15956 (N_15956,N_14673,N_13532);
and U15957 (N_15957,N_14358,N_13757);
nor U15958 (N_15958,N_14665,N_12908);
and U15959 (N_15959,N_12201,N_14687);
xnor U15960 (N_15960,N_14304,N_14440);
and U15961 (N_15961,N_12299,N_12233);
nor U15962 (N_15962,N_12081,N_12275);
nor U15963 (N_15963,N_14324,N_14856);
and U15964 (N_15964,N_13249,N_13130);
nor U15965 (N_15965,N_12470,N_12942);
xnor U15966 (N_15966,N_14864,N_12742);
xnor U15967 (N_15967,N_12460,N_13882);
nand U15968 (N_15968,N_14500,N_14111);
and U15969 (N_15969,N_14897,N_13064);
nor U15970 (N_15970,N_12401,N_13941);
nor U15971 (N_15971,N_12912,N_12630);
xor U15972 (N_15972,N_13797,N_14441);
xor U15973 (N_15973,N_14600,N_12240);
or U15974 (N_15974,N_12897,N_13150);
nand U15975 (N_15975,N_13934,N_12611);
or U15976 (N_15976,N_14034,N_13385);
nor U15977 (N_15977,N_12315,N_12992);
nand U15978 (N_15978,N_12956,N_12644);
xor U15979 (N_15979,N_12551,N_12873);
or U15980 (N_15980,N_13134,N_13050);
or U15981 (N_15981,N_14160,N_12365);
xnor U15982 (N_15982,N_13574,N_12600);
nor U15983 (N_15983,N_12628,N_14733);
and U15984 (N_15984,N_13171,N_13144);
and U15985 (N_15985,N_14948,N_12585);
and U15986 (N_15986,N_14460,N_13483);
and U15987 (N_15987,N_13055,N_13530);
and U15988 (N_15988,N_12978,N_12155);
nand U15989 (N_15989,N_14232,N_12008);
or U15990 (N_15990,N_14091,N_12352);
nand U15991 (N_15991,N_13969,N_12617);
xor U15992 (N_15992,N_14763,N_14650);
and U15993 (N_15993,N_14417,N_13905);
xor U15994 (N_15994,N_13344,N_12213);
nand U15995 (N_15995,N_12407,N_14451);
and U15996 (N_15996,N_12229,N_12396);
or U15997 (N_15997,N_13916,N_14224);
nor U15998 (N_15998,N_14243,N_12893);
xor U15999 (N_15999,N_14283,N_14377);
or U16000 (N_16000,N_12840,N_13432);
xnor U16001 (N_16001,N_12215,N_13276);
and U16002 (N_16002,N_14737,N_13899);
nand U16003 (N_16003,N_13537,N_14834);
nand U16004 (N_16004,N_14416,N_12028);
xnor U16005 (N_16005,N_13238,N_13048);
nor U16006 (N_16006,N_12069,N_12974);
or U16007 (N_16007,N_13494,N_13936);
xnor U16008 (N_16008,N_14617,N_12584);
nand U16009 (N_16009,N_14785,N_12906);
xnor U16010 (N_16010,N_13745,N_12589);
and U16011 (N_16011,N_14055,N_12872);
xnor U16012 (N_16012,N_14759,N_14443);
nor U16013 (N_16013,N_14214,N_13074);
nor U16014 (N_16014,N_14241,N_13234);
or U16015 (N_16015,N_14905,N_14821);
or U16016 (N_16016,N_13247,N_13439);
nor U16017 (N_16017,N_12870,N_13974);
and U16018 (N_16018,N_14193,N_13903);
nor U16019 (N_16019,N_13227,N_13502);
or U16020 (N_16020,N_14387,N_13328);
nand U16021 (N_16021,N_13791,N_13430);
nand U16022 (N_16022,N_12395,N_12116);
xor U16023 (N_16023,N_12713,N_12099);
nor U16024 (N_16024,N_12253,N_13163);
and U16025 (N_16025,N_12440,N_14775);
nor U16026 (N_16026,N_13260,N_12746);
nand U16027 (N_16027,N_14952,N_12898);
xnor U16028 (N_16028,N_13301,N_14885);
or U16029 (N_16029,N_13443,N_13805);
nor U16030 (N_16030,N_12854,N_12144);
and U16031 (N_16031,N_12572,N_12876);
and U16032 (N_16032,N_14188,N_13160);
nand U16033 (N_16033,N_13448,N_13761);
or U16034 (N_16034,N_13095,N_14732);
xor U16035 (N_16035,N_12784,N_12406);
xor U16036 (N_16036,N_14619,N_12419);
nand U16037 (N_16037,N_14121,N_12071);
or U16038 (N_16038,N_12859,N_13751);
xor U16039 (N_16039,N_12831,N_14772);
nor U16040 (N_16040,N_13847,N_13396);
nand U16041 (N_16041,N_14063,N_14445);
or U16042 (N_16042,N_13587,N_14329);
and U16043 (N_16043,N_14328,N_14166);
and U16044 (N_16044,N_13322,N_13759);
or U16045 (N_16045,N_14558,N_12587);
nand U16046 (N_16046,N_13164,N_13189);
nand U16047 (N_16047,N_12398,N_13334);
nand U16048 (N_16048,N_14765,N_14935);
or U16049 (N_16049,N_13360,N_12729);
or U16050 (N_16050,N_12337,N_12304);
or U16051 (N_16051,N_14896,N_13925);
and U16052 (N_16052,N_12638,N_13146);
nand U16053 (N_16053,N_14488,N_12659);
xor U16054 (N_16054,N_12372,N_14047);
xor U16055 (N_16055,N_14177,N_12163);
nor U16056 (N_16056,N_14138,N_13036);
or U16057 (N_16057,N_14671,N_12754);
xor U16058 (N_16058,N_14261,N_12462);
nand U16059 (N_16059,N_14643,N_13932);
and U16060 (N_16060,N_14836,N_12691);
and U16061 (N_16061,N_14588,N_13083);
and U16062 (N_16062,N_12671,N_12102);
nor U16063 (N_16063,N_13003,N_12106);
xnor U16064 (N_16064,N_14130,N_12450);
or U16065 (N_16065,N_12948,N_12989);
nand U16066 (N_16066,N_12583,N_12987);
and U16067 (N_16067,N_12814,N_14349);
nand U16068 (N_16068,N_13002,N_12686);
xor U16069 (N_16069,N_13417,N_14196);
nand U16070 (N_16070,N_14182,N_13851);
nor U16071 (N_16071,N_13875,N_12083);
nand U16072 (N_16072,N_14394,N_12841);
and U16073 (N_16073,N_13149,N_13688);
and U16074 (N_16074,N_14449,N_12853);
nand U16075 (N_16075,N_12566,N_12756);
and U16076 (N_16076,N_13086,N_13785);
or U16077 (N_16077,N_12143,N_14103);
nor U16078 (N_16078,N_13780,N_12452);
nor U16079 (N_16079,N_13732,N_12533);
or U16080 (N_16080,N_12051,N_13359);
and U16081 (N_16081,N_14644,N_12833);
or U16082 (N_16082,N_13858,N_13386);
nor U16083 (N_16083,N_12883,N_14101);
nor U16084 (N_16084,N_13464,N_13892);
and U16085 (N_16085,N_14609,N_12785);
nor U16086 (N_16086,N_14880,N_12961);
nand U16087 (N_16087,N_13681,N_13192);
xor U16088 (N_16088,N_13069,N_12197);
xnor U16089 (N_16089,N_14187,N_13244);
and U16090 (N_16090,N_13850,N_12982);
or U16091 (N_16091,N_14472,N_13828);
nand U16092 (N_16092,N_14001,N_13515);
nor U16093 (N_16093,N_14062,N_13544);
xor U16094 (N_16094,N_13827,N_14213);
nor U16095 (N_16095,N_13859,N_14290);
and U16096 (N_16096,N_13020,N_13317);
and U16097 (N_16097,N_14777,N_12964);
nand U16098 (N_16098,N_12500,N_14499);
and U16099 (N_16099,N_13397,N_13980);
or U16100 (N_16100,N_14940,N_13961);
or U16101 (N_16101,N_12916,N_13161);
nand U16102 (N_16102,N_13043,N_14057);
xor U16103 (N_16103,N_12328,N_12803);
nand U16104 (N_16104,N_12164,N_14565);
nand U16105 (N_16105,N_12648,N_14263);
xnor U16106 (N_16106,N_12516,N_14557);
and U16107 (N_16107,N_14410,N_14618);
nor U16108 (N_16108,N_12772,N_14281);
nand U16109 (N_16109,N_14738,N_13013);
and U16110 (N_16110,N_14434,N_14302);
and U16111 (N_16111,N_12665,N_13054);
and U16112 (N_16112,N_14668,N_12469);
nand U16113 (N_16113,N_14007,N_12925);
nand U16114 (N_16114,N_13066,N_12997);
xnor U16115 (N_16115,N_14240,N_14221);
xor U16116 (N_16116,N_14875,N_12894);
nand U16117 (N_16117,N_13568,N_13948);
nor U16118 (N_16118,N_12537,N_12280);
nand U16119 (N_16119,N_14537,N_12267);
nor U16120 (N_16120,N_12329,N_12157);
nor U16121 (N_16121,N_14512,N_14393);
nand U16122 (N_16122,N_14507,N_14118);
and U16123 (N_16123,N_14484,N_13433);
nand U16124 (N_16124,N_12342,N_12026);
xor U16125 (N_16125,N_13588,N_14998);
nand U16126 (N_16126,N_14204,N_12782);
and U16127 (N_16127,N_13314,N_12368);
nor U16128 (N_16128,N_14040,N_13646);
and U16129 (N_16129,N_14846,N_12663);
and U16130 (N_16130,N_14170,N_12199);
and U16131 (N_16131,N_14841,N_13928);
nand U16132 (N_16132,N_13937,N_13261);
xnor U16133 (N_16133,N_12279,N_14421);
and U16134 (N_16134,N_13099,N_13982);
or U16135 (N_16135,N_12735,N_12236);
nor U16136 (N_16136,N_14584,N_14580);
xnor U16137 (N_16137,N_14582,N_12410);
nor U16138 (N_16138,N_12186,N_14635);
nand U16139 (N_16139,N_13135,N_12618);
nor U16140 (N_16140,N_13887,N_13809);
nand U16141 (N_16141,N_12512,N_14987);
nor U16142 (N_16142,N_14181,N_12441);
and U16143 (N_16143,N_14115,N_13088);
and U16144 (N_16144,N_14419,N_13338);
nor U16145 (N_16145,N_12344,N_14715);
or U16146 (N_16146,N_14570,N_13484);
and U16147 (N_16147,N_12481,N_13339);
xor U16148 (N_16148,N_13459,N_14762);
nor U16149 (N_16149,N_14065,N_13720);
or U16150 (N_16150,N_13388,N_14818);
and U16151 (N_16151,N_13962,N_13910);
xor U16152 (N_16152,N_14080,N_12316);
nand U16153 (N_16153,N_12249,N_13659);
and U16154 (N_16154,N_13711,N_13803);
nand U16155 (N_16155,N_13343,N_14296);
nor U16156 (N_16156,N_13169,N_13648);
nor U16157 (N_16157,N_14038,N_14093);
nor U16158 (N_16158,N_12022,N_14469);
nor U16159 (N_16159,N_14519,N_13554);
nand U16160 (N_16160,N_14315,N_13526);
and U16161 (N_16161,N_12678,N_12224);
xnor U16162 (N_16162,N_12165,N_12196);
nand U16163 (N_16163,N_14153,N_12489);
nor U16164 (N_16164,N_14435,N_13810);
and U16165 (N_16165,N_14487,N_12035);
xor U16166 (N_16166,N_12427,N_14921);
nor U16167 (N_16167,N_13154,N_14984);
or U16168 (N_16168,N_13782,N_13282);
nand U16169 (N_16169,N_14989,N_12103);
nor U16170 (N_16170,N_14124,N_12604);
nor U16171 (N_16171,N_12609,N_13589);
nor U16172 (N_16172,N_13627,N_12612);
and U16173 (N_16173,N_13748,N_13818);
xor U16174 (N_16174,N_13063,N_12053);
nor U16175 (N_16175,N_12483,N_13289);
nor U16176 (N_16176,N_12598,N_14827);
and U16177 (N_16177,N_14185,N_12973);
xor U16178 (N_16178,N_13839,N_12882);
nand U16179 (N_16179,N_13405,N_14649);
xor U16180 (N_16180,N_13363,N_12847);
nor U16181 (N_16181,N_12412,N_12768);
nor U16182 (N_16182,N_12161,N_13614);
nand U16183 (N_16183,N_12272,N_13461);
xnor U16184 (N_16184,N_14611,N_14605);
and U16185 (N_16185,N_13861,N_14174);
or U16186 (N_16186,N_14823,N_14299);
and U16187 (N_16187,N_13985,N_12385);
nand U16188 (N_16188,N_14297,N_12891);
xor U16189 (N_16189,N_14740,N_14970);
and U16190 (N_16190,N_13008,N_14161);
or U16191 (N_16191,N_12140,N_13027);
nand U16192 (N_16192,N_12468,N_14021);
or U16193 (N_16193,N_14679,N_13037);
nand U16194 (N_16194,N_12487,N_14566);
and U16195 (N_16195,N_12737,N_13612);
nor U16196 (N_16196,N_14601,N_14003);
or U16197 (N_16197,N_13384,N_12767);
xor U16198 (N_16198,N_14968,N_12700);
nand U16199 (N_16199,N_14135,N_12383);
nand U16200 (N_16200,N_12523,N_13852);
nor U16201 (N_16201,N_12793,N_14878);
xnor U16202 (N_16202,N_13267,N_12787);
and U16203 (N_16203,N_13635,N_13193);
or U16204 (N_16204,N_13590,N_12209);
nor U16205 (N_16205,N_13101,N_12661);
xnor U16206 (N_16206,N_12844,N_13424);
xnor U16207 (N_16207,N_14934,N_13060);
xor U16208 (N_16208,N_12243,N_12682);
and U16209 (N_16209,N_13733,N_13853);
and U16210 (N_16210,N_14911,N_14074);
and U16211 (N_16211,N_14218,N_13584);
or U16212 (N_16212,N_13719,N_13068);
xor U16213 (N_16213,N_13022,N_12234);
nand U16214 (N_16214,N_12993,N_13940);
xor U16215 (N_16215,N_14351,N_12579);
and U16216 (N_16216,N_14848,N_12830);
xnor U16217 (N_16217,N_12062,N_14828);
or U16218 (N_16218,N_14430,N_12949);
and U16219 (N_16219,N_12738,N_13534);
and U16220 (N_16220,N_13323,N_12977);
and U16221 (N_16221,N_12491,N_12597);
nor U16222 (N_16222,N_12907,N_12471);
or U16223 (N_16223,N_12763,N_12309);
or U16224 (N_16224,N_14164,N_12581);
or U16225 (N_16225,N_12098,N_14126);
nor U16226 (N_16226,N_12950,N_13786);
nand U16227 (N_16227,N_13770,N_13677);
nor U16228 (N_16228,N_13040,N_14383);
nand U16229 (N_16229,N_14728,N_14171);
or U16230 (N_16230,N_13286,N_12621);
and U16231 (N_16231,N_12073,N_12301);
nand U16232 (N_16232,N_12067,N_14113);
or U16233 (N_16233,N_14787,N_13978);
nand U16234 (N_16234,N_14184,N_13678);
xnor U16235 (N_16235,N_14721,N_14050);
xnor U16236 (N_16236,N_14942,N_14039);
xnor U16237 (N_16237,N_13255,N_12097);
and U16238 (N_16238,N_12195,N_14444);
nand U16239 (N_16239,N_14386,N_14336);
nand U16240 (N_16240,N_14754,N_12824);
nand U16241 (N_16241,N_13229,N_14344);
and U16242 (N_16242,N_14167,N_12374);
nand U16243 (N_16243,N_13575,N_13922);
nor U16244 (N_16244,N_13606,N_12779);
nand U16245 (N_16245,N_14843,N_12699);
nor U16246 (N_16246,N_12716,N_12173);
nand U16247 (N_16247,N_13337,N_12387);
nor U16248 (N_16248,N_12544,N_12111);
and U16249 (N_16249,N_14112,N_13529);
nor U16250 (N_16250,N_12932,N_14573);
or U16251 (N_16251,N_14016,N_14325);
xor U16252 (N_16252,N_14494,N_12529);
xnor U16253 (N_16253,N_12520,N_12373);
nor U16254 (N_16254,N_14910,N_13658);
nor U16255 (N_16255,N_12185,N_14583);
and U16256 (N_16256,N_13028,N_13506);
xnor U16257 (N_16257,N_13218,N_13919);
nor U16258 (N_16258,N_12656,N_13913);
nor U16259 (N_16259,N_13355,N_14602);
nand U16260 (N_16260,N_12867,N_12160);
xnor U16261 (N_16261,N_13625,N_14044);
nand U16262 (N_16262,N_12629,N_12072);
nor U16263 (N_16263,N_14335,N_14516);
or U16264 (N_16264,N_13158,N_13297);
nor U16265 (N_16265,N_14119,N_14571);
or U16266 (N_16266,N_14518,N_13889);
and U16267 (N_16267,N_12745,N_13866);
and U16268 (N_16268,N_13880,N_13965);
or U16269 (N_16269,N_13608,N_14223);
nor U16270 (N_16270,N_13056,N_14331);
or U16271 (N_16271,N_12080,N_12019);
or U16272 (N_16272,N_14814,N_13474);
or U16273 (N_16273,N_14535,N_13690);
and U16274 (N_16274,N_14741,N_13781);
xnor U16275 (N_16275,N_14088,N_12310);
nand U16276 (N_16276,N_13225,N_14654);
or U16277 (N_16277,N_13148,N_13669);
nor U16278 (N_16278,N_13599,N_12578);
nand U16279 (N_16279,N_14918,N_13970);
and U16280 (N_16280,N_13924,N_14414);
nand U16281 (N_16281,N_12848,N_12860);
xnor U16282 (N_16282,N_14059,N_12945);
or U16283 (N_16283,N_14147,N_12834);
nand U16284 (N_16284,N_13888,N_14752);
and U16285 (N_16285,N_14724,N_13454);
nor U16286 (N_16286,N_12085,N_13820);
xor U16287 (N_16287,N_12139,N_13547);
nor U16288 (N_16288,N_14191,N_13779);
xor U16289 (N_16289,N_14095,N_14085);
xor U16290 (N_16290,N_12603,N_12341);
or U16291 (N_16291,N_12044,N_13621);
and U16292 (N_16292,N_14615,N_14210);
and U16293 (N_16293,N_13705,N_14076);
and U16294 (N_16294,N_14128,N_14810);
nor U16295 (N_16295,N_14468,N_12474);
nor U16296 (N_16296,N_13943,N_13991);
xnor U16297 (N_16297,N_13131,N_13383);
and U16298 (N_16298,N_12526,N_14280);
or U16299 (N_16299,N_14120,N_14798);
nor U16300 (N_16300,N_13886,N_13090);
nor U16301 (N_16301,N_13857,N_12232);
nor U16302 (N_16302,N_12172,N_12645);
xor U16303 (N_16303,N_12307,N_12692);
xnor U16304 (N_16304,N_14367,N_12818);
or U16305 (N_16305,N_14925,N_14154);
xnor U16306 (N_16306,N_13885,N_12170);
nor U16307 (N_16307,N_13664,N_12319);
or U16308 (N_16308,N_14288,N_14706);
xnor U16309 (N_16309,N_13179,N_13644);
nor U16310 (N_16310,N_13274,N_12640);
or U16311 (N_16311,N_12244,N_13224);
nor U16312 (N_16312,N_14669,N_14790);
nand U16313 (N_16313,N_14291,N_14750);
or U16314 (N_16314,N_12625,N_13840);
and U16315 (N_16315,N_13349,N_14985);
nor U16316 (N_16316,N_14452,N_14637);
xor U16317 (N_16317,N_12265,N_14915);
and U16318 (N_16318,N_12809,N_13636);
xnor U16319 (N_16319,N_13618,N_14197);
or U16320 (N_16320,N_13605,N_14459);
nor U16321 (N_16321,N_13817,N_13964);
nor U16322 (N_16322,N_14769,N_13750);
or U16323 (N_16323,N_12052,N_12688);
and U16324 (N_16324,N_13011,N_12343);
nand U16325 (N_16325,N_14656,N_14599);
nor U16326 (N_16326,N_14251,N_13634);
nand U16327 (N_16327,N_14012,N_12378);
or U16328 (N_16328,N_13398,N_12133);
nor U16329 (N_16329,N_12248,N_14190);
or U16330 (N_16330,N_12231,N_13416);
xor U16331 (N_16331,N_12259,N_13652);
nand U16332 (N_16332,N_12842,N_12312);
xor U16333 (N_16333,N_14964,N_13280);
and U16334 (N_16334,N_12015,N_14957);
and U16335 (N_16335,N_14357,N_14997);
and U16336 (N_16336,N_13296,N_13607);
nor U16337 (N_16337,N_12904,N_14924);
or U16338 (N_16338,N_13071,N_13807);
or U16339 (N_16339,N_14009,N_13438);
or U16340 (N_16340,N_14226,N_12857);
nand U16341 (N_16341,N_14874,N_13309);
nor U16342 (N_16342,N_12252,N_14045);
nor U16343 (N_16343,N_12066,N_13079);
nor U16344 (N_16344,N_14647,N_12033);
nor U16345 (N_16345,N_12510,N_13332);
xor U16346 (N_16346,N_13114,N_12525);
nand U16347 (N_16347,N_12004,N_13174);
or U16348 (N_16348,N_14590,N_13263);
or U16349 (N_16349,N_14033,N_14273);
or U16350 (N_16350,N_14099,N_13912);
and U16351 (N_16351,N_12998,N_12149);
and U16352 (N_16352,N_14252,N_13972);
nand U16353 (N_16353,N_14432,N_14838);
xor U16354 (N_16354,N_12592,N_12624);
and U16355 (N_16355,N_12696,N_13825);
and U16356 (N_16356,N_12527,N_14347);
xnor U16357 (N_16357,N_13246,N_13228);
nand U16358 (N_16358,N_13638,N_12417);
and U16359 (N_16359,N_14575,N_13971);
and U16360 (N_16360,N_13996,N_14708);
xnor U16361 (N_16361,N_12493,N_14249);
xnor U16362 (N_16362,N_14375,N_12190);
or U16363 (N_16363,N_12776,N_12881);
nor U16364 (N_16364,N_13760,N_13288);
and U16365 (N_16365,N_12135,N_14543);
nand U16366 (N_16366,N_13096,N_12087);
xor U16367 (N_16367,N_12550,N_12757);
xnor U16368 (N_16368,N_14567,N_14802);
nor U16369 (N_16369,N_14155,N_13749);
nor U16370 (N_16370,N_14253,N_12391);
or U16371 (N_16371,N_12730,N_14217);
nor U16372 (N_16372,N_12610,N_13837);
or U16373 (N_16373,N_14474,N_12118);
nand U16374 (N_16374,N_12032,N_13023);
or U16375 (N_16375,N_13696,N_12058);
and U16376 (N_16376,N_12068,N_12425);
or U16377 (N_16377,N_13740,N_14390);
nor U16378 (N_16378,N_14778,N_12762);
and U16379 (N_16379,N_12369,N_14424);
xor U16380 (N_16380,N_14220,N_12802);
nor U16381 (N_16381,N_13242,N_13493);
and U16382 (N_16382,N_13581,N_14075);
and U16383 (N_16383,N_14490,N_13173);
xnor U16384 (N_16384,N_12680,N_13680);
nand U16385 (N_16385,N_13736,N_14756);
or U16386 (N_16386,N_13329,N_14180);
nor U16387 (N_16387,N_14895,N_14620);
nand U16388 (N_16388,N_14714,N_14465);
and U16389 (N_16389,N_14264,N_12137);
xor U16390 (N_16390,N_13715,N_14279);
nor U16391 (N_16391,N_13829,N_13190);
nor U16392 (N_16392,N_12220,N_12508);
and U16393 (N_16393,N_12482,N_13053);
xor U16394 (N_16394,N_12180,N_14094);
or U16395 (N_16395,N_14986,N_14812);
or U16396 (N_16396,N_12877,N_14068);
xor U16397 (N_16397,N_13917,N_12515);
nor U16398 (N_16398,N_14116,N_14564);
nor U16399 (N_16399,N_12258,N_12524);
xor U16400 (N_16400,N_14676,N_14794);
nand U16401 (N_16401,N_12124,N_12476);
nand U16402 (N_16402,N_14289,N_12750);
nor U16403 (N_16403,N_13521,N_12174);
xor U16404 (N_16404,N_13414,N_13038);
or U16405 (N_16405,N_12513,N_12454);
nor U16406 (N_16406,N_12810,N_12345);
nor U16407 (N_16407,N_13109,N_14144);
nand U16408 (N_16408,N_13220,N_13672);
xnor U16409 (N_16409,N_13147,N_14699);
and U16410 (N_16410,N_14029,N_14152);
and U16411 (N_16411,N_12774,N_12546);
nand U16412 (N_16412,N_14346,N_14723);
nor U16413 (N_16413,N_12931,N_14234);
xnor U16414 (N_16414,N_12241,N_12559);
and U16415 (N_16415,N_12996,N_13527);
nand U16416 (N_16416,N_12188,N_14781);
nor U16417 (N_16417,N_14761,N_14780);
nor U16418 (N_16418,N_14342,N_12175);
xor U16419 (N_16419,N_12530,N_14604);
or U16420 (N_16420,N_13203,N_14385);
and U16421 (N_16421,N_12176,N_12866);
nand U16422 (N_16422,N_12984,N_12306);
nor U16423 (N_16423,N_13127,N_12075);
or U16424 (N_16424,N_13198,N_14678);
xnor U16425 (N_16425,N_12815,N_12014);
or U16426 (N_16426,N_14860,N_14332);
or U16427 (N_16427,N_12367,N_12187);
or U16428 (N_16428,N_14923,N_14809);
nand U16429 (N_16429,N_13139,N_13210);
and U16430 (N_16430,N_12217,N_14350);
or U16431 (N_16431,N_12246,N_13986);
nor U16432 (N_16432,N_14151,N_13401);
nor U16433 (N_16433,N_14379,N_12820);
nand U16434 (N_16434,N_14749,N_14764);
or U16435 (N_16435,N_12153,N_13085);
nand U16436 (N_16436,N_13126,N_14237);
nor U16437 (N_16437,N_14729,N_14100);
nor U16438 (N_16438,N_14744,N_14244);
nand U16439 (N_16439,N_14436,N_14854);
nand U16440 (N_16440,N_14278,N_13576);
nor U16441 (N_16441,N_12994,N_13087);
or U16442 (N_16442,N_13215,N_12235);
and U16443 (N_16443,N_12506,N_14423);
xnor U16444 (N_16444,N_13665,N_14140);
and U16445 (N_16445,N_13611,N_13212);
nor U16446 (N_16446,N_14064,N_12575);
nand U16447 (N_16447,N_13953,N_12979);
and U16448 (N_16448,N_14513,N_13469);
xor U16449 (N_16449,N_12552,N_13879);
or U16450 (N_16450,N_12012,N_13067);
nand U16451 (N_16451,N_14233,N_13516);
xor U16452 (N_16452,N_13990,N_12043);
and U16453 (N_16453,N_14141,N_12888);
xor U16454 (N_16454,N_12126,N_13743);
nor U16455 (N_16455,N_14917,N_13209);
nand U16456 (N_16456,N_13930,N_12752);
nand U16457 (N_16457,N_13789,N_12273);
and U16458 (N_16458,N_12753,N_12362);
nor U16459 (N_16459,N_14956,N_14962);
or U16460 (N_16460,N_12084,N_13254);
or U16461 (N_16461,N_12825,N_12554);
and U16462 (N_16462,N_13252,N_13159);
and U16463 (N_16463,N_14256,N_12426);
nor U16464 (N_16464,N_14020,N_12331);
xor U16465 (N_16465,N_14578,N_14146);
nor U16466 (N_16466,N_12711,N_12823);
and U16467 (N_16467,N_14018,N_14006);
nand U16468 (N_16468,N_13000,N_13216);
and U16469 (N_16469,N_14595,N_14718);
nand U16470 (N_16470,N_14666,N_12519);
nand U16471 (N_16471,N_13640,N_12413);
nand U16472 (N_16472,N_14122,N_13950);
and U16473 (N_16473,N_12239,N_13784);
or U16474 (N_16474,N_13485,N_14071);
nand U16475 (N_16475,N_13596,N_14680);
xor U16476 (N_16476,N_13704,N_12264);
or U16477 (N_16477,N_14624,N_13445);
or U16478 (N_16478,N_14483,N_12370);
xor U16479 (N_16479,N_14639,N_14887);
or U16480 (N_16480,N_14157,N_12386);
and U16481 (N_16481,N_14097,N_14725);
or U16482 (N_16482,N_13742,N_12480);
nor U16483 (N_16483,N_13849,N_12674);
nor U16484 (N_16484,N_12256,N_14550);
nor U16485 (N_16485,N_14495,N_13628);
or U16486 (N_16486,N_14707,N_13222);
nor U16487 (N_16487,N_14553,N_13045);
and U16488 (N_16488,N_13472,N_13265);
nand U16489 (N_16489,N_13467,N_13778);
nand U16490 (N_16490,N_14514,N_14510);
nor U16491 (N_16491,N_13046,N_12790);
nand U16492 (N_16492,N_13374,N_12851);
xor U16493 (N_16493,N_14453,N_14415);
nor U16494 (N_16494,N_14216,N_13219);
and U16495 (N_16495,N_12507,N_14194);
nand U16496 (N_16496,N_12178,N_12829);
or U16497 (N_16497,N_12858,N_12577);
xnor U16498 (N_16498,N_13519,N_12079);
xor U16499 (N_16499,N_12348,N_13318);
nand U16500 (N_16500,N_14623,N_14377);
and U16501 (N_16501,N_12859,N_13614);
nor U16502 (N_16502,N_13969,N_14954);
or U16503 (N_16503,N_13837,N_12589);
nand U16504 (N_16504,N_12373,N_14300);
xnor U16505 (N_16505,N_12409,N_12374);
nand U16506 (N_16506,N_13714,N_13471);
or U16507 (N_16507,N_14488,N_14235);
or U16508 (N_16508,N_12906,N_12786);
and U16509 (N_16509,N_13995,N_13066);
nand U16510 (N_16510,N_13882,N_12604);
xnor U16511 (N_16511,N_13720,N_13826);
nand U16512 (N_16512,N_12267,N_13248);
nor U16513 (N_16513,N_12011,N_13812);
and U16514 (N_16514,N_13020,N_12017);
xor U16515 (N_16515,N_14915,N_12404);
and U16516 (N_16516,N_13825,N_13815);
nor U16517 (N_16517,N_13961,N_13234);
nand U16518 (N_16518,N_12415,N_13527);
and U16519 (N_16519,N_12709,N_13904);
xor U16520 (N_16520,N_13393,N_12149);
and U16521 (N_16521,N_14930,N_13775);
nor U16522 (N_16522,N_14329,N_13758);
xnor U16523 (N_16523,N_13633,N_13329);
nor U16524 (N_16524,N_12662,N_14629);
nand U16525 (N_16525,N_14836,N_14299);
nand U16526 (N_16526,N_13277,N_14262);
nor U16527 (N_16527,N_13325,N_12142);
and U16528 (N_16528,N_12336,N_13155);
or U16529 (N_16529,N_14821,N_12572);
xor U16530 (N_16530,N_14813,N_14882);
nor U16531 (N_16531,N_12037,N_14696);
nor U16532 (N_16532,N_13493,N_14664);
and U16533 (N_16533,N_12288,N_13221);
or U16534 (N_16534,N_13823,N_13681);
nor U16535 (N_16535,N_13021,N_14738);
nand U16536 (N_16536,N_13354,N_14987);
nor U16537 (N_16537,N_13542,N_14544);
and U16538 (N_16538,N_14198,N_14000);
nand U16539 (N_16539,N_14160,N_13840);
nor U16540 (N_16540,N_13392,N_12797);
or U16541 (N_16541,N_14873,N_14463);
and U16542 (N_16542,N_14313,N_13904);
or U16543 (N_16543,N_12307,N_13893);
xor U16544 (N_16544,N_12936,N_12144);
and U16545 (N_16545,N_14404,N_14472);
or U16546 (N_16546,N_14606,N_12183);
and U16547 (N_16547,N_14246,N_14988);
nand U16548 (N_16548,N_14830,N_14642);
nand U16549 (N_16549,N_13148,N_12212);
nor U16550 (N_16550,N_14571,N_14848);
and U16551 (N_16551,N_13143,N_12652);
and U16552 (N_16552,N_14737,N_12980);
or U16553 (N_16553,N_14379,N_13970);
and U16554 (N_16554,N_12802,N_12724);
nor U16555 (N_16555,N_14949,N_14068);
nor U16556 (N_16556,N_13923,N_13641);
nor U16557 (N_16557,N_13355,N_12468);
or U16558 (N_16558,N_12779,N_12928);
and U16559 (N_16559,N_12348,N_12063);
nand U16560 (N_16560,N_12977,N_14718);
nor U16561 (N_16561,N_14013,N_14905);
nor U16562 (N_16562,N_13215,N_13235);
xor U16563 (N_16563,N_12412,N_12993);
xor U16564 (N_16564,N_13732,N_13269);
and U16565 (N_16565,N_14189,N_14316);
nor U16566 (N_16566,N_12836,N_12145);
or U16567 (N_16567,N_12850,N_14831);
and U16568 (N_16568,N_12400,N_14954);
nand U16569 (N_16569,N_12421,N_13201);
xnor U16570 (N_16570,N_13029,N_13329);
or U16571 (N_16571,N_14106,N_14012);
or U16572 (N_16572,N_14289,N_13683);
xnor U16573 (N_16573,N_14386,N_14562);
or U16574 (N_16574,N_12708,N_12623);
xor U16575 (N_16575,N_14916,N_13918);
nor U16576 (N_16576,N_13171,N_13076);
nand U16577 (N_16577,N_14020,N_14540);
nand U16578 (N_16578,N_12319,N_14999);
nor U16579 (N_16579,N_13539,N_12962);
or U16580 (N_16580,N_14335,N_14178);
nor U16581 (N_16581,N_14037,N_13699);
or U16582 (N_16582,N_12919,N_12932);
and U16583 (N_16583,N_12156,N_12665);
nand U16584 (N_16584,N_13041,N_13782);
xor U16585 (N_16585,N_12581,N_14399);
nand U16586 (N_16586,N_13290,N_12956);
nand U16587 (N_16587,N_13080,N_14241);
nand U16588 (N_16588,N_13729,N_13748);
and U16589 (N_16589,N_12728,N_13684);
and U16590 (N_16590,N_12025,N_13155);
xnor U16591 (N_16591,N_14412,N_13538);
nor U16592 (N_16592,N_13749,N_13665);
and U16593 (N_16593,N_12043,N_12688);
xor U16594 (N_16594,N_13726,N_13235);
or U16595 (N_16595,N_14645,N_13248);
nor U16596 (N_16596,N_12011,N_14217);
xnor U16597 (N_16597,N_14047,N_13262);
nor U16598 (N_16598,N_12013,N_12893);
nor U16599 (N_16599,N_12321,N_12124);
nand U16600 (N_16600,N_14603,N_12646);
and U16601 (N_16601,N_14031,N_13783);
xor U16602 (N_16602,N_12646,N_12924);
nor U16603 (N_16603,N_14415,N_13404);
nand U16604 (N_16604,N_12041,N_14822);
xor U16605 (N_16605,N_14167,N_14028);
or U16606 (N_16606,N_14500,N_14999);
nand U16607 (N_16607,N_13331,N_13557);
nand U16608 (N_16608,N_14196,N_13396);
and U16609 (N_16609,N_13701,N_14645);
xnor U16610 (N_16610,N_14703,N_12133);
nor U16611 (N_16611,N_14469,N_13480);
or U16612 (N_16612,N_13572,N_14083);
nor U16613 (N_16613,N_12031,N_13718);
or U16614 (N_16614,N_12982,N_14773);
and U16615 (N_16615,N_14057,N_14473);
or U16616 (N_16616,N_13182,N_13448);
xor U16617 (N_16617,N_13847,N_12145);
or U16618 (N_16618,N_14704,N_14263);
nand U16619 (N_16619,N_13813,N_13141);
or U16620 (N_16620,N_13095,N_14844);
xor U16621 (N_16621,N_12028,N_13629);
xnor U16622 (N_16622,N_13144,N_13830);
or U16623 (N_16623,N_12290,N_14254);
and U16624 (N_16624,N_12265,N_14327);
nand U16625 (N_16625,N_14809,N_12974);
or U16626 (N_16626,N_13641,N_14592);
nand U16627 (N_16627,N_14389,N_14459);
nor U16628 (N_16628,N_12125,N_14281);
nand U16629 (N_16629,N_13968,N_13209);
and U16630 (N_16630,N_13565,N_13113);
xor U16631 (N_16631,N_12526,N_12426);
xor U16632 (N_16632,N_13714,N_14582);
nor U16633 (N_16633,N_14483,N_14744);
and U16634 (N_16634,N_12909,N_14328);
and U16635 (N_16635,N_12442,N_13802);
or U16636 (N_16636,N_14631,N_13658);
nand U16637 (N_16637,N_14449,N_12976);
xor U16638 (N_16638,N_12165,N_12001);
and U16639 (N_16639,N_13116,N_13198);
xnor U16640 (N_16640,N_12937,N_13762);
nor U16641 (N_16641,N_13419,N_13782);
and U16642 (N_16642,N_13758,N_12216);
xor U16643 (N_16643,N_13693,N_13018);
or U16644 (N_16644,N_12389,N_12647);
or U16645 (N_16645,N_14079,N_13790);
xnor U16646 (N_16646,N_12089,N_14462);
xnor U16647 (N_16647,N_12889,N_12411);
and U16648 (N_16648,N_13541,N_13740);
nor U16649 (N_16649,N_12029,N_14004);
or U16650 (N_16650,N_12658,N_12219);
xor U16651 (N_16651,N_14610,N_12296);
xor U16652 (N_16652,N_13618,N_12103);
and U16653 (N_16653,N_12119,N_13062);
or U16654 (N_16654,N_13051,N_13010);
and U16655 (N_16655,N_12615,N_13785);
and U16656 (N_16656,N_12699,N_14810);
or U16657 (N_16657,N_14337,N_12295);
and U16658 (N_16658,N_12423,N_13168);
nor U16659 (N_16659,N_14598,N_14080);
nor U16660 (N_16660,N_13910,N_12340);
nand U16661 (N_16661,N_13022,N_12657);
nor U16662 (N_16662,N_12477,N_14973);
or U16663 (N_16663,N_14495,N_14524);
xnor U16664 (N_16664,N_12149,N_14375);
xor U16665 (N_16665,N_14123,N_12673);
nand U16666 (N_16666,N_12424,N_12989);
nor U16667 (N_16667,N_13284,N_12414);
and U16668 (N_16668,N_13104,N_12424);
nor U16669 (N_16669,N_14202,N_12958);
and U16670 (N_16670,N_12626,N_12320);
nand U16671 (N_16671,N_13420,N_14738);
and U16672 (N_16672,N_14770,N_12516);
nor U16673 (N_16673,N_12976,N_12746);
xnor U16674 (N_16674,N_13044,N_14305);
xnor U16675 (N_16675,N_14379,N_13950);
or U16676 (N_16676,N_13864,N_14071);
or U16677 (N_16677,N_13570,N_12043);
nor U16678 (N_16678,N_14775,N_12412);
or U16679 (N_16679,N_13636,N_12328);
or U16680 (N_16680,N_12132,N_12031);
and U16681 (N_16681,N_12397,N_12358);
nand U16682 (N_16682,N_12180,N_12768);
or U16683 (N_16683,N_14927,N_13941);
or U16684 (N_16684,N_12262,N_13690);
xor U16685 (N_16685,N_13174,N_13959);
xor U16686 (N_16686,N_14094,N_14888);
xnor U16687 (N_16687,N_14675,N_14269);
nor U16688 (N_16688,N_12523,N_13977);
xnor U16689 (N_16689,N_14376,N_14255);
nor U16690 (N_16690,N_14235,N_12329);
and U16691 (N_16691,N_13911,N_12269);
xor U16692 (N_16692,N_13219,N_14023);
nor U16693 (N_16693,N_13728,N_14695);
and U16694 (N_16694,N_14172,N_14645);
or U16695 (N_16695,N_12975,N_12215);
nand U16696 (N_16696,N_12860,N_13978);
nand U16697 (N_16697,N_14077,N_12827);
and U16698 (N_16698,N_13416,N_13420);
xnor U16699 (N_16699,N_14190,N_14383);
nand U16700 (N_16700,N_14898,N_13392);
nand U16701 (N_16701,N_14853,N_13274);
nand U16702 (N_16702,N_14354,N_13575);
xnor U16703 (N_16703,N_13175,N_14012);
and U16704 (N_16704,N_12951,N_13070);
nor U16705 (N_16705,N_12946,N_12613);
xor U16706 (N_16706,N_12367,N_13858);
or U16707 (N_16707,N_13806,N_14223);
nand U16708 (N_16708,N_12423,N_13641);
and U16709 (N_16709,N_12052,N_12967);
and U16710 (N_16710,N_12652,N_12157);
nor U16711 (N_16711,N_14800,N_14802);
nand U16712 (N_16712,N_13976,N_13907);
and U16713 (N_16713,N_12466,N_13362);
xnor U16714 (N_16714,N_13855,N_12033);
and U16715 (N_16715,N_13732,N_12742);
nand U16716 (N_16716,N_13144,N_12988);
xor U16717 (N_16717,N_12766,N_12145);
nand U16718 (N_16718,N_13911,N_14312);
or U16719 (N_16719,N_14716,N_13167);
xor U16720 (N_16720,N_12498,N_14600);
nor U16721 (N_16721,N_13526,N_14172);
or U16722 (N_16722,N_14921,N_12703);
and U16723 (N_16723,N_12200,N_14911);
nand U16724 (N_16724,N_13539,N_12913);
and U16725 (N_16725,N_13114,N_14391);
xor U16726 (N_16726,N_13827,N_12099);
and U16727 (N_16727,N_13909,N_14016);
or U16728 (N_16728,N_13384,N_14697);
nor U16729 (N_16729,N_12909,N_13001);
or U16730 (N_16730,N_13557,N_14628);
and U16731 (N_16731,N_14446,N_12790);
or U16732 (N_16732,N_12407,N_13958);
or U16733 (N_16733,N_12304,N_14527);
xor U16734 (N_16734,N_14893,N_12919);
nand U16735 (N_16735,N_12235,N_12679);
nor U16736 (N_16736,N_13586,N_14441);
and U16737 (N_16737,N_13662,N_13404);
nand U16738 (N_16738,N_12519,N_13790);
nor U16739 (N_16739,N_12705,N_13371);
xor U16740 (N_16740,N_12380,N_13487);
nor U16741 (N_16741,N_12423,N_13487);
nor U16742 (N_16742,N_14529,N_12581);
and U16743 (N_16743,N_12419,N_12218);
nand U16744 (N_16744,N_13542,N_14139);
or U16745 (N_16745,N_13891,N_14932);
or U16746 (N_16746,N_13520,N_12673);
nor U16747 (N_16747,N_12801,N_13531);
nand U16748 (N_16748,N_12206,N_14986);
nand U16749 (N_16749,N_14490,N_12244);
nor U16750 (N_16750,N_13290,N_13925);
xor U16751 (N_16751,N_14691,N_14126);
nand U16752 (N_16752,N_14625,N_13461);
nor U16753 (N_16753,N_14501,N_12136);
or U16754 (N_16754,N_13527,N_13348);
or U16755 (N_16755,N_14612,N_14290);
nor U16756 (N_16756,N_14593,N_12486);
xnor U16757 (N_16757,N_14004,N_14610);
xnor U16758 (N_16758,N_12738,N_13237);
xor U16759 (N_16759,N_12570,N_12675);
and U16760 (N_16760,N_13427,N_12416);
or U16761 (N_16761,N_13602,N_13601);
or U16762 (N_16762,N_14791,N_13722);
nand U16763 (N_16763,N_12980,N_14896);
xnor U16764 (N_16764,N_14420,N_13532);
xor U16765 (N_16765,N_13944,N_12838);
xnor U16766 (N_16766,N_12908,N_12245);
or U16767 (N_16767,N_14731,N_14358);
nand U16768 (N_16768,N_12138,N_12859);
xor U16769 (N_16769,N_13114,N_13623);
nand U16770 (N_16770,N_14587,N_14224);
nand U16771 (N_16771,N_13120,N_13639);
and U16772 (N_16772,N_14311,N_12187);
or U16773 (N_16773,N_13884,N_12292);
xor U16774 (N_16774,N_12780,N_14135);
xor U16775 (N_16775,N_14267,N_14917);
xor U16776 (N_16776,N_13203,N_14656);
or U16777 (N_16777,N_12219,N_13032);
xor U16778 (N_16778,N_12511,N_12730);
or U16779 (N_16779,N_12452,N_14153);
nor U16780 (N_16780,N_14107,N_12248);
and U16781 (N_16781,N_12856,N_12187);
nand U16782 (N_16782,N_13036,N_14740);
or U16783 (N_16783,N_14422,N_12158);
or U16784 (N_16784,N_14814,N_12898);
or U16785 (N_16785,N_13559,N_12116);
and U16786 (N_16786,N_12642,N_14969);
or U16787 (N_16787,N_13654,N_14365);
nor U16788 (N_16788,N_14915,N_12840);
nor U16789 (N_16789,N_13737,N_12025);
or U16790 (N_16790,N_14404,N_14351);
nor U16791 (N_16791,N_14320,N_12294);
and U16792 (N_16792,N_13297,N_12800);
or U16793 (N_16793,N_12739,N_14919);
and U16794 (N_16794,N_12132,N_12921);
nor U16795 (N_16795,N_12361,N_14262);
nand U16796 (N_16796,N_13596,N_13965);
or U16797 (N_16797,N_13594,N_14174);
nor U16798 (N_16798,N_13974,N_13720);
nor U16799 (N_16799,N_14099,N_12768);
and U16800 (N_16800,N_12865,N_14633);
or U16801 (N_16801,N_12726,N_13515);
and U16802 (N_16802,N_12830,N_13437);
xor U16803 (N_16803,N_12451,N_12119);
nand U16804 (N_16804,N_13567,N_13470);
xor U16805 (N_16805,N_12127,N_12407);
xnor U16806 (N_16806,N_12895,N_13176);
or U16807 (N_16807,N_14448,N_13402);
nand U16808 (N_16808,N_13215,N_14495);
xor U16809 (N_16809,N_13456,N_13064);
xor U16810 (N_16810,N_14035,N_12557);
nand U16811 (N_16811,N_12609,N_13413);
xor U16812 (N_16812,N_12358,N_13233);
or U16813 (N_16813,N_12470,N_13957);
nand U16814 (N_16814,N_14739,N_14713);
and U16815 (N_16815,N_12080,N_12030);
nor U16816 (N_16816,N_13746,N_12172);
or U16817 (N_16817,N_12399,N_13338);
nor U16818 (N_16818,N_12367,N_13124);
nor U16819 (N_16819,N_13693,N_14698);
and U16820 (N_16820,N_14138,N_12978);
xnor U16821 (N_16821,N_13841,N_13666);
nand U16822 (N_16822,N_14267,N_13155);
and U16823 (N_16823,N_12097,N_12128);
and U16824 (N_16824,N_13570,N_12023);
and U16825 (N_16825,N_13735,N_12035);
xor U16826 (N_16826,N_14797,N_14466);
nor U16827 (N_16827,N_14591,N_13166);
nand U16828 (N_16828,N_12477,N_14907);
and U16829 (N_16829,N_12612,N_13223);
or U16830 (N_16830,N_14792,N_13711);
or U16831 (N_16831,N_14237,N_12262);
and U16832 (N_16832,N_14430,N_12342);
or U16833 (N_16833,N_13388,N_13009);
xnor U16834 (N_16834,N_12067,N_14342);
nor U16835 (N_16835,N_13714,N_13844);
nand U16836 (N_16836,N_12759,N_13974);
and U16837 (N_16837,N_14105,N_12978);
nor U16838 (N_16838,N_12505,N_13747);
nand U16839 (N_16839,N_14835,N_12467);
nor U16840 (N_16840,N_13314,N_14307);
or U16841 (N_16841,N_13227,N_14821);
xnor U16842 (N_16842,N_14855,N_12637);
xnor U16843 (N_16843,N_12282,N_12160);
and U16844 (N_16844,N_12440,N_13807);
xor U16845 (N_16845,N_12666,N_14309);
and U16846 (N_16846,N_14255,N_12523);
and U16847 (N_16847,N_13892,N_12348);
xnor U16848 (N_16848,N_14137,N_13630);
and U16849 (N_16849,N_13928,N_14248);
xnor U16850 (N_16850,N_13192,N_12786);
xor U16851 (N_16851,N_13825,N_14130);
or U16852 (N_16852,N_14643,N_12392);
and U16853 (N_16853,N_13603,N_12444);
or U16854 (N_16854,N_12497,N_12361);
or U16855 (N_16855,N_14492,N_14442);
nand U16856 (N_16856,N_13281,N_14734);
nand U16857 (N_16857,N_12187,N_12759);
xor U16858 (N_16858,N_12294,N_14293);
xnor U16859 (N_16859,N_14552,N_13703);
nand U16860 (N_16860,N_14937,N_13637);
or U16861 (N_16861,N_12669,N_14349);
nand U16862 (N_16862,N_14475,N_12281);
xnor U16863 (N_16863,N_12090,N_12622);
and U16864 (N_16864,N_13661,N_14444);
and U16865 (N_16865,N_12631,N_12380);
xnor U16866 (N_16866,N_14306,N_13805);
nor U16867 (N_16867,N_14452,N_14409);
nor U16868 (N_16868,N_14683,N_14844);
or U16869 (N_16869,N_12374,N_12585);
xor U16870 (N_16870,N_13582,N_12830);
nor U16871 (N_16871,N_12931,N_12175);
xnor U16872 (N_16872,N_12882,N_12275);
xor U16873 (N_16873,N_14776,N_12902);
xnor U16874 (N_16874,N_14351,N_14666);
nor U16875 (N_16875,N_13920,N_13700);
nor U16876 (N_16876,N_13490,N_14185);
nor U16877 (N_16877,N_12502,N_12436);
and U16878 (N_16878,N_12710,N_14378);
or U16879 (N_16879,N_14022,N_12457);
nor U16880 (N_16880,N_14433,N_13719);
xor U16881 (N_16881,N_12796,N_12956);
nor U16882 (N_16882,N_14385,N_12348);
and U16883 (N_16883,N_13531,N_14630);
nand U16884 (N_16884,N_14278,N_13010);
xnor U16885 (N_16885,N_13271,N_14953);
xnor U16886 (N_16886,N_14981,N_14398);
xor U16887 (N_16887,N_12267,N_13337);
nor U16888 (N_16888,N_13107,N_13328);
or U16889 (N_16889,N_13926,N_12501);
xnor U16890 (N_16890,N_14219,N_13498);
or U16891 (N_16891,N_12868,N_14116);
nor U16892 (N_16892,N_14795,N_14154);
or U16893 (N_16893,N_12441,N_12007);
xnor U16894 (N_16894,N_13406,N_12777);
xnor U16895 (N_16895,N_13273,N_12421);
and U16896 (N_16896,N_13238,N_14349);
and U16897 (N_16897,N_12439,N_13198);
nor U16898 (N_16898,N_12216,N_12245);
or U16899 (N_16899,N_14426,N_12156);
nor U16900 (N_16900,N_14094,N_14624);
nor U16901 (N_16901,N_14038,N_12102);
nand U16902 (N_16902,N_12150,N_14785);
nor U16903 (N_16903,N_14661,N_14054);
nand U16904 (N_16904,N_13110,N_12575);
nand U16905 (N_16905,N_14736,N_13070);
xor U16906 (N_16906,N_12466,N_14643);
or U16907 (N_16907,N_12628,N_14841);
nand U16908 (N_16908,N_12817,N_13169);
or U16909 (N_16909,N_13695,N_12775);
nor U16910 (N_16910,N_13855,N_14571);
nor U16911 (N_16911,N_12119,N_14585);
nor U16912 (N_16912,N_14747,N_12721);
or U16913 (N_16913,N_13487,N_14525);
or U16914 (N_16914,N_14104,N_13756);
nor U16915 (N_16915,N_14239,N_13378);
nand U16916 (N_16916,N_12679,N_14678);
or U16917 (N_16917,N_14328,N_14244);
or U16918 (N_16918,N_14493,N_12226);
nand U16919 (N_16919,N_14094,N_14249);
or U16920 (N_16920,N_12069,N_14220);
xnor U16921 (N_16921,N_12760,N_13923);
and U16922 (N_16922,N_12660,N_12796);
and U16923 (N_16923,N_13504,N_12660);
or U16924 (N_16924,N_12863,N_14558);
nor U16925 (N_16925,N_14936,N_14023);
xnor U16926 (N_16926,N_13113,N_14897);
nand U16927 (N_16927,N_14097,N_14711);
nand U16928 (N_16928,N_14632,N_13181);
xor U16929 (N_16929,N_12837,N_12465);
or U16930 (N_16930,N_14357,N_12549);
xnor U16931 (N_16931,N_13928,N_14014);
xor U16932 (N_16932,N_13822,N_12811);
nor U16933 (N_16933,N_12890,N_12766);
nor U16934 (N_16934,N_14328,N_13950);
and U16935 (N_16935,N_13925,N_14198);
nand U16936 (N_16936,N_13599,N_13121);
nor U16937 (N_16937,N_12460,N_12731);
nand U16938 (N_16938,N_14319,N_14754);
nand U16939 (N_16939,N_14705,N_12128);
nand U16940 (N_16940,N_14985,N_13728);
xor U16941 (N_16941,N_14631,N_12687);
nand U16942 (N_16942,N_14362,N_13576);
or U16943 (N_16943,N_14298,N_13332);
and U16944 (N_16944,N_14157,N_13825);
or U16945 (N_16945,N_13573,N_13397);
xnor U16946 (N_16946,N_12345,N_14998);
nand U16947 (N_16947,N_14871,N_13147);
or U16948 (N_16948,N_14606,N_13834);
nor U16949 (N_16949,N_13410,N_14719);
and U16950 (N_16950,N_13721,N_14852);
nor U16951 (N_16951,N_12718,N_13913);
or U16952 (N_16952,N_14957,N_12094);
nand U16953 (N_16953,N_12527,N_12017);
nor U16954 (N_16954,N_12470,N_12762);
nand U16955 (N_16955,N_13820,N_12125);
nor U16956 (N_16956,N_14089,N_13059);
nor U16957 (N_16957,N_12776,N_12337);
nor U16958 (N_16958,N_13794,N_14599);
or U16959 (N_16959,N_13616,N_14744);
nor U16960 (N_16960,N_13105,N_14547);
or U16961 (N_16961,N_14205,N_12341);
nand U16962 (N_16962,N_14092,N_14837);
or U16963 (N_16963,N_13902,N_14006);
and U16964 (N_16964,N_14352,N_14095);
nor U16965 (N_16965,N_14427,N_13764);
nand U16966 (N_16966,N_13756,N_13224);
xnor U16967 (N_16967,N_14585,N_14694);
xnor U16968 (N_16968,N_14182,N_14554);
or U16969 (N_16969,N_14640,N_13324);
or U16970 (N_16970,N_13390,N_13451);
nor U16971 (N_16971,N_14184,N_14886);
nor U16972 (N_16972,N_13332,N_13136);
or U16973 (N_16973,N_14403,N_12913);
or U16974 (N_16974,N_13134,N_13763);
and U16975 (N_16975,N_12206,N_13335);
and U16976 (N_16976,N_13958,N_14431);
xnor U16977 (N_16977,N_13957,N_13702);
or U16978 (N_16978,N_13328,N_14598);
nor U16979 (N_16979,N_14884,N_13737);
nand U16980 (N_16980,N_13455,N_14531);
nand U16981 (N_16981,N_13002,N_12882);
or U16982 (N_16982,N_13196,N_12007);
nor U16983 (N_16983,N_14527,N_13324);
nor U16984 (N_16984,N_12865,N_14738);
or U16985 (N_16985,N_14610,N_14863);
nand U16986 (N_16986,N_12330,N_12307);
or U16987 (N_16987,N_14933,N_13328);
or U16988 (N_16988,N_13223,N_14221);
or U16989 (N_16989,N_14140,N_12710);
or U16990 (N_16990,N_13049,N_14932);
nor U16991 (N_16991,N_12598,N_14789);
nand U16992 (N_16992,N_12110,N_14781);
nor U16993 (N_16993,N_13019,N_14212);
and U16994 (N_16994,N_13693,N_14090);
or U16995 (N_16995,N_13025,N_13496);
xor U16996 (N_16996,N_12013,N_12553);
nand U16997 (N_16997,N_14997,N_13958);
nand U16998 (N_16998,N_13724,N_14746);
or U16999 (N_16999,N_14587,N_12715);
nand U17000 (N_17000,N_12271,N_13688);
or U17001 (N_17001,N_14786,N_14288);
nand U17002 (N_17002,N_13302,N_14038);
and U17003 (N_17003,N_13347,N_14416);
xor U17004 (N_17004,N_14942,N_14915);
and U17005 (N_17005,N_14895,N_14315);
nand U17006 (N_17006,N_12161,N_12016);
nor U17007 (N_17007,N_13097,N_12074);
or U17008 (N_17008,N_12657,N_12240);
xnor U17009 (N_17009,N_13580,N_14344);
nand U17010 (N_17010,N_12105,N_12583);
nor U17011 (N_17011,N_13981,N_13775);
nor U17012 (N_17012,N_13996,N_13363);
and U17013 (N_17013,N_13841,N_14084);
and U17014 (N_17014,N_12051,N_14480);
or U17015 (N_17015,N_12859,N_13791);
and U17016 (N_17016,N_14849,N_13525);
and U17017 (N_17017,N_12555,N_13970);
and U17018 (N_17018,N_14908,N_13705);
and U17019 (N_17019,N_12955,N_13942);
nor U17020 (N_17020,N_14381,N_12663);
or U17021 (N_17021,N_13098,N_14828);
xnor U17022 (N_17022,N_14424,N_13391);
nor U17023 (N_17023,N_12944,N_12732);
nor U17024 (N_17024,N_14093,N_14589);
xor U17025 (N_17025,N_14635,N_14686);
xnor U17026 (N_17026,N_12179,N_13327);
and U17027 (N_17027,N_14257,N_14873);
nand U17028 (N_17028,N_12077,N_13688);
xor U17029 (N_17029,N_12785,N_13235);
xnor U17030 (N_17030,N_12715,N_12217);
nor U17031 (N_17031,N_12794,N_14532);
or U17032 (N_17032,N_14642,N_12906);
nor U17033 (N_17033,N_12704,N_14478);
xor U17034 (N_17034,N_13500,N_13919);
and U17035 (N_17035,N_14942,N_14415);
nand U17036 (N_17036,N_13851,N_12159);
or U17037 (N_17037,N_12116,N_14979);
nor U17038 (N_17038,N_13582,N_12359);
nor U17039 (N_17039,N_12274,N_12204);
and U17040 (N_17040,N_14601,N_14566);
or U17041 (N_17041,N_14508,N_13422);
or U17042 (N_17042,N_12013,N_12403);
xor U17043 (N_17043,N_13487,N_13323);
or U17044 (N_17044,N_14797,N_12261);
xor U17045 (N_17045,N_13412,N_14077);
nor U17046 (N_17046,N_14350,N_13935);
and U17047 (N_17047,N_14741,N_13255);
and U17048 (N_17048,N_14231,N_13461);
nand U17049 (N_17049,N_13524,N_14884);
and U17050 (N_17050,N_12060,N_13824);
or U17051 (N_17051,N_13054,N_12790);
and U17052 (N_17052,N_14582,N_14153);
xor U17053 (N_17053,N_12915,N_13425);
xor U17054 (N_17054,N_12774,N_14898);
xor U17055 (N_17055,N_14636,N_12712);
or U17056 (N_17056,N_12191,N_14093);
nor U17057 (N_17057,N_13503,N_14263);
and U17058 (N_17058,N_12742,N_14810);
nor U17059 (N_17059,N_12371,N_13782);
nor U17060 (N_17060,N_12304,N_12490);
nor U17061 (N_17061,N_12042,N_13091);
xnor U17062 (N_17062,N_13109,N_13695);
nand U17063 (N_17063,N_13542,N_13653);
xnor U17064 (N_17064,N_14864,N_12859);
xnor U17065 (N_17065,N_14102,N_14027);
nor U17066 (N_17066,N_13459,N_12305);
xor U17067 (N_17067,N_14013,N_13358);
and U17068 (N_17068,N_14586,N_13267);
xor U17069 (N_17069,N_13704,N_12152);
xor U17070 (N_17070,N_13791,N_13179);
or U17071 (N_17071,N_12483,N_13270);
and U17072 (N_17072,N_13560,N_13971);
nor U17073 (N_17073,N_12499,N_13141);
nor U17074 (N_17074,N_13884,N_12522);
or U17075 (N_17075,N_14576,N_12242);
or U17076 (N_17076,N_14083,N_12503);
and U17077 (N_17077,N_13397,N_12979);
xnor U17078 (N_17078,N_14885,N_12247);
nor U17079 (N_17079,N_13794,N_12795);
nand U17080 (N_17080,N_12014,N_13940);
and U17081 (N_17081,N_13920,N_13433);
xnor U17082 (N_17082,N_13756,N_13458);
and U17083 (N_17083,N_12039,N_14494);
or U17084 (N_17084,N_13778,N_12559);
xnor U17085 (N_17085,N_14776,N_13826);
nand U17086 (N_17086,N_12234,N_14702);
nand U17087 (N_17087,N_12623,N_14584);
xnor U17088 (N_17088,N_13414,N_14966);
or U17089 (N_17089,N_12733,N_12652);
and U17090 (N_17090,N_12708,N_13862);
nor U17091 (N_17091,N_14271,N_14749);
and U17092 (N_17092,N_12881,N_13714);
xnor U17093 (N_17093,N_14543,N_13789);
nor U17094 (N_17094,N_14422,N_12024);
nor U17095 (N_17095,N_14033,N_13087);
nor U17096 (N_17096,N_12600,N_13031);
nor U17097 (N_17097,N_12332,N_13292);
and U17098 (N_17098,N_12161,N_13718);
and U17099 (N_17099,N_13434,N_12580);
and U17100 (N_17100,N_12708,N_12371);
or U17101 (N_17101,N_14726,N_14763);
or U17102 (N_17102,N_12590,N_14650);
nor U17103 (N_17103,N_13248,N_14493);
xnor U17104 (N_17104,N_13868,N_13454);
nand U17105 (N_17105,N_12394,N_13680);
xor U17106 (N_17106,N_12064,N_12747);
nand U17107 (N_17107,N_14992,N_12527);
and U17108 (N_17108,N_14889,N_13791);
and U17109 (N_17109,N_13377,N_13240);
and U17110 (N_17110,N_14399,N_13680);
xnor U17111 (N_17111,N_12058,N_13547);
nor U17112 (N_17112,N_14421,N_14595);
nand U17113 (N_17113,N_13156,N_14693);
or U17114 (N_17114,N_12545,N_14326);
or U17115 (N_17115,N_14089,N_14011);
or U17116 (N_17116,N_13317,N_13586);
and U17117 (N_17117,N_12264,N_13165);
nand U17118 (N_17118,N_14978,N_14216);
or U17119 (N_17119,N_12468,N_13221);
nand U17120 (N_17120,N_13643,N_13018);
nor U17121 (N_17121,N_14844,N_12133);
and U17122 (N_17122,N_13803,N_14245);
nor U17123 (N_17123,N_13726,N_12279);
xor U17124 (N_17124,N_13803,N_14861);
or U17125 (N_17125,N_14695,N_12248);
xnor U17126 (N_17126,N_14568,N_13590);
nand U17127 (N_17127,N_12715,N_12872);
nor U17128 (N_17128,N_13491,N_12864);
nor U17129 (N_17129,N_12972,N_13676);
nor U17130 (N_17130,N_13256,N_14958);
nor U17131 (N_17131,N_12726,N_12364);
nor U17132 (N_17132,N_12179,N_14790);
nand U17133 (N_17133,N_12016,N_14267);
nor U17134 (N_17134,N_14789,N_13969);
or U17135 (N_17135,N_13681,N_14569);
and U17136 (N_17136,N_14287,N_14420);
nand U17137 (N_17137,N_13961,N_13672);
xnor U17138 (N_17138,N_12779,N_13810);
and U17139 (N_17139,N_14486,N_14421);
nand U17140 (N_17140,N_13134,N_14936);
xor U17141 (N_17141,N_12514,N_13773);
xor U17142 (N_17142,N_13163,N_13858);
and U17143 (N_17143,N_13146,N_14133);
xnor U17144 (N_17144,N_13572,N_14803);
nand U17145 (N_17145,N_12512,N_12575);
nor U17146 (N_17146,N_12199,N_14038);
and U17147 (N_17147,N_14401,N_13243);
or U17148 (N_17148,N_13438,N_14098);
nor U17149 (N_17149,N_12462,N_13799);
nand U17150 (N_17150,N_12868,N_12761);
xor U17151 (N_17151,N_12076,N_13451);
xnor U17152 (N_17152,N_14895,N_12350);
nand U17153 (N_17153,N_12211,N_13266);
nand U17154 (N_17154,N_13762,N_12098);
xor U17155 (N_17155,N_13591,N_14375);
or U17156 (N_17156,N_12392,N_14738);
and U17157 (N_17157,N_13941,N_12429);
xnor U17158 (N_17158,N_12831,N_13892);
nand U17159 (N_17159,N_13959,N_13322);
and U17160 (N_17160,N_13169,N_12838);
or U17161 (N_17161,N_12024,N_14876);
or U17162 (N_17162,N_14696,N_12375);
nand U17163 (N_17163,N_12933,N_13982);
nor U17164 (N_17164,N_12559,N_14689);
or U17165 (N_17165,N_12483,N_14374);
xnor U17166 (N_17166,N_14121,N_12957);
or U17167 (N_17167,N_13335,N_14887);
and U17168 (N_17168,N_14802,N_12927);
nand U17169 (N_17169,N_12029,N_14794);
nand U17170 (N_17170,N_12833,N_12196);
or U17171 (N_17171,N_13231,N_14496);
nand U17172 (N_17172,N_14525,N_12746);
and U17173 (N_17173,N_13225,N_14887);
nor U17174 (N_17174,N_14222,N_13396);
xnor U17175 (N_17175,N_13776,N_13262);
nand U17176 (N_17176,N_14368,N_13155);
or U17177 (N_17177,N_12845,N_14663);
and U17178 (N_17178,N_13953,N_13807);
and U17179 (N_17179,N_14532,N_12144);
nand U17180 (N_17180,N_12071,N_12975);
xnor U17181 (N_17181,N_13798,N_12401);
nor U17182 (N_17182,N_14063,N_12621);
or U17183 (N_17183,N_14198,N_12137);
nand U17184 (N_17184,N_12278,N_14374);
or U17185 (N_17185,N_12930,N_12445);
and U17186 (N_17186,N_13465,N_14220);
nor U17187 (N_17187,N_12902,N_13355);
nand U17188 (N_17188,N_12918,N_13670);
or U17189 (N_17189,N_13250,N_12717);
or U17190 (N_17190,N_14698,N_13006);
xnor U17191 (N_17191,N_12307,N_12642);
nor U17192 (N_17192,N_13451,N_13284);
and U17193 (N_17193,N_12920,N_14011);
xor U17194 (N_17194,N_12454,N_13198);
and U17195 (N_17195,N_13760,N_12781);
or U17196 (N_17196,N_14604,N_13988);
and U17197 (N_17197,N_12791,N_14134);
nor U17198 (N_17198,N_14711,N_14553);
xnor U17199 (N_17199,N_14155,N_12314);
xor U17200 (N_17200,N_13615,N_12484);
nand U17201 (N_17201,N_14239,N_13980);
or U17202 (N_17202,N_14050,N_12482);
or U17203 (N_17203,N_12844,N_12373);
nor U17204 (N_17204,N_13919,N_14355);
xor U17205 (N_17205,N_12957,N_14126);
nand U17206 (N_17206,N_14235,N_14206);
xnor U17207 (N_17207,N_14380,N_13737);
xor U17208 (N_17208,N_14002,N_13058);
xor U17209 (N_17209,N_12839,N_12200);
nor U17210 (N_17210,N_14444,N_12333);
nand U17211 (N_17211,N_12545,N_13155);
or U17212 (N_17212,N_14139,N_13035);
or U17213 (N_17213,N_13413,N_13873);
xor U17214 (N_17214,N_12655,N_12336);
or U17215 (N_17215,N_14154,N_14874);
nor U17216 (N_17216,N_13915,N_14807);
xnor U17217 (N_17217,N_12854,N_14857);
or U17218 (N_17218,N_14494,N_14438);
xor U17219 (N_17219,N_14892,N_13554);
xor U17220 (N_17220,N_14880,N_13367);
xnor U17221 (N_17221,N_12161,N_14457);
or U17222 (N_17222,N_14268,N_14996);
nand U17223 (N_17223,N_12907,N_12192);
nand U17224 (N_17224,N_12457,N_12402);
and U17225 (N_17225,N_14681,N_12708);
nor U17226 (N_17226,N_14004,N_14064);
or U17227 (N_17227,N_14494,N_13286);
and U17228 (N_17228,N_14206,N_13206);
and U17229 (N_17229,N_12390,N_13081);
xor U17230 (N_17230,N_13507,N_13480);
or U17231 (N_17231,N_13048,N_12970);
and U17232 (N_17232,N_12722,N_13898);
or U17233 (N_17233,N_13142,N_13190);
nor U17234 (N_17234,N_14591,N_12655);
and U17235 (N_17235,N_13412,N_12945);
or U17236 (N_17236,N_14063,N_14751);
nor U17237 (N_17237,N_13057,N_13623);
xnor U17238 (N_17238,N_12528,N_12882);
nor U17239 (N_17239,N_14300,N_12756);
or U17240 (N_17240,N_12958,N_13258);
and U17241 (N_17241,N_13544,N_13614);
nand U17242 (N_17242,N_14188,N_13856);
nor U17243 (N_17243,N_13967,N_14674);
nand U17244 (N_17244,N_12225,N_14481);
or U17245 (N_17245,N_13349,N_14557);
or U17246 (N_17246,N_14457,N_13377);
or U17247 (N_17247,N_13927,N_13981);
nand U17248 (N_17248,N_12254,N_14044);
nor U17249 (N_17249,N_12491,N_13435);
and U17250 (N_17250,N_13758,N_14352);
and U17251 (N_17251,N_14251,N_14764);
nand U17252 (N_17252,N_14454,N_12594);
or U17253 (N_17253,N_12467,N_12458);
nand U17254 (N_17254,N_12348,N_14382);
or U17255 (N_17255,N_12439,N_12934);
or U17256 (N_17256,N_13719,N_14764);
xor U17257 (N_17257,N_12620,N_13775);
and U17258 (N_17258,N_13653,N_13777);
or U17259 (N_17259,N_13422,N_13003);
or U17260 (N_17260,N_13467,N_14198);
or U17261 (N_17261,N_13635,N_13812);
nand U17262 (N_17262,N_14852,N_12792);
nand U17263 (N_17263,N_14917,N_14592);
and U17264 (N_17264,N_13965,N_14278);
and U17265 (N_17265,N_12284,N_12021);
or U17266 (N_17266,N_13300,N_14752);
and U17267 (N_17267,N_13374,N_13394);
or U17268 (N_17268,N_14954,N_14280);
or U17269 (N_17269,N_12895,N_13403);
or U17270 (N_17270,N_13939,N_12035);
or U17271 (N_17271,N_14671,N_13677);
xnor U17272 (N_17272,N_14266,N_13028);
or U17273 (N_17273,N_13706,N_13103);
xor U17274 (N_17274,N_13158,N_14131);
nand U17275 (N_17275,N_14984,N_12297);
nand U17276 (N_17276,N_13697,N_14835);
and U17277 (N_17277,N_14108,N_14900);
xnor U17278 (N_17278,N_13294,N_14078);
and U17279 (N_17279,N_14506,N_12725);
xor U17280 (N_17280,N_14699,N_14518);
nand U17281 (N_17281,N_14735,N_12241);
or U17282 (N_17282,N_14394,N_12130);
nand U17283 (N_17283,N_14726,N_13403);
nor U17284 (N_17284,N_13141,N_13693);
and U17285 (N_17285,N_14180,N_14575);
nand U17286 (N_17286,N_13677,N_14644);
nand U17287 (N_17287,N_13332,N_12935);
xor U17288 (N_17288,N_13141,N_12652);
or U17289 (N_17289,N_14654,N_12673);
nand U17290 (N_17290,N_14117,N_14432);
xor U17291 (N_17291,N_14375,N_13098);
nor U17292 (N_17292,N_14648,N_12840);
or U17293 (N_17293,N_14703,N_12355);
and U17294 (N_17294,N_14688,N_14803);
xnor U17295 (N_17295,N_12275,N_12678);
nor U17296 (N_17296,N_13643,N_13182);
or U17297 (N_17297,N_14811,N_14024);
nand U17298 (N_17298,N_14522,N_14809);
xor U17299 (N_17299,N_14323,N_14765);
and U17300 (N_17300,N_12867,N_14198);
and U17301 (N_17301,N_14733,N_12107);
nor U17302 (N_17302,N_13374,N_12007);
nand U17303 (N_17303,N_14519,N_13172);
nand U17304 (N_17304,N_13275,N_13515);
nor U17305 (N_17305,N_12422,N_13521);
and U17306 (N_17306,N_12147,N_12175);
nand U17307 (N_17307,N_14387,N_13776);
and U17308 (N_17308,N_13032,N_14128);
nand U17309 (N_17309,N_13191,N_12280);
and U17310 (N_17310,N_13349,N_13270);
xor U17311 (N_17311,N_14303,N_13989);
xor U17312 (N_17312,N_12482,N_12985);
or U17313 (N_17313,N_12634,N_13460);
or U17314 (N_17314,N_13473,N_14206);
nor U17315 (N_17315,N_13936,N_14272);
and U17316 (N_17316,N_12282,N_13926);
xor U17317 (N_17317,N_13632,N_14709);
nor U17318 (N_17318,N_12159,N_12999);
nand U17319 (N_17319,N_12134,N_14411);
nor U17320 (N_17320,N_12269,N_12985);
or U17321 (N_17321,N_14668,N_13185);
and U17322 (N_17322,N_14453,N_12469);
xnor U17323 (N_17323,N_13840,N_12756);
or U17324 (N_17324,N_12460,N_12942);
and U17325 (N_17325,N_14816,N_14547);
nand U17326 (N_17326,N_13297,N_13825);
and U17327 (N_17327,N_12206,N_13575);
and U17328 (N_17328,N_13493,N_14850);
xor U17329 (N_17329,N_14721,N_12865);
or U17330 (N_17330,N_12309,N_12717);
nand U17331 (N_17331,N_14971,N_14284);
nor U17332 (N_17332,N_13275,N_14283);
xor U17333 (N_17333,N_14897,N_14321);
or U17334 (N_17334,N_12734,N_14129);
nor U17335 (N_17335,N_14918,N_12177);
or U17336 (N_17336,N_14971,N_12526);
nor U17337 (N_17337,N_14748,N_14891);
nor U17338 (N_17338,N_13685,N_14544);
and U17339 (N_17339,N_13649,N_14935);
and U17340 (N_17340,N_13828,N_12619);
nand U17341 (N_17341,N_13087,N_14061);
xor U17342 (N_17342,N_14006,N_13073);
nor U17343 (N_17343,N_13522,N_13295);
or U17344 (N_17344,N_13287,N_12569);
and U17345 (N_17345,N_13606,N_14672);
nand U17346 (N_17346,N_12987,N_14142);
xor U17347 (N_17347,N_12908,N_14756);
xor U17348 (N_17348,N_14207,N_14610);
xor U17349 (N_17349,N_13773,N_13379);
or U17350 (N_17350,N_12129,N_12104);
or U17351 (N_17351,N_12186,N_13612);
or U17352 (N_17352,N_14926,N_14821);
nor U17353 (N_17353,N_14807,N_13801);
and U17354 (N_17354,N_12922,N_14979);
and U17355 (N_17355,N_13195,N_14932);
and U17356 (N_17356,N_12291,N_14314);
nand U17357 (N_17357,N_12447,N_14845);
and U17358 (N_17358,N_12747,N_14226);
and U17359 (N_17359,N_12704,N_14190);
and U17360 (N_17360,N_13890,N_12888);
xnor U17361 (N_17361,N_12316,N_13227);
nor U17362 (N_17362,N_12644,N_12330);
nand U17363 (N_17363,N_12732,N_12279);
nor U17364 (N_17364,N_14850,N_12217);
xnor U17365 (N_17365,N_14297,N_14091);
xor U17366 (N_17366,N_12410,N_14721);
or U17367 (N_17367,N_12518,N_14757);
xnor U17368 (N_17368,N_12841,N_12625);
nor U17369 (N_17369,N_14232,N_12225);
nand U17370 (N_17370,N_13814,N_13448);
and U17371 (N_17371,N_14187,N_13456);
and U17372 (N_17372,N_12498,N_13217);
or U17373 (N_17373,N_12743,N_14143);
xnor U17374 (N_17374,N_13724,N_14638);
nor U17375 (N_17375,N_13171,N_14467);
or U17376 (N_17376,N_12463,N_13288);
or U17377 (N_17377,N_14081,N_12348);
xnor U17378 (N_17378,N_13540,N_13585);
nand U17379 (N_17379,N_12539,N_13244);
and U17380 (N_17380,N_12366,N_14129);
nand U17381 (N_17381,N_14073,N_13748);
xor U17382 (N_17382,N_12296,N_14547);
nand U17383 (N_17383,N_12211,N_14048);
nand U17384 (N_17384,N_12620,N_14310);
nand U17385 (N_17385,N_12117,N_14906);
nor U17386 (N_17386,N_12294,N_13167);
or U17387 (N_17387,N_13210,N_14481);
and U17388 (N_17388,N_12844,N_14305);
or U17389 (N_17389,N_13311,N_13468);
xnor U17390 (N_17390,N_13581,N_12542);
and U17391 (N_17391,N_14224,N_12626);
or U17392 (N_17392,N_14988,N_12161);
nand U17393 (N_17393,N_14793,N_14559);
and U17394 (N_17394,N_13524,N_14813);
or U17395 (N_17395,N_14876,N_12505);
nand U17396 (N_17396,N_12035,N_13639);
or U17397 (N_17397,N_13243,N_12446);
nand U17398 (N_17398,N_13388,N_12885);
and U17399 (N_17399,N_12253,N_14056);
or U17400 (N_17400,N_14870,N_14511);
and U17401 (N_17401,N_13601,N_13769);
xnor U17402 (N_17402,N_12786,N_13389);
nand U17403 (N_17403,N_14688,N_13184);
xor U17404 (N_17404,N_14491,N_12058);
xor U17405 (N_17405,N_14513,N_12735);
nand U17406 (N_17406,N_13997,N_13407);
nor U17407 (N_17407,N_12809,N_12575);
xnor U17408 (N_17408,N_12065,N_12069);
nand U17409 (N_17409,N_12154,N_14648);
nor U17410 (N_17410,N_13706,N_14740);
xor U17411 (N_17411,N_12083,N_12271);
xnor U17412 (N_17412,N_12707,N_14664);
or U17413 (N_17413,N_14070,N_12106);
and U17414 (N_17414,N_12784,N_13256);
nand U17415 (N_17415,N_12410,N_14155);
or U17416 (N_17416,N_14262,N_13906);
and U17417 (N_17417,N_12078,N_13455);
and U17418 (N_17418,N_12500,N_13854);
nor U17419 (N_17419,N_13290,N_13896);
nor U17420 (N_17420,N_13535,N_13543);
xnor U17421 (N_17421,N_14586,N_12462);
nand U17422 (N_17422,N_12817,N_12800);
xor U17423 (N_17423,N_13236,N_14530);
or U17424 (N_17424,N_13941,N_12380);
nor U17425 (N_17425,N_12732,N_14992);
nor U17426 (N_17426,N_13982,N_12979);
nor U17427 (N_17427,N_13817,N_14902);
xor U17428 (N_17428,N_14559,N_12644);
or U17429 (N_17429,N_13380,N_14014);
nand U17430 (N_17430,N_14015,N_12749);
or U17431 (N_17431,N_12759,N_13586);
nor U17432 (N_17432,N_12760,N_14904);
xnor U17433 (N_17433,N_14761,N_14205);
nor U17434 (N_17434,N_14507,N_14502);
or U17435 (N_17435,N_12836,N_12077);
nor U17436 (N_17436,N_12195,N_14914);
and U17437 (N_17437,N_12800,N_12123);
nand U17438 (N_17438,N_14769,N_14782);
nand U17439 (N_17439,N_12938,N_14915);
nand U17440 (N_17440,N_13718,N_14554);
and U17441 (N_17441,N_12976,N_14587);
xor U17442 (N_17442,N_12237,N_12260);
nand U17443 (N_17443,N_14939,N_14344);
and U17444 (N_17444,N_14505,N_13424);
xor U17445 (N_17445,N_12597,N_12193);
nor U17446 (N_17446,N_13929,N_14738);
xnor U17447 (N_17447,N_13373,N_13684);
xor U17448 (N_17448,N_13391,N_12911);
or U17449 (N_17449,N_12480,N_13199);
and U17450 (N_17450,N_12212,N_12996);
nor U17451 (N_17451,N_14766,N_14002);
or U17452 (N_17452,N_12327,N_12817);
and U17453 (N_17453,N_14629,N_12091);
and U17454 (N_17454,N_14317,N_14520);
and U17455 (N_17455,N_12773,N_13152);
nand U17456 (N_17456,N_12959,N_13382);
or U17457 (N_17457,N_13263,N_13818);
or U17458 (N_17458,N_13231,N_12222);
nor U17459 (N_17459,N_13222,N_14652);
nor U17460 (N_17460,N_12230,N_14645);
or U17461 (N_17461,N_14581,N_12654);
and U17462 (N_17462,N_12236,N_12110);
xnor U17463 (N_17463,N_12880,N_14493);
and U17464 (N_17464,N_12957,N_12680);
nor U17465 (N_17465,N_12385,N_14851);
or U17466 (N_17466,N_12271,N_13414);
xnor U17467 (N_17467,N_13702,N_12654);
and U17468 (N_17468,N_12539,N_14852);
nor U17469 (N_17469,N_13619,N_12348);
xnor U17470 (N_17470,N_13985,N_14350);
nand U17471 (N_17471,N_14242,N_13789);
xor U17472 (N_17472,N_12423,N_12236);
and U17473 (N_17473,N_12461,N_14019);
xnor U17474 (N_17474,N_13633,N_13655);
nor U17475 (N_17475,N_14903,N_13890);
xor U17476 (N_17476,N_13102,N_14833);
and U17477 (N_17477,N_13824,N_12928);
nor U17478 (N_17478,N_12945,N_13251);
xnor U17479 (N_17479,N_14634,N_13281);
nand U17480 (N_17480,N_12831,N_12893);
nand U17481 (N_17481,N_12017,N_14653);
xor U17482 (N_17482,N_12990,N_13022);
and U17483 (N_17483,N_14902,N_12145);
nor U17484 (N_17484,N_14891,N_12395);
or U17485 (N_17485,N_14303,N_12103);
and U17486 (N_17486,N_13830,N_14179);
xor U17487 (N_17487,N_12454,N_13299);
nor U17488 (N_17488,N_12625,N_13475);
or U17489 (N_17489,N_13681,N_12662);
or U17490 (N_17490,N_12949,N_14875);
and U17491 (N_17491,N_12661,N_14612);
and U17492 (N_17492,N_12058,N_12165);
or U17493 (N_17493,N_14587,N_14737);
nand U17494 (N_17494,N_13750,N_13019);
and U17495 (N_17495,N_13705,N_13323);
and U17496 (N_17496,N_12923,N_14147);
nor U17497 (N_17497,N_13482,N_13135);
or U17498 (N_17498,N_12446,N_14801);
nand U17499 (N_17499,N_12240,N_14012);
nor U17500 (N_17500,N_12228,N_14028);
and U17501 (N_17501,N_13176,N_12511);
nand U17502 (N_17502,N_13099,N_13188);
xor U17503 (N_17503,N_14356,N_13607);
nor U17504 (N_17504,N_14830,N_12123);
xnor U17505 (N_17505,N_14633,N_12939);
nand U17506 (N_17506,N_12816,N_12750);
nand U17507 (N_17507,N_12861,N_13757);
and U17508 (N_17508,N_14764,N_14133);
nand U17509 (N_17509,N_14325,N_12061);
nand U17510 (N_17510,N_14573,N_13453);
xnor U17511 (N_17511,N_14816,N_13818);
or U17512 (N_17512,N_12253,N_14301);
nand U17513 (N_17513,N_14448,N_13717);
nor U17514 (N_17514,N_13886,N_14874);
and U17515 (N_17515,N_12701,N_14587);
xor U17516 (N_17516,N_12404,N_12240);
or U17517 (N_17517,N_12278,N_14564);
or U17518 (N_17518,N_14438,N_14522);
xor U17519 (N_17519,N_12454,N_13108);
or U17520 (N_17520,N_13362,N_14099);
nand U17521 (N_17521,N_13485,N_14918);
and U17522 (N_17522,N_12311,N_13200);
nand U17523 (N_17523,N_14552,N_14688);
and U17524 (N_17524,N_14118,N_13906);
xnor U17525 (N_17525,N_13904,N_12065);
nor U17526 (N_17526,N_12203,N_13891);
xnor U17527 (N_17527,N_13849,N_14980);
nor U17528 (N_17528,N_13050,N_12198);
nor U17529 (N_17529,N_13351,N_12120);
and U17530 (N_17530,N_12754,N_14997);
nor U17531 (N_17531,N_14158,N_13200);
nand U17532 (N_17532,N_13005,N_12226);
or U17533 (N_17533,N_13510,N_14141);
or U17534 (N_17534,N_13368,N_14090);
xnor U17535 (N_17535,N_14590,N_14227);
nand U17536 (N_17536,N_12738,N_12239);
nor U17537 (N_17537,N_14574,N_13302);
nor U17538 (N_17538,N_13736,N_12850);
xor U17539 (N_17539,N_12267,N_13013);
and U17540 (N_17540,N_12378,N_13008);
and U17541 (N_17541,N_12271,N_12124);
and U17542 (N_17542,N_14114,N_14714);
or U17543 (N_17543,N_12225,N_14624);
nand U17544 (N_17544,N_12484,N_13911);
and U17545 (N_17545,N_13427,N_12222);
nand U17546 (N_17546,N_12167,N_14215);
xor U17547 (N_17547,N_14643,N_12050);
nor U17548 (N_17548,N_12978,N_14809);
nor U17549 (N_17549,N_12114,N_13299);
or U17550 (N_17550,N_12542,N_13610);
and U17551 (N_17551,N_12198,N_12350);
nor U17552 (N_17552,N_14800,N_13743);
nand U17553 (N_17553,N_12843,N_14064);
and U17554 (N_17554,N_14910,N_14005);
and U17555 (N_17555,N_13544,N_14538);
and U17556 (N_17556,N_14370,N_14527);
and U17557 (N_17557,N_12253,N_12564);
nor U17558 (N_17558,N_13367,N_14514);
xnor U17559 (N_17559,N_14676,N_13448);
or U17560 (N_17560,N_13079,N_13719);
and U17561 (N_17561,N_12631,N_14175);
and U17562 (N_17562,N_12906,N_13611);
nand U17563 (N_17563,N_13182,N_13404);
nand U17564 (N_17564,N_14277,N_13422);
nand U17565 (N_17565,N_14998,N_13420);
xor U17566 (N_17566,N_14954,N_12814);
and U17567 (N_17567,N_12674,N_12290);
xor U17568 (N_17568,N_12353,N_13989);
xor U17569 (N_17569,N_12307,N_12480);
nand U17570 (N_17570,N_14677,N_13410);
and U17571 (N_17571,N_12467,N_12172);
or U17572 (N_17572,N_14072,N_13805);
nor U17573 (N_17573,N_13970,N_14536);
nand U17574 (N_17574,N_12045,N_14395);
xnor U17575 (N_17575,N_12002,N_12140);
or U17576 (N_17576,N_12416,N_12007);
and U17577 (N_17577,N_13000,N_12474);
nand U17578 (N_17578,N_12846,N_12724);
and U17579 (N_17579,N_13027,N_12463);
nand U17580 (N_17580,N_13808,N_13586);
xnor U17581 (N_17581,N_14122,N_14230);
and U17582 (N_17582,N_13257,N_14028);
or U17583 (N_17583,N_14176,N_13939);
xor U17584 (N_17584,N_13435,N_14053);
or U17585 (N_17585,N_12791,N_14046);
nor U17586 (N_17586,N_13147,N_13743);
and U17587 (N_17587,N_12505,N_12996);
and U17588 (N_17588,N_14916,N_13425);
and U17589 (N_17589,N_14695,N_13608);
xnor U17590 (N_17590,N_12475,N_14672);
nand U17591 (N_17591,N_14027,N_12992);
and U17592 (N_17592,N_12743,N_14002);
and U17593 (N_17593,N_13317,N_14849);
nor U17594 (N_17594,N_12591,N_14983);
nor U17595 (N_17595,N_13765,N_12114);
xnor U17596 (N_17596,N_12554,N_13152);
nand U17597 (N_17597,N_12587,N_12753);
nor U17598 (N_17598,N_14202,N_13564);
nor U17599 (N_17599,N_14318,N_14719);
or U17600 (N_17600,N_14930,N_14767);
nand U17601 (N_17601,N_13269,N_12338);
and U17602 (N_17602,N_13255,N_14992);
and U17603 (N_17603,N_14380,N_12296);
or U17604 (N_17604,N_13947,N_12605);
and U17605 (N_17605,N_13619,N_14757);
and U17606 (N_17606,N_13005,N_12648);
and U17607 (N_17607,N_14647,N_12410);
nand U17608 (N_17608,N_12303,N_12129);
xnor U17609 (N_17609,N_12581,N_13711);
nor U17610 (N_17610,N_13020,N_12469);
and U17611 (N_17611,N_14103,N_14605);
nor U17612 (N_17612,N_13369,N_12340);
or U17613 (N_17613,N_13381,N_14117);
and U17614 (N_17614,N_13534,N_13338);
or U17615 (N_17615,N_14739,N_12854);
or U17616 (N_17616,N_14890,N_12058);
nand U17617 (N_17617,N_12987,N_12338);
xnor U17618 (N_17618,N_14893,N_13538);
or U17619 (N_17619,N_12416,N_13037);
and U17620 (N_17620,N_12947,N_14843);
or U17621 (N_17621,N_12067,N_13310);
xnor U17622 (N_17622,N_12883,N_14700);
and U17623 (N_17623,N_14944,N_13486);
xor U17624 (N_17624,N_14912,N_12176);
xnor U17625 (N_17625,N_12819,N_14395);
and U17626 (N_17626,N_12353,N_13125);
nor U17627 (N_17627,N_12320,N_13909);
and U17628 (N_17628,N_14419,N_14427);
or U17629 (N_17629,N_13037,N_12399);
or U17630 (N_17630,N_12650,N_13463);
nor U17631 (N_17631,N_14163,N_14872);
xor U17632 (N_17632,N_12690,N_13479);
xor U17633 (N_17633,N_14168,N_13906);
nor U17634 (N_17634,N_12247,N_14483);
or U17635 (N_17635,N_14850,N_13599);
nand U17636 (N_17636,N_13345,N_14467);
or U17637 (N_17637,N_12275,N_14911);
or U17638 (N_17638,N_13301,N_12468);
and U17639 (N_17639,N_12851,N_14409);
xnor U17640 (N_17640,N_12276,N_13275);
nand U17641 (N_17641,N_12349,N_12739);
or U17642 (N_17642,N_12617,N_13460);
nor U17643 (N_17643,N_13652,N_12501);
nor U17644 (N_17644,N_12340,N_14556);
nor U17645 (N_17645,N_12835,N_13712);
or U17646 (N_17646,N_13845,N_12061);
and U17647 (N_17647,N_14020,N_14367);
nor U17648 (N_17648,N_13059,N_13377);
xnor U17649 (N_17649,N_12674,N_13697);
nand U17650 (N_17650,N_14326,N_12479);
nand U17651 (N_17651,N_12299,N_13333);
nor U17652 (N_17652,N_12945,N_13309);
nor U17653 (N_17653,N_14207,N_12290);
nor U17654 (N_17654,N_14842,N_13670);
or U17655 (N_17655,N_12630,N_14048);
nand U17656 (N_17656,N_13045,N_12297);
nor U17657 (N_17657,N_13915,N_12540);
xnor U17658 (N_17658,N_12862,N_14558);
and U17659 (N_17659,N_14798,N_14484);
nand U17660 (N_17660,N_12567,N_13937);
xnor U17661 (N_17661,N_14521,N_14586);
nand U17662 (N_17662,N_13125,N_13732);
nor U17663 (N_17663,N_14098,N_12039);
nor U17664 (N_17664,N_13741,N_12701);
xor U17665 (N_17665,N_14097,N_12448);
xor U17666 (N_17666,N_12351,N_13124);
nand U17667 (N_17667,N_14315,N_14744);
nand U17668 (N_17668,N_14496,N_13783);
and U17669 (N_17669,N_12891,N_14059);
xor U17670 (N_17670,N_14621,N_12644);
xor U17671 (N_17671,N_13399,N_14698);
xnor U17672 (N_17672,N_12321,N_12510);
or U17673 (N_17673,N_12372,N_13691);
nand U17674 (N_17674,N_14361,N_12127);
and U17675 (N_17675,N_12353,N_12160);
or U17676 (N_17676,N_14453,N_12443);
xnor U17677 (N_17677,N_14686,N_12575);
nand U17678 (N_17678,N_13564,N_14425);
nor U17679 (N_17679,N_13319,N_12757);
xor U17680 (N_17680,N_13191,N_14435);
xor U17681 (N_17681,N_14531,N_14483);
xor U17682 (N_17682,N_13854,N_13604);
or U17683 (N_17683,N_13266,N_14788);
nor U17684 (N_17684,N_14274,N_12118);
xor U17685 (N_17685,N_14194,N_14454);
xnor U17686 (N_17686,N_13351,N_12067);
nor U17687 (N_17687,N_13361,N_14795);
and U17688 (N_17688,N_13214,N_14645);
nand U17689 (N_17689,N_12812,N_12214);
and U17690 (N_17690,N_12085,N_13691);
and U17691 (N_17691,N_14900,N_14603);
or U17692 (N_17692,N_14602,N_14236);
nor U17693 (N_17693,N_12035,N_14419);
nand U17694 (N_17694,N_13512,N_14196);
or U17695 (N_17695,N_12433,N_12970);
nor U17696 (N_17696,N_13632,N_14824);
or U17697 (N_17697,N_12417,N_14714);
xnor U17698 (N_17698,N_12630,N_14146);
or U17699 (N_17699,N_12020,N_14425);
and U17700 (N_17700,N_14831,N_12074);
nor U17701 (N_17701,N_13249,N_14480);
xor U17702 (N_17702,N_14849,N_13679);
nand U17703 (N_17703,N_12948,N_14654);
or U17704 (N_17704,N_13804,N_14181);
or U17705 (N_17705,N_13171,N_14880);
nand U17706 (N_17706,N_13060,N_14665);
nand U17707 (N_17707,N_14718,N_12062);
xnor U17708 (N_17708,N_13999,N_12288);
or U17709 (N_17709,N_12625,N_13234);
and U17710 (N_17710,N_12461,N_14601);
and U17711 (N_17711,N_12776,N_13534);
or U17712 (N_17712,N_14260,N_13657);
and U17713 (N_17713,N_13210,N_13089);
nor U17714 (N_17714,N_14505,N_12359);
nor U17715 (N_17715,N_13907,N_14547);
and U17716 (N_17716,N_13553,N_12682);
xnor U17717 (N_17717,N_14681,N_14548);
or U17718 (N_17718,N_13355,N_14048);
nor U17719 (N_17719,N_13308,N_13714);
xor U17720 (N_17720,N_13767,N_13323);
and U17721 (N_17721,N_13885,N_12797);
and U17722 (N_17722,N_13160,N_12960);
xor U17723 (N_17723,N_12170,N_13723);
or U17724 (N_17724,N_13846,N_12810);
xnor U17725 (N_17725,N_13779,N_12038);
and U17726 (N_17726,N_13231,N_13485);
xnor U17727 (N_17727,N_14460,N_12366);
xnor U17728 (N_17728,N_14733,N_14597);
and U17729 (N_17729,N_12422,N_14656);
nor U17730 (N_17730,N_13654,N_14808);
xnor U17731 (N_17731,N_12158,N_13994);
or U17732 (N_17732,N_12092,N_14805);
xor U17733 (N_17733,N_13891,N_12938);
nand U17734 (N_17734,N_13650,N_14516);
nand U17735 (N_17735,N_13672,N_13210);
and U17736 (N_17736,N_13080,N_13043);
and U17737 (N_17737,N_14675,N_12783);
nor U17738 (N_17738,N_13157,N_12141);
and U17739 (N_17739,N_14075,N_14061);
xnor U17740 (N_17740,N_13578,N_12045);
or U17741 (N_17741,N_13202,N_14520);
or U17742 (N_17742,N_14499,N_13700);
and U17743 (N_17743,N_14739,N_12692);
xnor U17744 (N_17744,N_12045,N_13914);
xor U17745 (N_17745,N_12036,N_13028);
nor U17746 (N_17746,N_14623,N_12495);
and U17747 (N_17747,N_12032,N_14020);
nor U17748 (N_17748,N_14679,N_13003);
or U17749 (N_17749,N_12917,N_14240);
xnor U17750 (N_17750,N_12201,N_12837);
and U17751 (N_17751,N_12643,N_14577);
and U17752 (N_17752,N_14108,N_12056);
nor U17753 (N_17753,N_14858,N_14432);
nand U17754 (N_17754,N_12646,N_13208);
nand U17755 (N_17755,N_14330,N_13185);
or U17756 (N_17756,N_14668,N_13571);
and U17757 (N_17757,N_13314,N_13971);
nand U17758 (N_17758,N_12698,N_13933);
nand U17759 (N_17759,N_13703,N_13386);
and U17760 (N_17760,N_12073,N_13761);
nor U17761 (N_17761,N_14262,N_13310);
nand U17762 (N_17762,N_13799,N_12995);
nand U17763 (N_17763,N_13985,N_12220);
and U17764 (N_17764,N_12375,N_12467);
and U17765 (N_17765,N_12784,N_13813);
or U17766 (N_17766,N_13196,N_12666);
or U17767 (N_17767,N_12431,N_14701);
nand U17768 (N_17768,N_12193,N_12569);
or U17769 (N_17769,N_13000,N_12954);
nand U17770 (N_17770,N_13290,N_13698);
or U17771 (N_17771,N_14234,N_14709);
nand U17772 (N_17772,N_14238,N_13899);
nor U17773 (N_17773,N_13466,N_13065);
xnor U17774 (N_17774,N_14597,N_13166);
nor U17775 (N_17775,N_12394,N_12584);
nor U17776 (N_17776,N_14316,N_12208);
or U17777 (N_17777,N_12544,N_13923);
xor U17778 (N_17778,N_14757,N_13087);
nand U17779 (N_17779,N_14674,N_12988);
and U17780 (N_17780,N_12731,N_13218);
or U17781 (N_17781,N_12237,N_13559);
nand U17782 (N_17782,N_13129,N_13240);
nor U17783 (N_17783,N_13842,N_14190);
and U17784 (N_17784,N_13773,N_14410);
nand U17785 (N_17785,N_12027,N_13519);
nand U17786 (N_17786,N_13228,N_12932);
nand U17787 (N_17787,N_12143,N_12576);
nand U17788 (N_17788,N_14566,N_12414);
and U17789 (N_17789,N_13522,N_14835);
and U17790 (N_17790,N_13219,N_14894);
nor U17791 (N_17791,N_12225,N_12512);
nor U17792 (N_17792,N_12126,N_14764);
and U17793 (N_17793,N_14870,N_12192);
xor U17794 (N_17794,N_12917,N_12899);
nor U17795 (N_17795,N_12099,N_14875);
nand U17796 (N_17796,N_13875,N_14902);
nor U17797 (N_17797,N_12646,N_12493);
or U17798 (N_17798,N_12280,N_14379);
or U17799 (N_17799,N_12540,N_12212);
xnor U17800 (N_17800,N_14654,N_12879);
or U17801 (N_17801,N_12916,N_14868);
xnor U17802 (N_17802,N_13030,N_12640);
and U17803 (N_17803,N_13599,N_13105);
nor U17804 (N_17804,N_13933,N_13385);
nor U17805 (N_17805,N_13914,N_12805);
nand U17806 (N_17806,N_12358,N_13212);
nor U17807 (N_17807,N_14083,N_13505);
or U17808 (N_17808,N_13447,N_12088);
or U17809 (N_17809,N_12467,N_12553);
nor U17810 (N_17810,N_13937,N_13212);
xnor U17811 (N_17811,N_12930,N_13649);
nor U17812 (N_17812,N_14342,N_12021);
xor U17813 (N_17813,N_14543,N_13787);
xor U17814 (N_17814,N_12914,N_14020);
and U17815 (N_17815,N_12552,N_14320);
nor U17816 (N_17816,N_14241,N_13880);
or U17817 (N_17817,N_12728,N_13918);
nor U17818 (N_17818,N_13470,N_14681);
nor U17819 (N_17819,N_12090,N_12231);
and U17820 (N_17820,N_14074,N_12346);
nand U17821 (N_17821,N_12304,N_13311);
xnor U17822 (N_17822,N_13075,N_14299);
nand U17823 (N_17823,N_14063,N_14657);
nand U17824 (N_17824,N_12429,N_13098);
xor U17825 (N_17825,N_12458,N_13547);
xor U17826 (N_17826,N_14015,N_12194);
nor U17827 (N_17827,N_14501,N_13258);
or U17828 (N_17828,N_12574,N_12146);
and U17829 (N_17829,N_12399,N_12060);
or U17830 (N_17830,N_12503,N_12513);
xor U17831 (N_17831,N_13636,N_12758);
nor U17832 (N_17832,N_12537,N_12351);
nand U17833 (N_17833,N_13785,N_13754);
nand U17834 (N_17834,N_13572,N_13003);
xnor U17835 (N_17835,N_13654,N_13791);
and U17836 (N_17836,N_13019,N_12660);
nand U17837 (N_17837,N_14204,N_13938);
or U17838 (N_17838,N_14857,N_12964);
nand U17839 (N_17839,N_12514,N_13846);
and U17840 (N_17840,N_12168,N_12493);
xnor U17841 (N_17841,N_12259,N_14065);
nor U17842 (N_17842,N_12458,N_13739);
or U17843 (N_17843,N_12763,N_14944);
nor U17844 (N_17844,N_14110,N_13088);
nand U17845 (N_17845,N_13384,N_14627);
and U17846 (N_17846,N_12210,N_12238);
and U17847 (N_17847,N_12243,N_13754);
or U17848 (N_17848,N_13351,N_14816);
or U17849 (N_17849,N_13136,N_12232);
nand U17850 (N_17850,N_13335,N_14124);
or U17851 (N_17851,N_13983,N_12360);
and U17852 (N_17852,N_12257,N_14935);
nand U17853 (N_17853,N_12115,N_14511);
nand U17854 (N_17854,N_13201,N_14721);
xor U17855 (N_17855,N_12324,N_14135);
nand U17856 (N_17856,N_12118,N_13533);
nor U17857 (N_17857,N_13228,N_12576);
xnor U17858 (N_17858,N_14243,N_13348);
xnor U17859 (N_17859,N_12137,N_14200);
xor U17860 (N_17860,N_12269,N_14501);
or U17861 (N_17861,N_12449,N_12558);
or U17862 (N_17862,N_14109,N_12019);
nor U17863 (N_17863,N_12263,N_13367);
or U17864 (N_17864,N_12678,N_13740);
and U17865 (N_17865,N_14641,N_13208);
nand U17866 (N_17866,N_13875,N_12481);
and U17867 (N_17867,N_12482,N_12013);
xnor U17868 (N_17868,N_12367,N_12435);
or U17869 (N_17869,N_13742,N_14961);
and U17870 (N_17870,N_14358,N_14490);
xnor U17871 (N_17871,N_12146,N_14585);
and U17872 (N_17872,N_12424,N_13851);
nand U17873 (N_17873,N_12041,N_13546);
xnor U17874 (N_17874,N_14535,N_13539);
xnor U17875 (N_17875,N_13583,N_12807);
and U17876 (N_17876,N_13740,N_13404);
nand U17877 (N_17877,N_14450,N_12429);
nor U17878 (N_17878,N_13090,N_12881);
nor U17879 (N_17879,N_13027,N_12172);
or U17880 (N_17880,N_12738,N_13695);
or U17881 (N_17881,N_14801,N_13163);
nand U17882 (N_17882,N_14457,N_12634);
nor U17883 (N_17883,N_14649,N_13036);
or U17884 (N_17884,N_13144,N_13820);
nand U17885 (N_17885,N_12193,N_14362);
or U17886 (N_17886,N_14665,N_13429);
nand U17887 (N_17887,N_12218,N_13735);
or U17888 (N_17888,N_14419,N_13352);
and U17889 (N_17889,N_13280,N_13176);
nor U17890 (N_17890,N_12805,N_13507);
or U17891 (N_17891,N_12787,N_14540);
nand U17892 (N_17892,N_13761,N_14391);
and U17893 (N_17893,N_13298,N_14172);
or U17894 (N_17894,N_13021,N_13851);
nor U17895 (N_17895,N_13287,N_12799);
or U17896 (N_17896,N_14891,N_13204);
nand U17897 (N_17897,N_12564,N_14434);
nor U17898 (N_17898,N_13089,N_14280);
xor U17899 (N_17899,N_12743,N_13932);
nand U17900 (N_17900,N_12872,N_14783);
xnor U17901 (N_17901,N_12094,N_12920);
or U17902 (N_17902,N_14018,N_12756);
nand U17903 (N_17903,N_12722,N_12536);
or U17904 (N_17904,N_14734,N_13434);
or U17905 (N_17905,N_12889,N_12884);
and U17906 (N_17906,N_13665,N_13527);
xnor U17907 (N_17907,N_13502,N_12306);
nand U17908 (N_17908,N_14032,N_13261);
and U17909 (N_17909,N_12001,N_14898);
nor U17910 (N_17910,N_14560,N_14192);
nor U17911 (N_17911,N_13126,N_13935);
or U17912 (N_17912,N_13359,N_12348);
or U17913 (N_17913,N_14631,N_13802);
nand U17914 (N_17914,N_13025,N_14579);
and U17915 (N_17915,N_12978,N_13099);
nor U17916 (N_17916,N_13627,N_14965);
xor U17917 (N_17917,N_14973,N_13676);
and U17918 (N_17918,N_13492,N_12292);
xor U17919 (N_17919,N_12341,N_12847);
and U17920 (N_17920,N_12938,N_14330);
nand U17921 (N_17921,N_12545,N_14850);
or U17922 (N_17922,N_12263,N_14044);
and U17923 (N_17923,N_12419,N_14545);
or U17924 (N_17924,N_12966,N_14026);
xor U17925 (N_17925,N_12665,N_14387);
and U17926 (N_17926,N_14077,N_12891);
nor U17927 (N_17927,N_12889,N_13474);
xor U17928 (N_17928,N_12489,N_14607);
nor U17929 (N_17929,N_13992,N_14995);
or U17930 (N_17930,N_13416,N_13116);
and U17931 (N_17931,N_12220,N_12032);
nor U17932 (N_17932,N_12829,N_12347);
nand U17933 (N_17933,N_14278,N_12985);
nand U17934 (N_17934,N_12796,N_13271);
nand U17935 (N_17935,N_13250,N_13300);
nand U17936 (N_17936,N_14042,N_14269);
nor U17937 (N_17937,N_14215,N_12784);
xnor U17938 (N_17938,N_13846,N_13618);
nand U17939 (N_17939,N_14168,N_12244);
or U17940 (N_17940,N_13062,N_13203);
or U17941 (N_17941,N_14657,N_12511);
and U17942 (N_17942,N_12435,N_12723);
xnor U17943 (N_17943,N_13974,N_12247);
nand U17944 (N_17944,N_14115,N_12153);
xnor U17945 (N_17945,N_13804,N_13337);
xnor U17946 (N_17946,N_12529,N_13525);
or U17947 (N_17947,N_14303,N_14016);
and U17948 (N_17948,N_13135,N_12576);
nor U17949 (N_17949,N_14558,N_13698);
and U17950 (N_17950,N_12923,N_14224);
nand U17951 (N_17951,N_14607,N_14759);
and U17952 (N_17952,N_14641,N_13451);
and U17953 (N_17953,N_14862,N_14461);
nand U17954 (N_17954,N_14501,N_14509);
or U17955 (N_17955,N_12223,N_13348);
and U17956 (N_17956,N_13333,N_12767);
nand U17957 (N_17957,N_12601,N_12799);
nor U17958 (N_17958,N_14738,N_13830);
xnor U17959 (N_17959,N_13323,N_12787);
xnor U17960 (N_17960,N_14617,N_14456);
and U17961 (N_17961,N_13134,N_12100);
nor U17962 (N_17962,N_14887,N_13497);
and U17963 (N_17963,N_14708,N_13978);
nor U17964 (N_17964,N_14561,N_12081);
nand U17965 (N_17965,N_14359,N_14011);
nand U17966 (N_17966,N_13700,N_12586);
or U17967 (N_17967,N_14377,N_13265);
nor U17968 (N_17968,N_13840,N_13552);
or U17969 (N_17969,N_12559,N_14812);
or U17970 (N_17970,N_14175,N_13342);
xnor U17971 (N_17971,N_13180,N_14413);
and U17972 (N_17972,N_12549,N_14429);
nand U17973 (N_17973,N_13246,N_14061);
xnor U17974 (N_17974,N_13883,N_14444);
nand U17975 (N_17975,N_14401,N_13013);
or U17976 (N_17976,N_14973,N_14816);
and U17977 (N_17977,N_13076,N_13877);
nand U17978 (N_17978,N_13675,N_14937);
nor U17979 (N_17979,N_12245,N_13975);
nor U17980 (N_17980,N_13684,N_14378);
or U17981 (N_17981,N_14931,N_14471);
and U17982 (N_17982,N_14635,N_12486);
or U17983 (N_17983,N_12477,N_14144);
and U17984 (N_17984,N_12142,N_14175);
or U17985 (N_17985,N_12475,N_12132);
or U17986 (N_17986,N_13361,N_12986);
and U17987 (N_17987,N_13777,N_12253);
nor U17988 (N_17988,N_14328,N_12555);
nor U17989 (N_17989,N_14700,N_14420);
or U17990 (N_17990,N_14525,N_14539);
nor U17991 (N_17991,N_14977,N_14815);
or U17992 (N_17992,N_14156,N_13562);
xnor U17993 (N_17993,N_12657,N_14058);
or U17994 (N_17994,N_13585,N_13203);
and U17995 (N_17995,N_12354,N_12797);
or U17996 (N_17996,N_13359,N_12185);
xnor U17997 (N_17997,N_14152,N_13200);
nand U17998 (N_17998,N_13155,N_14600);
or U17999 (N_17999,N_14309,N_14266);
or U18000 (N_18000,N_16709,N_16725);
nor U18001 (N_18001,N_17927,N_16255);
or U18002 (N_18002,N_15170,N_16933);
or U18003 (N_18003,N_17934,N_17545);
or U18004 (N_18004,N_16515,N_17039);
nand U18005 (N_18005,N_15660,N_16011);
nor U18006 (N_18006,N_16049,N_17506);
or U18007 (N_18007,N_16394,N_16270);
nand U18008 (N_18008,N_16641,N_16114);
nand U18009 (N_18009,N_16189,N_17003);
nand U18010 (N_18010,N_16617,N_16159);
nand U18011 (N_18011,N_16633,N_16964);
or U18012 (N_18012,N_16042,N_17301);
or U18013 (N_18013,N_16952,N_17219);
nor U18014 (N_18014,N_17200,N_16496);
or U18015 (N_18015,N_15398,N_16040);
or U18016 (N_18016,N_17754,N_16754);
and U18017 (N_18017,N_17243,N_16970);
and U18018 (N_18018,N_15132,N_15203);
or U18019 (N_18019,N_17220,N_16008);
and U18020 (N_18020,N_17151,N_15523);
nor U18021 (N_18021,N_16955,N_15618);
or U18022 (N_18022,N_17019,N_17153);
nand U18023 (N_18023,N_15179,N_16456);
nand U18024 (N_18024,N_16390,N_15668);
and U18025 (N_18025,N_17992,N_17907);
or U18026 (N_18026,N_16518,N_16358);
or U18027 (N_18027,N_16986,N_16648);
and U18028 (N_18028,N_16794,N_15727);
and U18029 (N_18029,N_15544,N_16561);
or U18030 (N_18030,N_16029,N_15961);
nor U18031 (N_18031,N_15886,N_16421);
nor U18032 (N_18032,N_17840,N_16027);
nor U18033 (N_18033,N_17702,N_15532);
or U18034 (N_18034,N_17511,N_17461);
nand U18035 (N_18035,N_16438,N_15837);
xnor U18036 (N_18036,N_15809,N_17224);
nand U18037 (N_18037,N_16424,N_15841);
xnor U18038 (N_18038,N_17403,N_17808);
or U18039 (N_18039,N_16742,N_16889);
nand U18040 (N_18040,N_17972,N_17267);
nor U18041 (N_18041,N_15745,N_16110);
or U18042 (N_18042,N_15555,N_16790);
nand U18043 (N_18043,N_17078,N_15232);
nor U18044 (N_18044,N_17662,N_15978);
nand U18045 (N_18045,N_17590,N_15976);
or U18046 (N_18046,N_15615,N_15317);
xnor U18047 (N_18047,N_17393,N_17346);
or U18048 (N_18048,N_17423,N_17124);
and U18049 (N_18049,N_15300,N_15396);
nor U18050 (N_18050,N_17179,N_17618);
nand U18051 (N_18051,N_15755,N_15207);
xor U18052 (N_18052,N_17080,N_15567);
or U18053 (N_18053,N_15401,N_16638);
nand U18054 (N_18054,N_16350,N_16890);
nor U18055 (N_18055,N_15492,N_16427);
or U18056 (N_18056,N_16582,N_16862);
nor U18057 (N_18057,N_16158,N_17190);
nand U18058 (N_18058,N_15891,N_15294);
and U18059 (N_18059,N_17593,N_16560);
and U18060 (N_18060,N_15698,N_16273);
and U18061 (N_18061,N_17572,N_16351);
or U18062 (N_18062,N_15487,N_15742);
nand U18063 (N_18063,N_15195,N_15919);
xor U18064 (N_18064,N_15551,N_17176);
or U18065 (N_18065,N_16398,N_17127);
and U18066 (N_18066,N_17141,N_15860);
xnor U18067 (N_18067,N_16010,N_15222);
and U18068 (N_18068,N_17717,N_16808);
nor U18069 (N_18069,N_17480,N_17299);
nor U18070 (N_18070,N_15547,N_15542);
and U18071 (N_18071,N_15554,N_16182);
xor U18072 (N_18072,N_16963,N_15906);
or U18073 (N_18073,N_16909,N_15849);
xor U18074 (N_18074,N_17390,N_15855);
nor U18075 (N_18075,N_15286,N_15172);
xor U18076 (N_18076,N_15691,N_16555);
and U18077 (N_18077,N_16167,N_16497);
or U18078 (N_18078,N_15356,N_16811);
nor U18079 (N_18079,N_16894,N_17362);
nand U18080 (N_18080,N_15751,N_16770);
nand U18081 (N_18081,N_17917,N_15921);
nand U18082 (N_18082,N_17880,N_15864);
nor U18083 (N_18083,N_17015,N_17115);
nor U18084 (N_18084,N_15139,N_17902);
xnor U18085 (N_18085,N_15832,N_15288);
or U18086 (N_18086,N_15955,N_17241);
xor U18087 (N_18087,N_15096,N_16702);
xor U18088 (N_18088,N_17690,N_15641);
xnor U18089 (N_18089,N_17007,N_16463);
xor U18090 (N_18090,N_16240,N_17057);
nand U18091 (N_18091,N_16141,N_15927);
or U18092 (N_18092,N_17746,N_15360);
nand U18093 (N_18093,N_16785,N_16195);
nor U18094 (N_18094,N_17231,N_17221);
or U18095 (N_18095,N_17077,N_15422);
xor U18096 (N_18096,N_15520,N_16198);
or U18097 (N_18097,N_17161,N_15722);
xor U18098 (N_18098,N_15406,N_15724);
and U18099 (N_18099,N_15901,N_15444);
nor U18100 (N_18100,N_15240,N_17488);
or U18101 (N_18101,N_17172,N_16651);
and U18102 (N_18102,N_15852,N_16342);
nand U18103 (N_18103,N_16052,N_16389);
nand U18104 (N_18104,N_16483,N_15163);
nor U18105 (N_18105,N_15024,N_16039);
and U18106 (N_18106,N_17610,N_17553);
xor U18107 (N_18107,N_16534,N_17722);
xor U18108 (N_18108,N_17806,N_17060);
xnor U18109 (N_18109,N_16715,N_15968);
nand U18110 (N_18110,N_15414,N_17277);
nand U18111 (N_18111,N_17298,N_16929);
and U18112 (N_18112,N_16054,N_15699);
nor U18113 (N_18113,N_16334,N_17276);
xor U18114 (N_18114,N_17058,N_15368);
xnor U18115 (N_18115,N_15078,N_17360);
and U18116 (N_18116,N_17912,N_17250);
xnor U18117 (N_18117,N_15201,N_15597);
or U18118 (N_18118,N_15256,N_15468);
nor U18119 (N_18119,N_17928,N_16938);
or U18120 (N_18120,N_16190,N_17351);
or U18121 (N_18121,N_17336,N_15452);
nor U18122 (N_18122,N_17048,N_15202);
and U18123 (N_18123,N_16896,N_17120);
nor U18124 (N_18124,N_15866,N_15223);
nand U18125 (N_18125,N_17434,N_16296);
xnor U18126 (N_18126,N_17929,N_16597);
nor U18127 (N_18127,N_17925,N_17409);
nor U18128 (N_18128,N_15051,N_16937);
xor U18129 (N_18129,N_17519,N_15609);
nor U18130 (N_18130,N_17159,N_17524);
nor U18131 (N_18131,N_15149,N_15788);
and U18132 (N_18132,N_16127,N_16876);
nand U18133 (N_18133,N_15090,N_16739);
or U18134 (N_18134,N_17897,N_17935);
nand U18135 (N_18135,N_17305,N_15416);
xor U18136 (N_18136,N_16936,N_17874);
or U18137 (N_18137,N_15244,N_15289);
nand U18138 (N_18138,N_17761,N_16913);
nor U18139 (N_18139,N_17122,N_15321);
nor U18140 (N_18140,N_15459,N_16466);
or U18141 (N_18141,N_17786,N_16769);
nor U18142 (N_18142,N_16053,N_17441);
or U18143 (N_18143,N_15226,N_15612);
or U18144 (N_18144,N_15228,N_15985);
xnor U18145 (N_18145,N_17338,N_17123);
or U18146 (N_18146,N_16418,N_15161);
xnor U18147 (N_18147,N_16679,N_17302);
or U18148 (N_18148,N_17232,N_15940);
nor U18149 (N_18149,N_15878,N_16917);
and U18150 (N_18150,N_16674,N_17967);
xnor U18151 (N_18151,N_16652,N_16532);
nor U18152 (N_18152,N_15266,N_15033);
and U18153 (N_18153,N_17713,N_15353);
xnor U18154 (N_18154,N_17566,N_17510);
or U18155 (N_18155,N_17879,N_16000);
or U18156 (N_18156,N_17333,N_15791);
and U18157 (N_18157,N_15009,N_16304);
nand U18158 (N_18158,N_16442,N_16412);
xor U18159 (N_18159,N_15141,N_17167);
nor U18160 (N_18160,N_17517,N_17832);
xnor U18161 (N_18161,N_15433,N_17429);
xor U18162 (N_18162,N_15050,N_16349);
nand U18163 (N_18163,N_15072,N_15524);
and U18164 (N_18164,N_15540,N_17865);
or U18165 (N_18165,N_16604,N_15227);
and U18166 (N_18166,N_17072,N_15405);
xor U18167 (N_18167,N_17777,N_17576);
and U18168 (N_18168,N_15109,N_16168);
nand U18169 (N_18169,N_15799,N_16206);
xor U18170 (N_18170,N_15498,N_16992);
nor U18171 (N_18171,N_15120,N_16043);
or U18172 (N_18172,N_16137,N_17960);
xnor U18173 (N_18173,N_16625,N_17317);
nor U18174 (N_18174,N_15596,N_16959);
and U18175 (N_18175,N_15086,N_16736);
and U18176 (N_18176,N_17392,N_17895);
and U18177 (N_18177,N_15477,N_16192);
nor U18178 (N_18178,N_17463,N_15404);
or U18179 (N_18179,N_17811,N_17814);
nor U18180 (N_18180,N_15510,N_16523);
and U18181 (N_18181,N_16869,N_16776);
nor U18182 (N_18182,N_15831,N_16209);
and U18183 (N_18183,N_17244,N_17182);
nand U18184 (N_18184,N_17582,N_16346);
or U18185 (N_18185,N_16121,N_15494);
and U18186 (N_18186,N_16289,N_17758);
nand U18187 (N_18187,N_17620,N_16512);
nor U18188 (N_18188,N_17196,N_17522);
xor U18189 (N_18189,N_15043,N_16612);
nor U18190 (N_18190,N_16145,N_16667);
or U18191 (N_18191,N_16672,N_15974);
nor U18192 (N_18192,N_15556,N_17165);
nand U18193 (N_18193,N_15638,N_16380);
or U18194 (N_18194,N_17813,N_15079);
nor U18195 (N_18195,N_16763,N_15795);
or U18196 (N_18196,N_16471,N_16336);
nand U18197 (N_18197,N_16149,N_17684);
nand U18198 (N_18198,N_15448,N_15601);
nor U18199 (N_18199,N_17860,N_17465);
or U18200 (N_18200,N_15100,N_17297);
or U18201 (N_18201,N_16552,N_17818);
xor U18202 (N_18202,N_17330,N_17347);
and U18203 (N_18203,N_16184,N_16975);
nand U18204 (N_18204,N_15943,N_16677);
and U18205 (N_18205,N_16060,N_17544);
and U18206 (N_18206,N_17263,N_17908);
nand U18207 (N_18207,N_16337,N_15177);
or U18208 (N_18208,N_15032,N_16269);
xor U18209 (N_18209,N_16096,N_16205);
or U18210 (N_18210,N_15663,N_16321);
nor U18211 (N_18211,N_17424,N_15165);
nor U18212 (N_18212,N_17410,N_15569);
and U18213 (N_18213,N_17552,N_16519);
and U18214 (N_18214,N_17686,N_17638);
nand U18215 (N_18215,N_17327,N_15765);
and U18216 (N_18216,N_15979,N_15390);
xnor U18217 (N_18217,N_16999,N_15187);
xor U18218 (N_18218,N_17111,N_15756);
and U18219 (N_18219,N_15284,N_17085);
and U18220 (N_18220,N_17676,N_16142);
nor U18221 (N_18221,N_15960,N_17567);
and U18222 (N_18222,N_15812,N_15140);
and U18223 (N_18223,N_17654,N_16001);
nor U18224 (N_18224,N_17926,N_15565);
and U18225 (N_18225,N_16341,N_15774);
xor U18226 (N_18226,N_15749,N_16958);
or U18227 (N_18227,N_16250,N_15453);
nor U18228 (N_18228,N_16684,N_15292);
xor U18229 (N_18229,N_16728,N_15215);
or U18230 (N_18230,N_16372,N_15903);
or U18231 (N_18231,N_16947,N_16177);
xnor U18232 (N_18232,N_17482,N_16690);
nor U18233 (N_18233,N_15212,N_17930);
or U18234 (N_18234,N_17872,N_15760);
or U18235 (N_18235,N_16095,N_16488);
or U18236 (N_18236,N_15330,N_15583);
or U18237 (N_18237,N_17851,N_17765);
xor U18238 (N_18238,N_17936,N_16792);
xor U18239 (N_18239,N_16017,N_15376);
or U18240 (N_18240,N_17665,N_15275);
xor U18241 (N_18241,N_17741,N_17841);
xnor U18242 (N_18242,N_16203,N_16226);
or U18243 (N_18243,N_17866,N_17720);
xor U18244 (N_18244,N_17822,N_17550);
nor U18245 (N_18245,N_15634,N_17303);
and U18246 (N_18246,N_15061,N_16038);
nand U18247 (N_18247,N_15265,N_16550);
nand U18248 (N_18248,N_17286,N_16824);
or U18249 (N_18249,N_17747,N_17599);
and U18250 (N_18250,N_17363,N_17331);
and U18251 (N_18251,N_15200,N_16375);
or U18252 (N_18252,N_17646,N_15074);
and U18253 (N_18253,N_17507,N_15006);
xnor U18254 (N_18254,N_16070,N_15683);
nor U18255 (N_18255,N_16924,N_17760);
nand U18256 (N_18256,N_15918,N_17442);
nor U18257 (N_18257,N_17024,N_16706);
xnor U18258 (N_18258,N_16018,N_16113);
xor U18259 (N_18259,N_16595,N_17460);
nor U18260 (N_18260,N_15123,N_15909);
or U18261 (N_18261,N_17495,N_16478);
nor U18262 (N_18262,N_16847,N_15216);
or U18263 (N_18263,N_17181,N_17364);
xnor U18264 (N_18264,N_17755,N_16707);
or U18265 (N_18265,N_17228,N_15470);
or U18266 (N_18266,N_15845,N_16084);
xor U18267 (N_18267,N_17933,N_16200);
nand U18268 (N_18268,N_17771,N_15714);
and U18269 (N_18269,N_15763,N_17177);
nor U18270 (N_18270,N_15382,N_16657);
nor U18271 (N_18271,N_16860,N_17361);
and U18272 (N_18272,N_17229,N_15121);
nor U18273 (N_18273,N_16546,N_16864);
nand U18274 (N_18274,N_17848,N_16535);
xnor U18275 (N_18275,N_15883,N_17382);
and U18276 (N_18276,N_17639,N_15311);
or U18277 (N_18277,N_15602,N_15824);
nand U18278 (N_18278,N_17581,N_16558);
nand U18279 (N_18279,N_17088,N_17957);
nor U18280 (N_18280,N_15594,N_15087);
and U18281 (N_18281,N_16248,N_17745);
and U18282 (N_18282,N_15528,N_16074);
xnor U18283 (N_18283,N_16571,N_16656);
or U18284 (N_18284,N_15944,N_17863);
xor U18285 (N_18285,N_16089,N_16368);
or U18286 (N_18286,N_15183,N_17201);
or U18287 (N_18287,N_17876,N_16883);
or U18288 (N_18288,N_15656,N_15859);
xnor U18289 (N_18289,N_15902,N_17752);
and U18290 (N_18290,N_16469,N_16099);
nand U18291 (N_18291,N_15255,N_15610);
xnor U18292 (N_18292,N_17262,N_16041);
or U18293 (N_18293,N_17595,N_17916);
or U18294 (N_18294,N_15920,N_16171);
and U18295 (N_18295,N_17574,N_15966);
or U18296 (N_18296,N_15060,N_17805);
xnor U18297 (N_18297,N_17032,N_15608);
or U18298 (N_18298,N_16157,N_17707);
xnor U18299 (N_18299,N_16888,N_17742);
xnor U18300 (N_18300,N_17559,N_15347);
xor U18301 (N_18301,N_17223,N_15996);
nor U18302 (N_18302,N_16034,N_16073);
xnor U18303 (N_18303,N_15213,N_17309);
nand U18304 (N_18304,N_16630,N_17809);
and U18305 (N_18305,N_17193,N_16735);
and U18306 (N_18306,N_15930,N_17738);
and U18307 (N_18307,N_15393,N_17171);
nand U18308 (N_18308,N_16576,N_15348);
nand U18309 (N_18309,N_17778,N_15178);
and U18310 (N_18310,N_17051,N_17207);
and U18311 (N_18311,N_17715,N_17973);
and U18312 (N_18312,N_17594,N_16697);
or U18313 (N_18313,N_17240,N_16379);
and U18314 (N_18314,N_15991,N_15616);
and U18315 (N_18315,N_17675,N_16570);
nor U18316 (N_18316,N_17473,N_16309);
nor U18317 (N_18317,N_16091,N_17425);
nor U18318 (N_18318,N_17601,N_15037);
or U18319 (N_18319,N_17970,N_15700);
nor U18320 (N_18320,N_17953,N_17197);
xnor U18321 (N_18321,N_16951,N_15913);
and U18322 (N_18322,N_17986,N_15890);
xor U18323 (N_18323,N_16646,N_17729);
nand U18324 (N_18324,N_17858,N_17401);
nor U18325 (N_18325,N_16082,N_17708);
nor U18326 (N_18326,N_17180,N_15999);
and U18327 (N_18327,N_16719,N_15900);
and U18328 (N_18328,N_16100,N_15243);
and U18329 (N_18329,N_17538,N_17107);
nand U18330 (N_18330,N_15426,N_16050);
or U18331 (N_18331,N_15512,N_15800);
xor U18332 (N_18332,N_17703,N_15154);
nand U18333 (N_18333,N_17353,N_17283);
xor U18334 (N_18334,N_17753,N_16968);
nor U18335 (N_18335,N_17527,N_17531);
or U18336 (N_18336,N_17896,N_16806);
and U18337 (N_18337,N_17468,N_15054);
xor U18338 (N_18338,N_15623,N_17047);
or U18339 (N_18339,N_17218,N_16631);
xor U18340 (N_18340,N_15075,N_17644);
or U18341 (N_18341,N_17561,N_17556);
and U18342 (N_18342,N_15108,N_15666);
nand U18343 (N_18343,N_16549,N_17640);
xnor U18344 (N_18344,N_15208,N_15062);
nand U18345 (N_18345,N_15118,N_16062);
nand U18346 (N_18346,N_17453,N_16148);
nor U18347 (N_18347,N_17609,N_16480);
nor U18348 (N_18348,N_15937,N_16536);
or U18349 (N_18349,N_16845,N_15392);
nand U18350 (N_18350,N_16985,N_17278);
nand U18351 (N_18351,N_16622,N_16830);
nor U18352 (N_18352,N_16542,N_17388);
nand U18353 (N_18353,N_16907,N_15586);
and U18354 (N_18354,N_16251,N_16102);
xor U18355 (N_18355,N_15709,N_15322);
nand U18356 (N_18356,N_17766,N_15785);
and U18357 (N_18357,N_17989,N_16670);
nor U18358 (N_18358,N_16044,N_15770);
and U18359 (N_18359,N_17154,N_16204);
nand U18360 (N_18360,N_17803,N_15533);
xor U18361 (N_18361,N_15296,N_16749);
nand U18362 (N_18362,N_15534,N_17189);
xnor U18363 (N_18363,N_17017,N_16283);
and U18364 (N_18364,N_15559,N_15325);
or U18365 (N_18365,N_15259,N_16780);
xor U18366 (N_18366,N_15989,N_17170);
nor U18367 (N_18367,N_15703,N_17018);
nand U18368 (N_18368,N_15914,N_17436);
xor U18369 (N_18369,N_16569,N_15097);
nor U18370 (N_18370,N_16410,N_15853);
and U18371 (N_18371,N_16333,N_16130);
nor U18372 (N_18372,N_17838,N_17526);
and U18373 (N_18373,N_17089,N_16843);
nand U18374 (N_18374,N_15950,N_16210);
and U18375 (N_18375,N_16014,N_16784);
xnor U18376 (N_18376,N_15112,N_15138);
xnor U18377 (N_18377,N_17118,N_17856);
or U18378 (N_18378,N_15245,N_15257);
and U18379 (N_18379,N_16281,N_17008);
or U18380 (N_18380,N_16948,N_15964);
nor U18381 (N_18381,N_16730,N_15478);
or U18382 (N_18382,N_16366,N_17090);
nand U18383 (N_18383,N_17270,N_15274);
or U18384 (N_18384,N_16880,N_15210);
or U18385 (N_18385,N_17615,N_16004);
and U18386 (N_18386,N_17097,N_17121);
nor U18387 (N_18387,N_15677,N_16691);
nor U18388 (N_18388,N_15354,N_15463);
xnor U18389 (N_18389,N_16152,N_15980);
or U18390 (N_18390,N_15219,N_17608);
or U18391 (N_18391,N_17381,N_15780);
or U18392 (N_18392,N_16923,N_17155);
xor U18393 (N_18393,N_16311,N_16867);
and U18394 (N_18394,N_17914,N_17312);
xor U18395 (N_18395,N_16766,N_17689);
and U18396 (N_18396,N_15184,N_16275);
and U18397 (N_18397,N_15735,N_17043);
or U18398 (N_18398,N_16545,N_16934);
nand U18399 (N_18399,N_17318,N_17021);
nor U18400 (N_18400,N_16188,N_15925);
or U18401 (N_18401,N_16729,N_16688);
nor U18402 (N_18402,N_16191,N_16287);
and U18403 (N_18403,N_16826,N_15643);
or U18404 (N_18404,N_17744,N_16821);
xor U18405 (N_18405,N_17990,N_16061);
or U18406 (N_18406,N_15005,N_17311);
and U18407 (N_18407,N_15142,N_15670);
nand U18408 (N_18408,N_16692,N_15496);
nand U18409 (N_18409,N_16288,N_17290);
nand U18410 (N_18410,N_17274,N_15590);
or U18411 (N_18411,N_17820,N_16957);
xor U18412 (N_18412,N_15821,N_17812);
nor U18413 (N_18413,N_15035,N_16922);
and U18414 (N_18414,N_16823,N_17178);
or U18415 (N_18415,N_17743,N_15797);
nor U18416 (N_18416,N_17625,N_17450);
and U18417 (N_18417,N_15664,N_15769);
nor U18418 (N_18418,N_15424,N_17762);
nor U18419 (N_18419,N_17963,N_17710);
or U18420 (N_18420,N_17259,N_16653);
and U18421 (N_18421,N_17328,N_16462);
nor U18422 (N_18422,N_17158,N_17040);
nor U18423 (N_18423,N_16915,N_17175);
nor U18424 (N_18424,N_15220,N_17621);
or U18425 (N_18425,N_15102,N_15829);
and U18426 (N_18426,N_15607,N_15803);
and U18427 (N_18427,N_15115,N_17281);
and U18428 (N_18428,N_15736,N_15897);
nand U18429 (N_18429,N_16978,N_15116);
nor U18430 (N_18430,N_16218,N_17310);
nor U18431 (N_18431,N_15151,N_17147);
nand U18432 (N_18432,N_16935,N_17092);
nand U18433 (N_18433,N_16954,N_15561);
or U18434 (N_18434,N_17604,N_15355);
or U18435 (N_18435,N_15907,N_15707);
and U18436 (N_18436,N_17308,N_17680);
or U18437 (N_18437,N_17651,N_17984);
nor U18438 (N_18438,N_17964,N_17073);
nand U18439 (N_18439,N_15268,N_15738);
and U18440 (N_18440,N_16639,N_16563);
and U18441 (N_18441,N_15372,N_16793);
xor U18442 (N_18442,N_15371,N_16698);
nand U18443 (N_18443,N_17248,N_16610);
or U18444 (N_18444,N_15467,N_15117);
or U18445 (N_18445,N_17801,N_16939);
nor U18446 (N_18446,N_15932,N_16768);
or U18447 (N_18447,N_16415,N_17988);
nor U18448 (N_18448,N_15378,N_17537);
or U18449 (N_18449,N_17135,N_15759);
nor U18450 (N_18450,N_15432,N_15816);
xnor U18451 (N_18451,N_15304,N_15145);
xor U18452 (N_18452,N_17408,N_17288);
or U18453 (N_18453,N_16263,N_16857);
xor U18454 (N_18454,N_15508,N_16352);
nor U18455 (N_18455,N_17864,N_15104);
nand U18456 (N_18456,N_16537,N_16391);
nand U18457 (N_18457,N_15858,N_15113);
nand U18458 (N_18458,N_16258,N_17455);
and U18459 (N_18459,N_15253,N_15085);
nand U18460 (N_18460,N_16249,N_16298);
or U18461 (N_18461,N_15928,N_16085);
xnor U18462 (N_18462,N_17013,N_15297);
and U18463 (N_18463,N_16506,N_15839);
nand U18464 (N_18464,N_16508,N_16165);
xnor U18465 (N_18465,N_16531,N_17104);
and U18466 (N_18466,N_15990,N_15495);
or U18467 (N_18467,N_16330,N_16755);
and U18468 (N_18468,N_17246,N_17899);
nor U18469 (N_18469,N_15877,N_17487);
nor U18470 (N_18470,N_16529,N_15538);
and U18471 (N_18471,N_17369,N_15209);
xor U18472 (N_18472,N_17046,N_16460);
and U18473 (N_18473,N_15513,N_16024);
nor U18474 (N_18474,N_15162,N_17975);
nand U18475 (N_18475,N_17323,N_16802);
nor U18476 (N_18476,N_15169,N_15680);
xor U18477 (N_18477,N_15553,N_15334);
xnor U18478 (N_18478,N_17406,N_17956);
nand U18479 (N_18479,N_16461,N_17705);
and U18480 (N_18480,N_15549,N_15229);
and U18481 (N_18481,N_17824,N_15341);
and U18482 (N_18482,N_17215,N_15970);
or U18483 (N_18483,N_16799,N_16107);
or U18484 (N_18484,N_15965,N_17448);
xnor U18485 (N_18485,N_15262,N_15929);
xor U18486 (N_18486,N_16694,N_15357);
nand U18487 (N_18487,N_15571,N_16429);
xnor U18488 (N_18488,N_17735,N_16406);
or U18489 (N_18489,N_15028,N_17284);
xnor U18490 (N_18490,N_15898,N_17205);
or U18491 (N_18491,N_17635,N_17560);
xnor U18492 (N_18492,N_15531,N_15580);
and U18493 (N_18493,N_16827,N_17113);
xor U18494 (N_18494,N_16919,N_15589);
xor U18495 (N_18495,N_15697,N_17920);
nor U18496 (N_18496,N_15572,N_17693);
xnor U18497 (N_18497,N_15904,N_15993);
nand U18498 (N_18498,N_15576,N_15499);
nor U18499 (N_18499,N_15713,N_17829);
xnor U18500 (N_18500,N_16164,N_16898);
and U18501 (N_18501,N_17422,N_16718);
xor U18502 (N_18502,N_15025,N_16960);
nand U18503 (N_18503,N_15817,N_15099);
or U18504 (N_18504,N_17139,N_16434);
nor U18505 (N_18505,N_15802,N_15715);
nand U18506 (N_18506,N_17130,N_15578);
nor U18507 (N_18507,N_16562,N_15048);
nor U18508 (N_18508,N_16435,N_17600);
or U18509 (N_18509,N_15529,N_16490);
xnor U18510 (N_18510,N_16910,N_17949);
xnor U18511 (N_18511,N_15777,N_17038);
and U18512 (N_18512,N_17993,N_16649);
nand U18513 (N_18513,N_17168,N_16282);
nand U18514 (N_18514,N_16431,N_17952);
nor U18515 (N_18515,N_15509,N_16155);
xor U18516 (N_18516,N_17066,N_17404);
or U18517 (N_18517,N_15389,N_17924);
nand U18518 (N_18518,N_16668,N_17358);
nor U18519 (N_18519,N_15194,N_15650);
nor U18520 (N_18520,N_15725,N_16405);
nand U18521 (N_18521,N_17669,N_17586);
xor U18522 (N_18522,N_16154,N_16838);
or U18523 (N_18523,N_16377,N_16274);
and U18524 (N_18524,N_15768,N_16186);
or U18525 (N_18525,N_16133,N_15339);
and U18526 (N_18526,N_15002,N_16411);
xor U18527 (N_18527,N_16637,N_15570);
nand U18528 (N_18528,N_16395,N_15316);
or U18529 (N_18529,N_16982,N_15279);
and U18530 (N_18530,N_17627,N_16795);
nor U18531 (N_18531,N_17208,N_15766);
nor U18532 (N_18532,N_15645,N_16176);
xor U18533 (N_18533,N_17850,N_15295);
and U18534 (N_18534,N_17557,N_17074);
or U18535 (N_18535,N_15176,N_16187);
nand U18536 (N_18536,N_17913,N_15310);
xor U18537 (N_18537,N_16605,N_15131);
xnor U18538 (N_18538,N_15862,N_17719);
nand U18539 (N_18539,N_17682,N_16773);
nor U18540 (N_18540,N_16814,N_16376);
and U18541 (N_18541,N_17691,N_15197);
nand U18542 (N_18542,N_15260,N_16738);
and U18543 (N_18543,N_15211,N_16733);
or U18544 (N_18544,N_15246,N_16547);
nand U18545 (N_18545,N_16884,N_17807);
nand U18546 (N_18546,N_17859,N_17109);
nand U18547 (N_18547,N_15977,N_16360);
nand U18548 (N_18548,N_15250,N_15536);
xor U18549 (N_18549,N_17452,N_17565);
and U18550 (N_18550,N_15704,N_17004);
xnor U18551 (N_18551,N_16172,N_16365);
xnor U18552 (N_18552,N_16608,N_16644);
and U18553 (N_18553,N_17134,N_16520);
xnor U18554 (N_18554,N_16930,N_16581);
and U18555 (N_18555,N_15899,N_16306);
nor U18556 (N_18556,N_15008,N_15367);
and U18557 (N_18557,N_16662,N_16477);
nand U18558 (N_18558,N_15026,N_17950);
or U18559 (N_18559,N_15427,N_16392);
nand U18560 (N_18560,N_15801,N_17444);
or U18561 (N_18561,N_16817,N_16362);
xor U18562 (N_18562,N_15894,N_16744);
or U18563 (N_18563,N_16385,N_17457);
xor U18564 (N_18564,N_16587,N_16627);
xor U18565 (N_18565,N_15204,N_17727);
and U18566 (N_18566,N_17998,N_16271);
xor U18567 (N_18567,N_15091,N_17343);
xnor U18568 (N_18568,N_15454,N_17030);
xor U18569 (N_18569,N_17905,N_17125);
xor U18570 (N_18570,N_15517,N_16144);
xnor U18571 (N_18571,N_16863,N_16789);
or U18572 (N_18572,N_17498,N_16993);
xnor U18573 (N_18573,N_17481,N_15484);
nand U18574 (N_18574,N_15397,N_16364);
and U18575 (N_18575,N_17010,N_17334);
nor U18576 (N_18576,N_16290,N_15375);
nand U18577 (N_18577,N_15464,N_15430);
xnor U18578 (N_18578,N_16804,N_16962);
xnor U18579 (N_18579,N_16032,N_17981);
or U18580 (N_18580,N_15254,N_17376);
or U18581 (N_18581,N_16498,N_17677);
nor U18582 (N_18582,N_17469,N_15474);
xnor U18583 (N_18583,N_17295,N_16063);
nand U18584 (N_18584,N_15481,N_17667);
nand U18585 (N_18585,N_16386,N_15038);
xnor U18586 (N_18586,N_16852,N_17633);
and U18587 (N_18587,N_16710,N_16714);
and U18588 (N_18588,N_16012,N_17339);
xnor U18589 (N_18589,N_16081,N_16783);
nor U18590 (N_18590,N_16021,N_16973);
and U18591 (N_18591,N_16800,N_15880);
or U18592 (N_18592,N_15055,N_15818);
nand U18593 (N_18593,N_15695,N_15125);
nand U18594 (N_18594,N_17551,N_15701);
nand U18595 (N_18595,N_16803,N_17245);
or U18596 (N_18596,N_17575,N_15535);
nand U18597 (N_18597,N_17187,N_15924);
xor U18598 (N_18598,N_17458,N_17796);
or U18599 (N_18599,N_17206,N_17792);
xnor U18600 (N_18600,N_17348,N_15543);
or U18601 (N_18601,N_17144,N_17937);
nand U18602 (N_18602,N_16829,N_17253);
nand U18603 (N_18603,N_16703,N_17878);
nor U18604 (N_18604,N_16327,N_17459);
xnor U18605 (N_18605,N_16556,N_15247);
nand U18606 (N_18606,N_17099,N_17294);
nor U18607 (N_18607,N_16874,N_16900);
nor U18608 (N_18608,N_17893,N_15566);
nand U18609 (N_18609,N_17623,N_16881);
nor U18610 (N_18610,N_17194,N_15122);
and U18611 (N_18611,N_15003,N_15873);
nand U18612 (N_18612,N_15385,N_15811);
nor U18613 (N_18613,N_17319,N_15483);
nor U18614 (N_18614,N_16227,N_16965);
or U18615 (N_18615,N_17505,N_17272);
nand U18616 (N_18616,N_17776,N_15633);
and U18617 (N_18617,N_15867,N_15486);
nor U18618 (N_18618,N_16443,N_16872);
nand U18619 (N_18619,N_17673,N_15719);
nor U18620 (N_18620,N_17462,N_15636);
and U18621 (N_18621,N_16199,N_16452);
xor U18622 (N_18622,N_17870,N_17543);
or U18623 (N_18623,N_15490,N_17374);
or U18624 (N_18624,N_16798,N_16578);
and U18625 (N_18625,N_17982,N_16426);
nor U18626 (N_18626,N_16717,N_16449);
xnor U18627 (N_18627,N_16318,N_17149);
xor U18628 (N_18628,N_17650,N_16640);
nor U18629 (N_18629,N_16378,N_16596);
and U18630 (N_18630,N_15447,N_16782);
or U18631 (N_18631,N_17923,N_16437);
xor U18632 (N_18632,N_17569,N_15190);
nor U18633 (N_18633,N_16276,N_17035);
nor U18634 (N_18634,N_17485,N_16116);
nand U18635 (N_18635,N_15711,N_16019);
and U18636 (N_18636,N_16680,N_15840);
xor U18637 (N_18637,N_17835,N_15599);
nor U18638 (N_18638,N_15331,N_16678);
xor U18639 (N_18639,N_15962,N_15741);
nor U18640 (N_18640,N_15935,N_17095);
xnor U18641 (N_18641,N_15624,N_15957);
nor U18642 (N_18642,N_17499,N_15539);
nor U18643 (N_18643,N_15063,N_15186);
nand U18644 (N_18644,N_15916,N_17721);
nor U18645 (N_18645,N_17324,N_15049);
and U18646 (N_18646,N_16256,N_16214);
nand U18647 (N_18647,N_16173,N_15473);
nand U18648 (N_18648,N_15750,N_17329);
xor U18649 (N_18649,N_15001,N_15748);
nor U18650 (N_18650,N_15861,N_17225);
and U18651 (N_18651,N_15865,N_15834);
nand U18652 (N_18652,N_15408,N_16538);
nand U18653 (N_18653,N_17653,N_16654);
and U18654 (N_18654,N_17587,N_17000);
nor U18655 (N_18655,N_16567,N_16465);
and U18656 (N_18656,N_17888,N_16945);
nor U18657 (N_18657,N_16745,N_17126);
nor U18658 (N_18658,N_15600,N_15754);
and U18659 (N_18659,N_16777,N_17414);
xnor U18660 (N_18660,N_16901,N_17054);
nand U18661 (N_18661,N_16601,N_15838);
nand U18662 (N_18662,N_16382,N_15198);
or U18663 (N_18663,N_17955,N_16925);
or U18664 (N_18664,N_17699,N_16179);
or U18665 (N_18665,N_17204,N_15655);
nand U18666 (N_18666,N_17849,N_16359);
or U18667 (N_18667,N_16075,N_15110);
xor U18668 (N_18668,N_17275,N_15130);
or U18669 (N_18669,N_17977,N_16967);
xor U18670 (N_18670,N_15874,N_17521);
nand U18671 (N_18671,N_15421,N_17211);
nand U18672 (N_18672,N_17022,N_17377);
nand U18673 (N_18673,N_15224,N_16583);
xnor U18674 (N_18674,N_17830,N_15548);
xnor U18675 (N_18675,N_16877,N_16231);
xor U18676 (N_18676,N_16485,N_15775);
nor U18677 (N_18677,N_17106,N_15628);
and U18678 (N_18678,N_17750,N_17887);
or U18679 (N_18679,N_15626,N_15042);
and U18680 (N_18680,N_15218,N_16517);
and U18681 (N_18681,N_15710,N_17475);
nand U18682 (N_18682,N_17968,N_15577);
and U18683 (N_18683,N_15733,N_15019);
nor U18684 (N_18684,N_15563,N_15587);
nor U18685 (N_18685,N_17921,N_15136);
nand U18686 (N_18686,N_17494,N_15456);
and U18687 (N_18687,N_17285,N_17002);
and U18688 (N_18688,N_15040,N_15439);
or U18689 (N_18689,N_15820,N_17940);
xor U18690 (N_18690,N_16305,N_15876);
and U18691 (N_18691,N_16400,N_16926);
xnor U18692 (N_18692,N_16354,N_16757);
or U18693 (N_18693,N_17020,N_15734);
nand U18694 (N_18694,N_15708,N_15205);
xor U18695 (N_18695,N_17663,N_16383);
xnor U18696 (N_18696,N_17428,N_17683);
nand U18697 (N_18697,N_16514,N_15269);
and U18698 (N_18698,N_16619,N_16457);
xor U18699 (N_18699,N_15155,N_15757);
xnor U18700 (N_18700,N_16740,N_16819);
nor U18701 (N_18701,N_15625,N_17611);
nor U18702 (N_18702,N_16634,N_17946);
nor U18703 (N_18703,N_15826,N_15252);
or U18704 (N_18704,N_17359,N_15689);
and U18705 (N_18705,N_17668,N_16373);
xnor U18706 (N_18706,N_17642,N_15942);
and U18707 (N_18707,N_15605,N_15409);
nor U18708 (N_18708,N_16067,N_15466);
nor U18709 (N_18709,N_16762,N_16722);
or U18710 (N_18710,N_15359,N_17780);
or U18711 (N_18711,N_16592,N_16201);
xnor U18712 (N_18712,N_16416,N_16300);
or U18713 (N_18713,N_17169,N_17315);
xor U18714 (N_18714,N_15661,N_16297);
or U18715 (N_18715,N_16510,N_15983);
or U18716 (N_18716,N_16139,N_16447);
nor U18717 (N_18717,N_17768,N_17589);
nand U18718 (N_18718,N_16430,N_15792);
nor U18719 (N_18719,N_16312,N_15667);
xnor U18720 (N_18720,N_15313,N_15654);
nor U18721 (N_18721,N_16574,N_17415);
nand U18722 (N_18722,N_17349,N_16059);
or U18723 (N_18723,N_16450,N_17724);
and U18724 (N_18724,N_16071,N_17129);
and U18725 (N_18725,N_17736,N_15248);
or U18726 (N_18726,N_16338,N_17260);
nor U18727 (N_18727,N_15217,N_17607);
xor U18728 (N_18728,N_16527,N_17700);
nor U18729 (N_18729,N_16006,N_15781);
xnor U18730 (N_18730,N_16642,N_15515);
or U18731 (N_18731,N_16588,N_15261);
or U18732 (N_18732,N_16202,N_17350);
nor U18733 (N_18733,N_15582,N_15758);
and U18734 (N_18734,N_15933,N_16262);
nor U18735 (N_18735,N_15997,N_15604);
nor U18736 (N_18736,N_15895,N_16245);
and U18737 (N_18737,N_15647,N_17235);
nor U18738 (N_18738,N_17230,N_15192);
xnor U18739 (N_18739,N_16976,N_17355);
nor U18740 (N_18740,N_15435,N_17588);
and U18741 (N_18741,N_16343,N_17026);
nand U18742 (N_18742,N_16147,N_15678);
and U18743 (N_18743,N_15181,N_17698);
xnor U18744 (N_18744,N_16586,N_15938);
or U18745 (N_18745,N_15391,N_16414);
nor U18746 (N_18746,N_16030,N_15568);
or U18747 (N_18747,N_16526,N_16150);
or U18748 (N_18748,N_17037,N_17366);
nand U18749 (N_18749,N_17539,N_17740);
nand U18750 (N_18750,N_17932,N_17597);
and U18751 (N_18751,N_16223,N_16833);
and U18752 (N_18752,N_17570,N_16685);
nand U18753 (N_18753,N_15794,N_17701);
xor U18754 (N_18754,N_16484,N_17542);
nor U18755 (N_18755,N_15762,N_15064);
and U18756 (N_18756,N_17289,N_15239);
and U18757 (N_18757,N_15098,N_16094);
nand U18758 (N_18758,N_17437,N_16225);
xor U18759 (N_18759,N_15241,N_17233);
nor U18760 (N_18760,N_16797,N_17300);
xnor U18761 (N_18761,N_17478,N_17951);
nor U18762 (N_18762,N_17630,N_16928);
xnor U18763 (N_18763,N_15819,N_15676);
nand U18764 (N_18764,N_17251,N_15737);
and U18765 (N_18765,N_17637,N_17657);
and U18766 (N_18766,N_15669,N_17445);
nor U18767 (N_18767,N_16384,N_16420);
nor U18768 (N_18768,N_15574,N_16720);
and U18769 (N_18769,N_16404,N_17877);
or U18770 (N_18770,N_17670,N_15830);
xor U18771 (N_18771,N_16241,N_17101);
and U18772 (N_18772,N_16990,N_17156);
and U18773 (N_18773,N_16682,N_17751);
xor U18774 (N_18774,N_17371,N_15868);
and U18775 (N_18775,N_16699,N_17027);
and U18776 (N_18776,N_15825,N_17476);
xnor U18777 (N_18777,N_17387,N_15303);
nand U18778 (N_18778,N_15995,N_15092);
and U18779 (N_18779,N_17426,N_16716);
nand U18780 (N_18780,N_17472,N_16325);
and U18781 (N_18781,N_17320,N_16079);
nor U18782 (N_18782,N_17810,N_17391);
or U18783 (N_18783,N_16319,N_16981);
nor U18784 (N_18784,N_16131,N_16988);
nand U18785 (N_18785,N_16228,N_15705);
and U18786 (N_18786,N_16551,N_16361);
xnor U18787 (N_18787,N_16303,N_17821);
xor U18788 (N_18788,N_16600,N_15501);
nor U18789 (N_18789,N_17939,N_17831);
nor U18790 (N_18790,N_17518,N_15752);
nand U18791 (N_18791,N_17352,N_16239);
nand U18792 (N_18792,N_16146,N_15946);
and U18793 (N_18793,N_15351,N_17540);
nand U18794 (N_18794,N_17432,N_15994);
and U18795 (N_18795,N_17728,N_15137);
and U18796 (N_18796,N_15363,N_17203);
nor U18797 (N_18797,N_15235,N_16669);
and U18798 (N_18798,N_15684,N_17103);
or U18799 (N_18799,N_15106,N_15236);
xor U18800 (N_18800,N_17198,N_17732);
or U18801 (N_18801,N_17834,N_17962);
or U18802 (N_18802,N_15617,N_16712);
nand U18803 (N_18803,N_15694,N_16242);
or U18804 (N_18804,N_15562,N_15693);
and U18805 (N_18805,N_15743,N_17029);
nor U18806 (N_18806,N_17282,N_15423);
xor U18807 (N_18807,N_16123,N_15462);
or U18808 (N_18808,N_15105,N_17915);
or U18809 (N_18809,N_16848,N_17764);
xor U18810 (N_18810,N_17596,N_17563);
xor U18811 (N_18811,N_16479,N_15127);
nand U18812 (N_18812,N_16835,N_16317);
nor U18813 (N_18813,N_15945,N_15067);
nor U18814 (N_18814,N_15744,N_17843);
nand U18815 (N_18815,N_15712,N_15731);
xnor U18816 (N_18816,N_16940,N_16841);
nor U18817 (N_18817,N_17733,N_15889);
nor U18818 (N_18818,N_17031,N_15394);
nor U18819 (N_18819,N_17116,N_17325);
nand U18820 (N_18820,N_16401,N_15308);
nor U18821 (N_18821,N_17692,N_17678);
and U18822 (N_18822,N_15682,N_15046);
xor U18823 (N_18823,N_15000,N_16128);
or U18824 (N_18824,N_16598,N_15281);
or U18825 (N_18825,N_16470,N_16161);
or U18826 (N_18826,N_17775,N_15129);
nand U18827 (N_18827,N_15383,N_15716);
and U18828 (N_18828,N_17449,N_16106);
and U18829 (N_18829,N_16388,N_16235);
or U18830 (N_18830,N_17784,N_17456);
nand U18831 (N_18831,N_16650,N_17273);
xor U18832 (N_18832,N_16774,N_16265);
nor U18833 (N_18833,N_16507,N_15998);
xnor U18834 (N_18834,N_15114,N_17628);
nand U18835 (N_18835,N_17999,N_17734);
nand U18836 (N_18836,N_15981,N_15635);
nor U18837 (N_18837,N_16513,N_17306);
xor U18838 (N_18838,N_16244,N_16068);
nor U18839 (N_18839,N_15639,N_15429);
xor U18840 (N_18840,N_16666,N_16895);
and U18841 (N_18841,N_16994,N_16613);
or U18842 (N_18842,N_17714,N_16875);
and U18843 (N_18843,N_16932,N_16611);
and U18844 (N_18844,N_17166,N_17005);
and U18845 (N_18845,N_15175,N_16849);
nand U18846 (N_18846,N_16760,N_15413);
nand U18847 (N_18847,N_16859,N_16181);
nand U18848 (N_18848,N_16476,N_15917);
nor U18849 (N_18849,N_15611,N_15657);
xnor U18850 (N_18850,N_17322,N_16897);
xnor U18851 (N_18851,N_16124,N_17344);
xnor U18852 (N_18852,N_16105,N_15352);
and U18853 (N_18853,N_16064,N_17909);
and U18854 (N_18854,N_17666,N_16246);
or U18855 (N_18855,N_15221,N_15338);
nand U18856 (N_18856,N_15789,N_17793);
and U18857 (N_18857,N_17602,N_15982);
and U18858 (N_18858,N_15640,N_15373);
or U18859 (N_18859,N_17484,N_15915);
and U18860 (N_18860,N_16232,N_15312);
or U18861 (N_18861,N_16101,N_17117);
xor U18862 (N_18862,N_16724,N_15975);
and U18863 (N_18863,N_17819,N_17407);
nand U18864 (N_18864,N_17997,N_17941);
and U18865 (N_18865,N_17247,N_16314);
or U18866 (N_18866,N_17430,N_16224);
nand U18867 (N_18867,N_16759,N_17649);
nor U18868 (N_18868,N_15761,N_16403);
or U18869 (N_18869,N_15144,N_16931);
or U18870 (N_18870,N_15786,N_15514);
xor U18871 (N_18871,N_15850,N_15199);
or U18872 (N_18872,N_16584,N_16454);
nor U18873 (N_18873,N_16455,N_15923);
or U18874 (N_18874,N_15337,N_15729);
nand U18875 (N_18875,N_17634,N_15521);
nand U18876 (N_18876,N_16340,N_16026);
or U18877 (N_18877,N_17405,N_15808);
or U18878 (N_18878,N_17656,N_17516);
or U18879 (N_18879,N_15431,N_15346);
xor U18880 (N_18880,N_17779,N_15896);
nand U18881 (N_18881,N_17548,N_17798);
nand U18882 (N_18882,N_16291,N_17739);
or U18883 (N_18883,N_16659,N_17862);
or U18884 (N_18884,N_16115,N_16093);
or U18885 (N_18885,N_16624,N_17316);
or U18886 (N_18886,N_17783,N_15546);
or U18887 (N_18887,N_17291,N_16260);
and U18888 (N_18888,N_16820,N_16647);
nand U18889 (N_18889,N_15362,N_15893);
and U18890 (N_18890,N_16916,N_17136);
xnor U18891 (N_18891,N_17056,N_16956);
xor U18892 (N_18892,N_15364,N_15076);
nand U18893 (N_18893,N_15084,N_16704);
xnor U18894 (N_18894,N_15306,N_17184);
nand U18895 (N_18895,N_17658,N_15012);
xor U18896 (N_18896,N_16886,N_17304);
or U18897 (N_18897,N_16329,N_17571);
nor U18898 (N_18898,N_15807,N_17420);
and U18899 (N_18899,N_17534,N_17471);
and U18900 (N_18900,N_16914,N_17183);
nor U18901 (N_18901,N_17791,N_15333);
nand U18902 (N_18902,N_15905,N_17398);
and U18903 (N_18903,N_17337,N_16013);
nand U18904 (N_18904,N_16015,N_16217);
or U18905 (N_18905,N_17884,N_15022);
and U18906 (N_18906,N_15119,N_17696);
and U18907 (N_18907,N_17500,N_17082);
nor U18908 (N_18908,N_16140,N_17643);
nor U18909 (N_18909,N_16502,N_16153);
or U18910 (N_18910,N_17969,N_16393);
nand U18911 (N_18911,N_17617,N_17023);
xnor U18912 (N_18912,N_17164,N_15967);
xor U18913 (N_18913,N_15646,N_17143);
xnor U18914 (N_18914,N_16593,N_16892);
xor U18915 (N_18915,N_17520,N_17655);
nor U18916 (N_18916,N_17059,N_16801);
nand U18917 (N_18917,N_15171,N_17787);
and U18918 (N_18918,N_16899,N_17261);
nand U18919 (N_18919,N_16156,N_17857);
xnor U18920 (N_18920,N_15835,N_15147);
or U18921 (N_18921,N_16681,N_16861);
or U18922 (N_18922,N_15280,N_16687);
or U18923 (N_18923,N_16125,N_17399);
or U18924 (N_18924,N_17264,N_15558);
and U18925 (N_18925,N_15591,N_16663);
nand U18926 (N_18926,N_16035,N_16363);
nor U18927 (N_18927,N_17191,N_15560);
xnor U18928 (N_18928,N_15101,N_17502);
or U18929 (N_18929,N_15148,N_15164);
nand U18930 (N_18930,N_17688,N_15776);
nor U18931 (N_18931,N_17493,N_15659);
and U18932 (N_18932,N_15649,N_17222);
nor U18933 (N_18933,N_15167,N_15692);
and U18934 (N_18934,N_17142,N_16222);
xnor U18935 (N_18935,N_16423,N_17062);
xnor U18936 (N_18936,N_17528,N_16525);
nor U18937 (N_18937,N_17174,N_17898);
nor U18938 (N_18938,N_15771,N_15343);
xor U18939 (N_18939,N_15395,N_16511);
xnor U18940 (N_18940,N_16174,N_16065);
xor U18941 (N_18941,N_15193,N_17825);
xnor U18942 (N_18942,N_16891,N_17055);
and U18943 (N_18943,N_17846,N_15277);
or U18944 (N_18944,N_15126,N_16844);
or U18945 (N_18945,N_16007,N_17983);
nor U18946 (N_18946,N_15159,N_17012);
nand U18947 (N_18947,N_17712,N_16169);
or U18948 (N_18948,N_16208,N_16104);
or U18949 (N_18949,N_15476,N_16175);
nand U18950 (N_18950,N_16772,N_15675);
xnor U18951 (N_18951,N_17354,N_16278);
xor U18952 (N_18952,N_15027,N_16557);
xnor U18953 (N_18953,N_17036,N_16098);
nand U18954 (N_18954,N_17852,N_16645);
nand U18955 (N_18955,N_17942,N_15238);
nor U18956 (N_18956,N_16229,N_15095);
and U18957 (N_18957,N_17087,N_15717);
or U18958 (N_18958,N_17292,N_16501);
or U18959 (N_18959,N_17647,N_16464);
xnor U18960 (N_18960,N_16815,N_17451);
and U18961 (N_18961,N_17332,N_16286);
xor U18962 (N_18962,N_16396,N_16989);
xnor U18963 (N_18963,N_15953,N_15941);
nand U18964 (N_18964,N_17959,N_16197);
xnor U18965 (N_18965,N_16323,N_15637);
and U18966 (N_18966,N_15282,N_17716);
and U18967 (N_18967,N_17071,N_15166);
or U18968 (N_18968,N_16216,N_15488);
and U18969 (N_18969,N_17001,N_17861);
xnor U18970 (N_18970,N_16591,N_15366);
nor U18971 (N_18971,N_17385,N_17365);
and U18972 (N_18972,N_16402,N_15593);
and U18973 (N_18973,N_15598,N_15047);
nor U18974 (N_18974,N_15482,N_17379);
nor U18975 (N_18975,N_15124,N_17961);
nor U18976 (N_18976,N_17794,N_17974);
or U18977 (N_18977,N_16045,N_16887);
or U18978 (N_18978,N_17947,N_15315);
xor U18979 (N_18979,N_16238,N_16446);
nor U18980 (N_18980,N_16746,N_17386);
nor U18981 (N_18981,N_17137,N_17938);
or U18982 (N_18982,N_17945,N_16310);
or U18983 (N_18983,N_15530,N_15278);
or U18984 (N_18984,N_15020,N_17427);
nand U18985 (N_18985,N_17695,N_17239);
or U18986 (N_18986,N_16564,N_16408);
or U18987 (N_18987,N_16135,N_15044);
nand U18988 (N_18988,N_15497,N_15089);
nor U18989 (N_18989,N_16301,N_16440);
or U18990 (N_18990,N_15685,N_16660);
nor U18991 (N_18991,N_17053,N_17530);
xor U18992 (N_18992,N_17533,N_16308);
xor U18993 (N_18993,N_15233,N_15237);
nor U18994 (N_18994,N_16675,N_15922);
and U18995 (N_18995,N_16002,N_15952);
or U18996 (N_18996,N_16328,N_15107);
nor U18997 (N_18997,N_15882,N_16996);
and U18998 (N_18998,N_15973,N_17867);
or U18999 (N_18999,N_16335,N_15778);
nand U19000 (N_19000,N_17257,N_15143);
and U19001 (N_19001,N_16138,N_15815);
nand U19002 (N_19002,N_15892,N_16565);
xnor U19003 (N_19003,N_16451,N_16834);
nor U19004 (N_19004,N_16737,N_16966);
and U19005 (N_19005,N_17202,N_16230);
nor U19006 (N_19006,N_16347,N_15081);
nor U19007 (N_19007,N_16467,N_15537);
nor U19008 (N_19008,N_15017,N_16129);
or U19009 (N_19009,N_16585,N_15805);
and U19010 (N_19010,N_17767,N_15671);
xor U19011 (N_19011,N_15450,N_17357);
xnor U19012 (N_19012,N_16163,N_16009);
xnor U19013 (N_19013,N_15672,N_16264);
nor U19014 (N_19014,N_17562,N_17948);
nor U19015 (N_19015,N_16355,N_16616);
nor U19016 (N_19016,N_16055,N_16953);
nand U19017 (N_19017,N_15336,N_17979);
xor U19018 (N_19018,N_16280,N_15440);
or U19019 (N_19019,N_17367,N_15326);
nand U19020 (N_19020,N_15690,N_17070);
nor U19021 (N_19021,N_17723,N_17496);
or U19022 (N_19022,N_17614,N_16655);
nand U19023 (N_19023,N_15088,N_16294);
xnor U19024 (N_19024,N_15706,N_17067);
and U19025 (N_19025,N_15485,N_15093);
nand U19026 (N_19026,N_17679,N_16912);
nand U19027 (N_19027,N_15302,N_17873);
and U19028 (N_19028,N_16635,N_17991);
and U19029 (N_19029,N_16357,N_16761);
nand U19030 (N_19030,N_17546,N_15272);
xnor U19031 (N_19031,N_17605,N_16528);
nor U19032 (N_19032,N_16458,N_17076);
or U19033 (N_19033,N_15045,N_16077);
and U19034 (N_19034,N_17828,N_17785);
xnor U19035 (N_19035,N_17254,N_16548);
xor U19036 (N_19036,N_15505,N_16850);
or U19037 (N_19037,N_16734,N_17236);
or U19038 (N_19038,N_16033,N_16522);
and U19039 (N_19039,N_15844,N_17906);
or U19040 (N_19040,N_17509,N_16721);
nand U19041 (N_19041,N_15258,N_15739);
nand U19042 (N_19042,N_16908,N_16732);
nor U19043 (N_19043,N_17006,N_16221);
xnor U19044 (N_19044,N_17064,N_16609);
nand U19045 (N_19045,N_17033,N_16832);
and U19046 (N_19046,N_16521,N_16031);
xor U19047 (N_19047,N_16178,N_15828);
or U19048 (N_19048,N_16998,N_15065);
or U19049 (N_19049,N_16213,N_16983);
or U19050 (N_19050,N_17894,N_17108);
and U19051 (N_19051,N_15936,N_17397);
and U19052 (N_19052,N_17173,N_17592);
or U19053 (N_19053,N_15827,N_17826);
or U19054 (N_19054,N_15992,N_17380);
nor U19055 (N_19055,N_16846,N_15073);
xor U19056 (N_19056,N_15374,N_16905);
nor U19057 (N_19057,N_16432,N_16858);
or U19058 (N_19058,N_16295,N_17718);
nand U19059 (N_19059,N_15379,N_17645);
and U19060 (N_19060,N_16371,N_16756);
and U19061 (N_19061,N_15415,N_15783);
nor U19062 (N_19062,N_15400,N_17891);
and U19063 (N_19063,N_17326,N_17466);
or U19064 (N_19064,N_15158,N_15327);
nand U19065 (N_19065,N_16166,N_17492);
xor U19066 (N_19066,N_16080,N_16233);
nor U19067 (N_19067,N_15290,N_17816);
and U19068 (N_19068,N_15822,N_16589);
nand U19069 (N_19069,N_17162,N_15299);
or U19070 (N_19070,N_15014,N_15287);
or U19071 (N_19071,N_15793,N_15443);
and U19072 (N_19072,N_17966,N_15361);
xnor U19073 (N_19073,N_15584,N_16132);
nand U19074 (N_19074,N_15370,N_16279);
xor U19075 (N_19075,N_17711,N_16428);
xor U19076 (N_19076,N_16344,N_16247);
nor U19077 (N_19077,N_15502,N_15631);
nand U19078 (N_19078,N_16051,N_15173);
xor U19079 (N_19079,N_16495,N_15058);
xnor U19080 (N_19080,N_16473,N_15234);
nand U19081 (N_19081,N_16487,N_15545);
or U19082 (N_19082,N_15445,N_17212);
nand U19083 (N_19083,N_16920,N_17084);
and U19084 (N_19084,N_15782,N_16316);
or U19085 (N_19085,N_15681,N_16903);
and U19086 (N_19086,N_15493,N_15688);
or U19087 (N_19087,N_16439,N_17697);
or U19088 (N_19088,N_15912,N_15412);
nand U19089 (N_19089,N_17335,N_16568);
and U19090 (N_19090,N_16628,N_15156);
nand U19091 (N_19091,N_15622,N_15934);
and U19092 (N_19092,N_15947,N_17146);
and U19093 (N_19093,N_15015,N_15779);
nand U19094 (N_19094,N_15350,N_17800);
nand U19095 (N_19095,N_16367,N_16087);
nand U19096 (N_19096,N_17886,N_15323);
nor U19097 (N_19097,N_15856,N_16658);
xor U19098 (N_19098,N_16056,N_15814);
or U19099 (N_19099,N_17868,N_16285);
and U19100 (N_19100,N_17370,N_17413);
nand U19101 (N_19101,N_15810,N_15931);
nor U19102 (N_19102,N_15887,N_15564);
or U19103 (N_19103,N_17624,N_16904);
xnor U19104 (N_19104,N_15455,N_15251);
or U19105 (N_19105,N_15291,N_15083);
nand U19106 (N_19106,N_16765,N_17501);
xnor U19107 (N_19107,N_15573,N_17631);
or U19108 (N_19108,N_16072,N_16796);
or U19109 (N_19109,N_15674,N_16969);
xnor U19110 (N_19110,N_15956,N_16831);
nand U19111 (N_19111,N_16324,N_17549);
nand U19112 (N_19112,N_16170,N_17474);
or U19113 (N_19113,N_15658,N_15740);
or U19114 (N_19114,N_16805,N_16991);
xor U19115 (N_19115,N_16865,N_15029);
xnor U19116 (N_19116,N_17844,N_17242);
nand U19117 (N_19117,N_15225,N_17226);
and U19118 (N_19118,N_17612,N_16407);
or U19119 (N_19119,N_16088,N_15465);
xnor U19120 (N_19120,N_15335,N_15094);
nor U19121 (N_19121,N_15442,N_15871);
and U19122 (N_19122,N_15851,N_15388);
and U19123 (N_19123,N_15526,N_17558);
nand U19124 (N_19124,N_17186,N_15951);
xnor U19125 (N_19125,N_17209,N_16836);
or U19126 (N_19126,N_15642,N_17028);
and U19127 (N_19127,N_16603,N_15753);
and U19128 (N_19128,N_16058,N_15857);
nand U19129 (N_19129,N_15673,N_15320);
or U19130 (N_19130,N_17439,N_17470);
nor U19131 (N_19131,N_15527,N_17447);
and U19132 (N_19132,N_17789,N_15911);
and U19133 (N_19133,N_16111,N_15702);
and U19134 (N_19134,N_17252,N_16016);
and U19135 (N_19135,N_16302,N_16623);
and U19136 (N_19136,N_16573,N_16828);
or U19137 (N_19137,N_15182,N_15369);
nor U19138 (N_19138,N_16870,N_15804);
xnor U19139 (N_19139,N_15848,N_17394);
or U19140 (N_19140,N_15939,N_16353);
nor U19141 (N_19141,N_16066,N_16499);
nor U19142 (N_19142,N_15263,N_15180);
or U19143 (N_19143,N_16036,N_15271);
nand U19144 (N_19144,N_16486,N_16902);
nor U19145 (N_19145,N_15847,N_16307);
xnor U19146 (N_19146,N_16599,N_16448);
and U19147 (N_19147,N_16661,N_15620);
and U19148 (N_19148,N_16322,N_15319);
and U19149 (N_19149,N_15128,N_16750);
nand U19150 (N_19150,N_17402,N_16022);
nor U19151 (N_19151,N_17837,N_15987);
nand U19152 (N_19152,N_17373,N_16553);
nor U19153 (N_19153,N_17616,N_16995);
or U19154 (N_19154,N_17603,N_17790);
or U19155 (N_19155,N_17145,N_17555);
and U19156 (N_19156,N_16533,N_16234);
nor U19157 (N_19157,N_16489,N_16313);
nor U19158 (N_19158,N_16693,N_16261);
xor U19159 (N_19159,N_16397,N_17591);
or U19160 (N_19160,N_15489,N_17815);
nor U19161 (N_19161,N_17079,N_17412);
nor U19162 (N_19162,N_16607,N_17613);
and U19163 (N_19163,N_17769,N_17131);
nor U19164 (N_19164,N_15196,N_15721);
or U19165 (N_19165,N_17195,N_17889);
and U19166 (N_19166,N_17314,N_17773);
and U19167 (N_19167,N_17788,N_16577);
xor U19168 (N_19168,N_15652,N_17454);
nand U19169 (N_19169,N_15031,N_17985);
xnor U19170 (N_19170,N_15653,N_17797);
and U19171 (N_19171,N_15071,N_16842);
and U19172 (N_19172,N_15457,N_17577);
and U19173 (N_19173,N_16083,N_17063);
nor U19174 (N_19174,N_16057,N_15723);
nor U19175 (N_19175,N_17980,N_17772);
nor U19176 (N_19176,N_15030,N_16705);
nand U19177 (N_19177,N_15231,N_15399);
nor U19178 (N_19178,N_17157,N_15541);
and U19179 (N_19179,N_16425,N_16758);
nand U19180 (N_19180,N_17681,N_15057);
nand U19181 (N_19181,N_17307,N_17188);
nand U19182 (N_19182,N_17083,N_17265);
xnor U19183 (N_19183,N_15614,N_17491);
nor U19184 (N_19184,N_17378,N_17995);
nand U19185 (N_19185,N_17598,N_17395);
nand U19186 (N_19186,N_17152,N_15613);
and U19187 (N_19187,N_17467,N_15410);
nand U19188 (N_19188,N_16253,N_15011);
nor U19189 (N_19189,N_17903,N_15080);
and U19190 (N_19190,N_16708,N_15627);
and U19191 (N_19191,N_15214,N_16180);
xnor U19192 (N_19192,N_15948,N_15230);
and U19193 (N_19193,N_16851,N_15686);
nand U19194 (N_19194,N_17554,N_16787);
nand U19195 (N_19195,N_16413,N_15842);
or U19196 (N_19196,N_15479,N_15507);
and U19197 (N_19197,N_16472,N_15550);
and U19198 (N_19198,N_15384,N_16807);
xor U19199 (N_19199,N_17050,N_15013);
nor U19200 (N_19200,N_17098,N_16284);
or U19201 (N_19201,N_17419,N_16906);
and U19202 (N_19202,N_16524,N_17140);
and U19203 (N_19203,N_15726,N_15679);
nand U19204 (N_19204,N_16977,N_17944);
and U19205 (N_19205,N_16117,N_16580);
nor U19206 (N_19206,N_17535,N_16541);
and U19207 (N_19207,N_17258,N_17034);
nand U19208 (N_19208,N_17573,N_15519);
nand U19209 (N_19209,N_17513,N_17431);
or U19210 (N_19210,N_16369,N_17287);
xnor U19211 (N_19211,N_16504,N_15034);
or U19212 (N_19212,N_17836,N_17014);
or U19213 (N_19213,N_16122,N_17910);
or U19214 (N_19214,N_16711,N_16259);
nand U19215 (N_19215,N_17749,N_17704);
nand U19216 (N_19216,N_16971,N_15157);
nand U19217 (N_19217,N_16212,N_15503);
nor U19218 (N_19218,N_17255,N_16387);
or U19219 (N_19219,N_16097,N_17266);
or U19220 (N_19220,N_17971,N_15772);
nand U19221 (N_19221,N_16731,N_15053);
nand U19222 (N_19222,N_15314,N_15836);
or U19223 (N_19223,N_16855,N_16332);
and U19224 (N_19224,N_17091,N_15506);
and U19225 (N_19225,N_16620,N_16118);
xnor U19226 (N_19226,N_17685,N_17606);
nor U19227 (N_19227,N_17296,N_16381);
or U19228 (N_19228,N_16813,N_16885);
nand U19229 (N_19229,N_17268,N_17508);
nand U19230 (N_19230,N_17238,N_16160);
and U19231 (N_19231,N_16812,N_17375);
or U19232 (N_19232,N_16539,N_16003);
and U19233 (N_19233,N_16109,N_17199);
or U19234 (N_19234,N_15746,N_17847);
and U19235 (N_19235,N_15767,N_16840);
and U19236 (N_19236,N_15285,N_15342);
and U19237 (N_19237,N_17435,N_17855);
and U19238 (N_19238,N_16492,N_15954);
nand U19239 (N_19239,N_17045,N_15134);
nor U19240 (N_19240,N_16193,N_17626);
nand U19241 (N_19241,N_17341,N_16664);
nand U19242 (N_19242,N_16331,N_16509);
nand U19243 (N_19243,N_15773,N_17632);
nand U19244 (N_19244,N_16069,N_16543);
and U19245 (N_19245,N_15972,N_17515);
and U19246 (N_19246,N_15016,N_15380);
nor U19247 (N_19247,N_16615,N_15813);
or U19248 (N_19248,N_16856,N_16326);
nand U19249 (N_19249,N_15242,N_16194);
or U19250 (N_19250,N_15875,N_16348);
or U19251 (N_19251,N_16871,N_17965);
and U19252 (N_19252,N_15276,N_15068);
nor U19253 (N_19253,N_15153,N_15511);
and U19254 (N_19254,N_16854,N_17804);
nor U19255 (N_19255,N_16701,N_17583);
nor U19256 (N_19256,N_17904,N_15843);
or U19257 (N_19257,N_16636,N_16530);
nand U19258 (N_19258,N_15798,N_16911);
and U19259 (N_19259,N_16540,N_15472);
or U19260 (N_19260,N_15328,N_17128);
nor U19261 (N_19261,N_15249,N_17433);
xor U19262 (N_19262,N_16162,N_15575);
or U19263 (N_19263,N_17875,N_17464);
nor U19264 (N_19264,N_17996,N_17823);
nand U19265 (N_19265,N_16944,N_15344);
nor U19266 (N_19266,N_17417,N_17853);
nor U19267 (N_19267,N_17486,N_17368);
xnor U19268 (N_19268,N_16879,N_16723);
and U19269 (N_19269,N_15619,N_17049);
and U19270 (N_19270,N_16868,N_15386);
and U19271 (N_19271,N_17578,N_16254);
or U19272 (N_19272,N_17795,N_17536);
nand U19273 (N_19273,N_17664,N_17781);
nand U19274 (N_19274,N_16980,N_16559);
nand U19275 (N_19275,N_15307,N_16134);
xnor U19276 (N_19276,N_16516,N_16853);
or U19277 (N_19277,N_15039,N_15881);
or U19278 (N_19278,N_16837,N_15437);
xnor U19279 (N_19279,N_16185,N_16788);
nor U19280 (N_19280,N_15888,N_17629);
nand U19281 (N_19281,N_15418,N_16572);
nor U19282 (N_19282,N_17081,N_15632);
or U19283 (N_19283,N_15133,N_15417);
xor U19284 (N_19284,N_16786,N_16809);
nand U19285 (N_19285,N_17132,N_17737);
or U19286 (N_19286,N_17514,N_16474);
or U19287 (N_19287,N_15588,N_16695);
or U19288 (N_19288,N_16503,N_17384);
xnor U19289 (N_19289,N_16267,N_15082);
or U19290 (N_19290,N_17102,N_15428);
nand U19291 (N_19291,N_15651,N_16046);
nor U19292 (N_19292,N_17210,N_16987);
nor U19293 (N_19293,N_17901,N_16779);
and U19294 (N_19294,N_15441,N_17086);
xor U19295 (N_19295,N_16544,N_17892);
or U19296 (N_19296,N_16676,N_15958);
or U19297 (N_19297,N_17882,N_17497);
nand U19298 (N_19298,N_15434,N_15784);
and U19299 (N_19299,N_16747,N_15581);
nand U19300 (N_19300,N_17249,N_16882);
nor U19301 (N_19301,N_17400,N_16494);
nand U19302 (N_19302,N_15069,N_16108);
nor U19303 (N_19303,N_17011,N_16339);
nor U19304 (N_19304,N_16626,N_15630);
and U19305 (N_19305,N_17052,N_15056);
nand U19306 (N_19306,N_16825,N_15696);
and U19307 (N_19307,N_16921,N_15884);
or U19308 (N_19308,N_17490,N_16103);
and U19309 (N_19309,N_15021,N_16614);
xnor U19310 (N_19310,N_16048,N_16942);
or U19311 (N_19311,N_15309,N_15324);
xnor U19312 (N_19312,N_17105,N_15036);
xor U19313 (N_19313,N_16025,N_17110);
and U19314 (N_19314,N_15010,N_15345);
or U19315 (N_19315,N_16590,N_16893);
nand U19316 (N_19316,N_17280,N_15425);
or U19317 (N_19317,N_16293,N_16092);
or U19318 (N_19318,N_15869,N_17911);
xor U19319 (N_19319,N_17525,N_17918);
xnor U19320 (N_19320,N_16775,N_16292);
nand U19321 (N_19321,N_15621,N_17383);
or U19322 (N_19322,N_15500,N_15665);
or U19323 (N_19323,N_17313,N_15365);
or U19324 (N_19324,N_17842,N_15518);
and U19325 (N_19325,N_16816,N_16207);
nand U19326 (N_19326,N_16500,N_15066);
nand U19327 (N_19327,N_15718,N_15206);
and U19328 (N_19328,N_16818,N_17041);
nand U19329 (N_19329,N_17321,N_17342);
xor U19330 (N_19330,N_17214,N_15522);
xor U19331 (N_19331,N_16315,N_15491);
or U19332 (N_19332,N_17641,N_16700);
or U19333 (N_19333,N_16023,N_15052);
and U19334 (N_19334,N_17416,N_17706);
nand U19335 (N_19335,N_17674,N_15267);
xnor U19336 (N_19336,N_17726,N_17133);
or U19337 (N_19337,N_16243,N_17730);
or U19338 (N_19338,N_15387,N_16949);
and U19339 (N_19339,N_17845,N_16028);
and U19340 (N_19340,N_17770,N_17523);
nor U19341 (N_19341,N_15971,N_16211);
or U19342 (N_19342,N_16444,N_16689);
xor U19343 (N_19343,N_16726,N_15160);
nand U19344 (N_19344,N_15959,N_15552);
xnor U19345 (N_19345,N_17636,N_15420);
nor U19346 (N_19346,N_15595,N_16236);
nand U19347 (N_19347,N_16778,N_16409);
nor U19348 (N_19348,N_16771,N_17396);
xnor U19349 (N_19349,N_15146,N_17418);
and U19350 (N_19350,N_17709,N_16665);
or U19351 (N_19351,N_16873,N_15969);
xor U19352 (N_19352,N_15984,N_17661);
or U19353 (N_19353,N_16417,N_16078);
and U19354 (N_19354,N_15174,N_17900);
nor U19355 (N_19355,N_16266,N_17479);
xor U19356 (N_19356,N_16374,N_16950);
xnor U19357 (N_19357,N_17672,N_17044);
and U19358 (N_19358,N_17075,N_16037);
or U19359 (N_19359,N_15018,N_15796);
nand U19360 (N_19360,N_17100,N_17547);
or U19361 (N_19361,N_16272,N_16791);
nand U19362 (N_19362,N_16579,N_16629);
and U19363 (N_19363,N_17839,N_17883);
nand U19364 (N_19364,N_17237,N_16839);
nand U19365 (N_19365,N_16086,N_16299);
and U19366 (N_19366,N_16120,N_17438);
nand U19367 (N_19367,N_16020,N_16237);
nand U19368 (N_19368,N_15438,N_16979);
or U19369 (N_19369,N_16126,N_17345);
and U19370 (N_19370,N_17541,N_15451);
xor U19371 (N_19371,N_17185,N_15381);
xnor U19372 (N_19372,N_17293,N_16866);
nor U19373 (N_19373,N_16696,N_17799);
nor U19374 (N_19374,N_17069,N_15449);
nor U19375 (N_19375,N_15041,N_15806);
xor U19376 (N_19376,N_15730,N_17564);
xnor U19377 (N_19377,N_15629,N_15790);
nand U19378 (N_19378,N_15648,N_16781);
xor U19379 (N_19379,N_17150,N_17652);
nor U19380 (N_19380,N_17093,N_15846);
and U19381 (N_19381,N_17477,N_16219);
nor U19382 (N_19382,N_17774,N_15525);
xor U19383 (N_19383,N_15301,N_15603);
xnor U19384 (N_19384,N_17213,N_15879);
or U19385 (N_19385,N_17096,N_15340);
nor U19386 (N_19386,N_15298,N_17919);
or U19387 (N_19387,N_15332,N_15854);
xor U19388 (N_19388,N_17748,N_15949);
nor U19389 (N_19389,N_16713,N_16810);
nand U19390 (N_19390,N_15475,N_17068);
or U19391 (N_19391,N_17922,N_15436);
and U19392 (N_19392,N_15833,N_16441);
nand U19393 (N_19393,N_17622,N_16997);
nand U19394 (N_19394,N_17446,N_17009);
and U19395 (N_19395,N_17958,N_15264);
or U19396 (N_19396,N_15460,N_16468);
or U19397 (N_19397,N_16215,N_17725);
or U19398 (N_19398,N_15377,N_17504);
or U19399 (N_19399,N_17148,N_16941);
xor U19400 (N_19400,N_16686,N_15403);
xnor U19401 (N_19401,N_17763,N_17759);
nand U19402 (N_19402,N_16748,N_17163);
or U19403 (N_19403,N_15407,N_16961);
xnor U19404 (N_19404,N_17192,N_15579);
xnor U19405 (N_19405,N_16433,N_17833);
and U19406 (N_19406,N_17094,N_17931);
nand U19407 (N_19407,N_16946,N_16422);
and U19408 (N_19408,N_16268,N_16878);
xnor U19409 (N_19409,N_17585,N_17356);
or U19410 (N_19410,N_16436,N_16764);
xor U19411 (N_19411,N_17782,N_17279);
nand U19412 (N_19412,N_16143,N_16621);
and U19413 (N_19413,N_15963,N_15150);
and U19414 (N_19414,N_16632,N_17269);
nor U19415 (N_19415,N_17757,N_16475);
nand U19416 (N_19416,N_17802,N_15446);
xor U19417 (N_19417,N_15191,N_17694);
or U19418 (N_19418,N_17976,N_17503);
xnor U19419 (N_19419,N_16671,N_17061);
nor U19420 (N_19420,N_17854,N_15273);
nor U19421 (N_19421,N_16151,N_17687);
and U19422 (N_19422,N_16345,N_17114);
xnor U19423 (N_19423,N_16277,N_17756);
xnor U19424 (N_19424,N_16399,N_15687);
or U19425 (N_19425,N_17372,N_15059);
xnor U19426 (N_19426,N_15644,N_15787);
nand U19427 (N_19427,N_17025,N_16943);
or U19428 (N_19428,N_16727,N_17112);
nor U19429 (N_19429,N_15185,N_16974);
nor U19430 (N_19430,N_16683,N_15988);
xnor U19431 (N_19431,N_15720,N_17016);
nand U19432 (N_19432,N_15402,N_15461);
xnor U19433 (N_19433,N_15023,N_15469);
nand U19434 (N_19434,N_16320,N_16743);
nand U19435 (N_19435,N_17532,N_17827);
and U19436 (N_19436,N_16112,N_17217);
or U19437 (N_19437,N_16984,N_16183);
or U19438 (N_19438,N_15926,N_16752);
nand U19439 (N_19439,N_15135,N_16491);
and U19440 (N_19440,N_17421,N_17987);
and U19441 (N_19441,N_15283,N_17881);
nand U19442 (N_19442,N_15411,N_15189);
xor U19443 (N_19443,N_17580,N_17234);
nand U19444 (N_19444,N_17443,N_17065);
nor U19445 (N_19445,N_17411,N_16767);
xnor U19446 (N_19446,N_17512,N_15863);
nand U19447 (N_19447,N_16575,N_15358);
nor U19448 (N_19448,N_17579,N_17817);
xor U19449 (N_19449,N_15004,N_15480);
nor U19450 (N_19450,N_16453,N_16972);
or U19451 (N_19451,N_16753,N_15318);
or U19452 (N_19452,N_16047,N_16751);
and U19453 (N_19453,N_17885,N_17568);
xor U19454 (N_19454,N_15516,N_17227);
nand U19455 (N_19455,N_17271,N_16643);
nand U19456 (N_19456,N_16606,N_17671);
xor U19457 (N_19457,N_17160,N_16554);
nor U19458 (N_19458,N_15728,N_17871);
xnor U19459 (N_19459,N_17660,N_17943);
nand U19460 (N_19460,N_16927,N_15111);
xor U19461 (N_19461,N_17483,N_15007);
nand U19462 (N_19462,N_15070,N_17389);
xor U19463 (N_19463,N_16741,N_17584);
and U19464 (N_19464,N_16918,N_16136);
nand U19465 (N_19465,N_16594,N_16822);
or U19466 (N_19466,N_16445,N_16370);
xnor U19467 (N_19467,N_17340,N_15504);
nand U19468 (N_19468,N_15270,N_16482);
or U19469 (N_19469,N_16252,N_16356);
nor U19470 (N_19470,N_15870,N_15305);
xor U19471 (N_19471,N_17731,N_15606);
xor U19472 (N_19472,N_16602,N_15908);
xnor U19473 (N_19473,N_17489,N_15152);
nand U19474 (N_19474,N_15458,N_17256);
xor U19475 (N_19475,N_15823,N_17869);
nand U19476 (N_19476,N_16005,N_15910);
nand U19477 (N_19477,N_15986,N_16090);
nand U19478 (N_19478,N_16220,N_17619);
and U19479 (N_19479,N_17440,N_16566);
nor U19480 (N_19480,N_17890,N_15168);
or U19481 (N_19481,N_16459,N_16076);
nand U19482 (N_19482,N_15293,N_16419);
and U19483 (N_19483,N_15764,N_15103);
and U19484 (N_19484,N_15471,N_15329);
or U19485 (N_19485,N_17659,N_17648);
and U19486 (N_19486,N_16481,N_15732);
nand U19487 (N_19487,N_15872,N_16618);
xnor U19488 (N_19488,N_17042,N_15747);
xor U19489 (N_19489,N_16505,N_15585);
nor U19490 (N_19490,N_15885,N_15188);
or U19491 (N_19491,N_16493,N_17216);
xnor U19492 (N_19492,N_15419,N_15592);
and U19493 (N_19493,N_15077,N_16119);
xor U19494 (N_19494,N_17138,N_17529);
or U19495 (N_19495,N_16257,N_17994);
nor U19496 (N_19496,N_15557,N_16196);
xnor U19497 (N_19497,N_15662,N_17119);
and U19498 (N_19498,N_16673,N_15349);
nand U19499 (N_19499,N_17978,N_17954);
and U19500 (N_19500,N_16858,N_17774);
nor U19501 (N_19501,N_16298,N_17823);
nor U19502 (N_19502,N_15968,N_15041);
or U19503 (N_19503,N_15908,N_15960);
nor U19504 (N_19504,N_15063,N_17601);
nand U19505 (N_19505,N_17381,N_16114);
nand U19506 (N_19506,N_17269,N_17811);
nand U19507 (N_19507,N_15886,N_17255);
or U19508 (N_19508,N_16288,N_16530);
xnor U19509 (N_19509,N_16143,N_16605);
nand U19510 (N_19510,N_15453,N_16872);
nor U19511 (N_19511,N_16598,N_15562);
and U19512 (N_19512,N_17718,N_17668);
nand U19513 (N_19513,N_17049,N_17034);
nor U19514 (N_19514,N_16441,N_16834);
and U19515 (N_19515,N_16049,N_15675);
or U19516 (N_19516,N_15301,N_17053);
or U19517 (N_19517,N_15250,N_17734);
nor U19518 (N_19518,N_15093,N_16506);
or U19519 (N_19519,N_16924,N_16324);
nand U19520 (N_19520,N_17839,N_17263);
nor U19521 (N_19521,N_16877,N_15417);
nor U19522 (N_19522,N_15526,N_17763);
nand U19523 (N_19523,N_17762,N_16652);
nand U19524 (N_19524,N_16066,N_16578);
and U19525 (N_19525,N_17937,N_15411);
or U19526 (N_19526,N_15523,N_16283);
and U19527 (N_19527,N_16290,N_16580);
nor U19528 (N_19528,N_16078,N_15627);
xnor U19529 (N_19529,N_17142,N_15379);
and U19530 (N_19530,N_17554,N_16807);
and U19531 (N_19531,N_15656,N_16290);
and U19532 (N_19532,N_15333,N_15489);
and U19533 (N_19533,N_16103,N_17162);
nor U19534 (N_19534,N_15820,N_15016);
or U19535 (N_19535,N_15245,N_17347);
or U19536 (N_19536,N_15309,N_16334);
nand U19537 (N_19537,N_17422,N_16983);
nand U19538 (N_19538,N_17005,N_17943);
xnor U19539 (N_19539,N_17799,N_15455);
or U19540 (N_19540,N_17477,N_15725);
nor U19541 (N_19541,N_16197,N_15557);
nand U19542 (N_19542,N_17131,N_15569);
xor U19543 (N_19543,N_16038,N_15560);
nand U19544 (N_19544,N_16744,N_15586);
or U19545 (N_19545,N_15948,N_16440);
xor U19546 (N_19546,N_17951,N_15872);
or U19547 (N_19547,N_16748,N_16441);
nand U19548 (N_19548,N_15229,N_16612);
nand U19549 (N_19549,N_16625,N_15119);
xor U19550 (N_19550,N_17093,N_16612);
or U19551 (N_19551,N_15786,N_16676);
nor U19552 (N_19552,N_15449,N_16078);
nor U19553 (N_19553,N_15962,N_16952);
xnor U19554 (N_19554,N_17462,N_17266);
xor U19555 (N_19555,N_16914,N_17493);
nand U19556 (N_19556,N_17973,N_16796);
xnor U19557 (N_19557,N_17417,N_17325);
nand U19558 (N_19558,N_17312,N_15093);
nor U19559 (N_19559,N_15906,N_15063);
nand U19560 (N_19560,N_17589,N_15169);
or U19561 (N_19561,N_17523,N_15536);
nand U19562 (N_19562,N_16905,N_15731);
nand U19563 (N_19563,N_15549,N_16120);
nor U19564 (N_19564,N_16033,N_16908);
nor U19565 (N_19565,N_15119,N_16729);
nor U19566 (N_19566,N_16565,N_16961);
xnor U19567 (N_19567,N_16976,N_17166);
nor U19568 (N_19568,N_17498,N_16581);
nor U19569 (N_19569,N_16824,N_15981);
nand U19570 (N_19570,N_16279,N_15582);
nand U19571 (N_19571,N_17066,N_17273);
or U19572 (N_19572,N_16304,N_17934);
or U19573 (N_19573,N_15821,N_16271);
nor U19574 (N_19574,N_17273,N_16626);
xnor U19575 (N_19575,N_16308,N_15300);
and U19576 (N_19576,N_16004,N_15286);
nand U19577 (N_19577,N_17239,N_16906);
xnor U19578 (N_19578,N_15807,N_15004);
nand U19579 (N_19579,N_15938,N_16092);
and U19580 (N_19580,N_17417,N_17891);
xor U19581 (N_19581,N_16076,N_15310);
or U19582 (N_19582,N_16953,N_16926);
and U19583 (N_19583,N_16393,N_15417);
and U19584 (N_19584,N_17502,N_17369);
and U19585 (N_19585,N_15786,N_17945);
or U19586 (N_19586,N_15798,N_15346);
nor U19587 (N_19587,N_17459,N_17046);
and U19588 (N_19588,N_17772,N_15533);
xnor U19589 (N_19589,N_17824,N_17703);
and U19590 (N_19590,N_16374,N_15959);
nand U19591 (N_19591,N_15860,N_17472);
and U19592 (N_19592,N_16845,N_16145);
xor U19593 (N_19593,N_16029,N_16313);
nor U19594 (N_19594,N_15763,N_16115);
and U19595 (N_19595,N_16013,N_16729);
nor U19596 (N_19596,N_15625,N_17328);
nand U19597 (N_19597,N_15189,N_15697);
nand U19598 (N_19598,N_17979,N_17357);
or U19599 (N_19599,N_17106,N_15548);
or U19600 (N_19600,N_15945,N_16299);
nor U19601 (N_19601,N_17574,N_15619);
nor U19602 (N_19602,N_15000,N_17725);
nor U19603 (N_19603,N_16589,N_17348);
nor U19604 (N_19604,N_15734,N_15547);
nand U19605 (N_19605,N_17315,N_17759);
and U19606 (N_19606,N_17245,N_17154);
or U19607 (N_19607,N_15651,N_17309);
xor U19608 (N_19608,N_17863,N_16606);
xnor U19609 (N_19609,N_16809,N_16909);
nand U19610 (N_19610,N_16287,N_16793);
nor U19611 (N_19611,N_15428,N_15385);
xor U19612 (N_19612,N_16848,N_16282);
nor U19613 (N_19613,N_16741,N_17311);
xor U19614 (N_19614,N_16207,N_17461);
nor U19615 (N_19615,N_16250,N_16624);
nor U19616 (N_19616,N_15135,N_16351);
or U19617 (N_19617,N_15318,N_16396);
and U19618 (N_19618,N_15709,N_16586);
and U19619 (N_19619,N_16411,N_17485);
xor U19620 (N_19620,N_15624,N_17836);
nand U19621 (N_19621,N_15286,N_16536);
nor U19622 (N_19622,N_17943,N_17143);
nand U19623 (N_19623,N_16985,N_17782);
or U19624 (N_19624,N_15140,N_15102);
or U19625 (N_19625,N_15189,N_15572);
nand U19626 (N_19626,N_15736,N_16204);
or U19627 (N_19627,N_15274,N_17438);
nor U19628 (N_19628,N_17990,N_16659);
and U19629 (N_19629,N_16892,N_15673);
nand U19630 (N_19630,N_15432,N_15226);
or U19631 (N_19631,N_16148,N_17850);
nor U19632 (N_19632,N_16463,N_15226);
nand U19633 (N_19633,N_17430,N_17485);
and U19634 (N_19634,N_17787,N_15676);
and U19635 (N_19635,N_16208,N_15538);
and U19636 (N_19636,N_15976,N_16690);
xor U19637 (N_19637,N_17093,N_15624);
nand U19638 (N_19638,N_17128,N_15253);
xnor U19639 (N_19639,N_16797,N_17292);
xnor U19640 (N_19640,N_15678,N_17431);
nand U19641 (N_19641,N_15315,N_16850);
and U19642 (N_19642,N_17135,N_17153);
xnor U19643 (N_19643,N_15868,N_15178);
xnor U19644 (N_19644,N_16084,N_15286);
nor U19645 (N_19645,N_16777,N_15437);
or U19646 (N_19646,N_15028,N_16041);
or U19647 (N_19647,N_16250,N_17313);
nor U19648 (N_19648,N_15543,N_16611);
and U19649 (N_19649,N_15874,N_15237);
and U19650 (N_19650,N_16969,N_17362);
nor U19651 (N_19651,N_15484,N_17196);
or U19652 (N_19652,N_16780,N_15147);
nor U19653 (N_19653,N_15483,N_15922);
nor U19654 (N_19654,N_17369,N_17217);
or U19655 (N_19655,N_16221,N_17000);
xnor U19656 (N_19656,N_15080,N_16671);
or U19657 (N_19657,N_15193,N_15702);
xnor U19658 (N_19658,N_17167,N_16714);
xor U19659 (N_19659,N_16601,N_15405);
or U19660 (N_19660,N_15925,N_15703);
xor U19661 (N_19661,N_17188,N_15774);
nand U19662 (N_19662,N_17399,N_16392);
and U19663 (N_19663,N_16778,N_16925);
xnor U19664 (N_19664,N_15863,N_17087);
nand U19665 (N_19665,N_17966,N_16364);
nor U19666 (N_19666,N_17423,N_17553);
nor U19667 (N_19667,N_17446,N_15340);
xnor U19668 (N_19668,N_15333,N_16832);
nor U19669 (N_19669,N_16005,N_15508);
nand U19670 (N_19670,N_16890,N_17578);
nand U19671 (N_19671,N_15024,N_16672);
and U19672 (N_19672,N_16193,N_16715);
and U19673 (N_19673,N_17899,N_16193);
and U19674 (N_19674,N_15359,N_15678);
nand U19675 (N_19675,N_17085,N_16143);
nor U19676 (N_19676,N_17310,N_15189);
nor U19677 (N_19677,N_15279,N_15753);
nor U19678 (N_19678,N_17665,N_15599);
nand U19679 (N_19679,N_17939,N_16473);
or U19680 (N_19680,N_16990,N_16706);
or U19681 (N_19681,N_16162,N_16857);
or U19682 (N_19682,N_15052,N_17515);
nor U19683 (N_19683,N_17059,N_15118);
and U19684 (N_19684,N_17459,N_15730);
or U19685 (N_19685,N_17816,N_17003);
and U19686 (N_19686,N_16958,N_15989);
or U19687 (N_19687,N_16403,N_16440);
nor U19688 (N_19688,N_17656,N_17964);
or U19689 (N_19689,N_17177,N_17604);
nor U19690 (N_19690,N_16728,N_16481);
xnor U19691 (N_19691,N_17461,N_16109);
nor U19692 (N_19692,N_16132,N_16736);
nand U19693 (N_19693,N_16927,N_16286);
nand U19694 (N_19694,N_17680,N_17860);
and U19695 (N_19695,N_17401,N_15147);
nor U19696 (N_19696,N_17664,N_15535);
or U19697 (N_19697,N_17405,N_16430);
xor U19698 (N_19698,N_16429,N_17993);
or U19699 (N_19699,N_15679,N_17742);
nand U19700 (N_19700,N_16602,N_15743);
xor U19701 (N_19701,N_16253,N_17810);
nand U19702 (N_19702,N_17340,N_17890);
nor U19703 (N_19703,N_15692,N_15376);
xnor U19704 (N_19704,N_16164,N_15894);
xnor U19705 (N_19705,N_15155,N_17111);
and U19706 (N_19706,N_17552,N_15509);
xor U19707 (N_19707,N_16613,N_16355);
nand U19708 (N_19708,N_17163,N_15525);
or U19709 (N_19709,N_15041,N_16436);
xor U19710 (N_19710,N_17412,N_15071);
xor U19711 (N_19711,N_16977,N_16029);
nand U19712 (N_19712,N_15561,N_17337);
or U19713 (N_19713,N_17084,N_17194);
xnor U19714 (N_19714,N_15632,N_17425);
nor U19715 (N_19715,N_15873,N_17290);
nand U19716 (N_19716,N_17616,N_15869);
nand U19717 (N_19717,N_17704,N_16324);
and U19718 (N_19718,N_17764,N_17573);
nand U19719 (N_19719,N_15685,N_16583);
xor U19720 (N_19720,N_17243,N_17000);
xor U19721 (N_19721,N_17402,N_17930);
nand U19722 (N_19722,N_15423,N_15285);
nand U19723 (N_19723,N_16868,N_15468);
or U19724 (N_19724,N_16992,N_15523);
nor U19725 (N_19725,N_17255,N_16774);
and U19726 (N_19726,N_15273,N_16943);
nor U19727 (N_19727,N_16564,N_17595);
nor U19728 (N_19728,N_16926,N_17753);
or U19729 (N_19729,N_15112,N_15552);
and U19730 (N_19730,N_17501,N_15694);
and U19731 (N_19731,N_16658,N_15127);
nor U19732 (N_19732,N_15275,N_16730);
xnor U19733 (N_19733,N_17592,N_16016);
xor U19734 (N_19734,N_16188,N_15931);
nor U19735 (N_19735,N_16484,N_16545);
and U19736 (N_19736,N_15075,N_17418);
or U19737 (N_19737,N_17629,N_17459);
nand U19738 (N_19738,N_16763,N_17360);
and U19739 (N_19739,N_16983,N_16914);
nor U19740 (N_19740,N_15663,N_15577);
and U19741 (N_19741,N_17638,N_17978);
and U19742 (N_19742,N_17679,N_16559);
and U19743 (N_19743,N_15491,N_16906);
or U19744 (N_19744,N_15467,N_16822);
or U19745 (N_19745,N_15419,N_15465);
or U19746 (N_19746,N_15087,N_15414);
nor U19747 (N_19747,N_17993,N_15456);
nand U19748 (N_19748,N_17710,N_17715);
xnor U19749 (N_19749,N_16919,N_16665);
nand U19750 (N_19750,N_17665,N_17748);
nand U19751 (N_19751,N_16064,N_16597);
nor U19752 (N_19752,N_15102,N_15264);
nand U19753 (N_19753,N_17343,N_15832);
xnor U19754 (N_19754,N_17321,N_17636);
and U19755 (N_19755,N_15316,N_15788);
and U19756 (N_19756,N_17156,N_17199);
xnor U19757 (N_19757,N_16661,N_16215);
and U19758 (N_19758,N_15314,N_16389);
or U19759 (N_19759,N_15255,N_17717);
and U19760 (N_19760,N_16095,N_17901);
nor U19761 (N_19761,N_17692,N_17375);
and U19762 (N_19762,N_15477,N_17330);
nand U19763 (N_19763,N_16746,N_17312);
nor U19764 (N_19764,N_16876,N_16265);
and U19765 (N_19765,N_16609,N_15407);
xor U19766 (N_19766,N_16135,N_15784);
or U19767 (N_19767,N_16131,N_17833);
and U19768 (N_19768,N_15640,N_17009);
and U19769 (N_19769,N_15556,N_17864);
and U19770 (N_19770,N_17648,N_17635);
and U19771 (N_19771,N_16729,N_17549);
xor U19772 (N_19772,N_17995,N_15007);
nand U19773 (N_19773,N_17872,N_15408);
nand U19774 (N_19774,N_17327,N_16952);
nor U19775 (N_19775,N_15834,N_17631);
nand U19776 (N_19776,N_17137,N_17178);
nand U19777 (N_19777,N_15945,N_17298);
xnor U19778 (N_19778,N_16070,N_15076);
or U19779 (N_19779,N_15828,N_16747);
and U19780 (N_19780,N_16576,N_16305);
or U19781 (N_19781,N_15322,N_16635);
and U19782 (N_19782,N_15483,N_17168);
xor U19783 (N_19783,N_15556,N_16938);
xnor U19784 (N_19784,N_15267,N_17158);
nor U19785 (N_19785,N_15167,N_15858);
and U19786 (N_19786,N_15439,N_16461);
nor U19787 (N_19787,N_15405,N_17218);
nand U19788 (N_19788,N_15631,N_15014);
and U19789 (N_19789,N_15566,N_16312);
nor U19790 (N_19790,N_16510,N_16611);
or U19791 (N_19791,N_17223,N_16300);
xor U19792 (N_19792,N_15481,N_15706);
nand U19793 (N_19793,N_17388,N_16292);
xor U19794 (N_19794,N_15271,N_17482);
or U19795 (N_19795,N_16520,N_17196);
or U19796 (N_19796,N_17877,N_17178);
nor U19797 (N_19797,N_17235,N_15756);
xor U19798 (N_19798,N_15353,N_15945);
nor U19799 (N_19799,N_15591,N_15878);
xnor U19800 (N_19800,N_16102,N_16710);
nor U19801 (N_19801,N_17289,N_17907);
xor U19802 (N_19802,N_15979,N_16477);
and U19803 (N_19803,N_17544,N_16650);
and U19804 (N_19804,N_15556,N_16804);
or U19805 (N_19805,N_17689,N_17320);
xnor U19806 (N_19806,N_16283,N_15199);
nor U19807 (N_19807,N_17775,N_17144);
and U19808 (N_19808,N_17330,N_17758);
nand U19809 (N_19809,N_16275,N_16770);
nor U19810 (N_19810,N_16773,N_16811);
or U19811 (N_19811,N_17933,N_17077);
nand U19812 (N_19812,N_15143,N_17898);
nor U19813 (N_19813,N_16800,N_17016);
and U19814 (N_19814,N_16470,N_17767);
nor U19815 (N_19815,N_15618,N_16309);
nand U19816 (N_19816,N_15107,N_16705);
and U19817 (N_19817,N_15043,N_16127);
nand U19818 (N_19818,N_15874,N_17566);
xnor U19819 (N_19819,N_17522,N_17851);
and U19820 (N_19820,N_16974,N_17582);
nor U19821 (N_19821,N_15087,N_15824);
xnor U19822 (N_19822,N_17620,N_17728);
and U19823 (N_19823,N_17959,N_15324);
nor U19824 (N_19824,N_16115,N_17826);
and U19825 (N_19825,N_17434,N_15440);
nand U19826 (N_19826,N_16911,N_15676);
and U19827 (N_19827,N_17549,N_17750);
or U19828 (N_19828,N_16194,N_16976);
and U19829 (N_19829,N_16767,N_17882);
xor U19830 (N_19830,N_16756,N_16491);
and U19831 (N_19831,N_15664,N_15024);
nand U19832 (N_19832,N_16390,N_16556);
nand U19833 (N_19833,N_17401,N_16613);
or U19834 (N_19834,N_15948,N_16039);
xnor U19835 (N_19835,N_16243,N_17148);
or U19836 (N_19836,N_16243,N_17774);
nor U19837 (N_19837,N_16476,N_15843);
xor U19838 (N_19838,N_16672,N_16138);
or U19839 (N_19839,N_16887,N_16219);
or U19840 (N_19840,N_15276,N_16978);
xor U19841 (N_19841,N_16478,N_15309);
and U19842 (N_19842,N_16191,N_15174);
nand U19843 (N_19843,N_17607,N_17330);
xor U19844 (N_19844,N_15420,N_17308);
nor U19845 (N_19845,N_16618,N_17536);
nand U19846 (N_19846,N_15196,N_15009);
and U19847 (N_19847,N_15116,N_16215);
and U19848 (N_19848,N_15684,N_15071);
or U19849 (N_19849,N_16863,N_16647);
xor U19850 (N_19850,N_16800,N_17265);
nand U19851 (N_19851,N_17430,N_15882);
nand U19852 (N_19852,N_16923,N_16667);
nor U19853 (N_19853,N_16775,N_16166);
nor U19854 (N_19854,N_15027,N_15086);
xnor U19855 (N_19855,N_15234,N_15909);
or U19856 (N_19856,N_17583,N_16705);
or U19857 (N_19857,N_17967,N_15735);
nand U19858 (N_19858,N_16386,N_16221);
nor U19859 (N_19859,N_16033,N_16273);
xnor U19860 (N_19860,N_16847,N_16588);
and U19861 (N_19861,N_16468,N_16399);
and U19862 (N_19862,N_17773,N_15137);
and U19863 (N_19863,N_17013,N_15817);
nand U19864 (N_19864,N_16444,N_16578);
and U19865 (N_19865,N_16043,N_15346);
nor U19866 (N_19866,N_15870,N_16109);
or U19867 (N_19867,N_15979,N_15889);
or U19868 (N_19868,N_16220,N_16365);
nor U19869 (N_19869,N_15090,N_16375);
or U19870 (N_19870,N_16049,N_15557);
nor U19871 (N_19871,N_17835,N_15452);
nor U19872 (N_19872,N_15894,N_17661);
nor U19873 (N_19873,N_15096,N_17485);
and U19874 (N_19874,N_15258,N_17884);
and U19875 (N_19875,N_16861,N_15874);
or U19876 (N_19876,N_17033,N_15193);
nand U19877 (N_19877,N_17080,N_17407);
or U19878 (N_19878,N_16399,N_15514);
or U19879 (N_19879,N_16661,N_15305);
or U19880 (N_19880,N_16643,N_17612);
or U19881 (N_19881,N_16804,N_16362);
and U19882 (N_19882,N_16141,N_15566);
or U19883 (N_19883,N_17496,N_17939);
xor U19884 (N_19884,N_16854,N_17871);
xor U19885 (N_19885,N_15339,N_15324);
nor U19886 (N_19886,N_15117,N_17816);
or U19887 (N_19887,N_15199,N_16566);
nor U19888 (N_19888,N_17396,N_16380);
nor U19889 (N_19889,N_17480,N_15483);
nand U19890 (N_19890,N_15989,N_16358);
nand U19891 (N_19891,N_16847,N_15395);
nor U19892 (N_19892,N_17383,N_15942);
and U19893 (N_19893,N_16635,N_15954);
xnor U19894 (N_19894,N_16312,N_15789);
and U19895 (N_19895,N_16579,N_17774);
xor U19896 (N_19896,N_16967,N_16307);
and U19897 (N_19897,N_16790,N_16865);
xnor U19898 (N_19898,N_17399,N_17030);
and U19899 (N_19899,N_16738,N_17795);
or U19900 (N_19900,N_17282,N_16004);
or U19901 (N_19901,N_16072,N_16353);
xnor U19902 (N_19902,N_17417,N_15978);
or U19903 (N_19903,N_16753,N_15087);
and U19904 (N_19904,N_15901,N_17058);
nor U19905 (N_19905,N_16040,N_17954);
nor U19906 (N_19906,N_15962,N_15701);
or U19907 (N_19907,N_16235,N_17531);
or U19908 (N_19908,N_17078,N_15617);
and U19909 (N_19909,N_16917,N_16314);
and U19910 (N_19910,N_15719,N_17759);
or U19911 (N_19911,N_16530,N_15027);
nand U19912 (N_19912,N_15777,N_15546);
nor U19913 (N_19913,N_16575,N_15695);
nor U19914 (N_19914,N_16919,N_17066);
nand U19915 (N_19915,N_16353,N_15643);
nor U19916 (N_19916,N_15077,N_17305);
nand U19917 (N_19917,N_15986,N_17737);
xnor U19918 (N_19918,N_15923,N_15106);
and U19919 (N_19919,N_17467,N_17393);
or U19920 (N_19920,N_16696,N_17980);
or U19921 (N_19921,N_15738,N_15999);
xor U19922 (N_19922,N_15780,N_16943);
or U19923 (N_19923,N_17460,N_15620);
and U19924 (N_19924,N_17069,N_16154);
nor U19925 (N_19925,N_17556,N_16012);
nor U19926 (N_19926,N_15253,N_17298);
or U19927 (N_19927,N_17202,N_15235);
xor U19928 (N_19928,N_15520,N_17305);
xnor U19929 (N_19929,N_17077,N_17883);
xnor U19930 (N_19930,N_17610,N_17983);
xnor U19931 (N_19931,N_17984,N_16716);
and U19932 (N_19932,N_15755,N_16261);
or U19933 (N_19933,N_17026,N_17164);
and U19934 (N_19934,N_16895,N_16456);
xnor U19935 (N_19935,N_17187,N_15640);
nor U19936 (N_19936,N_16253,N_16002);
xor U19937 (N_19937,N_16752,N_17456);
nor U19938 (N_19938,N_16088,N_17945);
xnor U19939 (N_19939,N_15642,N_17479);
or U19940 (N_19940,N_15381,N_15861);
nor U19941 (N_19941,N_15369,N_16846);
nor U19942 (N_19942,N_17776,N_15267);
nand U19943 (N_19943,N_16602,N_16990);
and U19944 (N_19944,N_15222,N_17870);
nor U19945 (N_19945,N_16357,N_17981);
or U19946 (N_19946,N_16530,N_17483);
xor U19947 (N_19947,N_17435,N_17337);
and U19948 (N_19948,N_17861,N_15014);
or U19949 (N_19949,N_16763,N_15937);
nor U19950 (N_19950,N_15098,N_16622);
nor U19951 (N_19951,N_15933,N_15650);
xnor U19952 (N_19952,N_16470,N_16239);
xnor U19953 (N_19953,N_17266,N_16975);
nor U19954 (N_19954,N_15819,N_15025);
nor U19955 (N_19955,N_17729,N_15600);
nand U19956 (N_19956,N_15610,N_16269);
nand U19957 (N_19957,N_15590,N_16478);
nor U19958 (N_19958,N_16694,N_15295);
and U19959 (N_19959,N_15867,N_17930);
nand U19960 (N_19960,N_17729,N_17572);
nor U19961 (N_19961,N_16342,N_15505);
nor U19962 (N_19962,N_15149,N_16980);
xnor U19963 (N_19963,N_17620,N_16664);
and U19964 (N_19964,N_17110,N_15898);
xor U19965 (N_19965,N_15626,N_17845);
xnor U19966 (N_19966,N_17272,N_17396);
xor U19967 (N_19967,N_15609,N_15248);
nand U19968 (N_19968,N_17980,N_17119);
and U19969 (N_19969,N_16019,N_16053);
or U19970 (N_19970,N_17293,N_17216);
nor U19971 (N_19971,N_16605,N_16406);
or U19972 (N_19972,N_17135,N_17673);
nor U19973 (N_19973,N_15767,N_17589);
nor U19974 (N_19974,N_17240,N_16037);
nor U19975 (N_19975,N_17201,N_15113);
nor U19976 (N_19976,N_17564,N_17528);
xnor U19977 (N_19977,N_15841,N_15843);
and U19978 (N_19978,N_17698,N_16229);
nor U19979 (N_19979,N_16246,N_16402);
or U19980 (N_19980,N_15037,N_15754);
or U19981 (N_19981,N_16186,N_16917);
xor U19982 (N_19982,N_16363,N_15222);
and U19983 (N_19983,N_15454,N_17521);
xnor U19984 (N_19984,N_17071,N_16783);
or U19985 (N_19985,N_16404,N_15288);
or U19986 (N_19986,N_17731,N_16871);
or U19987 (N_19987,N_16650,N_15949);
nand U19988 (N_19988,N_15142,N_15506);
or U19989 (N_19989,N_17953,N_15234);
xnor U19990 (N_19990,N_17226,N_17752);
xor U19991 (N_19991,N_15985,N_15930);
xnor U19992 (N_19992,N_15728,N_17428);
xnor U19993 (N_19993,N_16436,N_17849);
xor U19994 (N_19994,N_16263,N_15887);
or U19995 (N_19995,N_15417,N_17814);
xnor U19996 (N_19996,N_17428,N_17254);
or U19997 (N_19997,N_16996,N_15007);
nand U19998 (N_19998,N_16920,N_17464);
and U19999 (N_19999,N_15566,N_17008);
or U20000 (N_20000,N_17004,N_15564);
nand U20001 (N_20001,N_16866,N_16492);
nor U20002 (N_20002,N_16454,N_16738);
nor U20003 (N_20003,N_16695,N_17817);
nand U20004 (N_20004,N_17286,N_15163);
or U20005 (N_20005,N_16375,N_17036);
nor U20006 (N_20006,N_17197,N_17251);
nand U20007 (N_20007,N_15003,N_15087);
xor U20008 (N_20008,N_17902,N_15888);
nand U20009 (N_20009,N_16985,N_15468);
and U20010 (N_20010,N_15903,N_17694);
nor U20011 (N_20011,N_16768,N_16242);
xor U20012 (N_20012,N_16179,N_15611);
nor U20013 (N_20013,N_15339,N_16274);
nand U20014 (N_20014,N_17943,N_17177);
nor U20015 (N_20015,N_17718,N_15023);
or U20016 (N_20016,N_15027,N_15745);
or U20017 (N_20017,N_15657,N_15238);
or U20018 (N_20018,N_16296,N_17860);
nor U20019 (N_20019,N_15726,N_17573);
xor U20020 (N_20020,N_15172,N_17792);
nor U20021 (N_20021,N_16403,N_16364);
or U20022 (N_20022,N_16150,N_16255);
or U20023 (N_20023,N_17761,N_15458);
nor U20024 (N_20024,N_15317,N_15948);
or U20025 (N_20025,N_17227,N_16443);
xor U20026 (N_20026,N_16187,N_17584);
nand U20027 (N_20027,N_17567,N_16958);
nor U20028 (N_20028,N_16596,N_17120);
nand U20029 (N_20029,N_16308,N_17945);
or U20030 (N_20030,N_16318,N_15487);
nand U20031 (N_20031,N_16210,N_17688);
or U20032 (N_20032,N_17293,N_17024);
xnor U20033 (N_20033,N_15686,N_17895);
nor U20034 (N_20034,N_15556,N_15333);
or U20035 (N_20035,N_15253,N_16644);
or U20036 (N_20036,N_16367,N_17711);
and U20037 (N_20037,N_17669,N_16763);
and U20038 (N_20038,N_15245,N_15679);
xor U20039 (N_20039,N_15014,N_15952);
nand U20040 (N_20040,N_15029,N_16875);
xnor U20041 (N_20041,N_17438,N_16639);
nor U20042 (N_20042,N_15802,N_17112);
and U20043 (N_20043,N_15850,N_15745);
nor U20044 (N_20044,N_17292,N_17310);
xnor U20045 (N_20045,N_16582,N_15490);
nand U20046 (N_20046,N_16304,N_17013);
nand U20047 (N_20047,N_17629,N_17109);
and U20048 (N_20048,N_16320,N_16815);
or U20049 (N_20049,N_17108,N_16889);
nor U20050 (N_20050,N_17578,N_16856);
or U20051 (N_20051,N_17231,N_16831);
nand U20052 (N_20052,N_15433,N_15030);
or U20053 (N_20053,N_15078,N_17685);
and U20054 (N_20054,N_16189,N_16079);
nor U20055 (N_20055,N_16831,N_16985);
or U20056 (N_20056,N_16251,N_16338);
xnor U20057 (N_20057,N_17809,N_16493);
nor U20058 (N_20058,N_15940,N_15429);
and U20059 (N_20059,N_17478,N_15305);
xnor U20060 (N_20060,N_17004,N_15386);
or U20061 (N_20061,N_16367,N_16005);
nand U20062 (N_20062,N_16787,N_16024);
and U20063 (N_20063,N_16145,N_16249);
or U20064 (N_20064,N_16136,N_15074);
xor U20065 (N_20065,N_17538,N_16247);
nor U20066 (N_20066,N_16523,N_15916);
and U20067 (N_20067,N_15388,N_15133);
and U20068 (N_20068,N_15325,N_17805);
and U20069 (N_20069,N_16173,N_15449);
and U20070 (N_20070,N_17314,N_16783);
nand U20071 (N_20071,N_16759,N_16019);
xor U20072 (N_20072,N_16257,N_16314);
xor U20073 (N_20073,N_17690,N_17565);
nand U20074 (N_20074,N_15165,N_15914);
or U20075 (N_20075,N_15373,N_17765);
xor U20076 (N_20076,N_16729,N_16066);
or U20077 (N_20077,N_16394,N_15977);
and U20078 (N_20078,N_15756,N_17365);
nand U20079 (N_20079,N_17229,N_15656);
or U20080 (N_20080,N_17628,N_15285);
nand U20081 (N_20081,N_16894,N_17354);
and U20082 (N_20082,N_15953,N_15841);
nand U20083 (N_20083,N_16140,N_16462);
xnor U20084 (N_20084,N_16377,N_16141);
nor U20085 (N_20085,N_15410,N_17915);
xnor U20086 (N_20086,N_17003,N_17055);
or U20087 (N_20087,N_17632,N_15734);
nor U20088 (N_20088,N_17732,N_17536);
and U20089 (N_20089,N_15466,N_15407);
xor U20090 (N_20090,N_15395,N_17470);
xnor U20091 (N_20091,N_17020,N_16213);
and U20092 (N_20092,N_16749,N_15192);
nor U20093 (N_20093,N_16208,N_17255);
nor U20094 (N_20094,N_16443,N_17800);
nand U20095 (N_20095,N_17431,N_17692);
xnor U20096 (N_20096,N_17136,N_15816);
xnor U20097 (N_20097,N_15568,N_17747);
nand U20098 (N_20098,N_17904,N_17032);
nor U20099 (N_20099,N_17942,N_16370);
or U20100 (N_20100,N_17715,N_15840);
or U20101 (N_20101,N_16580,N_15279);
nor U20102 (N_20102,N_17001,N_16783);
nor U20103 (N_20103,N_15824,N_15046);
or U20104 (N_20104,N_15485,N_17637);
nor U20105 (N_20105,N_17834,N_16273);
and U20106 (N_20106,N_17015,N_15708);
nor U20107 (N_20107,N_17985,N_16254);
nand U20108 (N_20108,N_15004,N_17074);
xor U20109 (N_20109,N_17400,N_17278);
or U20110 (N_20110,N_15774,N_17714);
nor U20111 (N_20111,N_16963,N_15057);
xnor U20112 (N_20112,N_15635,N_17683);
xnor U20113 (N_20113,N_15701,N_17404);
nor U20114 (N_20114,N_15153,N_16705);
and U20115 (N_20115,N_17451,N_16120);
nand U20116 (N_20116,N_16059,N_16511);
xor U20117 (N_20117,N_17613,N_16159);
xor U20118 (N_20118,N_15977,N_16404);
nand U20119 (N_20119,N_17684,N_17727);
and U20120 (N_20120,N_15462,N_17584);
nand U20121 (N_20121,N_17649,N_16274);
nand U20122 (N_20122,N_15051,N_17872);
or U20123 (N_20123,N_15974,N_15519);
nand U20124 (N_20124,N_15868,N_15692);
nor U20125 (N_20125,N_17019,N_16614);
nor U20126 (N_20126,N_16505,N_15573);
nor U20127 (N_20127,N_16367,N_17052);
xor U20128 (N_20128,N_15287,N_17026);
and U20129 (N_20129,N_16875,N_16703);
or U20130 (N_20130,N_17592,N_17282);
or U20131 (N_20131,N_16511,N_15101);
or U20132 (N_20132,N_15423,N_16857);
xnor U20133 (N_20133,N_17771,N_17029);
and U20134 (N_20134,N_17582,N_16370);
or U20135 (N_20135,N_17825,N_15388);
xor U20136 (N_20136,N_16688,N_15981);
and U20137 (N_20137,N_17761,N_15700);
and U20138 (N_20138,N_16016,N_16548);
nor U20139 (N_20139,N_15160,N_17889);
nor U20140 (N_20140,N_17220,N_16974);
or U20141 (N_20141,N_15988,N_16477);
nor U20142 (N_20142,N_17134,N_17533);
nand U20143 (N_20143,N_15285,N_15907);
nor U20144 (N_20144,N_17326,N_15689);
nand U20145 (N_20145,N_16326,N_15202);
nor U20146 (N_20146,N_17083,N_17481);
or U20147 (N_20147,N_15231,N_15532);
xnor U20148 (N_20148,N_17252,N_16962);
nor U20149 (N_20149,N_17733,N_15425);
nand U20150 (N_20150,N_16069,N_16819);
nand U20151 (N_20151,N_16300,N_15318);
and U20152 (N_20152,N_15944,N_16893);
nor U20153 (N_20153,N_15463,N_15029);
xnor U20154 (N_20154,N_15252,N_16404);
and U20155 (N_20155,N_17700,N_17960);
nor U20156 (N_20156,N_16474,N_15594);
nor U20157 (N_20157,N_16982,N_15146);
xor U20158 (N_20158,N_17751,N_17673);
nand U20159 (N_20159,N_17668,N_16977);
or U20160 (N_20160,N_17728,N_16974);
nand U20161 (N_20161,N_15287,N_16866);
nor U20162 (N_20162,N_15594,N_15660);
and U20163 (N_20163,N_15150,N_17916);
and U20164 (N_20164,N_15216,N_15753);
xnor U20165 (N_20165,N_16322,N_17965);
xnor U20166 (N_20166,N_15103,N_17714);
nor U20167 (N_20167,N_16741,N_16692);
or U20168 (N_20168,N_15285,N_16181);
xor U20169 (N_20169,N_17277,N_15593);
and U20170 (N_20170,N_17769,N_16508);
and U20171 (N_20171,N_17286,N_15629);
and U20172 (N_20172,N_17313,N_15848);
nand U20173 (N_20173,N_15911,N_17023);
or U20174 (N_20174,N_16686,N_15787);
nor U20175 (N_20175,N_17735,N_17949);
nor U20176 (N_20176,N_16749,N_16971);
nand U20177 (N_20177,N_17076,N_17149);
nand U20178 (N_20178,N_15151,N_16156);
nor U20179 (N_20179,N_15609,N_16958);
and U20180 (N_20180,N_16253,N_17648);
nor U20181 (N_20181,N_15030,N_16860);
and U20182 (N_20182,N_17929,N_15050);
xor U20183 (N_20183,N_15282,N_15512);
xnor U20184 (N_20184,N_16010,N_17416);
or U20185 (N_20185,N_16488,N_15271);
or U20186 (N_20186,N_15365,N_17343);
or U20187 (N_20187,N_16198,N_17615);
and U20188 (N_20188,N_16119,N_17910);
nor U20189 (N_20189,N_15196,N_16007);
or U20190 (N_20190,N_15873,N_17213);
or U20191 (N_20191,N_17988,N_16162);
and U20192 (N_20192,N_15429,N_15432);
xor U20193 (N_20193,N_15838,N_15325);
nor U20194 (N_20194,N_17308,N_17506);
or U20195 (N_20195,N_15259,N_17458);
or U20196 (N_20196,N_16477,N_15296);
xor U20197 (N_20197,N_17491,N_16374);
nand U20198 (N_20198,N_16879,N_17927);
and U20199 (N_20199,N_15805,N_15639);
nor U20200 (N_20200,N_15914,N_17614);
or U20201 (N_20201,N_15243,N_16284);
xnor U20202 (N_20202,N_16375,N_16470);
xnor U20203 (N_20203,N_15845,N_17142);
or U20204 (N_20204,N_17540,N_15020);
xnor U20205 (N_20205,N_17678,N_16864);
xnor U20206 (N_20206,N_15161,N_15744);
nor U20207 (N_20207,N_16951,N_16523);
or U20208 (N_20208,N_16353,N_16660);
and U20209 (N_20209,N_16320,N_16976);
nand U20210 (N_20210,N_15304,N_17583);
nand U20211 (N_20211,N_17490,N_16883);
or U20212 (N_20212,N_17647,N_16088);
nand U20213 (N_20213,N_16027,N_15857);
xnor U20214 (N_20214,N_16768,N_16980);
or U20215 (N_20215,N_17597,N_17492);
nand U20216 (N_20216,N_15518,N_16664);
xnor U20217 (N_20217,N_17888,N_16901);
or U20218 (N_20218,N_17167,N_15419);
and U20219 (N_20219,N_15864,N_15296);
nand U20220 (N_20220,N_16562,N_15696);
nor U20221 (N_20221,N_17958,N_15617);
nand U20222 (N_20222,N_17352,N_16217);
xor U20223 (N_20223,N_17077,N_15446);
or U20224 (N_20224,N_16994,N_17140);
nand U20225 (N_20225,N_15710,N_16500);
and U20226 (N_20226,N_17185,N_17417);
and U20227 (N_20227,N_16213,N_15670);
or U20228 (N_20228,N_17495,N_16359);
nor U20229 (N_20229,N_17294,N_16304);
xnor U20230 (N_20230,N_15581,N_17541);
xnor U20231 (N_20231,N_17816,N_15850);
or U20232 (N_20232,N_16447,N_16115);
nand U20233 (N_20233,N_17680,N_15978);
and U20234 (N_20234,N_16618,N_17126);
and U20235 (N_20235,N_15813,N_17611);
and U20236 (N_20236,N_16316,N_17654);
or U20237 (N_20237,N_17238,N_16736);
nand U20238 (N_20238,N_15679,N_16556);
nor U20239 (N_20239,N_16200,N_17169);
xnor U20240 (N_20240,N_17765,N_17141);
nand U20241 (N_20241,N_16710,N_16807);
nand U20242 (N_20242,N_15603,N_17755);
nor U20243 (N_20243,N_15956,N_15246);
nand U20244 (N_20244,N_17400,N_15344);
and U20245 (N_20245,N_15347,N_16332);
or U20246 (N_20246,N_15120,N_15973);
or U20247 (N_20247,N_17468,N_15037);
nor U20248 (N_20248,N_17675,N_16181);
or U20249 (N_20249,N_16743,N_15331);
or U20250 (N_20250,N_15965,N_15295);
and U20251 (N_20251,N_17228,N_17226);
and U20252 (N_20252,N_15252,N_15899);
or U20253 (N_20253,N_17140,N_16704);
nand U20254 (N_20254,N_16440,N_15901);
and U20255 (N_20255,N_17019,N_15565);
nor U20256 (N_20256,N_17271,N_17935);
nand U20257 (N_20257,N_15735,N_15053);
and U20258 (N_20258,N_16562,N_16429);
and U20259 (N_20259,N_15498,N_16212);
xor U20260 (N_20260,N_15381,N_17512);
or U20261 (N_20261,N_15818,N_15582);
nor U20262 (N_20262,N_17910,N_16975);
or U20263 (N_20263,N_15895,N_15996);
nand U20264 (N_20264,N_16852,N_17739);
xnor U20265 (N_20265,N_15352,N_15921);
and U20266 (N_20266,N_16018,N_15449);
nor U20267 (N_20267,N_15237,N_15544);
and U20268 (N_20268,N_17999,N_16788);
nor U20269 (N_20269,N_17503,N_16058);
nor U20270 (N_20270,N_17560,N_17153);
or U20271 (N_20271,N_15281,N_17524);
xor U20272 (N_20272,N_17804,N_16601);
xor U20273 (N_20273,N_15177,N_17517);
xnor U20274 (N_20274,N_17659,N_16362);
nor U20275 (N_20275,N_17507,N_16650);
and U20276 (N_20276,N_16992,N_17503);
or U20277 (N_20277,N_15683,N_17579);
or U20278 (N_20278,N_16358,N_17802);
nor U20279 (N_20279,N_16951,N_17710);
xnor U20280 (N_20280,N_17853,N_16569);
xnor U20281 (N_20281,N_16127,N_16524);
nand U20282 (N_20282,N_16764,N_15774);
and U20283 (N_20283,N_16601,N_17441);
nand U20284 (N_20284,N_15670,N_17169);
xor U20285 (N_20285,N_15007,N_15072);
nor U20286 (N_20286,N_17305,N_15170);
nand U20287 (N_20287,N_17571,N_17740);
and U20288 (N_20288,N_16586,N_16309);
nand U20289 (N_20289,N_16693,N_17456);
nand U20290 (N_20290,N_15863,N_17173);
or U20291 (N_20291,N_17722,N_16825);
nand U20292 (N_20292,N_15013,N_15437);
nand U20293 (N_20293,N_16054,N_16502);
nand U20294 (N_20294,N_15290,N_17424);
nor U20295 (N_20295,N_15575,N_15480);
nor U20296 (N_20296,N_17919,N_16905);
and U20297 (N_20297,N_17222,N_15532);
xnor U20298 (N_20298,N_15371,N_17379);
nor U20299 (N_20299,N_16470,N_17048);
or U20300 (N_20300,N_15509,N_15900);
nand U20301 (N_20301,N_16483,N_16117);
xor U20302 (N_20302,N_17081,N_17004);
and U20303 (N_20303,N_16807,N_17242);
nor U20304 (N_20304,N_15045,N_16998);
or U20305 (N_20305,N_17555,N_15931);
or U20306 (N_20306,N_17831,N_15338);
nor U20307 (N_20307,N_16722,N_15541);
nand U20308 (N_20308,N_17302,N_16673);
nand U20309 (N_20309,N_17666,N_17618);
or U20310 (N_20310,N_15268,N_16049);
nor U20311 (N_20311,N_17636,N_17904);
and U20312 (N_20312,N_16574,N_16478);
nand U20313 (N_20313,N_17631,N_16323);
xnor U20314 (N_20314,N_17391,N_15396);
or U20315 (N_20315,N_15834,N_17260);
or U20316 (N_20316,N_15136,N_15882);
and U20317 (N_20317,N_15317,N_16922);
or U20318 (N_20318,N_16415,N_17716);
nor U20319 (N_20319,N_15405,N_15673);
nor U20320 (N_20320,N_16880,N_16849);
xor U20321 (N_20321,N_17984,N_17204);
or U20322 (N_20322,N_16763,N_17847);
xnor U20323 (N_20323,N_16113,N_17392);
xnor U20324 (N_20324,N_16270,N_17129);
or U20325 (N_20325,N_15393,N_17030);
and U20326 (N_20326,N_16538,N_15046);
or U20327 (N_20327,N_17404,N_17935);
or U20328 (N_20328,N_15387,N_15224);
nor U20329 (N_20329,N_16467,N_15896);
nor U20330 (N_20330,N_16654,N_16857);
nand U20331 (N_20331,N_17065,N_15935);
xnor U20332 (N_20332,N_17067,N_15833);
nor U20333 (N_20333,N_15185,N_16489);
nand U20334 (N_20334,N_16461,N_16922);
xor U20335 (N_20335,N_16098,N_17169);
nor U20336 (N_20336,N_16328,N_17231);
and U20337 (N_20337,N_15648,N_15208);
or U20338 (N_20338,N_17268,N_16277);
xor U20339 (N_20339,N_16334,N_17253);
nor U20340 (N_20340,N_16303,N_17296);
xnor U20341 (N_20341,N_17741,N_15029);
or U20342 (N_20342,N_16415,N_15221);
nor U20343 (N_20343,N_16024,N_15059);
or U20344 (N_20344,N_16865,N_16678);
and U20345 (N_20345,N_17196,N_15705);
nor U20346 (N_20346,N_17370,N_15286);
or U20347 (N_20347,N_16298,N_15307);
xnor U20348 (N_20348,N_17974,N_16424);
or U20349 (N_20349,N_16874,N_17571);
nor U20350 (N_20350,N_15174,N_17442);
nor U20351 (N_20351,N_15511,N_17539);
nor U20352 (N_20352,N_17225,N_17346);
and U20353 (N_20353,N_17146,N_17668);
xor U20354 (N_20354,N_15847,N_17092);
nand U20355 (N_20355,N_17870,N_16562);
xor U20356 (N_20356,N_17345,N_16999);
nand U20357 (N_20357,N_15246,N_17413);
and U20358 (N_20358,N_17428,N_17191);
and U20359 (N_20359,N_17464,N_15986);
xor U20360 (N_20360,N_16281,N_17752);
nand U20361 (N_20361,N_15646,N_15477);
xnor U20362 (N_20362,N_16202,N_16055);
nor U20363 (N_20363,N_17354,N_15675);
nand U20364 (N_20364,N_15382,N_15193);
xnor U20365 (N_20365,N_17169,N_16011);
nand U20366 (N_20366,N_15700,N_15668);
nand U20367 (N_20367,N_15886,N_16366);
or U20368 (N_20368,N_17362,N_15059);
and U20369 (N_20369,N_15791,N_16353);
nor U20370 (N_20370,N_15329,N_16518);
nor U20371 (N_20371,N_15274,N_16372);
nand U20372 (N_20372,N_17575,N_15194);
or U20373 (N_20373,N_15340,N_15662);
nor U20374 (N_20374,N_15757,N_17783);
or U20375 (N_20375,N_17313,N_16083);
nor U20376 (N_20376,N_17237,N_17420);
nor U20377 (N_20377,N_16740,N_16329);
and U20378 (N_20378,N_15355,N_15216);
or U20379 (N_20379,N_15285,N_17044);
nor U20380 (N_20380,N_16690,N_17607);
or U20381 (N_20381,N_15278,N_17701);
nand U20382 (N_20382,N_16963,N_16837);
xnor U20383 (N_20383,N_16757,N_17144);
nand U20384 (N_20384,N_17119,N_17518);
nor U20385 (N_20385,N_15859,N_16673);
nand U20386 (N_20386,N_15033,N_15248);
and U20387 (N_20387,N_16322,N_16801);
and U20388 (N_20388,N_16959,N_17790);
and U20389 (N_20389,N_16636,N_15961);
or U20390 (N_20390,N_15594,N_16921);
nand U20391 (N_20391,N_17955,N_16993);
and U20392 (N_20392,N_15188,N_16321);
xnor U20393 (N_20393,N_17844,N_15412);
and U20394 (N_20394,N_17098,N_16111);
and U20395 (N_20395,N_16639,N_17886);
or U20396 (N_20396,N_17198,N_15593);
xor U20397 (N_20397,N_17864,N_15220);
or U20398 (N_20398,N_16136,N_15432);
nand U20399 (N_20399,N_15230,N_17742);
or U20400 (N_20400,N_15368,N_17568);
nor U20401 (N_20401,N_17869,N_17438);
or U20402 (N_20402,N_16152,N_16779);
nand U20403 (N_20403,N_16714,N_16369);
and U20404 (N_20404,N_16811,N_17410);
and U20405 (N_20405,N_15477,N_15403);
xor U20406 (N_20406,N_16060,N_16272);
or U20407 (N_20407,N_16005,N_17077);
or U20408 (N_20408,N_17518,N_17578);
nand U20409 (N_20409,N_17463,N_17684);
xor U20410 (N_20410,N_16090,N_16291);
and U20411 (N_20411,N_16348,N_17341);
nor U20412 (N_20412,N_15373,N_17719);
nor U20413 (N_20413,N_17340,N_16142);
xor U20414 (N_20414,N_15987,N_17849);
and U20415 (N_20415,N_16622,N_16708);
nand U20416 (N_20416,N_16982,N_16120);
and U20417 (N_20417,N_15176,N_15944);
nand U20418 (N_20418,N_17679,N_15035);
xor U20419 (N_20419,N_15817,N_15244);
or U20420 (N_20420,N_15109,N_15332);
xnor U20421 (N_20421,N_15492,N_17111);
xor U20422 (N_20422,N_16237,N_15821);
nor U20423 (N_20423,N_16043,N_16471);
nor U20424 (N_20424,N_15598,N_17019);
nor U20425 (N_20425,N_16946,N_16914);
nor U20426 (N_20426,N_15208,N_15679);
nor U20427 (N_20427,N_16613,N_15197);
or U20428 (N_20428,N_15569,N_17646);
nor U20429 (N_20429,N_15732,N_16546);
and U20430 (N_20430,N_17687,N_17331);
and U20431 (N_20431,N_17204,N_16957);
and U20432 (N_20432,N_15929,N_17999);
nor U20433 (N_20433,N_16395,N_15393);
xnor U20434 (N_20434,N_16275,N_17340);
xnor U20435 (N_20435,N_17932,N_17968);
nor U20436 (N_20436,N_17195,N_16539);
xnor U20437 (N_20437,N_15254,N_15127);
xnor U20438 (N_20438,N_16933,N_17338);
nand U20439 (N_20439,N_17261,N_17410);
nand U20440 (N_20440,N_15987,N_16937);
or U20441 (N_20441,N_17279,N_17804);
xnor U20442 (N_20442,N_15884,N_17708);
xnor U20443 (N_20443,N_16871,N_15968);
xnor U20444 (N_20444,N_15672,N_15542);
nand U20445 (N_20445,N_16383,N_15227);
nor U20446 (N_20446,N_17423,N_15393);
xor U20447 (N_20447,N_15889,N_15895);
nand U20448 (N_20448,N_17147,N_16627);
nand U20449 (N_20449,N_15694,N_17118);
or U20450 (N_20450,N_16194,N_15101);
or U20451 (N_20451,N_17855,N_15733);
and U20452 (N_20452,N_16951,N_16598);
nor U20453 (N_20453,N_16511,N_15642);
nor U20454 (N_20454,N_15660,N_17251);
nor U20455 (N_20455,N_15382,N_16890);
xnor U20456 (N_20456,N_15393,N_15059);
nor U20457 (N_20457,N_16962,N_17367);
nand U20458 (N_20458,N_16583,N_17755);
nand U20459 (N_20459,N_15906,N_17573);
nand U20460 (N_20460,N_16567,N_17220);
and U20461 (N_20461,N_16184,N_17365);
xnor U20462 (N_20462,N_17163,N_17705);
nor U20463 (N_20463,N_15750,N_16254);
nor U20464 (N_20464,N_15205,N_15336);
or U20465 (N_20465,N_16249,N_16887);
xor U20466 (N_20466,N_16148,N_15795);
xnor U20467 (N_20467,N_16429,N_17987);
nand U20468 (N_20468,N_16908,N_17096);
nand U20469 (N_20469,N_15007,N_15539);
nand U20470 (N_20470,N_15835,N_15679);
or U20471 (N_20471,N_17470,N_15068);
nand U20472 (N_20472,N_17101,N_15377);
nor U20473 (N_20473,N_15204,N_15462);
nand U20474 (N_20474,N_17824,N_16889);
xnor U20475 (N_20475,N_15419,N_16566);
xor U20476 (N_20476,N_15783,N_16940);
nand U20477 (N_20477,N_16941,N_16298);
nand U20478 (N_20478,N_15057,N_16432);
and U20479 (N_20479,N_17553,N_17445);
and U20480 (N_20480,N_17842,N_16293);
xor U20481 (N_20481,N_17743,N_15834);
and U20482 (N_20482,N_16321,N_16111);
nand U20483 (N_20483,N_15636,N_17734);
nand U20484 (N_20484,N_15018,N_16201);
xnor U20485 (N_20485,N_16589,N_16305);
nand U20486 (N_20486,N_16484,N_17746);
nand U20487 (N_20487,N_17809,N_17341);
nand U20488 (N_20488,N_15744,N_15040);
nor U20489 (N_20489,N_17906,N_16544);
or U20490 (N_20490,N_16483,N_15166);
nor U20491 (N_20491,N_15550,N_17777);
nand U20492 (N_20492,N_17615,N_15408);
nor U20493 (N_20493,N_15919,N_17923);
and U20494 (N_20494,N_17831,N_15529);
xor U20495 (N_20495,N_17436,N_15915);
nand U20496 (N_20496,N_17799,N_16002);
and U20497 (N_20497,N_15323,N_16411);
nor U20498 (N_20498,N_15185,N_15578);
xor U20499 (N_20499,N_17617,N_17267);
nor U20500 (N_20500,N_16107,N_15728);
or U20501 (N_20501,N_15465,N_16061);
and U20502 (N_20502,N_16586,N_15832);
nor U20503 (N_20503,N_17841,N_17358);
or U20504 (N_20504,N_15255,N_17885);
nand U20505 (N_20505,N_15418,N_16214);
xnor U20506 (N_20506,N_15339,N_17241);
xnor U20507 (N_20507,N_16120,N_17252);
nor U20508 (N_20508,N_16405,N_17121);
xnor U20509 (N_20509,N_17337,N_15399);
and U20510 (N_20510,N_15797,N_16950);
and U20511 (N_20511,N_17631,N_15813);
nor U20512 (N_20512,N_16680,N_15400);
and U20513 (N_20513,N_15671,N_17554);
nand U20514 (N_20514,N_16601,N_17766);
nand U20515 (N_20515,N_17757,N_15447);
xnor U20516 (N_20516,N_16211,N_15162);
nor U20517 (N_20517,N_17357,N_15775);
nor U20518 (N_20518,N_16905,N_16646);
xor U20519 (N_20519,N_15512,N_17418);
or U20520 (N_20520,N_17008,N_17552);
or U20521 (N_20521,N_17476,N_15273);
or U20522 (N_20522,N_15147,N_17081);
or U20523 (N_20523,N_17577,N_15143);
and U20524 (N_20524,N_17042,N_15712);
nand U20525 (N_20525,N_15076,N_16094);
and U20526 (N_20526,N_16853,N_17956);
or U20527 (N_20527,N_15951,N_17601);
nand U20528 (N_20528,N_16292,N_17748);
nand U20529 (N_20529,N_16971,N_16977);
nor U20530 (N_20530,N_17943,N_17434);
and U20531 (N_20531,N_17967,N_16096);
or U20532 (N_20532,N_17514,N_17553);
nand U20533 (N_20533,N_17437,N_15871);
or U20534 (N_20534,N_17272,N_17961);
xor U20535 (N_20535,N_16271,N_17801);
and U20536 (N_20536,N_17794,N_16420);
and U20537 (N_20537,N_15066,N_16475);
and U20538 (N_20538,N_16145,N_16582);
and U20539 (N_20539,N_15292,N_17587);
nor U20540 (N_20540,N_17335,N_16886);
and U20541 (N_20541,N_16611,N_17627);
nand U20542 (N_20542,N_17433,N_15030);
xor U20543 (N_20543,N_16267,N_15580);
and U20544 (N_20544,N_15463,N_17502);
nand U20545 (N_20545,N_16159,N_17543);
or U20546 (N_20546,N_16616,N_17544);
nor U20547 (N_20547,N_17293,N_15887);
and U20548 (N_20548,N_15291,N_15404);
xnor U20549 (N_20549,N_15862,N_15078);
or U20550 (N_20550,N_17201,N_16706);
or U20551 (N_20551,N_16267,N_15674);
and U20552 (N_20552,N_15974,N_17440);
nand U20553 (N_20553,N_15701,N_17067);
xnor U20554 (N_20554,N_16665,N_16442);
nor U20555 (N_20555,N_17119,N_15794);
and U20556 (N_20556,N_17032,N_17160);
xor U20557 (N_20557,N_16750,N_17997);
nand U20558 (N_20558,N_17448,N_15964);
xor U20559 (N_20559,N_17551,N_17306);
nand U20560 (N_20560,N_15231,N_16366);
xnor U20561 (N_20561,N_16804,N_16108);
and U20562 (N_20562,N_16892,N_16524);
xor U20563 (N_20563,N_17740,N_15226);
and U20564 (N_20564,N_17959,N_15930);
nand U20565 (N_20565,N_15062,N_17269);
xor U20566 (N_20566,N_16488,N_15246);
and U20567 (N_20567,N_17688,N_15544);
nor U20568 (N_20568,N_15498,N_17567);
or U20569 (N_20569,N_16405,N_17848);
xnor U20570 (N_20570,N_17439,N_16919);
nand U20571 (N_20571,N_15983,N_16716);
xor U20572 (N_20572,N_15876,N_16251);
and U20573 (N_20573,N_16410,N_15754);
or U20574 (N_20574,N_16031,N_15687);
nand U20575 (N_20575,N_15991,N_16303);
or U20576 (N_20576,N_15764,N_16199);
and U20577 (N_20577,N_16742,N_16462);
and U20578 (N_20578,N_17155,N_17848);
nor U20579 (N_20579,N_15914,N_17531);
or U20580 (N_20580,N_16056,N_16128);
nand U20581 (N_20581,N_17866,N_17969);
nand U20582 (N_20582,N_16733,N_16490);
xor U20583 (N_20583,N_15644,N_16998);
nor U20584 (N_20584,N_15956,N_17398);
nand U20585 (N_20585,N_16326,N_15497);
nand U20586 (N_20586,N_17824,N_15912);
and U20587 (N_20587,N_16899,N_17253);
nor U20588 (N_20588,N_16090,N_17089);
xnor U20589 (N_20589,N_16283,N_17396);
xnor U20590 (N_20590,N_16666,N_17226);
nor U20591 (N_20591,N_16313,N_17385);
nor U20592 (N_20592,N_15733,N_15184);
nor U20593 (N_20593,N_17696,N_16990);
or U20594 (N_20594,N_15587,N_15684);
nor U20595 (N_20595,N_17634,N_15640);
or U20596 (N_20596,N_17146,N_17774);
and U20597 (N_20597,N_17140,N_17892);
nand U20598 (N_20598,N_17357,N_16839);
or U20599 (N_20599,N_15991,N_17459);
and U20600 (N_20600,N_16953,N_17878);
or U20601 (N_20601,N_17064,N_16931);
or U20602 (N_20602,N_17443,N_15108);
xor U20603 (N_20603,N_15475,N_17609);
or U20604 (N_20604,N_17766,N_16291);
nor U20605 (N_20605,N_15755,N_17707);
xnor U20606 (N_20606,N_15530,N_16642);
or U20607 (N_20607,N_15557,N_17012);
or U20608 (N_20608,N_17755,N_17201);
or U20609 (N_20609,N_17254,N_15450);
or U20610 (N_20610,N_16552,N_16485);
or U20611 (N_20611,N_16028,N_17088);
nor U20612 (N_20612,N_17454,N_15551);
nor U20613 (N_20613,N_16408,N_15374);
or U20614 (N_20614,N_16433,N_17014);
or U20615 (N_20615,N_15429,N_17754);
nor U20616 (N_20616,N_16971,N_17766);
and U20617 (N_20617,N_17013,N_16059);
or U20618 (N_20618,N_15955,N_15094);
nand U20619 (N_20619,N_16037,N_17816);
nand U20620 (N_20620,N_16246,N_16758);
nor U20621 (N_20621,N_17918,N_15465);
or U20622 (N_20622,N_15059,N_15753);
xor U20623 (N_20623,N_15343,N_16379);
and U20624 (N_20624,N_16079,N_15482);
xnor U20625 (N_20625,N_16904,N_16540);
nand U20626 (N_20626,N_16506,N_17886);
or U20627 (N_20627,N_16729,N_17003);
or U20628 (N_20628,N_15067,N_16080);
nor U20629 (N_20629,N_16164,N_16487);
xor U20630 (N_20630,N_17176,N_16325);
xnor U20631 (N_20631,N_15854,N_16241);
nand U20632 (N_20632,N_15924,N_17559);
nor U20633 (N_20633,N_16455,N_15003);
nand U20634 (N_20634,N_15112,N_17138);
or U20635 (N_20635,N_16649,N_17682);
and U20636 (N_20636,N_17534,N_16801);
nand U20637 (N_20637,N_16945,N_17354);
and U20638 (N_20638,N_17494,N_17225);
xor U20639 (N_20639,N_15682,N_15293);
or U20640 (N_20640,N_17440,N_15202);
or U20641 (N_20641,N_15210,N_17322);
or U20642 (N_20642,N_16533,N_17912);
xnor U20643 (N_20643,N_17432,N_16411);
nor U20644 (N_20644,N_15580,N_17500);
and U20645 (N_20645,N_15146,N_16708);
and U20646 (N_20646,N_17105,N_15059);
and U20647 (N_20647,N_15834,N_17110);
nor U20648 (N_20648,N_15781,N_16378);
xnor U20649 (N_20649,N_16140,N_17251);
nor U20650 (N_20650,N_17957,N_15565);
or U20651 (N_20651,N_17625,N_15792);
nand U20652 (N_20652,N_17432,N_16197);
xnor U20653 (N_20653,N_16374,N_15480);
and U20654 (N_20654,N_15678,N_15592);
xor U20655 (N_20655,N_15772,N_17101);
nor U20656 (N_20656,N_16793,N_15776);
nand U20657 (N_20657,N_17274,N_15346);
nand U20658 (N_20658,N_17935,N_17172);
xnor U20659 (N_20659,N_16673,N_17404);
xnor U20660 (N_20660,N_16021,N_16437);
or U20661 (N_20661,N_16012,N_17595);
nand U20662 (N_20662,N_17343,N_15759);
nor U20663 (N_20663,N_15572,N_15751);
xor U20664 (N_20664,N_16913,N_17964);
nand U20665 (N_20665,N_17545,N_17141);
xnor U20666 (N_20666,N_15762,N_17962);
nand U20667 (N_20667,N_15645,N_15404);
xnor U20668 (N_20668,N_17695,N_16203);
nand U20669 (N_20669,N_16688,N_15073);
xor U20670 (N_20670,N_16589,N_16189);
or U20671 (N_20671,N_15461,N_15639);
and U20672 (N_20672,N_17746,N_16595);
nand U20673 (N_20673,N_17639,N_15052);
nand U20674 (N_20674,N_17633,N_16012);
xnor U20675 (N_20675,N_15913,N_16318);
and U20676 (N_20676,N_16255,N_15409);
xor U20677 (N_20677,N_17594,N_15774);
or U20678 (N_20678,N_17201,N_17059);
xnor U20679 (N_20679,N_17915,N_17407);
xnor U20680 (N_20680,N_15912,N_16029);
nand U20681 (N_20681,N_16542,N_16681);
nor U20682 (N_20682,N_17021,N_15513);
and U20683 (N_20683,N_15461,N_16070);
or U20684 (N_20684,N_17218,N_15340);
or U20685 (N_20685,N_15871,N_17768);
xor U20686 (N_20686,N_15291,N_17059);
nor U20687 (N_20687,N_15274,N_16740);
nand U20688 (N_20688,N_17492,N_16917);
or U20689 (N_20689,N_15965,N_15562);
nor U20690 (N_20690,N_16220,N_17223);
and U20691 (N_20691,N_15950,N_15255);
and U20692 (N_20692,N_15844,N_15536);
or U20693 (N_20693,N_16051,N_17510);
xor U20694 (N_20694,N_15003,N_16973);
nand U20695 (N_20695,N_15962,N_15602);
nor U20696 (N_20696,N_17326,N_15850);
and U20697 (N_20697,N_17122,N_17574);
nor U20698 (N_20698,N_16577,N_15895);
or U20699 (N_20699,N_15742,N_15344);
nor U20700 (N_20700,N_15283,N_16553);
nor U20701 (N_20701,N_15665,N_15334);
or U20702 (N_20702,N_17963,N_16799);
nor U20703 (N_20703,N_16906,N_16506);
xor U20704 (N_20704,N_16464,N_17521);
nor U20705 (N_20705,N_16047,N_15757);
nor U20706 (N_20706,N_15075,N_16315);
or U20707 (N_20707,N_17532,N_17275);
nand U20708 (N_20708,N_16642,N_17180);
nand U20709 (N_20709,N_16635,N_17411);
xor U20710 (N_20710,N_17169,N_17084);
nand U20711 (N_20711,N_16376,N_15787);
or U20712 (N_20712,N_16459,N_17990);
xnor U20713 (N_20713,N_17588,N_15652);
nand U20714 (N_20714,N_17434,N_17124);
nand U20715 (N_20715,N_16160,N_15685);
or U20716 (N_20716,N_15307,N_17271);
or U20717 (N_20717,N_17489,N_16729);
nand U20718 (N_20718,N_15008,N_16109);
nor U20719 (N_20719,N_16659,N_16931);
nor U20720 (N_20720,N_17861,N_17538);
and U20721 (N_20721,N_17558,N_16811);
and U20722 (N_20722,N_16846,N_17101);
or U20723 (N_20723,N_15957,N_16312);
or U20724 (N_20724,N_17079,N_17136);
or U20725 (N_20725,N_16744,N_15435);
nand U20726 (N_20726,N_16650,N_15461);
and U20727 (N_20727,N_16913,N_15318);
and U20728 (N_20728,N_15740,N_17759);
and U20729 (N_20729,N_15777,N_17804);
nand U20730 (N_20730,N_16649,N_16885);
nor U20731 (N_20731,N_17395,N_15456);
xor U20732 (N_20732,N_17790,N_16632);
xnor U20733 (N_20733,N_16985,N_15490);
nand U20734 (N_20734,N_16868,N_15713);
or U20735 (N_20735,N_15941,N_15751);
xnor U20736 (N_20736,N_15156,N_16546);
and U20737 (N_20737,N_15925,N_15257);
nor U20738 (N_20738,N_16121,N_17097);
xor U20739 (N_20739,N_15854,N_16132);
nor U20740 (N_20740,N_17428,N_16926);
nor U20741 (N_20741,N_15925,N_17293);
nor U20742 (N_20742,N_15537,N_17152);
or U20743 (N_20743,N_15748,N_17109);
nor U20744 (N_20744,N_16494,N_16817);
nand U20745 (N_20745,N_17026,N_17209);
and U20746 (N_20746,N_15385,N_16619);
nand U20747 (N_20747,N_16375,N_16522);
nor U20748 (N_20748,N_16399,N_17010);
or U20749 (N_20749,N_15526,N_16803);
and U20750 (N_20750,N_17183,N_17077);
and U20751 (N_20751,N_15418,N_17187);
nor U20752 (N_20752,N_15086,N_15255);
xnor U20753 (N_20753,N_17438,N_15914);
nand U20754 (N_20754,N_17937,N_15294);
and U20755 (N_20755,N_16051,N_15759);
or U20756 (N_20756,N_15476,N_17573);
nand U20757 (N_20757,N_16909,N_15357);
nand U20758 (N_20758,N_15707,N_16055);
nand U20759 (N_20759,N_16862,N_15399);
xnor U20760 (N_20760,N_17368,N_16054);
and U20761 (N_20761,N_15407,N_17736);
or U20762 (N_20762,N_17525,N_17673);
and U20763 (N_20763,N_16046,N_15494);
xnor U20764 (N_20764,N_16454,N_15340);
and U20765 (N_20765,N_16850,N_16926);
nand U20766 (N_20766,N_16781,N_15775);
and U20767 (N_20767,N_17867,N_17810);
and U20768 (N_20768,N_16524,N_17782);
xor U20769 (N_20769,N_17072,N_16280);
xor U20770 (N_20770,N_17139,N_16270);
nand U20771 (N_20771,N_15689,N_17611);
nor U20772 (N_20772,N_16946,N_16792);
nand U20773 (N_20773,N_16789,N_16953);
and U20774 (N_20774,N_16804,N_17678);
nand U20775 (N_20775,N_15425,N_15393);
nor U20776 (N_20776,N_15696,N_17392);
nor U20777 (N_20777,N_16974,N_15885);
xnor U20778 (N_20778,N_15092,N_16462);
xnor U20779 (N_20779,N_17068,N_16352);
xnor U20780 (N_20780,N_15603,N_15033);
xor U20781 (N_20781,N_16414,N_17606);
nor U20782 (N_20782,N_15071,N_16303);
or U20783 (N_20783,N_16413,N_16825);
and U20784 (N_20784,N_17749,N_15530);
nor U20785 (N_20785,N_15887,N_15561);
nand U20786 (N_20786,N_17308,N_16474);
or U20787 (N_20787,N_15837,N_16326);
and U20788 (N_20788,N_15364,N_15175);
nand U20789 (N_20789,N_17364,N_17542);
and U20790 (N_20790,N_17357,N_17723);
nor U20791 (N_20791,N_17621,N_16380);
and U20792 (N_20792,N_16692,N_17471);
or U20793 (N_20793,N_16293,N_16391);
nand U20794 (N_20794,N_15804,N_16845);
nand U20795 (N_20795,N_17057,N_17445);
nor U20796 (N_20796,N_16337,N_16980);
nand U20797 (N_20797,N_16862,N_17643);
nor U20798 (N_20798,N_15790,N_15914);
and U20799 (N_20799,N_15290,N_15795);
nand U20800 (N_20800,N_16151,N_15989);
and U20801 (N_20801,N_17092,N_15472);
or U20802 (N_20802,N_17936,N_16344);
xnor U20803 (N_20803,N_16726,N_16764);
nand U20804 (N_20804,N_16957,N_17931);
or U20805 (N_20805,N_17032,N_16388);
nor U20806 (N_20806,N_16430,N_15547);
or U20807 (N_20807,N_17584,N_17129);
nor U20808 (N_20808,N_15777,N_16032);
nand U20809 (N_20809,N_16980,N_15666);
xnor U20810 (N_20810,N_16551,N_16400);
or U20811 (N_20811,N_17573,N_17153);
nand U20812 (N_20812,N_15407,N_17807);
xnor U20813 (N_20813,N_15213,N_17417);
nand U20814 (N_20814,N_17478,N_15499);
or U20815 (N_20815,N_16165,N_17432);
nor U20816 (N_20816,N_15183,N_15523);
or U20817 (N_20817,N_15396,N_17292);
nand U20818 (N_20818,N_17621,N_15674);
and U20819 (N_20819,N_17035,N_15291);
nand U20820 (N_20820,N_17456,N_17041);
nor U20821 (N_20821,N_16374,N_16988);
nand U20822 (N_20822,N_15873,N_15370);
or U20823 (N_20823,N_15038,N_17087);
or U20824 (N_20824,N_16459,N_15642);
or U20825 (N_20825,N_16999,N_15787);
and U20826 (N_20826,N_17139,N_15085);
or U20827 (N_20827,N_15318,N_17807);
or U20828 (N_20828,N_15451,N_15769);
and U20829 (N_20829,N_17338,N_15338);
or U20830 (N_20830,N_16820,N_15223);
nor U20831 (N_20831,N_15591,N_16579);
or U20832 (N_20832,N_15056,N_16473);
nand U20833 (N_20833,N_16452,N_17470);
or U20834 (N_20834,N_15044,N_16269);
nand U20835 (N_20835,N_15999,N_16113);
and U20836 (N_20836,N_15953,N_16204);
nor U20837 (N_20837,N_16539,N_15265);
and U20838 (N_20838,N_15452,N_16133);
nor U20839 (N_20839,N_16976,N_16127);
xnor U20840 (N_20840,N_15331,N_17565);
nand U20841 (N_20841,N_16247,N_17761);
nor U20842 (N_20842,N_17362,N_15310);
nand U20843 (N_20843,N_16296,N_16408);
nand U20844 (N_20844,N_16462,N_17336);
xor U20845 (N_20845,N_16206,N_15338);
or U20846 (N_20846,N_15528,N_15015);
xnor U20847 (N_20847,N_17942,N_17205);
nand U20848 (N_20848,N_16561,N_17795);
nand U20849 (N_20849,N_15200,N_16737);
nand U20850 (N_20850,N_15844,N_17185);
and U20851 (N_20851,N_16234,N_16553);
nor U20852 (N_20852,N_16947,N_16398);
xnor U20853 (N_20853,N_17278,N_16195);
and U20854 (N_20854,N_15665,N_16942);
nor U20855 (N_20855,N_15486,N_15576);
nand U20856 (N_20856,N_16156,N_17940);
nand U20857 (N_20857,N_15951,N_17206);
nor U20858 (N_20858,N_15168,N_15459);
nand U20859 (N_20859,N_17585,N_15426);
nor U20860 (N_20860,N_15119,N_15948);
xor U20861 (N_20861,N_15730,N_17221);
nor U20862 (N_20862,N_17900,N_16291);
or U20863 (N_20863,N_16974,N_16355);
xor U20864 (N_20864,N_15306,N_15822);
nor U20865 (N_20865,N_17512,N_15538);
nor U20866 (N_20866,N_16596,N_15105);
or U20867 (N_20867,N_15924,N_16228);
or U20868 (N_20868,N_15511,N_15583);
xor U20869 (N_20869,N_16810,N_16793);
nand U20870 (N_20870,N_16762,N_15787);
and U20871 (N_20871,N_15327,N_15069);
and U20872 (N_20872,N_15431,N_17887);
nor U20873 (N_20873,N_17011,N_15838);
xor U20874 (N_20874,N_17371,N_15524);
nand U20875 (N_20875,N_16236,N_16148);
nand U20876 (N_20876,N_17987,N_17274);
xnor U20877 (N_20877,N_17496,N_15892);
xnor U20878 (N_20878,N_17490,N_17547);
nor U20879 (N_20879,N_17281,N_16673);
and U20880 (N_20880,N_17147,N_15219);
nand U20881 (N_20881,N_16962,N_17993);
or U20882 (N_20882,N_17231,N_15176);
nand U20883 (N_20883,N_15428,N_17882);
and U20884 (N_20884,N_17635,N_16437);
or U20885 (N_20885,N_16499,N_15749);
nor U20886 (N_20886,N_15779,N_17100);
xnor U20887 (N_20887,N_16371,N_16735);
or U20888 (N_20888,N_16872,N_17376);
or U20889 (N_20889,N_16108,N_17407);
nand U20890 (N_20890,N_15674,N_17821);
nor U20891 (N_20891,N_16273,N_16329);
and U20892 (N_20892,N_15288,N_17262);
nand U20893 (N_20893,N_16531,N_15166);
nor U20894 (N_20894,N_17691,N_15248);
xor U20895 (N_20895,N_17406,N_16542);
nand U20896 (N_20896,N_16527,N_15821);
xnor U20897 (N_20897,N_15445,N_15168);
nor U20898 (N_20898,N_15665,N_15810);
xor U20899 (N_20899,N_15405,N_17641);
and U20900 (N_20900,N_16778,N_15959);
nand U20901 (N_20901,N_15389,N_16242);
or U20902 (N_20902,N_15655,N_15199);
or U20903 (N_20903,N_15368,N_16626);
or U20904 (N_20904,N_15681,N_17277);
xor U20905 (N_20905,N_15326,N_17922);
xor U20906 (N_20906,N_15164,N_17763);
and U20907 (N_20907,N_16200,N_17253);
or U20908 (N_20908,N_17684,N_17090);
nand U20909 (N_20909,N_15433,N_15967);
or U20910 (N_20910,N_15571,N_17886);
xor U20911 (N_20911,N_16947,N_16433);
nand U20912 (N_20912,N_16418,N_15262);
xnor U20913 (N_20913,N_16847,N_15628);
xnor U20914 (N_20914,N_16669,N_15291);
or U20915 (N_20915,N_17439,N_16923);
nand U20916 (N_20916,N_16475,N_15248);
or U20917 (N_20917,N_15398,N_17354);
nand U20918 (N_20918,N_16601,N_15921);
xor U20919 (N_20919,N_17772,N_17301);
nor U20920 (N_20920,N_16308,N_15916);
nor U20921 (N_20921,N_15513,N_15976);
xnor U20922 (N_20922,N_16557,N_16869);
nor U20923 (N_20923,N_16034,N_15208);
xor U20924 (N_20924,N_17832,N_17157);
nand U20925 (N_20925,N_16091,N_15577);
xor U20926 (N_20926,N_15897,N_16255);
nand U20927 (N_20927,N_15016,N_16148);
and U20928 (N_20928,N_17825,N_15116);
nor U20929 (N_20929,N_16037,N_16507);
nand U20930 (N_20930,N_16990,N_16104);
or U20931 (N_20931,N_15507,N_16520);
xor U20932 (N_20932,N_17330,N_16106);
nand U20933 (N_20933,N_17131,N_17139);
nand U20934 (N_20934,N_15368,N_17780);
or U20935 (N_20935,N_16449,N_17904);
nand U20936 (N_20936,N_15580,N_15336);
xor U20937 (N_20937,N_15666,N_17529);
nor U20938 (N_20938,N_17170,N_15727);
or U20939 (N_20939,N_16538,N_15666);
or U20940 (N_20940,N_16144,N_15114);
nand U20941 (N_20941,N_17503,N_15913);
nand U20942 (N_20942,N_15924,N_15733);
and U20943 (N_20943,N_16092,N_17201);
or U20944 (N_20944,N_17243,N_16721);
xor U20945 (N_20945,N_16705,N_15608);
nor U20946 (N_20946,N_16061,N_16284);
and U20947 (N_20947,N_16422,N_17555);
or U20948 (N_20948,N_15730,N_17773);
nor U20949 (N_20949,N_15792,N_16316);
and U20950 (N_20950,N_15227,N_15115);
or U20951 (N_20951,N_15159,N_16506);
nor U20952 (N_20952,N_16711,N_16155);
nand U20953 (N_20953,N_17092,N_16678);
xor U20954 (N_20954,N_17024,N_15062);
nand U20955 (N_20955,N_15902,N_15765);
or U20956 (N_20956,N_16626,N_17807);
and U20957 (N_20957,N_15275,N_15484);
and U20958 (N_20958,N_16063,N_16309);
and U20959 (N_20959,N_17717,N_15718);
nand U20960 (N_20960,N_15165,N_16892);
xnor U20961 (N_20961,N_17977,N_15793);
and U20962 (N_20962,N_15870,N_17099);
nand U20963 (N_20963,N_16184,N_17559);
nor U20964 (N_20964,N_17518,N_17989);
and U20965 (N_20965,N_15285,N_16195);
xnor U20966 (N_20966,N_16211,N_15127);
xor U20967 (N_20967,N_17104,N_16451);
nand U20968 (N_20968,N_17884,N_16255);
and U20969 (N_20969,N_16026,N_17577);
nand U20970 (N_20970,N_16635,N_16615);
nand U20971 (N_20971,N_16456,N_16187);
nand U20972 (N_20972,N_16197,N_15502);
and U20973 (N_20973,N_16855,N_16734);
xnor U20974 (N_20974,N_17620,N_17652);
xor U20975 (N_20975,N_15500,N_15920);
and U20976 (N_20976,N_15957,N_15998);
or U20977 (N_20977,N_16990,N_15720);
xor U20978 (N_20978,N_15662,N_17378);
and U20979 (N_20979,N_17596,N_16241);
xor U20980 (N_20980,N_15901,N_16212);
nor U20981 (N_20981,N_16278,N_15624);
and U20982 (N_20982,N_15604,N_15638);
xnor U20983 (N_20983,N_17037,N_17006);
nor U20984 (N_20984,N_17992,N_15906);
xnor U20985 (N_20985,N_16805,N_15695);
and U20986 (N_20986,N_16992,N_16102);
nor U20987 (N_20987,N_17533,N_15692);
xor U20988 (N_20988,N_16160,N_17685);
nor U20989 (N_20989,N_16583,N_15532);
or U20990 (N_20990,N_16678,N_15308);
and U20991 (N_20991,N_17970,N_15063);
xnor U20992 (N_20992,N_17156,N_17376);
and U20993 (N_20993,N_15680,N_15081);
and U20994 (N_20994,N_15144,N_15988);
nand U20995 (N_20995,N_15194,N_15870);
xnor U20996 (N_20996,N_15919,N_17197);
nor U20997 (N_20997,N_16173,N_16953);
nor U20998 (N_20998,N_17182,N_17043);
nand U20999 (N_20999,N_15113,N_16240);
nand U21000 (N_21000,N_18701,N_20650);
nor U21001 (N_21001,N_20099,N_20715);
or U21002 (N_21002,N_20980,N_19260);
and U21003 (N_21003,N_18746,N_19421);
xnor U21004 (N_21004,N_20087,N_20265);
nand U21005 (N_21005,N_19021,N_18188);
nor U21006 (N_21006,N_20954,N_18296);
or U21007 (N_21007,N_20981,N_18343);
and U21008 (N_21008,N_18186,N_20367);
or U21009 (N_21009,N_18462,N_20959);
and U21010 (N_21010,N_19961,N_18211);
and U21011 (N_21011,N_19453,N_19447);
nor U21012 (N_21012,N_18477,N_18481);
or U21013 (N_21013,N_20257,N_18148);
nand U21014 (N_21014,N_18530,N_19080);
nand U21015 (N_21015,N_18947,N_18932);
nor U21016 (N_21016,N_18442,N_20255);
xor U21017 (N_21017,N_18936,N_20978);
nand U21018 (N_21018,N_20784,N_19740);
or U21019 (N_21019,N_20997,N_19083);
nand U21020 (N_21020,N_18690,N_18771);
xor U21021 (N_21021,N_19849,N_18837);
and U21022 (N_21022,N_20609,N_20425);
nand U21023 (N_21023,N_18472,N_20931);
xnor U21024 (N_21024,N_20377,N_19201);
and U21025 (N_21025,N_20412,N_19382);
xor U21026 (N_21026,N_19488,N_20975);
xor U21027 (N_21027,N_19915,N_20334);
nand U21028 (N_21028,N_19725,N_20248);
xnor U21029 (N_21029,N_20688,N_18700);
xor U21030 (N_21030,N_19033,N_20707);
and U21031 (N_21031,N_18583,N_18512);
xor U21032 (N_21032,N_18585,N_20921);
xnor U21033 (N_21033,N_20607,N_18576);
or U21034 (N_21034,N_18480,N_18156);
xor U21035 (N_21035,N_19367,N_20328);
and U21036 (N_21036,N_19786,N_20471);
or U21037 (N_21037,N_20506,N_19994);
or U21038 (N_21038,N_19148,N_20811);
and U21039 (N_21039,N_19888,N_18820);
nor U21040 (N_21040,N_19236,N_19289);
xnor U21041 (N_21041,N_18678,N_19575);
xor U21042 (N_21042,N_18335,N_20705);
nor U21043 (N_21043,N_20354,N_20038);
nand U21044 (N_21044,N_18119,N_18282);
or U21045 (N_21045,N_20005,N_19244);
nor U21046 (N_21046,N_19403,N_20845);
and U21047 (N_21047,N_19733,N_18527);
nand U21048 (N_21048,N_18888,N_20774);
xor U21049 (N_21049,N_18078,N_18214);
and U21050 (N_21050,N_20379,N_18036);
nor U21051 (N_21051,N_20389,N_20962);
xor U21052 (N_21052,N_18274,N_19564);
nand U21053 (N_21053,N_18441,N_20837);
nand U21054 (N_21054,N_19895,N_19062);
xor U21055 (N_21055,N_18682,N_18229);
nand U21056 (N_21056,N_20368,N_20638);
nor U21057 (N_21057,N_20810,N_20970);
or U21058 (N_21058,N_18626,N_20591);
xor U21059 (N_21059,N_20376,N_19066);
nor U21060 (N_21060,N_18525,N_18909);
and U21061 (N_21061,N_19744,N_18065);
and U21062 (N_21062,N_18937,N_19206);
xnor U21063 (N_21063,N_19707,N_20017);
nor U21064 (N_21064,N_20292,N_18999);
or U21065 (N_21065,N_20472,N_20594);
nand U21066 (N_21066,N_18823,N_18278);
nand U21067 (N_21067,N_18336,N_19886);
xnor U21068 (N_21068,N_18658,N_20814);
or U21069 (N_21069,N_18747,N_18692);
or U21070 (N_21070,N_18557,N_19872);
nand U21071 (N_21071,N_19187,N_20671);
and U21072 (N_21072,N_19388,N_18548);
or U21073 (N_21073,N_19762,N_20485);
nand U21074 (N_21074,N_19373,N_18030);
xor U21075 (N_21075,N_18991,N_20022);
nor U21076 (N_21076,N_18327,N_20600);
nand U21077 (N_21077,N_20701,N_18509);
and U21078 (N_21078,N_20072,N_19253);
xnor U21079 (N_21079,N_19930,N_18653);
nor U21080 (N_21080,N_20631,N_19264);
or U21081 (N_21081,N_20436,N_19100);
xor U21082 (N_21082,N_18636,N_18190);
or U21083 (N_21083,N_20424,N_20362);
xnor U21084 (N_21084,N_19933,N_18052);
or U21085 (N_21085,N_19347,N_18633);
xnor U21086 (N_21086,N_20916,N_19739);
nor U21087 (N_21087,N_18147,N_19975);
nor U21088 (N_21088,N_19924,N_19379);
xnor U21089 (N_21089,N_18982,N_20491);
nor U21090 (N_21090,N_20855,N_19095);
and U21091 (N_21091,N_20236,N_19996);
nand U21092 (N_21092,N_20059,N_19225);
nand U21093 (N_21093,N_20805,N_19736);
nand U21094 (N_21094,N_18160,N_19919);
nand U21095 (N_21095,N_20341,N_20274);
nand U21096 (N_21096,N_20599,N_18814);
nor U21097 (N_21097,N_18985,N_18272);
or U21098 (N_21098,N_18169,N_18262);
nor U21099 (N_21099,N_19489,N_20026);
and U21100 (N_21100,N_20403,N_19880);
xor U21101 (N_21101,N_20596,N_18831);
xnor U21102 (N_21102,N_19598,N_18513);
and U21103 (N_21103,N_20699,N_19424);
and U21104 (N_21104,N_18025,N_20523);
and U21105 (N_21105,N_19109,N_20951);
xnor U21106 (N_21106,N_18801,N_20453);
or U21107 (N_21107,N_18136,N_20532);
and U21108 (N_21108,N_18604,N_19115);
nor U21109 (N_21109,N_20957,N_19011);
nor U21110 (N_21110,N_19916,N_19317);
nor U21111 (N_21111,N_20636,N_19013);
xor U21112 (N_21112,N_18780,N_20245);
xnor U21113 (N_21113,N_20181,N_20940);
xnor U21114 (N_21114,N_19061,N_18022);
or U21115 (N_21115,N_18582,N_20787);
nand U21116 (N_21116,N_18574,N_20849);
or U21117 (N_21117,N_20311,N_18080);
xor U21118 (N_21118,N_20298,N_19972);
and U21119 (N_21119,N_19511,N_19679);
and U21120 (N_21120,N_18993,N_19497);
and U21121 (N_21121,N_18688,N_19376);
or U21122 (N_21122,N_20289,N_18458);
nor U21123 (N_21123,N_20081,N_19577);
and U21124 (N_21124,N_20483,N_19071);
or U21125 (N_21125,N_20378,N_20366);
or U21126 (N_21126,N_19102,N_20608);
nand U21127 (N_21127,N_19413,N_18787);
and U21128 (N_21128,N_19398,N_19332);
and U21129 (N_21129,N_18459,N_20223);
nor U21130 (N_21130,N_20675,N_19491);
and U21131 (N_21131,N_19845,N_18643);
nor U21132 (N_21132,N_20309,N_19773);
nor U21133 (N_21133,N_18235,N_20383);
xnor U21134 (N_21134,N_19635,N_18028);
or U21135 (N_21135,N_18641,N_19416);
nor U21136 (N_21136,N_18351,N_19629);
and U21137 (N_21137,N_19111,N_20201);
nand U21138 (N_21138,N_19487,N_19638);
or U21139 (N_21139,N_18420,N_18573);
xor U21140 (N_21140,N_19908,N_18726);
or U21141 (N_21141,N_18245,N_19612);
nor U21142 (N_21142,N_18397,N_19454);
xnor U21143 (N_21143,N_19444,N_19706);
and U21144 (N_21144,N_19223,N_20348);
or U21145 (N_21145,N_20544,N_19392);
nand U21146 (N_21146,N_20509,N_18133);
and U21147 (N_21147,N_20006,N_19330);
nand U21148 (N_21148,N_20204,N_19094);
nand U21149 (N_21149,N_20729,N_20614);
or U21150 (N_21150,N_19999,N_18043);
xnor U21151 (N_21151,N_18804,N_20944);
nand U21152 (N_21152,N_19622,N_18452);
nor U21153 (N_21153,N_20155,N_20351);
and U21154 (N_21154,N_20286,N_19624);
nand U21155 (N_21155,N_20503,N_18146);
nor U21156 (N_21156,N_18998,N_20200);
or U21157 (N_21157,N_19351,N_20540);
and U21158 (N_21158,N_18528,N_18549);
and U21159 (N_21159,N_19568,N_20469);
nand U21160 (N_21160,N_18902,N_20674);
and U21161 (N_21161,N_20941,N_18349);
xnor U21162 (N_21162,N_20337,N_20007);
or U21163 (N_21163,N_20549,N_19466);
xnor U21164 (N_21164,N_18463,N_20199);
or U21165 (N_21165,N_18155,N_18066);
nor U21166 (N_21166,N_18341,N_20844);
nor U21167 (N_21167,N_18308,N_19586);
nor U21168 (N_21168,N_18627,N_19067);
nand U21169 (N_21169,N_18696,N_18830);
or U21170 (N_21170,N_19549,N_20990);
nor U21171 (N_21171,N_19121,N_19037);
xnor U21172 (N_21172,N_19580,N_20687);
or U21173 (N_21173,N_20069,N_18579);
xor U21174 (N_21174,N_19973,N_18038);
or U21175 (N_21175,N_19304,N_18051);
and U21176 (N_21176,N_19477,N_18824);
and U21177 (N_21177,N_18536,N_20495);
nand U21178 (N_21178,N_18491,N_18357);
xnor U21179 (N_21179,N_18802,N_20329);
or U21180 (N_21180,N_19688,N_20507);
and U21181 (N_21181,N_18176,N_18686);
xnor U21182 (N_21182,N_19172,N_20956);
or U21183 (N_21183,N_18957,N_19603);
and U21184 (N_21184,N_19667,N_19559);
nand U21185 (N_21185,N_19181,N_20075);
or U21186 (N_21186,N_18089,N_19976);
nand U21187 (N_21187,N_20039,N_20297);
nor U21188 (N_21188,N_19543,N_18163);
xor U21189 (N_21189,N_20794,N_19276);
xnor U21190 (N_21190,N_18847,N_18851);
and U21191 (N_21191,N_20382,N_20993);
nand U21192 (N_21192,N_20361,N_20347);
nor U21193 (N_21193,N_18942,N_19670);
nor U21194 (N_21194,N_19877,N_20691);
or U21195 (N_21195,N_18563,N_20313);
and U21196 (N_21196,N_20011,N_20876);
xor U21197 (N_21197,N_20719,N_19144);
and U21198 (N_21198,N_18446,N_18012);
nor U21199 (N_21199,N_20102,N_18005);
nor U21200 (N_21200,N_20212,N_18097);
nand U21201 (N_21201,N_18969,N_18488);
nand U21202 (N_21202,N_20879,N_18817);
or U21203 (N_21203,N_20709,N_20229);
or U21204 (N_21204,N_19584,N_18815);
and U21205 (N_21205,N_20175,N_18884);
nor U21206 (N_21206,N_19241,N_18974);
or U21207 (N_21207,N_18222,N_18453);
xnor U21208 (N_21208,N_18911,N_20371);
or U21209 (N_21209,N_18703,N_19325);
nor U21210 (N_21210,N_19215,N_19829);
nor U21211 (N_21211,N_19448,N_20098);
xor U21212 (N_21212,N_20791,N_19799);
or U21213 (N_21213,N_19793,N_19884);
nor U21214 (N_21214,N_18713,N_20909);
or U21215 (N_21215,N_20920,N_19778);
nand U21216 (N_21216,N_18590,N_19246);
and U21217 (N_21217,N_19309,N_20958);
or U21218 (N_21218,N_20898,N_20753);
xor U21219 (N_21219,N_19343,N_18535);
xnor U21220 (N_21220,N_19530,N_19834);
or U21221 (N_21221,N_18611,N_19393);
nor U21222 (N_21222,N_19469,N_18087);
nand U21223 (N_21223,N_18629,N_18032);
nand U21224 (N_21224,N_20977,N_20451);
or U21225 (N_21225,N_18224,N_19270);
and U21226 (N_21226,N_18580,N_20035);
nor U21227 (N_21227,N_19297,N_19257);
xor U21228 (N_21228,N_18927,N_19643);
nand U21229 (N_21229,N_18338,N_20883);
or U21230 (N_21230,N_19256,N_18923);
xor U21231 (N_21231,N_19105,N_20623);
nor U21232 (N_21232,N_20662,N_20530);
nand U21233 (N_21233,N_19230,N_19125);
and U21234 (N_21234,N_18873,N_18533);
xnor U21235 (N_21235,N_19213,N_20748);
and U21236 (N_21236,N_18892,N_20487);
nand U21237 (N_21237,N_18561,N_18587);
or U21238 (N_21238,N_20263,N_20013);
nand U21239 (N_21239,N_19027,N_18526);
xnor U21240 (N_21240,N_18717,N_18450);
nor U21241 (N_21241,N_19366,N_18129);
or U21242 (N_21242,N_20179,N_19914);
xnor U21243 (N_21243,N_19224,N_19988);
nand U21244 (N_21244,N_19651,N_20547);
or U21245 (N_21245,N_20801,N_18153);
and U21246 (N_21246,N_18073,N_19500);
and U21247 (N_21247,N_18182,N_18231);
nand U21248 (N_21248,N_20777,N_20324);
nand U21249 (N_21249,N_19294,N_18455);
nand U21250 (N_21250,N_19848,N_19952);
nand U21251 (N_21251,N_20654,N_20119);
nand U21252 (N_21252,N_19471,N_20987);
and U21253 (N_21253,N_18118,N_20074);
nand U21254 (N_21254,N_20936,N_19610);
and U21255 (N_21255,N_20942,N_20793);
nand U21256 (N_21256,N_20922,N_20796);
nor U21257 (N_21257,N_20349,N_20338);
nand U21258 (N_21258,N_20850,N_20408);
or U21259 (N_21259,N_20237,N_20374);
nor U21260 (N_21260,N_20032,N_19026);
or U21261 (N_21261,N_19771,N_20140);
nand U21262 (N_21262,N_19091,N_19426);
xor U21263 (N_21263,N_18705,N_18426);
nor U21264 (N_21264,N_18264,N_18346);
or U21265 (N_21265,N_18092,N_19616);
nor U21266 (N_21266,N_18061,N_19188);
nor U21267 (N_21267,N_19464,N_19173);
nand U21268 (N_21268,N_20208,N_20147);
and U21269 (N_21269,N_19024,N_20426);
nor U21270 (N_21270,N_18057,N_19182);
and U21271 (N_21271,N_20172,N_19307);
nand U21272 (N_21272,N_19402,N_19274);
and U21273 (N_21273,N_18139,N_18707);
nand U21274 (N_21274,N_19452,N_19969);
or U21275 (N_21275,N_20781,N_18236);
nor U21276 (N_21276,N_18875,N_20832);
or U21277 (N_21277,N_18174,N_20716);
and U21278 (N_21278,N_18638,N_20231);
nor U21279 (N_21279,N_20829,N_19287);
or U21280 (N_21280,N_20492,N_18828);
nor U21281 (N_21281,N_18017,N_19439);
nor U21282 (N_21282,N_18634,N_19846);
nor U21283 (N_21283,N_20431,N_18203);
or U21284 (N_21284,N_20443,N_20067);
nand U21285 (N_21285,N_19015,N_20734);
xnor U21286 (N_21286,N_19319,N_20124);
and U21287 (N_21287,N_20525,N_20937);
nand U21288 (N_21288,N_18261,N_18002);
nor U21289 (N_21289,N_19157,N_18449);
and U21290 (N_21290,N_20380,N_19650);
xnor U21291 (N_21291,N_19088,N_20375);
nand U21292 (N_21292,N_18595,N_20089);
or U21293 (N_21293,N_19904,N_19462);
nor U21294 (N_21294,N_18041,N_20021);
nor U21295 (N_21295,N_18623,N_20531);
nor U21296 (N_21296,N_20856,N_18009);
xnor U21297 (N_21297,N_20510,N_19073);
and U21298 (N_21298,N_20979,N_19672);
xor U21299 (N_21299,N_20282,N_20795);
nand U21300 (N_21300,N_18989,N_19698);
xnor U21301 (N_21301,N_19472,N_20184);
and U21302 (N_21302,N_19782,N_20104);
and U21303 (N_21303,N_19581,N_18408);
xnor U21304 (N_21304,N_18447,N_20740);
nor U21305 (N_21305,N_19434,N_19167);
nor U21306 (N_21306,N_19529,N_18113);
nand U21307 (N_21307,N_18644,N_20479);
xnor U21308 (N_21308,N_18496,N_20893);
nor U21309 (N_21309,N_19159,N_20157);
nor U21310 (N_21310,N_18433,N_19365);
xnor U21311 (N_21311,N_20611,N_19384);
and U21312 (N_21312,N_20296,N_19022);
or U21313 (N_21313,N_20198,N_18853);
nand U21314 (N_21314,N_19784,N_18244);
xor U21315 (N_21315,N_20809,N_18288);
nor U21316 (N_21316,N_18173,N_20452);
or U21317 (N_21317,N_20584,N_19150);
nand U21318 (N_21318,N_18598,N_18166);
and U21319 (N_21319,N_18414,N_18651);
or U21320 (N_21320,N_18482,N_20217);
and U21321 (N_21321,N_19284,N_19763);
nand U21322 (N_21322,N_18001,N_19751);
nand U21323 (N_21323,N_18791,N_18469);
nor U21324 (N_21324,N_19619,N_19712);
xnor U21325 (N_21325,N_19611,N_18945);
nor U21326 (N_21326,N_20877,N_19503);
and U21327 (N_21327,N_19138,N_20533);
nor U21328 (N_21328,N_18374,N_19582);
nor U21329 (N_21329,N_18870,N_20618);
xnor U21330 (N_21330,N_18592,N_18609);
and U21331 (N_21331,N_19548,N_20249);
or U21332 (N_21332,N_20449,N_18323);
nor U21333 (N_21333,N_18287,N_18101);
xnor U21334 (N_21334,N_18781,N_18130);
and U21335 (N_21335,N_18532,N_20346);
nand U21336 (N_21336,N_19820,N_19524);
or U21337 (N_21337,N_19291,N_20148);
nand U21338 (N_21338,N_20456,N_18935);
and U21339 (N_21339,N_18708,N_18096);
nor U21340 (N_21340,N_19790,N_18265);
and U21341 (N_21341,N_18310,N_20244);
and U21342 (N_21342,N_18733,N_18213);
xor U21343 (N_21343,N_20446,N_20496);
and U21344 (N_21344,N_19345,N_18861);
nand U21345 (N_21345,N_19627,N_18751);
and U21346 (N_21346,N_18271,N_20385);
or U21347 (N_21347,N_20935,N_20321);
nor U21348 (N_21348,N_18732,N_19713);
and U21349 (N_21349,N_20156,N_19777);
nand U21350 (N_21350,N_18309,N_20842);
and U21351 (N_21351,N_20352,N_19551);
xnor U21352 (N_21352,N_19867,N_20222);
or U21353 (N_21353,N_20894,N_18880);
and U21354 (N_21354,N_18887,N_18578);
or U21355 (N_21355,N_20275,N_19387);
xor U21356 (N_21356,N_20142,N_19669);
and U21357 (N_21357,N_18984,N_18545);
xor U21358 (N_21358,N_19016,N_20955);
xnor U21359 (N_21359,N_19571,N_18042);
or U21360 (N_21360,N_19708,N_18559);
nor U21361 (N_21361,N_19843,N_18725);
nor U21362 (N_21362,N_18445,N_20463);
or U21363 (N_21363,N_19866,N_18050);
and U21364 (N_21364,N_18220,N_20888);
and U21365 (N_21365,N_18276,N_19760);
nand U21366 (N_21366,N_19288,N_18739);
or U21367 (N_21367,N_18874,N_18767);
nand U21368 (N_21368,N_18508,N_20640);
and U21369 (N_21369,N_18786,N_20397);
nor U21370 (N_21370,N_20224,N_19131);
xor U21371 (N_21371,N_19463,N_18370);
xnor U21372 (N_21372,N_18172,N_18813);
or U21373 (N_21373,N_18293,N_19864);
or U21374 (N_21374,N_20350,N_19517);
nor U21375 (N_21375,N_20852,N_20384);
and U21376 (N_21376,N_19767,N_19953);
nand U21377 (N_21377,N_18840,N_18869);
nand U21378 (N_21378,N_18109,N_20713);
and U21379 (N_21379,N_18313,N_19252);
xor U21380 (N_21380,N_20939,N_18177);
nand U21381 (N_21381,N_19401,N_18511);
nand U21382 (N_21382,N_18689,N_18342);
nor U21383 (N_21383,N_19749,N_19496);
nor U21384 (N_21384,N_18056,N_20667);
or U21385 (N_21385,N_18444,N_19711);
and U21386 (N_21386,N_19639,N_18350);
nand U21387 (N_21387,N_18962,N_19110);
nor U21388 (N_21388,N_20043,N_19427);
nand U21389 (N_21389,N_19684,N_18208);
and U21390 (N_21390,N_18094,N_19630);
and U21391 (N_21391,N_18972,N_20372);
nand U21392 (N_21392,N_19197,N_18081);
xnor U21393 (N_21393,N_19789,N_20735);
or U21394 (N_21394,N_20731,N_18591);
or U21395 (N_21395,N_20808,N_19179);
nor U21396 (N_21396,N_19852,N_18669);
or U21397 (N_21397,N_20127,N_20702);
nand U21398 (N_21398,N_20566,N_18683);
or U21399 (N_21399,N_19889,N_19894);
or U21400 (N_21400,N_19657,N_19579);
and U21401 (N_21401,N_18337,N_20615);
or U21402 (N_21402,N_20154,N_18108);
or U21403 (N_21403,N_19572,N_18033);
or U21404 (N_21404,N_18018,N_18646);
and U21405 (N_21405,N_19455,N_19300);
xnor U21406 (N_21406,N_19007,N_20111);
or U21407 (N_21407,N_18670,N_19836);
xnor U21408 (N_21408,N_20863,N_18484);
nand U21409 (N_21409,N_19126,N_20214);
xor U21410 (N_21410,N_19879,N_18956);
or U21411 (N_21411,N_19911,N_19534);
xnor U21412 (N_21412,N_18008,N_19608);
and U21413 (N_21413,N_19565,N_19090);
and U21414 (N_21414,N_18523,N_20191);
nand U21415 (N_21415,N_20875,N_18493);
and U21416 (N_21416,N_19556,N_19231);
and U21417 (N_21417,N_19419,N_18389);
or U21418 (N_21418,N_19028,N_20370);
nand U21419 (N_21419,N_18534,N_20441);
or U21420 (N_21420,N_19944,N_18090);
and U21421 (N_21421,N_19951,N_19470);
or U21422 (N_21422,N_20874,N_18316);
xor U21423 (N_21423,N_18663,N_18552);
xor U21424 (N_21424,N_18454,N_19178);
or U21425 (N_21425,N_20092,N_19128);
or U21426 (N_21426,N_18483,N_19386);
nand U21427 (N_21427,N_19003,N_20151);
nand U21428 (N_21428,N_18436,N_18344);
or U21429 (N_21429,N_19788,N_19456);
and U21430 (N_21430,N_18404,N_19898);
and U21431 (N_21431,N_18200,N_18601);
nand U21432 (N_21432,N_20919,N_18886);
nand U21433 (N_21433,N_19589,N_19342);
or U21434 (N_21434,N_20840,N_20992);
nand U21435 (N_21435,N_20024,N_19585);
and U21436 (N_21436,N_19907,N_20839);
or U21437 (N_21437,N_19747,N_20235);
or U21438 (N_21438,N_18011,N_18320);
and U21439 (N_21439,N_19748,N_18248);
nand U21440 (N_21440,N_19897,N_18777);
or U21441 (N_21441,N_18883,N_20268);
xnor U21442 (N_21442,N_18857,N_18062);
nand U21443 (N_21443,N_20381,N_20995);
nor U21444 (N_21444,N_19647,N_18330);
nor U21445 (N_21445,N_18893,N_19974);
xnor U21446 (N_21446,N_20910,N_20115);
or U21447 (N_21447,N_19312,N_19314);
xor U21448 (N_21448,N_20945,N_20878);
or U21449 (N_21449,N_19561,N_19839);
nand U21450 (N_21450,N_19085,N_18460);
xnor U21451 (N_21451,N_18219,N_20188);
nand U21452 (N_21452,N_18571,N_18765);
and U21453 (N_21453,N_18635,N_18014);
or U21454 (N_21454,N_20467,N_19910);
nor U21455 (N_21455,N_19406,N_18471);
nor U21456 (N_21456,N_19368,N_18671);
nor U21457 (N_21457,N_18753,N_19353);
nand U21458 (N_21458,N_20029,N_19631);
nor U21459 (N_21459,N_18518,N_20225);
nand U21460 (N_21460,N_18685,N_20972);
xor U21461 (N_21461,N_19927,N_20514);
or U21462 (N_21462,N_19958,N_19675);
and U21463 (N_21463,N_18209,N_18976);
xnor U21464 (N_21464,N_19163,N_20080);
and U21465 (N_21465,N_20143,N_19282);
and U21466 (N_21466,N_20927,N_19086);
nand U21467 (N_21467,N_18154,N_19117);
nand U21468 (N_21468,N_20393,N_18864);
and U21469 (N_21469,N_19268,N_19438);
nand U21470 (N_21470,N_18400,N_18560);
and U21471 (N_21471,N_20813,N_20798);
xnor U21472 (N_21472,N_18656,N_20565);
or U21473 (N_21473,N_18237,N_20195);
and U21474 (N_21474,N_19687,N_19449);
or U21475 (N_21475,N_19104,N_20247);
and U21476 (N_21476,N_20867,N_18630);
or U21477 (N_21477,N_18364,N_20516);
or U21478 (N_21478,N_20266,N_19702);
xor U21479 (N_21479,N_18915,N_19059);
and U21480 (N_21480,N_19508,N_18827);
nor U21481 (N_21481,N_19533,N_18825);
nor U21482 (N_21482,N_18137,N_20925);
nor U21483 (N_21483,N_20527,N_18267);
or U21484 (N_21484,N_20129,N_20714);
xor U21485 (N_21485,N_20588,N_20415);
and U21486 (N_21486,N_18632,N_19132);
or U21487 (N_21487,N_19233,N_18805);
nor U21488 (N_21488,N_19058,N_19507);
and U21489 (N_21489,N_20333,N_20851);
or U21490 (N_21490,N_20345,N_20901);
nand U21491 (N_21491,N_20278,N_20088);
nor U21492 (N_21492,N_19074,N_19254);
nor U21493 (N_21493,N_19315,N_20256);
nor U21494 (N_21494,N_20316,N_19337);
or U21495 (N_21495,N_19475,N_18046);
nand U21496 (N_21496,N_18240,N_18562);
xnor U21497 (N_21497,N_20799,N_19106);
nand U21498 (N_21498,N_19468,N_18866);
and U21499 (N_21499,N_20578,N_19542);
nor U21500 (N_21500,N_19302,N_19029);
and U21501 (N_21501,N_20163,N_19005);
and U21502 (N_21502,N_20420,N_18834);
or U21503 (N_21503,N_19296,N_19193);
xor U21504 (N_21504,N_19823,N_19779);
or U21505 (N_21505,N_19764,N_18619);
nand U21506 (N_21506,N_18207,N_18440);
nand U21507 (N_21507,N_20853,N_20363);
or U21508 (N_21508,N_19754,N_18158);
and U21509 (N_21509,N_18067,N_18439);
xor U21510 (N_21510,N_19522,N_20947);
nor U21511 (N_21511,N_20930,N_19756);
xor U21512 (N_21512,N_19576,N_19092);
nand U21513 (N_21513,N_19941,N_18958);
nand U21514 (N_21514,N_20086,N_20335);
xnor U21515 (N_21515,N_20180,N_20399);
and U21516 (N_21516,N_20949,N_18256);
xor U21517 (N_21517,N_18218,N_20008);
nor U21518 (N_21518,N_20246,N_20196);
and U21519 (N_21519,N_18970,N_18498);
nand U21520 (N_21520,N_20183,N_19937);
nor U21521 (N_21521,N_19593,N_18138);
or U21522 (N_21522,N_19262,N_20529);
nor U21523 (N_21523,N_18419,N_20106);
or U21524 (N_21524,N_18808,N_18183);
nor U21525 (N_21525,N_20892,N_20693);
or U21526 (N_21526,N_19514,N_19804);
xnor U21527 (N_21527,N_20756,N_20053);
nor U21528 (N_21528,N_19617,N_19597);
or U21529 (N_21529,N_20182,N_20511);
or U21530 (N_21530,N_20331,N_20816);
and U21531 (N_21531,N_19437,N_19642);
nand U21532 (N_21532,N_18111,N_20698);
or U21533 (N_21533,N_18740,N_19202);
and U21534 (N_21534,N_19541,N_20645);
and U21535 (N_21535,N_18555,N_19506);
or U21536 (N_21536,N_18238,N_19012);
nand U21537 (N_21537,N_20652,N_18451);
or U21538 (N_21538,N_18735,N_18944);
and U21539 (N_21539,N_19535,N_20557);
nand U21540 (N_21540,N_19259,N_20218);
nor U21541 (N_21541,N_19335,N_19634);
or U21542 (N_21542,N_19936,N_20232);
nand U21543 (N_21543,N_18675,N_19636);
and U21544 (N_21544,N_18943,N_19162);
nand U21545 (N_21545,N_19285,N_20918);
nand U21546 (N_21546,N_20771,N_18639);
nand U21547 (N_21547,N_18565,N_18551);
or U21548 (N_21548,N_19440,N_18766);
nor U21549 (N_21549,N_20827,N_20595);
nor U21550 (N_21550,N_19155,N_20033);
and U21551 (N_21551,N_18225,N_18312);
nand U21552 (N_21552,N_19982,N_18843);
xor U21553 (N_21553,N_19991,N_20685);
nor U21554 (N_21554,N_19806,N_19665);
nor U21555 (N_21555,N_18004,N_19774);
nand U21556 (N_21556,N_18736,N_19054);
xnor U21557 (N_21557,N_20964,N_18305);
and U21558 (N_21558,N_19478,N_19097);
or U21559 (N_21559,N_19526,N_18194);
and U21560 (N_21560,N_20788,N_18912);
xor U21561 (N_21561,N_18247,N_18546);
or U21562 (N_21562,N_19135,N_19513);
nor U21563 (N_21563,N_19093,N_19045);
nor U21564 (N_21564,N_19794,N_18384);
nand U21565 (N_21565,N_19422,N_18858);
xnor U21566 (N_21566,N_18354,N_20066);
nor U21567 (N_21567,N_18233,N_19661);
or U21568 (N_21568,N_19905,N_18134);
xor U21569 (N_21569,N_18243,N_20190);
xor U21570 (N_21570,N_18919,N_18811);
nand U21571 (N_21571,N_20745,N_20897);
or U21572 (N_21572,N_20342,N_18833);
nand U21573 (N_21573,N_19383,N_20136);
or U21574 (N_21574,N_20911,N_20160);
nand U21575 (N_21575,N_19978,N_19130);
nor U21576 (N_21576,N_20090,N_20974);
and U21577 (N_21577,N_18045,N_19137);
nand U21578 (N_21578,N_20736,N_19145);
nand U21579 (N_21579,N_20470,N_18665);
nor U21580 (N_21580,N_18783,N_19710);
nor U21581 (N_21581,N_19940,N_19495);
and U21582 (N_21582,N_19175,N_18189);
and U21583 (N_21583,N_18179,N_19676);
nor U21584 (N_21584,N_20421,N_20783);
and U21585 (N_21585,N_20015,N_20488);
and U21586 (N_21586,N_18121,N_19412);
nand U21587 (N_21587,N_19531,N_18939);
xor U21588 (N_21588,N_20679,N_18849);
nor U21589 (N_21589,N_18161,N_18401);
nand U21590 (N_21590,N_19239,N_18728);
nand U21591 (N_21591,N_18047,N_18818);
nor U21592 (N_21592,N_19854,N_18467);
or U21593 (N_21593,N_20681,N_18901);
xnor U21594 (N_21594,N_18468,N_19573);
and U21595 (N_21595,N_18301,N_20520);
xor U21596 (N_21596,N_18704,N_19108);
and U21597 (N_21597,N_19047,N_20128);
nor U21598 (N_21598,N_20482,N_19222);
and U21599 (N_21599,N_18764,N_18844);
or U21600 (N_21600,N_19605,N_20648);
nor U21601 (N_21601,N_20985,N_20272);
xnor U21602 (N_21602,N_18519,N_19211);
or U21603 (N_21603,N_20454,N_19525);
or U21604 (N_21604,N_18149,N_20830);
nand U21605 (N_21605,N_20435,N_20187);
or U21606 (N_21606,N_20302,N_18910);
or U21607 (N_21607,N_18319,N_20766);
nand U21608 (N_21608,N_18687,N_19435);
and U21609 (N_21609,N_18140,N_19360);
nor U21610 (N_21610,N_19680,N_19546);
xnor U21611 (N_21611,N_20114,N_19646);
nor U21612 (N_21612,N_20613,N_18292);
nand U21613 (N_21613,N_18882,N_18461);
nor U21614 (N_21614,N_19391,N_18596);
or U21615 (N_21615,N_18540,N_20281);
and U21616 (N_21616,N_18524,N_19780);
or U21617 (N_21617,N_18588,N_19008);
and U21618 (N_21618,N_18879,N_18151);
nand U21619 (N_21619,N_18421,N_19258);
or U21620 (N_21620,N_20121,N_20933);
xor U21621 (N_21621,N_18345,N_19423);
and U21622 (N_21622,N_18645,N_20433);
nor U21623 (N_21623,N_20310,N_18900);
nand U21624 (N_21624,N_19357,N_19051);
nor U21625 (N_21625,N_19519,N_20998);
or U21626 (N_21626,N_20401,N_20680);
xnor U21627 (N_21627,N_20301,N_20678);
xor U21628 (N_21628,N_18607,N_19243);
nor U21629 (N_21629,N_19286,N_18785);
and U21630 (N_21630,N_18929,N_20097);
nand U21631 (N_21631,N_18662,N_18885);
or U21632 (N_21632,N_19425,N_19114);
or U21633 (N_21633,N_19658,N_19662);
and U21634 (N_21634,N_19014,N_19429);
nand U21635 (N_21635,N_19563,N_20085);
nor U21636 (N_21636,N_20489,N_19826);
and U21637 (N_21637,N_19633,N_18898);
and U21638 (N_21638,N_19832,N_20094);
nand U21639 (N_21639,N_18795,N_18495);
nor U21640 (N_21640,N_20480,N_18198);
nand U21641 (N_21641,N_18616,N_19160);
xnor U21642 (N_21642,N_18822,N_18378);
and U21643 (N_21643,N_18920,N_20513);
or U21644 (N_21644,N_19023,N_18904);
nand U21645 (N_21645,N_19295,N_19204);
nor U21646 (N_21646,N_20084,N_18379);
nand U21647 (N_21647,N_19686,N_19890);
nand U21648 (N_21648,N_20580,N_20541);
nand U21649 (N_21649,N_18916,N_19544);
nor U21650 (N_21650,N_20019,N_18409);
nand U21651 (N_21651,N_19874,N_19119);
xnor U21652 (N_21652,N_19983,N_20885);
xor U21653 (N_21653,N_20881,N_20490);
nand U21654 (N_21654,N_19746,N_20010);
nand U21655 (N_21655,N_19833,N_18144);
xnor U21656 (N_21656,N_19903,N_20473);
xor U21657 (N_21657,N_18114,N_18907);
nor U21658 (N_21658,N_18842,N_18721);
xnor U21659 (N_21659,N_19745,N_20288);
nand U21660 (N_21660,N_18277,N_20498);
xnor U21661 (N_21661,N_19123,N_19775);
and U21662 (N_21662,N_18412,N_20259);
nand U21663 (N_21663,N_18128,N_18784);
nand U21664 (N_21664,N_19813,N_20724);
nand U21665 (N_21665,N_20826,N_20770);
xor U21666 (N_21666,N_18284,N_20044);
and U21667 (N_21667,N_18505,N_19737);
nor U21668 (N_21668,N_19934,N_19420);
xnor U21669 (N_21669,N_19355,N_19742);
xnor U21670 (N_21670,N_20576,N_19267);
and U21671 (N_21671,N_19065,N_19394);
and U21672 (N_21672,N_18698,N_19498);
xor U21673 (N_21673,N_18326,N_18127);
xor U21674 (N_21674,N_19313,N_20060);
nand U21675 (N_21675,N_19263,N_19168);
nand U21676 (N_21676,N_18143,N_20821);
nand U21677 (N_21677,N_19063,N_18387);
and U21678 (N_21678,N_20590,N_19140);
nand U21679 (N_21679,N_20620,N_20760);
nand U21680 (N_21680,N_20508,N_18395);
or U21681 (N_21681,N_19928,N_18069);
nand U21682 (N_21682,N_19685,N_18654);
or U21683 (N_21683,N_19965,N_20439);
nor U21684 (N_21684,N_20889,N_18978);
xor U21685 (N_21685,N_20858,N_18352);
nor U21686 (N_21686,N_18329,N_18720);
or U21687 (N_21687,N_20928,N_18259);
and U21688 (N_21688,N_19174,N_19995);
nor U21689 (N_21689,N_19395,N_20670);
or U21690 (N_21690,N_20167,N_19810);
nand U21691 (N_21691,N_18353,N_18075);
or U21692 (N_21692,N_18709,N_20475);
nand U21693 (N_21693,N_18088,N_20134);
nand U21694 (N_21694,N_19555,N_19043);
nor U21695 (N_21695,N_19860,N_19010);
nand U21696 (N_21696,N_19626,N_20061);
nand U21697 (N_21697,N_19129,N_19553);
nand U21698 (N_21698,N_18193,N_19855);
and U21699 (N_21699,N_20538,N_19652);
xnor U21700 (N_21700,N_20130,N_20323);
and U21701 (N_21701,N_20697,N_18744);
or U21702 (N_21702,N_18380,N_18602);
nor U21703 (N_21703,N_20836,N_18933);
and U21704 (N_21704,N_20146,N_20150);
xnor U21705 (N_21705,N_19732,N_19798);
nor U21706 (N_21706,N_20812,N_19671);
nand U21707 (N_21707,N_19981,N_18980);
nor U21708 (N_21708,N_18572,N_18760);
nor U21709 (N_21709,N_20912,N_18191);
or U21710 (N_21710,N_18295,N_18807);
xnor U21711 (N_21711,N_19663,N_19459);
xor U21712 (N_21712,N_20336,N_20737);
xor U21713 (N_21713,N_18470,N_19308);
or U21714 (N_21714,N_19031,N_20800);
nand U21715 (N_21715,N_20854,N_20656);
nand U21716 (N_21716,N_20581,N_18365);
nor U21717 (N_21717,N_20637,N_20665);
nand U21718 (N_21718,N_18167,N_19220);
xnor U21719 (N_21719,N_20141,N_19283);
or U21720 (N_21720,N_18321,N_18895);
xnor U21721 (N_21721,N_19446,N_18543);
nand U21722 (N_21722,N_18841,N_18928);
xnor U21723 (N_21723,N_19795,N_18093);
and U21724 (N_21724,N_19056,N_20644);
nand U21725 (N_21725,N_20332,N_20828);
xnor U21726 (N_21726,N_19637,N_18748);
xor U21727 (N_21727,N_19004,N_19141);
and U21728 (N_21728,N_18681,N_18606);
or U21729 (N_21729,N_20669,N_19346);
nor U21730 (N_21730,N_19666,N_20261);
and U21731 (N_21731,N_19184,N_18135);
nor U21732 (N_21732,N_18250,N_18377);
xnor U21733 (N_21733,N_18599,N_18230);
xnor U21734 (N_21734,N_19363,N_20107);
nand U21735 (N_21735,N_19876,N_20045);
or U21736 (N_21736,N_18044,N_19409);
xor U21737 (N_21737,N_19787,N_19070);
or U21738 (N_21738,N_18099,N_18021);
nand U21739 (N_21739,N_18727,N_18881);
nand U21740 (N_21740,N_20561,N_19574);
nor U21741 (N_21741,N_19523,N_18624);
nand U21742 (N_21742,N_20994,N_19923);
nor U21743 (N_21743,N_18878,N_19505);
nor U21744 (N_21744,N_18965,N_20712);
xnor U21745 (N_21745,N_19596,N_18106);
nand U21746 (N_21746,N_18184,N_20461);
xor U21747 (N_21747,N_19232,N_18862);
and U21748 (N_21748,N_19840,N_18438);
xor U21749 (N_21749,N_19192,N_18968);
and U21750 (N_21750,N_19293,N_20240);
and U21751 (N_21751,N_18854,N_18564);
and U21752 (N_21752,N_20861,N_18202);
xor U21753 (N_21753,N_18649,N_18504);
or U21754 (N_21754,N_19053,N_18415);
nand U21755 (N_21755,N_19838,N_20859);
xor U21756 (N_21756,N_19414,N_18375);
or U21757 (N_21757,N_18115,N_19199);
nand U21758 (N_21758,N_20857,N_19089);
nor U21759 (N_21759,N_19191,N_19251);
xor U21760 (N_21760,N_18263,N_18275);
xnor U21761 (N_21761,N_19177,N_20700);
nor U21762 (N_21762,N_18997,N_19583);
xnor U21763 (N_21763,N_19699,N_18059);
xnor U21764 (N_21764,N_20234,N_19545);
nand U21765 (N_21765,N_19156,N_20899);
nand U21766 (N_21766,N_19537,N_20907);
and U21767 (N_21767,N_18537,N_19521);
or U21768 (N_21768,N_18790,N_19501);
xor U21769 (N_21769,N_20264,N_20579);
nor U21770 (N_21770,N_20989,N_20986);
nand U21771 (N_21771,N_20391,N_20720);
and U21772 (N_21772,N_20915,N_18076);
nor U21773 (N_21773,N_20792,N_18960);
and U21774 (N_21774,N_18637,N_18672);
nor U21775 (N_21775,N_18196,N_19692);
xor U21776 (N_21776,N_19417,N_18423);
xor U21777 (N_21777,N_19796,N_19587);
xnor U21778 (N_21778,N_20673,N_19757);
nor U21779 (N_21779,N_19209,N_20023);
or U21780 (N_21780,N_19098,N_19602);
and U21781 (N_21781,N_20546,N_18399);
or U21782 (N_21782,N_20474,N_20305);
or U21783 (N_21783,N_20704,N_18605);
and U21784 (N_21784,N_20083,N_20759);
and U21785 (N_21785,N_19766,N_20241);
nand U21786 (N_21786,N_20071,N_20062);
nor U21787 (N_21787,N_19479,N_18625);
and U21788 (N_21788,N_18810,N_20502);
or U21789 (N_21789,N_18570,N_19887);
xor U21790 (N_21790,N_19539,N_18903);
or U21791 (N_21791,N_19176,N_20582);
xor U21792 (N_21792,N_18494,N_20824);
and U21793 (N_21793,N_18489,N_19279);
and U21794 (N_21794,N_18948,N_18967);
xnor U21795 (N_21795,N_18210,N_18131);
xor U21796 (N_21796,N_19431,N_20717);
nor U21797 (N_21797,N_20118,N_18072);
or U21798 (N_21798,N_18058,N_20924);
nand U21799 (N_21799,N_20790,N_18953);
or U21800 (N_21800,N_19590,N_20260);
and U21801 (N_21801,N_20220,N_20575);
nand U21802 (N_21802,N_19722,N_19042);
and U21803 (N_21803,N_18417,N_20135);
xnor U21804 (N_21804,N_19492,N_19985);
xor U21805 (N_21805,N_19957,N_19993);
xnor U21806 (N_21806,N_19229,N_20616);
nand U21807 (N_21807,N_20552,N_19772);
nor U21808 (N_21808,N_20782,N_20056);
and U21809 (N_21809,N_18091,N_19189);
nand U21810 (N_21810,N_19428,N_20563);
nand U21811 (N_21811,N_19389,N_20786);
nand U21812 (N_21812,N_20754,N_20173);
xor U21813 (N_21813,N_18026,N_20870);
xor U21814 (N_21814,N_18930,N_19683);
or U21815 (N_21815,N_20279,N_18877);
xor U21816 (N_21816,N_18302,N_19929);
xnor U21817 (N_21817,N_20238,N_18859);
and U21818 (N_21818,N_19120,N_20983);
and U21819 (N_21819,N_18197,N_20322);
xnor U21820 (N_21820,N_20768,N_20197);
or U21821 (N_21821,N_18914,N_19025);
xnor U21822 (N_21822,N_18431,N_19250);
nand U21823 (N_21823,N_20486,N_19805);
xnor U21824 (N_21824,N_18283,N_18141);
nor U21825 (N_21825,N_18204,N_19613);
nand U21826 (N_21826,N_19557,N_18215);
and U21827 (N_21827,N_20168,N_20230);
nand U21828 (N_21828,N_18315,N_20070);
nor U21829 (N_21829,N_18661,N_20055);
and U21830 (N_21830,N_20049,N_19305);
nand U21831 (N_21831,N_19984,N_20545);
nand U21832 (N_21832,N_19913,N_18950);
or U21833 (N_21833,N_20835,N_19743);
and U21834 (N_21834,N_18279,N_19112);
or U21835 (N_21835,N_20948,N_19032);
and U21836 (N_21836,N_20779,N_19358);
nand U21837 (N_21837,N_20553,N_19482);
and U21838 (N_21838,N_19474,N_19938);
nand U21839 (N_21839,N_19298,N_20526);
or U21840 (N_21840,N_18897,N_18613);
and U21841 (N_21841,N_19380,N_20633);
or U21842 (N_21842,N_18782,N_18547);
xor U21843 (N_21843,N_18702,N_20619);
nand U21844 (N_21844,N_19249,N_18386);
xnor U21845 (N_21845,N_20568,N_20250);
nand U21846 (N_21846,N_20030,N_20866);
and U21847 (N_21847,N_20524,N_20054);
xnor U21848 (N_21848,N_19050,N_18797);
xor U21849 (N_21849,N_19001,N_20110);
or U21850 (N_21850,N_20239,N_20419);
nor U21851 (N_21851,N_18934,N_19364);
xor U21852 (N_21852,N_19018,N_20537);
xor U21853 (N_21853,N_19136,N_20763);
or U21854 (N_21854,N_19458,N_20430);
nor U21855 (N_21855,N_19761,N_20554);
xor U21856 (N_21856,N_19660,N_18836);
nand U21857 (N_21857,N_19306,N_19681);
nand U21858 (N_21858,N_18855,N_18355);
nor U21859 (N_21859,N_19900,N_19436);
xnor U21860 (N_21860,N_20395,N_18185);
xor U21861 (N_21861,N_19127,N_20999);
or U21862 (N_21862,N_20388,N_20226);
or U21863 (N_21863,N_18667,N_18693);
and U21864 (N_21864,N_18752,N_19377);
nor U21865 (N_21865,N_18098,N_19678);
xnor U21866 (N_21866,N_19165,N_20117);
or U21867 (N_21867,N_19547,N_20612);
nor U21868 (N_21868,N_18922,N_18360);
nand U21869 (N_21869,N_19715,N_19516);
nand U21870 (N_21870,N_20460,N_19705);
and U21871 (N_21871,N_20818,N_19800);
and U21872 (N_21872,N_19361,N_19831);
and U21873 (N_21873,N_18071,N_19277);
nor U21874 (N_21874,N_20914,N_19035);
nor U21875 (N_21875,N_18759,N_18199);
or U21876 (N_21876,N_18290,N_20418);
or U21877 (N_21877,N_19532,N_18383);
xor U21878 (N_21878,N_18159,N_18657);
or U21879 (N_21879,N_18221,N_20589);
and U21880 (N_21880,N_18049,N_20276);
and U21881 (N_21881,N_19195,N_18103);
or U21882 (N_21882,N_19340,N_20186);
xnor U21883 (N_21883,N_19857,N_20884);
and U21884 (N_21884,N_18990,N_20373);
and U21885 (N_21885,N_20887,N_19133);
nor U21886 (N_21886,N_20762,N_20315);
or U21887 (N_21887,N_19101,N_20886);
and U21888 (N_21888,N_18234,N_19408);
nor U21889 (N_21889,N_18756,N_19081);
nor U21890 (N_21890,N_18567,N_19139);
nor U21891 (N_21891,N_20749,N_20138);
nor U21892 (N_21892,N_19871,N_18577);
xnor U21893 (N_21893,N_20484,N_19170);
nand U21894 (N_21894,N_18515,N_20598);
nand U21895 (N_21895,N_20539,N_18120);
xor U21896 (N_21896,N_20494,N_20233);
nand U21897 (N_21897,N_19560,N_18116);
xnor U21898 (N_21898,N_18334,N_19323);
xor U21899 (N_21899,N_20176,N_20052);
xnor U21900 (N_21900,N_18706,N_20517);
nand U21901 (N_21901,N_18206,N_19902);
or U21902 (N_21902,N_19460,N_18223);
and U21903 (N_21903,N_18422,N_19483);
nor U21904 (N_21904,N_20676,N_20284);
or U21905 (N_21905,N_19801,N_20457);
nand U21906 (N_21906,N_20755,N_18178);
nor U21907 (N_21907,N_18612,N_20819);
nor U21908 (N_21908,N_20192,N_20882);
or U21909 (N_21909,N_18876,N_18371);
nor U21910 (N_21910,N_20703,N_19000);
or U21911 (N_21911,N_20610,N_20091);
or U21912 (N_21912,N_19240,N_20535);
xor U21913 (N_21913,N_19341,N_20360);
and U21914 (N_21914,N_20603,N_19099);
and U21915 (N_21915,N_20550,N_20077);
nand U21916 (N_21916,N_20057,N_18655);
xnor U21917 (N_21917,N_18659,N_19947);
xor U21918 (N_21918,N_20846,N_19569);
nand U21919 (N_21919,N_18027,N_20295);
and U21920 (N_21920,N_20048,N_20743);
nor U21921 (N_21921,N_18542,N_19356);
xor U21922 (N_21922,N_20410,N_18994);
and U21923 (N_21923,N_19219,N_20621);
nor U21924 (N_21924,N_19235,N_19194);
nor U21925 (N_21925,N_19896,N_20661);
nor U21926 (N_21926,N_18816,N_20658);
xnor U21927 (N_21927,N_20725,N_19628);
nand U21928 (N_21928,N_19512,N_18428);
nor U21929 (N_21929,N_20666,N_18520);
nand U21930 (N_21930,N_18896,N_19538);
and U21931 (N_21931,N_19079,N_20923);
and U21932 (N_21932,N_20560,N_20569);
or U21933 (N_21933,N_18964,N_20442);
xnor U21934 (N_21934,N_20971,N_18095);
and U21935 (N_21935,N_20726,N_19275);
or U21936 (N_21936,N_19690,N_19765);
xnor U21937 (N_21937,N_20004,N_19709);
and U21938 (N_21938,N_19695,N_20402);
xor U21939 (N_21939,N_18110,N_20105);
or U21940 (N_21940,N_19087,N_20583);
or U21941 (N_21941,N_20162,N_19693);
or U21942 (N_21942,N_20982,N_19724);
and U21943 (N_21943,N_19212,N_19374);
xor U21944 (N_21944,N_20317,N_19149);
or U21945 (N_21945,N_20327,N_18289);
nor U21946 (N_21946,N_18754,N_19266);
nor U21947 (N_21947,N_18340,N_18000);
nor U21948 (N_21948,N_18792,N_18499);
or U21949 (N_21949,N_18722,N_20215);
nand U21950 (N_21950,N_20570,N_20177);
or U21951 (N_21951,N_20628,N_18743);
nand U21952 (N_21952,N_18443,N_19339);
or U21953 (N_21953,N_18788,N_19835);
nand U21954 (N_21954,N_20521,N_19166);
or U21955 (N_21955,N_19570,N_20394);
nor U21956 (N_21956,N_19301,N_18405);
and U21957 (N_21957,N_19604,N_20051);
nand U21958 (N_21958,N_18324,N_18029);
xnor U21959 (N_21959,N_19623,N_20789);
nand U21960 (N_21960,N_19404,N_20558);
nand U21961 (N_21961,N_18048,N_18304);
xor U21962 (N_21962,N_18325,N_19971);
nand U21963 (N_21963,N_18846,N_20710);
xor U21964 (N_21964,N_19390,N_20174);
nor U21965 (N_21965,N_18737,N_19461);
nand U21966 (N_21966,N_19960,N_18677);
and U21967 (N_21967,N_19731,N_18541);
and U21968 (N_21968,N_19935,N_19451);
or U21969 (N_21969,N_20020,N_20820);
nand U21970 (N_21970,N_18773,N_19959);
and U21971 (N_21971,N_19039,N_19484);
xnor U21972 (N_21972,N_20751,N_19901);
and U21973 (N_21973,N_18850,N_18684);
nor U21974 (N_21974,N_18906,N_19333);
and U21975 (N_21975,N_18954,N_18382);
nor U21976 (N_21976,N_18486,N_18971);
xor U21977 (N_21977,N_18652,N_18232);
nor U21978 (N_21978,N_18988,N_19807);
nor U21979 (N_21979,N_20325,N_20690);
nand U21980 (N_21980,N_18077,N_18674);
xnor U21981 (N_21981,N_18517,N_19348);
or U21982 (N_21982,N_20775,N_19645);
xnor U21983 (N_21983,N_19407,N_19618);
nor U21984 (N_21984,N_20455,N_19714);
nor U21985 (N_21985,N_18150,N_20953);
and U21986 (N_21986,N_20834,N_18286);
nor U21987 (N_21987,N_18889,N_19510);
nor U21988 (N_21988,N_20358,N_20205);
or U21989 (N_21989,N_18531,N_19237);
nor U21990 (N_21990,N_18676,N_19118);
and U21991 (N_21991,N_18863,N_20677);
xor U21992 (N_21992,N_18122,N_20585);
or U21993 (N_21993,N_20862,N_20314);
or U21994 (N_21994,N_19980,N_20254);
xnor U21995 (N_21995,N_18941,N_19811);
and U21996 (N_21996,N_20169,N_20293);
xor U21997 (N_21997,N_19649,N_19316);
and U21998 (N_21998,N_18403,N_19963);
or U21999 (N_21999,N_20804,N_18297);
nor U22000 (N_22000,N_19190,N_18544);
and U22001 (N_22001,N_19970,N_18280);
nand U22002 (N_22002,N_18757,N_18085);
or U22003 (N_22003,N_18252,N_19741);
and U22004 (N_22004,N_20116,N_18829);
xnor U22005 (N_22005,N_18908,N_18745);
nand U22006 (N_22006,N_20908,N_20872);
nand U22007 (N_22007,N_20559,N_20145);
xor U22008 (N_22008,N_19977,N_20158);
xnor U22009 (N_22009,N_19878,N_18554);
or U22010 (N_22010,N_20414,N_18411);
xnor U22011 (N_22011,N_18617,N_20732);
nand U22012 (N_22012,N_19734,N_19964);
or U22013 (N_22013,N_18848,N_19824);
and U22014 (N_22014,N_19885,N_20423);
and U22015 (N_22015,N_20392,N_18506);
or U22016 (N_22016,N_19481,N_19396);
nand U22017 (N_22017,N_20440,N_19278);
and U22018 (N_22018,N_18475,N_19020);
xnor U22019 (N_22019,N_18640,N_18152);
xor U22020 (N_22020,N_19040,N_18987);
nor U22021 (N_22021,N_19290,N_20068);
or U22022 (N_22022,N_19052,N_19750);
or U22023 (N_22023,N_20404,N_19329);
xor U22024 (N_22024,N_19311,N_18393);
xor U22025 (N_22025,N_18614,N_19853);
or U22026 (N_22026,N_18285,N_18125);
or U22027 (N_22027,N_19324,N_19410);
and U22028 (N_22028,N_19677,N_18258);
nor U22029 (N_22029,N_18890,N_19075);
and U22030 (N_22030,N_18664,N_19792);
and U22031 (N_22031,N_19552,N_19255);
nand U22032 (N_22032,N_20050,N_18868);
nand U22033 (N_22033,N_20966,N_19467);
xnor U22034 (N_22034,N_18778,N_19735);
xnor U22035 (N_22035,N_19036,N_18020);
nand U22036 (N_22036,N_19443,N_18407);
nor U22037 (N_22037,N_19615,N_19850);
xor U22038 (N_22038,N_20692,N_19248);
xnor U22039 (N_22039,N_20016,N_18852);
xnor U22040 (N_22040,N_20562,N_20159);
or U22041 (N_22041,N_19485,N_18860);
nand U22042 (N_22042,N_19815,N_18755);
and U22043 (N_22043,N_18977,N_18100);
xor U22044 (N_22044,N_20312,N_20002);
xnor U22045 (N_22045,N_20967,N_19499);
xor U22046 (N_22046,N_20757,N_20253);
or U22047 (N_22047,N_19385,N_19142);
xor U22048 (N_22048,N_18832,N_20164);
xor U22049 (N_22049,N_19520,N_20895);
xor U22050 (N_22050,N_18013,N_19998);
and U22051 (N_22051,N_19147,N_20758);
nor U22052 (N_22052,N_19445,N_20803);
xnor U22053 (N_22053,N_19060,N_18750);
xnor U22054 (N_22054,N_20642,N_19169);
xor U22055 (N_22055,N_20593,N_18983);
xor U22056 (N_22056,N_20340,N_19718);
nand U22057 (N_22057,N_19518,N_19226);
xnor U22058 (N_22058,N_19945,N_18584);
xnor U22059 (N_22059,N_18145,N_19567);
xnor U22060 (N_22060,N_18251,N_19700);
nor U22061 (N_22061,N_18938,N_20624);
nor U22062 (N_22062,N_20125,N_19851);
nor U22063 (N_22063,N_20663,N_20133);
nand U22064 (N_22064,N_20126,N_19528);
or U22065 (N_22065,N_19668,N_20058);
nor U22066 (N_22066,N_18003,N_18918);
and U22067 (N_22067,N_19186,N_20326);
or U22068 (N_22068,N_19769,N_20718);
or U22069 (N_22069,N_20630,N_19917);
nor U22070 (N_22070,N_19844,N_20041);
nor U22071 (N_22071,N_19034,N_20078);
and U22072 (N_22072,N_18729,N_20727);
nand U22073 (N_22073,N_20767,N_20228);
nand U22074 (N_22074,N_19228,N_19990);
xor U22075 (N_22075,N_18996,N_18742);
xnor U22076 (N_22076,N_20991,N_19606);
and U22077 (N_22077,N_19227,N_18306);
xnor U22078 (N_22078,N_20300,N_18253);
xnor U22079 (N_22079,N_20843,N_18775);
xnor U22080 (N_22080,N_20708,N_20865);
and U22081 (N_22081,N_20063,N_18157);
nand U22082 (N_22082,N_19962,N_20906);
and U22083 (N_22083,N_19809,N_19218);
nand U22084 (N_22084,N_19803,N_20873);
and U22085 (N_22085,N_19621,N_20211);
nand U22086 (N_22086,N_20095,N_19334);
xor U22087 (N_22087,N_20132,N_18913);
or U22088 (N_22088,N_19359,N_19490);
xor U22089 (N_22089,N_20641,N_19465);
nor U22090 (N_22090,N_18694,N_20306);
and U22091 (N_22091,N_19701,N_20258);
xnor U22092 (N_22092,N_18107,N_18856);
xnor U22093 (N_22093,N_18464,N_20318);
xor U22094 (N_22094,N_19473,N_18255);
nor U22095 (N_22095,N_19942,N_19967);
or U22096 (N_22096,N_19825,N_18239);
nand U22097 (N_22097,N_20028,N_19153);
or U22098 (N_22098,N_19949,N_19869);
nand U22099 (N_22099,N_18558,N_18951);
nand U22100 (N_22100,N_19540,N_20904);
xnor U22101 (N_22101,N_20476,N_19728);
nand U22102 (N_22102,N_18917,N_20988);
nand U22103 (N_22103,N_19899,N_18180);
or U22104 (N_22104,N_19922,N_20462);
xnor U22105 (N_22105,N_20776,N_20120);
nand U22106 (N_22106,N_20046,N_20601);
or U22107 (N_22107,N_20926,N_19261);
and U22108 (N_22108,N_18650,N_20343);
or U22109 (N_22109,N_19783,N_18064);
nand U22110 (N_22110,N_20073,N_20291);
nor U22111 (N_22111,N_19415,N_20429);
xnor U22112 (N_22112,N_19208,N_18719);
and U22113 (N_22113,N_18054,N_20574);
nor U22114 (N_22114,N_20555,N_20387);
xor U22115 (N_22115,N_18510,N_20152);
or U22116 (N_22116,N_19183,N_18966);
and U22117 (N_22117,N_19870,N_19595);
nor U22118 (N_22118,N_20499,N_18269);
xor U22119 (N_22119,N_20459,N_18608);
nand U22120 (N_22120,N_19956,N_20413);
nand U22121 (N_22121,N_18254,N_20518);
or U22122 (N_22122,N_18758,N_18691);
nor U22123 (N_22123,N_19143,N_18961);
nor U22124 (N_22124,N_19113,N_18812);
nand U22125 (N_22125,N_18622,N_18835);
nor U22126 (N_22126,N_18921,N_18478);
nor U22127 (N_22127,N_18273,N_20303);
and U22128 (N_22128,N_19411,N_20357);
nand U22129 (N_22129,N_20625,N_20353);
nand U22130 (N_22130,N_20193,N_18410);
or U22131 (N_22131,N_20409,N_20769);
nor U22132 (N_22132,N_18838,N_18170);
nand U22133 (N_22133,N_18647,N_18806);
nor U22134 (N_22134,N_19819,N_20018);
xnor U22135 (N_22135,N_20112,N_18741);
xnor U22136 (N_22136,N_18126,N_19797);
nor U22137 (N_22137,N_18435,N_20113);
nor U22138 (N_22138,N_19932,N_18175);
nor U22139 (N_22139,N_20744,N_20108);
nand U22140 (N_22140,N_20014,N_18104);
and U22141 (N_22141,N_20780,N_19566);
and U22142 (N_22142,N_18738,N_19493);
or U22143 (N_22143,N_19430,N_18362);
xor U22144 (N_22144,N_20400,N_20262);
nor U22145 (N_22145,N_19375,N_18332);
xor U22146 (N_22146,N_20761,N_20695);
nor U22147 (N_22147,N_20504,N_19273);
nand U22148 (N_22148,N_18368,N_18597);
and U22149 (N_22149,N_20267,N_20900);
nor U22150 (N_22150,N_20100,N_20438);
xor U22151 (N_22151,N_20210,N_18734);
or U22152 (N_22152,N_20428,N_18006);
nand U22153 (N_22153,N_20466,N_19161);
nand U22154 (N_22154,N_19217,N_19591);
nand U22155 (N_22155,N_18074,N_18724);
or U22156 (N_22156,N_18621,N_19450);
xor U22157 (N_22157,N_18718,N_18361);
nand U22158 (N_22158,N_20891,N_18187);
xor U22159 (N_22159,N_18241,N_18473);
xor U22160 (N_22160,N_20806,N_18249);
or U22161 (N_22161,N_19931,N_20686);
xor U22162 (N_22162,N_19554,N_19030);
or U22163 (N_22163,N_20407,N_20500);
and U22164 (N_22164,N_20597,N_20093);
xor U22165 (N_22165,N_18770,N_20505);
or U22166 (N_22166,N_19019,N_18796);
xor U22167 (N_22167,N_19327,N_18959);
nand U22168 (N_22168,N_18083,N_19755);
nor U22169 (N_22169,N_19017,N_19048);
nand U22170 (N_22170,N_19906,N_19781);
or U22171 (N_22171,N_19827,N_18434);
or U22172 (N_22172,N_20634,N_19818);
or U22173 (N_22173,N_20047,N_20880);
nand U22174 (N_22174,N_19146,N_19247);
and U22175 (N_22175,N_20271,N_19078);
xor U22176 (N_22176,N_18949,N_20001);
nand U22177 (N_22177,N_18416,N_18396);
nor U22178 (N_22178,N_18749,N_18016);
nor U22179 (N_22179,N_19196,N_20655);
and U22180 (N_22180,N_20564,N_18164);
nor U22181 (N_22181,N_20721,N_20481);
or U22182 (N_22182,N_18610,N_18242);
and U22183 (N_22183,N_19720,N_18392);
nand U22184 (N_22184,N_19271,N_18774);
or U22185 (N_22185,N_19578,N_18437);
xnor U22186 (N_22186,N_20207,N_19752);
xor U22187 (N_22187,N_18600,N_18731);
and U22188 (N_22188,N_18124,N_18299);
xor U22189 (N_22189,N_20448,N_20752);
and U22190 (N_22190,N_19550,N_18359);
nor U22191 (N_22191,N_18763,N_18712);
nor U22192 (N_22192,N_20706,N_19955);
nor U22193 (N_22193,N_19654,N_20369);
xor U22194 (N_22194,N_20653,N_19644);
xnor U22195 (N_22195,N_19370,N_19234);
and U22196 (N_22196,N_20209,N_20009);
nor U22197 (N_22197,N_19600,N_20627);
xor U22198 (N_22198,N_20178,N_20365);
nor U22199 (N_22199,N_20445,N_20573);
and U22200 (N_22200,N_18266,N_19399);
nand U22201 (N_22201,N_19369,N_19920);
or U22202 (N_22202,N_18789,N_20577);
and U22203 (N_22203,N_19837,N_18986);
and U22204 (N_22204,N_18566,N_19527);
and U22205 (N_22205,N_19704,N_18086);
xnor U22206 (N_22206,N_20534,N_18339);
xnor U22207 (N_22207,N_18894,N_20202);
or U22208 (N_22208,N_20963,N_20528);
and U22209 (N_22209,N_20270,N_20398);
or U22210 (N_22210,N_19817,N_18448);
nand U22211 (N_22211,N_19986,N_20356);
or U22212 (N_22212,N_20101,N_18373);
nor U22213 (N_22213,N_19659,N_20320);
nor U22214 (N_22214,N_18593,N_18680);
nor U22215 (N_22215,N_19349,N_18192);
nand U22216 (N_22216,N_18024,N_18666);
and U22217 (N_22217,N_19558,N_19152);
or U22218 (N_22218,N_19269,N_20664);
and U22219 (N_22219,N_20950,N_18068);
or U22220 (N_22220,N_20739,N_19405);
and U22221 (N_22221,N_19918,N_18322);
nor U22222 (N_22222,N_18695,N_20405);
and U22223 (N_22223,N_20076,N_18117);
xor U22224 (N_22224,N_20968,N_18500);
or U22225 (N_22225,N_19068,N_20773);
and U22226 (N_22226,N_18257,N_18516);
or U22227 (N_22227,N_20493,N_20189);
and U22228 (N_22228,N_20817,N_18779);
nor U22229 (N_22229,N_18648,N_18385);
xnor U22230 (N_22230,N_19893,N_19682);
or U22231 (N_22231,N_20280,N_19814);
nand U22232 (N_22232,N_18429,N_19057);
xor U22233 (N_22233,N_18946,N_20617);
xnor U22234 (N_22234,N_18331,N_19154);
nor U22235 (N_22235,N_20605,N_20283);
xnor U22236 (N_22236,N_19044,N_19344);
nand U22237 (N_22237,N_18586,N_19703);
xor U22238 (N_22238,N_18673,N_18398);
nand U22239 (N_22239,N_20622,N_18699);
nor U22240 (N_22240,N_19791,N_20432);
nand U22241 (N_22241,N_19372,N_18457);
nand U22242 (N_22242,N_18212,N_20294);
nor U22243 (N_22243,N_20542,N_20161);
nand U22244 (N_22244,N_18679,N_20185);
nor U22245 (N_22245,N_19077,N_20478);
xnor U22246 (N_22246,N_18538,N_20344);
xnor U22247 (N_22247,N_18697,N_18466);
and U22248 (N_22248,N_18366,N_19084);
and U22249 (N_22249,N_20890,N_19822);
nor U22250 (N_22250,N_20797,N_20123);
and U22251 (N_22251,N_20359,N_20728);
nor U22252 (N_22252,N_18102,N_20548);
xor U22253 (N_22253,N_20287,N_20444);
or U22254 (N_22254,N_19442,N_18620);
xnor U22255 (N_22255,N_19950,N_18490);
nor U22256 (N_22256,N_20683,N_19354);
xor U22257 (N_22257,N_18776,N_20902);
or U22258 (N_22258,N_20515,N_19921);
nand U22259 (N_22259,N_18037,N_20390);
and U22260 (N_22260,N_18082,N_18456);
xnor U22261 (N_22261,N_19842,N_19331);
and U22262 (N_22262,N_20213,N_18594);
nor U22263 (N_22263,N_18317,N_18363);
nor U22264 (N_22264,N_19318,N_19694);
or U22265 (N_22265,N_20905,N_20003);
nand U22266 (N_22266,N_20696,N_19076);
nand U22267 (N_22267,N_20031,N_19203);
and U22268 (N_22268,N_20847,N_19009);
or U22269 (N_22269,N_19338,N_20868);
xor U22270 (N_22270,N_19946,N_19759);
nor U22271 (N_22271,N_19989,N_20543);
and U22272 (N_22272,N_20034,N_18975);
xnor U22273 (N_22273,N_20864,N_20646);
xnor U22274 (N_22274,N_20497,N_19504);
nor U22275 (N_22275,N_20684,N_19303);
or U22276 (N_22276,N_20984,N_19515);
nor U22277 (N_22277,N_20733,N_19891);
nor U22278 (N_22278,N_20871,N_19134);
nor U22279 (N_22279,N_19726,N_20917);
or U22280 (N_22280,N_20450,N_18575);
nand U22281 (N_22281,N_19859,N_18522);
xor U22282 (N_22282,N_19509,N_19164);
xnor U22283 (N_22283,N_19381,N_19002);
nand U22284 (N_22284,N_20657,N_20969);
nor U22285 (N_22285,N_19418,N_20242);
xor U22286 (N_22286,N_19862,N_18318);
and U22287 (N_22287,N_20946,N_20252);
xor U22288 (N_22288,N_20308,N_18798);
and U22289 (N_22289,N_18550,N_19948);
xor U22290 (N_22290,N_20778,N_20170);
and U22291 (N_22291,N_18227,N_19776);
and U22292 (N_22292,N_20036,N_20723);
xor U22293 (N_22293,N_18427,N_19655);
xnor U22294 (N_22294,N_18226,N_20411);
nor U22295 (N_22295,N_19785,N_20465);
and U22296 (N_22296,N_20464,N_19588);
or U22297 (N_22297,N_18010,N_20722);
or U22298 (N_22298,N_19648,N_19664);
and U22299 (N_22299,N_19292,N_20822);
and U22300 (N_22300,N_19875,N_19046);
or U22301 (N_22301,N_20903,N_20694);
and U22302 (N_22302,N_19350,N_20659);
nand U22303 (N_22303,N_18819,N_19494);
nand U22304 (N_22304,N_20406,N_18503);
or U22305 (N_22305,N_19730,N_19758);
or U22306 (N_22306,N_20572,N_18487);
or U22307 (N_22307,N_20587,N_20943);
xnor U22308 (N_22308,N_18539,N_18369);
and U22309 (N_22309,N_20416,N_19216);
nor U22310 (N_22310,N_18430,N_18981);
nand U22311 (N_22311,N_18867,N_20689);
or U22312 (N_22312,N_20825,N_20750);
nand U22313 (N_22313,N_18217,N_20815);
nand U22314 (N_22314,N_19432,N_18132);
or U22315 (N_22315,N_20319,N_19601);
or U22316 (N_22316,N_20711,N_19987);
nor U22317 (N_22317,N_18201,N_19214);
nor U22318 (N_22318,N_18413,N_18298);
or U22319 (N_22319,N_19674,N_19858);
or U22320 (N_22320,N_20166,N_20647);
and U22321 (N_22321,N_19502,N_19966);
nor U22322 (N_22322,N_18372,N_20746);
xor U22323 (N_22323,N_20139,N_20522);
nor U22324 (N_22324,N_20730,N_20802);
or U22325 (N_22325,N_20079,N_18181);
nor U22326 (N_22326,N_19352,N_18123);
and U22327 (N_22327,N_18391,N_19620);
xor U22328 (N_22328,N_20082,N_19943);
xnor U22329 (N_22329,N_18281,N_20243);
or U22330 (N_22330,N_18501,N_18955);
nor U22331 (N_22331,N_18845,N_19242);
or U22332 (N_22332,N_20285,N_19265);
nand U22333 (N_22333,N_18497,N_18216);
and U22334 (N_22334,N_20592,N_18710);
xnor U22335 (N_22335,N_19116,N_19336);
or U22336 (N_22336,N_20848,N_19939);
and U22337 (N_22337,N_20571,N_20932);
or U22338 (N_22338,N_18716,N_18768);
or U22339 (N_22339,N_18060,N_19562);
or U22340 (N_22340,N_20064,N_20396);
nor U22341 (N_22341,N_20913,N_18418);
nand U22342 (N_22342,N_18007,N_18940);
and U22343 (N_22343,N_20299,N_19049);
and U22344 (N_22344,N_18821,N_19640);
or U22345 (N_22345,N_18642,N_20273);
nand U22346 (N_22346,N_19378,N_19055);
nand U22347 (N_22347,N_18270,N_20153);
and U22348 (N_22348,N_18376,N_20606);
xor U22349 (N_22349,N_19753,N_20838);
or U22350 (N_22350,N_18963,N_19821);
and U22351 (N_22351,N_19041,N_20660);
and U22352 (N_22352,N_18926,N_18063);
xor U22353 (N_22353,N_19124,N_20194);
or U22354 (N_22354,N_20501,N_20896);
and U22355 (N_22355,N_19082,N_18556);
xor U22356 (N_22356,N_19362,N_20458);
xor U22357 (N_22357,N_20417,N_20519);
xnor U22358 (N_22358,N_19397,N_18347);
nor U22359 (N_22359,N_20764,N_18381);
xor U22360 (N_22360,N_19006,N_20037);
nand U22361 (N_22361,N_18660,N_19828);
and U22362 (N_22362,N_18031,N_20096);
nor U22363 (N_22363,N_18479,N_19599);
nor U22364 (N_22364,N_18040,N_18171);
or U22365 (N_22365,N_19614,N_19816);
and U22366 (N_22366,N_19861,N_18307);
nor U22367 (N_22367,N_19868,N_20643);
and U22368 (N_22368,N_20668,N_19038);
and U22369 (N_22369,N_20149,N_18589);
or U22370 (N_22370,N_19238,N_20772);
and U22371 (N_22371,N_20437,N_19594);
xnor U22372 (N_22372,N_19863,N_19841);
and U22373 (N_22373,N_18931,N_18714);
xor U22374 (N_22374,N_20144,N_18529);
nand U22375 (N_22375,N_18311,N_20602);
nor U22376 (N_22376,N_19198,N_18205);
xnor U22377 (N_22377,N_20040,N_20277);
and U22378 (N_22378,N_18402,N_18521);
nor U22379 (N_22379,N_18162,N_18979);
or U22380 (N_22380,N_18055,N_19609);
and U22381 (N_22381,N_18924,N_18668);
nand U22382 (N_22382,N_20290,N_19856);
or U22383 (N_22383,N_18761,N_18872);
nand U22384 (N_22384,N_19245,N_19925);
nor U22385 (N_22385,N_19727,N_20386);
and U22386 (N_22386,N_19691,N_20938);
or U22387 (N_22387,N_19696,N_19656);
or U22388 (N_22388,N_20065,N_20833);
or U22389 (N_22389,N_19185,N_18039);
or U22390 (N_22390,N_20304,N_18260);
nor U22391 (N_22391,N_20447,N_20227);
nor U22392 (N_22392,N_18314,N_19433);
nand U22393 (N_22393,N_20339,N_19069);
and U22394 (N_22394,N_20841,N_19729);
nand U22395 (N_22395,N_19926,N_18070);
or U22396 (N_22396,N_20934,N_18291);
or U22397 (N_22397,N_19480,N_18715);
nand U22398 (N_22398,N_19321,N_19812);
and U22399 (N_22399,N_18992,N_18952);
or U22400 (N_22400,N_18476,N_19322);
xnor U22401 (N_22401,N_18569,N_19122);
xnor U22402 (N_22402,N_19400,N_20649);
or U22403 (N_22403,N_19721,N_19536);
and U22404 (N_22404,N_18084,N_19954);
nor U22405 (N_22405,N_19768,N_19476);
nor U22406 (N_22406,N_19205,N_20929);
or U22407 (N_22407,N_18973,N_20364);
nand U22408 (N_22408,N_19107,N_19909);
or U22409 (N_22409,N_18891,N_20171);
and U22410 (N_22410,N_18865,N_18465);
and U22411 (N_22411,N_20629,N_18492);
xnor U22412 (N_22412,N_20122,N_18019);
or U22413 (N_22413,N_20131,N_20556);
nand U22414 (N_22414,N_18905,N_20434);
xor U22415 (N_22415,N_18034,N_19653);
and U22416 (N_22416,N_18142,N_18474);
nor U22417 (N_22417,N_20672,N_20738);
or U22418 (N_22418,N_18772,N_18507);
xor U22419 (N_22419,N_18300,N_19689);
nand U22420 (N_22420,N_18390,N_18328);
nand U22421 (N_22421,N_19486,N_18388);
nor U22422 (N_22422,N_18826,N_18871);
xor U22423 (N_22423,N_20632,N_18333);
nand U22424 (N_22424,N_18581,N_18246);
and U22425 (N_22425,N_20042,N_18553);
or U22426 (N_22426,N_19881,N_20567);
nor U22427 (N_22427,N_19770,N_18432);
xnor U22428 (N_22428,N_19310,N_18035);
and U22429 (N_22429,N_18367,N_20996);
nor U22430 (N_22430,N_18053,N_20961);
or U22431 (N_22431,N_18762,N_20355);
or U22432 (N_22432,N_18800,N_18023);
or U22433 (N_22433,N_18168,N_19716);
xnor U22434 (N_22434,N_19719,N_20103);
nor U22435 (N_22435,N_19207,N_18268);
nand U22436 (N_22436,N_19592,N_18015);
nand U22437 (N_22437,N_18165,N_20586);
or U22438 (N_22438,N_20512,N_18615);
nand U22439 (N_22439,N_20869,N_18502);
nand U22440 (N_22440,N_20269,N_18794);
and U22441 (N_22441,N_19992,N_18394);
xor U22442 (N_22442,N_19210,N_19873);
nand U22443 (N_22443,N_20973,N_20965);
and U22444 (N_22444,N_19180,N_20330);
nand U22445 (N_22445,N_19723,N_18793);
nor U22446 (N_22446,N_19103,N_19882);
or U22447 (N_22447,N_20219,N_20807);
and U22448 (N_22448,N_20682,N_20027);
nand U22449 (N_22449,N_18799,N_18348);
and U22450 (N_22450,N_20976,N_20741);
xor U22451 (N_22451,N_18105,N_20251);
nor U22452 (N_22452,N_20536,N_19328);
and U22453 (N_22453,N_18769,N_20427);
nor U22454 (N_22454,N_18723,N_20742);
nor U22455 (N_22455,N_20025,N_19912);
and U22456 (N_22456,N_20551,N_19457);
nand U22457 (N_22457,N_18303,N_18079);
nor U22458 (N_22458,N_18730,N_18356);
or U22459 (N_22459,N_19883,N_19441);
nand U22460 (N_22460,N_18406,N_19808);
xnor U22461 (N_22461,N_18628,N_18485);
and U22462 (N_22462,N_19625,N_20477);
or U22463 (N_22463,N_19371,N_18711);
and U22464 (N_22464,N_20635,N_19717);
nand U22465 (N_22465,N_18809,N_20109);
or U22466 (N_22466,N_20960,N_18568);
nand U22467 (N_22467,N_18631,N_19607);
xor U22468 (N_22468,N_20651,N_18603);
nor U22469 (N_22469,N_20785,N_20203);
nand U22470 (N_22470,N_19299,N_18228);
nor U22471 (N_22471,N_20468,N_18294);
xnor U22472 (N_22472,N_19968,N_19072);
xor U22473 (N_22473,N_20765,N_20626);
nand U22474 (N_22474,N_20221,N_19632);
or U22475 (N_22475,N_20165,N_19802);
nor U22476 (N_22476,N_20952,N_19641);
xor U22477 (N_22477,N_20216,N_18358);
nand U22478 (N_22478,N_20307,N_19171);
xor U22479 (N_22479,N_20639,N_19830);
or U22480 (N_22480,N_20206,N_19326);
and U22481 (N_22481,N_18425,N_20012);
nand U22482 (N_22482,N_20831,N_20137);
xor U22483 (N_22483,N_19221,N_19151);
nor U22484 (N_22484,N_19738,N_19697);
nand U22485 (N_22485,N_20747,N_19979);
nand U22486 (N_22486,N_18803,N_19200);
nand U22487 (N_22487,N_19997,N_19096);
nand U22488 (N_22488,N_20604,N_20422);
nand U22489 (N_22489,N_19272,N_18618);
nor U22490 (N_22490,N_19158,N_18839);
and U22491 (N_22491,N_18195,N_18514);
nand U22492 (N_22492,N_19865,N_19847);
and U22493 (N_22493,N_19280,N_19281);
nor U22494 (N_22494,N_20860,N_19892);
or U22495 (N_22495,N_18925,N_20823);
xnor U22496 (N_22496,N_19320,N_18424);
nor U22497 (N_22497,N_19673,N_18112);
or U22498 (N_22498,N_19064,N_18899);
nand U22499 (N_22499,N_20000,N_18995);
xnor U22500 (N_22500,N_19651,N_18860);
xor U22501 (N_22501,N_18358,N_18185);
and U22502 (N_22502,N_18563,N_18544);
xnor U22503 (N_22503,N_18719,N_18402);
nor U22504 (N_22504,N_20684,N_20963);
nor U22505 (N_22505,N_18989,N_19193);
or U22506 (N_22506,N_20652,N_20339);
nand U22507 (N_22507,N_18458,N_19630);
or U22508 (N_22508,N_20097,N_18030);
and U22509 (N_22509,N_18808,N_20888);
nor U22510 (N_22510,N_18926,N_20356);
nor U22511 (N_22511,N_18516,N_18209);
and U22512 (N_22512,N_19276,N_18138);
nand U22513 (N_22513,N_19426,N_20243);
or U22514 (N_22514,N_19994,N_20646);
or U22515 (N_22515,N_20333,N_19382);
and U22516 (N_22516,N_18099,N_18653);
xor U22517 (N_22517,N_20691,N_18399);
nand U22518 (N_22518,N_20184,N_19893);
nand U22519 (N_22519,N_18113,N_18285);
nand U22520 (N_22520,N_18019,N_19721);
xnor U22521 (N_22521,N_19346,N_20907);
nor U22522 (N_22522,N_18030,N_19632);
or U22523 (N_22523,N_19183,N_19096);
or U22524 (N_22524,N_18838,N_19162);
and U22525 (N_22525,N_18695,N_20257);
nand U22526 (N_22526,N_20071,N_20143);
nor U22527 (N_22527,N_19469,N_18500);
nand U22528 (N_22528,N_19025,N_20861);
and U22529 (N_22529,N_18019,N_20438);
and U22530 (N_22530,N_19430,N_20601);
and U22531 (N_22531,N_19317,N_18805);
xor U22532 (N_22532,N_20872,N_19822);
xor U22533 (N_22533,N_20889,N_18803);
and U22534 (N_22534,N_19164,N_18235);
nor U22535 (N_22535,N_18589,N_20509);
nand U22536 (N_22536,N_19207,N_20642);
or U22537 (N_22537,N_18072,N_19582);
nand U22538 (N_22538,N_20373,N_19051);
and U22539 (N_22539,N_20217,N_19109);
xor U22540 (N_22540,N_18151,N_18243);
nor U22541 (N_22541,N_19836,N_18160);
xor U22542 (N_22542,N_19827,N_19277);
nor U22543 (N_22543,N_18575,N_20389);
or U22544 (N_22544,N_19839,N_20329);
nand U22545 (N_22545,N_20648,N_20570);
nand U22546 (N_22546,N_20551,N_20414);
xor U22547 (N_22547,N_18371,N_19584);
nor U22548 (N_22548,N_18164,N_18975);
and U22549 (N_22549,N_18884,N_20806);
nand U22550 (N_22550,N_19622,N_20340);
nand U22551 (N_22551,N_20069,N_19301);
nand U22552 (N_22552,N_18049,N_19129);
nor U22553 (N_22553,N_18310,N_20308);
nand U22554 (N_22554,N_19546,N_20320);
and U22555 (N_22555,N_19690,N_19660);
nand U22556 (N_22556,N_19961,N_20732);
nor U22557 (N_22557,N_20230,N_20482);
nor U22558 (N_22558,N_19719,N_19099);
xor U22559 (N_22559,N_19722,N_20021);
nor U22560 (N_22560,N_18479,N_19534);
nor U22561 (N_22561,N_18952,N_19331);
nand U22562 (N_22562,N_18387,N_20082);
xor U22563 (N_22563,N_19410,N_19207);
or U22564 (N_22564,N_20059,N_19755);
and U22565 (N_22565,N_20647,N_19826);
or U22566 (N_22566,N_19180,N_19380);
and U22567 (N_22567,N_19885,N_18276);
or U22568 (N_22568,N_19451,N_18324);
xnor U22569 (N_22569,N_18262,N_19187);
nor U22570 (N_22570,N_19580,N_18736);
nor U22571 (N_22571,N_20746,N_19053);
and U22572 (N_22572,N_20474,N_19513);
nor U22573 (N_22573,N_19634,N_18673);
nor U22574 (N_22574,N_18282,N_18303);
xor U22575 (N_22575,N_19872,N_20586);
nand U22576 (N_22576,N_20211,N_20634);
or U22577 (N_22577,N_20759,N_18184);
nand U22578 (N_22578,N_18542,N_19449);
nand U22579 (N_22579,N_18691,N_19525);
xor U22580 (N_22580,N_19262,N_18094);
nor U22581 (N_22581,N_18292,N_20918);
and U22582 (N_22582,N_19512,N_18420);
or U22583 (N_22583,N_20410,N_18685);
or U22584 (N_22584,N_19311,N_18915);
nand U22585 (N_22585,N_18122,N_20596);
or U22586 (N_22586,N_19968,N_20896);
nand U22587 (N_22587,N_20248,N_18674);
nor U22588 (N_22588,N_20832,N_20431);
xnor U22589 (N_22589,N_19687,N_18745);
nor U22590 (N_22590,N_18417,N_19485);
nand U22591 (N_22591,N_18049,N_18411);
nand U22592 (N_22592,N_18349,N_19169);
nand U22593 (N_22593,N_20255,N_20207);
nor U22594 (N_22594,N_18052,N_20665);
or U22595 (N_22595,N_18428,N_18100);
and U22596 (N_22596,N_20133,N_20556);
nor U22597 (N_22597,N_19596,N_20938);
and U22598 (N_22598,N_19931,N_19041);
and U22599 (N_22599,N_20243,N_18872);
xor U22600 (N_22600,N_18457,N_20264);
and U22601 (N_22601,N_20694,N_20689);
nand U22602 (N_22602,N_18502,N_18760);
nor U22603 (N_22603,N_18752,N_18091);
xnor U22604 (N_22604,N_18323,N_20389);
and U22605 (N_22605,N_18124,N_19745);
nand U22606 (N_22606,N_20887,N_18282);
xnor U22607 (N_22607,N_18368,N_19274);
nor U22608 (N_22608,N_18898,N_20516);
or U22609 (N_22609,N_20245,N_19940);
xnor U22610 (N_22610,N_20708,N_18286);
nand U22611 (N_22611,N_19583,N_18529);
or U22612 (N_22612,N_20832,N_19487);
nand U22613 (N_22613,N_19992,N_19168);
and U22614 (N_22614,N_18234,N_18701);
xnor U22615 (N_22615,N_19869,N_20418);
or U22616 (N_22616,N_18375,N_19432);
xor U22617 (N_22617,N_18927,N_18287);
or U22618 (N_22618,N_19632,N_19556);
nor U22619 (N_22619,N_18186,N_19631);
nand U22620 (N_22620,N_18308,N_18079);
nor U22621 (N_22621,N_20554,N_19756);
nor U22622 (N_22622,N_19788,N_18678);
and U22623 (N_22623,N_18861,N_18282);
nand U22624 (N_22624,N_19441,N_18686);
nand U22625 (N_22625,N_20330,N_20726);
nand U22626 (N_22626,N_19566,N_18951);
xor U22627 (N_22627,N_18660,N_19098);
xor U22628 (N_22628,N_19136,N_18128);
nand U22629 (N_22629,N_18798,N_20108);
nor U22630 (N_22630,N_20650,N_18075);
nand U22631 (N_22631,N_18157,N_20980);
nand U22632 (N_22632,N_18202,N_20562);
or U22633 (N_22633,N_19513,N_18569);
or U22634 (N_22634,N_18289,N_20797);
xor U22635 (N_22635,N_20827,N_20004);
and U22636 (N_22636,N_20243,N_20726);
or U22637 (N_22637,N_19932,N_18338);
xnor U22638 (N_22638,N_18068,N_20920);
or U22639 (N_22639,N_20803,N_19199);
and U22640 (N_22640,N_20860,N_19724);
nor U22641 (N_22641,N_19761,N_20002);
xor U22642 (N_22642,N_18368,N_18106);
nand U22643 (N_22643,N_18625,N_19107);
or U22644 (N_22644,N_18044,N_18698);
and U22645 (N_22645,N_19935,N_18345);
xnor U22646 (N_22646,N_19290,N_18835);
or U22647 (N_22647,N_20468,N_18453);
or U22648 (N_22648,N_18491,N_20173);
xnor U22649 (N_22649,N_20525,N_20063);
nor U22650 (N_22650,N_18777,N_18038);
nor U22651 (N_22651,N_19516,N_20872);
nor U22652 (N_22652,N_19322,N_19495);
nor U22653 (N_22653,N_19607,N_19129);
or U22654 (N_22654,N_18567,N_20097);
xor U22655 (N_22655,N_19801,N_20343);
xnor U22656 (N_22656,N_19834,N_19928);
or U22657 (N_22657,N_20743,N_20803);
or U22658 (N_22658,N_20899,N_19586);
nand U22659 (N_22659,N_20494,N_18059);
or U22660 (N_22660,N_20838,N_19404);
nor U22661 (N_22661,N_19495,N_20223);
nor U22662 (N_22662,N_20941,N_19689);
and U22663 (N_22663,N_19300,N_18877);
or U22664 (N_22664,N_20024,N_18460);
and U22665 (N_22665,N_19355,N_20844);
xor U22666 (N_22666,N_20101,N_19604);
nor U22667 (N_22667,N_19113,N_19219);
or U22668 (N_22668,N_20074,N_20851);
and U22669 (N_22669,N_19719,N_18271);
or U22670 (N_22670,N_18948,N_19565);
or U22671 (N_22671,N_19699,N_19224);
xor U22672 (N_22672,N_19082,N_19190);
and U22673 (N_22673,N_18356,N_18055);
nand U22674 (N_22674,N_19869,N_20611);
and U22675 (N_22675,N_20823,N_18334);
or U22676 (N_22676,N_19067,N_18258);
and U22677 (N_22677,N_19763,N_18226);
and U22678 (N_22678,N_20648,N_18337);
and U22679 (N_22679,N_20020,N_20389);
nand U22680 (N_22680,N_19777,N_20589);
or U22681 (N_22681,N_20939,N_19653);
and U22682 (N_22682,N_18071,N_20206);
xnor U22683 (N_22683,N_19854,N_19954);
or U22684 (N_22684,N_20042,N_18095);
xnor U22685 (N_22685,N_19446,N_18929);
xnor U22686 (N_22686,N_19252,N_18129);
and U22687 (N_22687,N_18167,N_18376);
and U22688 (N_22688,N_20327,N_20139);
or U22689 (N_22689,N_18922,N_20362);
nor U22690 (N_22690,N_18283,N_19078);
and U22691 (N_22691,N_20763,N_19654);
and U22692 (N_22692,N_19997,N_19469);
nand U22693 (N_22693,N_19247,N_20110);
and U22694 (N_22694,N_20706,N_18115);
and U22695 (N_22695,N_20526,N_19472);
and U22696 (N_22696,N_20726,N_19000);
or U22697 (N_22697,N_19950,N_18373);
nand U22698 (N_22698,N_20106,N_18607);
xnor U22699 (N_22699,N_20955,N_20139);
or U22700 (N_22700,N_18386,N_20171);
and U22701 (N_22701,N_18408,N_19299);
and U22702 (N_22702,N_19435,N_20330);
and U22703 (N_22703,N_18178,N_18456);
or U22704 (N_22704,N_18311,N_18151);
or U22705 (N_22705,N_19473,N_18377);
and U22706 (N_22706,N_19597,N_20066);
or U22707 (N_22707,N_19129,N_20256);
or U22708 (N_22708,N_18668,N_18629);
nor U22709 (N_22709,N_18980,N_20571);
xnor U22710 (N_22710,N_19238,N_20318);
and U22711 (N_22711,N_19762,N_18467);
nor U22712 (N_22712,N_20546,N_20206);
and U22713 (N_22713,N_18668,N_19792);
and U22714 (N_22714,N_20898,N_20629);
nand U22715 (N_22715,N_20531,N_19070);
and U22716 (N_22716,N_19003,N_20627);
or U22717 (N_22717,N_20146,N_19082);
xor U22718 (N_22718,N_19814,N_18279);
nand U22719 (N_22719,N_20093,N_19926);
and U22720 (N_22720,N_18982,N_20376);
nor U22721 (N_22721,N_19167,N_20476);
or U22722 (N_22722,N_19259,N_18292);
nor U22723 (N_22723,N_20075,N_20703);
nor U22724 (N_22724,N_18657,N_18513);
nand U22725 (N_22725,N_20734,N_18880);
or U22726 (N_22726,N_20629,N_20437);
or U22727 (N_22727,N_19697,N_20467);
xor U22728 (N_22728,N_18830,N_20243);
and U22729 (N_22729,N_20677,N_18064);
and U22730 (N_22730,N_18306,N_18949);
nor U22731 (N_22731,N_18802,N_19186);
nand U22732 (N_22732,N_18154,N_20480);
xor U22733 (N_22733,N_20579,N_18854);
xnor U22734 (N_22734,N_20176,N_19938);
xnor U22735 (N_22735,N_20468,N_19284);
and U22736 (N_22736,N_20140,N_19549);
or U22737 (N_22737,N_18417,N_19640);
and U22738 (N_22738,N_19987,N_18199);
or U22739 (N_22739,N_19524,N_20029);
nor U22740 (N_22740,N_19209,N_20830);
nor U22741 (N_22741,N_19577,N_18908);
xor U22742 (N_22742,N_18164,N_19222);
xor U22743 (N_22743,N_18195,N_19243);
nor U22744 (N_22744,N_19268,N_18094);
nor U22745 (N_22745,N_19017,N_20201);
xor U22746 (N_22746,N_18777,N_18949);
nor U22747 (N_22747,N_20248,N_20611);
nor U22748 (N_22748,N_20988,N_18731);
nor U22749 (N_22749,N_19736,N_20722);
xor U22750 (N_22750,N_20683,N_20234);
xor U22751 (N_22751,N_18456,N_20078);
nand U22752 (N_22752,N_19908,N_18340);
and U22753 (N_22753,N_18998,N_18248);
nand U22754 (N_22754,N_20547,N_18370);
and U22755 (N_22755,N_20056,N_19931);
xnor U22756 (N_22756,N_18685,N_19882);
nor U22757 (N_22757,N_20757,N_18240);
nor U22758 (N_22758,N_18009,N_19123);
xor U22759 (N_22759,N_18314,N_20087);
or U22760 (N_22760,N_20636,N_18245);
xnor U22761 (N_22761,N_20994,N_20770);
nand U22762 (N_22762,N_18141,N_20661);
nor U22763 (N_22763,N_18045,N_18491);
xor U22764 (N_22764,N_19046,N_18784);
nand U22765 (N_22765,N_19759,N_18149);
nor U22766 (N_22766,N_19333,N_18101);
xnor U22767 (N_22767,N_19989,N_19606);
nand U22768 (N_22768,N_19938,N_18661);
or U22769 (N_22769,N_19608,N_20794);
xnor U22770 (N_22770,N_18190,N_20582);
or U22771 (N_22771,N_20678,N_18425);
nand U22772 (N_22772,N_19605,N_18293);
or U22773 (N_22773,N_19818,N_19683);
nand U22774 (N_22774,N_20439,N_20336);
nor U22775 (N_22775,N_20041,N_20665);
xor U22776 (N_22776,N_18295,N_18351);
nor U22777 (N_22777,N_18595,N_20636);
xnor U22778 (N_22778,N_19788,N_19124);
or U22779 (N_22779,N_18936,N_20134);
or U22780 (N_22780,N_19983,N_18079);
xor U22781 (N_22781,N_20072,N_20280);
nand U22782 (N_22782,N_18418,N_19730);
nor U22783 (N_22783,N_18073,N_18072);
nor U22784 (N_22784,N_20779,N_18291);
and U22785 (N_22785,N_18183,N_19961);
nand U22786 (N_22786,N_19177,N_19068);
and U22787 (N_22787,N_20957,N_19224);
xnor U22788 (N_22788,N_20194,N_20603);
or U22789 (N_22789,N_18853,N_20357);
xnor U22790 (N_22790,N_19182,N_18556);
or U22791 (N_22791,N_20644,N_20711);
or U22792 (N_22792,N_19976,N_18755);
nor U22793 (N_22793,N_19046,N_20453);
xnor U22794 (N_22794,N_18331,N_19593);
nand U22795 (N_22795,N_18604,N_18878);
nand U22796 (N_22796,N_20474,N_18727);
or U22797 (N_22797,N_19858,N_19921);
nand U22798 (N_22798,N_19229,N_18869);
xor U22799 (N_22799,N_19086,N_18863);
and U22800 (N_22800,N_18243,N_18473);
and U22801 (N_22801,N_19292,N_20117);
and U22802 (N_22802,N_20390,N_19862);
and U22803 (N_22803,N_19022,N_20274);
or U22804 (N_22804,N_18505,N_18708);
and U22805 (N_22805,N_20368,N_19154);
nand U22806 (N_22806,N_18797,N_20860);
and U22807 (N_22807,N_20019,N_20753);
nor U22808 (N_22808,N_19952,N_20787);
nor U22809 (N_22809,N_19749,N_18118);
and U22810 (N_22810,N_19617,N_19167);
nor U22811 (N_22811,N_19186,N_19371);
nor U22812 (N_22812,N_19704,N_20062);
nor U22813 (N_22813,N_19443,N_19488);
or U22814 (N_22814,N_20373,N_19403);
nand U22815 (N_22815,N_20425,N_18689);
nand U22816 (N_22816,N_19807,N_20706);
or U22817 (N_22817,N_18282,N_19268);
and U22818 (N_22818,N_18589,N_20962);
xnor U22819 (N_22819,N_19552,N_19664);
or U22820 (N_22820,N_18672,N_19571);
xor U22821 (N_22821,N_20898,N_20444);
nand U22822 (N_22822,N_20559,N_18148);
xnor U22823 (N_22823,N_18672,N_19741);
nor U22824 (N_22824,N_20731,N_19779);
xnor U22825 (N_22825,N_20478,N_19503);
nor U22826 (N_22826,N_19068,N_18505);
and U22827 (N_22827,N_20978,N_18689);
nand U22828 (N_22828,N_19340,N_18072);
and U22829 (N_22829,N_20351,N_19822);
nor U22830 (N_22830,N_19580,N_19185);
nand U22831 (N_22831,N_20197,N_19053);
or U22832 (N_22832,N_18087,N_20777);
or U22833 (N_22833,N_20500,N_18713);
xnor U22834 (N_22834,N_19209,N_20708);
xnor U22835 (N_22835,N_20605,N_19880);
nand U22836 (N_22836,N_18084,N_18729);
or U22837 (N_22837,N_19556,N_20725);
or U22838 (N_22838,N_19437,N_19958);
nor U22839 (N_22839,N_18085,N_19117);
and U22840 (N_22840,N_18585,N_18498);
or U22841 (N_22841,N_20938,N_19267);
nand U22842 (N_22842,N_20198,N_20635);
and U22843 (N_22843,N_20436,N_20543);
xnor U22844 (N_22844,N_20096,N_19262);
and U22845 (N_22845,N_20997,N_18893);
or U22846 (N_22846,N_20454,N_18956);
and U22847 (N_22847,N_19936,N_19655);
or U22848 (N_22848,N_18722,N_18617);
xor U22849 (N_22849,N_18705,N_19668);
xnor U22850 (N_22850,N_18275,N_18253);
and U22851 (N_22851,N_19138,N_19283);
nand U22852 (N_22852,N_19616,N_19544);
or U22853 (N_22853,N_18588,N_20740);
and U22854 (N_22854,N_20120,N_20955);
or U22855 (N_22855,N_19469,N_20032);
nand U22856 (N_22856,N_20042,N_20692);
or U22857 (N_22857,N_18196,N_20225);
or U22858 (N_22858,N_18334,N_18356);
or U22859 (N_22859,N_19616,N_19410);
nor U22860 (N_22860,N_20607,N_19663);
nand U22861 (N_22861,N_18884,N_19212);
nand U22862 (N_22862,N_18333,N_18941);
xor U22863 (N_22863,N_18246,N_19985);
or U22864 (N_22864,N_19596,N_18081);
nand U22865 (N_22865,N_20530,N_19484);
and U22866 (N_22866,N_19725,N_18604);
and U22867 (N_22867,N_19924,N_18303);
xor U22868 (N_22868,N_18909,N_19721);
nand U22869 (N_22869,N_20347,N_19335);
and U22870 (N_22870,N_20041,N_18755);
or U22871 (N_22871,N_20575,N_20616);
nor U22872 (N_22872,N_18677,N_20906);
or U22873 (N_22873,N_20755,N_19955);
nor U22874 (N_22874,N_19078,N_20352);
nor U22875 (N_22875,N_20140,N_18791);
and U22876 (N_22876,N_19962,N_19791);
or U22877 (N_22877,N_19993,N_20203);
nand U22878 (N_22878,N_18184,N_18595);
nor U22879 (N_22879,N_20853,N_19801);
or U22880 (N_22880,N_20205,N_18784);
nand U22881 (N_22881,N_20409,N_20535);
xnor U22882 (N_22882,N_18340,N_19479);
nand U22883 (N_22883,N_18269,N_20835);
nand U22884 (N_22884,N_18458,N_19716);
nor U22885 (N_22885,N_19674,N_19088);
nand U22886 (N_22886,N_18110,N_19841);
or U22887 (N_22887,N_18844,N_19130);
xnor U22888 (N_22888,N_20565,N_20076);
and U22889 (N_22889,N_20226,N_18572);
nand U22890 (N_22890,N_18625,N_20118);
and U22891 (N_22891,N_20294,N_19838);
and U22892 (N_22892,N_18791,N_20671);
nor U22893 (N_22893,N_18924,N_18356);
xnor U22894 (N_22894,N_19333,N_18144);
xor U22895 (N_22895,N_18507,N_19314);
xor U22896 (N_22896,N_18098,N_19676);
and U22897 (N_22897,N_18662,N_18908);
or U22898 (N_22898,N_18718,N_19520);
nand U22899 (N_22899,N_20507,N_18656);
nor U22900 (N_22900,N_18440,N_19198);
xor U22901 (N_22901,N_20504,N_18101);
and U22902 (N_22902,N_18941,N_19101);
and U22903 (N_22903,N_19093,N_19772);
nand U22904 (N_22904,N_18848,N_20375);
nand U22905 (N_22905,N_20546,N_20127);
and U22906 (N_22906,N_19642,N_19793);
or U22907 (N_22907,N_18876,N_20186);
xnor U22908 (N_22908,N_20379,N_18625);
nor U22909 (N_22909,N_19661,N_18745);
and U22910 (N_22910,N_19523,N_18174);
and U22911 (N_22911,N_20234,N_19783);
nor U22912 (N_22912,N_20277,N_19747);
xnor U22913 (N_22913,N_20711,N_18282);
and U22914 (N_22914,N_18985,N_20103);
xor U22915 (N_22915,N_19632,N_19446);
xnor U22916 (N_22916,N_20069,N_18135);
nor U22917 (N_22917,N_19942,N_19235);
xor U22918 (N_22918,N_20139,N_18485);
xor U22919 (N_22919,N_19616,N_20722);
and U22920 (N_22920,N_19275,N_18928);
and U22921 (N_22921,N_19787,N_18945);
xnor U22922 (N_22922,N_20250,N_19973);
xor U22923 (N_22923,N_20881,N_18836);
and U22924 (N_22924,N_20383,N_19278);
nor U22925 (N_22925,N_19514,N_20771);
nor U22926 (N_22926,N_20904,N_18614);
and U22927 (N_22927,N_19933,N_20938);
and U22928 (N_22928,N_18179,N_19098);
or U22929 (N_22929,N_19831,N_20052);
nand U22930 (N_22930,N_20076,N_19669);
xnor U22931 (N_22931,N_20841,N_20394);
nand U22932 (N_22932,N_20482,N_20880);
nor U22933 (N_22933,N_18449,N_20306);
nand U22934 (N_22934,N_19851,N_19598);
nor U22935 (N_22935,N_20782,N_19563);
or U22936 (N_22936,N_20582,N_18320);
nand U22937 (N_22937,N_18384,N_19277);
nor U22938 (N_22938,N_18527,N_19790);
xnor U22939 (N_22939,N_20240,N_19605);
nor U22940 (N_22940,N_19413,N_18091);
nand U22941 (N_22941,N_18877,N_19372);
nand U22942 (N_22942,N_20795,N_18004);
nand U22943 (N_22943,N_19909,N_20251);
nand U22944 (N_22944,N_18862,N_18724);
nor U22945 (N_22945,N_18378,N_18727);
nand U22946 (N_22946,N_20686,N_20613);
nor U22947 (N_22947,N_18532,N_20786);
xnor U22948 (N_22948,N_20996,N_20318);
nand U22949 (N_22949,N_18934,N_20544);
nor U22950 (N_22950,N_19812,N_20127);
xnor U22951 (N_22951,N_19740,N_20958);
or U22952 (N_22952,N_19942,N_18525);
nor U22953 (N_22953,N_20565,N_19574);
xor U22954 (N_22954,N_19642,N_19459);
or U22955 (N_22955,N_20816,N_18872);
nor U22956 (N_22956,N_20015,N_20644);
or U22957 (N_22957,N_20074,N_20460);
xnor U22958 (N_22958,N_19148,N_19614);
or U22959 (N_22959,N_18623,N_18215);
and U22960 (N_22960,N_18783,N_20779);
nor U22961 (N_22961,N_20891,N_20459);
nor U22962 (N_22962,N_20846,N_18484);
nor U22963 (N_22963,N_18009,N_20367);
or U22964 (N_22964,N_19648,N_18398);
xor U22965 (N_22965,N_19201,N_18370);
or U22966 (N_22966,N_18157,N_19892);
or U22967 (N_22967,N_20507,N_19530);
nor U22968 (N_22968,N_18827,N_20347);
nor U22969 (N_22969,N_20741,N_19291);
and U22970 (N_22970,N_19239,N_18050);
xnor U22971 (N_22971,N_19864,N_18736);
nand U22972 (N_22972,N_18259,N_18115);
and U22973 (N_22973,N_19462,N_19931);
nor U22974 (N_22974,N_20822,N_20475);
nand U22975 (N_22975,N_20726,N_20295);
xnor U22976 (N_22976,N_19300,N_18503);
xnor U22977 (N_22977,N_20609,N_19921);
or U22978 (N_22978,N_19974,N_19896);
nor U22979 (N_22979,N_20721,N_20922);
nor U22980 (N_22980,N_18159,N_19481);
nor U22981 (N_22981,N_19521,N_20576);
nand U22982 (N_22982,N_20614,N_20193);
nand U22983 (N_22983,N_19391,N_20044);
or U22984 (N_22984,N_19936,N_18809);
nor U22985 (N_22985,N_20619,N_20454);
xnor U22986 (N_22986,N_18540,N_20474);
and U22987 (N_22987,N_18992,N_19531);
nor U22988 (N_22988,N_19255,N_19002);
or U22989 (N_22989,N_20505,N_19762);
xnor U22990 (N_22990,N_18467,N_18554);
or U22991 (N_22991,N_20387,N_18704);
xor U22992 (N_22992,N_18197,N_19651);
or U22993 (N_22993,N_20304,N_19661);
or U22994 (N_22994,N_18229,N_18663);
or U22995 (N_22995,N_20023,N_19255);
nor U22996 (N_22996,N_19687,N_20081);
nor U22997 (N_22997,N_20198,N_19292);
or U22998 (N_22998,N_20326,N_20909);
nor U22999 (N_22999,N_19313,N_19256);
nand U23000 (N_23000,N_20593,N_18504);
nand U23001 (N_23001,N_20739,N_19466);
nor U23002 (N_23002,N_20357,N_18130);
or U23003 (N_23003,N_18049,N_20834);
nor U23004 (N_23004,N_19939,N_20263);
nor U23005 (N_23005,N_18310,N_18479);
xor U23006 (N_23006,N_20196,N_19654);
and U23007 (N_23007,N_19045,N_20920);
nor U23008 (N_23008,N_18292,N_20250);
nand U23009 (N_23009,N_18941,N_18349);
or U23010 (N_23010,N_19223,N_20571);
xor U23011 (N_23011,N_18434,N_19108);
nand U23012 (N_23012,N_20302,N_19541);
xor U23013 (N_23013,N_18353,N_19245);
xor U23014 (N_23014,N_18149,N_18050);
nor U23015 (N_23015,N_20563,N_20693);
and U23016 (N_23016,N_20780,N_19738);
nor U23017 (N_23017,N_20414,N_18201);
nand U23018 (N_23018,N_18421,N_20139);
or U23019 (N_23019,N_20475,N_20957);
xnor U23020 (N_23020,N_19550,N_18233);
nand U23021 (N_23021,N_19737,N_20559);
nand U23022 (N_23022,N_19828,N_18829);
nand U23023 (N_23023,N_18368,N_20807);
and U23024 (N_23024,N_19949,N_20810);
xnor U23025 (N_23025,N_19469,N_19789);
nand U23026 (N_23026,N_19138,N_20343);
and U23027 (N_23027,N_19927,N_19925);
xnor U23028 (N_23028,N_18202,N_20539);
nand U23029 (N_23029,N_20994,N_18724);
xor U23030 (N_23030,N_20156,N_18820);
nor U23031 (N_23031,N_20039,N_18714);
and U23032 (N_23032,N_19773,N_19829);
xor U23033 (N_23033,N_19864,N_19921);
and U23034 (N_23034,N_19563,N_19134);
or U23035 (N_23035,N_19269,N_20382);
nor U23036 (N_23036,N_18899,N_18708);
and U23037 (N_23037,N_18607,N_19019);
xnor U23038 (N_23038,N_18376,N_19261);
or U23039 (N_23039,N_19808,N_20504);
and U23040 (N_23040,N_19294,N_20997);
and U23041 (N_23041,N_19426,N_18820);
and U23042 (N_23042,N_20059,N_18894);
xor U23043 (N_23043,N_18025,N_18658);
or U23044 (N_23044,N_20732,N_18018);
nand U23045 (N_23045,N_19883,N_20816);
nand U23046 (N_23046,N_18714,N_19956);
and U23047 (N_23047,N_19459,N_18256);
nor U23048 (N_23048,N_19173,N_20427);
or U23049 (N_23049,N_20251,N_18588);
and U23050 (N_23050,N_20026,N_18358);
nor U23051 (N_23051,N_20968,N_18004);
and U23052 (N_23052,N_18640,N_19852);
xnor U23053 (N_23053,N_18672,N_20184);
or U23054 (N_23054,N_20907,N_18278);
nor U23055 (N_23055,N_19359,N_18404);
and U23056 (N_23056,N_19230,N_20539);
xnor U23057 (N_23057,N_18002,N_19008);
xnor U23058 (N_23058,N_19299,N_20582);
xnor U23059 (N_23059,N_19427,N_20977);
nor U23060 (N_23060,N_18016,N_20445);
or U23061 (N_23061,N_20519,N_20541);
nand U23062 (N_23062,N_20355,N_20487);
nor U23063 (N_23063,N_20827,N_19145);
nor U23064 (N_23064,N_18953,N_18153);
nor U23065 (N_23065,N_19136,N_19310);
xnor U23066 (N_23066,N_19666,N_19363);
xor U23067 (N_23067,N_20984,N_20155);
or U23068 (N_23068,N_18930,N_19089);
or U23069 (N_23069,N_20859,N_18998);
nor U23070 (N_23070,N_18769,N_18460);
nand U23071 (N_23071,N_19387,N_18566);
and U23072 (N_23072,N_19911,N_18937);
and U23073 (N_23073,N_20651,N_19592);
nand U23074 (N_23074,N_20530,N_20897);
or U23075 (N_23075,N_20278,N_20743);
and U23076 (N_23076,N_18880,N_18977);
nand U23077 (N_23077,N_19493,N_20939);
nor U23078 (N_23078,N_20332,N_18450);
xnor U23079 (N_23079,N_20875,N_18449);
nand U23080 (N_23080,N_19529,N_18451);
nor U23081 (N_23081,N_19244,N_18976);
and U23082 (N_23082,N_19222,N_18358);
nor U23083 (N_23083,N_20297,N_18535);
nand U23084 (N_23084,N_20101,N_19130);
xor U23085 (N_23085,N_18627,N_19744);
nand U23086 (N_23086,N_20805,N_18939);
nor U23087 (N_23087,N_19281,N_18130);
or U23088 (N_23088,N_18839,N_18305);
nor U23089 (N_23089,N_18047,N_20524);
xnor U23090 (N_23090,N_20027,N_18984);
or U23091 (N_23091,N_18073,N_20151);
nand U23092 (N_23092,N_20151,N_19748);
or U23093 (N_23093,N_20961,N_19715);
nor U23094 (N_23094,N_20037,N_20169);
nor U23095 (N_23095,N_19352,N_18506);
nand U23096 (N_23096,N_18237,N_20677);
nor U23097 (N_23097,N_18612,N_18235);
nor U23098 (N_23098,N_20367,N_19525);
nor U23099 (N_23099,N_19585,N_18406);
nor U23100 (N_23100,N_19411,N_20716);
xnor U23101 (N_23101,N_18431,N_19103);
nand U23102 (N_23102,N_20630,N_18982);
nor U23103 (N_23103,N_20844,N_19659);
and U23104 (N_23104,N_20365,N_19935);
nand U23105 (N_23105,N_20666,N_18357);
nor U23106 (N_23106,N_18680,N_19831);
and U23107 (N_23107,N_20704,N_19591);
nand U23108 (N_23108,N_18711,N_19624);
or U23109 (N_23109,N_18334,N_18493);
nand U23110 (N_23110,N_19171,N_20208);
xor U23111 (N_23111,N_20259,N_20967);
and U23112 (N_23112,N_18489,N_18670);
nor U23113 (N_23113,N_19688,N_20876);
nand U23114 (N_23114,N_18616,N_20330);
and U23115 (N_23115,N_19425,N_19028);
xor U23116 (N_23116,N_18260,N_20154);
or U23117 (N_23117,N_19551,N_19141);
xor U23118 (N_23118,N_18020,N_19865);
or U23119 (N_23119,N_19629,N_20220);
nor U23120 (N_23120,N_19370,N_18893);
and U23121 (N_23121,N_20528,N_19075);
nor U23122 (N_23122,N_20306,N_18594);
xnor U23123 (N_23123,N_20452,N_18625);
nor U23124 (N_23124,N_18397,N_20100);
xnor U23125 (N_23125,N_18411,N_19187);
or U23126 (N_23126,N_18309,N_19832);
and U23127 (N_23127,N_19094,N_20929);
nor U23128 (N_23128,N_18067,N_20578);
nor U23129 (N_23129,N_18522,N_20444);
and U23130 (N_23130,N_18491,N_18718);
nor U23131 (N_23131,N_19761,N_20150);
and U23132 (N_23132,N_20374,N_18499);
nor U23133 (N_23133,N_18488,N_20597);
nand U23134 (N_23134,N_18102,N_19086);
xor U23135 (N_23135,N_20650,N_19591);
nor U23136 (N_23136,N_19022,N_19225);
and U23137 (N_23137,N_20812,N_20274);
nand U23138 (N_23138,N_19902,N_19099);
xor U23139 (N_23139,N_20354,N_19185);
and U23140 (N_23140,N_19400,N_19083);
or U23141 (N_23141,N_19193,N_19314);
nor U23142 (N_23142,N_20893,N_20054);
nand U23143 (N_23143,N_20226,N_19357);
and U23144 (N_23144,N_18725,N_18452);
nand U23145 (N_23145,N_18662,N_19724);
nor U23146 (N_23146,N_18487,N_19351);
nand U23147 (N_23147,N_19782,N_20273);
xor U23148 (N_23148,N_20687,N_18521);
or U23149 (N_23149,N_19352,N_20403);
nor U23150 (N_23150,N_19765,N_20882);
and U23151 (N_23151,N_20768,N_19317);
or U23152 (N_23152,N_18528,N_19972);
nand U23153 (N_23153,N_18559,N_20582);
or U23154 (N_23154,N_19113,N_18213);
xnor U23155 (N_23155,N_20639,N_18158);
or U23156 (N_23156,N_19001,N_19662);
nand U23157 (N_23157,N_19913,N_19370);
xnor U23158 (N_23158,N_19980,N_20780);
nand U23159 (N_23159,N_20454,N_18595);
xnor U23160 (N_23160,N_18527,N_20445);
xnor U23161 (N_23161,N_18601,N_19992);
and U23162 (N_23162,N_19432,N_19488);
nand U23163 (N_23163,N_18506,N_20176);
xor U23164 (N_23164,N_19696,N_18988);
xor U23165 (N_23165,N_19193,N_18183);
nor U23166 (N_23166,N_20096,N_20864);
nand U23167 (N_23167,N_20787,N_19150);
or U23168 (N_23168,N_18026,N_18692);
xnor U23169 (N_23169,N_19731,N_20087);
xnor U23170 (N_23170,N_19176,N_19918);
and U23171 (N_23171,N_18724,N_19980);
and U23172 (N_23172,N_19447,N_18757);
or U23173 (N_23173,N_19130,N_19315);
nor U23174 (N_23174,N_20805,N_19523);
xnor U23175 (N_23175,N_18800,N_18778);
xnor U23176 (N_23176,N_18460,N_18859);
or U23177 (N_23177,N_20114,N_19885);
or U23178 (N_23178,N_20007,N_20889);
nand U23179 (N_23179,N_19112,N_20392);
and U23180 (N_23180,N_18320,N_19774);
and U23181 (N_23181,N_20501,N_18410);
and U23182 (N_23182,N_19420,N_20456);
nor U23183 (N_23183,N_19532,N_18573);
nand U23184 (N_23184,N_20736,N_18991);
and U23185 (N_23185,N_20061,N_20227);
and U23186 (N_23186,N_18291,N_20827);
or U23187 (N_23187,N_19709,N_18016);
xnor U23188 (N_23188,N_20933,N_19415);
and U23189 (N_23189,N_18177,N_20084);
nor U23190 (N_23190,N_18231,N_18514);
or U23191 (N_23191,N_19986,N_19863);
or U23192 (N_23192,N_18975,N_18242);
nand U23193 (N_23193,N_18455,N_19559);
xor U23194 (N_23194,N_20424,N_19993);
nor U23195 (N_23195,N_18850,N_20433);
xor U23196 (N_23196,N_20418,N_20293);
nor U23197 (N_23197,N_18607,N_18518);
and U23198 (N_23198,N_19167,N_18421);
or U23199 (N_23199,N_19732,N_18050);
nor U23200 (N_23200,N_20484,N_19590);
nand U23201 (N_23201,N_18344,N_18234);
and U23202 (N_23202,N_18178,N_18360);
nand U23203 (N_23203,N_18577,N_20478);
or U23204 (N_23204,N_18984,N_18326);
xnor U23205 (N_23205,N_20760,N_18217);
and U23206 (N_23206,N_18486,N_19885);
nor U23207 (N_23207,N_20410,N_20057);
and U23208 (N_23208,N_18326,N_20949);
and U23209 (N_23209,N_20474,N_19233);
nand U23210 (N_23210,N_18357,N_20733);
nor U23211 (N_23211,N_19309,N_19197);
xnor U23212 (N_23212,N_18898,N_18560);
xnor U23213 (N_23213,N_20558,N_19904);
nand U23214 (N_23214,N_20249,N_18191);
xor U23215 (N_23215,N_20790,N_20619);
and U23216 (N_23216,N_20161,N_20367);
or U23217 (N_23217,N_20845,N_19021);
nor U23218 (N_23218,N_19557,N_19718);
nand U23219 (N_23219,N_18937,N_20363);
and U23220 (N_23220,N_20793,N_18616);
xor U23221 (N_23221,N_19030,N_18896);
xor U23222 (N_23222,N_20345,N_20915);
xnor U23223 (N_23223,N_18412,N_20540);
xor U23224 (N_23224,N_19423,N_18275);
xor U23225 (N_23225,N_18619,N_20834);
nand U23226 (N_23226,N_20364,N_19344);
xnor U23227 (N_23227,N_20309,N_19585);
xor U23228 (N_23228,N_18857,N_19224);
nand U23229 (N_23229,N_20700,N_20732);
nor U23230 (N_23230,N_19225,N_20992);
nand U23231 (N_23231,N_19089,N_20041);
nor U23232 (N_23232,N_19213,N_20424);
nand U23233 (N_23233,N_20220,N_18590);
xnor U23234 (N_23234,N_20946,N_18947);
nand U23235 (N_23235,N_18818,N_20887);
nand U23236 (N_23236,N_20089,N_18621);
and U23237 (N_23237,N_20839,N_20115);
or U23238 (N_23238,N_18782,N_18757);
and U23239 (N_23239,N_19644,N_19518);
and U23240 (N_23240,N_18983,N_18609);
and U23241 (N_23241,N_20567,N_19927);
or U23242 (N_23242,N_18228,N_19072);
nor U23243 (N_23243,N_18905,N_19553);
and U23244 (N_23244,N_18219,N_20459);
and U23245 (N_23245,N_18413,N_19046);
and U23246 (N_23246,N_18022,N_20364);
nand U23247 (N_23247,N_19961,N_20003);
nor U23248 (N_23248,N_20689,N_20963);
and U23249 (N_23249,N_19153,N_19999);
nor U23250 (N_23250,N_18284,N_20364);
or U23251 (N_23251,N_18719,N_18729);
xnor U23252 (N_23252,N_20642,N_19556);
xor U23253 (N_23253,N_20881,N_19779);
and U23254 (N_23254,N_18139,N_19948);
and U23255 (N_23255,N_20249,N_20538);
or U23256 (N_23256,N_18930,N_20924);
or U23257 (N_23257,N_19489,N_20384);
or U23258 (N_23258,N_19968,N_20691);
nor U23259 (N_23259,N_19043,N_20806);
nand U23260 (N_23260,N_19013,N_19214);
nor U23261 (N_23261,N_18451,N_20042);
or U23262 (N_23262,N_18071,N_19679);
and U23263 (N_23263,N_20228,N_18518);
and U23264 (N_23264,N_20324,N_19567);
xor U23265 (N_23265,N_18823,N_18984);
nand U23266 (N_23266,N_20857,N_19215);
nor U23267 (N_23267,N_18920,N_18461);
or U23268 (N_23268,N_19397,N_19952);
xor U23269 (N_23269,N_18060,N_19715);
xnor U23270 (N_23270,N_18205,N_19164);
xor U23271 (N_23271,N_18763,N_19164);
or U23272 (N_23272,N_19408,N_19997);
xor U23273 (N_23273,N_19806,N_20559);
xnor U23274 (N_23274,N_18194,N_20703);
xor U23275 (N_23275,N_19381,N_18276);
and U23276 (N_23276,N_18253,N_18222);
nand U23277 (N_23277,N_18302,N_18509);
and U23278 (N_23278,N_20858,N_20013);
or U23279 (N_23279,N_18395,N_19127);
nor U23280 (N_23280,N_19419,N_18284);
xor U23281 (N_23281,N_18296,N_19767);
and U23282 (N_23282,N_18940,N_20833);
nand U23283 (N_23283,N_19340,N_18226);
and U23284 (N_23284,N_18645,N_19849);
nand U23285 (N_23285,N_18246,N_18404);
or U23286 (N_23286,N_20387,N_20640);
or U23287 (N_23287,N_19318,N_19287);
nor U23288 (N_23288,N_18363,N_20665);
xor U23289 (N_23289,N_20455,N_20836);
nor U23290 (N_23290,N_18819,N_19690);
nor U23291 (N_23291,N_19612,N_18707);
nand U23292 (N_23292,N_19352,N_18070);
xor U23293 (N_23293,N_20139,N_19351);
nor U23294 (N_23294,N_20550,N_18970);
and U23295 (N_23295,N_19490,N_18828);
xnor U23296 (N_23296,N_18942,N_19703);
and U23297 (N_23297,N_19274,N_18625);
nor U23298 (N_23298,N_19136,N_19808);
xor U23299 (N_23299,N_20528,N_18635);
or U23300 (N_23300,N_18177,N_19072);
nand U23301 (N_23301,N_20023,N_20866);
xor U23302 (N_23302,N_19499,N_18456);
nor U23303 (N_23303,N_18201,N_18527);
and U23304 (N_23304,N_19880,N_19313);
xnor U23305 (N_23305,N_20742,N_20773);
nor U23306 (N_23306,N_19441,N_18053);
nor U23307 (N_23307,N_18587,N_20469);
xnor U23308 (N_23308,N_19977,N_19040);
or U23309 (N_23309,N_20870,N_19606);
nand U23310 (N_23310,N_19620,N_18663);
and U23311 (N_23311,N_19594,N_18904);
and U23312 (N_23312,N_18704,N_20467);
nor U23313 (N_23313,N_20195,N_18053);
xnor U23314 (N_23314,N_18422,N_19290);
xor U23315 (N_23315,N_18504,N_20711);
and U23316 (N_23316,N_18402,N_19192);
and U23317 (N_23317,N_19590,N_20105);
nand U23318 (N_23318,N_19659,N_20179);
nor U23319 (N_23319,N_20552,N_18943);
or U23320 (N_23320,N_20836,N_20198);
and U23321 (N_23321,N_18165,N_19950);
nand U23322 (N_23322,N_18546,N_20030);
nor U23323 (N_23323,N_20174,N_20506);
xor U23324 (N_23324,N_18815,N_19861);
or U23325 (N_23325,N_18569,N_18982);
xnor U23326 (N_23326,N_18702,N_19402);
nand U23327 (N_23327,N_18213,N_19749);
nor U23328 (N_23328,N_18615,N_19688);
and U23329 (N_23329,N_19360,N_20963);
and U23330 (N_23330,N_19659,N_19585);
nor U23331 (N_23331,N_18774,N_19891);
and U23332 (N_23332,N_19262,N_18128);
nand U23333 (N_23333,N_19537,N_19881);
nand U23334 (N_23334,N_20896,N_18464);
and U23335 (N_23335,N_19028,N_18354);
xor U23336 (N_23336,N_18850,N_20084);
and U23337 (N_23337,N_19952,N_19015);
xnor U23338 (N_23338,N_19368,N_19900);
nand U23339 (N_23339,N_18167,N_18956);
nand U23340 (N_23340,N_19455,N_18126);
xnor U23341 (N_23341,N_20876,N_19985);
xnor U23342 (N_23342,N_18371,N_19244);
and U23343 (N_23343,N_18363,N_19682);
nand U23344 (N_23344,N_19023,N_19221);
xor U23345 (N_23345,N_20767,N_20970);
nand U23346 (N_23346,N_18799,N_20306);
xor U23347 (N_23347,N_19124,N_18450);
nand U23348 (N_23348,N_20371,N_19337);
and U23349 (N_23349,N_20979,N_18575);
and U23350 (N_23350,N_19660,N_18353);
nor U23351 (N_23351,N_19219,N_19392);
and U23352 (N_23352,N_20565,N_19311);
or U23353 (N_23353,N_19206,N_20214);
nor U23354 (N_23354,N_18435,N_19358);
or U23355 (N_23355,N_18968,N_19052);
nand U23356 (N_23356,N_19809,N_18978);
nor U23357 (N_23357,N_20950,N_19424);
or U23358 (N_23358,N_18681,N_20745);
nand U23359 (N_23359,N_18154,N_18206);
and U23360 (N_23360,N_20713,N_20183);
and U23361 (N_23361,N_18123,N_19182);
nand U23362 (N_23362,N_18870,N_19583);
nand U23363 (N_23363,N_19054,N_19943);
nor U23364 (N_23364,N_19939,N_19210);
and U23365 (N_23365,N_20791,N_20177);
nor U23366 (N_23366,N_18719,N_19034);
nor U23367 (N_23367,N_18044,N_19948);
or U23368 (N_23368,N_20812,N_19204);
nand U23369 (N_23369,N_20785,N_20648);
or U23370 (N_23370,N_20855,N_19889);
or U23371 (N_23371,N_19872,N_19708);
or U23372 (N_23372,N_18779,N_19979);
and U23373 (N_23373,N_19317,N_19600);
and U23374 (N_23374,N_18651,N_18394);
nor U23375 (N_23375,N_19717,N_20702);
xor U23376 (N_23376,N_18615,N_19321);
nor U23377 (N_23377,N_20481,N_19930);
or U23378 (N_23378,N_19887,N_18652);
nand U23379 (N_23379,N_19233,N_20649);
nand U23380 (N_23380,N_18492,N_18122);
or U23381 (N_23381,N_20774,N_18451);
xnor U23382 (N_23382,N_18381,N_19572);
xnor U23383 (N_23383,N_19968,N_18812);
nand U23384 (N_23384,N_20491,N_19424);
nor U23385 (N_23385,N_19181,N_18580);
and U23386 (N_23386,N_19999,N_18308);
or U23387 (N_23387,N_19485,N_20448);
nand U23388 (N_23388,N_19608,N_20310);
or U23389 (N_23389,N_18719,N_18811);
nand U23390 (N_23390,N_18595,N_19755);
nand U23391 (N_23391,N_18679,N_20239);
nor U23392 (N_23392,N_20840,N_18205);
xor U23393 (N_23393,N_20680,N_19704);
or U23394 (N_23394,N_20826,N_19375);
or U23395 (N_23395,N_18824,N_18087);
or U23396 (N_23396,N_20358,N_19337);
xor U23397 (N_23397,N_18757,N_18854);
nand U23398 (N_23398,N_19927,N_19075);
or U23399 (N_23399,N_20634,N_18780);
and U23400 (N_23400,N_18367,N_18665);
or U23401 (N_23401,N_18306,N_20540);
and U23402 (N_23402,N_18321,N_20394);
nand U23403 (N_23403,N_20524,N_20815);
or U23404 (N_23404,N_18594,N_20900);
nand U23405 (N_23405,N_19560,N_19584);
xor U23406 (N_23406,N_20398,N_19399);
xor U23407 (N_23407,N_18781,N_18184);
or U23408 (N_23408,N_18624,N_18240);
and U23409 (N_23409,N_18830,N_18371);
and U23410 (N_23410,N_20579,N_20718);
and U23411 (N_23411,N_19457,N_20495);
xor U23412 (N_23412,N_18685,N_19907);
nor U23413 (N_23413,N_20826,N_18676);
nand U23414 (N_23414,N_20659,N_19089);
or U23415 (N_23415,N_19773,N_20147);
xnor U23416 (N_23416,N_20034,N_20512);
and U23417 (N_23417,N_20467,N_18625);
nor U23418 (N_23418,N_18307,N_18704);
xnor U23419 (N_23419,N_19811,N_19631);
nor U23420 (N_23420,N_20766,N_20569);
nor U23421 (N_23421,N_18240,N_18373);
xnor U23422 (N_23422,N_18003,N_18426);
and U23423 (N_23423,N_19242,N_18517);
or U23424 (N_23424,N_18867,N_19698);
and U23425 (N_23425,N_19980,N_20437);
nand U23426 (N_23426,N_20415,N_20590);
xnor U23427 (N_23427,N_18978,N_19463);
and U23428 (N_23428,N_20296,N_19881);
or U23429 (N_23429,N_20224,N_20471);
nand U23430 (N_23430,N_20363,N_18040);
and U23431 (N_23431,N_18665,N_18691);
or U23432 (N_23432,N_18307,N_20104);
or U23433 (N_23433,N_19976,N_20788);
or U23434 (N_23434,N_19540,N_18749);
nand U23435 (N_23435,N_19764,N_20678);
or U23436 (N_23436,N_19960,N_20356);
or U23437 (N_23437,N_20569,N_19165);
xnor U23438 (N_23438,N_19804,N_20200);
or U23439 (N_23439,N_19499,N_18103);
xnor U23440 (N_23440,N_20922,N_20327);
and U23441 (N_23441,N_18193,N_18071);
xor U23442 (N_23442,N_18528,N_19794);
nor U23443 (N_23443,N_20519,N_18822);
nand U23444 (N_23444,N_19713,N_19271);
or U23445 (N_23445,N_18346,N_20667);
and U23446 (N_23446,N_19759,N_19509);
nor U23447 (N_23447,N_18570,N_20531);
nor U23448 (N_23448,N_18451,N_19104);
nand U23449 (N_23449,N_18891,N_18058);
or U23450 (N_23450,N_19445,N_20960);
or U23451 (N_23451,N_18956,N_19126);
nor U23452 (N_23452,N_18246,N_18688);
and U23453 (N_23453,N_19821,N_19711);
xnor U23454 (N_23454,N_18676,N_18194);
or U23455 (N_23455,N_20429,N_19526);
nand U23456 (N_23456,N_19514,N_20514);
nand U23457 (N_23457,N_18392,N_18457);
nor U23458 (N_23458,N_18663,N_19726);
and U23459 (N_23459,N_20168,N_19752);
nand U23460 (N_23460,N_19202,N_20238);
nor U23461 (N_23461,N_18011,N_19535);
or U23462 (N_23462,N_18731,N_18284);
nand U23463 (N_23463,N_18657,N_20919);
nor U23464 (N_23464,N_19244,N_20246);
xnor U23465 (N_23465,N_19349,N_18912);
nand U23466 (N_23466,N_18578,N_19326);
xnor U23467 (N_23467,N_20138,N_20238);
or U23468 (N_23468,N_18987,N_18220);
xor U23469 (N_23469,N_20851,N_20297);
nand U23470 (N_23470,N_18508,N_18263);
xnor U23471 (N_23471,N_18889,N_19696);
and U23472 (N_23472,N_19322,N_18107);
or U23473 (N_23473,N_19693,N_20095);
nor U23474 (N_23474,N_18516,N_20428);
xor U23475 (N_23475,N_20494,N_19772);
nand U23476 (N_23476,N_20856,N_19469);
and U23477 (N_23477,N_19932,N_19923);
xor U23478 (N_23478,N_19941,N_18455);
nand U23479 (N_23479,N_19667,N_20655);
and U23480 (N_23480,N_20130,N_20604);
and U23481 (N_23481,N_20352,N_18177);
or U23482 (N_23482,N_19533,N_19704);
nor U23483 (N_23483,N_18360,N_18414);
xnor U23484 (N_23484,N_20374,N_20042);
or U23485 (N_23485,N_18916,N_18128);
xnor U23486 (N_23486,N_19496,N_19644);
nand U23487 (N_23487,N_20551,N_19978);
or U23488 (N_23488,N_18296,N_18636);
nor U23489 (N_23489,N_20152,N_20213);
xor U23490 (N_23490,N_18655,N_20055);
and U23491 (N_23491,N_19191,N_20612);
nand U23492 (N_23492,N_19526,N_18346);
xor U23493 (N_23493,N_20195,N_18803);
nor U23494 (N_23494,N_19846,N_19512);
xnor U23495 (N_23495,N_20399,N_20702);
xnor U23496 (N_23496,N_20882,N_18094);
xor U23497 (N_23497,N_18338,N_18105);
and U23498 (N_23498,N_18540,N_20018);
nand U23499 (N_23499,N_18703,N_18214);
xor U23500 (N_23500,N_18530,N_20596);
nor U23501 (N_23501,N_19507,N_20769);
or U23502 (N_23502,N_20582,N_18203);
or U23503 (N_23503,N_20980,N_20945);
nor U23504 (N_23504,N_18222,N_18433);
and U23505 (N_23505,N_20072,N_18146);
and U23506 (N_23506,N_19036,N_19150);
nor U23507 (N_23507,N_18648,N_19219);
or U23508 (N_23508,N_18123,N_20933);
xor U23509 (N_23509,N_19879,N_18999);
xor U23510 (N_23510,N_18808,N_20649);
nor U23511 (N_23511,N_19268,N_18474);
or U23512 (N_23512,N_18610,N_18903);
nor U23513 (N_23513,N_18577,N_18206);
and U23514 (N_23514,N_20393,N_20208);
xnor U23515 (N_23515,N_20815,N_20768);
nand U23516 (N_23516,N_19533,N_19420);
or U23517 (N_23517,N_19824,N_18040);
xor U23518 (N_23518,N_18082,N_18446);
nand U23519 (N_23519,N_19540,N_18487);
nor U23520 (N_23520,N_18712,N_19395);
and U23521 (N_23521,N_18484,N_18858);
nand U23522 (N_23522,N_20182,N_19548);
nor U23523 (N_23523,N_18479,N_18745);
and U23524 (N_23524,N_19201,N_20656);
nand U23525 (N_23525,N_18101,N_19237);
or U23526 (N_23526,N_19051,N_18448);
and U23527 (N_23527,N_20720,N_20864);
and U23528 (N_23528,N_20242,N_18841);
nand U23529 (N_23529,N_19733,N_19758);
or U23530 (N_23530,N_20736,N_19815);
nand U23531 (N_23531,N_18520,N_19098);
nand U23532 (N_23532,N_18328,N_19951);
nor U23533 (N_23533,N_18654,N_20367);
or U23534 (N_23534,N_19470,N_20369);
xor U23535 (N_23535,N_19132,N_20341);
or U23536 (N_23536,N_19355,N_18743);
nor U23537 (N_23537,N_19500,N_20066);
and U23538 (N_23538,N_20369,N_19861);
nand U23539 (N_23539,N_18103,N_19822);
and U23540 (N_23540,N_20976,N_19186);
nand U23541 (N_23541,N_18023,N_18404);
or U23542 (N_23542,N_20571,N_20082);
nand U23543 (N_23543,N_19648,N_18311);
nor U23544 (N_23544,N_19546,N_20537);
and U23545 (N_23545,N_18150,N_20579);
nor U23546 (N_23546,N_19635,N_19053);
nor U23547 (N_23547,N_18929,N_19315);
or U23548 (N_23548,N_20332,N_19925);
xnor U23549 (N_23549,N_18480,N_18000);
nor U23550 (N_23550,N_20297,N_20997);
or U23551 (N_23551,N_20664,N_18432);
and U23552 (N_23552,N_19734,N_18406);
xor U23553 (N_23553,N_19298,N_20348);
xor U23554 (N_23554,N_19948,N_18529);
or U23555 (N_23555,N_20586,N_18068);
nand U23556 (N_23556,N_18865,N_18369);
and U23557 (N_23557,N_20745,N_18773);
nand U23558 (N_23558,N_19645,N_18817);
nor U23559 (N_23559,N_19198,N_19108);
nor U23560 (N_23560,N_20801,N_20655);
xor U23561 (N_23561,N_19925,N_20095);
xor U23562 (N_23562,N_18081,N_20816);
xnor U23563 (N_23563,N_20369,N_18917);
nand U23564 (N_23564,N_18387,N_18011);
or U23565 (N_23565,N_18126,N_18538);
or U23566 (N_23566,N_18945,N_18517);
nor U23567 (N_23567,N_18611,N_19976);
xnor U23568 (N_23568,N_18581,N_20697);
or U23569 (N_23569,N_19896,N_18410);
nor U23570 (N_23570,N_18294,N_20561);
and U23571 (N_23571,N_18345,N_18093);
nand U23572 (N_23572,N_19321,N_19994);
nand U23573 (N_23573,N_18876,N_20532);
or U23574 (N_23574,N_20087,N_19084);
xor U23575 (N_23575,N_20933,N_18809);
and U23576 (N_23576,N_18425,N_20628);
nor U23577 (N_23577,N_18060,N_18691);
nand U23578 (N_23578,N_19418,N_18303);
or U23579 (N_23579,N_20445,N_20183);
or U23580 (N_23580,N_19405,N_19328);
nand U23581 (N_23581,N_18237,N_19130);
nor U23582 (N_23582,N_19256,N_20266);
or U23583 (N_23583,N_18661,N_19333);
xnor U23584 (N_23584,N_19022,N_19098);
nor U23585 (N_23585,N_20140,N_20057);
or U23586 (N_23586,N_20346,N_19547);
and U23587 (N_23587,N_19130,N_20568);
nand U23588 (N_23588,N_19147,N_18709);
and U23589 (N_23589,N_19466,N_19844);
nand U23590 (N_23590,N_18624,N_20291);
or U23591 (N_23591,N_18078,N_19656);
nor U23592 (N_23592,N_19756,N_20857);
nor U23593 (N_23593,N_20751,N_18006);
xor U23594 (N_23594,N_19483,N_18026);
nand U23595 (N_23595,N_20398,N_18407);
and U23596 (N_23596,N_18372,N_18258);
or U23597 (N_23597,N_20254,N_20842);
xnor U23598 (N_23598,N_19905,N_20930);
xnor U23599 (N_23599,N_18134,N_19391);
nand U23600 (N_23600,N_19789,N_18497);
nor U23601 (N_23601,N_18683,N_20185);
and U23602 (N_23602,N_18797,N_20195);
or U23603 (N_23603,N_20188,N_18222);
nor U23604 (N_23604,N_19375,N_19799);
nor U23605 (N_23605,N_20657,N_20428);
and U23606 (N_23606,N_20899,N_18649);
nand U23607 (N_23607,N_18676,N_18224);
nor U23608 (N_23608,N_18413,N_19914);
or U23609 (N_23609,N_19033,N_20649);
nor U23610 (N_23610,N_19141,N_20824);
nor U23611 (N_23611,N_18958,N_19209);
nand U23612 (N_23612,N_20966,N_19738);
nand U23613 (N_23613,N_19395,N_20461);
nand U23614 (N_23614,N_19212,N_20763);
or U23615 (N_23615,N_20398,N_18484);
nor U23616 (N_23616,N_19010,N_19502);
nor U23617 (N_23617,N_18077,N_18191);
nor U23618 (N_23618,N_20442,N_20831);
nand U23619 (N_23619,N_18516,N_20378);
nor U23620 (N_23620,N_18250,N_19001);
and U23621 (N_23621,N_20841,N_18876);
or U23622 (N_23622,N_19188,N_19098);
nand U23623 (N_23623,N_19123,N_18595);
or U23624 (N_23624,N_18854,N_18732);
nand U23625 (N_23625,N_20971,N_19085);
nand U23626 (N_23626,N_18488,N_18367);
nor U23627 (N_23627,N_20791,N_18336);
xnor U23628 (N_23628,N_19338,N_19007);
nand U23629 (N_23629,N_20288,N_20273);
or U23630 (N_23630,N_18007,N_19317);
nand U23631 (N_23631,N_20559,N_20416);
nand U23632 (N_23632,N_20180,N_20945);
nand U23633 (N_23633,N_18564,N_18481);
or U23634 (N_23634,N_20728,N_18892);
and U23635 (N_23635,N_18229,N_20930);
or U23636 (N_23636,N_20753,N_19511);
or U23637 (N_23637,N_19728,N_20544);
and U23638 (N_23638,N_19400,N_18090);
xnor U23639 (N_23639,N_20320,N_18643);
or U23640 (N_23640,N_20473,N_19317);
and U23641 (N_23641,N_18959,N_19210);
nor U23642 (N_23642,N_18891,N_18216);
nor U23643 (N_23643,N_18665,N_20333);
and U23644 (N_23644,N_18289,N_20374);
nand U23645 (N_23645,N_20873,N_18822);
and U23646 (N_23646,N_19836,N_18649);
xor U23647 (N_23647,N_20231,N_19702);
or U23648 (N_23648,N_19076,N_20432);
or U23649 (N_23649,N_20842,N_18110);
nand U23650 (N_23650,N_18340,N_20692);
or U23651 (N_23651,N_18013,N_18140);
nor U23652 (N_23652,N_19399,N_20857);
and U23653 (N_23653,N_19904,N_18573);
xnor U23654 (N_23654,N_19470,N_18225);
or U23655 (N_23655,N_19643,N_18723);
and U23656 (N_23656,N_19039,N_20884);
nor U23657 (N_23657,N_18163,N_18950);
or U23658 (N_23658,N_19377,N_19722);
xor U23659 (N_23659,N_18971,N_19693);
nor U23660 (N_23660,N_19592,N_19578);
nand U23661 (N_23661,N_19704,N_18082);
xor U23662 (N_23662,N_20808,N_19390);
nand U23663 (N_23663,N_19697,N_19510);
nand U23664 (N_23664,N_18634,N_20412);
nand U23665 (N_23665,N_20534,N_18173);
nand U23666 (N_23666,N_19614,N_19305);
or U23667 (N_23667,N_18028,N_20502);
nand U23668 (N_23668,N_19420,N_18384);
and U23669 (N_23669,N_19354,N_19400);
nand U23670 (N_23670,N_18165,N_19216);
and U23671 (N_23671,N_18910,N_20145);
and U23672 (N_23672,N_19087,N_18591);
nor U23673 (N_23673,N_20257,N_20273);
nor U23674 (N_23674,N_19367,N_19633);
nor U23675 (N_23675,N_18148,N_18177);
and U23676 (N_23676,N_20077,N_19789);
nand U23677 (N_23677,N_18929,N_18930);
or U23678 (N_23678,N_20889,N_19359);
nand U23679 (N_23679,N_19594,N_19785);
or U23680 (N_23680,N_19774,N_19056);
xor U23681 (N_23681,N_20637,N_20519);
nor U23682 (N_23682,N_19308,N_19388);
nor U23683 (N_23683,N_19205,N_20141);
and U23684 (N_23684,N_18924,N_18781);
nor U23685 (N_23685,N_19980,N_19154);
xor U23686 (N_23686,N_20693,N_19862);
and U23687 (N_23687,N_18372,N_18522);
and U23688 (N_23688,N_18203,N_18968);
nor U23689 (N_23689,N_19045,N_20087);
and U23690 (N_23690,N_20630,N_19420);
and U23691 (N_23691,N_18642,N_20503);
nor U23692 (N_23692,N_19661,N_18223);
or U23693 (N_23693,N_19358,N_20680);
and U23694 (N_23694,N_20986,N_18486);
and U23695 (N_23695,N_19304,N_18701);
or U23696 (N_23696,N_20433,N_19875);
and U23697 (N_23697,N_19891,N_19580);
xor U23698 (N_23698,N_20242,N_20154);
nor U23699 (N_23699,N_19316,N_19481);
nor U23700 (N_23700,N_18401,N_20846);
nor U23701 (N_23701,N_20929,N_19722);
nor U23702 (N_23702,N_18167,N_19908);
xnor U23703 (N_23703,N_18192,N_20027);
and U23704 (N_23704,N_20817,N_20858);
nand U23705 (N_23705,N_19692,N_18877);
and U23706 (N_23706,N_20910,N_20963);
xor U23707 (N_23707,N_18528,N_19764);
and U23708 (N_23708,N_18065,N_18225);
nor U23709 (N_23709,N_20856,N_18699);
xnor U23710 (N_23710,N_20385,N_19370);
nor U23711 (N_23711,N_18597,N_20098);
xor U23712 (N_23712,N_20525,N_18614);
nand U23713 (N_23713,N_18027,N_20287);
nor U23714 (N_23714,N_19428,N_18514);
and U23715 (N_23715,N_20924,N_19804);
or U23716 (N_23716,N_18179,N_18640);
and U23717 (N_23717,N_19851,N_20170);
and U23718 (N_23718,N_19258,N_19868);
nand U23719 (N_23719,N_19666,N_18653);
nand U23720 (N_23720,N_20549,N_20769);
and U23721 (N_23721,N_18027,N_18748);
nand U23722 (N_23722,N_18491,N_20669);
nand U23723 (N_23723,N_20044,N_18632);
and U23724 (N_23724,N_19238,N_18929);
nor U23725 (N_23725,N_20514,N_19836);
nor U23726 (N_23726,N_18870,N_20257);
nor U23727 (N_23727,N_18740,N_18961);
xnor U23728 (N_23728,N_18047,N_19881);
or U23729 (N_23729,N_20882,N_19477);
and U23730 (N_23730,N_20927,N_19583);
xnor U23731 (N_23731,N_20205,N_19259);
and U23732 (N_23732,N_18780,N_20766);
or U23733 (N_23733,N_18961,N_18812);
nor U23734 (N_23734,N_19177,N_18575);
nand U23735 (N_23735,N_18892,N_18507);
nor U23736 (N_23736,N_18672,N_19097);
nor U23737 (N_23737,N_19280,N_19947);
xor U23738 (N_23738,N_19360,N_18852);
nand U23739 (N_23739,N_20107,N_19234);
or U23740 (N_23740,N_20870,N_20467);
nor U23741 (N_23741,N_18235,N_19567);
or U23742 (N_23742,N_18801,N_19635);
and U23743 (N_23743,N_18477,N_18984);
nor U23744 (N_23744,N_20850,N_19836);
nand U23745 (N_23745,N_19968,N_20198);
nor U23746 (N_23746,N_20680,N_19376);
xor U23747 (N_23747,N_19645,N_20992);
and U23748 (N_23748,N_20033,N_19924);
xnor U23749 (N_23749,N_19857,N_20825);
and U23750 (N_23750,N_20417,N_19990);
nor U23751 (N_23751,N_20356,N_19635);
or U23752 (N_23752,N_19078,N_19783);
nor U23753 (N_23753,N_20042,N_19996);
xnor U23754 (N_23754,N_20729,N_20436);
xnor U23755 (N_23755,N_19271,N_20876);
nor U23756 (N_23756,N_18831,N_18235);
or U23757 (N_23757,N_19071,N_19885);
nand U23758 (N_23758,N_20384,N_19417);
and U23759 (N_23759,N_18138,N_20572);
nor U23760 (N_23760,N_18282,N_19924);
xnor U23761 (N_23761,N_19281,N_19421);
nor U23762 (N_23762,N_19296,N_20258);
xnor U23763 (N_23763,N_19612,N_18970);
nand U23764 (N_23764,N_20014,N_18218);
xor U23765 (N_23765,N_20156,N_19506);
and U23766 (N_23766,N_20958,N_19725);
xor U23767 (N_23767,N_19766,N_20701);
and U23768 (N_23768,N_18550,N_18011);
xor U23769 (N_23769,N_18398,N_19988);
nand U23770 (N_23770,N_20663,N_20168);
and U23771 (N_23771,N_20593,N_20112);
nor U23772 (N_23772,N_20483,N_20253);
and U23773 (N_23773,N_19803,N_18709);
and U23774 (N_23774,N_20992,N_19032);
and U23775 (N_23775,N_18351,N_19343);
or U23776 (N_23776,N_18814,N_19216);
nor U23777 (N_23777,N_19625,N_19675);
nand U23778 (N_23778,N_18492,N_19450);
or U23779 (N_23779,N_18571,N_19237);
or U23780 (N_23780,N_19119,N_20974);
xnor U23781 (N_23781,N_18588,N_20148);
and U23782 (N_23782,N_20184,N_19763);
nor U23783 (N_23783,N_18373,N_20047);
nor U23784 (N_23784,N_20278,N_19953);
nand U23785 (N_23785,N_19926,N_19151);
xor U23786 (N_23786,N_20081,N_18759);
nand U23787 (N_23787,N_18826,N_19251);
nand U23788 (N_23788,N_18440,N_18988);
and U23789 (N_23789,N_20350,N_20673);
nor U23790 (N_23790,N_18469,N_18621);
nand U23791 (N_23791,N_19363,N_20306);
nand U23792 (N_23792,N_18253,N_19476);
nand U23793 (N_23793,N_18251,N_19962);
and U23794 (N_23794,N_19140,N_19052);
nor U23795 (N_23795,N_18905,N_20991);
nor U23796 (N_23796,N_18807,N_20157);
nand U23797 (N_23797,N_19149,N_19768);
and U23798 (N_23798,N_18121,N_19799);
or U23799 (N_23799,N_18510,N_19996);
or U23800 (N_23800,N_19605,N_19400);
nor U23801 (N_23801,N_20212,N_19496);
nand U23802 (N_23802,N_20549,N_20309);
or U23803 (N_23803,N_18545,N_19847);
xnor U23804 (N_23804,N_19899,N_20735);
nor U23805 (N_23805,N_20165,N_19502);
or U23806 (N_23806,N_20659,N_20246);
nor U23807 (N_23807,N_19513,N_18874);
nor U23808 (N_23808,N_20507,N_20913);
nor U23809 (N_23809,N_18743,N_19635);
nor U23810 (N_23810,N_19266,N_19374);
and U23811 (N_23811,N_19485,N_19318);
or U23812 (N_23812,N_18985,N_18930);
and U23813 (N_23813,N_19727,N_19234);
nand U23814 (N_23814,N_20984,N_19553);
and U23815 (N_23815,N_20181,N_20826);
and U23816 (N_23816,N_19687,N_18024);
nand U23817 (N_23817,N_20510,N_19410);
and U23818 (N_23818,N_18612,N_20234);
xnor U23819 (N_23819,N_19112,N_20768);
nor U23820 (N_23820,N_19680,N_20264);
nor U23821 (N_23821,N_20409,N_19699);
or U23822 (N_23822,N_19138,N_18486);
and U23823 (N_23823,N_19006,N_19356);
xor U23824 (N_23824,N_18381,N_19667);
or U23825 (N_23825,N_18942,N_19615);
and U23826 (N_23826,N_20593,N_20838);
nand U23827 (N_23827,N_18361,N_20217);
nor U23828 (N_23828,N_18552,N_20007);
xnor U23829 (N_23829,N_18158,N_20939);
nor U23830 (N_23830,N_19918,N_20468);
or U23831 (N_23831,N_18966,N_19128);
nor U23832 (N_23832,N_20017,N_19589);
or U23833 (N_23833,N_19094,N_20403);
nor U23834 (N_23834,N_19511,N_20380);
or U23835 (N_23835,N_18942,N_18122);
nand U23836 (N_23836,N_19493,N_19783);
xnor U23837 (N_23837,N_20589,N_20567);
nand U23838 (N_23838,N_19664,N_20964);
nor U23839 (N_23839,N_20129,N_18630);
xor U23840 (N_23840,N_19630,N_20729);
or U23841 (N_23841,N_19350,N_18155);
or U23842 (N_23842,N_19222,N_18085);
nand U23843 (N_23843,N_20969,N_18274);
nand U23844 (N_23844,N_19837,N_19254);
nor U23845 (N_23845,N_20301,N_20807);
and U23846 (N_23846,N_20465,N_20705);
and U23847 (N_23847,N_19357,N_20799);
or U23848 (N_23848,N_20061,N_18062);
nor U23849 (N_23849,N_20286,N_20080);
or U23850 (N_23850,N_18264,N_19861);
xor U23851 (N_23851,N_19099,N_20096);
xor U23852 (N_23852,N_19757,N_19313);
or U23853 (N_23853,N_19213,N_18587);
and U23854 (N_23854,N_20070,N_20847);
or U23855 (N_23855,N_18165,N_18291);
and U23856 (N_23856,N_19771,N_18967);
or U23857 (N_23857,N_18685,N_20129);
nand U23858 (N_23858,N_20269,N_19542);
or U23859 (N_23859,N_20721,N_18786);
xnor U23860 (N_23860,N_18026,N_20590);
nor U23861 (N_23861,N_20237,N_18549);
and U23862 (N_23862,N_20871,N_19722);
nand U23863 (N_23863,N_18780,N_19212);
or U23864 (N_23864,N_20527,N_19205);
and U23865 (N_23865,N_20971,N_18548);
nor U23866 (N_23866,N_19979,N_18549);
xnor U23867 (N_23867,N_19619,N_18579);
nand U23868 (N_23868,N_19839,N_19783);
and U23869 (N_23869,N_18212,N_20728);
xnor U23870 (N_23870,N_20877,N_18683);
xor U23871 (N_23871,N_19014,N_20178);
nand U23872 (N_23872,N_20126,N_18656);
nor U23873 (N_23873,N_19233,N_19600);
nand U23874 (N_23874,N_18592,N_19641);
xnor U23875 (N_23875,N_19958,N_19670);
or U23876 (N_23876,N_20600,N_18082);
nand U23877 (N_23877,N_20076,N_18615);
and U23878 (N_23878,N_18489,N_20183);
nor U23879 (N_23879,N_19914,N_20515);
xnor U23880 (N_23880,N_18108,N_18146);
xor U23881 (N_23881,N_19732,N_18055);
nand U23882 (N_23882,N_19514,N_19661);
or U23883 (N_23883,N_20694,N_19784);
nand U23884 (N_23884,N_18410,N_20507);
or U23885 (N_23885,N_18107,N_20624);
xnor U23886 (N_23886,N_20064,N_19208);
and U23887 (N_23887,N_18951,N_18637);
or U23888 (N_23888,N_20854,N_18084);
nand U23889 (N_23889,N_18399,N_20447);
nor U23890 (N_23890,N_19217,N_18811);
nor U23891 (N_23891,N_19352,N_20161);
nor U23892 (N_23892,N_18170,N_20970);
xnor U23893 (N_23893,N_20964,N_20231);
or U23894 (N_23894,N_18546,N_19446);
and U23895 (N_23895,N_20216,N_19643);
xor U23896 (N_23896,N_19696,N_20165);
xnor U23897 (N_23897,N_20343,N_20089);
xor U23898 (N_23898,N_20004,N_18444);
nand U23899 (N_23899,N_20136,N_20929);
xor U23900 (N_23900,N_18952,N_20348);
xor U23901 (N_23901,N_19474,N_20704);
or U23902 (N_23902,N_20775,N_18230);
or U23903 (N_23903,N_18218,N_19374);
nor U23904 (N_23904,N_18073,N_18995);
nand U23905 (N_23905,N_19436,N_20234);
or U23906 (N_23906,N_18651,N_20196);
or U23907 (N_23907,N_19332,N_18665);
or U23908 (N_23908,N_20350,N_18922);
or U23909 (N_23909,N_20316,N_20243);
nand U23910 (N_23910,N_19000,N_19556);
nand U23911 (N_23911,N_19078,N_19205);
and U23912 (N_23912,N_19569,N_20101);
nor U23913 (N_23913,N_18805,N_20491);
or U23914 (N_23914,N_18206,N_20039);
and U23915 (N_23915,N_20942,N_18908);
nand U23916 (N_23916,N_20122,N_20950);
nor U23917 (N_23917,N_20449,N_19024);
and U23918 (N_23918,N_19197,N_19948);
and U23919 (N_23919,N_20613,N_19200);
xnor U23920 (N_23920,N_18801,N_18071);
nor U23921 (N_23921,N_18972,N_19633);
and U23922 (N_23922,N_20643,N_19794);
and U23923 (N_23923,N_19889,N_20989);
and U23924 (N_23924,N_19651,N_18810);
and U23925 (N_23925,N_18433,N_19219);
and U23926 (N_23926,N_20102,N_18994);
nand U23927 (N_23927,N_18963,N_18153);
nand U23928 (N_23928,N_20316,N_18984);
or U23929 (N_23929,N_20085,N_20707);
and U23930 (N_23930,N_20260,N_18852);
nor U23931 (N_23931,N_20826,N_20872);
or U23932 (N_23932,N_20937,N_19892);
or U23933 (N_23933,N_18719,N_19309);
xnor U23934 (N_23934,N_18827,N_20834);
or U23935 (N_23935,N_20306,N_20422);
nand U23936 (N_23936,N_18365,N_19903);
nor U23937 (N_23937,N_19959,N_20948);
nor U23938 (N_23938,N_18863,N_19906);
or U23939 (N_23939,N_20679,N_18071);
nand U23940 (N_23940,N_20898,N_20083);
nor U23941 (N_23941,N_18342,N_18468);
and U23942 (N_23942,N_19886,N_20466);
nand U23943 (N_23943,N_20054,N_18163);
xor U23944 (N_23944,N_20164,N_18591);
and U23945 (N_23945,N_18811,N_20296);
nand U23946 (N_23946,N_20181,N_20928);
nor U23947 (N_23947,N_18154,N_20680);
xor U23948 (N_23948,N_20502,N_19832);
and U23949 (N_23949,N_19977,N_18521);
and U23950 (N_23950,N_20023,N_19339);
xnor U23951 (N_23951,N_20502,N_18707);
nand U23952 (N_23952,N_20368,N_18123);
and U23953 (N_23953,N_20299,N_18378);
and U23954 (N_23954,N_20960,N_19097);
nand U23955 (N_23955,N_18375,N_20579);
nand U23956 (N_23956,N_20595,N_19897);
nand U23957 (N_23957,N_19457,N_20054);
and U23958 (N_23958,N_18764,N_20425);
xor U23959 (N_23959,N_18199,N_20864);
nor U23960 (N_23960,N_18409,N_20094);
xnor U23961 (N_23961,N_20254,N_19588);
or U23962 (N_23962,N_20240,N_19982);
and U23963 (N_23963,N_19334,N_20542);
xor U23964 (N_23964,N_18878,N_20187);
xor U23965 (N_23965,N_18880,N_19526);
xor U23966 (N_23966,N_19470,N_18036);
and U23967 (N_23967,N_19665,N_20075);
nor U23968 (N_23968,N_19164,N_19866);
xnor U23969 (N_23969,N_18306,N_20208);
and U23970 (N_23970,N_19913,N_18090);
nand U23971 (N_23971,N_18908,N_19020);
or U23972 (N_23972,N_19573,N_19902);
xnor U23973 (N_23973,N_19337,N_19767);
xnor U23974 (N_23974,N_19880,N_20941);
nand U23975 (N_23975,N_20424,N_19386);
xor U23976 (N_23976,N_19585,N_19917);
nor U23977 (N_23977,N_18663,N_20153);
nand U23978 (N_23978,N_18898,N_18446);
nor U23979 (N_23979,N_19644,N_19838);
nand U23980 (N_23980,N_19338,N_20121);
or U23981 (N_23981,N_20823,N_20356);
xnor U23982 (N_23982,N_20118,N_19835);
or U23983 (N_23983,N_20435,N_19697);
xor U23984 (N_23984,N_19056,N_18506);
nor U23985 (N_23985,N_18744,N_20433);
or U23986 (N_23986,N_19303,N_18191);
and U23987 (N_23987,N_18467,N_20988);
and U23988 (N_23988,N_20041,N_20928);
and U23989 (N_23989,N_18181,N_18416);
and U23990 (N_23990,N_18665,N_20128);
or U23991 (N_23991,N_20415,N_18972);
nand U23992 (N_23992,N_20004,N_19212);
or U23993 (N_23993,N_19834,N_19290);
and U23994 (N_23994,N_20655,N_18146);
or U23995 (N_23995,N_19816,N_20637);
xor U23996 (N_23996,N_18708,N_19802);
or U23997 (N_23997,N_18930,N_20519);
or U23998 (N_23998,N_18542,N_18343);
or U23999 (N_23999,N_20119,N_20152);
or U24000 (N_24000,N_22180,N_21944);
and U24001 (N_24001,N_22772,N_23013);
xnor U24002 (N_24002,N_21815,N_22474);
nor U24003 (N_24003,N_22659,N_23058);
nand U24004 (N_24004,N_23457,N_21332);
and U24005 (N_24005,N_23305,N_23880);
nor U24006 (N_24006,N_22977,N_22355);
nor U24007 (N_24007,N_23154,N_22909);
nor U24008 (N_24008,N_21164,N_23486);
nor U24009 (N_24009,N_22538,N_23766);
or U24010 (N_24010,N_21061,N_23502);
or U24011 (N_24011,N_21005,N_22848);
nand U24012 (N_24012,N_21328,N_22370);
xor U24013 (N_24013,N_23842,N_21729);
nor U24014 (N_24014,N_23854,N_21468);
or U24015 (N_24015,N_21206,N_21720);
or U24016 (N_24016,N_21900,N_21349);
xnor U24017 (N_24017,N_23315,N_22012);
or U24018 (N_24018,N_23840,N_21634);
and U24019 (N_24019,N_21963,N_22974);
nor U24020 (N_24020,N_23417,N_22630);
nor U24021 (N_24021,N_21416,N_22762);
and U24022 (N_24022,N_21135,N_22827);
and U24023 (N_24023,N_23487,N_21489);
or U24024 (N_24024,N_21772,N_22737);
or U24025 (N_24025,N_23292,N_23957);
nor U24026 (N_24026,N_21060,N_21214);
nand U24027 (N_24027,N_22542,N_21483);
nor U24028 (N_24028,N_22577,N_21934);
nor U24029 (N_24029,N_22555,N_23334);
or U24030 (N_24030,N_23931,N_23538);
nor U24031 (N_24031,N_21422,N_23145);
nand U24032 (N_24032,N_22479,N_22778);
and U24033 (N_24033,N_23994,N_22371);
and U24034 (N_24034,N_23375,N_22655);
or U24035 (N_24035,N_23934,N_23970);
or U24036 (N_24036,N_21566,N_23727);
or U24037 (N_24037,N_22065,N_21556);
or U24038 (N_24038,N_22249,N_23000);
xnor U24039 (N_24039,N_22080,N_23271);
or U24040 (N_24040,N_23675,N_22712);
nor U24041 (N_24041,N_21210,N_23998);
nand U24042 (N_24042,N_21993,N_23924);
nor U24043 (N_24043,N_23965,N_21001);
nor U24044 (N_24044,N_22450,N_21724);
nor U24045 (N_24045,N_23303,N_23193);
nand U24046 (N_24046,N_22026,N_23796);
nand U24047 (N_24047,N_21896,N_21192);
or U24048 (N_24048,N_21694,N_21590);
xor U24049 (N_24049,N_21335,N_23626);
xor U24050 (N_24050,N_23606,N_22968);
xnor U24051 (N_24051,N_22586,N_22616);
xor U24052 (N_24052,N_21317,N_22907);
nand U24053 (N_24053,N_21235,N_22412);
and U24054 (N_24054,N_21107,N_22821);
xnor U24055 (N_24055,N_22188,N_23878);
nand U24056 (N_24056,N_22162,N_21809);
nor U24057 (N_24057,N_23564,N_23231);
xor U24058 (N_24058,N_23191,N_22843);
nand U24059 (N_24059,N_23425,N_23782);
or U24060 (N_24060,N_23337,N_22683);
and U24061 (N_24061,N_23648,N_23990);
nand U24062 (N_24062,N_23577,N_21516);
nor U24063 (N_24063,N_22866,N_23959);
xnor U24064 (N_24064,N_22047,N_21254);
nor U24065 (N_24065,N_23379,N_22501);
and U24066 (N_24066,N_23644,N_23165);
nor U24067 (N_24067,N_22276,N_22265);
xor U24068 (N_24068,N_23918,N_23465);
or U24069 (N_24069,N_21293,N_22031);
and U24070 (N_24070,N_22987,N_23411);
xnor U24071 (N_24071,N_22918,N_22988);
or U24072 (N_24072,N_23049,N_23696);
nor U24073 (N_24073,N_22819,N_23055);
xor U24074 (N_24074,N_22956,N_22477);
and U24075 (N_24075,N_23911,N_21383);
xnor U24076 (N_24076,N_21817,N_23006);
nand U24077 (N_24077,N_22032,N_22131);
nand U24078 (N_24078,N_22269,N_21597);
xor U24079 (N_24079,N_21668,N_22947);
xnor U24080 (N_24080,N_22675,N_22602);
xnor U24081 (N_24081,N_23537,N_21904);
xor U24082 (N_24082,N_23557,N_23076);
xnor U24083 (N_24083,N_21946,N_21725);
and U24084 (N_24084,N_23177,N_22013);
nand U24085 (N_24085,N_23532,N_23304);
nor U24086 (N_24086,N_21956,N_21825);
nor U24087 (N_24087,N_21042,N_22944);
or U24088 (N_24088,N_23229,N_22802);
xor U24089 (N_24089,N_21831,N_23124);
nand U24090 (N_24090,N_23956,N_21881);
and U24091 (N_24091,N_23484,N_21111);
and U24092 (N_24092,N_21712,N_22615);
nor U24093 (N_24093,N_22279,N_22315);
and U24094 (N_24094,N_22749,N_23438);
xnor U24095 (N_24095,N_22658,N_22585);
xnor U24096 (N_24096,N_22543,N_23244);
nand U24097 (N_24097,N_21929,N_23674);
nor U24098 (N_24098,N_22251,N_21237);
nand U24099 (N_24099,N_21050,N_23901);
or U24100 (N_24100,N_21924,N_21666);
nor U24101 (N_24101,N_21909,N_23308);
or U24102 (N_24102,N_21802,N_22268);
nor U24103 (N_24103,N_23104,N_23655);
nand U24104 (N_24104,N_23961,N_22148);
xnor U24105 (N_24105,N_23389,N_22407);
xor U24106 (N_24106,N_21594,N_23364);
xnor U24107 (N_24107,N_23706,N_22088);
xnor U24108 (N_24108,N_21083,N_21721);
xnor U24109 (N_24109,N_21550,N_21770);
nand U24110 (N_24110,N_23159,N_23687);
or U24111 (N_24111,N_23640,N_23715);
or U24112 (N_24112,N_23050,N_21910);
xor U24113 (N_24113,N_22054,N_21188);
and U24114 (N_24114,N_21189,N_21346);
and U24115 (N_24115,N_22770,N_23637);
xnor U24116 (N_24116,N_21275,N_21264);
xor U24117 (N_24117,N_21620,N_22816);
or U24118 (N_24118,N_23102,N_21742);
nor U24119 (N_24119,N_23651,N_23386);
and U24120 (N_24120,N_23689,N_23157);
or U24121 (N_24121,N_22533,N_23171);
or U24122 (N_24122,N_23398,N_23097);
nor U24123 (N_24123,N_23784,N_22610);
nand U24124 (N_24124,N_22512,N_22916);
nor U24125 (N_24125,N_21600,N_23678);
xor U24126 (N_24126,N_21280,N_22900);
nor U24127 (N_24127,N_21120,N_22879);
and U24128 (N_24128,N_21090,N_21052);
xnor U24129 (N_24129,N_21173,N_21760);
or U24130 (N_24130,N_23493,N_21213);
nand U24131 (N_24131,N_23984,N_22614);
nand U24132 (N_24132,N_23581,N_23570);
nand U24133 (N_24133,N_21907,N_23716);
or U24134 (N_24134,N_22419,N_22536);
and U24135 (N_24135,N_21967,N_21466);
or U24136 (N_24136,N_22911,N_23643);
nand U24137 (N_24137,N_23295,N_22984);
and U24138 (N_24138,N_21057,N_22851);
xnor U24139 (N_24139,N_22862,N_21857);
nand U24140 (N_24140,N_21239,N_21696);
nor U24141 (N_24141,N_21244,N_21726);
nor U24142 (N_24142,N_23693,N_22068);
or U24143 (N_24143,N_21657,N_22850);
xor U24144 (N_24144,N_21064,N_21314);
nor U24145 (N_24145,N_21906,N_22449);
nand U24146 (N_24146,N_21345,N_21402);
xor U24147 (N_24147,N_21571,N_22203);
or U24148 (N_24148,N_21592,N_21059);
nor U24149 (N_24149,N_22828,N_22522);
nor U24150 (N_24150,N_23201,N_22183);
nor U24151 (N_24151,N_21846,N_23627);
xnor U24152 (N_24152,N_23933,N_21688);
nand U24153 (N_24153,N_23472,N_22334);
or U24154 (N_24154,N_23014,N_22651);
xor U24155 (N_24155,N_22596,N_21096);
nand U24156 (N_24156,N_22137,N_23714);
or U24157 (N_24157,N_23742,N_22669);
or U24158 (N_24158,N_22840,N_21800);
xnor U24159 (N_24159,N_23945,N_22353);
and U24160 (N_24160,N_22794,N_22223);
nand U24161 (N_24161,N_21948,N_21609);
nor U24162 (N_24162,N_21599,N_23819);
nor U24163 (N_24163,N_21893,N_21236);
or U24164 (N_24164,N_21957,N_22402);
and U24165 (N_24165,N_23483,N_22689);
or U24166 (N_24166,N_22405,N_21409);
nor U24167 (N_24167,N_21663,N_22073);
xnor U24168 (N_24168,N_23414,N_21397);
or U24169 (N_24169,N_21415,N_22566);
or U24170 (N_24170,N_21584,N_21326);
or U24171 (N_24171,N_21698,N_23153);
xnor U24172 (N_24172,N_23514,N_21185);
and U24173 (N_24173,N_22520,N_21912);
nor U24174 (N_24174,N_21358,N_23407);
nand U24175 (N_24175,N_21308,N_22923);
nor U24176 (N_24176,N_23041,N_22896);
nor U24177 (N_24177,N_21253,N_23515);
nand U24178 (N_24178,N_21020,N_21921);
nor U24179 (N_24179,N_23915,N_23089);
nor U24180 (N_24180,N_21341,N_23978);
or U24181 (N_24181,N_21552,N_21465);
nor U24182 (N_24182,N_22006,N_22375);
or U24183 (N_24183,N_22933,N_22225);
xor U24184 (N_24184,N_21865,N_22460);
and U24185 (N_24185,N_21676,N_22519);
xnor U24186 (N_24186,N_23353,N_23437);
xor U24187 (N_24187,N_22788,N_22789);
xnor U24188 (N_24188,N_21304,N_21361);
xnor U24189 (N_24189,N_22679,N_21453);
and U24190 (N_24190,N_21240,N_22835);
or U24191 (N_24191,N_22563,N_22343);
nor U24192 (N_24192,N_22677,N_22463);
and U24193 (N_24193,N_21227,N_23738);
xnor U24194 (N_24194,N_23078,N_22248);
or U24195 (N_24195,N_21311,N_23845);
and U24196 (N_24196,N_21582,N_23613);
or U24197 (N_24197,N_22965,N_22574);
nand U24198 (N_24198,N_21961,N_23694);
nand U24199 (N_24199,N_22832,N_22457);
xor U24200 (N_24200,N_21137,N_22886);
xnor U24201 (N_24201,N_22898,N_23061);
nor U24202 (N_24202,N_23241,N_23416);
or U24203 (N_24203,N_23633,N_21231);
nand U24204 (N_24204,N_21348,N_22147);
nor U24205 (N_24205,N_22901,N_23953);
nor U24206 (N_24206,N_22885,N_21419);
xnor U24207 (N_24207,N_23596,N_22880);
xor U24208 (N_24208,N_22876,N_23008);
xnor U24209 (N_24209,N_21932,N_22417);
xnor U24210 (N_24210,N_23068,N_21740);
and U24211 (N_24211,N_22786,N_22009);
nand U24212 (N_24212,N_23307,N_23833);
xnor U24213 (N_24213,N_21854,N_22409);
nor U24214 (N_24214,N_21834,N_23293);
and U24215 (N_24215,N_23419,N_21498);
nand U24216 (N_24216,N_21565,N_21751);
or U24217 (N_24217,N_22200,N_22143);
nand U24218 (N_24218,N_22261,N_22650);
nand U24219 (N_24219,N_23453,N_21216);
or U24220 (N_24220,N_22979,N_22314);
or U24221 (N_24221,N_22600,N_22090);
xnor U24222 (N_24222,N_23942,N_23677);
nor U24223 (N_24223,N_22608,N_23340);
or U24224 (N_24224,N_21215,N_22042);
nand U24225 (N_24225,N_21297,N_22513);
nor U24226 (N_24226,N_23958,N_22685);
and U24227 (N_24227,N_23296,N_21462);
or U24228 (N_24228,N_21132,N_22515);
or U24229 (N_24229,N_21719,N_22124);
xnor U24230 (N_24230,N_21505,N_23128);
and U24231 (N_24231,N_21562,N_21438);
or U24232 (N_24232,N_22497,N_22922);
nand U24233 (N_24233,N_23018,N_22485);
nor U24234 (N_24234,N_23310,N_23943);
xnor U24235 (N_24235,N_21257,N_21178);
nand U24236 (N_24236,N_22410,N_21521);
and U24237 (N_24237,N_21493,N_22550);
nand U24238 (N_24238,N_23332,N_21174);
or U24239 (N_24239,N_23559,N_22189);
and U24240 (N_24240,N_23974,N_22699);
and U24241 (N_24241,N_22633,N_23243);
nand U24242 (N_24242,N_23300,N_22861);
xor U24243 (N_24243,N_22713,N_21820);
or U24244 (N_24244,N_22233,N_22473);
and U24245 (N_24245,N_22528,N_22817);
and U24246 (N_24246,N_23800,N_21141);
xnor U24247 (N_24247,N_23807,N_23822);
and U24248 (N_24248,N_21618,N_22111);
nand U24249 (N_24249,N_21777,N_22403);
nor U24250 (N_24250,N_21350,N_22842);
and U24251 (N_24251,N_22038,N_23489);
xor U24252 (N_24252,N_23654,N_21169);
xnor U24253 (N_24253,N_22108,N_23922);
nand U24254 (N_24254,N_23075,N_22101);
and U24255 (N_24255,N_23753,N_21212);
nor U24256 (N_24256,N_22604,N_21097);
xnor U24257 (N_24257,N_23470,N_21014);
and U24258 (N_24258,N_21601,N_21832);
xor U24259 (N_24259,N_23544,N_21838);
nand U24260 (N_24260,N_22426,N_23764);
nand U24261 (N_24261,N_23370,N_22465);
nor U24262 (N_24262,N_22167,N_23125);
and U24263 (N_24263,N_23792,N_21593);
and U24264 (N_24264,N_22682,N_23259);
nor U24265 (N_24265,N_23030,N_22505);
nor U24266 (N_24266,N_22270,N_21794);
and U24267 (N_24267,N_22316,N_21852);
nand U24268 (N_24268,N_22197,N_21119);
or U24269 (N_24269,N_23447,N_21951);
or U24270 (N_24270,N_21261,N_23434);
or U24271 (N_24271,N_23762,N_21140);
xnor U24272 (N_24272,N_22171,N_23914);
and U24273 (N_24273,N_22389,N_21568);
nor U24274 (N_24274,N_22164,N_21327);
nor U24275 (N_24275,N_21177,N_23503);
and U24276 (N_24276,N_21378,N_21025);
nor U24277 (N_24277,N_21660,N_23598);
nor U24278 (N_24278,N_22396,N_23034);
or U24279 (N_24279,N_22741,N_21232);
or U24280 (N_24280,N_21970,N_22573);
xnor U24281 (N_24281,N_23712,N_21157);
nand U24282 (N_24282,N_21058,N_22572);
xnor U24283 (N_24283,N_23848,N_21673);
xor U24284 (N_24284,N_22309,N_22415);
nor U24285 (N_24285,N_21614,N_22684);
xnor U24286 (N_24286,N_22481,N_23939);
or U24287 (N_24287,N_22235,N_22652);
nand U24288 (N_24288,N_21445,N_21190);
nor U24289 (N_24289,N_23492,N_22982);
nor U24290 (N_24290,N_22387,N_23667);
and U24291 (N_24291,N_21977,N_23987);
xor U24292 (N_24292,N_23316,N_21204);
nor U24293 (N_24293,N_21197,N_23067);
nand U24294 (N_24294,N_23136,N_23299);
nor U24295 (N_24295,N_21360,N_21707);
nor U24296 (N_24296,N_21596,N_21766);
and U24297 (N_24297,N_23263,N_22349);
nand U24298 (N_24298,N_22322,N_22997);
nor U24299 (N_24299,N_21863,N_21022);
nand U24300 (N_24300,N_22062,N_22673);
or U24301 (N_24301,N_23117,N_23488);
and U24302 (N_24302,N_23586,N_23169);
nand U24303 (N_24303,N_23226,N_22765);
and U24304 (N_24304,N_22339,N_23402);
xor U24305 (N_24305,N_23383,N_22037);
nor U24306 (N_24306,N_22694,N_23906);
or U24307 (N_24307,N_21905,N_21155);
and U24308 (N_24308,N_21708,N_22480);
nand U24309 (N_24309,N_22932,N_22635);
nor U24310 (N_24310,N_23002,N_22333);
nand U24311 (N_24311,N_21091,N_23108);
nand U24312 (N_24312,N_22425,N_22284);
nor U24313 (N_24313,N_23812,N_22844);
and U24314 (N_24314,N_22022,N_22763);
xnor U24315 (N_24315,N_23988,N_23948);
nand U24316 (N_24316,N_22136,N_23035);
and U24317 (N_24317,N_22064,N_22970);
and U24318 (N_24318,N_23040,N_23755);
and U24319 (N_24319,N_21196,N_22191);
nand U24320 (N_24320,N_23856,N_23944);
xor U24321 (N_24321,N_21262,N_22045);
xor U24322 (N_24322,N_21911,N_23929);
nor U24323 (N_24323,N_22499,N_21381);
nand U24324 (N_24324,N_21558,N_21417);
and U24325 (N_24325,N_23350,N_21903);
nor U24326 (N_24326,N_23589,N_21675);
and U24327 (N_24327,N_21535,N_21495);
and U24328 (N_24328,N_21006,N_23883);
nor U24329 (N_24329,N_23342,N_21645);
nor U24330 (N_24330,N_21960,N_23546);
or U24331 (N_24331,N_21123,N_21723);
nand U24332 (N_24332,N_23042,N_22949);
xor U24333 (N_24333,N_23092,N_21291);
xor U24334 (N_24334,N_22920,N_21952);
nand U24335 (N_24335,N_22498,N_22422);
nor U24336 (N_24336,N_22967,N_21063);
and U24337 (N_24337,N_22895,N_22263);
or U24338 (N_24338,N_23384,N_23032);
nand U24339 (N_24339,N_23597,N_23960);
or U24340 (N_24340,N_21363,N_21610);
xnor U24341 (N_24341,N_23657,N_21224);
xor U24342 (N_24342,N_22447,N_21303);
or U24343 (N_24343,N_23257,N_21321);
nor U24344 (N_24344,N_22527,N_21843);
and U24345 (N_24345,N_23767,N_23232);
xor U24346 (N_24346,N_21106,N_22312);
xnor U24347 (N_24347,N_22039,N_22166);
xnor U24348 (N_24348,N_22307,N_21643);
nand U24349 (N_24349,N_22790,N_22808);
or U24350 (N_24350,N_23397,N_22989);
and U24351 (N_24351,N_21251,N_21969);
and U24352 (N_24352,N_22603,N_21194);
nor U24353 (N_24353,N_22751,N_21138);
or U24354 (N_24354,N_22597,N_23528);
nor U24355 (N_24355,N_23699,N_21773);
and U24356 (N_24356,N_23795,N_23190);
and U24357 (N_24357,N_22636,N_22133);
xnor U24358 (N_24358,N_22113,N_23963);
nand U24359 (N_24359,N_22648,N_23358);
xor U24360 (N_24360,N_23357,N_21856);
nand U24361 (N_24361,N_23695,N_21805);
and U24362 (N_24362,N_21671,N_23382);
xor U24363 (N_24363,N_22913,N_21522);
or U24364 (N_24364,N_23572,N_23641);
and U24365 (N_24365,N_21529,N_22362);
or U24366 (N_24366,N_22123,N_22461);
and U24367 (N_24367,N_21743,N_23571);
nand U24368 (N_24368,N_22390,N_23107);
xnor U24369 (N_24369,N_23155,N_23517);
and U24370 (N_24370,N_21472,N_23608);
and U24371 (N_24371,N_22381,N_21575);
xnor U24372 (N_24372,N_23940,N_22072);
nand U24373 (N_24373,N_22411,N_22357);
nor U24374 (N_24374,N_22545,N_21736);
nor U24375 (N_24375,N_23853,N_23805);
and U24376 (N_24376,N_21113,N_21756);
and U24377 (N_24377,N_21539,N_21233);
nor U24378 (N_24378,N_22548,N_23801);
xor U24379 (N_24379,N_22490,N_21441);
nor U24380 (N_24380,N_23343,N_23480);
nor U24381 (N_24381,N_22871,N_22187);
nand U24382 (N_24382,N_21109,N_23583);
nor U24383 (N_24383,N_21283,N_21023);
xor U24384 (N_24384,N_22019,N_21690);
and U24385 (N_24385,N_23832,N_21268);
xor U24386 (N_24386,N_22823,N_22326);
nor U24387 (N_24387,N_22116,N_21325);
and U24388 (N_24388,N_21356,N_22508);
and U24389 (N_24389,N_23967,N_23290);
xnor U24390 (N_24390,N_23843,N_23621);
nor U24391 (N_24391,N_23951,N_23007);
and U24392 (N_24392,N_21016,N_23786);
nand U24393 (N_24393,N_21249,N_22937);
or U24394 (N_24394,N_22611,N_23436);
and U24395 (N_24395,N_21950,N_21474);
and U24396 (N_24396,N_21744,N_21979);
or U24397 (N_24397,N_23509,N_22506);
and U24398 (N_24398,N_21928,N_23863);
and U24399 (N_24399,N_23279,N_23802);
and U24400 (N_24400,N_22331,N_22882);
and U24401 (N_24401,N_21890,N_22864);
nor U24402 (N_24402,N_22406,N_21036);
or U24403 (N_24403,N_22173,N_21028);
and U24404 (N_24404,N_21144,N_23427);
xnor U24405 (N_24405,N_22094,N_22190);
nand U24406 (N_24406,N_21876,N_23467);
or U24407 (N_24407,N_22742,N_23700);
nor U24408 (N_24408,N_22814,N_21983);
nand U24409 (N_24409,N_21242,N_22945);
and U24410 (N_24410,N_23200,N_23697);
nor U24411 (N_24411,N_21316,N_23276);
xor U24412 (N_24412,N_22126,N_21991);
nand U24413 (N_24413,N_22551,N_23870);
nand U24414 (N_24414,N_21718,N_21589);
nand U24415 (N_24415,N_23199,N_22239);
xnor U24416 (N_24416,N_22714,N_23806);
nor U24417 (N_24417,N_23661,N_23839);
or U24418 (N_24418,N_21450,N_23713);
nor U24419 (N_24419,N_23558,N_21633);
or U24420 (N_24420,N_23444,N_22238);
nor U24421 (N_24421,N_23935,N_21923);
xor U24422 (N_24422,N_23685,N_23829);
nor U24423 (N_24423,N_23979,N_23494);
xor U24424 (N_24424,N_21702,N_23019);
nand U24425 (N_24425,N_23827,N_21473);
or U24426 (N_24426,N_21201,N_21156);
and U24427 (N_24427,N_23745,N_23248);
nor U24428 (N_24428,N_23808,N_21373);
xnor U24429 (N_24429,N_21256,N_23680);
and U24430 (N_24430,N_23445,N_22360);
nor U24431 (N_24431,N_21246,N_21502);
nand U24432 (N_24432,N_23512,N_21027);
xnor U24433 (N_24433,N_21570,N_21585);
and U24434 (N_24434,N_23650,N_21658);
and U24435 (N_24435,N_22569,N_23875);
or U24436 (N_24436,N_22324,N_21258);
and U24437 (N_24437,N_21554,N_23036);
nor U24438 (N_24438,N_22277,N_23252);
xor U24439 (N_24439,N_21630,N_21999);
nand U24440 (N_24440,N_22386,N_23775);
nand U24441 (N_24441,N_21420,N_22975);
nand U24442 (N_24442,N_21376,N_23850);
nor U24443 (N_24443,N_21282,N_21228);
or U24444 (N_24444,N_23455,N_21300);
nor U24445 (N_24445,N_23964,N_21211);
nor U24446 (N_24446,N_21433,N_21414);
and U24447 (N_24447,N_21017,N_21377);
nor U24448 (N_24448,N_23575,N_22336);
nor U24449 (N_24449,N_21305,N_23099);
and U24450 (N_24450,N_23681,N_22385);
or U24451 (N_24451,N_22969,N_22549);
nor U24452 (N_24452,N_22732,N_21833);
and U24453 (N_24453,N_22983,N_23993);
nor U24454 (N_24454,N_22264,N_21333);
or U24455 (N_24455,N_21222,N_22283);
xnor U24456 (N_24456,N_23268,N_23098);
nand U24457 (N_24457,N_23356,N_23972);
and U24458 (N_24458,N_21919,N_21813);
nand U24459 (N_24459,N_21705,N_23253);
nand U24460 (N_24460,N_22016,N_23454);
nor U24461 (N_24461,N_21741,N_22745);
or U24462 (N_24462,N_23214,N_23496);
nand U24463 (N_24463,N_23485,N_22752);
nor U24464 (N_24464,N_21301,N_23463);
or U24465 (N_24465,N_23120,N_22467);
and U24466 (N_24466,N_22154,N_22274);
xnor U24467 (N_24467,N_22294,N_23505);
or U24468 (N_24468,N_23218,N_22592);
and U24469 (N_24469,N_23312,N_21292);
or U24470 (N_24470,N_23789,N_22060);
and U24471 (N_24471,N_22860,N_22210);
xor U24472 (N_24472,N_23614,N_21804);
nand U24473 (N_24473,N_23996,N_23701);
nor U24474 (N_24474,N_21738,N_22792);
nand U24475 (N_24475,N_22972,N_23410);
and U24476 (N_24476,N_21478,N_21176);
and U24477 (N_24477,N_23527,N_23717);
xor U24478 (N_24478,N_23146,N_22129);
and U24479 (N_24479,N_21623,N_22962);
nor U24480 (N_24480,N_23004,N_22346);
nor U24481 (N_24481,N_22423,N_23217);
xor U24482 (N_24482,N_23913,N_22328);
nor U24483 (N_24483,N_22489,N_22374);
nor U24484 (N_24484,N_21873,N_23834);
and U24485 (N_24485,N_23639,N_21713);
xnor U24486 (N_24486,N_23511,N_23448);
nand U24487 (N_24487,N_21886,N_21287);
nand U24488 (N_24488,N_23736,N_22622);
nand U24489 (N_24489,N_23429,N_23413);
or U24490 (N_24490,N_22342,N_23794);
or U24491 (N_24491,N_21093,N_21870);
and U24492 (N_24492,N_23404,N_21078);
nor U24493 (N_24493,N_23023,N_22856);
xnor U24494 (N_24494,N_21652,N_23652);
or U24495 (N_24495,N_21024,N_22537);
and U24496 (N_24496,N_21986,N_23287);
nor U24497 (N_24497,N_23743,N_23121);
xor U24498 (N_24498,N_22934,N_21267);
nor U24499 (N_24499,N_21576,N_23275);
or U24500 (N_24500,N_22702,N_21531);
and U24501 (N_24501,N_23844,N_21758);
or U24502 (N_24502,N_21342,N_21965);
or U24503 (N_24503,N_22395,N_23326);
xnor U24504 (N_24504,N_23301,N_21755);
xnor U24505 (N_24505,N_21868,N_21560);
xor U24506 (N_24506,N_21686,N_21647);
or U24507 (N_24507,N_21094,N_22579);
or U24508 (N_24508,N_23240,N_22291);
nor U24509 (N_24509,N_21079,N_23372);
xnor U24510 (N_24510,N_23450,N_21700);
nor U24511 (N_24511,N_21380,N_23531);
nor U24512 (N_24512,N_23520,N_21737);
nor U24513 (N_24513,N_23380,N_23314);
xnor U24514 (N_24514,N_21199,N_23524);
nor U24515 (N_24515,N_23424,N_21747);
nand U24516 (N_24516,N_21161,N_23874);
or U24517 (N_24517,N_23084,N_21954);
or U24518 (N_24518,N_23735,N_22767);
and U24519 (N_24519,N_23282,N_22416);
nand U24520 (N_24520,N_21761,N_21082);
nand U24521 (N_24521,N_22335,N_22785);
or U24522 (N_24522,N_23313,N_23066);
or U24523 (N_24523,N_22085,N_23751);
nand U24524 (N_24524,N_23223,N_22950);
nand U24525 (N_24525,N_21163,N_21980);
xnor U24526 (N_24526,N_22253,N_21801);
xor U24527 (N_24527,N_23368,N_22289);
xor U24528 (N_24528,N_21467,N_22259);
nand U24529 (N_24529,N_23896,N_21114);
xor U24530 (N_24530,N_23711,N_22155);
or U24531 (N_24531,N_22071,N_21278);
and U24532 (N_24532,N_23603,N_22948);
nand U24533 (N_24533,N_22867,N_21229);
or U24534 (N_24534,N_23950,N_21959);
nor U24535 (N_24535,N_21851,N_21208);
xnor U24536 (N_24536,N_21021,N_23879);
xor U24537 (N_24537,N_23975,N_21167);
or U24538 (N_24538,N_23325,N_23044);
nand U24539 (N_24539,N_22014,N_23973);
nor U24540 (N_24540,N_22858,N_23270);
nor U24541 (N_24541,N_23865,N_23065);
nor U24542 (N_24542,N_21624,N_22696);
or U24543 (N_24543,N_21730,N_22354);
and U24544 (N_24544,N_22966,N_21336);
or U24545 (N_24545,N_23861,N_23362);
xnor U24546 (N_24546,N_21627,N_22830);
and U24547 (N_24547,N_21835,N_23473);
and U24548 (N_24548,N_22942,N_23164);
nand U24549 (N_24549,N_21309,N_22340);
nor U24550 (N_24550,N_21115,N_23760);
or U24551 (N_24551,N_23665,N_22228);
xor U24552 (N_24552,N_21930,N_23636);
xnor U24553 (N_24553,N_21693,N_23899);
nand U24554 (N_24554,N_23012,N_23607);
or U24555 (N_24555,N_23726,N_23947);
nand U24556 (N_24556,N_22833,N_22906);
xor U24557 (N_24557,N_21644,N_22557);
xnor U24558 (N_24558,N_22161,N_21136);
xnor U24559 (N_24559,N_21538,N_23280);
xor U24560 (N_24560,N_21265,N_22626);
and U24561 (N_24561,N_22800,N_22372);
xor U24562 (N_24562,N_22925,N_21032);
and U24563 (N_24563,N_22888,N_22546);
nor U24564 (N_24564,N_23771,N_22178);
nand U24565 (N_24565,N_23284,N_22097);
or U24566 (N_24566,N_23811,N_21661);
and U24567 (N_24567,N_22981,N_21127);
nand U24568 (N_24568,N_22475,N_23818);
xor U24569 (N_24569,N_21653,N_22719);
or U24570 (N_24570,N_21112,N_22872);
nor U24571 (N_24571,N_22120,N_23617);
or U24572 (N_24572,N_23646,N_22275);
nand U24573 (N_24573,N_21260,N_21029);
nand U24574 (N_24574,N_22096,N_21049);
nand U24575 (N_24575,N_22282,N_22793);
nand U24576 (N_24576,N_23476,N_22991);
nand U24577 (N_24577,N_22653,N_22067);
xnor U24578 (N_24578,N_22027,N_23837);
or U24579 (N_24579,N_22380,N_21013);
nor U24580 (N_24580,N_23638,N_22055);
or U24581 (N_24581,N_23553,N_23590);
or U24582 (N_24582,N_23087,N_23803);
or U24583 (N_24583,N_23186,N_23148);
nor U24584 (N_24584,N_23867,N_23176);
and U24585 (N_24585,N_22773,N_23909);
nand U24586 (N_24586,N_21683,N_23756);
and U24587 (N_24587,N_22838,N_21966);
nor U24588 (N_24588,N_23926,N_22028);
or U24589 (N_24589,N_22236,N_21793);
nor U24590 (N_24590,N_22695,N_21774);
nor U24591 (N_24591,N_21824,N_23228);
nand U24592 (N_24592,N_22706,N_21818);
or U24593 (N_24593,N_23912,N_21147);
nand U24594 (N_24594,N_21862,N_22262);
nor U24595 (N_24595,N_23768,N_21494);
or U24596 (N_24596,N_22529,N_21089);
and U24597 (N_24597,N_22008,N_22996);
nand U24598 (N_24598,N_22358,N_21302);
or U24599 (N_24599,N_22050,N_22007);
nand U24600 (N_24600,N_22930,N_21323);
or U24601 (N_24601,N_23338,N_23195);
nand U24602 (N_24602,N_21563,N_22927);
xor U24603 (N_24603,N_22666,N_21551);
nand U24604 (N_24604,N_21754,N_21479);
xnor U24605 (N_24605,N_21710,N_23698);
or U24606 (N_24606,N_22383,N_21543);
nand U24607 (N_24607,N_22951,N_22365);
and U24608 (N_24608,N_21715,N_22992);
nand U24609 (N_24609,N_21913,N_22753);
nor U24610 (N_24610,N_21252,N_23855);
nor U24611 (N_24611,N_21180,N_22562);
and U24612 (N_24612,N_23890,N_23348);
xnor U24613 (N_24613,N_23123,N_23080);
nor U24614 (N_24614,N_23202,N_21860);
nand U24615 (N_24615,N_23734,N_21577);
nand U24616 (N_24616,N_23134,N_23359);
nand U24617 (N_24617,N_23816,N_21814);
nor U24618 (N_24618,N_21750,N_23298);
xnor U24619 (N_24619,N_22017,N_22735);
nor U24620 (N_24620,N_23908,N_23788);
nand U24621 (N_24621,N_23741,N_23830);
and U24622 (N_24622,N_21299,N_22320);
nand U24623 (N_24623,N_21674,N_21247);
nand U24624 (N_24624,N_21972,N_22290);
or U24625 (N_24625,N_22523,N_21126);
and U24626 (N_24626,N_22725,N_22280);
or U24627 (N_24627,N_22103,N_22672);
nand U24628 (N_24628,N_22338,N_23769);
and U24629 (N_24629,N_21488,N_21583);
and U24630 (N_24630,N_22069,N_23432);
and U24631 (N_24631,N_22717,N_23311);
or U24632 (N_24632,N_23462,N_23645);
nor U24633 (N_24633,N_23147,N_23053);
or U24634 (N_24634,N_22754,N_23302);
nand U24635 (N_24635,N_23401,N_21423);
nor U24636 (N_24636,N_22547,N_21612);
xor U24637 (N_24637,N_21035,N_23849);
nor U24638 (N_24638,N_23222,N_23037);
xor U24639 (N_24639,N_21307,N_22146);
nor U24640 (N_24640,N_22931,N_23746);
and U24641 (N_24641,N_21273,N_21476);
nand U24642 (N_24642,N_23221,N_21731);
nand U24643 (N_24643,N_22213,N_23921);
and U24644 (N_24644,N_23181,N_22980);
and U24645 (N_24645,N_23500,N_23668);
or U24646 (N_24646,N_22588,N_22158);
nor U24647 (N_24647,N_23601,N_21015);
and U24648 (N_24648,N_22217,N_22511);
xor U24649 (N_24649,N_22304,N_23459);
and U24650 (N_24650,N_22825,N_21128);
and U24651 (N_24651,N_23897,N_23872);
and U24652 (N_24652,N_21621,N_21399);
nand U24653 (N_24653,N_21679,N_21891);
or U24654 (N_24654,N_22718,N_21687);
and U24655 (N_24655,N_23090,N_21243);
and U24656 (N_24656,N_22722,N_23130);
xor U24657 (N_24657,N_23022,N_23043);
or U24658 (N_24658,N_21578,N_22791);
or U24659 (N_24659,N_23618,N_23466);
or U24660 (N_24660,N_21110,N_22746);
nor U24661 (N_24661,N_22516,N_22787);
nor U24662 (N_24662,N_22130,N_21352);
and U24663 (N_24663,N_21631,N_22105);
nor U24664 (N_24664,N_22676,N_21102);
nand U24665 (N_24665,N_21775,N_23167);
xor U24666 (N_24666,N_23916,N_22640);
xor U24667 (N_24667,N_22642,N_21389);
nor U24668 (N_24668,N_21520,N_22493);
nand U24669 (N_24669,N_21867,N_22119);
nand U24670 (N_24670,N_21672,N_23420);
nand U24671 (N_24671,N_21555,N_22526);
nand U24672 (N_24672,N_21709,N_23966);
nor U24673 (N_24673,N_21629,N_21532);
and U24674 (N_24674,N_23903,N_23156);
nand U24675 (N_24675,N_21162,N_21691);
xnor U24676 (N_24676,N_23750,N_23773);
and U24677 (N_24677,N_23622,N_23094);
nor U24678 (N_24678,N_22418,N_23374);
nor U24679 (N_24679,N_21711,N_22540);
and U24680 (N_24680,N_23220,N_22468);
xor U24681 (N_24681,N_21084,N_21369);
nor U24682 (N_24682,N_21528,N_22628);
nor U24683 (N_24683,N_21481,N_22311);
and U24684 (N_24684,N_23530,N_21622);
xor U24685 (N_24685,N_21628,N_22337);
nand U24686 (N_24686,N_21191,N_23027);
nor U24687 (N_24687,N_22869,N_23971);
nor U24688 (N_24688,N_23235,N_21685);
or U24689 (N_24689,N_23649,N_23482);
or U24690 (N_24690,N_21134,N_22492);
xor U24691 (N_24691,N_22114,N_21044);
nor U24692 (N_24692,N_21319,N_22205);
or U24693 (N_24693,N_21101,N_23518);
xor U24694 (N_24694,N_23905,N_23219);
xor U24695 (N_24695,N_21998,N_21048);
and U24696 (N_24696,N_23534,N_21008);
nand U24697 (N_24697,N_23250,N_22589);
nand U24698 (N_24698,N_23258,N_22029);
xnor U24699 (N_24699,N_23183,N_22344);
nor U24700 (N_24700,N_21418,N_22889);
xnor U24701 (N_24701,N_23451,N_21888);
xor U24702 (N_24702,N_22429,N_23692);
and U24703 (N_24703,N_22903,N_21706);
xnor U24704 (N_24704,N_22078,N_21037);
or U24705 (N_24705,N_22394,N_23452);
nor U24706 (N_24706,N_23900,N_23831);
nand U24707 (N_24707,N_22285,N_21461);
nor U24708 (N_24708,N_23980,N_22246);
nor U24709 (N_24709,N_22341,N_21810);
or U24710 (N_24710,N_21179,N_21812);
xor U24711 (N_24711,N_22472,N_21581);
or U24712 (N_24712,N_21393,N_21534);
nor U24713 (N_24713,N_21442,N_21816);
or U24714 (N_24714,N_22617,N_23992);
and U24715 (N_24715,N_23140,N_22744);
and U24716 (N_24716,N_22656,N_23024);
xnor U24717 (N_24717,N_22809,N_23281);
nand U24718 (N_24718,N_21330,N_21444);
nand U24719 (N_24719,N_23209,N_23112);
xor U24720 (N_24720,N_21981,N_21186);
xnor U24721 (N_24721,N_23765,N_23859);
nand U24722 (N_24722,N_23937,N_21000);
and U24723 (N_24723,N_21047,N_22194);
nand U24724 (N_24724,N_21051,N_22568);
nor U24725 (N_24725,N_22700,N_22297);
and U24726 (N_24726,N_21917,N_21763);
nand U24727 (N_24727,N_21103,N_22110);
and U24728 (N_24728,N_23776,N_23249);
nand U24729 (N_24729,N_23560,N_22641);
and U24730 (N_24730,N_21315,N_21382);
and U24731 (N_24731,N_23196,N_22567);
xnor U24732 (N_24732,N_23858,N_22952);
nand U24733 (N_24733,N_22193,N_23723);
or U24734 (N_24734,N_22446,N_21436);
and U24735 (N_24735,N_23498,N_22764);
nor U24736 (N_24736,N_23175,N_23391);
or U24737 (N_24737,N_22359,N_23331);
nor U24738 (N_24738,N_21785,N_22807);
and U24739 (N_24739,N_22897,N_21806);
xnor U24740 (N_24740,N_22075,N_23932);
xnor U24741 (N_24741,N_23101,N_22707);
nor U24742 (N_24742,N_21811,N_21054);
xnor U24743 (N_24743,N_21789,N_22728);
and U24744 (N_24744,N_22936,N_22040);
and U24745 (N_24745,N_21403,N_23917);
nand U24746 (N_24746,N_21281,N_22051);
xnor U24747 (N_24747,N_21682,N_23541);
xor U24748 (N_24748,N_21497,N_22929);
nor U24749 (N_24749,N_23260,N_23783);
nor U24750 (N_24750,N_21613,N_21411);
nand U24751 (N_24751,N_21739,N_21294);
nand U24752 (N_24752,N_23385,N_22820);
nor U24753 (N_24753,N_22919,N_21068);
or U24754 (N_24754,N_22414,N_23461);
or U24755 (N_24755,N_21787,N_21887);
xnor U24756 (N_24756,N_22935,N_21975);
nor U24757 (N_24757,N_22165,N_21276);
nor U24758 (N_24758,N_21407,N_22151);
nand U24759 (N_24759,N_23763,N_23272);
and U24760 (N_24760,N_22803,N_23860);
xor U24761 (N_24761,N_21649,N_22660);
nand U24762 (N_24762,N_22959,N_21408);
nand U24763 (N_24763,N_22591,N_22115);
nor U24764 (N_24764,N_22873,N_22605);
and U24765 (N_24765,N_21221,N_23441);
xor U24766 (N_24766,N_22716,N_23591);
or U24767 (N_24767,N_21394,N_22220);
and U24768 (N_24768,N_21648,N_21245);
or U24769 (N_24769,N_22964,N_21518);
xor U24770 (N_24770,N_23605,N_23083);
nand U24771 (N_24771,N_23611,N_22452);
xor U24772 (N_24772,N_23409,N_23045);
nor U24773 (N_24773,N_21121,N_22323);
nand U24774 (N_24774,N_22163,N_23095);
xor U24775 (N_24775,N_21153,N_22798);
nor U24776 (N_24776,N_23609,N_21219);
and U24777 (N_24777,N_23977,N_21455);
and U24778 (N_24778,N_22757,N_23739);
nor U24779 (N_24779,N_23469,N_23892);
nor U24780 (N_24780,N_23737,N_22680);
and U24781 (N_24781,N_22571,N_23519);
nand U24782 (N_24782,N_21588,N_21318);
nor U24783 (N_24783,N_23624,N_23203);
nand U24784 (N_24784,N_22521,N_22464);
nor U24785 (N_24785,N_21031,N_22145);
nor U24786 (N_24786,N_21925,N_21343);
nand U24787 (N_24787,N_22606,N_21486);
nand U24788 (N_24788,N_22993,N_21840);
nor U24789 (N_24789,N_23522,N_21655);
and U24790 (N_24790,N_23096,N_23852);
xor U24791 (N_24791,N_22905,N_23170);
nor U24792 (N_24792,N_23330,N_22525);
nand U24793 (N_24793,N_23406,N_23902);
nand U24794 (N_24794,N_21310,N_23390);
nand U24795 (N_24795,N_23399,N_22043);
xnor U24796 (N_24796,N_21768,N_21605);
nor U24797 (N_24797,N_21181,N_23205);
xnor U24798 (N_24798,N_21591,N_23785);
and U24799 (N_24799,N_22292,N_22688);
nand U24800 (N_24800,N_23632,N_21019);
xor U24801 (N_24801,N_21175,N_21171);
nand U24802 (N_24802,N_23659,N_21159);
xnor U24803 (N_24803,N_21749,N_21011);
xnor U24804 (N_24804,N_21874,N_21359);
nand U24805 (N_24805,N_23594,N_23187);
or U24806 (N_24806,N_22703,N_23017);
xor U24807 (N_24807,N_22318,N_23554);
nor U24808 (N_24808,N_22690,N_21065);
or U24809 (N_24809,N_21902,N_21734);
nand U24810 (N_24810,N_21365,N_22021);
or U24811 (N_24811,N_23592,N_22231);
nor U24812 (N_24812,N_22644,N_23690);
and U24813 (N_24813,N_23904,N_23192);
nand U24814 (N_24814,N_22859,N_22207);
and U24815 (N_24815,N_22963,N_22098);
xnor U24816 (N_24816,N_21372,N_22774);
or U24817 (N_24817,N_22025,N_22186);
or U24818 (N_24818,N_23110,N_22532);
nand U24819 (N_24819,N_23266,N_21198);
xor U24820 (N_24820,N_22091,N_21041);
nor U24821 (N_24821,N_23113,N_22795);
nand U24822 (N_24822,N_23930,N_21182);
or U24823 (N_24823,N_23625,N_22112);
xnor U24824 (N_24824,N_23568,N_21916);
xnor U24825 (N_24825,N_21861,N_21482);
nor U24826 (N_24826,N_22796,N_22229);
nand U24827 (N_24827,N_21586,N_22368);
nand U24828 (N_24828,N_23962,N_22976);
or U24829 (N_24829,N_23799,N_21490);
nor U24830 (N_24830,N_23684,N_21458);
and U24831 (N_24831,N_23732,N_23162);
xnor U24832 (N_24832,N_23551,N_22321);
xnor U24833 (N_24833,N_22215,N_21546);
xnor U24834 (N_24834,N_21125,N_21871);
nand U24835 (N_24835,N_23479,N_21574);
and U24836 (N_24836,N_21637,N_21512);
or U24837 (N_24837,N_22500,N_22582);
nand U24838 (N_24838,N_23683,N_22482);
nor U24839 (N_24839,N_22665,N_21650);
xnor U24840 (N_24840,N_23206,N_23804);
nor U24841 (N_24841,N_21943,N_22720);
nor U24842 (N_24842,N_22070,N_23671);
nor U24843 (N_24843,N_23576,N_21428);
nor U24844 (N_24844,N_22845,N_21547);
xor U24845 (N_24845,N_21602,N_21764);
nand U24846 (N_24846,N_21427,N_21003);
or U24847 (N_24847,N_21043,N_22564);
and U24848 (N_24848,N_21313,N_22201);
or U24849 (N_24849,N_21351,N_23319);
or U24850 (N_24850,N_22836,N_21839);
and U24851 (N_24851,N_22398,N_21259);
nand U24852 (N_24852,N_21587,N_22424);
and U24853 (N_24853,N_22863,N_21898);
xor U24854 (N_24854,N_22868,N_22724);
nor U24855 (N_24855,N_23122,N_22240);
nand U24856 (N_24856,N_21798,N_23197);
xor U24857 (N_24857,N_23133,N_23664);
nor U24858 (N_24858,N_21517,N_22288);
nand U24859 (N_24859,N_23707,N_22241);
xor U24860 (N_24860,N_22487,N_22232);
or U24861 (N_24861,N_23215,N_23082);
or U24862 (N_24862,N_21340,N_21945);
or U24863 (N_24863,N_21619,N_23277);
nand U24864 (N_24864,N_22899,N_21680);
and U24865 (N_24865,N_23919,N_23446);
nor U24866 (N_24866,N_21880,N_22781);
nor U24867 (N_24867,N_21329,N_21026);
nor U24868 (N_24868,N_22476,N_23744);
xnor U24869 (N_24869,N_23086,N_23274);
nand U24870 (N_24870,N_22444,N_22104);
or U24871 (N_24871,N_21279,N_21099);
and U24872 (N_24872,N_21200,N_23291);
nor U24873 (N_24873,N_21579,N_23660);
nor U24874 (N_24874,N_22364,N_23793);
and U24875 (N_24875,N_21974,N_22329);
nand U24876 (N_24876,N_23118,N_22199);
or U24877 (N_24877,N_21819,N_22295);
nor U24878 (N_24878,N_23225,N_23143);
nor U24879 (N_24879,N_22150,N_22704);
or U24880 (N_24880,N_21608,N_22804);
nor U24881 (N_24881,N_22607,N_23821);
or U24882 (N_24882,N_23373,N_22541);
and U24883 (N_24883,N_23610,N_21298);
or U24884 (N_24884,N_22462,N_23138);
or U24885 (N_24885,N_22243,N_21362);
and U24886 (N_24886,N_21218,N_23616);
nor U24887 (N_24887,N_23421,N_23048);
nand U24888 (N_24888,N_23920,N_23499);
nand U24889 (N_24889,N_23846,N_22442);
nand U24890 (N_24890,N_23207,N_21166);
nand U24891 (N_24891,N_21331,N_23369);
nor U24892 (N_24892,N_23072,N_22076);
xnor U24893 (N_24893,N_23779,N_22401);
or U24894 (N_24894,N_22544,N_22938);
and U24895 (N_24895,N_21073,N_22260);
nand U24896 (N_24896,N_21823,N_21053);
or U24897 (N_24897,N_23306,N_21781);
xnor U24898 (N_24898,N_23567,N_21938);
or U24899 (N_24899,N_22000,N_23388);
nor U24900 (N_24900,N_21782,N_21845);
nand U24901 (N_24901,N_22599,N_22247);
nor U24902 (N_24902,N_21540,N_21475);
or U24903 (N_24903,N_21496,N_22503);
and U24904 (N_24904,N_23393,N_22435);
and U24905 (N_24905,N_22459,N_21446);
and U24906 (N_24906,N_23910,N_22769);
nand U24907 (N_24907,N_21384,N_22961);
nor U24908 (N_24908,N_21988,N_22917);
nand U24909 (N_24909,N_21220,N_21987);
nor U24910 (N_24910,N_23976,N_23286);
xnor U24911 (N_24911,N_21745,N_21439);
or U24912 (N_24912,N_22756,N_23329);
or U24913 (N_24913,N_23543,N_23851);
nand U24914 (N_24914,N_23724,N_23995);
nor U24915 (N_24915,N_22049,N_23333);
xnor U24916 (N_24916,N_23267,N_21548);
nand U24917 (N_24917,N_21753,N_21425);
nor U24918 (N_24918,N_22160,N_21791);
nand U24919 (N_24919,N_22244,N_22400);
nand U24920 (N_24920,N_22504,N_22731);
nand U24921 (N_24921,N_22061,N_23893);
xnor U24922 (N_24922,N_23168,N_23825);
xor U24923 (N_24923,N_21447,N_21677);
nor U24924 (N_24924,N_23513,N_22747);
xnor U24925 (N_24925,N_23728,N_21487);
nand U24926 (N_24926,N_23208,N_21536);
and U24927 (N_24927,N_22729,N_23490);
nand U24928 (N_24928,N_21172,N_21697);
and U24929 (N_24929,N_22035,N_23814);
nor U24930 (N_24930,N_22377,N_21762);
and U24931 (N_24931,N_23781,N_22940);
or U24932 (N_24932,N_22875,N_23857);
or U24933 (N_24933,N_22625,N_23381);
nor U24934 (N_24934,N_22760,N_21296);
nor U24935 (N_24935,N_22293,N_22553);
xnor U24936 (N_24936,N_22030,N_23236);
nor U24937 (N_24937,N_23535,N_23230);
nand U24938 (N_24938,N_23415,N_23545);
or U24939 (N_24939,N_23059,N_21430);
nor U24940 (N_24940,N_22454,N_23378);
and U24941 (N_24941,N_21728,N_21238);
nand U24942 (N_24942,N_21841,N_22637);
xnor U24943 (N_24943,N_23439,N_22443);
nor U24944 (N_24944,N_23720,N_23163);
or U24945 (N_24945,N_22595,N_22388);
nand U24946 (N_24946,N_22083,N_21055);
xnor U24947 (N_24947,N_22583,N_21129);
or U24948 (N_24948,N_23265,N_23815);
nor U24949 (N_24949,N_23491,N_23820);
and U24950 (N_24950,N_23602,N_21116);
nor U24951 (N_24951,N_22530,N_23578);
or U24952 (N_24952,N_23536,N_21205);
xor U24953 (N_24953,N_21701,N_22033);
xnor U24954 (N_24954,N_22005,N_21337);
or U24955 (N_24955,N_22834,N_23841);
nand U24956 (N_24956,N_21285,N_22034);
nand U24957 (N_24957,N_22351,N_23709);
and U24958 (N_24958,N_23923,N_22420);
and U24959 (N_24959,N_23708,N_22855);
and U24960 (N_24960,N_21767,N_22384);
xnor U24961 (N_24961,N_22726,N_22518);
or U24962 (N_24962,N_22779,N_23579);
xnor U24963 (N_24963,N_23710,N_21778);
nor U24964 (N_24964,N_23881,N_21412);
and U24965 (N_24965,N_21410,N_22159);
or U24966 (N_24966,N_22978,N_22184);
xor U24967 (N_24967,N_22870,N_23351);
nand U24968 (N_24968,N_23888,N_23887);
nor U24969 (N_24969,N_22631,N_22638);
or U24970 (N_24970,N_22634,N_23345);
or U24971 (N_24971,N_23731,N_21885);
xnor U24972 (N_24972,N_23132,N_21312);
xnor U24973 (N_24973,N_22079,N_23623);
nand U24974 (N_24974,N_22681,N_22084);
nor U24975 (N_24975,N_22392,N_23216);
xnor U24976 (N_24976,N_21933,N_21746);
nor U24977 (N_24977,N_21398,N_23925);
or U24978 (N_24978,N_23021,N_22004);
and U24979 (N_24979,N_23179,N_21122);
or U24980 (N_24980,N_21792,N_22750);
xor U24981 (N_24981,N_22813,N_21821);
nand U24982 (N_24982,N_23748,N_23547);
or U24983 (N_24983,N_23497,N_23983);
xor U24984 (N_24984,N_21405,N_22258);
xnor U24985 (N_24985,N_23426,N_23777);
nand U24986 (N_24986,N_22001,N_21484);
nand U24987 (N_24987,N_21504,N_21150);
or U24988 (N_24988,N_22471,N_21388);
and U24989 (N_24989,N_21470,N_23422);
xnor U24990 (N_24990,N_21670,N_22924);
nand U24991 (N_24991,N_23288,N_21779);
xor U24992 (N_24992,N_22185,N_21828);
xor U24993 (N_24993,N_23327,N_23588);
xnor U24994 (N_24994,N_21580,N_23428);
nand U24995 (N_24995,N_23100,N_22327);
nand U24996 (N_24996,N_22587,N_22369);
and U24997 (N_24997,N_22620,N_21124);
nor U24998 (N_24998,N_23770,N_21836);
and U24999 (N_24999,N_21266,N_21374);
xor U25000 (N_25000,N_21632,N_23106);
or U25001 (N_25001,N_23985,N_21353);
nor U25002 (N_25002,N_21667,N_21776);
nor U25003 (N_25003,N_23733,N_23255);
nor U25004 (N_25004,N_23064,N_23721);
or U25005 (N_25005,N_22134,N_21636);
nand U25006 (N_25006,N_22739,N_21086);
nand U25007 (N_25007,N_23245,N_23079);
or U25008 (N_25008,N_23025,N_22439);
nor U25009 (N_25009,N_23982,N_21962);
and U25010 (N_25010,N_22325,N_22910);
nand U25011 (N_25011,N_23355,N_22960);
and U25012 (N_25012,N_23289,N_23349);
and U25013 (N_25013,N_22436,N_22469);
xnor U25014 (N_25014,N_21733,N_23239);
or U25015 (N_25015,N_21401,N_22887);
nor U25016 (N_25016,N_23435,N_22619);
nor U25017 (N_25017,N_23149,N_23224);
nor U25018 (N_25018,N_23456,N_22491);
nor U25019 (N_25019,N_21878,N_21914);
or U25020 (N_25020,N_22149,N_22252);
and U25021 (N_25021,N_22715,N_23178);
and U25022 (N_25022,N_21092,N_22382);
or U25023 (N_25023,N_23352,N_21822);
and U25024 (N_25024,N_21995,N_22748);
or U25025 (N_25025,N_23673,N_21844);
nor U25026 (N_25026,N_23449,N_21413);
and U25027 (N_25027,N_21390,N_22106);
xnor U25028 (N_25028,N_22663,N_21526);
nor U25029 (N_25029,N_23862,N_22488);
xnor U25030 (N_25030,N_22797,N_23180);
xor U25031 (N_25031,N_21651,N_22196);
nor U25032 (N_25032,N_21344,N_21976);
nor U25033 (N_25033,N_23403,N_23679);
and U25034 (N_25034,N_21872,N_23204);
or U25035 (N_25035,N_21477,N_23620);
xor U25036 (N_25036,N_23754,N_21030);
and U25037 (N_25037,N_21936,N_23151);
xnor U25038 (N_25038,N_21997,N_21424);
nor U25039 (N_25039,N_22273,N_23246);
xnor U25040 (N_25040,N_23184,N_21982);
or U25041 (N_25041,N_22723,N_21984);
nand U25042 (N_25042,N_22140,N_23261);
and U25043 (N_25043,N_23028,N_21146);
nand U25044 (N_25044,N_21664,N_21195);
and U25045 (N_25045,N_22534,N_21931);
and U25046 (N_25046,N_21148,N_22784);
nor U25047 (N_25047,N_22953,N_21463);
nand U25048 (N_25048,N_21525,N_21074);
or U25049 (N_25049,N_22456,N_22912);
or U25050 (N_25050,N_22234,N_22806);
nand U25051 (N_25051,N_21339,N_22531);
nand U25052 (N_25052,N_23869,N_21511);
xor U25053 (N_25053,N_21796,N_21783);
nand U25054 (N_25054,N_21371,N_21426);
or U25055 (N_25055,N_22507,N_22278);
and U25056 (N_25056,N_22811,N_23539);
xor U25057 (N_25057,N_22366,N_21607);
xor U25058 (N_25058,N_22198,N_22379);
or U25059 (N_25059,N_21567,N_23631);
and U25060 (N_25060,N_23105,N_22632);
nor U25061 (N_25061,N_21151,N_21527);
or U25062 (N_25062,N_21404,N_22755);
xnor U25063 (N_25063,N_22775,N_23936);
nor U25064 (N_25064,N_22121,N_22559);
or U25065 (N_25065,N_22727,N_21735);
xnor U25066 (N_25066,N_23057,N_21429);
or U25067 (N_25067,N_22670,N_22299);
or U25068 (N_25068,N_21347,N_21842);
xor U25069 (N_25069,N_23033,N_23894);
and U25070 (N_25070,N_21646,N_22003);
and U25071 (N_25071,N_23521,N_23468);
or U25072 (N_25072,N_23672,N_23269);
xor U25073 (N_25073,N_21072,N_21722);
xnor U25074 (N_25074,N_22928,N_21443);
or U25075 (N_25075,N_22561,N_21953);
or U25076 (N_25076,N_21149,N_22230);
and U25077 (N_25077,N_22393,N_22486);
or U25078 (N_25078,N_23772,N_23111);
or U25079 (N_25079,N_21850,N_21250);
or U25080 (N_25080,N_22440,N_22053);
xnor U25081 (N_25081,N_22074,N_22330);
xor U25082 (N_25082,N_22853,N_21320);
xor U25083 (N_25083,N_21454,N_23759);
xnor U25084 (N_25084,N_21662,N_21207);
xor U25085 (N_25085,N_21509,N_22570);
nor U25086 (N_25086,N_22086,N_21826);
nor U25087 (N_25087,N_21732,N_22458);
nor U25088 (N_25088,N_21448,N_23251);
nor U25089 (N_25089,N_22127,N_22857);
nand U25090 (N_25090,N_22759,N_21338);
or U25091 (N_25091,N_21184,N_22580);
or U25092 (N_25092,N_21431,N_23119);
and U25093 (N_25093,N_21449,N_21692);
and U25094 (N_25094,N_21139,N_21615);
or U25095 (N_25095,N_21748,N_22892);
xor U25096 (N_25096,N_21544,N_22046);
or U25097 (N_25097,N_22177,N_23172);
and U25098 (N_25098,N_22052,N_23320);
nand U25099 (N_25099,N_22308,N_22376);
or U25100 (N_25100,N_21075,N_22662);
or U25101 (N_25101,N_23991,N_23131);
and U25102 (N_25102,N_22301,N_23647);
or U25103 (N_25103,N_23341,N_23273);
and U25104 (N_25104,N_23876,N_23566);
and U25105 (N_25105,N_22300,N_22915);
nand U25106 (N_25106,N_23052,N_22302);
nand U25107 (N_25107,N_21513,N_23109);
nor U25108 (N_25108,N_23073,N_22224);
and U25109 (N_25109,N_21289,N_23871);
and U25110 (N_25110,N_21717,N_21598);
and U25111 (N_25111,N_22361,N_22609);
nand U25112 (N_25112,N_22138,N_22287);
nor U25113 (N_25113,N_22209,N_21456);
and U25114 (N_25114,N_21897,N_22466);
or U25115 (N_25115,N_23774,N_22846);
nor U25116 (N_25116,N_21949,N_21223);
xnor U25117 (N_25117,N_23365,N_21366);
or U25118 (N_25118,N_22643,N_22661);
or U25119 (N_25119,N_21654,N_21895);
nand U25120 (N_25120,N_23722,N_22831);
nor U25121 (N_25121,N_21866,N_22777);
nor U25122 (N_25122,N_23460,N_22733);
nor U25123 (N_25123,N_23443,N_22413);
and U25124 (N_25124,N_23628,N_23077);
nand U25125 (N_25125,N_23656,N_21611);
nand U25126 (N_25126,N_23582,N_23464);
xnor U25127 (N_25127,N_22350,N_23703);
and U25128 (N_25128,N_23242,N_21877);
nor U25129 (N_25129,N_23026,N_22266);
nor U25130 (N_25130,N_23091,N_23328);
and U25131 (N_25131,N_21117,N_22168);
nor U25132 (N_25132,N_21572,N_22226);
and U25133 (N_25133,N_23526,N_22157);
nor U25134 (N_25134,N_22494,N_21703);
and U25135 (N_25135,N_21545,N_21635);
xnor U25136 (N_25136,N_21780,N_21853);
and U25137 (N_25137,N_21869,N_22495);
xnor U25138 (N_25138,N_21131,N_22957);
nor U25139 (N_25139,N_21071,N_21922);
nand U25140 (N_25140,N_23020,N_23046);
nor U25141 (N_25141,N_21012,N_23635);
xor U25142 (N_25142,N_23471,N_21009);
nand U25143 (N_25143,N_21271,N_22122);
or U25144 (N_25144,N_23600,N_21421);
nand U25145 (N_25145,N_21606,N_21533);
nor U25146 (N_25146,N_23069,N_21187);
nand U25147 (N_25147,N_21209,N_23752);
or U25148 (N_25148,N_23321,N_21883);
xor U25149 (N_25149,N_23038,N_23477);
or U25150 (N_25150,N_21002,N_22738);
or U25151 (N_25151,N_23676,N_21143);
xnor U25152 (N_25152,N_22099,N_21480);
xnor U25153 (N_25153,N_23552,N_22908);
nor U25154 (N_25154,N_23166,N_23010);
or U25155 (N_25155,N_23981,N_23548);
xor U25156 (N_25156,N_22399,N_22448);
and U25157 (N_25157,N_21847,N_21056);
nor U25158 (N_25158,N_22883,N_23344);
nor U25159 (N_25159,N_21915,N_22227);
or U25160 (N_25160,N_22363,N_23550);
nor U25161 (N_25161,N_21395,N_21859);
nor U25162 (N_25162,N_22593,N_21018);
and U25163 (N_25163,N_22510,N_21158);
or U25164 (N_25164,N_21322,N_21908);
or U25165 (N_25165,N_23688,N_21152);
and U25166 (N_25166,N_21435,N_22613);
or U25167 (N_25167,N_21040,N_21656);
nand U25168 (N_25168,N_23740,N_23009);
xnor U25169 (N_25169,N_21973,N_23523);
nor U25170 (N_25170,N_23686,N_23630);
or U25171 (N_25171,N_23507,N_21226);
xor U25172 (N_25172,N_23824,N_21364);
nor U25173 (N_25173,N_23285,N_23440);
nand U25174 (N_25174,N_22010,N_22219);
or U25175 (N_25175,N_23895,N_21926);
or U25176 (N_25176,N_23160,N_21515);
or U25177 (N_25177,N_23927,N_21786);
nand U25178 (N_25178,N_21500,N_23070);
or U25179 (N_25179,N_22397,N_22576);
nand U25180 (N_25180,N_21769,N_21324);
or U25181 (N_25181,N_21894,N_21638);
nand U25182 (N_25182,N_22208,N_22601);
nor U25183 (N_25183,N_21968,N_21154);
xor U25184 (N_25184,N_22740,N_23144);
and U25185 (N_25185,N_22558,N_23847);
nor U25186 (N_25186,N_23946,N_23574);
nand U25187 (N_25187,N_23347,N_22771);
or U25188 (N_25188,N_21508,N_22878);
nor U25189 (N_25189,N_21641,N_22849);
and U25190 (N_25190,N_23563,N_21081);
xor U25191 (N_25191,N_22687,N_23394);
xnor U25192 (N_25192,N_21039,N_23584);
xor U25193 (N_25193,N_23371,N_22093);
and U25194 (N_25194,N_23873,N_22761);
or U25195 (N_25195,N_23780,N_23889);
and U25196 (N_25196,N_22847,N_23474);
and U25197 (N_25197,N_23001,N_21942);
or U25198 (N_25198,N_22678,N_22478);
nor U25199 (N_25199,N_22627,N_22671);
xnor U25200 (N_25200,N_22954,N_21994);
and U25201 (N_25201,N_21202,N_23658);
nor U25202 (N_25202,N_23081,N_22087);
or U25203 (N_25203,N_21375,N_23619);
and U25204 (N_25204,N_22594,N_21255);
nand U25205 (N_25205,N_21130,N_23324);
nor U25206 (N_25206,N_22175,N_21168);
xor U25207 (N_25207,N_22095,N_22250);
nand U25208 (N_25208,N_23555,N_22552);
and U25209 (N_25209,N_22884,N_22139);
nor U25210 (N_25210,N_21958,N_22192);
and U25211 (N_25211,N_21704,N_22144);
and U25212 (N_25212,N_23533,N_22995);
nand U25213 (N_25213,N_22701,N_21573);
or U25214 (N_25214,N_22955,N_23297);
nor U25215 (N_25215,N_22306,N_22657);
nor U25216 (N_25216,N_23396,N_21432);
xor U25217 (N_25217,N_23828,N_23256);
nor U25218 (N_25218,N_22310,N_22710);
xnor U25219 (N_25219,N_22170,N_22036);
or U25220 (N_25220,N_22612,N_23005);
nand U25221 (N_25221,N_21684,N_22092);
xor U25222 (N_25222,N_22204,N_23405);
or U25223 (N_25223,N_21370,N_22271);
or U25224 (N_25224,N_22812,N_23189);
nand U25225 (N_25225,N_23798,N_22810);
xnor U25226 (N_25226,N_23884,N_21807);
and U25227 (N_25227,N_22998,N_22891);
and U25228 (N_25228,N_21935,N_23354);
and U25229 (N_25229,N_23093,N_22893);
nand U25230 (N_25230,N_21080,N_23367);
nor U25231 (N_25231,N_21626,N_22082);
or U25232 (N_25232,N_23986,N_23247);
nand U25233 (N_25233,N_23254,N_22483);
xor U25234 (N_25234,N_22211,N_21459);
or U25235 (N_25235,N_21884,N_22286);
and U25236 (N_25236,N_22081,N_23211);
xor U25237 (N_25237,N_22865,N_23051);
nand U25238 (N_25238,N_22408,N_21971);
nand U25239 (N_25239,N_22169,N_21118);
or U25240 (N_25240,N_22839,N_22345);
or U25241 (N_25241,N_21989,N_23141);
nand U25242 (N_25242,N_23790,N_23999);
xnor U25243 (N_25243,N_23758,N_21665);
nand U25244 (N_25244,N_22218,N_21460);
xor U25245 (N_25245,N_23054,N_23088);
nor U25246 (N_25246,N_23823,N_22041);
and U25247 (N_25247,N_21457,N_23836);
or U25248 (N_25248,N_21659,N_21033);
and U25249 (N_25249,N_22222,N_21537);
and U25250 (N_25250,N_22216,N_21803);
nand U25251 (N_25251,N_23016,N_23283);
or U25252 (N_25252,N_21625,N_23761);
and U25253 (N_25253,N_22356,N_21990);
or U25254 (N_25254,N_23729,N_21387);
and U25255 (N_25255,N_22941,N_22697);
xnor U25256 (N_25256,N_22195,N_23126);
or U25257 (N_25257,N_23562,N_22142);
and U25258 (N_25258,N_21464,N_23137);
or U25259 (N_25259,N_21955,N_21062);
xnor U25260 (N_25260,N_23510,N_23949);
or U25261 (N_25261,N_22367,N_23294);
and U25262 (N_25262,N_21542,N_22667);
nand U25263 (N_25263,N_21165,N_21277);
and U25264 (N_25264,N_23114,N_21108);
and U25265 (N_25265,N_21485,N_22881);
or U25266 (N_25266,N_22135,N_22254);
or U25267 (N_25267,N_23565,N_22059);
xor U25268 (N_25268,N_23952,N_21530);
xnor U25269 (N_25269,N_21217,N_23718);
and U25270 (N_25270,N_23778,N_21788);
and U25271 (N_25271,N_21889,N_22066);
or U25272 (N_25272,N_22470,N_22431);
or U25273 (N_25273,N_21295,N_23481);
or U25274 (N_25274,N_21830,N_21145);
nand U25275 (N_25275,N_22373,N_22674);
and U25276 (N_25276,N_22581,N_21355);
xor U25277 (N_25277,N_22441,N_23395);
and U25278 (N_25278,N_23691,N_21104);
xnor U25279 (N_25279,N_21837,N_22214);
or U25280 (N_25280,N_21864,N_22958);
and U25281 (N_25281,N_22453,N_21765);
nor U25282 (N_25282,N_21992,N_23194);
and U25283 (N_25283,N_21503,N_21334);
nand U25284 (N_25284,N_21400,N_23882);
xnor U25285 (N_25285,N_21270,N_22890);
or U25286 (N_25286,N_21357,N_23540);
nand U25287 (N_25287,N_21392,N_21947);
or U25288 (N_25288,N_22780,N_23408);
xnor U25289 (N_25289,N_22645,N_22629);
nand U25290 (N_25290,N_23213,N_21985);
and U25291 (N_25291,N_22242,N_21379);
nand U25292 (N_25292,N_22939,N_22044);
or U25293 (N_25293,N_22433,N_21434);
or U25294 (N_25294,N_22852,N_23237);
nand U25295 (N_25295,N_22693,N_21437);
and U25296 (N_25296,N_21892,N_22826);
nand U25297 (N_25297,N_21286,N_21452);
nand U25298 (N_25298,N_23525,N_22646);
nor U25299 (N_25299,N_23360,N_22319);
and U25300 (N_25300,N_21561,N_21689);
nand U25301 (N_25301,N_22801,N_22023);
nand U25302 (N_25302,N_23115,N_23278);
and U25303 (N_25303,N_23504,N_22590);
xor U25304 (N_25304,N_23085,N_23423);
nor U25305 (N_25305,N_22624,N_23835);
nor U25306 (N_25306,N_21034,N_22109);
xor U25307 (N_25307,N_21604,N_21105);
or U25308 (N_25308,N_23392,N_21727);
or U25309 (N_25309,N_23886,N_21170);
nor U25310 (N_25310,N_23430,N_23318);
nand U25311 (N_25311,N_21098,N_23264);
xnor U25312 (N_25312,N_23063,N_22874);
or U25313 (N_25313,N_23478,N_23011);
and U25314 (N_25314,N_22783,N_23663);
or U25315 (N_25315,N_22709,N_21085);
and U25316 (N_25316,N_23135,N_22202);
nand U25317 (N_25317,N_23062,N_23725);
nor U25318 (N_25318,N_21193,N_22766);
nand U25319 (N_25319,N_21784,N_22181);
and U25320 (N_25320,N_22221,N_23029);
and U25321 (N_25321,N_22445,N_23182);
xnor U25322 (N_25322,N_22427,N_22539);
nand U25323 (N_25323,N_21541,N_23682);
nor U25324 (N_25324,N_22206,N_22584);
nand U25325 (N_25325,N_23615,N_23662);
nor U25326 (N_25326,N_21368,N_23704);
and U25327 (N_25327,N_22815,N_23653);
xnor U25328 (N_25328,N_22654,N_21920);
and U25329 (N_25329,N_22313,N_23074);
nand U25330 (N_25330,N_23139,N_22172);
nand U25331 (N_25331,N_22296,N_22305);
nand U25332 (N_25332,N_22999,N_23549);
nor U25333 (N_25333,N_21603,N_21385);
nor U25334 (N_25334,N_23864,N_21849);
nand U25335 (N_25335,N_23047,N_21901);
nand U25336 (N_25336,N_22132,N_21183);
nor U25337 (N_25337,N_23387,N_22179);
and U25338 (N_25338,N_21406,N_22768);
nand U25339 (N_25339,N_22267,N_22298);
and U25340 (N_25340,N_21284,N_23400);
nor U25341 (N_25341,N_23666,N_23938);
xnor U25342 (N_25342,N_23366,N_22743);
nand U25343 (N_25343,N_21510,N_23928);
nor U25344 (N_25344,N_22514,N_23442);
or U25345 (N_25345,N_21681,N_22272);
nor U25346 (N_25346,N_22818,N_23898);
or U25347 (N_25347,N_22332,N_21699);
xor U25348 (N_25348,N_21076,N_21095);
or U25349 (N_25349,N_22575,N_23826);
nand U25350 (N_25350,N_23198,N_21501);
xor U25351 (N_25351,N_22058,N_22484);
nand U25352 (N_25352,N_22902,N_22437);
and U25353 (N_25353,N_21272,N_22565);
or U25354 (N_25354,N_21918,N_21616);
nor U25355 (N_25355,N_21549,N_23317);
nor U25356 (N_25356,N_22141,N_23031);
xor U25357 (N_25357,N_22926,N_21492);
nand U25358 (N_25358,N_21288,N_21499);
xnor U25359 (N_25359,N_22317,N_21506);
nand U25360 (N_25360,N_23969,N_22782);
and U25361 (N_25361,N_23749,N_22107);
and U25362 (N_25362,N_23604,N_21640);
nor U25363 (N_25363,N_23702,N_21595);
nor U25364 (N_25364,N_21882,N_22153);
xor U25365 (N_25365,N_22020,N_22535);
nand U25366 (N_25366,N_23056,N_21996);
nor U25367 (N_25367,N_21386,N_21491);
nor U25368 (N_25368,N_23506,N_22117);
and U25369 (N_25369,N_23941,N_21524);
nand U25370 (N_25370,N_23495,N_21927);
xnor U25371 (N_25371,N_23877,N_21642);
nand U25372 (N_25372,N_23907,N_21440);
xnor U25373 (N_25373,N_23599,N_22647);
xor U25374 (N_25374,N_23116,N_21160);
xor U25375 (N_25375,N_23634,N_22623);
nor U25376 (N_25376,N_23152,N_21939);
or U25377 (N_25377,N_23015,N_23561);
nand U25378 (N_25378,N_21087,N_21274);
nor U25379 (N_25379,N_23127,N_21354);
nand U25380 (N_25380,N_22102,N_22002);
nor U25381 (N_25381,N_21617,N_23791);
nand U25382 (N_25382,N_21046,N_21230);
or U25383 (N_25383,N_21678,N_21759);
and U25384 (N_25384,N_21451,N_22509);
nor U25385 (N_25385,N_22245,N_21069);
nand U25386 (N_25386,N_23705,N_22455);
and U25387 (N_25387,N_22303,N_23868);
nor U25388 (N_25388,N_21203,N_21557);
and U25389 (N_25389,N_21225,N_21553);
nor U25390 (N_25390,N_23377,N_22255);
and U25391 (N_25391,N_21559,N_23585);
nand U25392 (N_25392,N_21142,N_23508);
or U25393 (N_25393,N_22237,N_23757);
xor U25394 (N_25394,N_23339,N_23809);
or U25395 (N_25395,N_23669,N_22943);
and U25396 (N_25396,N_22281,N_21066);
or U25397 (N_25397,N_22822,N_21855);
and U25398 (N_25398,N_22618,N_23501);
nand U25399 (N_25399,N_21306,N_23212);
nand U25400 (N_25400,N_23573,N_22156);
nand U25401 (N_25401,N_23580,N_21771);
and U25402 (N_25402,N_21808,N_23150);
nor U25403 (N_25403,N_22011,N_22496);
xor U25404 (N_25404,N_23629,N_22971);
nor U25405 (N_25405,N_21070,N_23719);
and U25406 (N_25406,N_22877,N_22799);
nor U25407 (N_25407,N_21716,N_22352);
and U25408 (N_25408,N_22705,N_22421);
and U25409 (N_25409,N_21899,N_23817);
nand U25410 (N_25410,N_21010,N_22736);
xor U25411 (N_25411,N_23516,N_22946);
and U25412 (N_25412,N_22994,N_21858);
nor U25413 (N_25413,N_21100,N_23233);
and U25414 (N_25414,N_21757,N_22824);
or U25415 (N_25415,N_23968,N_21507);
nand U25416 (N_25416,N_21827,N_21290);
or U25417 (N_25417,N_22554,N_21519);
nand U25418 (N_25418,N_21875,N_21523);
and U25419 (N_25419,N_22434,N_21241);
xor U25420 (N_25420,N_22089,N_22118);
and U25421 (N_25421,N_23747,N_22432);
xor U25422 (N_25422,N_22174,N_22057);
nand U25423 (N_25423,N_23787,N_22560);
or U25424 (N_25424,N_21941,N_23997);
nor U25425 (N_25425,N_22015,N_22664);
xor U25426 (N_25426,N_23458,N_22598);
nand U25427 (N_25427,N_22711,N_22698);
nor U25428 (N_25428,N_23003,N_22152);
nand U25429 (N_25429,N_21269,N_21940);
nor U25430 (N_25430,N_23039,N_21077);
and U25431 (N_25431,N_23569,N_21067);
nand U25432 (N_25432,N_23309,N_23361);
nand U25433 (N_25433,N_23529,N_22128);
nand U25434 (N_25434,N_21004,N_22024);
xor U25435 (N_25435,N_23431,N_22708);
nand U25436 (N_25436,N_22430,N_22100);
and U25437 (N_25437,N_23323,N_23174);
or U25438 (N_25438,N_22973,N_21007);
and U25439 (N_25439,N_23262,N_22805);
or U25440 (N_25440,N_22056,N_21088);
nor U25441 (N_25441,N_22212,N_23238);
or U25442 (N_25442,N_22894,N_23363);
xor U25443 (N_25443,N_23813,N_21879);
and U25444 (N_25444,N_23838,N_22986);
nor U25445 (N_25445,N_21639,N_22776);
or U25446 (N_25446,N_22348,N_21799);
xnor U25447 (N_25447,N_21829,N_23234);
and U25448 (N_25448,N_23542,N_21038);
or U25449 (N_25449,N_23161,N_23587);
xor U25450 (N_25450,N_23060,N_22985);
or U25451 (N_25451,N_22692,N_22758);
nand U25452 (N_25452,N_22649,N_23954);
xor U25453 (N_25453,N_22517,N_21564);
nand U25454 (N_25454,N_21937,N_22829);
and U25455 (N_25455,N_22721,N_21795);
and U25456 (N_25456,N_22428,N_21752);
and U25457 (N_25457,N_22904,N_22347);
or U25458 (N_25458,N_22257,N_23955);
and U25459 (N_25459,N_23185,N_23989);
xnor U25460 (N_25460,N_22018,N_22691);
xor U25461 (N_25461,N_21978,N_23593);
nor U25462 (N_25462,N_22077,N_23335);
nand U25463 (N_25463,N_22451,N_23642);
or U25464 (N_25464,N_22176,N_21391);
nand U25465 (N_25465,N_23891,N_22621);
and U25466 (N_25466,N_22837,N_21714);
xor U25467 (N_25467,N_22502,N_23142);
or U25468 (N_25468,N_23556,N_22914);
xor U25469 (N_25469,N_22730,N_23885);
or U25470 (N_25470,N_21133,N_23188);
nor U25471 (N_25471,N_21695,N_23412);
and U25472 (N_25472,N_22841,N_21263);
and U25473 (N_25473,N_23475,N_21471);
xnor U25474 (N_25474,N_22404,N_22854);
xor U25475 (N_25475,N_22921,N_22556);
or U25476 (N_25476,N_21790,N_22639);
nor U25477 (N_25477,N_21669,N_22686);
nor U25478 (N_25478,N_21569,N_23670);
nand U25479 (N_25479,N_23227,N_23797);
and U25480 (N_25480,N_21248,N_22125);
nor U25481 (N_25481,N_23129,N_23158);
xor U25482 (N_25482,N_23103,N_21848);
or U25483 (N_25483,N_23336,N_23173);
nand U25484 (N_25484,N_23433,N_21234);
nor U25485 (N_25485,N_21514,N_23595);
and U25486 (N_25486,N_23866,N_21469);
and U25487 (N_25487,N_23346,N_21797);
or U25488 (N_25488,N_23612,N_21045);
and U25489 (N_25489,N_22391,N_21367);
or U25490 (N_25490,N_22378,N_23810);
or U25491 (N_25491,N_23418,N_21396);
or U25492 (N_25492,N_22734,N_23730);
or U25493 (N_25493,N_22990,N_21964);
nor U25494 (N_25494,N_23376,N_22048);
and U25495 (N_25495,N_22438,N_23322);
xor U25496 (N_25496,N_23210,N_22063);
and U25497 (N_25497,N_22524,N_22578);
nand U25498 (N_25498,N_23071,N_22668);
and U25499 (N_25499,N_22182,N_22256);
and U25500 (N_25500,N_23220,N_22848);
and U25501 (N_25501,N_21320,N_23686);
or U25502 (N_25502,N_23518,N_23216);
and U25503 (N_25503,N_22141,N_21187);
and U25504 (N_25504,N_21079,N_21205);
nor U25505 (N_25505,N_23215,N_21617);
nand U25506 (N_25506,N_21483,N_22847);
xnor U25507 (N_25507,N_21924,N_23275);
and U25508 (N_25508,N_21061,N_23555);
nand U25509 (N_25509,N_23734,N_23411);
and U25510 (N_25510,N_22530,N_22035);
nor U25511 (N_25511,N_21000,N_21328);
and U25512 (N_25512,N_21303,N_21902);
xnor U25513 (N_25513,N_22841,N_21973);
nand U25514 (N_25514,N_21869,N_21637);
nor U25515 (N_25515,N_23979,N_23110);
nand U25516 (N_25516,N_21962,N_21326);
nand U25517 (N_25517,N_21127,N_21920);
nor U25518 (N_25518,N_23896,N_22785);
nand U25519 (N_25519,N_21891,N_22768);
and U25520 (N_25520,N_22554,N_22325);
nor U25521 (N_25521,N_22309,N_22522);
and U25522 (N_25522,N_23395,N_21864);
or U25523 (N_25523,N_21998,N_23064);
or U25524 (N_25524,N_23042,N_21454);
nor U25525 (N_25525,N_22652,N_22601);
nor U25526 (N_25526,N_23448,N_21994);
nor U25527 (N_25527,N_22146,N_23319);
xor U25528 (N_25528,N_22126,N_23115);
xor U25529 (N_25529,N_23948,N_23814);
or U25530 (N_25530,N_23889,N_21357);
or U25531 (N_25531,N_21822,N_23655);
nand U25532 (N_25532,N_21130,N_22803);
xor U25533 (N_25533,N_23401,N_22450);
nor U25534 (N_25534,N_22330,N_22588);
nand U25535 (N_25535,N_22062,N_21707);
nor U25536 (N_25536,N_23498,N_23543);
or U25537 (N_25537,N_23621,N_21766);
xnor U25538 (N_25538,N_22406,N_23228);
nand U25539 (N_25539,N_22035,N_21294);
or U25540 (N_25540,N_21224,N_22463);
or U25541 (N_25541,N_22669,N_23856);
or U25542 (N_25542,N_23067,N_23080);
and U25543 (N_25543,N_21487,N_21062);
nand U25544 (N_25544,N_22794,N_21242);
nand U25545 (N_25545,N_21249,N_22706);
nand U25546 (N_25546,N_22332,N_23790);
nor U25547 (N_25547,N_23087,N_21804);
nor U25548 (N_25548,N_22278,N_21731);
xnor U25549 (N_25549,N_22362,N_21482);
and U25550 (N_25550,N_23931,N_22872);
and U25551 (N_25551,N_22995,N_23661);
nor U25552 (N_25552,N_23161,N_21023);
and U25553 (N_25553,N_22733,N_23770);
and U25554 (N_25554,N_21622,N_23784);
and U25555 (N_25555,N_23404,N_21092);
xnor U25556 (N_25556,N_22711,N_21234);
nand U25557 (N_25557,N_23528,N_21588);
xor U25558 (N_25558,N_21516,N_21735);
xnor U25559 (N_25559,N_22759,N_21081);
nand U25560 (N_25560,N_21605,N_22202);
xnor U25561 (N_25561,N_23015,N_22303);
nor U25562 (N_25562,N_23805,N_23353);
nand U25563 (N_25563,N_22901,N_23209);
nand U25564 (N_25564,N_22187,N_21467);
nor U25565 (N_25565,N_22478,N_22636);
xnor U25566 (N_25566,N_23709,N_21379);
and U25567 (N_25567,N_22518,N_21847);
and U25568 (N_25568,N_23895,N_23718);
and U25569 (N_25569,N_23897,N_21132);
or U25570 (N_25570,N_23040,N_21393);
nand U25571 (N_25571,N_23788,N_21032);
and U25572 (N_25572,N_21048,N_23481);
or U25573 (N_25573,N_23234,N_22116);
and U25574 (N_25574,N_22847,N_21454);
and U25575 (N_25575,N_22755,N_21908);
nand U25576 (N_25576,N_21767,N_22609);
nand U25577 (N_25577,N_21429,N_23305);
nand U25578 (N_25578,N_21718,N_23698);
nand U25579 (N_25579,N_23661,N_22426);
and U25580 (N_25580,N_21669,N_22746);
and U25581 (N_25581,N_23711,N_21383);
nor U25582 (N_25582,N_23677,N_23036);
nand U25583 (N_25583,N_23836,N_23529);
or U25584 (N_25584,N_23802,N_22066);
nand U25585 (N_25585,N_21711,N_22602);
and U25586 (N_25586,N_21305,N_22484);
xor U25587 (N_25587,N_21563,N_21681);
xor U25588 (N_25588,N_21921,N_21983);
and U25589 (N_25589,N_23057,N_23113);
and U25590 (N_25590,N_22116,N_21550);
and U25591 (N_25591,N_22638,N_21943);
nand U25592 (N_25592,N_23810,N_21685);
nor U25593 (N_25593,N_22064,N_21860);
or U25594 (N_25594,N_21270,N_23229);
or U25595 (N_25595,N_22589,N_23103);
xnor U25596 (N_25596,N_21138,N_22957);
xnor U25597 (N_25597,N_22199,N_23391);
xnor U25598 (N_25598,N_21117,N_23048);
nor U25599 (N_25599,N_23042,N_21955);
xnor U25600 (N_25600,N_21467,N_21531);
nand U25601 (N_25601,N_23514,N_23553);
or U25602 (N_25602,N_23819,N_21191);
xnor U25603 (N_25603,N_21821,N_23505);
or U25604 (N_25604,N_21024,N_22799);
or U25605 (N_25605,N_23171,N_22077);
nand U25606 (N_25606,N_21998,N_22929);
and U25607 (N_25607,N_23587,N_21546);
or U25608 (N_25608,N_23243,N_21386);
nand U25609 (N_25609,N_21710,N_23610);
or U25610 (N_25610,N_22122,N_22437);
xnor U25611 (N_25611,N_22693,N_23437);
xnor U25612 (N_25612,N_21590,N_22084);
and U25613 (N_25613,N_23479,N_22056);
nand U25614 (N_25614,N_23085,N_22248);
nand U25615 (N_25615,N_21432,N_21868);
and U25616 (N_25616,N_22613,N_21217);
or U25617 (N_25617,N_23230,N_23279);
and U25618 (N_25618,N_21046,N_22523);
and U25619 (N_25619,N_21476,N_23976);
nand U25620 (N_25620,N_23513,N_22808);
xor U25621 (N_25621,N_22037,N_21332);
nand U25622 (N_25622,N_21794,N_22882);
and U25623 (N_25623,N_21573,N_23476);
xnor U25624 (N_25624,N_22505,N_23552);
xor U25625 (N_25625,N_21677,N_23976);
or U25626 (N_25626,N_22013,N_22172);
nor U25627 (N_25627,N_23194,N_21273);
nand U25628 (N_25628,N_22423,N_21103);
nor U25629 (N_25629,N_21862,N_21327);
xor U25630 (N_25630,N_21518,N_21382);
xnor U25631 (N_25631,N_22912,N_23478);
or U25632 (N_25632,N_22440,N_23890);
nand U25633 (N_25633,N_22284,N_21932);
nand U25634 (N_25634,N_23163,N_22285);
nor U25635 (N_25635,N_23183,N_22393);
nand U25636 (N_25636,N_22737,N_23521);
and U25637 (N_25637,N_22305,N_21477);
xor U25638 (N_25638,N_22023,N_23809);
nand U25639 (N_25639,N_23237,N_22587);
xnor U25640 (N_25640,N_22972,N_23169);
and U25641 (N_25641,N_23618,N_23632);
and U25642 (N_25642,N_22339,N_22578);
xnor U25643 (N_25643,N_22171,N_21800);
nand U25644 (N_25644,N_22251,N_22945);
and U25645 (N_25645,N_21746,N_22120);
nor U25646 (N_25646,N_23164,N_21384);
nand U25647 (N_25647,N_21371,N_22688);
and U25648 (N_25648,N_22347,N_23896);
xor U25649 (N_25649,N_23043,N_21629);
or U25650 (N_25650,N_21421,N_21520);
nand U25651 (N_25651,N_21328,N_23823);
nor U25652 (N_25652,N_22892,N_22897);
or U25653 (N_25653,N_23844,N_23682);
nand U25654 (N_25654,N_23152,N_22503);
nor U25655 (N_25655,N_21913,N_21554);
or U25656 (N_25656,N_23597,N_22374);
xor U25657 (N_25657,N_22653,N_23939);
nand U25658 (N_25658,N_22754,N_22944);
or U25659 (N_25659,N_23526,N_23361);
nor U25660 (N_25660,N_21277,N_21044);
xor U25661 (N_25661,N_23183,N_21530);
xnor U25662 (N_25662,N_23945,N_22060);
or U25663 (N_25663,N_23519,N_22622);
nor U25664 (N_25664,N_22670,N_21796);
and U25665 (N_25665,N_21398,N_21410);
nor U25666 (N_25666,N_23526,N_23969);
xnor U25667 (N_25667,N_21715,N_23833);
nor U25668 (N_25668,N_23950,N_23627);
or U25669 (N_25669,N_21686,N_23159);
nand U25670 (N_25670,N_22334,N_21781);
nor U25671 (N_25671,N_23588,N_23409);
nand U25672 (N_25672,N_23760,N_23123);
or U25673 (N_25673,N_22147,N_22189);
xnor U25674 (N_25674,N_23307,N_21916);
xor U25675 (N_25675,N_23382,N_22451);
xnor U25676 (N_25676,N_21634,N_22329);
and U25677 (N_25677,N_23883,N_23256);
xor U25678 (N_25678,N_21622,N_23930);
or U25679 (N_25679,N_23071,N_23687);
or U25680 (N_25680,N_22730,N_22867);
xnor U25681 (N_25681,N_22531,N_23698);
and U25682 (N_25682,N_21211,N_21554);
nor U25683 (N_25683,N_22835,N_22245);
or U25684 (N_25684,N_23646,N_23148);
and U25685 (N_25685,N_22893,N_23214);
nand U25686 (N_25686,N_21344,N_22790);
xor U25687 (N_25687,N_21480,N_22711);
and U25688 (N_25688,N_21597,N_21593);
nor U25689 (N_25689,N_23379,N_22091);
nor U25690 (N_25690,N_22648,N_23292);
and U25691 (N_25691,N_21123,N_22850);
nor U25692 (N_25692,N_22295,N_23237);
xnor U25693 (N_25693,N_21377,N_23994);
nand U25694 (N_25694,N_21769,N_22697);
and U25695 (N_25695,N_22907,N_23898);
and U25696 (N_25696,N_23924,N_21764);
nor U25697 (N_25697,N_23237,N_22513);
and U25698 (N_25698,N_21854,N_21070);
or U25699 (N_25699,N_22325,N_21904);
and U25700 (N_25700,N_22678,N_22576);
nand U25701 (N_25701,N_21879,N_23555);
and U25702 (N_25702,N_21016,N_21882);
or U25703 (N_25703,N_22210,N_23588);
nand U25704 (N_25704,N_23994,N_23919);
nor U25705 (N_25705,N_23423,N_22591);
and U25706 (N_25706,N_21067,N_23605);
nor U25707 (N_25707,N_22344,N_23212);
nand U25708 (N_25708,N_23782,N_22606);
xor U25709 (N_25709,N_21180,N_21181);
nand U25710 (N_25710,N_22657,N_23669);
xor U25711 (N_25711,N_22393,N_23321);
or U25712 (N_25712,N_21874,N_23557);
xor U25713 (N_25713,N_23345,N_22450);
nand U25714 (N_25714,N_21628,N_21749);
xnor U25715 (N_25715,N_22442,N_21222);
and U25716 (N_25716,N_23815,N_22092);
nor U25717 (N_25717,N_23778,N_21944);
xor U25718 (N_25718,N_23393,N_21035);
nand U25719 (N_25719,N_23897,N_22296);
nor U25720 (N_25720,N_22853,N_21811);
xor U25721 (N_25721,N_22452,N_21229);
nand U25722 (N_25722,N_21314,N_22317);
nand U25723 (N_25723,N_23000,N_21640);
nand U25724 (N_25724,N_22779,N_21080);
nand U25725 (N_25725,N_22529,N_22362);
nor U25726 (N_25726,N_22061,N_22488);
or U25727 (N_25727,N_21182,N_21958);
and U25728 (N_25728,N_23277,N_23055);
or U25729 (N_25729,N_21506,N_21375);
and U25730 (N_25730,N_22634,N_23220);
nor U25731 (N_25731,N_22761,N_23564);
and U25732 (N_25732,N_21894,N_21910);
nand U25733 (N_25733,N_22456,N_22308);
nand U25734 (N_25734,N_21172,N_21482);
or U25735 (N_25735,N_21171,N_21298);
or U25736 (N_25736,N_21943,N_22466);
and U25737 (N_25737,N_22734,N_21488);
nand U25738 (N_25738,N_23427,N_21687);
xnor U25739 (N_25739,N_21798,N_21511);
nand U25740 (N_25740,N_23284,N_23728);
xnor U25741 (N_25741,N_21849,N_23249);
or U25742 (N_25742,N_22376,N_22738);
and U25743 (N_25743,N_21784,N_23277);
xnor U25744 (N_25744,N_22988,N_21216);
and U25745 (N_25745,N_21095,N_23295);
and U25746 (N_25746,N_22681,N_22734);
xor U25747 (N_25747,N_21729,N_21893);
or U25748 (N_25748,N_22412,N_23339);
and U25749 (N_25749,N_22041,N_22567);
xor U25750 (N_25750,N_23817,N_21167);
nand U25751 (N_25751,N_22176,N_23857);
nand U25752 (N_25752,N_23168,N_23107);
nor U25753 (N_25753,N_22713,N_23971);
nand U25754 (N_25754,N_21040,N_23649);
nand U25755 (N_25755,N_23995,N_21376);
or U25756 (N_25756,N_21258,N_21280);
nand U25757 (N_25757,N_21165,N_23213);
nor U25758 (N_25758,N_23656,N_22039);
nand U25759 (N_25759,N_23667,N_22233);
xnor U25760 (N_25760,N_23352,N_23940);
and U25761 (N_25761,N_22422,N_22839);
xnor U25762 (N_25762,N_21265,N_23934);
nor U25763 (N_25763,N_23054,N_21793);
nor U25764 (N_25764,N_23989,N_23887);
and U25765 (N_25765,N_21225,N_22606);
and U25766 (N_25766,N_23866,N_23892);
nand U25767 (N_25767,N_23622,N_22482);
xor U25768 (N_25768,N_23135,N_21302);
nand U25769 (N_25769,N_22584,N_23004);
nand U25770 (N_25770,N_22487,N_22387);
nand U25771 (N_25771,N_21509,N_22173);
and U25772 (N_25772,N_22721,N_23775);
nand U25773 (N_25773,N_21458,N_23813);
nand U25774 (N_25774,N_21289,N_22023);
and U25775 (N_25775,N_21197,N_23501);
nor U25776 (N_25776,N_22615,N_21151);
nor U25777 (N_25777,N_23502,N_22881);
or U25778 (N_25778,N_22859,N_23320);
xnor U25779 (N_25779,N_22652,N_22965);
nand U25780 (N_25780,N_23519,N_21291);
and U25781 (N_25781,N_23584,N_22571);
nand U25782 (N_25782,N_21291,N_23105);
or U25783 (N_25783,N_23051,N_22700);
xnor U25784 (N_25784,N_21074,N_21547);
xnor U25785 (N_25785,N_22019,N_21490);
xor U25786 (N_25786,N_23332,N_22057);
and U25787 (N_25787,N_22575,N_22826);
or U25788 (N_25788,N_22554,N_23158);
xnor U25789 (N_25789,N_21587,N_22837);
or U25790 (N_25790,N_21398,N_22488);
or U25791 (N_25791,N_23947,N_23078);
xor U25792 (N_25792,N_21054,N_21246);
or U25793 (N_25793,N_23080,N_23610);
or U25794 (N_25794,N_21729,N_21488);
or U25795 (N_25795,N_22502,N_22586);
nor U25796 (N_25796,N_23526,N_21409);
nand U25797 (N_25797,N_22038,N_22456);
nor U25798 (N_25798,N_22951,N_23421);
xor U25799 (N_25799,N_22027,N_23242);
and U25800 (N_25800,N_21175,N_22877);
and U25801 (N_25801,N_22876,N_22211);
xor U25802 (N_25802,N_21835,N_23574);
nand U25803 (N_25803,N_23761,N_21088);
xor U25804 (N_25804,N_22897,N_23759);
nor U25805 (N_25805,N_23949,N_23545);
or U25806 (N_25806,N_21545,N_22116);
or U25807 (N_25807,N_21807,N_21394);
nand U25808 (N_25808,N_22027,N_21892);
xor U25809 (N_25809,N_23700,N_23588);
nand U25810 (N_25810,N_22211,N_23387);
nand U25811 (N_25811,N_21236,N_21174);
xor U25812 (N_25812,N_22598,N_23341);
nand U25813 (N_25813,N_23835,N_23869);
xnor U25814 (N_25814,N_23052,N_22150);
or U25815 (N_25815,N_22210,N_22744);
or U25816 (N_25816,N_22989,N_21869);
nor U25817 (N_25817,N_23705,N_22088);
or U25818 (N_25818,N_21868,N_21988);
and U25819 (N_25819,N_22137,N_21514);
nor U25820 (N_25820,N_22223,N_22236);
xnor U25821 (N_25821,N_23147,N_22456);
or U25822 (N_25822,N_21096,N_22224);
xor U25823 (N_25823,N_22183,N_22407);
nor U25824 (N_25824,N_22390,N_22274);
and U25825 (N_25825,N_22868,N_21426);
nor U25826 (N_25826,N_23181,N_23443);
nand U25827 (N_25827,N_21073,N_21262);
or U25828 (N_25828,N_22421,N_22860);
and U25829 (N_25829,N_21990,N_22432);
xor U25830 (N_25830,N_23079,N_22409);
nand U25831 (N_25831,N_22671,N_22378);
or U25832 (N_25832,N_21154,N_21289);
nand U25833 (N_25833,N_22548,N_23530);
nor U25834 (N_25834,N_21636,N_21642);
nand U25835 (N_25835,N_22998,N_22063);
or U25836 (N_25836,N_21223,N_22308);
xor U25837 (N_25837,N_22055,N_23081);
nor U25838 (N_25838,N_21044,N_23870);
or U25839 (N_25839,N_23993,N_22554);
nand U25840 (N_25840,N_21544,N_23604);
nor U25841 (N_25841,N_21911,N_21655);
or U25842 (N_25842,N_23494,N_21515);
or U25843 (N_25843,N_22076,N_21302);
and U25844 (N_25844,N_21536,N_23684);
or U25845 (N_25845,N_23075,N_22092);
and U25846 (N_25846,N_23498,N_22007);
nor U25847 (N_25847,N_21742,N_21158);
or U25848 (N_25848,N_23931,N_23488);
and U25849 (N_25849,N_23485,N_21767);
nand U25850 (N_25850,N_22682,N_23909);
xor U25851 (N_25851,N_21742,N_22680);
xor U25852 (N_25852,N_22153,N_21660);
nor U25853 (N_25853,N_21940,N_23900);
xnor U25854 (N_25854,N_22496,N_22407);
nor U25855 (N_25855,N_22528,N_22256);
and U25856 (N_25856,N_23460,N_23946);
or U25857 (N_25857,N_23504,N_21554);
xnor U25858 (N_25858,N_22800,N_22042);
nand U25859 (N_25859,N_23217,N_21870);
nor U25860 (N_25860,N_23367,N_23243);
and U25861 (N_25861,N_21517,N_22600);
xor U25862 (N_25862,N_22903,N_23564);
nand U25863 (N_25863,N_23367,N_23130);
and U25864 (N_25864,N_23509,N_22054);
or U25865 (N_25865,N_22766,N_23728);
or U25866 (N_25866,N_21809,N_22803);
or U25867 (N_25867,N_23606,N_21456);
nand U25868 (N_25868,N_23863,N_23151);
or U25869 (N_25869,N_21985,N_22950);
nor U25870 (N_25870,N_22151,N_22627);
or U25871 (N_25871,N_21665,N_22427);
and U25872 (N_25872,N_23305,N_22051);
or U25873 (N_25873,N_21898,N_21748);
or U25874 (N_25874,N_23733,N_23723);
xor U25875 (N_25875,N_22092,N_22155);
and U25876 (N_25876,N_23936,N_22152);
or U25877 (N_25877,N_23697,N_23755);
or U25878 (N_25878,N_21348,N_23323);
nand U25879 (N_25879,N_23249,N_22049);
or U25880 (N_25880,N_22742,N_22823);
or U25881 (N_25881,N_23009,N_21146);
xnor U25882 (N_25882,N_22361,N_21244);
xnor U25883 (N_25883,N_23286,N_21758);
xor U25884 (N_25884,N_22374,N_23357);
and U25885 (N_25885,N_21237,N_22974);
nor U25886 (N_25886,N_21899,N_21111);
or U25887 (N_25887,N_22712,N_21022);
and U25888 (N_25888,N_22848,N_22612);
and U25889 (N_25889,N_22727,N_22970);
and U25890 (N_25890,N_21695,N_22404);
nor U25891 (N_25891,N_23975,N_22286);
or U25892 (N_25892,N_22787,N_21016);
or U25893 (N_25893,N_22663,N_22474);
nand U25894 (N_25894,N_23054,N_21047);
xor U25895 (N_25895,N_23599,N_23358);
nor U25896 (N_25896,N_23447,N_23575);
nand U25897 (N_25897,N_23804,N_22082);
xor U25898 (N_25898,N_21185,N_21312);
and U25899 (N_25899,N_23944,N_21005);
nand U25900 (N_25900,N_22718,N_21361);
or U25901 (N_25901,N_22752,N_21544);
and U25902 (N_25902,N_23698,N_22748);
xnor U25903 (N_25903,N_23409,N_22524);
xnor U25904 (N_25904,N_23568,N_23062);
xnor U25905 (N_25905,N_21247,N_23585);
or U25906 (N_25906,N_22427,N_21833);
or U25907 (N_25907,N_22965,N_21240);
xnor U25908 (N_25908,N_21065,N_22392);
and U25909 (N_25909,N_21083,N_23369);
or U25910 (N_25910,N_22888,N_21055);
nand U25911 (N_25911,N_23790,N_21517);
or U25912 (N_25912,N_22487,N_21490);
nand U25913 (N_25913,N_23366,N_22784);
nand U25914 (N_25914,N_23392,N_22111);
nor U25915 (N_25915,N_23096,N_23918);
xor U25916 (N_25916,N_21771,N_21786);
or U25917 (N_25917,N_23768,N_23274);
xor U25918 (N_25918,N_22658,N_23734);
xnor U25919 (N_25919,N_23175,N_21481);
nor U25920 (N_25920,N_23093,N_23701);
nand U25921 (N_25921,N_23643,N_21409);
nand U25922 (N_25922,N_23307,N_21964);
and U25923 (N_25923,N_22915,N_23035);
nor U25924 (N_25924,N_21490,N_23529);
xnor U25925 (N_25925,N_21272,N_22504);
nand U25926 (N_25926,N_21074,N_23613);
nor U25927 (N_25927,N_23735,N_22281);
nor U25928 (N_25928,N_23356,N_22003);
xor U25929 (N_25929,N_23469,N_21525);
or U25930 (N_25930,N_23549,N_21855);
or U25931 (N_25931,N_23283,N_22035);
nor U25932 (N_25932,N_23138,N_21053);
nand U25933 (N_25933,N_22178,N_21456);
xnor U25934 (N_25934,N_21554,N_23951);
nor U25935 (N_25935,N_22788,N_22185);
or U25936 (N_25936,N_22280,N_23710);
and U25937 (N_25937,N_22416,N_23043);
nor U25938 (N_25938,N_22902,N_21189);
and U25939 (N_25939,N_22006,N_21475);
nor U25940 (N_25940,N_23194,N_22389);
and U25941 (N_25941,N_21566,N_21945);
xor U25942 (N_25942,N_22193,N_22534);
nor U25943 (N_25943,N_21365,N_23734);
and U25944 (N_25944,N_23969,N_22383);
nand U25945 (N_25945,N_23714,N_22003);
nor U25946 (N_25946,N_22804,N_22795);
and U25947 (N_25947,N_23025,N_21474);
nor U25948 (N_25948,N_21525,N_22722);
xnor U25949 (N_25949,N_23721,N_21413);
and U25950 (N_25950,N_22537,N_23153);
or U25951 (N_25951,N_23376,N_23221);
nand U25952 (N_25952,N_22246,N_21527);
and U25953 (N_25953,N_21560,N_21016);
nand U25954 (N_25954,N_22435,N_22417);
or U25955 (N_25955,N_21713,N_21547);
or U25956 (N_25956,N_23426,N_21805);
nor U25957 (N_25957,N_22851,N_22063);
xnor U25958 (N_25958,N_21995,N_23621);
nor U25959 (N_25959,N_21419,N_21461);
and U25960 (N_25960,N_23197,N_23957);
and U25961 (N_25961,N_22500,N_21264);
nor U25962 (N_25962,N_22490,N_21878);
or U25963 (N_25963,N_23435,N_22155);
or U25964 (N_25964,N_21816,N_21431);
nand U25965 (N_25965,N_23336,N_23563);
or U25966 (N_25966,N_22825,N_22319);
nor U25967 (N_25967,N_22951,N_23172);
nor U25968 (N_25968,N_22990,N_22690);
nand U25969 (N_25969,N_21709,N_21453);
or U25970 (N_25970,N_21190,N_21027);
nor U25971 (N_25971,N_22557,N_21849);
nand U25972 (N_25972,N_21871,N_22517);
and U25973 (N_25973,N_22006,N_21904);
nor U25974 (N_25974,N_23392,N_21884);
or U25975 (N_25975,N_21029,N_21319);
and U25976 (N_25976,N_22013,N_21166);
nand U25977 (N_25977,N_23639,N_21054);
or U25978 (N_25978,N_21801,N_21548);
nor U25979 (N_25979,N_23514,N_23450);
or U25980 (N_25980,N_23952,N_21971);
nor U25981 (N_25981,N_23946,N_23681);
or U25982 (N_25982,N_21300,N_21584);
nor U25983 (N_25983,N_22578,N_23993);
nand U25984 (N_25984,N_23160,N_22210);
nand U25985 (N_25985,N_23322,N_21057);
nor U25986 (N_25986,N_21347,N_23251);
nand U25987 (N_25987,N_21004,N_22721);
nor U25988 (N_25988,N_22213,N_21456);
xor U25989 (N_25989,N_22436,N_21587);
nor U25990 (N_25990,N_21572,N_21746);
xnor U25991 (N_25991,N_22357,N_22639);
nor U25992 (N_25992,N_22130,N_21648);
nor U25993 (N_25993,N_21159,N_21592);
xnor U25994 (N_25994,N_22598,N_21765);
xor U25995 (N_25995,N_21826,N_21112);
nor U25996 (N_25996,N_22269,N_23843);
or U25997 (N_25997,N_22001,N_23233);
nor U25998 (N_25998,N_23694,N_22846);
xnor U25999 (N_25999,N_23312,N_22825);
and U26000 (N_26000,N_21442,N_23398);
nor U26001 (N_26001,N_23193,N_23223);
nand U26002 (N_26002,N_23022,N_21716);
or U26003 (N_26003,N_22141,N_22721);
nor U26004 (N_26004,N_23187,N_21467);
xor U26005 (N_26005,N_23797,N_23504);
nand U26006 (N_26006,N_23178,N_21996);
xor U26007 (N_26007,N_23759,N_21802);
nand U26008 (N_26008,N_23289,N_23996);
and U26009 (N_26009,N_23823,N_21388);
nand U26010 (N_26010,N_21143,N_23719);
and U26011 (N_26011,N_21919,N_23706);
xnor U26012 (N_26012,N_23622,N_22208);
and U26013 (N_26013,N_21443,N_21947);
nor U26014 (N_26014,N_22181,N_21143);
xor U26015 (N_26015,N_22767,N_23561);
nor U26016 (N_26016,N_23904,N_22664);
nand U26017 (N_26017,N_23444,N_21699);
xnor U26018 (N_26018,N_23557,N_23683);
nor U26019 (N_26019,N_21418,N_23303);
or U26020 (N_26020,N_22656,N_23896);
nand U26021 (N_26021,N_21518,N_21961);
or U26022 (N_26022,N_21357,N_22821);
or U26023 (N_26023,N_22612,N_21226);
nor U26024 (N_26024,N_21241,N_23077);
nor U26025 (N_26025,N_21792,N_23142);
nor U26026 (N_26026,N_22684,N_21327);
xnor U26027 (N_26027,N_22552,N_23703);
xnor U26028 (N_26028,N_23957,N_22743);
or U26029 (N_26029,N_22701,N_21893);
xnor U26030 (N_26030,N_21269,N_22133);
xor U26031 (N_26031,N_21002,N_23006);
xor U26032 (N_26032,N_21401,N_23901);
and U26033 (N_26033,N_22176,N_22486);
nor U26034 (N_26034,N_21626,N_21576);
xor U26035 (N_26035,N_23555,N_23006);
xnor U26036 (N_26036,N_23849,N_23653);
nand U26037 (N_26037,N_21432,N_23892);
and U26038 (N_26038,N_22658,N_21779);
nor U26039 (N_26039,N_23424,N_22295);
nor U26040 (N_26040,N_23685,N_22781);
and U26041 (N_26041,N_22183,N_21779);
nor U26042 (N_26042,N_21000,N_22338);
nor U26043 (N_26043,N_21079,N_21373);
nor U26044 (N_26044,N_21192,N_22795);
nor U26045 (N_26045,N_21056,N_22937);
xor U26046 (N_26046,N_21888,N_22665);
nor U26047 (N_26047,N_23759,N_22457);
and U26048 (N_26048,N_23762,N_22850);
nand U26049 (N_26049,N_21061,N_21493);
and U26050 (N_26050,N_22498,N_22838);
nand U26051 (N_26051,N_21451,N_21440);
xor U26052 (N_26052,N_22299,N_23520);
and U26053 (N_26053,N_22905,N_22582);
xnor U26054 (N_26054,N_22862,N_21641);
xor U26055 (N_26055,N_22611,N_22039);
and U26056 (N_26056,N_23060,N_23444);
or U26057 (N_26057,N_23091,N_21585);
and U26058 (N_26058,N_22160,N_22202);
or U26059 (N_26059,N_21468,N_22152);
xnor U26060 (N_26060,N_22291,N_23563);
nand U26061 (N_26061,N_23368,N_22933);
or U26062 (N_26062,N_21659,N_21891);
or U26063 (N_26063,N_21256,N_21316);
nand U26064 (N_26064,N_23428,N_22561);
xnor U26065 (N_26065,N_21447,N_22676);
nand U26066 (N_26066,N_23897,N_21386);
and U26067 (N_26067,N_22179,N_23499);
xnor U26068 (N_26068,N_21796,N_23515);
or U26069 (N_26069,N_23400,N_23872);
nor U26070 (N_26070,N_23640,N_22308);
nand U26071 (N_26071,N_23212,N_21612);
and U26072 (N_26072,N_22217,N_22433);
nor U26073 (N_26073,N_23498,N_23358);
nand U26074 (N_26074,N_22132,N_22220);
nor U26075 (N_26075,N_21877,N_21572);
xor U26076 (N_26076,N_21581,N_21449);
xnor U26077 (N_26077,N_23223,N_21354);
nor U26078 (N_26078,N_23449,N_21287);
or U26079 (N_26079,N_21305,N_23203);
nand U26080 (N_26080,N_22420,N_23787);
and U26081 (N_26081,N_23957,N_23525);
xor U26082 (N_26082,N_21473,N_22717);
xor U26083 (N_26083,N_22344,N_23799);
and U26084 (N_26084,N_23148,N_22977);
or U26085 (N_26085,N_22639,N_22260);
and U26086 (N_26086,N_22442,N_21377);
nand U26087 (N_26087,N_23331,N_23753);
nand U26088 (N_26088,N_22652,N_21217);
nand U26089 (N_26089,N_23882,N_21467);
or U26090 (N_26090,N_21097,N_22277);
and U26091 (N_26091,N_23009,N_23503);
nand U26092 (N_26092,N_23421,N_21368);
nor U26093 (N_26093,N_21181,N_23399);
or U26094 (N_26094,N_23893,N_22540);
or U26095 (N_26095,N_22849,N_23588);
nor U26096 (N_26096,N_23084,N_22188);
or U26097 (N_26097,N_22624,N_21144);
or U26098 (N_26098,N_23900,N_22786);
or U26099 (N_26099,N_22035,N_22911);
or U26100 (N_26100,N_21138,N_23649);
nor U26101 (N_26101,N_23463,N_22165);
nand U26102 (N_26102,N_21942,N_21493);
nor U26103 (N_26103,N_23367,N_23607);
xnor U26104 (N_26104,N_21848,N_23693);
and U26105 (N_26105,N_21728,N_23033);
and U26106 (N_26106,N_22616,N_23817);
and U26107 (N_26107,N_22284,N_21264);
nand U26108 (N_26108,N_22221,N_23711);
nand U26109 (N_26109,N_23214,N_23704);
or U26110 (N_26110,N_21335,N_22419);
or U26111 (N_26111,N_23013,N_23543);
nand U26112 (N_26112,N_23873,N_21015);
or U26113 (N_26113,N_21553,N_23725);
nand U26114 (N_26114,N_22356,N_23864);
or U26115 (N_26115,N_22992,N_22923);
nand U26116 (N_26116,N_21861,N_23578);
nand U26117 (N_26117,N_23554,N_23810);
xnor U26118 (N_26118,N_22821,N_22460);
nor U26119 (N_26119,N_22064,N_23622);
nor U26120 (N_26120,N_21806,N_22784);
or U26121 (N_26121,N_21858,N_23776);
nor U26122 (N_26122,N_21925,N_23576);
or U26123 (N_26123,N_23619,N_23595);
nor U26124 (N_26124,N_23268,N_21371);
xnor U26125 (N_26125,N_21899,N_23785);
nor U26126 (N_26126,N_21279,N_21481);
and U26127 (N_26127,N_23329,N_23188);
nor U26128 (N_26128,N_21331,N_22197);
xnor U26129 (N_26129,N_21058,N_21865);
or U26130 (N_26130,N_22434,N_22407);
and U26131 (N_26131,N_23021,N_22910);
xnor U26132 (N_26132,N_22326,N_22762);
and U26133 (N_26133,N_23521,N_23976);
xor U26134 (N_26134,N_22368,N_21742);
or U26135 (N_26135,N_23574,N_21322);
or U26136 (N_26136,N_21982,N_21306);
nor U26137 (N_26137,N_21810,N_21989);
nor U26138 (N_26138,N_21432,N_23773);
nor U26139 (N_26139,N_22810,N_23545);
xor U26140 (N_26140,N_23661,N_21728);
or U26141 (N_26141,N_22449,N_22344);
and U26142 (N_26142,N_21343,N_23582);
xnor U26143 (N_26143,N_22218,N_22272);
and U26144 (N_26144,N_23768,N_22899);
nor U26145 (N_26145,N_21143,N_22260);
nand U26146 (N_26146,N_23940,N_23065);
or U26147 (N_26147,N_23289,N_21952);
and U26148 (N_26148,N_23389,N_21761);
nor U26149 (N_26149,N_23811,N_21177);
xor U26150 (N_26150,N_22095,N_23219);
nor U26151 (N_26151,N_23524,N_21546);
nand U26152 (N_26152,N_23516,N_22433);
nand U26153 (N_26153,N_23824,N_23831);
nor U26154 (N_26154,N_23399,N_23190);
and U26155 (N_26155,N_22793,N_21849);
nor U26156 (N_26156,N_21304,N_23851);
xnor U26157 (N_26157,N_22411,N_22039);
or U26158 (N_26158,N_22237,N_22574);
xnor U26159 (N_26159,N_23442,N_21537);
nor U26160 (N_26160,N_23503,N_21226);
or U26161 (N_26161,N_22483,N_21587);
or U26162 (N_26162,N_23304,N_22585);
nor U26163 (N_26163,N_21599,N_22287);
or U26164 (N_26164,N_21391,N_22725);
and U26165 (N_26165,N_23306,N_23388);
nand U26166 (N_26166,N_21894,N_21181);
and U26167 (N_26167,N_23816,N_21216);
and U26168 (N_26168,N_23847,N_23644);
xnor U26169 (N_26169,N_23439,N_21598);
nor U26170 (N_26170,N_21263,N_22574);
nand U26171 (N_26171,N_23750,N_22370);
nor U26172 (N_26172,N_23425,N_22849);
or U26173 (N_26173,N_21087,N_23457);
nand U26174 (N_26174,N_22626,N_23804);
and U26175 (N_26175,N_23747,N_22227);
or U26176 (N_26176,N_22005,N_22940);
xnor U26177 (N_26177,N_22538,N_23754);
nand U26178 (N_26178,N_21346,N_23485);
and U26179 (N_26179,N_21748,N_23008);
or U26180 (N_26180,N_21744,N_21460);
nor U26181 (N_26181,N_21581,N_22487);
nor U26182 (N_26182,N_23960,N_21415);
and U26183 (N_26183,N_23043,N_21284);
or U26184 (N_26184,N_22028,N_23833);
nand U26185 (N_26185,N_21350,N_22552);
xor U26186 (N_26186,N_23222,N_21742);
xnor U26187 (N_26187,N_23853,N_22889);
or U26188 (N_26188,N_22958,N_21077);
nor U26189 (N_26189,N_21403,N_22042);
and U26190 (N_26190,N_23789,N_21893);
and U26191 (N_26191,N_23064,N_22743);
and U26192 (N_26192,N_22310,N_22906);
nor U26193 (N_26193,N_21735,N_23834);
xnor U26194 (N_26194,N_21535,N_21314);
xor U26195 (N_26195,N_23006,N_23806);
nand U26196 (N_26196,N_22682,N_21562);
nor U26197 (N_26197,N_23846,N_21090);
nor U26198 (N_26198,N_23728,N_22433);
nand U26199 (N_26199,N_21356,N_22239);
and U26200 (N_26200,N_21758,N_23427);
nand U26201 (N_26201,N_21761,N_22148);
and U26202 (N_26202,N_23577,N_23710);
and U26203 (N_26203,N_22041,N_22403);
nor U26204 (N_26204,N_23918,N_21721);
nor U26205 (N_26205,N_22183,N_21308);
nand U26206 (N_26206,N_23874,N_23462);
or U26207 (N_26207,N_23286,N_23439);
xnor U26208 (N_26208,N_23555,N_22038);
nand U26209 (N_26209,N_22655,N_21500);
and U26210 (N_26210,N_23295,N_22415);
nand U26211 (N_26211,N_21511,N_22866);
nor U26212 (N_26212,N_22728,N_21834);
nand U26213 (N_26213,N_21300,N_21928);
and U26214 (N_26214,N_21569,N_23149);
and U26215 (N_26215,N_21518,N_23837);
or U26216 (N_26216,N_21502,N_23315);
nor U26217 (N_26217,N_23559,N_21691);
xnor U26218 (N_26218,N_21375,N_22808);
and U26219 (N_26219,N_21649,N_22379);
nand U26220 (N_26220,N_22701,N_23971);
xnor U26221 (N_26221,N_21107,N_23175);
nand U26222 (N_26222,N_22529,N_21042);
or U26223 (N_26223,N_21001,N_23479);
and U26224 (N_26224,N_23735,N_23258);
nor U26225 (N_26225,N_22445,N_21324);
nand U26226 (N_26226,N_22814,N_23043);
or U26227 (N_26227,N_21913,N_21711);
xnor U26228 (N_26228,N_21868,N_23706);
nor U26229 (N_26229,N_23180,N_23721);
nand U26230 (N_26230,N_21279,N_23924);
and U26231 (N_26231,N_23282,N_23138);
or U26232 (N_26232,N_22366,N_21617);
or U26233 (N_26233,N_22989,N_22766);
xor U26234 (N_26234,N_22446,N_22261);
nand U26235 (N_26235,N_21905,N_23777);
nor U26236 (N_26236,N_22829,N_21906);
or U26237 (N_26237,N_22040,N_22306);
nor U26238 (N_26238,N_23364,N_23110);
xor U26239 (N_26239,N_21579,N_23825);
nor U26240 (N_26240,N_22226,N_21767);
and U26241 (N_26241,N_22098,N_21954);
and U26242 (N_26242,N_22156,N_23165);
nor U26243 (N_26243,N_22379,N_21948);
nand U26244 (N_26244,N_21484,N_21364);
nand U26245 (N_26245,N_21430,N_21877);
nand U26246 (N_26246,N_21840,N_23037);
nor U26247 (N_26247,N_22303,N_21971);
xnor U26248 (N_26248,N_23641,N_23000);
nand U26249 (N_26249,N_21100,N_21689);
nand U26250 (N_26250,N_21114,N_23183);
nand U26251 (N_26251,N_22249,N_21594);
and U26252 (N_26252,N_23814,N_22679);
nor U26253 (N_26253,N_21167,N_22377);
nor U26254 (N_26254,N_21778,N_21104);
and U26255 (N_26255,N_21404,N_21258);
nand U26256 (N_26256,N_23849,N_23399);
xnor U26257 (N_26257,N_21419,N_23543);
nand U26258 (N_26258,N_21244,N_22360);
nor U26259 (N_26259,N_23623,N_21895);
and U26260 (N_26260,N_22493,N_23476);
nor U26261 (N_26261,N_23723,N_22002);
xnor U26262 (N_26262,N_21246,N_22788);
or U26263 (N_26263,N_21972,N_22485);
and U26264 (N_26264,N_23373,N_23699);
and U26265 (N_26265,N_22361,N_22479);
nor U26266 (N_26266,N_23342,N_22418);
nor U26267 (N_26267,N_21477,N_22368);
nand U26268 (N_26268,N_21478,N_23686);
and U26269 (N_26269,N_22721,N_23830);
or U26270 (N_26270,N_23851,N_23929);
nand U26271 (N_26271,N_23760,N_21119);
nand U26272 (N_26272,N_23306,N_22225);
nand U26273 (N_26273,N_21152,N_22896);
or U26274 (N_26274,N_23164,N_22951);
and U26275 (N_26275,N_23335,N_22180);
or U26276 (N_26276,N_23110,N_22652);
xor U26277 (N_26277,N_21185,N_22926);
nor U26278 (N_26278,N_21725,N_23944);
or U26279 (N_26279,N_23916,N_22729);
xor U26280 (N_26280,N_22586,N_22443);
xor U26281 (N_26281,N_23294,N_23142);
or U26282 (N_26282,N_23574,N_22303);
nand U26283 (N_26283,N_22614,N_22681);
and U26284 (N_26284,N_22742,N_22326);
or U26285 (N_26285,N_21192,N_22144);
nor U26286 (N_26286,N_22019,N_23612);
xor U26287 (N_26287,N_21422,N_23913);
and U26288 (N_26288,N_22130,N_21594);
and U26289 (N_26289,N_23045,N_22241);
or U26290 (N_26290,N_22223,N_23104);
nor U26291 (N_26291,N_23698,N_22267);
or U26292 (N_26292,N_22234,N_22889);
and U26293 (N_26293,N_21030,N_21651);
nand U26294 (N_26294,N_23244,N_23183);
nand U26295 (N_26295,N_22511,N_23274);
nand U26296 (N_26296,N_21522,N_23988);
or U26297 (N_26297,N_21385,N_21856);
nand U26298 (N_26298,N_23082,N_22674);
nor U26299 (N_26299,N_23866,N_23893);
nor U26300 (N_26300,N_21020,N_21573);
xnor U26301 (N_26301,N_21229,N_23041);
and U26302 (N_26302,N_23715,N_23519);
nor U26303 (N_26303,N_23222,N_21367);
nor U26304 (N_26304,N_21421,N_22051);
nand U26305 (N_26305,N_21468,N_21543);
nor U26306 (N_26306,N_23357,N_21654);
and U26307 (N_26307,N_23018,N_22315);
nor U26308 (N_26308,N_22860,N_21178);
xnor U26309 (N_26309,N_22630,N_21602);
nand U26310 (N_26310,N_23688,N_23377);
and U26311 (N_26311,N_22291,N_21542);
nand U26312 (N_26312,N_23073,N_21172);
xnor U26313 (N_26313,N_23106,N_21189);
xor U26314 (N_26314,N_21654,N_22650);
or U26315 (N_26315,N_22157,N_21008);
xor U26316 (N_26316,N_22574,N_23663);
xnor U26317 (N_26317,N_21442,N_22279);
and U26318 (N_26318,N_22735,N_22600);
nand U26319 (N_26319,N_22564,N_22534);
nand U26320 (N_26320,N_21335,N_23477);
or U26321 (N_26321,N_21024,N_22040);
or U26322 (N_26322,N_21909,N_22093);
xor U26323 (N_26323,N_21756,N_21631);
xor U26324 (N_26324,N_22913,N_22088);
nand U26325 (N_26325,N_22329,N_23215);
nor U26326 (N_26326,N_23613,N_21700);
and U26327 (N_26327,N_23586,N_23765);
and U26328 (N_26328,N_21809,N_21338);
or U26329 (N_26329,N_23265,N_22995);
nor U26330 (N_26330,N_22954,N_23474);
xnor U26331 (N_26331,N_22052,N_23678);
nor U26332 (N_26332,N_21843,N_21244);
and U26333 (N_26333,N_23118,N_22802);
or U26334 (N_26334,N_22561,N_21274);
and U26335 (N_26335,N_21316,N_21788);
xnor U26336 (N_26336,N_21785,N_23827);
or U26337 (N_26337,N_22505,N_22560);
xnor U26338 (N_26338,N_22368,N_22837);
nand U26339 (N_26339,N_23238,N_21971);
or U26340 (N_26340,N_23985,N_23790);
nand U26341 (N_26341,N_22671,N_22790);
xor U26342 (N_26342,N_21224,N_21022);
or U26343 (N_26343,N_22038,N_21237);
xnor U26344 (N_26344,N_21416,N_23453);
nand U26345 (N_26345,N_22936,N_21800);
nand U26346 (N_26346,N_23980,N_21600);
nand U26347 (N_26347,N_22682,N_23385);
or U26348 (N_26348,N_21601,N_21264);
and U26349 (N_26349,N_22548,N_21043);
and U26350 (N_26350,N_22923,N_21142);
or U26351 (N_26351,N_22910,N_22695);
and U26352 (N_26352,N_22434,N_23715);
and U26353 (N_26353,N_22379,N_21366);
nor U26354 (N_26354,N_21322,N_22774);
or U26355 (N_26355,N_22921,N_21550);
nand U26356 (N_26356,N_21545,N_23101);
xnor U26357 (N_26357,N_23072,N_23333);
and U26358 (N_26358,N_23205,N_22138);
or U26359 (N_26359,N_21059,N_21893);
and U26360 (N_26360,N_22464,N_21373);
nor U26361 (N_26361,N_23002,N_21237);
xnor U26362 (N_26362,N_21053,N_22984);
nor U26363 (N_26363,N_22650,N_21318);
xnor U26364 (N_26364,N_21836,N_23445);
xor U26365 (N_26365,N_22469,N_22779);
or U26366 (N_26366,N_21153,N_23987);
xor U26367 (N_26367,N_23996,N_23128);
nand U26368 (N_26368,N_21263,N_21219);
or U26369 (N_26369,N_23684,N_22955);
xor U26370 (N_26370,N_21167,N_21792);
nand U26371 (N_26371,N_23598,N_21663);
xnor U26372 (N_26372,N_23305,N_21637);
nand U26373 (N_26373,N_21224,N_22252);
and U26374 (N_26374,N_22968,N_23910);
and U26375 (N_26375,N_21189,N_23186);
nor U26376 (N_26376,N_23545,N_21466);
nand U26377 (N_26377,N_21851,N_21862);
nand U26378 (N_26378,N_22765,N_22567);
nor U26379 (N_26379,N_23646,N_23890);
and U26380 (N_26380,N_21267,N_22447);
nor U26381 (N_26381,N_22456,N_21343);
nand U26382 (N_26382,N_22921,N_23786);
and U26383 (N_26383,N_21429,N_23635);
xor U26384 (N_26384,N_21816,N_22652);
nand U26385 (N_26385,N_21673,N_22438);
and U26386 (N_26386,N_22957,N_23947);
xor U26387 (N_26387,N_23269,N_21837);
or U26388 (N_26388,N_22080,N_21603);
and U26389 (N_26389,N_21001,N_23296);
nor U26390 (N_26390,N_21826,N_21721);
xnor U26391 (N_26391,N_23790,N_21658);
xor U26392 (N_26392,N_21511,N_21761);
nor U26393 (N_26393,N_23745,N_21161);
and U26394 (N_26394,N_23545,N_21976);
nor U26395 (N_26395,N_21463,N_21260);
xnor U26396 (N_26396,N_23510,N_22156);
xnor U26397 (N_26397,N_21029,N_23068);
and U26398 (N_26398,N_22020,N_22921);
nor U26399 (N_26399,N_23653,N_21131);
xor U26400 (N_26400,N_21809,N_23334);
nand U26401 (N_26401,N_21034,N_23606);
or U26402 (N_26402,N_23245,N_23726);
xor U26403 (N_26403,N_21630,N_23324);
nor U26404 (N_26404,N_23412,N_23270);
nor U26405 (N_26405,N_23558,N_21143);
nor U26406 (N_26406,N_23367,N_23013);
nor U26407 (N_26407,N_22351,N_22209);
and U26408 (N_26408,N_21627,N_21183);
nand U26409 (N_26409,N_22003,N_21456);
or U26410 (N_26410,N_21201,N_23183);
nand U26411 (N_26411,N_23916,N_23771);
and U26412 (N_26412,N_23463,N_22031);
nand U26413 (N_26413,N_23328,N_23115);
and U26414 (N_26414,N_22529,N_21054);
nand U26415 (N_26415,N_21587,N_22564);
nor U26416 (N_26416,N_21082,N_22192);
or U26417 (N_26417,N_23465,N_21759);
or U26418 (N_26418,N_22455,N_23124);
nor U26419 (N_26419,N_21630,N_23239);
nand U26420 (N_26420,N_22051,N_22838);
and U26421 (N_26421,N_23321,N_23966);
xnor U26422 (N_26422,N_23430,N_23115);
and U26423 (N_26423,N_23728,N_21440);
nor U26424 (N_26424,N_21816,N_21476);
nand U26425 (N_26425,N_22446,N_22411);
xor U26426 (N_26426,N_23217,N_22282);
or U26427 (N_26427,N_22456,N_22613);
nor U26428 (N_26428,N_23329,N_21782);
xor U26429 (N_26429,N_22997,N_22206);
or U26430 (N_26430,N_23748,N_22548);
nor U26431 (N_26431,N_23939,N_21415);
xnor U26432 (N_26432,N_21261,N_23098);
xor U26433 (N_26433,N_22110,N_23740);
nand U26434 (N_26434,N_21166,N_23149);
nor U26435 (N_26435,N_21138,N_22496);
nand U26436 (N_26436,N_22122,N_23751);
and U26437 (N_26437,N_22422,N_23739);
xnor U26438 (N_26438,N_21875,N_22010);
nor U26439 (N_26439,N_23488,N_22766);
and U26440 (N_26440,N_22369,N_23349);
nor U26441 (N_26441,N_22727,N_23257);
nand U26442 (N_26442,N_21292,N_23268);
xnor U26443 (N_26443,N_23226,N_23078);
and U26444 (N_26444,N_23836,N_21719);
nand U26445 (N_26445,N_23910,N_21067);
nor U26446 (N_26446,N_22296,N_22859);
or U26447 (N_26447,N_21550,N_22340);
xnor U26448 (N_26448,N_23806,N_22816);
or U26449 (N_26449,N_22266,N_21297);
xor U26450 (N_26450,N_23961,N_23455);
xnor U26451 (N_26451,N_22037,N_23359);
xnor U26452 (N_26452,N_22470,N_22110);
nand U26453 (N_26453,N_23860,N_23159);
xor U26454 (N_26454,N_23661,N_22288);
nor U26455 (N_26455,N_22664,N_21399);
nor U26456 (N_26456,N_23487,N_22983);
nor U26457 (N_26457,N_22868,N_23424);
nand U26458 (N_26458,N_22610,N_23508);
and U26459 (N_26459,N_23752,N_22624);
nand U26460 (N_26460,N_22329,N_22735);
xor U26461 (N_26461,N_21399,N_22996);
and U26462 (N_26462,N_22801,N_22299);
and U26463 (N_26463,N_23339,N_22324);
nor U26464 (N_26464,N_23594,N_21703);
xnor U26465 (N_26465,N_23572,N_21097);
nand U26466 (N_26466,N_23386,N_23059);
nor U26467 (N_26467,N_22067,N_21169);
nor U26468 (N_26468,N_21582,N_22515);
nand U26469 (N_26469,N_23948,N_21150);
and U26470 (N_26470,N_21180,N_23446);
nor U26471 (N_26471,N_21597,N_21734);
xor U26472 (N_26472,N_22769,N_21496);
nand U26473 (N_26473,N_23287,N_21314);
xnor U26474 (N_26474,N_21269,N_21932);
or U26475 (N_26475,N_22989,N_22996);
nor U26476 (N_26476,N_21611,N_21727);
xor U26477 (N_26477,N_23433,N_22822);
nor U26478 (N_26478,N_23806,N_21293);
nand U26479 (N_26479,N_21645,N_21764);
nor U26480 (N_26480,N_21999,N_22477);
or U26481 (N_26481,N_23219,N_21659);
xor U26482 (N_26482,N_23470,N_23756);
and U26483 (N_26483,N_21484,N_23225);
nor U26484 (N_26484,N_21944,N_23121);
and U26485 (N_26485,N_23530,N_22836);
xor U26486 (N_26486,N_23534,N_22383);
nor U26487 (N_26487,N_23812,N_23909);
nand U26488 (N_26488,N_21892,N_22912);
and U26489 (N_26489,N_22560,N_23884);
or U26490 (N_26490,N_21132,N_21775);
or U26491 (N_26491,N_23328,N_22016);
and U26492 (N_26492,N_21552,N_23597);
or U26493 (N_26493,N_23418,N_22974);
xnor U26494 (N_26494,N_23574,N_23525);
nand U26495 (N_26495,N_23262,N_22807);
nand U26496 (N_26496,N_22939,N_23736);
xor U26497 (N_26497,N_22392,N_22987);
nor U26498 (N_26498,N_23988,N_22383);
or U26499 (N_26499,N_21872,N_22357);
or U26500 (N_26500,N_23261,N_23034);
nand U26501 (N_26501,N_22440,N_21099);
or U26502 (N_26502,N_22631,N_23070);
xor U26503 (N_26503,N_21211,N_23894);
xor U26504 (N_26504,N_23491,N_23406);
nand U26505 (N_26505,N_22431,N_22394);
xor U26506 (N_26506,N_23980,N_21840);
xor U26507 (N_26507,N_23704,N_21135);
or U26508 (N_26508,N_23307,N_23918);
and U26509 (N_26509,N_23478,N_21577);
or U26510 (N_26510,N_22572,N_23080);
nand U26511 (N_26511,N_22694,N_23757);
nand U26512 (N_26512,N_22209,N_22998);
or U26513 (N_26513,N_22084,N_23219);
nand U26514 (N_26514,N_23036,N_21442);
or U26515 (N_26515,N_22584,N_21251);
xor U26516 (N_26516,N_21363,N_21759);
and U26517 (N_26517,N_21985,N_21560);
nor U26518 (N_26518,N_22867,N_22631);
or U26519 (N_26519,N_22941,N_23726);
xor U26520 (N_26520,N_23044,N_21622);
or U26521 (N_26521,N_22637,N_23412);
xor U26522 (N_26522,N_21501,N_22843);
xnor U26523 (N_26523,N_22646,N_22698);
or U26524 (N_26524,N_22043,N_23331);
and U26525 (N_26525,N_21807,N_21708);
nand U26526 (N_26526,N_23285,N_22104);
and U26527 (N_26527,N_21018,N_22545);
nor U26528 (N_26528,N_23217,N_21535);
or U26529 (N_26529,N_21922,N_21636);
xnor U26530 (N_26530,N_21116,N_23889);
and U26531 (N_26531,N_23194,N_22295);
nand U26532 (N_26532,N_23650,N_21890);
nor U26533 (N_26533,N_21671,N_21696);
and U26534 (N_26534,N_23410,N_22661);
nand U26535 (N_26535,N_22798,N_22042);
nor U26536 (N_26536,N_21634,N_23123);
nand U26537 (N_26537,N_21360,N_23736);
xor U26538 (N_26538,N_22134,N_21915);
xor U26539 (N_26539,N_22293,N_21162);
xor U26540 (N_26540,N_23073,N_23940);
nor U26541 (N_26541,N_23644,N_22049);
or U26542 (N_26542,N_23320,N_23424);
or U26543 (N_26543,N_22147,N_21211);
or U26544 (N_26544,N_23956,N_22423);
xor U26545 (N_26545,N_22761,N_21395);
xor U26546 (N_26546,N_22267,N_22890);
xnor U26547 (N_26547,N_23959,N_21449);
and U26548 (N_26548,N_21902,N_23417);
nand U26549 (N_26549,N_22059,N_23090);
nor U26550 (N_26550,N_21806,N_23130);
nor U26551 (N_26551,N_22547,N_22652);
or U26552 (N_26552,N_22717,N_23806);
nor U26553 (N_26553,N_23337,N_21083);
or U26554 (N_26554,N_22722,N_21373);
nor U26555 (N_26555,N_21154,N_23342);
nor U26556 (N_26556,N_21456,N_22796);
and U26557 (N_26557,N_21406,N_21014);
nand U26558 (N_26558,N_22548,N_23471);
nand U26559 (N_26559,N_21782,N_21319);
and U26560 (N_26560,N_23446,N_22109);
nor U26561 (N_26561,N_23022,N_22698);
nor U26562 (N_26562,N_22068,N_22377);
nor U26563 (N_26563,N_22912,N_22116);
and U26564 (N_26564,N_22104,N_21069);
nand U26565 (N_26565,N_21865,N_22005);
xor U26566 (N_26566,N_22383,N_21110);
nor U26567 (N_26567,N_23102,N_22228);
or U26568 (N_26568,N_22349,N_21613);
and U26569 (N_26569,N_21162,N_21173);
nand U26570 (N_26570,N_21428,N_22569);
nor U26571 (N_26571,N_23194,N_23477);
or U26572 (N_26572,N_22585,N_23340);
nor U26573 (N_26573,N_21332,N_22408);
xor U26574 (N_26574,N_22670,N_21994);
xor U26575 (N_26575,N_22589,N_23356);
and U26576 (N_26576,N_22545,N_23851);
or U26577 (N_26577,N_21462,N_23852);
and U26578 (N_26578,N_21784,N_22796);
xor U26579 (N_26579,N_23797,N_22984);
nor U26580 (N_26580,N_22356,N_22556);
nor U26581 (N_26581,N_22130,N_21839);
and U26582 (N_26582,N_22982,N_21021);
nor U26583 (N_26583,N_23518,N_21267);
nand U26584 (N_26584,N_22884,N_21428);
and U26585 (N_26585,N_23451,N_22953);
nand U26586 (N_26586,N_21924,N_22078);
xnor U26587 (N_26587,N_22200,N_23037);
nor U26588 (N_26588,N_22378,N_21533);
or U26589 (N_26589,N_22939,N_22678);
and U26590 (N_26590,N_23249,N_21520);
or U26591 (N_26591,N_21793,N_22461);
nor U26592 (N_26592,N_23783,N_23734);
or U26593 (N_26593,N_22322,N_22839);
xor U26594 (N_26594,N_22397,N_22007);
xnor U26595 (N_26595,N_21665,N_22986);
or U26596 (N_26596,N_23026,N_21708);
and U26597 (N_26597,N_21865,N_21110);
and U26598 (N_26598,N_22457,N_23956);
xnor U26599 (N_26599,N_22631,N_22271);
and U26600 (N_26600,N_23580,N_21903);
nand U26601 (N_26601,N_22002,N_22818);
nand U26602 (N_26602,N_21577,N_23174);
xnor U26603 (N_26603,N_22666,N_21591);
and U26604 (N_26604,N_22730,N_21336);
nor U26605 (N_26605,N_23545,N_23020);
xnor U26606 (N_26606,N_22745,N_21016);
xor U26607 (N_26607,N_22091,N_21867);
xnor U26608 (N_26608,N_22412,N_21440);
and U26609 (N_26609,N_22326,N_21058);
or U26610 (N_26610,N_23125,N_21920);
and U26611 (N_26611,N_23519,N_23448);
and U26612 (N_26612,N_22900,N_21875);
nor U26613 (N_26613,N_22336,N_22234);
or U26614 (N_26614,N_23684,N_22845);
nor U26615 (N_26615,N_22692,N_23490);
nand U26616 (N_26616,N_21616,N_22321);
nand U26617 (N_26617,N_22233,N_22046);
and U26618 (N_26618,N_22668,N_22103);
or U26619 (N_26619,N_21352,N_21287);
and U26620 (N_26620,N_21207,N_22735);
xnor U26621 (N_26621,N_22981,N_22536);
nor U26622 (N_26622,N_23776,N_22142);
or U26623 (N_26623,N_23789,N_23811);
xnor U26624 (N_26624,N_22144,N_22365);
and U26625 (N_26625,N_23897,N_21666);
nand U26626 (N_26626,N_23746,N_22541);
and U26627 (N_26627,N_23468,N_21461);
nor U26628 (N_26628,N_21331,N_22906);
xnor U26629 (N_26629,N_22976,N_23129);
or U26630 (N_26630,N_22281,N_21293);
and U26631 (N_26631,N_21207,N_21501);
xor U26632 (N_26632,N_21945,N_23249);
nand U26633 (N_26633,N_21594,N_22633);
and U26634 (N_26634,N_22063,N_23594);
xor U26635 (N_26635,N_22460,N_21384);
or U26636 (N_26636,N_22501,N_22293);
or U26637 (N_26637,N_21151,N_22250);
xor U26638 (N_26638,N_21508,N_21091);
or U26639 (N_26639,N_22148,N_22544);
nor U26640 (N_26640,N_21187,N_22517);
xor U26641 (N_26641,N_22350,N_21762);
or U26642 (N_26642,N_23975,N_22786);
xor U26643 (N_26643,N_22153,N_22531);
nor U26644 (N_26644,N_22472,N_23047);
or U26645 (N_26645,N_22587,N_21756);
nand U26646 (N_26646,N_22155,N_21161);
xnor U26647 (N_26647,N_21813,N_22004);
or U26648 (N_26648,N_21693,N_23664);
or U26649 (N_26649,N_22525,N_22043);
or U26650 (N_26650,N_21256,N_21153);
and U26651 (N_26651,N_22673,N_21043);
xnor U26652 (N_26652,N_22640,N_22222);
and U26653 (N_26653,N_21621,N_22056);
xnor U26654 (N_26654,N_21934,N_21340);
and U26655 (N_26655,N_21144,N_21015);
or U26656 (N_26656,N_22392,N_23253);
nand U26657 (N_26657,N_22671,N_22410);
and U26658 (N_26658,N_22032,N_22533);
nand U26659 (N_26659,N_21217,N_23164);
and U26660 (N_26660,N_22056,N_23191);
or U26661 (N_26661,N_23246,N_22787);
or U26662 (N_26662,N_21059,N_23852);
nor U26663 (N_26663,N_23925,N_23276);
xor U26664 (N_26664,N_22066,N_22111);
and U26665 (N_26665,N_22877,N_21086);
nor U26666 (N_26666,N_21522,N_22493);
nor U26667 (N_26667,N_23098,N_23253);
nand U26668 (N_26668,N_22511,N_22611);
nor U26669 (N_26669,N_23479,N_23572);
nor U26670 (N_26670,N_23147,N_23991);
nor U26671 (N_26671,N_23776,N_23964);
or U26672 (N_26672,N_21596,N_21223);
and U26673 (N_26673,N_23907,N_23115);
nor U26674 (N_26674,N_22858,N_22658);
xnor U26675 (N_26675,N_23184,N_22706);
or U26676 (N_26676,N_23530,N_21766);
or U26677 (N_26677,N_21530,N_21397);
and U26678 (N_26678,N_21915,N_23355);
xor U26679 (N_26679,N_21607,N_22893);
or U26680 (N_26680,N_21216,N_23971);
nand U26681 (N_26681,N_21300,N_22498);
and U26682 (N_26682,N_21626,N_23687);
xor U26683 (N_26683,N_23849,N_23206);
nor U26684 (N_26684,N_21697,N_22742);
xnor U26685 (N_26685,N_23778,N_23945);
nor U26686 (N_26686,N_23307,N_21893);
nand U26687 (N_26687,N_21834,N_21744);
or U26688 (N_26688,N_23486,N_22586);
nand U26689 (N_26689,N_22300,N_23229);
nand U26690 (N_26690,N_21713,N_23878);
and U26691 (N_26691,N_22065,N_21068);
nor U26692 (N_26692,N_23398,N_23183);
nor U26693 (N_26693,N_23885,N_23533);
and U26694 (N_26694,N_23470,N_23894);
and U26695 (N_26695,N_23842,N_21195);
nand U26696 (N_26696,N_23999,N_23886);
nand U26697 (N_26697,N_22334,N_21208);
nor U26698 (N_26698,N_23334,N_23126);
and U26699 (N_26699,N_23768,N_22078);
nand U26700 (N_26700,N_21529,N_21861);
or U26701 (N_26701,N_23701,N_21054);
or U26702 (N_26702,N_23234,N_22160);
nand U26703 (N_26703,N_22385,N_22037);
xor U26704 (N_26704,N_21452,N_23665);
nand U26705 (N_26705,N_21441,N_22336);
nand U26706 (N_26706,N_21558,N_23913);
xor U26707 (N_26707,N_22291,N_22987);
nor U26708 (N_26708,N_23885,N_22354);
or U26709 (N_26709,N_21004,N_21508);
xor U26710 (N_26710,N_22162,N_21415);
or U26711 (N_26711,N_21675,N_22608);
and U26712 (N_26712,N_22372,N_23995);
xor U26713 (N_26713,N_22659,N_21222);
nor U26714 (N_26714,N_23887,N_21426);
xnor U26715 (N_26715,N_21094,N_22985);
xnor U26716 (N_26716,N_22752,N_22611);
xnor U26717 (N_26717,N_21502,N_23256);
xnor U26718 (N_26718,N_22711,N_22781);
and U26719 (N_26719,N_23478,N_21626);
xnor U26720 (N_26720,N_22584,N_23409);
xnor U26721 (N_26721,N_22014,N_22026);
or U26722 (N_26722,N_22349,N_22049);
xor U26723 (N_26723,N_21925,N_21905);
or U26724 (N_26724,N_21149,N_21225);
xor U26725 (N_26725,N_21543,N_23192);
xnor U26726 (N_26726,N_21547,N_23540);
nand U26727 (N_26727,N_21130,N_23405);
nand U26728 (N_26728,N_23042,N_23108);
or U26729 (N_26729,N_22705,N_22804);
and U26730 (N_26730,N_21867,N_21591);
and U26731 (N_26731,N_22588,N_22742);
nor U26732 (N_26732,N_22753,N_21634);
or U26733 (N_26733,N_23768,N_23884);
and U26734 (N_26734,N_23689,N_21289);
nand U26735 (N_26735,N_21314,N_23527);
nor U26736 (N_26736,N_22324,N_21922);
or U26737 (N_26737,N_23491,N_22937);
or U26738 (N_26738,N_21014,N_22432);
and U26739 (N_26739,N_22345,N_21975);
xnor U26740 (N_26740,N_21150,N_22708);
nand U26741 (N_26741,N_21745,N_22907);
nor U26742 (N_26742,N_21540,N_22340);
xnor U26743 (N_26743,N_22387,N_23254);
nand U26744 (N_26744,N_21854,N_23340);
and U26745 (N_26745,N_21312,N_22335);
or U26746 (N_26746,N_23900,N_23472);
xor U26747 (N_26747,N_22339,N_21622);
and U26748 (N_26748,N_23718,N_21951);
and U26749 (N_26749,N_22491,N_22042);
nor U26750 (N_26750,N_21506,N_23430);
and U26751 (N_26751,N_23700,N_22473);
and U26752 (N_26752,N_21862,N_22460);
or U26753 (N_26753,N_22589,N_21450);
or U26754 (N_26754,N_22967,N_21163);
and U26755 (N_26755,N_22852,N_23055);
nand U26756 (N_26756,N_21977,N_23210);
or U26757 (N_26757,N_21305,N_22471);
nand U26758 (N_26758,N_23034,N_23326);
nor U26759 (N_26759,N_22799,N_22913);
and U26760 (N_26760,N_21620,N_23228);
and U26761 (N_26761,N_21528,N_23076);
xor U26762 (N_26762,N_22955,N_22523);
nor U26763 (N_26763,N_23459,N_23716);
and U26764 (N_26764,N_21121,N_21947);
and U26765 (N_26765,N_23911,N_23145);
xor U26766 (N_26766,N_21688,N_23092);
xor U26767 (N_26767,N_22981,N_22637);
nor U26768 (N_26768,N_23159,N_23366);
and U26769 (N_26769,N_23852,N_21549);
or U26770 (N_26770,N_22171,N_22362);
and U26771 (N_26771,N_22653,N_21896);
nor U26772 (N_26772,N_23805,N_22968);
nor U26773 (N_26773,N_23678,N_22282);
and U26774 (N_26774,N_23329,N_22575);
and U26775 (N_26775,N_22780,N_22209);
nand U26776 (N_26776,N_22459,N_21880);
nand U26777 (N_26777,N_21933,N_21604);
and U26778 (N_26778,N_22698,N_22248);
nor U26779 (N_26779,N_22666,N_21115);
and U26780 (N_26780,N_22840,N_22005);
nand U26781 (N_26781,N_22079,N_23013);
nor U26782 (N_26782,N_21864,N_21992);
and U26783 (N_26783,N_23654,N_23605);
and U26784 (N_26784,N_22338,N_22726);
nor U26785 (N_26785,N_21641,N_23359);
xnor U26786 (N_26786,N_23298,N_21282);
and U26787 (N_26787,N_22874,N_21467);
or U26788 (N_26788,N_23474,N_22958);
nand U26789 (N_26789,N_22519,N_23365);
xnor U26790 (N_26790,N_21710,N_21455);
nor U26791 (N_26791,N_22704,N_22450);
nand U26792 (N_26792,N_21713,N_21073);
nand U26793 (N_26793,N_23041,N_22490);
nor U26794 (N_26794,N_22261,N_23694);
or U26795 (N_26795,N_21961,N_22283);
nor U26796 (N_26796,N_22531,N_23681);
nand U26797 (N_26797,N_23611,N_23957);
nor U26798 (N_26798,N_22064,N_22015);
and U26799 (N_26799,N_22330,N_23415);
nor U26800 (N_26800,N_23495,N_22082);
and U26801 (N_26801,N_23665,N_22691);
nand U26802 (N_26802,N_21559,N_22468);
nand U26803 (N_26803,N_22500,N_22489);
nor U26804 (N_26804,N_22479,N_23014);
and U26805 (N_26805,N_23108,N_23591);
nand U26806 (N_26806,N_21432,N_21182);
nand U26807 (N_26807,N_23514,N_23942);
nand U26808 (N_26808,N_22304,N_21756);
nor U26809 (N_26809,N_21207,N_21675);
xnor U26810 (N_26810,N_23238,N_22652);
nor U26811 (N_26811,N_21156,N_21792);
nor U26812 (N_26812,N_22324,N_22004);
and U26813 (N_26813,N_22072,N_23650);
or U26814 (N_26814,N_21226,N_23186);
or U26815 (N_26815,N_23595,N_21674);
nor U26816 (N_26816,N_21297,N_21415);
and U26817 (N_26817,N_22166,N_23539);
xnor U26818 (N_26818,N_23470,N_22477);
nor U26819 (N_26819,N_21346,N_22102);
nand U26820 (N_26820,N_23835,N_23721);
nand U26821 (N_26821,N_22618,N_23428);
nand U26822 (N_26822,N_22629,N_23601);
and U26823 (N_26823,N_22304,N_23391);
and U26824 (N_26824,N_22203,N_23124);
and U26825 (N_26825,N_22031,N_21518);
nand U26826 (N_26826,N_22697,N_22230);
and U26827 (N_26827,N_21317,N_23614);
xnor U26828 (N_26828,N_22422,N_22776);
nor U26829 (N_26829,N_23332,N_23905);
xnor U26830 (N_26830,N_23806,N_22832);
nand U26831 (N_26831,N_21530,N_23553);
or U26832 (N_26832,N_23563,N_22254);
xor U26833 (N_26833,N_22644,N_21152);
nor U26834 (N_26834,N_23598,N_23208);
nor U26835 (N_26835,N_23533,N_23214);
nor U26836 (N_26836,N_21995,N_22361);
xnor U26837 (N_26837,N_23508,N_23269);
or U26838 (N_26838,N_22530,N_22293);
and U26839 (N_26839,N_23784,N_21981);
xor U26840 (N_26840,N_22377,N_23634);
xnor U26841 (N_26841,N_21075,N_22626);
xnor U26842 (N_26842,N_21156,N_21447);
or U26843 (N_26843,N_22505,N_23796);
xor U26844 (N_26844,N_23553,N_22077);
or U26845 (N_26845,N_23231,N_22302);
nor U26846 (N_26846,N_21397,N_21111);
xor U26847 (N_26847,N_22348,N_23988);
nor U26848 (N_26848,N_23737,N_22366);
or U26849 (N_26849,N_22471,N_21207);
and U26850 (N_26850,N_23378,N_22648);
nor U26851 (N_26851,N_22899,N_21939);
nand U26852 (N_26852,N_23655,N_23051);
and U26853 (N_26853,N_21251,N_23647);
nor U26854 (N_26854,N_23817,N_21272);
or U26855 (N_26855,N_23595,N_23546);
xnor U26856 (N_26856,N_22280,N_21463);
or U26857 (N_26857,N_22917,N_23753);
and U26858 (N_26858,N_21048,N_21927);
or U26859 (N_26859,N_23821,N_22340);
and U26860 (N_26860,N_21053,N_23802);
and U26861 (N_26861,N_22044,N_23067);
or U26862 (N_26862,N_23124,N_21833);
nor U26863 (N_26863,N_22479,N_22954);
xor U26864 (N_26864,N_23245,N_21144);
nor U26865 (N_26865,N_21680,N_22561);
and U26866 (N_26866,N_21064,N_23122);
xnor U26867 (N_26867,N_22156,N_21152);
nor U26868 (N_26868,N_21385,N_23762);
or U26869 (N_26869,N_21486,N_22285);
nor U26870 (N_26870,N_22109,N_22639);
and U26871 (N_26871,N_21313,N_23200);
nor U26872 (N_26872,N_22571,N_23254);
xnor U26873 (N_26873,N_21020,N_21431);
or U26874 (N_26874,N_22597,N_22252);
xor U26875 (N_26875,N_22752,N_22614);
xor U26876 (N_26876,N_21538,N_21345);
or U26877 (N_26877,N_21995,N_21777);
or U26878 (N_26878,N_23362,N_22770);
nand U26879 (N_26879,N_22452,N_21397);
nand U26880 (N_26880,N_21585,N_22997);
xor U26881 (N_26881,N_22484,N_23954);
and U26882 (N_26882,N_21872,N_21790);
nand U26883 (N_26883,N_21456,N_22490);
or U26884 (N_26884,N_22140,N_23823);
xnor U26885 (N_26885,N_23183,N_21232);
or U26886 (N_26886,N_23943,N_21955);
or U26887 (N_26887,N_23792,N_21139);
xnor U26888 (N_26888,N_22804,N_21715);
and U26889 (N_26889,N_22519,N_23978);
or U26890 (N_26890,N_22212,N_21397);
or U26891 (N_26891,N_23998,N_23096);
nand U26892 (N_26892,N_23427,N_21557);
xnor U26893 (N_26893,N_23017,N_23982);
nand U26894 (N_26894,N_23776,N_21081);
and U26895 (N_26895,N_21184,N_21422);
or U26896 (N_26896,N_23388,N_21735);
or U26897 (N_26897,N_23723,N_22798);
xor U26898 (N_26898,N_23663,N_23456);
and U26899 (N_26899,N_22181,N_22080);
or U26900 (N_26900,N_21345,N_21200);
xnor U26901 (N_26901,N_21915,N_21443);
nor U26902 (N_26902,N_23650,N_21134);
nor U26903 (N_26903,N_22235,N_23756);
nor U26904 (N_26904,N_21513,N_23456);
nor U26905 (N_26905,N_23100,N_23720);
or U26906 (N_26906,N_23254,N_22158);
nand U26907 (N_26907,N_21097,N_23249);
xnor U26908 (N_26908,N_23273,N_23508);
and U26909 (N_26909,N_22984,N_22072);
nor U26910 (N_26910,N_22873,N_23216);
or U26911 (N_26911,N_22786,N_22967);
xnor U26912 (N_26912,N_23314,N_21705);
and U26913 (N_26913,N_22938,N_21348);
xor U26914 (N_26914,N_21634,N_23948);
and U26915 (N_26915,N_21513,N_22240);
and U26916 (N_26916,N_23837,N_23608);
and U26917 (N_26917,N_21587,N_23846);
nor U26918 (N_26918,N_23617,N_21295);
and U26919 (N_26919,N_23444,N_21937);
and U26920 (N_26920,N_23610,N_23195);
or U26921 (N_26921,N_21381,N_21525);
xnor U26922 (N_26922,N_21233,N_21486);
nor U26923 (N_26923,N_22601,N_21760);
nand U26924 (N_26924,N_21781,N_23031);
xnor U26925 (N_26925,N_23507,N_21270);
nor U26926 (N_26926,N_22315,N_21942);
or U26927 (N_26927,N_23328,N_23252);
nor U26928 (N_26928,N_21145,N_23899);
nand U26929 (N_26929,N_23273,N_21241);
xor U26930 (N_26930,N_21345,N_23549);
or U26931 (N_26931,N_21657,N_22011);
nand U26932 (N_26932,N_21949,N_21541);
nor U26933 (N_26933,N_21784,N_22730);
nand U26934 (N_26934,N_21396,N_21473);
nand U26935 (N_26935,N_22469,N_21395);
nand U26936 (N_26936,N_21274,N_23028);
and U26937 (N_26937,N_21232,N_23708);
or U26938 (N_26938,N_21322,N_23761);
or U26939 (N_26939,N_21315,N_23537);
xor U26940 (N_26940,N_22866,N_21355);
nor U26941 (N_26941,N_23731,N_23697);
or U26942 (N_26942,N_21598,N_21253);
nor U26943 (N_26943,N_23216,N_23401);
nor U26944 (N_26944,N_21538,N_21258);
and U26945 (N_26945,N_22053,N_23855);
or U26946 (N_26946,N_22627,N_22490);
nand U26947 (N_26947,N_23949,N_22673);
xnor U26948 (N_26948,N_21651,N_22156);
or U26949 (N_26949,N_21954,N_23252);
or U26950 (N_26950,N_23131,N_22409);
and U26951 (N_26951,N_22292,N_21726);
and U26952 (N_26952,N_21026,N_23100);
nor U26953 (N_26953,N_23499,N_23566);
and U26954 (N_26954,N_22789,N_21708);
nand U26955 (N_26955,N_23438,N_22294);
nand U26956 (N_26956,N_23495,N_21180);
and U26957 (N_26957,N_22057,N_22967);
nor U26958 (N_26958,N_22086,N_21105);
and U26959 (N_26959,N_21930,N_21017);
or U26960 (N_26960,N_23188,N_21373);
or U26961 (N_26961,N_22680,N_21647);
and U26962 (N_26962,N_21890,N_23689);
or U26963 (N_26963,N_21797,N_21791);
and U26964 (N_26964,N_23238,N_21069);
nand U26965 (N_26965,N_21285,N_23017);
nand U26966 (N_26966,N_21307,N_23424);
nand U26967 (N_26967,N_23270,N_22875);
and U26968 (N_26968,N_22183,N_23022);
and U26969 (N_26969,N_21965,N_21474);
or U26970 (N_26970,N_21513,N_23103);
xnor U26971 (N_26971,N_22887,N_22835);
nand U26972 (N_26972,N_21186,N_22945);
and U26973 (N_26973,N_22920,N_23556);
xnor U26974 (N_26974,N_23565,N_23954);
xor U26975 (N_26975,N_23102,N_22609);
or U26976 (N_26976,N_21962,N_23833);
and U26977 (N_26977,N_22310,N_22703);
xor U26978 (N_26978,N_21824,N_22894);
nand U26979 (N_26979,N_22970,N_22574);
nand U26980 (N_26980,N_23784,N_21241);
or U26981 (N_26981,N_21061,N_22266);
nand U26982 (N_26982,N_23170,N_22916);
nand U26983 (N_26983,N_23872,N_23561);
and U26984 (N_26984,N_23790,N_22954);
and U26985 (N_26985,N_21239,N_21145);
and U26986 (N_26986,N_23381,N_22965);
nand U26987 (N_26987,N_22478,N_22654);
and U26988 (N_26988,N_21768,N_22372);
or U26989 (N_26989,N_23153,N_23020);
and U26990 (N_26990,N_23113,N_21691);
and U26991 (N_26991,N_22092,N_21010);
nor U26992 (N_26992,N_22300,N_23992);
nor U26993 (N_26993,N_22465,N_23622);
and U26994 (N_26994,N_23340,N_21864);
and U26995 (N_26995,N_23611,N_21068);
nor U26996 (N_26996,N_22802,N_21224);
and U26997 (N_26997,N_22888,N_21688);
nor U26998 (N_26998,N_21553,N_21804);
xnor U26999 (N_26999,N_22469,N_21479);
nand U27000 (N_27000,N_25824,N_24703);
nor U27001 (N_27001,N_25938,N_25095);
and U27002 (N_27002,N_26249,N_24952);
xor U27003 (N_27003,N_25925,N_24058);
or U27004 (N_27004,N_24579,N_25948);
nor U27005 (N_27005,N_24720,N_26415);
nor U27006 (N_27006,N_24965,N_24646);
xor U27007 (N_27007,N_26259,N_25662);
or U27008 (N_27008,N_25754,N_26204);
nor U27009 (N_27009,N_26084,N_24786);
nand U27010 (N_27010,N_26920,N_25955);
nand U27011 (N_27011,N_25335,N_25597);
or U27012 (N_27012,N_25803,N_24233);
nand U27013 (N_27013,N_24298,N_25959);
xor U27014 (N_27014,N_26975,N_25254);
xnor U27015 (N_27015,N_24966,N_24679);
nor U27016 (N_27016,N_26927,N_24582);
nand U27017 (N_27017,N_26760,N_24062);
xor U27018 (N_27018,N_25999,N_24235);
nand U27019 (N_27019,N_25247,N_24307);
nand U27020 (N_27020,N_25638,N_25892);
xor U27021 (N_27021,N_26307,N_25550);
and U27022 (N_27022,N_25471,N_24516);
or U27023 (N_27023,N_26248,N_24749);
xor U27024 (N_27024,N_24261,N_26352);
and U27025 (N_27025,N_24434,N_26202);
nand U27026 (N_27026,N_26147,N_26491);
nor U27027 (N_27027,N_25812,N_26325);
xor U27028 (N_27028,N_26376,N_24179);
nand U27029 (N_27029,N_25272,N_26501);
nor U27030 (N_27030,N_24659,N_25120);
nand U27031 (N_27031,N_25053,N_25267);
nand U27032 (N_27032,N_25571,N_25210);
nand U27033 (N_27033,N_26126,N_25664);
xnor U27034 (N_27034,N_24685,N_25054);
and U27035 (N_27035,N_25307,N_24736);
nand U27036 (N_27036,N_24610,N_25167);
and U27037 (N_27037,N_25286,N_24936);
or U27038 (N_27038,N_24573,N_24551);
and U27039 (N_27039,N_24077,N_24841);
nand U27040 (N_27040,N_24008,N_26161);
nand U27041 (N_27041,N_26590,N_24539);
nor U27042 (N_27042,N_26324,N_26390);
nand U27043 (N_27043,N_26203,N_24323);
or U27044 (N_27044,N_25699,N_24276);
and U27045 (N_27045,N_25215,N_26518);
and U27046 (N_27046,N_24324,N_24175);
nor U27047 (N_27047,N_24207,N_25278);
nor U27048 (N_27048,N_26093,N_26574);
nor U27049 (N_27049,N_24466,N_26237);
or U27050 (N_27050,N_24110,N_26326);
nand U27051 (N_27051,N_25381,N_25972);
nor U27052 (N_27052,N_26672,N_24524);
and U27053 (N_27053,N_24231,N_25728);
xor U27054 (N_27054,N_25726,N_24648);
nor U27055 (N_27055,N_24721,N_24758);
and U27056 (N_27056,N_24407,N_24433);
or U27057 (N_27057,N_25020,N_26253);
xor U27058 (N_27058,N_25069,N_26659);
nand U27059 (N_27059,N_26452,N_26860);
nand U27060 (N_27060,N_25917,N_26804);
nand U27061 (N_27061,N_25178,N_25640);
and U27062 (N_27062,N_25332,N_26757);
and U27063 (N_27063,N_25601,N_25637);
nor U27064 (N_27064,N_26532,N_25139);
nor U27065 (N_27065,N_25371,N_25880);
and U27066 (N_27066,N_24205,N_25829);
or U27067 (N_27067,N_26981,N_25872);
or U27068 (N_27068,N_26886,N_26377);
nor U27069 (N_27069,N_26740,N_26961);
and U27070 (N_27070,N_25791,N_26064);
xor U27071 (N_27071,N_26081,N_24288);
xnor U27072 (N_27072,N_24894,N_25870);
nand U27073 (N_27073,N_26615,N_24701);
nor U27074 (N_27074,N_26314,N_24764);
and U27075 (N_27075,N_26152,N_25559);
xnor U27076 (N_27076,N_25137,N_25249);
and U27077 (N_27077,N_24742,N_24732);
and U27078 (N_27078,N_24018,N_25469);
nand U27079 (N_27079,N_24413,N_26617);
or U27080 (N_27080,N_24396,N_24939);
nand U27081 (N_27081,N_25374,N_26030);
xor U27082 (N_27082,N_24373,N_26356);
and U27083 (N_27083,N_25626,N_24193);
xnor U27084 (N_27084,N_26512,N_24740);
nand U27085 (N_27085,N_26543,N_26427);
nand U27086 (N_27086,N_25441,N_24994);
xnor U27087 (N_27087,N_26934,N_26255);
nand U27088 (N_27088,N_24349,N_26669);
and U27089 (N_27089,N_25825,N_24509);
nor U27090 (N_27090,N_25881,N_24174);
xor U27091 (N_27091,N_26406,N_24831);
and U27092 (N_27092,N_26507,N_25453);
nor U27093 (N_27093,N_25182,N_24791);
nor U27094 (N_27094,N_26190,N_25067);
xor U27095 (N_27095,N_26137,N_26162);
xnor U27096 (N_27096,N_25265,N_26799);
xnor U27097 (N_27097,N_25416,N_26751);
nand U27098 (N_27098,N_25670,N_25544);
xnor U27099 (N_27099,N_25352,N_26720);
or U27100 (N_27100,N_25276,N_26213);
xor U27101 (N_27101,N_25147,N_26422);
nand U27102 (N_27102,N_26301,N_26242);
xor U27103 (N_27103,N_24618,N_25867);
nand U27104 (N_27104,N_24441,N_25968);
xor U27105 (N_27105,N_24541,N_24596);
and U27106 (N_27106,N_26527,N_24617);
and U27107 (N_27107,N_25903,N_24086);
nand U27108 (N_27108,N_24908,N_26509);
nand U27109 (N_27109,N_24655,N_24960);
or U27110 (N_27110,N_24003,N_26941);
nand U27111 (N_27111,N_24989,N_25848);
xor U27112 (N_27112,N_24036,N_26191);
nand U27113 (N_27113,N_25906,N_25214);
and U27114 (N_27114,N_25168,N_24023);
and U27115 (N_27115,N_26401,N_26002);
or U27116 (N_27116,N_26447,N_25011);
and U27117 (N_27117,N_25992,N_24107);
or U27118 (N_27118,N_24739,N_24801);
or U27119 (N_27119,N_24904,N_25465);
and U27120 (N_27120,N_24126,N_24605);
xnor U27121 (N_27121,N_25455,N_25016);
xnor U27122 (N_27122,N_25783,N_25749);
nor U27123 (N_27123,N_24654,N_25582);
nor U27124 (N_27124,N_24247,N_25108);
nor U27125 (N_27125,N_24998,N_25945);
nand U27126 (N_27126,N_26776,N_26115);
xnor U27127 (N_27127,N_25190,N_26613);
xor U27128 (N_27128,N_25826,N_26304);
or U27129 (N_27129,N_26297,N_24977);
nand U27130 (N_27130,N_26652,N_26550);
xor U27131 (N_27131,N_26537,N_24280);
xor U27132 (N_27132,N_24395,N_25440);
xnor U27133 (N_27133,N_25962,N_26719);
and U27134 (N_27134,N_25390,N_25226);
or U27135 (N_27135,N_24306,N_24465);
nor U27136 (N_27136,N_26344,N_25394);
nor U27137 (N_27137,N_24978,N_26027);
nor U27138 (N_27138,N_26578,N_26750);
xor U27139 (N_27139,N_24278,N_25415);
xor U27140 (N_27140,N_24526,N_24845);
or U27141 (N_27141,N_24528,N_26591);
xor U27142 (N_27142,N_26756,N_25162);
nor U27143 (N_27143,N_26627,N_26494);
and U27144 (N_27144,N_25532,N_26890);
and U27145 (N_27145,N_26705,N_25346);
xnor U27146 (N_27146,N_24025,N_24042);
or U27147 (N_27147,N_24871,N_24419);
xor U27148 (N_27148,N_26303,N_24300);
xnor U27149 (N_27149,N_24302,N_25409);
or U27150 (N_27150,N_24265,N_24729);
and U27151 (N_27151,N_25629,N_26646);
and U27152 (N_27152,N_24249,N_24702);
nor U27153 (N_27153,N_25093,N_26783);
nor U27154 (N_27154,N_24151,N_26539);
nand U27155 (N_27155,N_25688,N_24420);
nor U27156 (N_27156,N_26817,N_25882);
or U27157 (N_27157,N_26038,N_24669);
nor U27158 (N_27158,N_26440,N_24435);
and U27159 (N_27159,N_26536,N_24052);
and U27160 (N_27160,N_24754,N_26108);
nand U27161 (N_27161,N_26540,N_24012);
nor U27162 (N_27162,N_25943,N_24398);
and U27163 (N_27163,N_25443,N_24511);
xnor U27164 (N_27164,N_24422,N_25654);
or U27165 (N_27165,N_24044,N_25540);
or U27166 (N_27166,N_24519,N_25492);
and U27167 (N_27167,N_25539,N_25007);
nand U27168 (N_27168,N_25036,N_26694);
nand U27169 (N_27169,N_24309,N_25823);
nand U27170 (N_27170,N_26748,N_24860);
and U27171 (N_27171,N_26319,N_25133);
nand U27172 (N_27172,N_26355,N_26071);
and U27173 (N_27173,N_25623,N_25169);
nand U27174 (N_27174,N_26604,N_24079);
nand U27175 (N_27175,N_24337,N_26306);
xor U27176 (N_27176,N_26291,N_25865);
and U27177 (N_27177,N_26809,N_25555);
xnor U27178 (N_27178,N_25407,N_26962);
nor U27179 (N_27179,N_25336,N_26565);
or U27180 (N_27180,N_24499,N_26272);
and U27181 (N_27181,N_25197,N_26519);
xnor U27182 (N_27182,N_24687,N_26883);
and U27183 (N_27183,N_24218,N_24898);
nand U27184 (N_27184,N_24345,N_24899);
and U27185 (N_27185,N_25103,N_25625);
and U27186 (N_27186,N_26568,N_25362);
xor U27187 (N_27187,N_24271,N_26025);
xor U27188 (N_27188,N_25996,N_25705);
nor U27189 (N_27189,N_24827,N_25836);
or U27190 (N_27190,N_24514,N_26090);
nand U27191 (N_27191,N_25546,N_26774);
nand U27192 (N_27192,N_24240,N_26786);
nor U27193 (N_27193,N_24990,N_25293);
or U27194 (N_27194,N_25126,N_24521);
and U27195 (N_27195,N_26921,N_26978);
nand U27196 (N_27196,N_26982,N_26881);
or U27197 (N_27197,N_26160,N_26368);
nor U27198 (N_27198,N_25909,N_26770);
or U27199 (N_27199,N_25157,N_24672);
xor U27200 (N_27200,N_24201,N_24838);
or U27201 (N_27201,N_26983,N_24048);
nand U27202 (N_27202,N_25551,N_26431);
nor U27203 (N_27203,N_26577,N_25375);
nand U27204 (N_27204,N_24730,N_26647);
and U27205 (N_27205,N_26214,N_24070);
or U27206 (N_27206,N_26937,N_24093);
and U27207 (N_27207,N_24105,N_26096);
xor U27208 (N_27208,N_24628,N_25835);
and U27209 (N_27209,N_26369,N_25413);
nand U27210 (N_27210,N_24725,N_26693);
nor U27211 (N_27211,N_26278,N_25482);
or U27212 (N_27212,N_26793,N_26383);
nand U27213 (N_27213,N_26360,N_24762);
nor U27214 (N_27214,N_26648,N_24131);
and U27215 (N_27215,N_25635,N_24212);
nor U27216 (N_27216,N_24559,N_26818);
and U27217 (N_27217,N_25149,N_25518);
and U27218 (N_27218,N_25119,N_25475);
nand U27219 (N_27219,N_24316,N_26286);
xor U27220 (N_27220,N_25869,N_25758);
and U27221 (N_27221,N_24456,N_24745);
nor U27222 (N_27222,N_24092,N_25245);
nand U27223 (N_27223,N_25639,N_24439);
nor U27224 (N_27224,N_26544,N_25195);
and U27225 (N_27225,N_24892,N_25048);
nand U27226 (N_27226,N_26347,N_24080);
and U27227 (N_27227,N_26097,N_24180);
nor U27228 (N_27228,N_24158,N_26396);
nand U27229 (N_27229,N_25176,N_24747);
nor U27230 (N_27230,N_25402,N_24479);
nand U27231 (N_27231,N_24492,N_24774);
nand U27232 (N_27232,N_26337,N_25766);
or U27233 (N_27233,N_25599,N_25656);
or U27234 (N_27234,N_25859,N_25275);
nor U27235 (N_27235,N_25682,N_24252);
or U27236 (N_27236,N_24597,N_24505);
or U27237 (N_27237,N_24792,N_24026);
xnor U27238 (N_27238,N_26063,N_24947);
nor U27239 (N_27239,N_25460,N_25291);
nor U27240 (N_27240,N_24870,N_25813);
and U27241 (N_27241,N_26479,N_24517);
nor U27242 (N_27242,N_26414,N_25260);
xnor U27243 (N_27243,N_24440,N_24621);
xor U27244 (N_27244,N_24583,N_26183);
xor U27245 (N_27245,N_24763,N_25023);
xnor U27246 (N_27246,N_24431,N_26623);
or U27247 (N_27247,N_26877,N_24810);
nand U27248 (N_27248,N_25145,N_24882);
or U27249 (N_27249,N_24748,N_26492);
or U27250 (N_27250,N_25521,N_26432);
xor U27251 (N_27251,N_24384,N_25185);
nor U27252 (N_27252,N_26503,N_26022);
nand U27253 (N_27253,N_24983,N_26716);
and U27254 (N_27254,N_24301,N_24377);
and U27255 (N_27255,N_25724,N_24735);
nand U27256 (N_27256,N_24075,N_25083);
or U27257 (N_27257,N_24194,N_25568);
xnor U27258 (N_27258,N_26239,N_25595);
nor U27259 (N_27259,N_24906,N_26234);
nand U27260 (N_27260,N_25944,N_26245);
or U27261 (N_27261,N_24255,N_25557);
xor U27262 (N_27262,N_24177,N_24447);
nor U27263 (N_27263,N_25498,N_26007);
xor U27264 (N_27264,N_25849,N_25367);
nor U27265 (N_27265,N_26892,N_25014);
xor U27266 (N_27266,N_26382,N_25747);
or U27267 (N_27267,N_24046,N_26262);
and U27268 (N_27268,N_24136,N_24397);
xnor U27269 (N_27269,N_24826,N_26661);
xnor U27270 (N_27270,N_26820,N_26634);
and U27271 (N_27271,N_25043,N_24344);
nor U27272 (N_27272,N_25030,N_25129);
and U27273 (N_27273,N_26714,N_25364);
nor U27274 (N_27274,N_24608,N_25667);
and U27275 (N_27275,N_26362,N_25932);
nor U27276 (N_27276,N_24051,N_26821);
xnor U27277 (N_27277,N_26515,N_26510);
or U27278 (N_27278,N_24881,N_26562);
and U27279 (N_27279,N_25243,N_24173);
xnor U27280 (N_27280,N_26233,N_24495);
nor U27281 (N_27281,N_26739,N_26749);
or U27282 (N_27282,N_26640,N_24626);
nand U27283 (N_27283,N_26708,N_24032);
or U27284 (N_27284,N_25894,N_24449);
and U27285 (N_27285,N_24925,N_26736);
nor U27286 (N_27286,N_26588,N_25039);
nor U27287 (N_27287,N_25833,N_24733);
or U27288 (N_27288,N_24340,N_26358);
or U27289 (N_27289,N_25353,N_24015);
and U27290 (N_27290,N_25918,N_26206);
or U27291 (N_27291,N_26080,N_25154);
nor U27292 (N_27292,N_25049,N_24753);
nor U27293 (N_27293,N_24320,N_25001);
nand U27294 (N_27294,N_24497,N_24922);
xor U27295 (N_27295,N_25669,N_25850);
or U27296 (N_27296,N_24338,N_26192);
and U27297 (N_27297,N_24006,N_26989);
nand U27298 (N_27298,N_25148,N_25731);
nor U27299 (N_27299,N_25319,N_25960);
or U27300 (N_27300,N_25564,N_26200);
nor U27301 (N_27301,N_24141,N_24816);
nand U27302 (N_27302,N_26318,N_24043);
or U27303 (N_27303,N_26970,N_24727);
and U27304 (N_27304,N_24888,N_24601);
or U27305 (N_27305,N_26472,N_26180);
xor U27306 (N_27306,N_24198,N_24461);
xor U27307 (N_27307,N_24536,N_26410);
nor U27308 (N_27308,N_26828,N_24555);
and U27309 (N_27309,N_25743,N_26878);
or U27310 (N_27310,N_25574,N_25285);
or U27311 (N_27311,N_26730,N_25752);
nand U27312 (N_27312,N_24852,N_25224);
or U27313 (N_27313,N_25658,N_24948);
or U27314 (N_27314,N_26316,N_25627);
xnor U27315 (N_27315,N_24157,N_24619);
and U27316 (N_27316,N_26834,N_24707);
nand U27317 (N_27317,N_25923,N_26687);
nand U27318 (N_27318,N_24981,N_25101);
xor U27319 (N_27319,N_25290,N_25552);
xor U27320 (N_27320,N_25107,N_24038);
and U27321 (N_27321,N_24661,N_26681);
or U27322 (N_27322,N_26944,N_24371);
or U27323 (N_27323,N_24854,N_25745);
xor U27324 (N_27324,N_25655,N_25099);
or U27325 (N_27325,N_26849,N_24895);
or U27326 (N_27326,N_25366,N_25143);
nand U27327 (N_27327,N_24066,N_26618);
and U27328 (N_27328,N_26541,N_24907);
xnor U27329 (N_27329,N_25261,N_24625);
nor U27330 (N_27330,N_26182,N_26292);
nand U27331 (N_27331,N_25642,N_24567);
and U27332 (N_27332,N_24432,N_25250);
nand U27333 (N_27333,N_25058,N_26046);
xor U27334 (N_27334,N_26762,N_25802);
xor U27335 (N_27335,N_25419,N_25790);
nand U27336 (N_27336,N_25983,N_25700);
nor U27337 (N_27337,N_24788,N_26656);
and U27338 (N_27338,N_25828,N_24078);
nor U27339 (N_27339,N_24129,N_24743);
and U27340 (N_27340,N_24532,N_25288);
and U27341 (N_27341,N_24171,N_25671);
nor U27342 (N_27342,N_25221,N_25619);
or U27343 (N_27343,N_24600,N_25109);
and U27344 (N_27344,N_25831,N_25665);
xnor U27345 (N_27345,N_26187,N_26232);
nor U27346 (N_27346,N_25462,N_25504);
or U27347 (N_27347,N_25038,N_25273);
nand U27348 (N_27348,N_25920,N_24314);
nor U27349 (N_27349,N_26898,N_25712);
xnor U27350 (N_27350,N_25222,N_25239);
xor U27351 (N_27351,N_24564,N_26626);
or U27352 (N_27352,N_24269,N_26620);
xnor U27353 (N_27353,N_25989,N_26043);
xnor U27354 (N_27354,N_26622,N_24970);
xor U27355 (N_27355,N_25796,N_26439);
nor U27356 (N_27356,N_25596,N_25350);
xnor U27357 (N_27357,N_24357,N_26671);
nor U27358 (N_27358,N_24114,N_25526);
and U27359 (N_27359,N_25572,N_24484);
or U27360 (N_27360,N_26058,N_25957);
xnor U27361 (N_27361,N_26228,N_26308);
nor U27362 (N_27362,N_24122,N_24570);
and U27363 (N_27363,N_24752,N_25488);
or U27364 (N_27364,N_26380,N_26149);
nor U27365 (N_27365,N_25569,N_24404);
nor U27366 (N_27366,N_25683,N_24322);
or U27367 (N_27367,N_25991,N_26350);
or U27368 (N_27368,N_24670,N_25768);
nand U27369 (N_27369,N_25156,N_25716);
or U27370 (N_27370,N_26741,N_25691);
nand U27371 (N_27371,N_26449,N_26123);
or U27372 (N_27372,N_25904,N_25949);
nand U27373 (N_27373,N_24210,N_24379);
xor U27374 (N_27374,N_24355,N_24408);
nor U27375 (N_27375,N_25964,N_24225);
xor U27376 (N_27376,N_26504,N_24128);
or U27377 (N_27377,N_25301,N_26289);
or U27378 (N_27378,N_25090,N_25377);
nand U27379 (N_27379,N_25287,N_25021);
nand U27380 (N_27380,N_25248,N_26702);
or U27381 (N_27381,N_26059,N_25610);
xnor U27382 (N_27382,N_25031,N_25675);
xnor U27383 (N_27383,N_24694,N_26379);
or U27384 (N_27384,N_25476,N_24427);
and U27385 (N_27385,N_25725,N_25958);
or U27386 (N_27386,N_24784,N_24928);
and U27387 (N_27387,N_26967,N_24459);
nand U27388 (N_27388,N_24571,N_24958);
nor U27389 (N_27389,N_26181,N_24411);
and U27390 (N_27390,N_25305,N_24972);
nor U27391 (N_27391,N_26143,N_25392);
xnor U27392 (N_27392,N_24217,N_25842);
nand U27393 (N_27393,N_24724,N_24176);
xor U27394 (N_27394,N_25891,N_26900);
or U27395 (N_27395,N_25485,N_24489);
nor U27396 (N_27396,N_26384,N_24089);
xnor U27397 (N_27397,N_26779,N_25317);
and U27398 (N_27398,N_25383,N_25577);
or U27399 (N_27399,N_26017,N_25755);
and U27400 (N_27400,N_24319,N_26679);
nor U27401 (N_27401,N_25044,N_24961);
xnor U27402 (N_27402,N_24417,N_24256);
or U27403 (N_27403,N_26435,N_26098);
nor U27404 (N_27404,N_25269,N_25528);
and U27405 (N_27405,N_25098,N_24964);
nand U27406 (N_27406,N_25040,N_24623);
nor U27407 (N_27407,N_25029,N_25592);
or U27408 (N_27408,N_26960,N_26986);
xor U27409 (N_27409,N_24676,N_24189);
and U27410 (N_27410,N_24488,N_25458);
nor U27411 (N_27411,N_26990,N_26794);
nand U27412 (N_27412,N_25138,N_25928);
and U27413 (N_27413,N_26609,N_25282);
nor U27414 (N_27414,N_25424,N_25834);
and U27415 (N_27415,N_25255,N_24656);
xnor U27416 (N_27416,N_26474,N_26759);
nand U27417 (N_27417,N_26522,N_26870);
and U27418 (N_27418,N_26199,N_24560);
xor U27419 (N_27419,N_25063,N_26631);
nor U27420 (N_27420,N_25448,N_24468);
or U27421 (N_27421,N_24806,N_25961);
or U27422 (N_27422,N_24400,N_26542);
and U27423 (N_27423,N_26805,N_25379);
and U27424 (N_27424,N_25857,N_24372);
nand U27425 (N_27425,N_25295,N_24808);
xnor U27426 (N_27426,N_25082,N_26822);
and U27427 (N_27427,N_25591,N_25771);
xor U27428 (N_27428,N_26930,N_24649);
nand U27429 (N_27429,N_26997,N_24169);
or U27430 (N_27430,N_26103,N_24968);
nor U27431 (N_27431,N_25203,N_25707);
xnor U27432 (N_27432,N_25751,N_26438);
nand U27433 (N_27433,N_26680,N_25034);
and U27434 (N_27434,N_24836,N_24140);
nand U27435 (N_27435,N_26611,N_26221);
and U27436 (N_27436,N_25463,N_25838);
nor U27437 (N_27437,N_24506,N_25950);
nor U27438 (N_27438,N_25888,N_26049);
nand U27439 (N_27439,N_26351,N_25765);
xor U27440 (N_27440,N_24234,N_26582);
nand U27441 (N_27441,N_26469,N_24139);
and U27442 (N_27442,N_24024,N_24056);
or U27443 (N_27443,N_25432,N_25589);
nor U27444 (N_27444,N_26125,N_25438);
nor U27445 (N_27445,N_26295,N_24835);
or U27446 (N_27446,N_26140,N_24190);
or U27447 (N_27447,N_24274,N_24029);
nor U27448 (N_27448,N_26545,N_24443);
nand U27449 (N_27449,N_25084,N_26457);
nor U27450 (N_27450,N_26312,N_26745);
nand U27451 (N_27451,N_25519,N_24647);
or U27452 (N_27452,N_25788,N_25505);
or U27453 (N_27453,N_24199,N_24941);
nor U27454 (N_27454,N_24267,N_25418);
or U27455 (N_27455,N_24704,N_24381);
nand U27456 (N_27456,N_25708,N_26461);
nor U27457 (N_27457,N_25934,N_26775);
nand U27458 (N_27458,N_24033,N_25180);
or U27459 (N_27459,N_26475,N_26529);
nor U27460 (N_27460,N_26905,N_25815);
nand U27461 (N_27461,N_24460,N_26386);
and U27462 (N_27462,N_24437,N_25114);
or U27463 (N_27463,N_26994,N_24250);
or U27464 (N_27464,N_24867,N_25296);
and U27465 (N_27465,N_25117,N_24452);
nor U27466 (N_27466,N_24430,N_25780);
or U27467 (N_27467,N_25748,N_26330);
nand U27468 (N_27468,N_24911,N_26737);
and U27469 (N_27469,N_26548,N_26910);
xnor U27470 (N_27470,N_26211,N_25358);
and U27471 (N_27471,N_24368,N_24412);
nor U27472 (N_27472,N_24285,N_25809);
nand U27473 (N_27473,N_26315,N_25511);
nand U27474 (N_27474,N_24039,N_25543);
nor U27475 (N_27475,N_26244,N_26616);
nor U27476 (N_27476,N_25693,N_24469);
nor U27477 (N_27477,N_26048,N_26130);
nor U27478 (N_27478,N_26019,N_26302);
nor U27479 (N_27479,N_26629,N_24927);
nand U27480 (N_27480,N_24979,N_26381);
nor U27481 (N_27481,N_26867,N_26830);
xor U27482 (N_27482,N_25562,N_25118);
or U27483 (N_27483,N_24475,N_25115);
and U27484 (N_27484,N_25150,N_25643);
xnor U27485 (N_27485,N_26850,N_24232);
nand U27486 (N_27486,N_26594,N_26484);
nand U27487 (N_27487,N_26015,N_24878);
nand U27488 (N_27488,N_24790,N_25294);
nand U27489 (N_27489,N_24991,N_26412);
and U27490 (N_27490,N_25620,N_26556);
xnor U27491 (N_27491,N_25901,N_24581);
xor U27492 (N_27492,N_26339,N_25611);
nor U27493 (N_27493,N_24765,N_24620);
and U27494 (N_27494,N_26225,N_24147);
or U27495 (N_27495,N_26333,N_24354);
nor U27496 (N_27496,N_26782,N_25628);
or U27497 (N_27497,N_24457,N_25009);
or U27498 (N_27498,N_26338,N_26639);
nand U27499 (N_27499,N_24442,N_25986);
xnor U27500 (N_27500,N_26095,N_26801);
xor U27501 (N_27501,N_26606,N_24668);
nand U27502 (N_27502,N_26842,N_24746);
and U27503 (N_27503,N_24538,N_24680);
nand U27504 (N_27504,N_25000,N_24108);
nor U27505 (N_27505,N_26089,N_25380);
or U27506 (N_27506,N_26882,N_25895);
or U27507 (N_27507,N_25580,N_25914);
nor U27508 (N_27508,N_25819,N_25738);
xnor U27509 (N_27509,N_25079,N_26713);
nand U27510 (N_27510,N_24840,N_24616);
xor U27511 (N_27511,N_25345,N_25410);
or U27512 (N_27512,N_25799,N_25516);
or U27513 (N_27513,N_25616,N_26988);
nor U27514 (N_27514,N_26122,N_25204);
nand U27515 (N_27515,N_24168,N_24304);
nand U27516 (N_27516,N_26141,N_25696);
xor U27517 (N_27517,N_24789,N_26426);
nand U27518 (N_27518,N_25188,N_25985);
and U27519 (N_27519,N_24604,N_26938);
or U27520 (N_27520,N_24099,N_26642);
and U27521 (N_27521,N_24635,N_24318);
or U27522 (N_27522,N_25795,N_26145);
and U27523 (N_27523,N_24244,N_24919);
xor U27524 (N_27524,N_26706,N_24364);
and U27525 (N_27525,N_24508,N_25617);
or U27526 (N_27526,N_24612,N_24638);
nand U27527 (N_27527,N_24374,N_26018);
and U27528 (N_27528,N_25404,N_26328);
and U27529 (N_27529,N_25342,N_25411);
or U27530 (N_27530,N_25744,N_25878);
or U27531 (N_27531,N_26744,N_26045);
or U27532 (N_27532,N_24553,N_24281);
nor U27533 (N_27533,N_25680,N_24470);
nor U27534 (N_27534,N_25171,N_24289);
or U27535 (N_27535,N_26798,N_24496);
nor U27536 (N_27536,N_25365,N_24926);
or U27537 (N_27537,N_26709,N_26632);
or U27538 (N_27538,N_26964,N_24013);
or U27539 (N_27539,N_25710,N_26392);
nor U27540 (N_27540,N_26743,N_26271);
nand U27541 (N_27541,N_26275,N_26458);
and U27542 (N_27542,N_25979,N_26624);
nor U27543 (N_27543,N_25408,N_24418);
xor U27544 (N_27544,N_25360,N_25401);
or U27545 (N_27545,N_24054,N_26558);
and U27546 (N_27546,N_26400,N_25863);
or U27547 (N_27547,N_26601,N_25633);
nor U27548 (N_27548,N_26662,N_25321);
or U27549 (N_27549,N_26075,N_24812);
nor U27550 (N_27550,N_25232,N_24940);
xor U27551 (N_27551,N_25263,N_24719);
and U27552 (N_27552,N_26188,N_24577);
nand U27553 (N_27553,N_24876,N_25449);
nand U27554 (N_27554,N_26733,N_24510);
nand U27555 (N_27555,N_24303,N_24486);
nand U27556 (N_27556,N_24277,N_24462);
xor U27557 (N_27557,N_25385,N_24104);
nor U27558 (N_27558,N_26142,N_24081);
xnor U27559 (N_27559,N_25217,N_26021);
xnor U27560 (N_27560,N_24133,N_26735);
and U27561 (N_27561,N_24877,N_25756);
and U27562 (N_27562,N_25209,N_26766);
xnor U27563 (N_27563,N_25131,N_25930);
nand U27564 (N_27564,N_24444,N_25166);
nand U27565 (N_27565,N_26193,N_25370);
or U27566 (N_27566,N_24049,N_25422);
xor U27567 (N_27567,N_26718,N_24116);
xnor U27568 (N_27568,N_26581,N_25333);
and U27569 (N_27569,N_24260,N_24557);
nor U27570 (N_27570,N_25727,N_26692);
nand U27571 (N_27571,N_26409,N_26943);
and U27572 (N_27572,N_26120,N_25739);
nand U27573 (N_27573,N_25668,N_24705);
or U27574 (N_27574,N_25778,N_26957);
xor U27575 (N_27575,N_24220,N_25234);
xor U27576 (N_27576,N_25847,N_24242);
or U27577 (N_27577,N_26322,N_26649);
nor U27578 (N_27578,N_26072,N_26223);
or U27579 (N_27579,N_25478,N_26273);
or U27580 (N_27580,N_25467,N_24376);
nor U27581 (N_27581,N_24627,N_25206);
xnor U27582 (N_27582,N_24677,N_24865);
or U27583 (N_27583,N_26560,N_26079);
xor U27584 (N_27584,N_26240,N_25937);
or U27585 (N_27585,N_24561,N_25889);
and U27586 (N_27586,N_25399,N_25531);
nor U27587 (N_27587,N_26290,N_24683);
and U27588 (N_27588,N_26991,N_25630);
and U27589 (N_27589,N_26712,N_26062);
or U27590 (N_27590,N_25614,N_25225);
nand U27591 (N_27591,N_26592,N_25736);
xor U27592 (N_27592,N_26270,N_24473);
xor U27593 (N_27593,N_26175,N_24405);
or U27594 (N_27594,N_26664,N_24215);
or U27595 (N_27595,N_26690,N_25702);
nor U27596 (N_27596,N_24545,N_26825);
and U27597 (N_27597,N_26287,N_26901);
nand U27598 (N_27598,N_25240,N_24639);
xnor U27599 (N_27599,N_25158,N_24161);
and U27600 (N_27600,N_24858,N_25946);
nand U27601 (N_27601,N_24653,N_26250);
nand U27602 (N_27602,N_26628,N_24558);
xnor U27603 (N_27603,N_24706,N_24578);
or U27604 (N_27604,N_26012,N_24599);
xnor U27605 (N_27605,N_24264,N_24750);
xnor U27606 (N_27606,N_26885,N_26243);
and U27607 (N_27607,N_26972,N_25292);
or U27608 (N_27608,N_26218,N_24438);
or U27609 (N_27609,N_25740,N_24195);
and U27610 (N_27610,N_24820,N_25657);
nand U27611 (N_27611,N_25650,N_25774);
or U27612 (N_27612,N_25052,N_24057);
nand U27613 (N_27613,N_24019,N_25233);
nor U27614 (N_27614,N_25721,N_26677);
and U27615 (N_27615,N_26446,N_26482);
xor U27616 (N_27616,N_24035,N_24986);
nor U27617 (N_27617,N_26112,N_26968);
nor U27618 (N_27618,N_26777,N_26466);
xnor U27619 (N_27619,N_24848,N_26230);
xor U27620 (N_27620,N_25205,N_24315);
nor U27621 (N_27621,N_24305,N_25420);
or U27622 (N_27622,N_24296,N_26831);
or U27623 (N_27623,N_26700,N_25644);
or U27624 (N_27624,N_26554,N_24014);
and U27625 (N_27625,N_24918,N_24535);
xnor U27626 (N_27626,N_25770,N_25057);
nor U27627 (N_27627,N_26060,N_25161);
xor U27628 (N_27628,N_25760,N_24544);
xnor U27629 (N_27629,N_26153,N_25536);
and U27630 (N_27630,N_24310,N_24971);
and U27631 (N_27631,N_25941,N_24985);
nor U27632 (N_27632,N_26389,N_25347);
and U27633 (N_27633,N_24450,N_24166);
nand U27634 (N_27634,N_25843,N_26463);
xnor U27635 (N_27635,N_26995,N_24088);
xnor U27636 (N_27636,N_26945,N_25284);
and U27637 (N_27637,N_25837,N_25105);
nand U27638 (N_27638,N_26139,N_26425);
nand U27639 (N_27639,N_26088,N_26605);
nor U27640 (N_27640,N_26772,N_25522);
or U27641 (N_27641,N_25741,N_26488);
nand U27642 (N_27642,N_26916,N_26465);
xor U27643 (N_27643,N_26932,N_25003);
nor U27644 (N_27644,N_25684,N_24485);
nand U27645 (N_27645,N_24547,N_25315);
or U27646 (N_27646,N_26946,N_25337);
or U27647 (N_27647,N_25908,N_24708);
xnor U27648 (N_27648,N_24768,N_24290);
xnor U27649 (N_27649,N_26041,N_25609);
nor U27650 (N_27650,N_25587,N_24766);
nor U27651 (N_27651,N_24756,N_24165);
or U27652 (N_27652,N_24453,N_26138);
or U27653 (N_27653,N_25885,N_24295);
xor U27654 (N_27654,N_26023,N_25216);
nand U27655 (N_27655,N_26231,N_25186);
nand U27656 (N_27656,N_26441,N_25343);
xnor U27657 (N_27657,N_25879,N_25600);
nand U27658 (N_27658,N_26923,N_24363);
and U27659 (N_27659,N_26430,N_26359);
nand U27660 (N_27660,N_24525,N_24580);
nor U27661 (N_27661,N_24351,N_24294);
nor U27662 (N_27662,N_25207,N_24287);
nor U27663 (N_27663,N_25874,N_25887);
nor U27664 (N_27664,N_25134,N_26336);
or U27665 (N_27665,N_26210,N_26033);
and U27666 (N_27666,N_25223,N_26641);
xor U27667 (N_27667,N_24331,N_25554);
nand U27668 (N_27668,N_24575,N_25856);
nor U27669 (N_27669,N_26929,N_26477);
or U27670 (N_27670,N_24996,N_26987);
xor U27671 (N_27671,N_25076,N_24109);
nor U27672 (N_27672,N_26939,N_26154);
nor U27673 (N_27673,N_25583,N_25106);
nand U27674 (N_27674,N_24987,N_25066);
or U27675 (N_27675,N_26169,N_26454);
nor U27676 (N_27676,N_24778,N_26654);
xnor U27677 (N_27677,N_25088,N_26031);
and U27678 (N_27678,N_26067,N_25527);
and U27679 (N_27679,N_24772,N_25974);
or U27680 (N_27680,N_25454,N_25737);
xnor U27681 (N_27681,N_24693,N_24803);
or U27682 (N_27682,N_25012,N_26555);
xor U27683 (N_27683,N_24258,N_24113);
or U27684 (N_27684,N_25855,N_26971);
nor U27685 (N_27685,N_24084,N_25534);
or U27686 (N_27686,N_24362,N_26101);
nand U27687 (N_27687,N_25875,N_25382);
nor U27688 (N_27688,N_25452,N_24591);
nand U27689 (N_27689,N_24641,N_25236);
and U27690 (N_27690,N_24675,N_26734);
nor U27691 (N_27691,N_24236,N_24115);
nand U27692 (N_27692,N_25077,N_24537);
and U27693 (N_27693,N_26612,N_24481);
nor U27694 (N_27694,N_24799,N_26596);
nand U27695 (N_27695,N_25303,N_26535);
and U27696 (N_27696,N_24903,N_25864);
nor U27697 (N_27697,N_24216,N_24651);
nor U27698 (N_27698,N_24083,N_24471);
nor U27699 (N_27699,N_24010,N_26954);
or U27700 (N_27700,N_26177,N_25165);
and U27701 (N_27701,N_25081,N_24905);
xor U27702 (N_27702,N_26841,N_25689);
xnor U27703 (N_27703,N_26151,N_26811);
xnor U27704 (N_27704,N_25024,N_24910);
and U27705 (N_27705,N_25877,N_25348);
xnor U27706 (N_27706,N_26950,N_24500);
nor U27707 (N_27707,N_24185,N_26172);
xor U27708 (N_27708,N_26194,N_24134);
and U27709 (N_27709,N_25074,N_26114);
or U27710 (N_27710,N_26753,N_26305);
or U27711 (N_27711,N_26111,N_25313);
nor U27712 (N_27712,N_24698,N_24238);
and U27713 (N_27713,N_26497,N_26586);
or U27714 (N_27714,N_25384,N_24507);
xnor U27715 (N_27715,N_26703,N_25973);
and U27716 (N_27716,N_24710,N_24843);
nand U27717 (N_27717,N_26561,N_25018);
nor U27718 (N_27718,N_26580,N_25805);
xor U27719 (N_27719,N_25387,N_24097);
nor U27720 (N_27720,N_25395,N_26293);
nand U27721 (N_27721,N_24491,N_26092);
xor U27722 (N_27722,N_26404,N_26829);
or U27723 (N_27723,N_24498,N_25590);
nor U27724 (N_27724,N_24266,N_26424);
nand U27725 (N_27725,N_25530,N_25541);
nand U27726 (N_27726,N_25159,N_26437);
and U27727 (N_27727,N_26129,N_26732);
and U27728 (N_27728,N_26603,N_26668);
nor U27729 (N_27729,N_26197,N_24916);
nor U27730 (N_27730,N_26678,N_25331);
nor U27731 (N_27731,N_25775,N_26564);
nand U27732 (N_27732,N_24980,N_25798);
and U27733 (N_27733,N_26666,N_25915);
xor U27734 (N_27734,N_25339,N_24375);
or U27735 (N_27735,N_24744,N_25378);
and U27736 (N_27736,N_25152,N_25116);
xnor U27737 (N_27737,N_25567,N_24251);
or U27738 (N_27738,N_26839,N_24336);
nand U27739 (N_27739,N_24182,N_24847);
and U27740 (N_27740,N_26670,N_24502);
or U27741 (N_27741,N_26363,N_24283);
and U27742 (N_27742,N_25677,N_25087);
xor U27743 (N_27743,N_24999,N_24248);
nor U27744 (N_27744,N_24642,N_26908);
or U27745 (N_27745,N_25320,N_26788);
nor U27746 (N_27746,N_26704,N_25852);
nor U27747 (N_27747,N_25376,N_26803);
or U27748 (N_27748,N_26636,N_26299);
and U27749 (N_27749,N_25723,N_25047);
nor U27750 (N_27750,N_24394,N_25229);
nand U27751 (N_27751,N_24206,N_26915);
nor U27752 (N_27752,N_24253,N_26832);
or U27753 (N_27753,N_25561,N_26335);
nor U27754 (N_27754,N_26996,N_25091);
or U27755 (N_27755,N_25976,N_26715);
and U27756 (N_27756,N_26625,N_25674);
xor U27757 (N_27757,N_26855,N_26133);
nor U27758 (N_27758,N_25757,N_25817);
nand U27759 (N_27759,N_24385,N_25868);
nand U27760 (N_27760,N_25808,N_26320);
and U27761 (N_27761,N_26455,N_26016);
nand U27762 (N_27762,N_24246,N_24667);
and U27763 (N_27763,N_24779,N_26104);
xor U27764 (N_27764,N_25839,N_25919);
nor U27765 (N_27765,N_24167,N_26005);
or U27766 (N_27766,N_26117,N_24650);
xnor U27767 (N_27767,N_24192,N_24121);
or U27768 (N_27768,N_26050,N_25268);
and U27769 (N_27769,N_24429,N_24124);
xnor U27770 (N_27770,N_26598,N_26963);
or U27771 (N_27771,N_24699,N_26589);
nor U27772 (N_27772,N_25200,N_24594);
and U27773 (N_27773,N_24782,N_24487);
or U27774 (N_27774,N_25198,N_24490);
nor U27775 (N_27775,N_24333,N_25316);
nor U27776 (N_27776,N_24938,N_25912);
or U27777 (N_27777,N_24603,N_24976);
nand U27778 (N_27778,N_25495,N_26513);
and U27779 (N_27779,N_26094,N_26848);
or U27780 (N_27780,N_25061,N_26675);
and U27781 (N_27781,N_24822,N_25995);
and U27782 (N_27782,N_25351,N_24783);
nor U27783 (N_27783,N_26493,N_24312);
or U27784 (N_27784,N_24636,N_25451);
xor U27785 (N_27785,N_25988,N_25841);
or U27786 (N_27786,N_26003,N_26847);
or U27787 (N_27787,N_25388,N_24663);
nand U27788 (N_27788,N_25283,N_25698);
nand U27789 (N_27789,N_24067,N_26317);
and U27790 (N_27790,N_25494,N_25396);
and U27791 (N_27791,N_25132,N_25496);
nor U27792 (N_27792,N_26168,N_25818);
or U27793 (N_27793,N_26282,N_26166);
nand U27794 (N_27794,N_25368,N_25298);
xnor U27795 (N_27795,N_25262,N_24386);
nor U27796 (N_27796,N_25816,N_26370);
xor U27797 (N_27797,N_26266,N_25753);
or U27798 (N_27798,N_25538,N_26345);
or U27799 (N_27799,N_25328,N_24884);
and U27800 (N_27800,N_24334,N_25533);
and U27801 (N_27801,N_25761,N_25006);
nand U27802 (N_27802,N_24464,N_25936);
and U27803 (N_27803,N_24674,N_26076);
xor U27804 (N_27804,N_24458,N_25902);
xnor U27805 (N_27805,N_26039,N_25663);
xnor U27806 (N_27806,N_26926,N_24091);
and U27807 (N_27807,N_25279,N_24901);
and U27808 (N_27808,N_25046,N_26116);
xnor U27809 (N_27809,N_25421,N_26837);
and U27810 (N_27810,N_24120,N_26483);
and U27811 (N_27811,N_26195,N_25735);
and U27812 (N_27812,N_24098,N_26029);
nor U27813 (N_27813,N_26405,N_25035);
xor U27814 (N_27814,N_25706,N_24348);
xnor U27815 (N_27815,N_25022,N_26858);
nor U27816 (N_27816,N_24482,N_25442);
and U27817 (N_27817,N_24162,N_25025);
nor U27818 (N_27818,N_25606,N_25647);
xor U27819 (N_27819,N_26288,N_25456);
and U27820 (N_27820,N_25372,N_25238);
and U27821 (N_27821,N_26102,N_24243);
nand U27822 (N_27822,N_24223,N_25136);
nor U27823 (N_27823,N_26595,N_26723);
xnor U27824 (N_27824,N_24992,N_26013);
or U27825 (N_27825,N_25220,N_24914);
and U27826 (N_27826,N_26567,N_25330);
nand U27827 (N_27827,N_25998,N_26091);
or U27828 (N_27828,N_25579,N_25982);
and U27829 (N_27829,N_26280,N_24837);
and U27830 (N_27830,N_25581,N_26797);
and U27831 (N_27831,N_25326,N_25615);
nor U27832 (N_27832,N_24082,N_25501);
nand U27833 (N_27833,N_24818,N_25952);
and U27834 (N_27834,N_26109,N_24797);
or U27835 (N_27835,N_26563,N_25078);
nor U27836 (N_27836,N_24863,N_25211);
nor U27837 (N_27837,N_25164,N_25406);
or U27838 (N_27838,N_24588,N_24630);
or U27839 (N_27839,N_26879,N_26913);
nand U27840 (N_27840,N_26635,N_26802);
nand U27841 (N_27841,N_25742,N_26787);
nand U27842 (N_27842,N_24000,N_24700);
and U27843 (N_27843,N_25886,N_26696);
and U27844 (N_27844,N_24152,N_26645);
nor U27845 (N_27845,N_25762,N_24872);
nor U27846 (N_27846,N_25242,N_25306);
xnor U27847 (N_27847,N_24222,N_25830);
nand U27848 (N_27848,N_24945,N_24853);
and U27849 (N_27849,N_24226,N_26936);
and U27850 (N_27850,N_26294,N_26808);
xnor U27851 (N_27851,N_25094,N_24445);
nor U27852 (N_27852,N_24929,N_24540);
and U27853 (N_27853,N_26485,N_26600);
nand U27854 (N_27854,N_24263,N_24891);
nor U27855 (N_27855,N_25704,N_26526);
and U27856 (N_27856,N_26443,N_26663);
xor U27857 (N_27857,N_26052,N_25434);
nor U27858 (N_27858,N_26973,N_25356);
xnor U27859 (N_27859,N_25070,N_26053);
nand U27860 (N_27860,N_24533,N_26309);
or U27861 (N_27861,N_25068,N_25773);
nand U27862 (N_27862,N_24020,N_26506);
nor U27863 (N_27863,N_25545,N_26450);
nand U27864 (N_27864,N_24153,N_25871);
xor U27865 (N_27865,N_25430,N_25202);
nor U27866 (N_27866,N_26131,N_24912);
nor U27867 (N_27867,N_24030,N_26445);
xnor U27868 (N_27868,N_24137,N_26495);
nand U27869 (N_27869,N_25905,N_26918);
or U27870 (N_27870,N_26148,N_24241);
or U27871 (N_27871,N_25714,N_24428);
nor U27872 (N_27872,N_24074,N_26444);
nand U27873 (N_27873,N_24566,N_24472);
and U27874 (N_27874,N_25065,N_25690);
and U27875 (N_27875,N_25777,N_24406);
xnor U27876 (N_27876,N_25898,N_25827);
xnor U27877 (N_27877,N_26557,N_24609);
nor U27878 (N_27878,N_24237,N_24085);
or U27879 (N_27879,N_25032,N_26710);
nand U27880 (N_27880,N_26695,N_25310);
or U27881 (N_27881,N_26408,N_24330);
or U27882 (N_27882,N_25270,N_26375);
nand U27883 (N_27883,N_24311,N_25523);
or U27884 (N_27884,N_26418,N_26619);
nand U27885 (N_27885,N_25794,N_26311);
nor U27886 (N_27886,N_25503,N_24493);
and U27887 (N_27887,N_25722,N_25361);
and U27888 (N_27888,N_25271,N_24326);
or U27889 (N_27889,N_25102,N_26650);
and U27890 (N_27890,N_26593,N_24286);
nor U27891 (N_27891,N_24793,N_26869);
nand U27892 (N_27892,N_24741,N_25769);
and U27893 (N_27893,N_26816,N_25840);
and U27894 (N_27894,N_26024,N_25355);
nand U27895 (N_27895,N_26156,N_25258);
and U27896 (N_27896,N_24664,N_25942);
and U27897 (N_27897,N_26252,N_26951);
nor U27898 (N_27898,N_24100,N_24598);
or U27899 (N_27899,N_24829,N_25549);
xor U27900 (N_27900,N_24426,N_25652);
xnor U27901 (N_27901,N_25340,N_25951);
nand U27902 (N_27902,N_25008,N_24392);
nand U27903 (N_27903,N_26725,N_26276);
and U27904 (N_27904,N_26711,N_26579);
and U27905 (N_27905,N_24781,N_25431);
and U27906 (N_27906,N_26471,N_26843);
and U27907 (N_27907,N_24144,N_26442);
or U27908 (N_27908,N_25160,N_26150);
or U27909 (N_27909,N_24146,N_25575);
or U27910 (N_27910,N_26087,N_25608);
and U27911 (N_27911,N_26502,N_24503);
or U27912 (N_27912,N_26113,N_26836);
nand U27913 (N_27913,N_24476,N_25459);
nor U27914 (N_27914,N_26947,N_25692);
xor U27915 (N_27915,N_26505,N_25427);
nor U27916 (N_27916,N_24673,N_24695);
nand U27917 (N_27917,N_24589,N_25140);
or U27918 (N_27918,N_26784,N_26416);
xnor U27919 (N_27919,N_25701,N_26313);
and U27920 (N_27920,N_24213,N_24817);
nand U27921 (N_27921,N_26569,N_24202);
nor U27922 (N_27922,N_26546,N_24522);
or U27923 (N_27923,N_25730,N_25899);
nor U27924 (N_27924,N_24962,N_24714);
xor U27925 (N_27925,N_24886,N_24632);
xnor U27926 (N_27926,N_24613,N_24224);
xor U27927 (N_27927,N_24920,N_24425);
or U27928 (N_27928,N_24204,N_25585);
or U27929 (N_27929,N_24897,N_26768);
nor U27930 (N_27930,N_24982,N_24291);
and U27931 (N_27931,N_25804,N_24529);
nand U27932 (N_27932,N_26896,N_25042);
nand U27933 (N_27933,N_24527,N_26931);
nand U27934 (N_27934,N_25883,N_24221);
and U27935 (N_27935,N_24949,N_26835);
and U27936 (N_27936,N_24007,N_26201);
and U27937 (N_27937,N_24053,N_26217);
and U27938 (N_27938,N_26357,N_25929);
nor U27939 (N_27939,N_24842,N_26366);
nand U27940 (N_27940,N_25967,N_26584);
nand U27941 (N_27941,N_26959,N_25311);
or U27942 (N_27942,N_25318,N_24678);
nand U27943 (N_27943,N_26608,N_25661);
and U27944 (N_27944,N_25845,N_24856);
xnor U27945 (N_27945,N_25327,N_25907);
xor U27946 (N_27946,N_26917,N_25792);
nand U27947 (N_27947,N_24387,N_24769);
or U27948 (N_27948,N_25064,N_25594);
nor U27949 (N_27949,N_24050,N_24154);
and U27950 (N_27950,N_26260,N_25993);
nand U27951 (N_27951,N_26824,N_25497);
xor U27952 (N_27952,N_25947,N_24463);
and U27953 (N_27953,N_25900,N_26220);
or U27954 (N_27954,N_25096,N_24722);
nor U27955 (N_27955,N_24313,N_26660);
nor U27956 (N_27956,N_25612,N_26912);
or U27957 (N_27957,N_24988,N_24359);
nand U27958 (N_27958,N_24821,N_26928);
or U27959 (N_27959,N_25218,N_26124);
xnor U27960 (N_27960,N_24102,N_25274);
and U27961 (N_27961,N_26044,N_24550);
xnor U27962 (N_27962,N_25971,N_26771);
and U27963 (N_27963,N_24543,N_25785);
xor U27964 (N_27964,N_25547,N_24200);
or U27965 (N_27965,N_25593,N_26796);
or U27966 (N_27966,N_26953,N_25264);
and U27967 (N_27967,N_26105,N_26795);
xor U27968 (N_27968,N_26897,N_26676);
xnor U27969 (N_27969,N_26857,N_26658);
nor U27970 (N_27970,N_24370,N_25553);
and U27971 (N_27971,N_26321,N_25931);
xor U27972 (N_27972,N_24771,N_24515);
nand U27973 (N_27973,N_26178,N_24424);
nand U27974 (N_27974,N_24688,N_24859);
and U27975 (N_27975,N_24552,N_25417);
nand U27976 (N_27976,N_25252,N_26790);
and U27977 (N_27977,N_24513,N_24072);
and U27978 (N_27978,N_26865,N_24896);
xnor U27979 (N_27979,N_24542,N_26346);
nand U27980 (N_27980,N_24393,N_25359);
xor U27981 (N_27981,N_25241,N_26353);
and U27982 (N_27982,N_24900,N_26559);
nor U27983 (N_27983,N_26785,N_24819);
xnor U27984 (N_27984,N_24414,N_26533);
nor U27985 (N_27985,N_26815,N_24520);
and U27986 (N_27986,N_24587,N_25219);
or U27987 (N_27987,N_26247,N_25235);
and U27988 (N_27988,N_24935,N_24761);
nor U27989 (N_27989,N_24002,N_24880);
or U27990 (N_27990,N_26525,N_24930);
nor U27991 (N_27991,N_26037,N_26413);
nand U27992 (N_27992,N_24963,N_25028);
or U27993 (N_27993,N_24055,N_24186);
nor U27994 (N_27994,N_25369,N_25266);
nand U27995 (N_27995,N_25524,N_26851);
xor U27996 (N_27996,N_24040,N_26573);
and U27997 (N_27997,N_24209,N_26521);
nand U27998 (N_27998,N_26070,N_26066);
and U27999 (N_27999,N_24814,N_24751);
and U28000 (N_28000,N_26571,N_25660);
and U28001 (N_28001,N_25821,N_26873);
nand U28002 (N_28002,N_25994,N_26899);
and U28003 (N_28003,N_26726,N_24329);
nand U28004 (N_28004,N_24069,N_26599);
xnor U28005 (N_28005,N_24713,N_24825);
or U28006 (N_28006,N_25019,N_25776);
and U28007 (N_28007,N_25470,N_24523);
or U28008 (N_28008,N_26864,N_24448);
nor U28009 (N_28009,N_26838,N_25786);
nand U28010 (N_28010,N_25715,N_26000);
nand U28011 (N_28011,N_25151,N_25113);
nand U28012 (N_28012,N_26456,N_24005);
nor U28013 (N_28013,N_25517,N_24001);
and U28014 (N_28014,N_26436,N_26773);
or U28015 (N_28015,N_26417,N_26186);
and U28016 (N_28016,N_24849,N_24697);
or U28017 (N_28017,N_24282,N_25194);
or U28018 (N_28018,N_24068,N_25558);
nand U28019 (N_28019,N_25779,N_25515);
nand U28020 (N_28020,N_26840,N_25341);
or U28021 (N_28021,N_26258,N_25508);
or U28022 (N_28022,N_26421,N_25560);
nor U28023 (N_28023,N_26085,N_24353);
or U28024 (N_28024,N_25026,N_26862);
nand U28025 (N_28025,N_26398,N_26906);
nand U28026 (N_28026,N_24572,N_26597);
nand U28027 (N_28027,N_26999,N_26992);
xnor U28028 (N_28028,N_24755,N_24953);
or U28029 (N_28029,N_26955,N_26285);
or U28030 (N_28030,N_24760,N_24273);
nand U28031 (N_28031,N_26174,N_26065);
nand U28032 (N_28032,N_24923,N_24188);
nor U28033 (N_28033,N_26009,N_24293);
and U28034 (N_28034,N_26697,N_26976);
nor U28035 (N_28035,N_26216,N_25033);
nand U28036 (N_28036,N_24954,N_24268);
and U28037 (N_28037,N_26042,N_26570);
nor U28038 (N_28038,N_26159,N_26256);
nor U28039 (N_28039,N_26184,N_26683);
or U28040 (N_28040,N_26106,N_24833);
and U28041 (N_28041,N_26004,N_26429);
xnor U28042 (N_28042,N_25709,N_25890);
and U28043 (N_28043,N_26423,N_24614);
nand U28044 (N_28044,N_26852,N_24270);
nor U28045 (N_28045,N_26800,N_24028);
nor U28046 (N_28046,N_24454,N_26395);
or U28047 (N_28047,N_24640,N_24873);
nor U28048 (N_28048,N_25309,N_24602);
or U28049 (N_28049,N_26020,N_25851);
xor U28050 (N_28050,N_24811,N_24512);
or U28051 (N_28051,N_26428,N_25121);
nand U28052 (N_28052,N_25426,N_25474);
nand U28053 (N_28053,N_24037,N_24142);
nor U28054 (N_28054,N_25312,N_26170);
xnor U28055 (N_28055,N_24451,N_25576);
nand U28056 (N_28056,N_25782,N_24347);
xnor U28057 (N_28057,N_26478,N_25578);
and U28058 (N_28058,N_25429,N_26277);
and U28059 (N_28059,N_26026,N_24586);
xor U28060 (N_28060,N_25334,N_25174);
nand U28061 (N_28061,N_26128,N_26673);
nand U28062 (N_28062,N_25259,N_25537);
and U28063 (N_28063,N_26100,N_24574);
or U28064 (N_28064,N_26402,N_25977);
nor U28065 (N_28065,N_26682,N_24973);
or U28066 (N_28066,N_24717,N_26054);
xnor U28067 (N_28067,N_26107,N_24777);
nor U28068 (N_28068,N_24780,N_25896);
or U28069 (N_28069,N_26157,N_24622);
nor U28070 (N_28070,N_24665,N_25787);
nand U28071 (N_28071,N_25289,N_26158);
nand U28072 (N_28072,N_24164,N_24467);
nand U28073 (N_28073,N_26763,N_26998);
nor U28074 (N_28074,N_24718,N_26607);
xnor U28075 (N_28075,N_25112,N_26517);
and U28076 (N_28076,N_25325,N_24027);
xnor U28077 (N_28077,N_24807,N_26185);
and U28078 (N_28078,N_25457,N_24950);
and U28079 (N_28079,N_26394,N_26083);
and U28080 (N_28080,N_26985,N_25566);
nand U28081 (N_28081,N_24230,N_25423);
and U28082 (N_28082,N_26977,N_24690);
and U28083 (N_28083,N_26894,N_25354);
nand U28084 (N_28084,N_25784,N_26880);
nor U28085 (N_28085,N_26268,N_25542);
nor U28086 (N_28086,N_26827,N_25695);
nor U28087 (N_28087,N_24585,N_26806);
or U28088 (N_28088,N_26956,N_24890);
and U28089 (N_28089,N_24211,N_26035);
xor U28090 (N_28090,N_26643,N_25323);
and U28091 (N_28091,N_24361,N_24366);
or U28092 (N_28092,N_26585,N_25338);
nand U28093 (N_28093,N_24531,N_25997);
nand U28094 (N_28094,N_25123,N_25391);
or U28095 (N_28095,N_25189,N_25846);
nand U28096 (N_28096,N_26378,N_24862);
and U28097 (N_28097,N_26728,N_24546);
nand U28098 (N_28098,N_24061,N_26189);
nand U28099 (N_28099,N_25125,N_24804);
or U28100 (N_28100,N_25080,N_26086);
xor U28101 (N_28101,N_25231,N_26872);
nor U28102 (N_28102,N_25685,N_24239);
and U28103 (N_28103,N_25933,N_24208);
nor U28104 (N_28104,N_24378,N_26331);
xor U28105 (N_28105,N_26332,N_24738);
nor U28106 (N_28106,N_25257,N_25772);
and U28107 (N_28107,N_26689,N_24399);
and U28108 (N_28108,N_24767,N_24103);
xor U28109 (N_28109,N_24629,N_24090);
nand U28110 (N_28110,N_26387,N_24956);
xnor U28111 (N_28111,N_24117,N_26235);
nor U28112 (N_28112,N_26399,N_26844);
nor U28113 (N_28113,N_24480,N_24045);
and U28114 (N_28114,N_26419,N_26826);
or U28115 (N_28115,N_25956,N_25277);
nand U28116 (N_28116,N_26846,N_26348);
nand U28117 (N_28117,N_24004,N_26343);
nor U28118 (N_28118,N_25428,N_24662);
xnor U28119 (N_28119,N_25092,N_24073);
or U28120 (N_28120,N_26888,N_24681);
or U28121 (N_28121,N_25666,N_24272);
nor U28122 (N_28122,N_25072,N_25713);
nor U28123 (N_28123,N_25412,N_24135);
nor U28124 (N_28124,N_26819,N_26397);
nand U28125 (N_28125,N_24415,N_26665);
nor U28126 (N_28126,N_24118,N_24868);
and U28127 (N_28127,N_25636,N_26907);
or U28128 (N_28128,N_25393,N_24297);
nor U28129 (N_28129,N_26530,N_25201);
xor U28130 (N_28130,N_25797,N_26110);
nand U28131 (N_28131,N_25510,N_25681);
or U28132 (N_28132,N_25085,N_24388);
xor U28133 (N_28133,N_24159,N_25980);
or U28134 (N_28134,N_24125,N_25910);
nor U28135 (N_28135,N_25844,N_24254);
nor U28136 (N_28136,N_25984,N_24576);
or U28137 (N_28137,N_24723,N_25445);
xor U28138 (N_28138,N_24974,N_26121);
xor U28139 (N_28139,N_25481,N_26281);
nor U28140 (N_28140,N_26476,N_25718);
nor U28141 (N_28141,N_24183,N_26904);
nor U28142 (N_28142,N_26729,N_24684);
and U28143 (N_28143,N_26298,N_25622);
and U28144 (N_28144,N_24339,N_25400);
and U28145 (N_28145,N_24369,N_25056);
nor U28146 (N_28146,N_25687,N_24145);
nor U28147 (N_28147,N_26467,N_26633);
xnor U28148 (N_28148,N_26340,N_25940);
nor U28149 (N_28149,N_25059,N_25322);
xnor U28150 (N_28150,N_26969,N_26006);
xnor U28151 (N_28151,N_24637,N_25173);
nand U28152 (N_28152,N_25489,N_26300);
xor U28153 (N_28153,N_25764,N_26979);
nand U28154 (N_28154,N_24932,N_25978);
or U28155 (N_28155,N_24728,N_25122);
and U28156 (N_28156,N_25060,N_24391);
and U28157 (N_28157,N_24328,N_25447);
xor U28158 (N_28158,N_26224,N_26069);
xor U28159 (N_28159,N_26651,N_24590);
xor U28160 (N_28160,N_26948,N_25866);
and U28161 (N_28161,N_26264,N_26874);
or U28162 (N_28162,N_25860,N_26699);
and U28163 (N_28163,N_26077,N_24389);
and U28164 (N_28164,N_26621,N_24584);
xor U28165 (N_28165,N_24795,N_26040);
or U28166 (N_28166,N_24196,N_26136);
xor U28167 (N_28167,N_26388,N_24155);
and U28168 (N_28168,N_25732,N_25135);
nand U28169 (N_28169,N_26528,N_24615);
and U28170 (N_28170,N_24352,N_25004);
nand U28171 (N_28171,N_24150,N_25002);
and U28172 (N_28172,N_26765,N_25924);
nor U28173 (N_28173,N_24944,N_24022);
nand U28174 (N_28174,N_24607,N_26755);
or U28175 (N_28175,N_26364,N_25142);
nand U28176 (N_28176,N_24997,N_26547);
or U28177 (N_28177,N_25763,N_24197);
nand U28178 (N_28178,N_26385,N_26144);
xor U28179 (N_28179,N_25607,N_26630);
and U28180 (N_28180,N_25493,N_26919);
nand U28181 (N_28181,N_25911,N_24593);
xor U28182 (N_28182,N_24643,N_25807);
nand U28183 (N_28183,N_26911,N_24130);
or U28184 (N_28184,N_25357,N_25734);
and U28185 (N_28185,N_25916,N_25717);
xnor U28186 (N_28186,N_25403,N_25506);
and U28187 (N_28187,N_24409,N_25965);
and U28188 (N_28188,N_26895,N_25963);
nand U28189 (N_28189,N_26499,N_25750);
and U28190 (N_28190,N_26207,N_26284);
nor U28191 (N_28191,N_24184,N_26717);
nand U28192 (N_28192,N_26032,N_26176);
or U28193 (N_28193,N_26587,N_24889);
nor U28194 (N_28194,N_25646,N_26367);
and U28195 (N_28195,N_25651,N_25177);
xnor U28196 (N_28196,N_26411,N_25344);
and U28197 (N_28197,N_25621,N_25013);
or U28198 (N_28198,N_24382,N_26498);
nand U28199 (N_28199,N_24815,N_25473);
xor U28200 (N_28200,N_24955,N_24696);
nor U28201 (N_28201,N_26707,N_25953);
xor U28202 (N_28202,N_26922,N_24770);
nor U28203 (N_28203,N_26135,N_25172);
nand U28204 (N_28204,N_25097,N_26372);
nor U28205 (N_28205,N_24106,N_24156);
xor U28206 (N_28206,N_26891,N_25759);
and U28207 (N_28207,N_25486,N_25535);
nor U28208 (N_28208,N_26420,N_25990);
xor U28209 (N_28209,N_25811,N_25144);
and U28210 (N_28210,N_26727,N_24321);
nor U28211 (N_28211,N_25502,N_26473);
xor U28212 (N_28212,N_24317,N_24279);
xnor U28213 (N_28213,N_26993,N_25632);
or U28214 (N_28214,N_24682,N_24096);
xor U28215 (N_28215,N_26257,N_25487);
or U28216 (N_28216,N_26296,N_25089);
xnor U28217 (N_28217,N_25922,N_24358);
nand U28218 (N_28218,N_24346,N_24299);
nor U28219 (N_28219,N_26198,N_24734);
nor U28220 (N_28220,N_25349,N_24711);
and U28221 (N_28221,N_26082,N_25570);
or U28222 (N_28222,N_25653,N_26572);
nand U28223 (N_28223,N_26814,N_24094);
xnor U28224 (N_28224,N_24401,N_24933);
and U28225 (N_28225,N_24562,N_25686);
xor U28226 (N_28226,N_26254,N_24203);
or U28227 (N_28227,N_26391,N_25939);
xnor U28228 (N_28228,N_24111,N_25329);
xnor U28229 (N_28229,N_25073,N_25832);
or U28230 (N_28230,N_24455,N_24946);
nand U28231 (N_28231,N_24967,N_25179);
or U28232 (N_28232,N_25789,N_25363);
nor U28233 (N_28233,N_25897,N_26470);
nor U28234 (N_28234,N_26238,N_25499);
or U28235 (N_28235,N_26361,N_25184);
and U28236 (N_28236,N_26171,N_26868);
nor U28237 (N_28237,N_26553,N_26952);
or U28238 (N_28238,N_26655,N_24834);
xor U28239 (N_28239,N_25822,N_25436);
nor U28240 (N_28240,N_25062,N_26792);
xnor U28241 (N_28241,N_25075,N_24796);
or U28242 (N_28242,N_24101,N_25548);
xnor U28243 (N_28243,N_24644,N_25230);
or U28244 (N_28244,N_25500,N_24658);
or U28245 (N_28245,N_24556,N_25884);
and U28246 (N_28246,N_26500,N_25170);
xor U28247 (N_28247,N_25037,N_25810);
nor U28248 (N_28248,N_24846,N_24262);
and U28249 (N_28249,N_24380,N_24402);
nand U28250 (N_28250,N_24016,N_25645);
xnor U28251 (N_28251,N_25598,N_25479);
or U28252 (N_28252,N_24360,N_26219);
nor U28253 (N_28253,N_25302,N_25767);
nor U28254 (N_28254,N_25191,N_25913);
nor U28255 (N_28255,N_25800,N_25017);
and U28256 (N_28256,N_26859,N_25425);
or U28257 (N_28257,N_26011,N_24563);
or U28258 (N_28258,N_24606,N_26520);
nor U28259 (N_28259,N_25648,N_26468);
nor U28260 (N_28260,N_26055,N_25005);
nor U28261 (N_28261,N_25175,N_26481);
nor U28262 (N_28262,N_24951,N_26966);
nand U28263 (N_28263,N_26688,N_25071);
or U28264 (N_28264,N_26686,N_25746);
and U28265 (N_28265,N_25854,N_26887);
and U28266 (N_28266,N_24645,N_24245);
xnor U28267 (N_28267,N_26173,N_24993);
nor U28268 (N_28268,N_26241,N_26451);
xnor U28269 (N_28269,N_25584,N_26229);
nand U28270 (N_28270,N_26747,N_25876);
or U28271 (N_28271,N_26496,N_25703);
xnor U28272 (N_28272,N_26731,N_26767);
and U28273 (N_28273,N_25975,N_24857);
nor U28274 (N_28274,N_26434,N_24844);
nor U28275 (N_28275,N_26807,N_24931);
nor U28276 (N_28276,N_25104,N_25227);
nand U28277 (N_28277,N_25954,N_26167);
nand U28278 (N_28278,N_24327,N_25634);
xor U28279 (N_28279,N_25446,N_26761);
nor U28280 (N_28280,N_26373,N_24219);
and U28281 (N_28281,N_25373,N_24759);
xor U28282 (N_28282,N_26812,N_25719);
nand U28283 (N_28283,N_24686,N_26269);
or U28284 (N_28284,N_24474,N_26914);
xnor U28285 (N_28285,N_25146,N_24416);
or U28286 (N_28286,N_26924,N_26222);
nand U28287 (N_28287,N_26010,N_25314);
nor U28288 (N_28288,N_26267,N_24995);
nand U28289 (N_28289,N_24975,N_26942);
nor U28290 (N_28290,N_25659,N_26722);
and U28291 (N_28291,N_24595,N_25468);
or U28292 (N_28292,N_25010,N_24477);
nor U28293 (N_28293,N_25208,N_24132);
nand U28294 (N_28294,N_25861,N_24805);
nor U28295 (N_28295,N_26984,N_25086);
nor U28296 (N_28296,N_26134,N_26323);
or U28297 (N_28297,N_26549,N_24119);
xnor U28298 (N_28298,N_26925,N_26854);
nor U28299 (N_28299,N_24148,N_26813);
or U28300 (N_28300,N_24172,N_25987);
xor U28301 (N_28301,N_24390,N_25299);
xnor U28302 (N_28302,N_24800,N_26538);
and U28303 (N_28303,N_26861,N_26576);
nor U28304 (N_28304,N_24624,N_24383);
nand U28305 (N_28305,N_25280,N_25297);
nor U28306 (N_28306,N_26061,N_24802);
nand U28307 (N_28307,N_26371,N_24187);
nor U28308 (N_28308,N_26460,N_26462);
and U28309 (N_28309,N_25304,N_25124);
xor U28310 (N_28310,N_25212,N_25801);
nand U28311 (N_28311,N_24436,N_25507);
or U28312 (N_28312,N_25141,N_26486);
or U28313 (N_28313,N_25130,N_26552);
or U28314 (N_28314,N_25935,N_25246);
nand U28315 (N_28315,N_26853,N_25586);
nand U28316 (N_28316,N_24178,N_26127);
nand U28317 (N_28317,N_26164,N_24501);
nand U28318 (N_28318,N_26856,N_26742);
or U28319 (N_28319,N_25490,N_24569);
or U28320 (N_28320,N_25100,N_24902);
or U28321 (N_28321,N_25676,N_25480);
nor U28322 (N_28322,N_25820,N_26246);
or U28323 (N_28323,N_25389,N_24071);
and U28324 (N_28324,N_26354,N_24798);
nor U28325 (N_28325,N_24611,N_24851);
nand U28326 (N_28326,N_26889,N_25300);
nand U28327 (N_28327,N_24828,N_26653);
nand U28328 (N_28328,N_26863,N_26283);
xor U28329 (N_28329,N_26845,N_24554);
or U28330 (N_28330,N_26327,N_25155);
xor U28331 (N_28331,N_25253,N_25237);
and U28332 (N_28332,N_26551,N_25256);
or U28333 (N_28333,N_26393,N_26310);
nor U28334 (N_28334,N_25624,N_26637);
or U28335 (N_28335,N_26099,N_25444);
nor U28336 (N_28336,N_26163,N_24356);
nor U28337 (N_28337,N_24112,N_26146);
nor U28338 (N_28338,N_24017,N_24087);
nand U28339 (N_28339,N_25433,N_25439);
nand U28340 (N_28340,N_25414,N_26236);
and U28341 (N_28341,N_24969,N_24059);
nand U28342 (N_28342,N_26001,N_26884);
nand U28343 (N_28343,N_25981,N_25525);
and U28344 (N_28344,N_25450,N_25853);
nor U28345 (N_28345,N_24534,N_24652);
or U28346 (N_28346,N_25969,N_26667);
nor U28347 (N_28347,N_25565,N_26487);
and U28348 (N_28348,N_24915,N_26657);
or U28349 (N_28349,N_26464,N_24866);
and U28350 (N_28350,N_26684,N_26132);
or U28351 (N_28351,N_24921,N_26754);
or U28352 (N_28352,N_24229,N_24832);
nor U28353 (N_28353,N_26209,N_24660);
nor U28354 (N_28354,N_26056,N_24259);
or U28355 (N_28355,N_26701,N_26036);
or U28356 (N_28356,N_24214,N_25970);
nor U28357 (N_28357,N_24689,N_24031);
or U28358 (N_28358,N_25464,N_24731);
or U28359 (N_28359,N_25127,N_24160);
or U28360 (N_28360,N_24787,N_26119);
xnor U28361 (N_28361,N_26489,N_24666);
and U28362 (N_28362,N_24478,N_24034);
or U28363 (N_28363,N_26902,N_25604);
and U28364 (N_28364,N_26374,N_26215);
or U28365 (N_28365,N_25110,N_26155);
or U28366 (N_28366,N_26078,N_26871);
or U28367 (N_28367,N_25397,N_26602);
or U28368 (N_28368,N_26329,N_26047);
nand U28369 (N_28369,N_24913,N_24343);
nand U28370 (N_28370,N_26480,N_26738);
and U28371 (N_28371,N_26909,N_24634);
and U28372 (N_28372,N_24893,N_25613);
or U28373 (N_28373,N_26674,N_24937);
and U28374 (N_28374,N_26940,N_24883);
or U28375 (N_28375,N_25153,N_26949);
or U28376 (N_28376,N_24421,N_26212);
nand U28377 (N_28377,N_25045,N_24592);
xnor U28378 (N_28378,N_24021,N_24095);
nor U28379 (N_28379,N_24341,N_26514);
nand U28380 (N_28380,N_24446,N_24138);
nand U28381 (N_28381,N_26205,N_24942);
or U28382 (N_28382,N_25729,N_26508);
xnor U28383 (N_28383,N_24850,N_24885);
and U28384 (N_28384,N_26196,N_25588);
and U28385 (N_28385,N_24325,N_25649);
xor U28386 (N_28386,N_25720,N_25618);
and U28387 (N_28387,N_25694,N_26403);
nor U28388 (N_28388,N_24127,N_24410);
nor U28389 (N_28389,N_25193,N_26523);
xor U28390 (N_28390,N_26511,N_25921);
xnor U28391 (N_28391,N_26698,N_26566);
or U28392 (N_28392,N_25405,N_25244);
and U28393 (N_28393,N_26014,N_25697);
nor U28394 (N_28394,N_26875,N_26524);
and U28395 (N_28395,N_26644,N_24143);
nor U28396 (N_28396,N_24824,N_25862);
nand U28397 (N_28397,N_26342,N_25673);
xnor U28398 (N_28398,N_24284,N_26893);
and U28399 (N_28399,N_25050,N_26721);
nand U28400 (N_28400,N_25483,N_25927);
or U28401 (N_28401,N_25196,N_26791);
nor U28402 (N_28402,N_25573,N_25484);
nand U28403 (N_28403,N_25183,N_26227);
xnor U28404 (N_28404,N_24163,N_25672);
or U28405 (N_28405,N_25509,N_24342);
and U28406 (N_28406,N_24855,N_24909);
or U28407 (N_28407,N_26165,N_26833);
and U28408 (N_28408,N_24041,N_26866);
or U28409 (N_28409,N_24861,N_25966);
and U28410 (N_28410,N_24332,N_24504);
nor U28411 (N_28411,N_24170,N_24813);
nand U28412 (N_28412,N_24726,N_26781);
and U28413 (N_28413,N_26407,N_25041);
and U28414 (N_28414,N_25602,N_26459);
or U28415 (N_28415,N_25603,N_26778);
or U28416 (N_28416,N_26685,N_25251);
xor U28417 (N_28417,N_24874,N_25128);
or U28418 (N_28418,N_24227,N_24149);
nand U28419 (N_28419,N_25491,N_25514);
xnor U28420 (N_28420,N_26534,N_24065);
nand U28421 (N_28421,N_24737,N_25398);
nor U28422 (N_28422,N_25926,N_24483);
and U28423 (N_28423,N_25631,N_26758);
nand U28424 (N_28424,N_26034,N_26279);
and U28425 (N_28425,N_26780,N_26365);
and U28426 (N_28426,N_24809,N_24060);
and U28427 (N_28427,N_24076,N_26965);
or U28428 (N_28428,N_24257,N_24712);
and U28429 (N_28429,N_25733,N_24423);
and U28430 (N_28430,N_24875,N_26179);
nand U28431 (N_28431,N_24365,N_26516);
and U28432 (N_28432,N_26903,N_26610);
or U28433 (N_28433,N_25199,N_26263);
nor U28434 (N_28434,N_24011,N_26974);
and U28435 (N_28435,N_26226,N_24657);
and U28436 (N_28436,N_25213,N_25641);
and U28437 (N_28437,N_24123,N_26074);
xor U28438 (N_28438,N_26614,N_25781);
nand U28439 (N_28439,N_24864,N_24009);
nor U28440 (N_28440,N_26764,N_25678);
or U28441 (N_28441,N_25529,N_24715);
xor U28442 (N_28442,N_25711,N_24794);
or U28443 (N_28443,N_25873,N_26448);
nor U28444 (N_28444,N_24823,N_24403);
or U28445 (N_28445,N_24064,N_24549);
or U28446 (N_28446,N_25111,N_24757);
xnor U28447 (N_28447,N_24181,N_25466);
and U28448 (N_28448,N_24773,N_24350);
nor U28449 (N_28449,N_24063,N_24633);
nor U28450 (N_28450,N_25556,N_25520);
or U28451 (N_28451,N_26933,N_24275);
and U28452 (N_28452,N_26453,N_26531);
xnor U28453 (N_28453,N_24292,N_24308);
xnor U28454 (N_28454,N_24887,N_26208);
nand U28455 (N_28455,N_25386,N_26980);
nor U28456 (N_28456,N_26746,N_25187);
xnor U28457 (N_28457,N_24530,N_24494);
nand U28458 (N_28458,N_25308,N_26575);
nand U28459 (N_28459,N_25228,N_25435);
xor U28460 (N_28460,N_24228,N_24934);
nand U28461 (N_28461,N_24367,N_26265);
nor U28462 (N_28462,N_25512,N_26724);
xor U28463 (N_28463,N_24924,N_26028);
nor U28464 (N_28464,N_24839,N_26691);
or U28465 (N_28465,N_26008,N_24692);
xor U28466 (N_28466,N_25806,N_26823);
and U28467 (N_28467,N_24917,N_26057);
nor U28468 (N_28468,N_25181,N_26810);
and U28469 (N_28469,N_25027,N_24869);
or U28470 (N_28470,N_26073,N_25192);
or U28471 (N_28471,N_26638,N_25461);
and U28472 (N_28472,N_26433,N_24775);
xnor U28473 (N_28473,N_25472,N_26251);
or U28474 (N_28474,N_26583,N_24191);
xnor U28475 (N_28475,N_24830,N_24631);
nand U28476 (N_28476,N_25793,N_25563);
nor U28477 (N_28477,N_25513,N_24691);
nand U28478 (N_28478,N_25858,N_26068);
nand U28479 (N_28479,N_26274,N_24957);
nand U28480 (N_28480,N_26341,N_25814);
xor U28481 (N_28481,N_24879,N_25163);
xnor U28482 (N_28482,N_25051,N_24671);
nor U28483 (N_28483,N_25477,N_26051);
nand U28484 (N_28484,N_26349,N_24716);
and U28485 (N_28485,N_26752,N_26118);
or U28486 (N_28486,N_24709,N_26958);
nor U28487 (N_28487,N_24785,N_24047);
nor U28488 (N_28488,N_24959,N_26490);
and U28489 (N_28489,N_25015,N_25605);
nor U28490 (N_28490,N_24518,N_25893);
xor U28491 (N_28491,N_25055,N_25324);
and U28492 (N_28492,N_26334,N_26261);
nand U28493 (N_28493,N_25437,N_24548);
xor U28494 (N_28494,N_26935,N_25679);
nor U28495 (N_28495,N_24984,N_24568);
nor U28496 (N_28496,N_26769,N_24565);
xnor U28497 (N_28497,N_24943,N_24776);
nand U28498 (N_28498,N_26789,N_24335);
nor U28499 (N_28499,N_26876,N_25281);
and U28500 (N_28500,N_24488,N_26136);
nor U28501 (N_28501,N_25175,N_24323);
or U28502 (N_28502,N_25226,N_24106);
or U28503 (N_28503,N_24036,N_24187);
xnor U28504 (N_28504,N_25549,N_26211);
and U28505 (N_28505,N_24966,N_24045);
or U28506 (N_28506,N_25289,N_26326);
xnor U28507 (N_28507,N_26075,N_26473);
nor U28508 (N_28508,N_24756,N_25630);
nor U28509 (N_28509,N_25411,N_26003);
nand U28510 (N_28510,N_25590,N_26705);
xor U28511 (N_28511,N_25074,N_24671);
xor U28512 (N_28512,N_25510,N_24716);
and U28513 (N_28513,N_24316,N_26065);
and U28514 (N_28514,N_25968,N_24462);
and U28515 (N_28515,N_25703,N_26806);
xnor U28516 (N_28516,N_26501,N_26141);
nand U28517 (N_28517,N_25691,N_24814);
and U28518 (N_28518,N_26854,N_26608);
or U28519 (N_28519,N_25056,N_26905);
xnor U28520 (N_28520,N_26662,N_24940);
and U28521 (N_28521,N_24818,N_24029);
xor U28522 (N_28522,N_26966,N_25275);
xnor U28523 (N_28523,N_26444,N_24931);
nand U28524 (N_28524,N_24243,N_26928);
or U28525 (N_28525,N_26145,N_25924);
and U28526 (N_28526,N_25537,N_25372);
nor U28527 (N_28527,N_26714,N_25029);
nand U28528 (N_28528,N_24764,N_24123);
nor U28529 (N_28529,N_24133,N_26643);
and U28530 (N_28530,N_26947,N_25698);
nor U28531 (N_28531,N_26155,N_24123);
xnor U28532 (N_28532,N_24437,N_24369);
xnor U28533 (N_28533,N_24129,N_26479);
xor U28534 (N_28534,N_26554,N_26159);
nor U28535 (N_28535,N_24615,N_24660);
nand U28536 (N_28536,N_24071,N_25564);
nand U28537 (N_28537,N_26355,N_24747);
nand U28538 (N_28538,N_26831,N_25926);
or U28539 (N_28539,N_26794,N_24538);
nor U28540 (N_28540,N_26084,N_26567);
and U28541 (N_28541,N_25587,N_25487);
and U28542 (N_28542,N_24892,N_25021);
nor U28543 (N_28543,N_24524,N_24218);
and U28544 (N_28544,N_24311,N_25899);
and U28545 (N_28545,N_26243,N_24942);
and U28546 (N_28546,N_26823,N_24061);
or U28547 (N_28547,N_24588,N_24260);
or U28548 (N_28548,N_25866,N_25381);
or U28549 (N_28549,N_24034,N_24010);
nand U28550 (N_28550,N_25242,N_25145);
nor U28551 (N_28551,N_25774,N_25040);
xnor U28552 (N_28552,N_26316,N_26771);
and U28553 (N_28553,N_25569,N_24466);
and U28554 (N_28554,N_26670,N_25632);
and U28555 (N_28555,N_25127,N_26910);
or U28556 (N_28556,N_24782,N_24980);
or U28557 (N_28557,N_26727,N_25154);
or U28558 (N_28558,N_26946,N_24476);
or U28559 (N_28559,N_25890,N_24499);
or U28560 (N_28560,N_25712,N_26189);
or U28561 (N_28561,N_26957,N_25704);
or U28562 (N_28562,N_26676,N_25848);
nor U28563 (N_28563,N_24377,N_25864);
nor U28564 (N_28564,N_24958,N_25189);
and U28565 (N_28565,N_24627,N_25162);
nand U28566 (N_28566,N_26620,N_24874);
nand U28567 (N_28567,N_26042,N_25526);
nand U28568 (N_28568,N_26494,N_26332);
xor U28569 (N_28569,N_26938,N_26368);
nand U28570 (N_28570,N_26541,N_26203);
or U28571 (N_28571,N_25005,N_26607);
nor U28572 (N_28572,N_26939,N_24083);
nor U28573 (N_28573,N_24819,N_24447);
and U28574 (N_28574,N_24252,N_24800);
nand U28575 (N_28575,N_24136,N_26222);
xor U28576 (N_28576,N_25848,N_24515);
or U28577 (N_28577,N_25944,N_24544);
nor U28578 (N_28578,N_25589,N_26146);
and U28579 (N_28579,N_26561,N_26930);
xor U28580 (N_28580,N_25059,N_25163);
xor U28581 (N_28581,N_24425,N_25238);
xor U28582 (N_28582,N_24778,N_25965);
xnor U28583 (N_28583,N_24915,N_24077);
or U28584 (N_28584,N_25577,N_24071);
nand U28585 (N_28585,N_25197,N_26571);
or U28586 (N_28586,N_25642,N_26113);
nand U28587 (N_28587,N_25891,N_25920);
or U28588 (N_28588,N_24172,N_25226);
nand U28589 (N_28589,N_24832,N_26589);
and U28590 (N_28590,N_26952,N_25721);
or U28591 (N_28591,N_25491,N_24436);
xor U28592 (N_28592,N_26373,N_25410);
nand U28593 (N_28593,N_24007,N_26563);
and U28594 (N_28594,N_24801,N_25141);
nand U28595 (N_28595,N_26703,N_24484);
nand U28596 (N_28596,N_24979,N_24056);
nor U28597 (N_28597,N_26426,N_25062);
and U28598 (N_28598,N_25808,N_25313);
nand U28599 (N_28599,N_26435,N_26650);
nor U28600 (N_28600,N_25610,N_24079);
or U28601 (N_28601,N_26170,N_25436);
nand U28602 (N_28602,N_24853,N_25577);
nand U28603 (N_28603,N_24768,N_25964);
xnor U28604 (N_28604,N_26203,N_24336);
nand U28605 (N_28605,N_26127,N_24951);
nand U28606 (N_28606,N_24526,N_26466);
nand U28607 (N_28607,N_24758,N_24799);
nand U28608 (N_28608,N_24564,N_25818);
xnor U28609 (N_28609,N_24625,N_26944);
xor U28610 (N_28610,N_26035,N_26819);
xor U28611 (N_28611,N_25095,N_25288);
and U28612 (N_28612,N_26130,N_24040);
xnor U28613 (N_28613,N_26872,N_25594);
or U28614 (N_28614,N_25799,N_25390);
nor U28615 (N_28615,N_24698,N_25569);
xor U28616 (N_28616,N_24541,N_24858);
and U28617 (N_28617,N_26927,N_25410);
nor U28618 (N_28618,N_24477,N_24370);
nand U28619 (N_28619,N_25972,N_24427);
nand U28620 (N_28620,N_25855,N_24447);
and U28621 (N_28621,N_26709,N_26910);
nor U28622 (N_28622,N_26443,N_24196);
nor U28623 (N_28623,N_26860,N_25037);
nand U28624 (N_28624,N_26099,N_25251);
nand U28625 (N_28625,N_24260,N_25022);
or U28626 (N_28626,N_24401,N_25436);
nand U28627 (N_28627,N_24664,N_25674);
xnor U28628 (N_28628,N_26041,N_25140);
and U28629 (N_28629,N_25456,N_24701);
xor U28630 (N_28630,N_24113,N_25327);
nor U28631 (N_28631,N_25438,N_26064);
xnor U28632 (N_28632,N_25694,N_25974);
and U28633 (N_28633,N_26640,N_24395);
nand U28634 (N_28634,N_25131,N_24484);
nor U28635 (N_28635,N_24029,N_25810);
xor U28636 (N_28636,N_26892,N_25906);
nor U28637 (N_28637,N_25364,N_26473);
nand U28638 (N_28638,N_24942,N_26554);
and U28639 (N_28639,N_24194,N_26859);
and U28640 (N_28640,N_25363,N_26198);
xnor U28641 (N_28641,N_26833,N_24763);
nor U28642 (N_28642,N_24002,N_26353);
and U28643 (N_28643,N_26087,N_24140);
nand U28644 (N_28644,N_25471,N_25796);
xnor U28645 (N_28645,N_24423,N_26099);
nand U28646 (N_28646,N_24223,N_25179);
or U28647 (N_28647,N_24695,N_24167);
nor U28648 (N_28648,N_25627,N_26518);
xor U28649 (N_28649,N_25463,N_26285);
nor U28650 (N_28650,N_25224,N_24275);
and U28651 (N_28651,N_24315,N_24345);
or U28652 (N_28652,N_26517,N_26069);
and U28653 (N_28653,N_26334,N_25983);
or U28654 (N_28654,N_24617,N_24524);
and U28655 (N_28655,N_24195,N_24817);
xor U28656 (N_28656,N_26238,N_24629);
or U28657 (N_28657,N_24117,N_26011);
nand U28658 (N_28658,N_24635,N_24627);
and U28659 (N_28659,N_25807,N_26995);
xnor U28660 (N_28660,N_26772,N_25817);
nor U28661 (N_28661,N_24235,N_25138);
and U28662 (N_28662,N_26134,N_26801);
xor U28663 (N_28663,N_24619,N_26192);
xnor U28664 (N_28664,N_25225,N_24824);
or U28665 (N_28665,N_26245,N_26819);
xor U28666 (N_28666,N_26019,N_24318);
or U28667 (N_28667,N_25748,N_26707);
xor U28668 (N_28668,N_25313,N_24399);
or U28669 (N_28669,N_25585,N_24294);
and U28670 (N_28670,N_25265,N_25576);
nand U28671 (N_28671,N_26206,N_25356);
or U28672 (N_28672,N_24513,N_26258);
nor U28673 (N_28673,N_26741,N_26458);
nor U28674 (N_28674,N_25499,N_26732);
and U28675 (N_28675,N_24753,N_26879);
nor U28676 (N_28676,N_26708,N_26412);
nor U28677 (N_28677,N_24201,N_25783);
nand U28678 (N_28678,N_25863,N_25899);
and U28679 (N_28679,N_25250,N_24514);
and U28680 (N_28680,N_25529,N_26330);
xnor U28681 (N_28681,N_24340,N_26804);
or U28682 (N_28682,N_24132,N_25212);
nor U28683 (N_28683,N_25523,N_26211);
nand U28684 (N_28684,N_25923,N_25709);
and U28685 (N_28685,N_24339,N_24183);
nand U28686 (N_28686,N_24792,N_25340);
or U28687 (N_28687,N_25221,N_26747);
nand U28688 (N_28688,N_26115,N_24277);
nor U28689 (N_28689,N_26891,N_25150);
xor U28690 (N_28690,N_24106,N_25127);
and U28691 (N_28691,N_26516,N_24989);
or U28692 (N_28692,N_26979,N_24962);
or U28693 (N_28693,N_25780,N_25731);
nand U28694 (N_28694,N_24589,N_25306);
or U28695 (N_28695,N_24664,N_24367);
xnor U28696 (N_28696,N_25020,N_25811);
and U28697 (N_28697,N_26152,N_24885);
nand U28698 (N_28698,N_26615,N_24858);
xnor U28699 (N_28699,N_26268,N_26073);
nand U28700 (N_28700,N_25910,N_24855);
and U28701 (N_28701,N_25486,N_26621);
and U28702 (N_28702,N_24081,N_26088);
nand U28703 (N_28703,N_25233,N_25504);
nor U28704 (N_28704,N_24752,N_24180);
nor U28705 (N_28705,N_24145,N_26314);
nor U28706 (N_28706,N_24447,N_25888);
and U28707 (N_28707,N_26099,N_26993);
and U28708 (N_28708,N_26815,N_25266);
and U28709 (N_28709,N_25916,N_24589);
xor U28710 (N_28710,N_25936,N_24579);
and U28711 (N_28711,N_26544,N_26214);
nand U28712 (N_28712,N_25093,N_25370);
and U28713 (N_28713,N_24467,N_26050);
or U28714 (N_28714,N_24943,N_24817);
and U28715 (N_28715,N_25185,N_26427);
nor U28716 (N_28716,N_26151,N_25139);
or U28717 (N_28717,N_24411,N_26887);
xor U28718 (N_28718,N_24475,N_26795);
or U28719 (N_28719,N_25311,N_24784);
and U28720 (N_28720,N_24646,N_25003);
nand U28721 (N_28721,N_25365,N_26475);
and U28722 (N_28722,N_24362,N_26205);
or U28723 (N_28723,N_24255,N_25164);
nor U28724 (N_28724,N_25055,N_26650);
and U28725 (N_28725,N_26064,N_26568);
nand U28726 (N_28726,N_25114,N_24993);
or U28727 (N_28727,N_26475,N_25337);
and U28728 (N_28728,N_25617,N_24875);
nor U28729 (N_28729,N_26136,N_26652);
and U28730 (N_28730,N_24391,N_25262);
nand U28731 (N_28731,N_26702,N_24354);
nor U28732 (N_28732,N_24071,N_24383);
nor U28733 (N_28733,N_26254,N_25601);
or U28734 (N_28734,N_24107,N_25875);
xnor U28735 (N_28735,N_25841,N_24240);
xnor U28736 (N_28736,N_25188,N_25876);
nand U28737 (N_28737,N_26894,N_24396);
nor U28738 (N_28738,N_25158,N_24230);
nand U28739 (N_28739,N_24003,N_26923);
and U28740 (N_28740,N_25594,N_24303);
and U28741 (N_28741,N_26680,N_25541);
nor U28742 (N_28742,N_24342,N_24074);
xor U28743 (N_28743,N_26342,N_26240);
and U28744 (N_28744,N_25779,N_24118);
and U28745 (N_28745,N_25304,N_24947);
or U28746 (N_28746,N_24526,N_26401);
xor U28747 (N_28747,N_25201,N_25958);
nand U28748 (N_28748,N_25651,N_25044);
and U28749 (N_28749,N_26860,N_25623);
nand U28750 (N_28750,N_26022,N_26365);
nor U28751 (N_28751,N_24894,N_25907);
xor U28752 (N_28752,N_25539,N_24445);
nand U28753 (N_28753,N_25668,N_25346);
xnor U28754 (N_28754,N_25896,N_25379);
or U28755 (N_28755,N_25604,N_24538);
and U28756 (N_28756,N_25760,N_24185);
and U28757 (N_28757,N_26692,N_24749);
nand U28758 (N_28758,N_24115,N_25911);
nand U28759 (N_28759,N_24182,N_25069);
nand U28760 (N_28760,N_25135,N_25589);
or U28761 (N_28761,N_25841,N_25161);
nand U28762 (N_28762,N_24179,N_26183);
and U28763 (N_28763,N_24396,N_26773);
xor U28764 (N_28764,N_24321,N_25456);
nor U28765 (N_28765,N_26993,N_26399);
and U28766 (N_28766,N_24792,N_24368);
or U28767 (N_28767,N_25861,N_25909);
and U28768 (N_28768,N_24022,N_24972);
nor U28769 (N_28769,N_24187,N_26350);
and U28770 (N_28770,N_26660,N_24845);
and U28771 (N_28771,N_24146,N_26592);
nand U28772 (N_28772,N_25445,N_24603);
nand U28773 (N_28773,N_25580,N_25024);
and U28774 (N_28774,N_24737,N_26481);
nor U28775 (N_28775,N_26598,N_24330);
and U28776 (N_28776,N_24582,N_24621);
xor U28777 (N_28777,N_24316,N_25894);
and U28778 (N_28778,N_25115,N_26140);
nor U28779 (N_28779,N_24539,N_26738);
and U28780 (N_28780,N_25395,N_24151);
xnor U28781 (N_28781,N_26301,N_26682);
nor U28782 (N_28782,N_25876,N_24781);
or U28783 (N_28783,N_26854,N_26103);
xor U28784 (N_28784,N_25765,N_25200);
or U28785 (N_28785,N_24516,N_25093);
nand U28786 (N_28786,N_26491,N_26802);
and U28787 (N_28787,N_25254,N_26706);
or U28788 (N_28788,N_25988,N_26697);
nand U28789 (N_28789,N_25561,N_24042);
nand U28790 (N_28790,N_25078,N_24632);
nor U28791 (N_28791,N_24228,N_25835);
xnor U28792 (N_28792,N_26698,N_25754);
nand U28793 (N_28793,N_25091,N_24974);
nor U28794 (N_28794,N_25991,N_24324);
nor U28795 (N_28795,N_26361,N_24117);
xnor U28796 (N_28796,N_24459,N_26886);
or U28797 (N_28797,N_25958,N_24705);
and U28798 (N_28798,N_26713,N_26932);
nor U28799 (N_28799,N_24467,N_25768);
and U28800 (N_28800,N_25482,N_26088);
xor U28801 (N_28801,N_26521,N_26601);
nor U28802 (N_28802,N_26407,N_25325);
nor U28803 (N_28803,N_24001,N_24441);
and U28804 (N_28804,N_26124,N_26799);
xnor U28805 (N_28805,N_25627,N_24679);
or U28806 (N_28806,N_24363,N_25064);
and U28807 (N_28807,N_25771,N_25976);
xnor U28808 (N_28808,N_25763,N_26667);
nand U28809 (N_28809,N_24861,N_26747);
or U28810 (N_28810,N_24269,N_26711);
or U28811 (N_28811,N_26069,N_25281);
and U28812 (N_28812,N_24936,N_26527);
or U28813 (N_28813,N_25135,N_26447);
and U28814 (N_28814,N_24860,N_26234);
nor U28815 (N_28815,N_26225,N_24649);
and U28816 (N_28816,N_26132,N_26370);
xor U28817 (N_28817,N_25896,N_25209);
nand U28818 (N_28818,N_26348,N_25704);
nand U28819 (N_28819,N_25678,N_25723);
or U28820 (N_28820,N_25725,N_26122);
nand U28821 (N_28821,N_26922,N_24358);
nor U28822 (N_28822,N_25704,N_26449);
nand U28823 (N_28823,N_26161,N_24674);
and U28824 (N_28824,N_25668,N_26115);
and U28825 (N_28825,N_24056,N_24835);
and U28826 (N_28826,N_26879,N_26022);
nand U28827 (N_28827,N_26290,N_26574);
xor U28828 (N_28828,N_25039,N_25903);
nand U28829 (N_28829,N_26275,N_26726);
and U28830 (N_28830,N_26569,N_25475);
and U28831 (N_28831,N_26486,N_24221);
and U28832 (N_28832,N_24457,N_26110);
and U28833 (N_28833,N_25960,N_24549);
nand U28834 (N_28834,N_26531,N_25542);
xnor U28835 (N_28835,N_25535,N_25378);
nand U28836 (N_28836,N_24849,N_24105);
nor U28837 (N_28837,N_24237,N_24350);
xor U28838 (N_28838,N_25845,N_25216);
or U28839 (N_28839,N_24129,N_25555);
xnor U28840 (N_28840,N_25956,N_26731);
nand U28841 (N_28841,N_26565,N_26387);
xnor U28842 (N_28842,N_26317,N_26326);
xor U28843 (N_28843,N_24809,N_24346);
nor U28844 (N_28844,N_24641,N_24786);
nor U28845 (N_28845,N_24768,N_25770);
nor U28846 (N_28846,N_24520,N_25197);
and U28847 (N_28847,N_24888,N_25825);
and U28848 (N_28848,N_26365,N_25675);
nand U28849 (N_28849,N_25544,N_26453);
nor U28850 (N_28850,N_24725,N_25910);
or U28851 (N_28851,N_24408,N_26742);
and U28852 (N_28852,N_24931,N_26614);
or U28853 (N_28853,N_24905,N_25878);
or U28854 (N_28854,N_24762,N_25147);
xor U28855 (N_28855,N_25719,N_24018);
nand U28856 (N_28856,N_26726,N_26465);
or U28857 (N_28857,N_25016,N_24624);
nor U28858 (N_28858,N_25174,N_26735);
nand U28859 (N_28859,N_26488,N_25294);
nand U28860 (N_28860,N_25025,N_24478);
xnor U28861 (N_28861,N_25683,N_24659);
nand U28862 (N_28862,N_26964,N_25143);
or U28863 (N_28863,N_25475,N_25356);
or U28864 (N_28864,N_25923,N_26631);
nand U28865 (N_28865,N_24191,N_25080);
or U28866 (N_28866,N_24368,N_25430);
nor U28867 (N_28867,N_24374,N_26331);
or U28868 (N_28868,N_26292,N_26474);
nor U28869 (N_28869,N_25622,N_24126);
nor U28870 (N_28870,N_24819,N_26667);
and U28871 (N_28871,N_26488,N_25316);
nor U28872 (N_28872,N_24975,N_25079);
and U28873 (N_28873,N_25174,N_25122);
or U28874 (N_28874,N_25331,N_26462);
or U28875 (N_28875,N_24986,N_24287);
nor U28876 (N_28876,N_26475,N_25519);
xnor U28877 (N_28877,N_24606,N_25368);
nand U28878 (N_28878,N_26152,N_25097);
and U28879 (N_28879,N_25541,N_24753);
or U28880 (N_28880,N_25408,N_26156);
xor U28881 (N_28881,N_26860,N_26614);
or U28882 (N_28882,N_24701,N_25790);
xnor U28883 (N_28883,N_25608,N_25235);
and U28884 (N_28884,N_25707,N_26806);
nand U28885 (N_28885,N_26701,N_26729);
and U28886 (N_28886,N_25195,N_26770);
nand U28887 (N_28887,N_25933,N_24281);
nand U28888 (N_28888,N_25444,N_26104);
or U28889 (N_28889,N_25409,N_26165);
nor U28890 (N_28890,N_26012,N_25404);
or U28891 (N_28891,N_25534,N_26039);
xnor U28892 (N_28892,N_24568,N_25179);
xor U28893 (N_28893,N_25984,N_25016);
nor U28894 (N_28894,N_25731,N_25876);
xnor U28895 (N_28895,N_24562,N_24560);
and U28896 (N_28896,N_25341,N_24789);
nor U28897 (N_28897,N_24187,N_25371);
xnor U28898 (N_28898,N_24254,N_24931);
nor U28899 (N_28899,N_24167,N_24956);
or U28900 (N_28900,N_26851,N_25815);
nor U28901 (N_28901,N_25539,N_26987);
xor U28902 (N_28902,N_25377,N_24491);
nor U28903 (N_28903,N_25919,N_24489);
xnor U28904 (N_28904,N_25105,N_25291);
xor U28905 (N_28905,N_25846,N_25836);
xnor U28906 (N_28906,N_26635,N_25948);
nor U28907 (N_28907,N_26686,N_25988);
nand U28908 (N_28908,N_24551,N_25376);
or U28909 (N_28909,N_26719,N_24945);
or U28910 (N_28910,N_24439,N_25136);
nand U28911 (N_28911,N_24908,N_25137);
and U28912 (N_28912,N_24669,N_26644);
and U28913 (N_28913,N_24761,N_26190);
nor U28914 (N_28914,N_26931,N_26337);
or U28915 (N_28915,N_24262,N_25269);
nand U28916 (N_28916,N_25675,N_26853);
nand U28917 (N_28917,N_24871,N_26433);
and U28918 (N_28918,N_26287,N_26695);
or U28919 (N_28919,N_25720,N_26650);
nor U28920 (N_28920,N_26317,N_25228);
and U28921 (N_28921,N_26034,N_24311);
or U28922 (N_28922,N_24496,N_24974);
nand U28923 (N_28923,N_25666,N_24137);
nor U28924 (N_28924,N_25706,N_24559);
and U28925 (N_28925,N_24849,N_25588);
xnor U28926 (N_28926,N_26119,N_25170);
and U28927 (N_28927,N_24555,N_25444);
nand U28928 (N_28928,N_26371,N_24555);
and U28929 (N_28929,N_24455,N_25295);
xor U28930 (N_28930,N_25517,N_25349);
xnor U28931 (N_28931,N_25679,N_25172);
nand U28932 (N_28932,N_25750,N_26807);
nand U28933 (N_28933,N_25932,N_24148);
nor U28934 (N_28934,N_24032,N_24895);
nand U28935 (N_28935,N_25015,N_24202);
xnor U28936 (N_28936,N_24051,N_24611);
and U28937 (N_28937,N_24857,N_26739);
or U28938 (N_28938,N_24439,N_26746);
and U28939 (N_28939,N_24350,N_26328);
xnor U28940 (N_28940,N_26779,N_26620);
nand U28941 (N_28941,N_25356,N_26387);
xor U28942 (N_28942,N_26646,N_26326);
and U28943 (N_28943,N_26442,N_24594);
nand U28944 (N_28944,N_25561,N_26662);
nand U28945 (N_28945,N_26645,N_26897);
nand U28946 (N_28946,N_24967,N_26989);
nand U28947 (N_28947,N_25197,N_26697);
nand U28948 (N_28948,N_24372,N_24544);
nand U28949 (N_28949,N_24258,N_25967);
and U28950 (N_28950,N_26631,N_24585);
nand U28951 (N_28951,N_24320,N_26809);
and U28952 (N_28952,N_25637,N_24819);
or U28953 (N_28953,N_25661,N_24727);
xnor U28954 (N_28954,N_24538,N_26416);
nand U28955 (N_28955,N_24767,N_26522);
xor U28956 (N_28956,N_24977,N_25247);
xor U28957 (N_28957,N_26583,N_26753);
and U28958 (N_28958,N_26803,N_25908);
or U28959 (N_28959,N_24440,N_24011);
nand U28960 (N_28960,N_24591,N_24379);
xnor U28961 (N_28961,N_26396,N_26149);
nand U28962 (N_28962,N_26910,N_24785);
nor U28963 (N_28963,N_24358,N_25112);
nor U28964 (N_28964,N_26955,N_24715);
and U28965 (N_28965,N_24966,N_26475);
nor U28966 (N_28966,N_25988,N_24411);
nor U28967 (N_28967,N_26802,N_26211);
and U28968 (N_28968,N_25774,N_25455);
nor U28969 (N_28969,N_25534,N_26687);
xor U28970 (N_28970,N_25197,N_24093);
or U28971 (N_28971,N_24333,N_26821);
or U28972 (N_28972,N_24901,N_26082);
xor U28973 (N_28973,N_24690,N_24898);
and U28974 (N_28974,N_26758,N_24544);
nor U28975 (N_28975,N_24053,N_25905);
and U28976 (N_28976,N_25979,N_26718);
nand U28977 (N_28977,N_26284,N_25296);
and U28978 (N_28978,N_26829,N_26399);
xor U28979 (N_28979,N_24378,N_24616);
nor U28980 (N_28980,N_26032,N_24954);
nand U28981 (N_28981,N_25872,N_24756);
and U28982 (N_28982,N_26331,N_25645);
nand U28983 (N_28983,N_24504,N_24868);
and U28984 (N_28984,N_26698,N_25736);
nor U28985 (N_28985,N_25000,N_26966);
nand U28986 (N_28986,N_24832,N_26156);
nand U28987 (N_28987,N_25585,N_25676);
xnor U28988 (N_28988,N_25726,N_25173);
nor U28989 (N_28989,N_24523,N_24738);
nor U28990 (N_28990,N_26504,N_24436);
and U28991 (N_28991,N_24547,N_26877);
xnor U28992 (N_28992,N_24886,N_25594);
nand U28993 (N_28993,N_24850,N_24708);
xnor U28994 (N_28994,N_25348,N_26264);
nor U28995 (N_28995,N_24780,N_24675);
or U28996 (N_28996,N_26142,N_26847);
or U28997 (N_28997,N_24021,N_24809);
nand U28998 (N_28998,N_24502,N_25454);
or U28999 (N_28999,N_26806,N_24664);
xor U29000 (N_29000,N_25590,N_26305);
or U29001 (N_29001,N_25935,N_26227);
or U29002 (N_29002,N_24545,N_26299);
xnor U29003 (N_29003,N_26598,N_25736);
nand U29004 (N_29004,N_24582,N_24842);
or U29005 (N_29005,N_24716,N_25099);
nand U29006 (N_29006,N_26739,N_24525);
and U29007 (N_29007,N_25631,N_26972);
xnor U29008 (N_29008,N_25235,N_26472);
nand U29009 (N_29009,N_26484,N_24612);
nand U29010 (N_29010,N_26459,N_24609);
nor U29011 (N_29011,N_24033,N_26864);
and U29012 (N_29012,N_26095,N_25907);
nor U29013 (N_29013,N_26467,N_24064);
xnor U29014 (N_29014,N_24368,N_25636);
or U29015 (N_29015,N_26755,N_24304);
nand U29016 (N_29016,N_24923,N_25645);
and U29017 (N_29017,N_24672,N_25460);
nor U29018 (N_29018,N_26086,N_26612);
nor U29019 (N_29019,N_26761,N_24943);
and U29020 (N_29020,N_26690,N_25625);
nand U29021 (N_29021,N_25423,N_26738);
and U29022 (N_29022,N_24220,N_25039);
and U29023 (N_29023,N_26542,N_25956);
or U29024 (N_29024,N_24493,N_25567);
and U29025 (N_29025,N_26759,N_24398);
xnor U29026 (N_29026,N_26986,N_25337);
xor U29027 (N_29027,N_25558,N_25399);
or U29028 (N_29028,N_24732,N_26205);
or U29029 (N_29029,N_24727,N_26210);
xnor U29030 (N_29030,N_24135,N_25963);
or U29031 (N_29031,N_25965,N_25987);
xnor U29032 (N_29032,N_26536,N_26947);
or U29033 (N_29033,N_26719,N_25703);
and U29034 (N_29034,N_26767,N_24631);
or U29035 (N_29035,N_26216,N_26441);
and U29036 (N_29036,N_24575,N_26344);
xnor U29037 (N_29037,N_26623,N_25340);
nand U29038 (N_29038,N_25798,N_24814);
and U29039 (N_29039,N_24367,N_26331);
or U29040 (N_29040,N_24799,N_25954);
xor U29041 (N_29041,N_26703,N_25365);
or U29042 (N_29042,N_25311,N_24100);
xor U29043 (N_29043,N_25220,N_26578);
and U29044 (N_29044,N_25475,N_26010);
xor U29045 (N_29045,N_25272,N_26899);
nand U29046 (N_29046,N_26233,N_25362);
or U29047 (N_29047,N_24668,N_26084);
xor U29048 (N_29048,N_26363,N_25092);
xor U29049 (N_29049,N_25102,N_26363);
or U29050 (N_29050,N_25617,N_25569);
nor U29051 (N_29051,N_25456,N_24577);
nor U29052 (N_29052,N_26236,N_26954);
and U29053 (N_29053,N_24003,N_25140);
nand U29054 (N_29054,N_25606,N_24253);
xnor U29055 (N_29055,N_24185,N_24212);
nor U29056 (N_29056,N_25489,N_26321);
and U29057 (N_29057,N_26543,N_25893);
and U29058 (N_29058,N_24263,N_24005);
or U29059 (N_29059,N_24720,N_25380);
and U29060 (N_29060,N_25507,N_26595);
nand U29061 (N_29061,N_24518,N_24000);
or U29062 (N_29062,N_25107,N_26583);
nor U29063 (N_29063,N_26001,N_24774);
and U29064 (N_29064,N_26584,N_26041);
nand U29065 (N_29065,N_25053,N_24360);
xnor U29066 (N_29066,N_26357,N_25595);
nand U29067 (N_29067,N_26169,N_24211);
nand U29068 (N_29068,N_26340,N_25111);
and U29069 (N_29069,N_25726,N_26482);
and U29070 (N_29070,N_25621,N_26179);
and U29071 (N_29071,N_26386,N_26670);
nor U29072 (N_29072,N_26172,N_25173);
or U29073 (N_29073,N_25207,N_25660);
or U29074 (N_29074,N_24536,N_25032);
nor U29075 (N_29075,N_26586,N_25960);
or U29076 (N_29076,N_25287,N_25071);
nor U29077 (N_29077,N_25993,N_26866);
nand U29078 (N_29078,N_25473,N_26118);
or U29079 (N_29079,N_26990,N_25476);
nand U29080 (N_29080,N_26944,N_26530);
or U29081 (N_29081,N_25344,N_25291);
xnor U29082 (N_29082,N_25807,N_26893);
nand U29083 (N_29083,N_24581,N_26042);
xnor U29084 (N_29084,N_26440,N_26205);
and U29085 (N_29085,N_24353,N_25759);
and U29086 (N_29086,N_24824,N_26960);
nand U29087 (N_29087,N_26832,N_24464);
or U29088 (N_29088,N_24728,N_24310);
and U29089 (N_29089,N_24899,N_24995);
nor U29090 (N_29090,N_25298,N_25447);
or U29091 (N_29091,N_25295,N_25126);
or U29092 (N_29092,N_24954,N_24911);
nand U29093 (N_29093,N_25834,N_26152);
and U29094 (N_29094,N_24617,N_24964);
and U29095 (N_29095,N_25939,N_24011);
or U29096 (N_29096,N_24676,N_25463);
or U29097 (N_29097,N_25698,N_24529);
and U29098 (N_29098,N_25802,N_25706);
nor U29099 (N_29099,N_25318,N_24923);
or U29100 (N_29100,N_25913,N_24534);
or U29101 (N_29101,N_26956,N_26136);
and U29102 (N_29102,N_25944,N_26399);
and U29103 (N_29103,N_26703,N_26121);
xor U29104 (N_29104,N_26176,N_24152);
and U29105 (N_29105,N_25211,N_25373);
and U29106 (N_29106,N_26177,N_24370);
or U29107 (N_29107,N_26324,N_24818);
nor U29108 (N_29108,N_24928,N_25964);
xnor U29109 (N_29109,N_26397,N_26138);
or U29110 (N_29110,N_26036,N_24125);
xnor U29111 (N_29111,N_26912,N_25125);
nand U29112 (N_29112,N_25556,N_25191);
nand U29113 (N_29113,N_24821,N_25709);
xor U29114 (N_29114,N_24371,N_25927);
nor U29115 (N_29115,N_24384,N_26393);
or U29116 (N_29116,N_26897,N_24110);
xnor U29117 (N_29117,N_26443,N_26717);
nor U29118 (N_29118,N_24492,N_25915);
nand U29119 (N_29119,N_24834,N_26145);
xor U29120 (N_29120,N_24904,N_25937);
xnor U29121 (N_29121,N_25967,N_24257);
nand U29122 (N_29122,N_25917,N_26529);
nor U29123 (N_29123,N_24275,N_26423);
and U29124 (N_29124,N_26396,N_24358);
and U29125 (N_29125,N_24179,N_26210);
and U29126 (N_29126,N_26815,N_25777);
and U29127 (N_29127,N_25877,N_25744);
or U29128 (N_29128,N_26697,N_24010);
xor U29129 (N_29129,N_26842,N_25739);
nand U29130 (N_29130,N_26925,N_25737);
and U29131 (N_29131,N_24434,N_25030);
nand U29132 (N_29132,N_24240,N_25256);
xor U29133 (N_29133,N_24076,N_24957);
nor U29134 (N_29134,N_24271,N_24269);
or U29135 (N_29135,N_26717,N_24289);
or U29136 (N_29136,N_26020,N_26084);
nand U29137 (N_29137,N_24244,N_24704);
nor U29138 (N_29138,N_25152,N_25689);
xor U29139 (N_29139,N_25397,N_26623);
and U29140 (N_29140,N_24005,N_24733);
or U29141 (N_29141,N_25657,N_24894);
nand U29142 (N_29142,N_25813,N_25560);
xor U29143 (N_29143,N_26027,N_24850);
or U29144 (N_29144,N_25844,N_25980);
nor U29145 (N_29145,N_25339,N_26903);
nor U29146 (N_29146,N_26243,N_26329);
and U29147 (N_29147,N_26050,N_24746);
nand U29148 (N_29148,N_26532,N_25348);
nor U29149 (N_29149,N_25138,N_25786);
nand U29150 (N_29150,N_24501,N_24917);
or U29151 (N_29151,N_24857,N_26628);
nor U29152 (N_29152,N_24414,N_25189);
or U29153 (N_29153,N_24550,N_24644);
xnor U29154 (N_29154,N_24165,N_25761);
nand U29155 (N_29155,N_25773,N_26767);
or U29156 (N_29156,N_25087,N_26619);
or U29157 (N_29157,N_24396,N_26366);
nand U29158 (N_29158,N_25817,N_26826);
nand U29159 (N_29159,N_25509,N_25185);
and U29160 (N_29160,N_25312,N_25501);
and U29161 (N_29161,N_25705,N_24753);
nand U29162 (N_29162,N_24430,N_26896);
nand U29163 (N_29163,N_26729,N_25249);
or U29164 (N_29164,N_25559,N_25662);
xor U29165 (N_29165,N_25744,N_24322);
xnor U29166 (N_29166,N_26369,N_24004);
xnor U29167 (N_29167,N_25961,N_25196);
xnor U29168 (N_29168,N_26867,N_24922);
or U29169 (N_29169,N_24375,N_24200);
nor U29170 (N_29170,N_24118,N_25827);
nand U29171 (N_29171,N_26410,N_24218);
or U29172 (N_29172,N_25216,N_25125);
and U29173 (N_29173,N_26689,N_25351);
or U29174 (N_29174,N_26599,N_25939);
nand U29175 (N_29175,N_25709,N_26330);
nor U29176 (N_29176,N_26585,N_24415);
nand U29177 (N_29177,N_25118,N_26038);
or U29178 (N_29178,N_24122,N_25319);
nand U29179 (N_29179,N_24366,N_24848);
nor U29180 (N_29180,N_26148,N_25515);
and U29181 (N_29181,N_24319,N_25537);
and U29182 (N_29182,N_24916,N_25583);
xor U29183 (N_29183,N_26126,N_24934);
xnor U29184 (N_29184,N_24185,N_24199);
and U29185 (N_29185,N_25235,N_25658);
nand U29186 (N_29186,N_25645,N_24739);
and U29187 (N_29187,N_25922,N_26488);
nand U29188 (N_29188,N_24275,N_24209);
nand U29189 (N_29189,N_25894,N_26727);
nor U29190 (N_29190,N_25671,N_24936);
nand U29191 (N_29191,N_26708,N_25808);
nor U29192 (N_29192,N_26641,N_25030);
nand U29193 (N_29193,N_24418,N_24220);
and U29194 (N_29194,N_24969,N_24995);
nand U29195 (N_29195,N_24938,N_26661);
nor U29196 (N_29196,N_26826,N_25728);
xnor U29197 (N_29197,N_24221,N_26750);
nor U29198 (N_29198,N_26477,N_26628);
or U29199 (N_29199,N_26884,N_24205);
xor U29200 (N_29200,N_25888,N_25098);
and U29201 (N_29201,N_25412,N_24243);
nor U29202 (N_29202,N_25000,N_24909);
nand U29203 (N_29203,N_26717,N_26767);
and U29204 (N_29204,N_25826,N_26292);
xor U29205 (N_29205,N_26921,N_24510);
nor U29206 (N_29206,N_24964,N_24331);
or U29207 (N_29207,N_24157,N_25755);
xor U29208 (N_29208,N_26976,N_24521);
nand U29209 (N_29209,N_26452,N_24070);
and U29210 (N_29210,N_26362,N_26084);
xor U29211 (N_29211,N_26876,N_26618);
and U29212 (N_29212,N_25303,N_26480);
nand U29213 (N_29213,N_25580,N_25775);
and U29214 (N_29214,N_25365,N_26886);
or U29215 (N_29215,N_26722,N_24894);
and U29216 (N_29216,N_25897,N_26113);
or U29217 (N_29217,N_24507,N_24056);
nand U29218 (N_29218,N_25685,N_26801);
nand U29219 (N_29219,N_25251,N_25452);
xnor U29220 (N_29220,N_26371,N_25596);
nor U29221 (N_29221,N_25090,N_24270);
xor U29222 (N_29222,N_26186,N_26467);
xor U29223 (N_29223,N_25681,N_25267);
and U29224 (N_29224,N_26320,N_25385);
xor U29225 (N_29225,N_26345,N_26963);
nand U29226 (N_29226,N_25277,N_26001);
xor U29227 (N_29227,N_26319,N_25901);
nor U29228 (N_29228,N_25190,N_24812);
xnor U29229 (N_29229,N_24012,N_25461);
and U29230 (N_29230,N_25095,N_25603);
and U29231 (N_29231,N_24536,N_25783);
nor U29232 (N_29232,N_26667,N_25909);
nor U29233 (N_29233,N_26291,N_24593);
and U29234 (N_29234,N_26004,N_25118);
and U29235 (N_29235,N_24068,N_24345);
nand U29236 (N_29236,N_25779,N_25643);
xor U29237 (N_29237,N_25321,N_26235);
nor U29238 (N_29238,N_24995,N_25768);
nand U29239 (N_29239,N_25001,N_26221);
nand U29240 (N_29240,N_26975,N_26769);
nand U29241 (N_29241,N_26701,N_25782);
or U29242 (N_29242,N_24876,N_26796);
nand U29243 (N_29243,N_26901,N_26011);
nor U29244 (N_29244,N_25968,N_24012);
or U29245 (N_29245,N_25837,N_25174);
nor U29246 (N_29246,N_26571,N_25442);
nor U29247 (N_29247,N_24318,N_24490);
nor U29248 (N_29248,N_24550,N_24945);
and U29249 (N_29249,N_25979,N_26436);
nor U29250 (N_29250,N_24578,N_25785);
nor U29251 (N_29251,N_25480,N_26261);
xnor U29252 (N_29252,N_24186,N_26704);
xor U29253 (N_29253,N_25607,N_25876);
xor U29254 (N_29254,N_25467,N_25648);
nor U29255 (N_29255,N_26548,N_24272);
and U29256 (N_29256,N_25334,N_24757);
xor U29257 (N_29257,N_25258,N_24911);
or U29258 (N_29258,N_24899,N_24532);
or U29259 (N_29259,N_25944,N_26742);
nor U29260 (N_29260,N_25472,N_25148);
or U29261 (N_29261,N_24980,N_26333);
nand U29262 (N_29262,N_25456,N_24546);
xnor U29263 (N_29263,N_24344,N_26502);
nor U29264 (N_29264,N_26285,N_25702);
nand U29265 (N_29265,N_26019,N_26805);
nand U29266 (N_29266,N_24358,N_25778);
xnor U29267 (N_29267,N_25235,N_24655);
nor U29268 (N_29268,N_25614,N_25558);
nor U29269 (N_29269,N_24658,N_24426);
nor U29270 (N_29270,N_24590,N_26601);
nand U29271 (N_29271,N_26532,N_24984);
or U29272 (N_29272,N_26874,N_25555);
nand U29273 (N_29273,N_24476,N_26991);
xnor U29274 (N_29274,N_26609,N_24746);
nor U29275 (N_29275,N_26085,N_24619);
nor U29276 (N_29276,N_26681,N_26616);
or U29277 (N_29277,N_24212,N_26142);
and U29278 (N_29278,N_26068,N_24628);
nor U29279 (N_29279,N_25310,N_25215);
or U29280 (N_29280,N_24537,N_24285);
or U29281 (N_29281,N_26291,N_25481);
xnor U29282 (N_29282,N_25342,N_25024);
xor U29283 (N_29283,N_25883,N_26237);
nor U29284 (N_29284,N_25539,N_26585);
xor U29285 (N_29285,N_24599,N_25260);
or U29286 (N_29286,N_25417,N_26655);
xnor U29287 (N_29287,N_24664,N_25467);
or U29288 (N_29288,N_24021,N_24257);
or U29289 (N_29289,N_25696,N_24765);
nor U29290 (N_29290,N_25748,N_24898);
nor U29291 (N_29291,N_24328,N_25477);
or U29292 (N_29292,N_25015,N_24123);
or U29293 (N_29293,N_26041,N_25700);
xor U29294 (N_29294,N_25813,N_24157);
or U29295 (N_29295,N_26087,N_24569);
nor U29296 (N_29296,N_26521,N_25349);
nand U29297 (N_29297,N_25864,N_24711);
and U29298 (N_29298,N_24853,N_24926);
or U29299 (N_29299,N_26280,N_24771);
nor U29300 (N_29300,N_24724,N_25458);
xor U29301 (N_29301,N_26218,N_25813);
or U29302 (N_29302,N_24143,N_24340);
nor U29303 (N_29303,N_25313,N_26513);
xnor U29304 (N_29304,N_26283,N_25985);
nor U29305 (N_29305,N_24644,N_26212);
xnor U29306 (N_29306,N_26893,N_25180);
or U29307 (N_29307,N_24620,N_25758);
and U29308 (N_29308,N_24220,N_26208);
nor U29309 (N_29309,N_26073,N_25660);
nand U29310 (N_29310,N_24046,N_25909);
or U29311 (N_29311,N_25796,N_26954);
or U29312 (N_29312,N_25042,N_24725);
nor U29313 (N_29313,N_24384,N_25477);
and U29314 (N_29314,N_25778,N_25330);
and U29315 (N_29315,N_26883,N_24903);
nor U29316 (N_29316,N_25054,N_24239);
or U29317 (N_29317,N_24766,N_24774);
xor U29318 (N_29318,N_24607,N_25384);
and U29319 (N_29319,N_24751,N_26260);
and U29320 (N_29320,N_25308,N_24649);
or U29321 (N_29321,N_25690,N_24407);
or U29322 (N_29322,N_26355,N_25474);
nor U29323 (N_29323,N_26011,N_24152);
and U29324 (N_29324,N_26565,N_26648);
nand U29325 (N_29325,N_26462,N_26145);
nor U29326 (N_29326,N_25471,N_26907);
nand U29327 (N_29327,N_25534,N_26876);
and U29328 (N_29328,N_26213,N_25178);
or U29329 (N_29329,N_26737,N_24260);
and U29330 (N_29330,N_24828,N_24500);
and U29331 (N_29331,N_24963,N_24447);
xnor U29332 (N_29332,N_25298,N_26996);
nor U29333 (N_29333,N_25620,N_24620);
xor U29334 (N_29334,N_24543,N_25399);
and U29335 (N_29335,N_26289,N_24581);
and U29336 (N_29336,N_25925,N_26860);
or U29337 (N_29337,N_26152,N_26704);
xnor U29338 (N_29338,N_24907,N_24946);
xor U29339 (N_29339,N_26191,N_24407);
nor U29340 (N_29340,N_24626,N_25348);
or U29341 (N_29341,N_26715,N_25063);
or U29342 (N_29342,N_25270,N_26508);
or U29343 (N_29343,N_25246,N_25102);
nand U29344 (N_29344,N_24561,N_24901);
or U29345 (N_29345,N_24709,N_25142);
nand U29346 (N_29346,N_25506,N_25127);
nand U29347 (N_29347,N_25942,N_24577);
nor U29348 (N_29348,N_26298,N_26941);
nand U29349 (N_29349,N_25372,N_24320);
xnor U29350 (N_29350,N_26462,N_26805);
nand U29351 (N_29351,N_26579,N_25273);
nand U29352 (N_29352,N_24394,N_26408);
nor U29353 (N_29353,N_26679,N_26456);
nor U29354 (N_29354,N_25198,N_25614);
or U29355 (N_29355,N_24965,N_26782);
or U29356 (N_29356,N_25933,N_25806);
or U29357 (N_29357,N_24772,N_26239);
and U29358 (N_29358,N_25708,N_24688);
xor U29359 (N_29359,N_26605,N_26590);
nor U29360 (N_29360,N_26497,N_24124);
nor U29361 (N_29361,N_25529,N_25357);
or U29362 (N_29362,N_26178,N_24680);
and U29363 (N_29363,N_25618,N_26437);
or U29364 (N_29364,N_26000,N_25610);
and U29365 (N_29365,N_24672,N_26176);
nor U29366 (N_29366,N_24175,N_26725);
and U29367 (N_29367,N_25452,N_24977);
and U29368 (N_29368,N_24735,N_25747);
nand U29369 (N_29369,N_24354,N_26258);
or U29370 (N_29370,N_25914,N_25824);
nand U29371 (N_29371,N_25002,N_24949);
nand U29372 (N_29372,N_25032,N_25515);
nor U29373 (N_29373,N_24530,N_24920);
or U29374 (N_29374,N_24682,N_25337);
nand U29375 (N_29375,N_25179,N_26138);
and U29376 (N_29376,N_26701,N_26900);
nor U29377 (N_29377,N_26853,N_25133);
nand U29378 (N_29378,N_26448,N_26424);
and U29379 (N_29379,N_25719,N_25032);
or U29380 (N_29380,N_24860,N_25758);
and U29381 (N_29381,N_26994,N_24178);
or U29382 (N_29382,N_26936,N_25167);
or U29383 (N_29383,N_25704,N_26387);
and U29384 (N_29384,N_25843,N_26204);
nand U29385 (N_29385,N_24809,N_24530);
or U29386 (N_29386,N_26622,N_25585);
and U29387 (N_29387,N_25027,N_24427);
nand U29388 (N_29388,N_26800,N_26094);
and U29389 (N_29389,N_26009,N_26530);
and U29390 (N_29390,N_26456,N_25747);
nand U29391 (N_29391,N_24425,N_25987);
nand U29392 (N_29392,N_26300,N_26112);
and U29393 (N_29393,N_26496,N_24352);
and U29394 (N_29394,N_26358,N_24492);
xnor U29395 (N_29395,N_25027,N_26015);
nand U29396 (N_29396,N_24837,N_25061);
or U29397 (N_29397,N_24973,N_26375);
nor U29398 (N_29398,N_25179,N_24390);
and U29399 (N_29399,N_26142,N_24979);
xor U29400 (N_29400,N_25167,N_25727);
or U29401 (N_29401,N_25435,N_24200);
xnor U29402 (N_29402,N_26140,N_26250);
nand U29403 (N_29403,N_25072,N_25674);
nor U29404 (N_29404,N_24609,N_24666);
and U29405 (N_29405,N_24552,N_25234);
or U29406 (N_29406,N_24345,N_25480);
nor U29407 (N_29407,N_26069,N_24422);
nor U29408 (N_29408,N_26257,N_25496);
nor U29409 (N_29409,N_25460,N_26703);
nor U29410 (N_29410,N_25771,N_25301);
xor U29411 (N_29411,N_24143,N_24270);
or U29412 (N_29412,N_26978,N_24135);
nand U29413 (N_29413,N_24764,N_25849);
or U29414 (N_29414,N_24410,N_26222);
nand U29415 (N_29415,N_24602,N_24939);
xor U29416 (N_29416,N_25376,N_26788);
xnor U29417 (N_29417,N_25894,N_24647);
and U29418 (N_29418,N_24220,N_26797);
or U29419 (N_29419,N_24192,N_24263);
xnor U29420 (N_29420,N_26153,N_25302);
and U29421 (N_29421,N_24930,N_25892);
or U29422 (N_29422,N_24048,N_25079);
nor U29423 (N_29423,N_24936,N_26546);
nand U29424 (N_29424,N_25855,N_26743);
nor U29425 (N_29425,N_24338,N_25535);
xnor U29426 (N_29426,N_24460,N_26451);
or U29427 (N_29427,N_24656,N_25194);
xor U29428 (N_29428,N_24746,N_25823);
nor U29429 (N_29429,N_24641,N_25749);
and U29430 (N_29430,N_25552,N_24827);
and U29431 (N_29431,N_24993,N_24840);
nand U29432 (N_29432,N_25106,N_26094);
nand U29433 (N_29433,N_26682,N_25494);
nand U29434 (N_29434,N_24649,N_26996);
nor U29435 (N_29435,N_24203,N_26972);
or U29436 (N_29436,N_25387,N_26857);
or U29437 (N_29437,N_25374,N_24181);
or U29438 (N_29438,N_24015,N_25494);
xor U29439 (N_29439,N_25611,N_24007);
nand U29440 (N_29440,N_25952,N_24457);
and U29441 (N_29441,N_24305,N_24061);
nor U29442 (N_29442,N_26678,N_25434);
nand U29443 (N_29443,N_26503,N_24647);
or U29444 (N_29444,N_24696,N_25980);
nand U29445 (N_29445,N_24549,N_26565);
xor U29446 (N_29446,N_25600,N_25630);
nor U29447 (N_29447,N_25491,N_25767);
nand U29448 (N_29448,N_26140,N_25042);
nor U29449 (N_29449,N_25772,N_25095);
nor U29450 (N_29450,N_26036,N_25250);
nor U29451 (N_29451,N_24655,N_26877);
and U29452 (N_29452,N_25126,N_26284);
or U29453 (N_29453,N_24863,N_24234);
and U29454 (N_29454,N_26572,N_26262);
xnor U29455 (N_29455,N_24146,N_26413);
and U29456 (N_29456,N_25925,N_26971);
and U29457 (N_29457,N_26397,N_26017);
or U29458 (N_29458,N_26048,N_25039);
and U29459 (N_29459,N_25553,N_24369);
nor U29460 (N_29460,N_26087,N_25230);
nor U29461 (N_29461,N_24375,N_24827);
or U29462 (N_29462,N_26650,N_25283);
nand U29463 (N_29463,N_24328,N_24294);
xor U29464 (N_29464,N_26401,N_24939);
nand U29465 (N_29465,N_25592,N_24571);
or U29466 (N_29466,N_26677,N_26493);
nor U29467 (N_29467,N_26960,N_25554);
nor U29468 (N_29468,N_24191,N_24434);
nand U29469 (N_29469,N_24900,N_26202);
nor U29470 (N_29470,N_25109,N_26860);
or U29471 (N_29471,N_24959,N_26277);
nor U29472 (N_29472,N_24867,N_25664);
nand U29473 (N_29473,N_26530,N_25465);
and U29474 (N_29474,N_25039,N_26343);
and U29475 (N_29475,N_25075,N_26523);
xor U29476 (N_29476,N_25692,N_24283);
and U29477 (N_29477,N_25941,N_26594);
and U29478 (N_29478,N_24123,N_24503);
nand U29479 (N_29479,N_26982,N_24841);
or U29480 (N_29480,N_24439,N_24121);
nor U29481 (N_29481,N_24544,N_26257);
nor U29482 (N_29482,N_25366,N_26577);
and U29483 (N_29483,N_25158,N_24552);
nand U29484 (N_29484,N_24934,N_25357);
nor U29485 (N_29485,N_24937,N_25069);
and U29486 (N_29486,N_25507,N_24296);
or U29487 (N_29487,N_26956,N_26429);
nor U29488 (N_29488,N_24674,N_25647);
and U29489 (N_29489,N_24640,N_26050);
xnor U29490 (N_29490,N_26832,N_25786);
nor U29491 (N_29491,N_26641,N_25436);
nor U29492 (N_29492,N_24468,N_25465);
and U29493 (N_29493,N_26915,N_26889);
or U29494 (N_29494,N_25909,N_24744);
xor U29495 (N_29495,N_25054,N_24397);
nor U29496 (N_29496,N_24098,N_24523);
nor U29497 (N_29497,N_25725,N_24552);
nand U29498 (N_29498,N_25720,N_24500);
or U29499 (N_29499,N_26393,N_26931);
and U29500 (N_29500,N_25654,N_24235);
or U29501 (N_29501,N_24484,N_25003);
or U29502 (N_29502,N_24646,N_24172);
and U29503 (N_29503,N_25596,N_25546);
nand U29504 (N_29504,N_24582,N_26788);
nor U29505 (N_29505,N_25423,N_25375);
or U29506 (N_29506,N_25148,N_24240);
or U29507 (N_29507,N_24811,N_26951);
xor U29508 (N_29508,N_24424,N_24333);
nand U29509 (N_29509,N_24495,N_26424);
nand U29510 (N_29510,N_26869,N_26848);
or U29511 (N_29511,N_25021,N_26501);
nor U29512 (N_29512,N_24898,N_24596);
or U29513 (N_29513,N_26285,N_24155);
nand U29514 (N_29514,N_26640,N_26661);
nand U29515 (N_29515,N_25846,N_26249);
nand U29516 (N_29516,N_26478,N_25483);
xor U29517 (N_29517,N_25249,N_26447);
and U29518 (N_29518,N_25070,N_24690);
and U29519 (N_29519,N_26448,N_25470);
nand U29520 (N_29520,N_26832,N_26404);
nor U29521 (N_29521,N_24627,N_25759);
nand U29522 (N_29522,N_25651,N_26601);
xor U29523 (N_29523,N_26004,N_25936);
and U29524 (N_29524,N_24366,N_26852);
xnor U29525 (N_29525,N_26301,N_24699);
xor U29526 (N_29526,N_26470,N_25956);
nor U29527 (N_29527,N_24032,N_24771);
and U29528 (N_29528,N_24490,N_24150);
nor U29529 (N_29529,N_24854,N_25546);
and U29530 (N_29530,N_26610,N_25973);
or U29531 (N_29531,N_26066,N_26385);
and U29532 (N_29532,N_26186,N_24068);
xor U29533 (N_29533,N_25634,N_25636);
or U29534 (N_29534,N_24818,N_24729);
nor U29535 (N_29535,N_26057,N_25232);
nor U29536 (N_29536,N_25625,N_26937);
nand U29537 (N_29537,N_25731,N_25931);
nor U29538 (N_29538,N_25200,N_25785);
or U29539 (N_29539,N_25264,N_26510);
or U29540 (N_29540,N_26078,N_24920);
xor U29541 (N_29541,N_26334,N_25087);
nand U29542 (N_29542,N_26700,N_25374);
and U29543 (N_29543,N_25320,N_25232);
nand U29544 (N_29544,N_26477,N_24788);
and U29545 (N_29545,N_24432,N_26238);
and U29546 (N_29546,N_25886,N_24190);
nor U29547 (N_29547,N_26137,N_26766);
nand U29548 (N_29548,N_24066,N_25694);
or U29549 (N_29549,N_26478,N_26623);
nor U29550 (N_29550,N_25537,N_24650);
or U29551 (N_29551,N_25944,N_26194);
xnor U29552 (N_29552,N_25731,N_26666);
nand U29553 (N_29553,N_26782,N_26405);
or U29554 (N_29554,N_25488,N_24569);
nor U29555 (N_29555,N_24809,N_25615);
nor U29556 (N_29556,N_25926,N_26289);
and U29557 (N_29557,N_25907,N_24522);
and U29558 (N_29558,N_24398,N_24313);
or U29559 (N_29559,N_26961,N_25998);
nor U29560 (N_29560,N_26687,N_24986);
nor U29561 (N_29561,N_26510,N_25667);
nand U29562 (N_29562,N_25229,N_26992);
and U29563 (N_29563,N_26633,N_25251);
nand U29564 (N_29564,N_26039,N_24641);
or U29565 (N_29565,N_25918,N_26200);
nor U29566 (N_29566,N_25014,N_26370);
nor U29567 (N_29567,N_25772,N_26806);
nand U29568 (N_29568,N_26486,N_24560);
xor U29569 (N_29569,N_25049,N_25026);
nand U29570 (N_29570,N_26210,N_26275);
or U29571 (N_29571,N_26901,N_26110);
xnor U29572 (N_29572,N_25833,N_24345);
xnor U29573 (N_29573,N_26456,N_24437);
xor U29574 (N_29574,N_26462,N_25117);
or U29575 (N_29575,N_26553,N_26336);
nand U29576 (N_29576,N_26423,N_26242);
xnor U29577 (N_29577,N_24767,N_24791);
nor U29578 (N_29578,N_25870,N_25717);
xor U29579 (N_29579,N_26466,N_24950);
nor U29580 (N_29580,N_25810,N_24488);
xor U29581 (N_29581,N_24612,N_25174);
nand U29582 (N_29582,N_25230,N_26435);
xnor U29583 (N_29583,N_24100,N_26197);
or U29584 (N_29584,N_24288,N_25139);
xnor U29585 (N_29585,N_25816,N_24453);
or U29586 (N_29586,N_24983,N_25725);
nand U29587 (N_29587,N_26469,N_26370);
nor U29588 (N_29588,N_25507,N_25325);
nand U29589 (N_29589,N_24415,N_25424);
nand U29590 (N_29590,N_26964,N_25572);
nor U29591 (N_29591,N_24242,N_24790);
nand U29592 (N_29592,N_24564,N_24810);
nor U29593 (N_29593,N_24559,N_24790);
xor U29594 (N_29594,N_24431,N_25505);
nor U29595 (N_29595,N_26571,N_25043);
nand U29596 (N_29596,N_24178,N_24196);
xnor U29597 (N_29597,N_26394,N_25263);
nand U29598 (N_29598,N_24889,N_26650);
nand U29599 (N_29599,N_24262,N_24855);
xnor U29600 (N_29600,N_26794,N_24771);
or U29601 (N_29601,N_24015,N_26737);
nand U29602 (N_29602,N_26165,N_26458);
nand U29603 (N_29603,N_25290,N_26735);
or U29604 (N_29604,N_26334,N_24530);
xnor U29605 (N_29605,N_24351,N_26347);
nand U29606 (N_29606,N_24529,N_24599);
nand U29607 (N_29607,N_26940,N_26667);
nand U29608 (N_29608,N_24908,N_25172);
nor U29609 (N_29609,N_24287,N_25465);
nor U29610 (N_29610,N_26522,N_24755);
nand U29611 (N_29611,N_24159,N_25034);
nor U29612 (N_29612,N_26601,N_24121);
nand U29613 (N_29613,N_24541,N_26297);
xnor U29614 (N_29614,N_26686,N_26581);
xnor U29615 (N_29615,N_25591,N_26391);
nand U29616 (N_29616,N_25989,N_24324);
nor U29617 (N_29617,N_26671,N_25718);
nor U29618 (N_29618,N_25546,N_25173);
or U29619 (N_29619,N_26123,N_24314);
nand U29620 (N_29620,N_24137,N_25260);
nand U29621 (N_29621,N_24420,N_26784);
and U29622 (N_29622,N_24145,N_24021);
nand U29623 (N_29623,N_25789,N_26720);
and U29624 (N_29624,N_25518,N_24841);
nor U29625 (N_29625,N_26365,N_24362);
or U29626 (N_29626,N_24171,N_24802);
xnor U29627 (N_29627,N_26963,N_26878);
nand U29628 (N_29628,N_26569,N_25212);
nor U29629 (N_29629,N_24980,N_24313);
xor U29630 (N_29630,N_26243,N_24832);
nor U29631 (N_29631,N_25734,N_26616);
nor U29632 (N_29632,N_25053,N_25951);
xnor U29633 (N_29633,N_26411,N_24641);
nand U29634 (N_29634,N_25857,N_25328);
nand U29635 (N_29635,N_24089,N_25844);
and U29636 (N_29636,N_25529,N_26789);
nand U29637 (N_29637,N_25753,N_25349);
nor U29638 (N_29638,N_25087,N_25904);
or U29639 (N_29639,N_25699,N_24623);
nand U29640 (N_29640,N_24704,N_25069);
and U29641 (N_29641,N_26644,N_26698);
xor U29642 (N_29642,N_26299,N_25277);
or U29643 (N_29643,N_24686,N_24909);
nand U29644 (N_29644,N_24504,N_24199);
nand U29645 (N_29645,N_26373,N_25892);
xor U29646 (N_29646,N_24503,N_25296);
xor U29647 (N_29647,N_24143,N_26144);
nand U29648 (N_29648,N_25317,N_26263);
or U29649 (N_29649,N_25306,N_24049);
or U29650 (N_29650,N_25946,N_24537);
and U29651 (N_29651,N_24268,N_26461);
nor U29652 (N_29652,N_25491,N_25708);
and U29653 (N_29653,N_24716,N_25541);
nor U29654 (N_29654,N_24220,N_25923);
nand U29655 (N_29655,N_25818,N_26370);
nand U29656 (N_29656,N_25858,N_26170);
and U29657 (N_29657,N_26147,N_24624);
xnor U29658 (N_29658,N_26268,N_25139);
nand U29659 (N_29659,N_24618,N_24864);
or U29660 (N_29660,N_25155,N_26080);
xor U29661 (N_29661,N_24693,N_26319);
and U29662 (N_29662,N_24361,N_26589);
nand U29663 (N_29663,N_26023,N_25492);
and U29664 (N_29664,N_26951,N_24791);
nand U29665 (N_29665,N_26149,N_24177);
nand U29666 (N_29666,N_24826,N_24569);
nor U29667 (N_29667,N_24030,N_24535);
nand U29668 (N_29668,N_24594,N_26874);
xor U29669 (N_29669,N_24560,N_25917);
nor U29670 (N_29670,N_25742,N_25471);
nor U29671 (N_29671,N_24489,N_25090);
nor U29672 (N_29672,N_25481,N_24611);
xor U29673 (N_29673,N_24849,N_24521);
xor U29674 (N_29674,N_26940,N_25713);
and U29675 (N_29675,N_24011,N_24040);
xnor U29676 (N_29676,N_26396,N_25358);
and U29677 (N_29677,N_24039,N_24281);
nand U29678 (N_29678,N_26499,N_26805);
or U29679 (N_29679,N_24669,N_24423);
nand U29680 (N_29680,N_25927,N_24496);
xor U29681 (N_29681,N_26109,N_24315);
and U29682 (N_29682,N_26618,N_26770);
or U29683 (N_29683,N_26038,N_26772);
xor U29684 (N_29684,N_24336,N_24646);
nand U29685 (N_29685,N_24967,N_24290);
nand U29686 (N_29686,N_26353,N_25277);
nand U29687 (N_29687,N_26726,N_25220);
nand U29688 (N_29688,N_24663,N_26539);
and U29689 (N_29689,N_25974,N_26231);
nor U29690 (N_29690,N_24407,N_25622);
nor U29691 (N_29691,N_24930,N_24514);
xor U29692 (N_29692,N_25934,N_25587);
or U29693 (N_29693,N_25440,N_24664);
or U29694 (N_29694,N_26544,N_24021);
or U29695 (N_29695,N_25079,N_26680);
nor U29696 (N_29696,N_25901,N_26561);
nand U29697 (N_29697,N_26601,N_24181);
or U29698 (N_29698,N_24875,N_26702);
nor U29699 (N_29699,N_26140,N_24864);
nor U29700 (N_29700,N_24627,N_24421);
nand U29701 (N_29701,N_24948,N_25997);
xor U29702 (N_29702,N_24603,N_26722);
xor U29703 (N_29703,N_25321,N_26360);
nand U29704 (N_29704,N_24387,N_24426);
and U29705 (N_29705,N_24655,N_25065);
or U29706 (N_29706,N_24940,N_26670);
xor U29707 (N_29707,N_24447,N_26447);
or U29708 (N_29708,N_26676,N_26840);
or U29709 (N_29709,N_26120,N_24737);
or U29710 (N_29710,N_26807,N_26414);
or U29711 (N_29711,N_24001,N_24668);
and U29712 (N_29712,N_25542,N_26057);
and U29713 (N_29713,N_25430,N_26248);
or U29714 (N_29714,N_24833,N_26151);
nor U29715 (N_29715,N_26888,N_25580);
and U29716 (N_29716,N_26012,N_24385);
and U29717 (N_29717,N_25958,N_26672);
nor U29718 (N_29718,N_26741,N_24810);
or U29719 (N_29719,N_26381,N_25590);
nor U29720 (N_29720,N_25065,N_26814);
xor U29721 (N_29721,N_25696,N_24186);
or U29722 (N_29722,N_26607,N_26622);
xnor U29723 (N_29723,N_24679,N_25918);
xnor U29724 (N_29724,N_24652,N_25437);
nor U29725 (N_29725,N_24209,N_25290);
and U29726 (N_29726,N_26666,N_25663);
xor U29727 (N_29727,N_24725,N_26471);
nor U29728 (N_29728,N_24519,N_26894);
nand U29729 (N_29729,N_26256,N_25411);
xor U29730 (N_29730,N_24450,N_25607);
xnor U29731 (N_29731,N_24910,N_25233);
nor U29732 (N_29732,N_26734,N_24270);
and U29733 (N_29733,N_24776,N_26380);
xor U29734 (N_29734,N_24617,N_25844);
and U29735 (N_29735,N_26561,N_24151);
and U29736 (N_29736,N_26429,N_24788);
xor U29737 (N_29737,N_26585,N_24589);
and U29738 (N_29738,N_26851,N_24767);
xor U29739 (N_29739,N_26897,N_26881);
xnor U29740 (N_29740,N_26813,N_26675);
xnor U29741 (N_29741,N_26375,N_26159);
nor U29742 (N_29742,N_25423,N_24383);
xor U29743 (N_29743,N_25474,N_24725);
or U29744 (N_29744,N_26493,N_25644);
nor U29745 (N_29745,N_24397,N_25607);
xor U29746 (N_29746,N_26198,N_26175);
xor U29747 (N_29747,N_24439,N_25831);
and U29748 (N_29748,N_25601,N_24530);
xnor U29749 (N_29749,N_26500,N_25080);
nor U29750 (N_29750,N_26475,N_24623);
xnor U29751 (N_29751,N_24282,N_24692);
and U29752 (N_29752,N_24999,N_24592);
nor U29753 (N_29753,N_24287,N_25575);
nand U29754 (N_29754,N_24932,N_25047);
xor U29755 (N_29755,N_26589,N_24290);
and U29756 (N_29756,N_26974,N_26419);
nor U29757 (N_29757,N_24336,N_26614);
xor U29758 (N_29758,N_25862,N_24046);
and U29759 (N_29759,N_26111,N_24095);
xnor U29760 (N_29760,N_24964,N_24652);
and U29761 (N_29761,N_26258,N_26221);
or U29762 (N_29762,N_24498,N_24819);
nor U29763 (N_29763,N_25270,N_25417);
xor U29764 (N_29764,N_25351,N_26901);
nand U29765 (N_29765,N_26728,N_26210);
and U29766 (N_29766,N_25759,N_26168);
and U29767 (N_29767,N_25485,N_26725);
xor U29768 (N_29768,N_25042,N_26514);
nor U29769 (N_29769,N_26166,N_24513);
nor U29770 (N_29770,N_24904,N_25981);
or U29771 (N_29771,N_24020,N_25659);
xnor U29772 (N_29772,N_24460,N_26620);
xor U29773 (N_29773,N_25921,N_26967);
or U29774 (N_29774,N_26847,N_24430);
nor U29775 (N_29775,N_26577,N_25570);
xor U29776 (N_29776,N_25743,N_25732);
nand U29777 (N_29777,N_26960,N_26244);
or U29778 (N_29778,N_25848,N_24878);
and U29779 (N_29779,N_24065,N_25804);
or U29780 (N_29780,N_25278,N_25150);
nand U29781 (N_29781,N_25633,N_26865);
nand U29782 (N_29782,N_24695,N_24001);
and U29783 (N_29783,N_25471,N_26623);
xor U29784 (N_29784,N_24838,N_26342);
nor U29785 (N_29785,N_25734,N_24859);
or U29786 (N_29786,N_26007,N_24487);
nand U29787 (N_29787,N_25009,N_26915);
or U29788 (N_29788,N_24515,N_24667);
nand U29789 (N_29789,N_26828,N_25164);
or U29790 (N_29790,N_25374,N_25574);
xor U29791 (N_29791,N_26105,N_25952);
nor U29792 (N_29792,N_25270,N_24517);
nor U29793 (N_29793,N_26974,N_25044);
nor U29794 (N_29794,N_25389,N_24626);
xnor U29795 (N_29795,N_25906,N_26756);
and U29796 (N_29796,N_25404,N_24233);
or U29797 (N_29797,N_26186,N_26675);
and U29798 (N_29798,N_24993,N_26196);
nor U29799 (N_29799,N_25366,N_25484);
nor U29800 (N_29800,N_24971,N_24640);
or U29801 (N_29801,N_25110,N_24054);
nor U29802 (N_29802,N_26109,N_26842);
nor U29803 (N_29803,N_25163,N_24817);
xor U29804 (N_29804,N_24303,N_25454);
or U29805 (N_29805,N_24016,N_26282);
and U29806 (N_29806,N_25838,N_26680);
nand U29807 (N_29807,N_25610,N_24076);
xor U29808 (N_29808,N_25114,N_24004);
or U29809 (N_29809,N_24907,N_24712);
xnor U29810 (N_29810,N_24612,N_25231);
nand U29811 (N_29811,N_25249,N_24116);
xor U29812 (N_29812,N_24254,N_24164);
nand U29813 (N_29813,N_24456,N_24799);
and U29814 (N_29814,N_24736,N_25897);
nor U29815 (N_29815,N_24248,N_25632);
and U29816 (N_29816,N_25447,N_25409);
nand U29817 (N_29817,N_24920,N_25326);
nand U29818 (N_29818,N_25310,N_26332);
and U29819 (N_29819,N_26450,N_25578);
nand U29820 (N_29820,N_26506,N_25260);
xor U29821 (N_29821,N_26106,N_25693);
and U29822 (N_29822,N_24822,N_24048);
and U29823 (N_29823,N_26162,N_24173);
and U29824 (N_29824,N_24002,N_25873);
and U29825 (N_29825,N_26044,N_24812);
nand U29826 (N_29826,N_25946,N_24626);
nand U29827 (N_29827,N_24555,N_26366);
nor U29828 (N_29828,N_25865,N_24669);
nand U29829 (N_29829,N_26540,N_26838);
xor U29830 (N_29830,N_25009,N_25301);
and U29831 (N_29831,N_25209,N_25161);
nand U29832 (N_29832,N_24866,N_25984);
nand U29833 (N_29833,N_26109,N_25493);
nor U29834 (N_29834,N_25844,N_26984);
nand U29835 (N_29835,N_24455,N_26718);
nand U29836 (N_29836,N_26685,N_24141);
xor U29837 (N_29837,N_24272,N_25031);
xor U29838 (N_29838,N_26403,N_25455);
or U29839 (N_29839,N_26166,N_26307);
and U29840 (N_29840,N_25266,N_24082);
xor U29841 (N_29841,N_24803,N_26346);
nand U29842 (N_29842,N_25214,N_24390);
nand U29843 (N_29843,N_25776,N_26060);
nand U29844 (N_29844,N_25740,N_24054);
xor U29845 (N_29845,N_24457,N_25746);
xnor U29846 (N_29846,N_25354,N_25411);
or U29847 (N_29847,N_26147,N_25289);
nor U29848 (N_29848,N_25856,N_24433);
or U29849 (N_29849,N_25854,N_26720);
and U29850 (N_29850,N_24996,N_24850);
nand U29851 (N_29851,N_26609,N_26334);
or U29852 (N_29852,N_24528,N_25502);
and U29853 (N_29853,N_25725,N_26974);
and U29854 (N_29854,N_24073,N_25832);
nand U29855 (N_29855,N_24682,N_24802);
xor U29856 (N_29856,N_24166,N_25522);
nor U29857 (N_29857,N_24130,N_25996);
or U29858 (N_29858,N_24974,N_25748);
or U29859 (N_29859,N_24057,N_25815);
nor U29860 (N_29860,N_26007,N_24090);
or U29861 (N_29861,N_26304,N_25633);
xnor U29862 (N_29862,N_26594,N_26903);
nand U29863 (N_29863,N_26693,N_25323);
or U29864 (N_29864,N_24023,N_24198);
or U29865 (N_29865,N_25168,N_24551);
nand U29866 (N_29866,N_24145,N_26134);
nand U29867 (N_29867,N_26394,N_24460);
xor U29868 (N_29868,N_24771,N_26580);
or U29869 (N_29869,N_24768,N_26059);
xnor U29870 (N_29870,N_25697,N_25781);
xnor U29871 (N_29871,N_26107,N_26294);
nor U29872 (N_29872,N_25483,N_25501);
nand U29873 (N_29873,N_25741,N_24190);
nor U29874 (N_29874,N_26410,N_26934);
or U29875 (N_29875,N_25599,N_26097);
nor U29876 (N_29876,N_26894,N_26044);
and U29877 (N_29877,N_24321,N_26864);
nor U29878 (N_29878,N_25266,N_24838);
and U29879 (N_29879,N_24339,N_24127);
xor U29880 (N_29880,N_24027,N_26197);
nor U29881 (N_29881,N_25141,N_25434);
or U29882 (N_29882,N_25124,N_24318);
nor U29883 (N_29883,N_24486,N_24573);
nor U29884 (N_29884,N_24227,N_25519);
or U29885 (N_29885,N_25943,N_25896);
xnor U29886 (N_29886,N_24669,N_25732);
nand U29887 (N_29887,N_25181,N_25563);
nor U29888 (N_29888,N_25474,N_25653);
and U29889 (N_29889,N_26641,N_25579);
nand U29890 (N_29890,N_26026,N_24917);
xnor U29891 (N_29891,N_25392,N_26248);
and U29892 (N_29892,N_24913,N_24420);
nor U29893 (N_29893,N_25329,N_24232);
xor U29894 (N_29894,N_25931,N_26165);
nor U29895 (N_29895,N_25614,N_24174);
nand U29896 (N_29896,N_24107,N_26718);
nand U29897 (N_29897,N_26171,N_25256);
nor U29898 (N_29898,N_26744,N_24612);
and U29899 (N_29899,N_26267,N_24169);
and U29900 (N_29900,N_26103,N_24729);
nor U29901 (N_29901,N_24330,N_25676);
nand U29902 (N_29902,N_25063,N_24680);
and U29903 (N_29903,N_26295,N_24853);
nand U29904 (N_29904,N_25165,N_26928);
xor U29905 (N_29905,N_25470,N_24596);
nor U29906 (N_29906,N_24959,N_25231);
nor U29907 (N_29907,N_24099,N_26006);
or U29908 (N_29908,N_25625,N_26077);
nor U29909 (N_29909,N_25856,N_25500);
nand U29910 (N_29910,N_24165,N_25864);
nand U29911 (N_29911,N_24458,N_24120);
xnor U29912 (N_29912,N_26686,N_24150);
and U29913 (N_29913,N_25143,N_26881);
nand U29914 (N_29914,N_25934,N_25561);
and U29915 (N_29915,N_25716,N_24174);
xor U29916 (N_29916,N_25654,N_25988);
xnor U29917 (N_29917,N_24550,N_24048);
or U29918 (N_29918,N_26262,N_25808);
and U29919 (N_29919,N_24911,N_25586);
xor U29920 (N_29920,N_26013,N_25740);
xnor U29921 (N_29921,N_24459,N_24817);
and U29922 (N_29922,N_24828,N_24507);
and U29923 (N_29923,N_24812,N_26334);
or U29924 (N_29924,N_24270,N_26342);
or U29925 (N_29925,N_24937,N_26250);
nand U29926 (N_29926,N_24027,N_25817);
xnor U29927 (N_29927,N_24797,N_25349);
nand U29928 (N_29928,N_25974,N_24179);
and U29929 (N_29929,N_25496,N_24464);
and U29930 (N_29930,N_25759,N_26179);
nor U29931 (N_29931,N_24761,N_24106);
or U29932 (N_29932,N_24093,N_26747);
and U29933 (N_29933,N_25138,N_26487);
xor U29934 (N_29934,N_24792,N_26055);
or U29935 (N_29935,N_25740,N_26714);
nor U29936 (N_29936,N_24571,N_26838);
nor U29937 (N_29937,N_24948,N_26586);
xor U29938 (N_29938,N_26524,N_26017);
xor U29939 (N_29939,N_25965,N_26521);
xnor U29940 (N_29940,N_26568,N_25494);
or U29941 (N_29941,N_24107,N_24055);
nand U29942 (N_29942,N_24035,N_26796);
nand U29943 (N_29943,N_24160,N_25517);
nor U29944 (N_29944,N_24369,N_26911);
and U29945 (N_29945,N_26026,N_24942);
nor U29946 (N_29946,N_25512,N_26906);
xnor U29947 (N_29947,N_24448,N_25449);
nor U29948 (N_29948,N_26064,N_25382);
nor U29949 (N_29949,N_24375,N_24278);
or U29950 (N_29950,N_26973,N_25051);
xnor U29951 (N_29951,N_26462,N_26207);
xnor U29952 (N_29952,N_24246,N_25324);
or U29953 (N_29953,N_25789,N_26045);
and U29954 (N_29954,N_26622,N_25027);
and U29955 (N_29955,N_26267,N_26625);
xnor U29956 (N_29956,N_25637,N_26567);
and U29957 (N_29957,N_25622,N_26297);
xor U29958 (N_29958,N_26211,N_25586);
nand U29959 (N_29959,N_24764,N_25944);
nand U29960 (N_29960,N_25769,N_24024);
xor U29961 (N_29961,N_24296,N_25325);
xor U29962 (N_29962,N_25921,N_25517);
nor U29963 (N_29963,N_24754,N_26292);
nor U29964 (N_29964,N_25642,N_25236);
nor U29965 (N_29965,N_24452,N_26965);
nand U29966 (N_29966,N_24993,N_26652);
xnor U29967 (N_29967,N_25938,N_25779);
xor U29968 (N_29968,N_25440,N_26604);
nor U29969 (N_29969,N_26079,N_24086);
and U29970 (N_29970,N_25900,N_25562);
nand U29971 (N_29971,N_24412,N_26593);
nand U29972 (N_29972,N_25943,N_25325);
xor U29973 (N_29973,N_24087,N_26845);
and U29974 (N_29974,N_25839,N_26705);
nor U29975 (N_29975,N_25276,N_24224);
and U29976 (N_29976,N_25275,N_25152);
and U29977 (N_29977,N_25448,N_26740);
nor U29978 (N_29978,N_25015,N_26299);
nor U29979 (N_29979,N_26724,N_25692);
nand U29980 (N_29980,N_25263,N_24519);
nor U29981 (N_29981,N_24021,N_25888);
and U29982 (N_29982,N_25577,N_24674);
or U29983 (N_29983,N_26051,N_25618);
and U29984 (N_29984,N_24488,N_26546);
nor U29985 (N_29985,N_25058,N_26445);
or U29986 (N_29986,N_26687,N_26011);
xor U29987 (N_29987,N_24058,N_26943);
nor U29988 (N_29988,N_25141,N_26167);
nand U29989 (N_29989,N_25044,N_26047);
or U29990 (N_29990,N_25364,N_26276);
xor U29991 (N_29991,N_25555,N_26200);
nand U29992 (N_29992,N_25113,N_25506);
nand U29993 (N_29993,N_24725,N_26237);
nor U29994 (N_29994,N_24125,N_26842);
xnor U29995 (N_29995,N_25028,N_26259);
nand U29996 (N_29996,N_24727,N_26774);
or U29997 (N_29997,N_26136,N_25208);
nand U29998 (N_29998,N_26859,N_24554);
and U29999 (N_29999,N_24465,N_26588);
nor UO_0 (O_0,N_28367,N_28938);
nor UO_1 (O_1,N_27273,N_27798);
xor UO_2 (O_2,N_27698,N_27958);
nand UO_3 (O_3,N_29161,N_27948);
nand UO_4 (O_4,N_28679,N_28566);
xor UO_5 (O_5,N_29006,N_29024);
nand UO_6 (O_6,N_29295,N_29102);
nand UO_7 (O_7,N_29289,N_27704);
xor UO_8 (O_8,N_28258,N_27239);
nand UO_9 (O_9,N_27506,N_29101);
and UO_10 (O_10,N_29713,N_27579);
nand UO_11 (O_11,N_29346,N_27565);
or UO_12 (O_12,N_29103,N_28098);
and UO_13 (O_13,N_28345,N_28958);
and UO_14 (O_14,N_27288,N_27102);
nor UO_15 (O_15,N_28822,N_28494);
nor UO_16 (O_16,N_27540,N_27258);
and UO_17 (O_17,N_29555,N_28721);
nor UO_18 (O_18,N_27525,N_29091);
nor UO_19 (O_19,N_27402,N_29473);
or UO_20 (O_20,N_28633,N_27117);
and UO_21 (O_21,N_29232,N_27635);
nor UO_22 (O_22,N_29076,N_28615);
xnor UO_23 (O_23,N_28217,N_28265);
nand UO_24 (O_24,N_28834,N_29418);
nand UO_25 (O_25,N_27602,N_29347);
xnor UO_26 (O_26,N_27189,N_29335);
xnor UO_27 (O_27,N_29435,N_28038);
nor UO_28 (O_28,N_28002,N_28324);
nand UO_29 (O_29,N_29797,N_27765);
nor UO_30 (O_30,N_28982,N_28313);
nand UO_31 (O_31,N_29953,N_29805);
or UO_32 (O_32,N_29446,N_27379);
nor UO_33 (O_33,N_28851,N_27970);
xnor UO_34 (O_34,N_27995,N_28144);
or UO_35 (O_35,N_29707,N_28832);
and UO_36 (O_36,N_27904,N_27663);
and UO_37 (O_37,N_29959,N_28348);
and UO_38 (O_38,N_28584,N_28638);
and UO_39 (O_39,N_27289,N_28937);
nor UO_40 (O_40,N_28435,N_27697);
or UO_41 (O_41,N_29643,N_28473);
nor UO_42 (O_42,N_27768,N_28527);
and UO_43 (O_43,N_27243,N_27639);
or UO_44 (O_44,N_28541,N_28409);
xor UO_45 (O_45,N_28316,N_28155);
xnor UO_46 (O_46,N_28802,N_29297);
nor UO_47 (O_47,N_28942,N_28526);
nor UO_48 (O_48,N_27286,N_27888);
xnor UO_49 (O_49,N_28768,N_27574);
nor UO_50 (O_50,N_28852,N_27595);
or UO_51 (O_51,N_29382,N_28547);
and UO_52 (O_52,N_27305,N_27363);
and UO_53 (O_53,N_28051,N_28126);
and UO_54 (O_54,N_27311,N_28075);
nand UO_55 (O_55,N_27984,N_27673);
xnor UO_56 (O_56,N_28684,N_29256);
and UO_57 (O_57,N_28119,N_28833);
xor UO_58 (O_58,N_27365,N_28025);
and UO_59 (O_59,N_28077,N_27324);
nand UO_60 (O_60,N_27309,N_27790);
nand UO_61 (O_61,N_28796,N_29300);
nand UO_62 (O_62,N_28891,N_28425);
and UO_63 (O_63,N_27781,N_29921);
or UO_64 (O_64,N_28629,N_28718);
nor UO_65 (O_65,N_29552,N_28790);
nand UO_66 (O_66,N_29238,N_28442);
or UO_67 (O_67,N_27800,N_29119);
and UO_68 (O_68,N_28818,N_29618);
or UO_69 (O_69,N_28397,N_28807);
nand UO_70 (O_70,N_27035,N_29367);
xnor UO_71 (O_71,N_27213,N_29170);
nor UO_72 (O_72,N_29833,N_28900);
nor UO_73 (O_73,N_27617,N_29026);
and UO_74 (O_74,N_29392,N_29225);
xor UO_75 (O_75,N_28582,N_29812);
xor UO_76 (O_76,N_27822,N_27632);
and UO_77 (O_77,N_28377,N_27393);
nand UO_78 (O_78,N_28734,N_27333);
nand UO_79 (O_79,N_28018,N_28107);
nor UO_80 (O_80,N_28996,N_28339);
and UO_81 (O_81,N_29796,N_27714);
or UO_82 (O_82,N_27631,N_27915);
and UO_83 (O_83,N_27348,N_27813);
and UO_84 (O_84,N_27121,N_27621);
nor UO_85 (O_85,N_29730,N_27657);
and UO_86 (O_86,N_28487,N_28167);
xnor UO_87 (O_87,N_27486,N_29989);
nand UO_88 (O_88,N_27655,N_27173);
or UO_89 (O_89,N_29031,N_28291);
or UO_90 (O_90,N_29700,N_28088);
nand UO_91 (O_91,N_28800,N_29742);
and UO_92 (O_92,N_27523,N_29889);
or UO_93 (O_93,N_27537,N_29692);
or UO_94 (O_94,N_28656,N_27116);
and UO_95 (O_95,N_27476,N_29041);
nand UO_96 (O_96,N_28248,N_29158);
or UO_97 (O_97,N_27505,N_27844);
xor UO_98 (O_98,N_29985,N_29913);
xnor UO_99 (O_99,N_28955,N_28207);
and UO_100 (O_100,N_27508,N_29563);
nand UO_101 (O_101,N_29818,N_27404);
nand UO_102 (O_102,N_28616,N_29981);
and UO_103 (O_103,N_27222,N_28137);
nor UO_104 (O_104,N_27108,N_28559);
nand UO_105 (O_105,N_28598,N_27923);
nand UO_106 (O_106,N_28784,N_28285);
or UO_107 (O_107,N_29512,N_29670);
and UO_108 (O_108,N_28024,N_28223);
and UO_109 (O_109,N_28558,N_29544);
xnor UO_110 (O_110,N_28497,N_29665);
or UO_111 (O_111,N_27088,N_27753);
and UO_112 (O_112,N_29301,N_28754);
nor UO_113 (O_113,N_29129,N_28522);
or UO_114 (O_114,N_29058,N_27566);
nor UO_115 (O_115,N_28694,N_28774);
xnor UO_116 (O_116,N_28564,N_28429);
and UO_117 (O_117,N_29570,N_28720);
nand UO_118 (O_118,N_29716,N_27864);
xor UO_119 (O_119,N_28404,N_28132);
nor UO_120 (O_120,N_27067,N_29595);
xnor UO_121 (O_121,N_27019,N_29711);
and UO_122 (O_122,N_29004,N_27648);
xor UO_123 (O_123,N_28163,N_29896);
nand UO_124 (O_124,N_29747,N_27316);
nor UO_125 (O_125,N_29467,N_29630);
nand UO_126 (O_126,N_28118,N_29503);
xor UO_127 (O_127,N_27827,N_28978);
nor UO_128 (O_128,N_29649,N_28658);
nand UO_129 (O_129,N_28214,N_28446);
nand UO_130 (O_130,N_27453,N_28444);
xnor UO_131 (O_131,N_28931,N_29083);
xnor UO_132 (O_132,N_27164,N_27887);
and UO_133 (O_133,N_29694,N_28538);
nor UO_134 (O_134,N_29380,N_27496);
nor UO_135 (O_135,N_27025,N_27469);
nand UO_136 (O_136,N_27747,N_29815);
nor UO_137 (O_137,N_29152,N_29086);
or UO_138 (O_138,N_28260,N_29881);
nand UO_139 (O_139,N_28640,N_27352);
nor UO_140 (O_140,N_27122,N_28460);
xnor UO_141 (O_141,N_28114,N_29729);
nand UO_142 (O_142,N_29837,N_28927);
or UO_143 (O_143,N_29991,N_28950);
or UO_144 (O_144,N_29764,N_27694);
xnor UO_145 (O_145,N_28687,N_29343);
xnor UO_146 (O_146,N_28773,N_29982);
xnor UO_147 (O_147,N_27332,N_29847);
nor UO_148 (O_148,N_29314,N_28850);
xnor UO_149 (O_149,N_27702,N_28352);
xor UO_150 (O_150,N_29299,N_28874);
or UO_151 (O_151,N_27172,N_28231);
and UO_152 (O_152,N_28635,N_29931);
or UO_153 (O_153,N_28110,N_28310);
nor UO_154 (O_154,N_28935,N_29506);
or UO_155 (O_155,N_29371,N_28235);
nor UO_156 (O_156,N_28856,N_29614);
and UO_157 (O_157,N_28337,N_27950);
and UO_158 (O_158,N_28142,N_27170);
or UO_159 (O_159,N_27290,N_27128);
nor UO_160 (O_160,N_27489,N_27852);
or UO_161 (O_161,N_29691,N_29903);
xor UO_162 (O_162,N_27903,N_29140);
nand UO_163 (O_163,N_27291,N_28432);
and UO_164 (O_164,N_27658,N_28454);
nand UO_165 (O_165,N_29949,N_29112);
nor UO_166 (O_166,N_27608,N_29012);
xnor UO_167 (O_167,N_28863,N_29302);
nor UO_168 (O_168,N_28783,N_27878);
nor UO_169 (O_169,N_29217,N_28924);
nand UO_170 (O_170,N_27115,N_28692);
xor UO_171 (O_171,N_27487,N_27778);
or UO_172 (O_172,N_28458,N_29693);
and UO_173 (O_173,N_27840,N_28325);
nand UO_174 (O_174,N_29702,N_29378);
nand UO_175 (O_175,N_28908,N_29211);
xor UO_176 (O_176,N_27004,N_27780);
or UO_177 (O_177,N_27089,N_29278);
xnor UO_178 (O_178,N_29125,N_28866);
and UO_179 (O_179,N_27362,N_27132);
and UO_180 (O_180,N_29735,N_28683);
nand UO_181 (O_181,N_29843,N_27622);
or UO_182 (O_182,N_27819,N_27816);
and UO_183 (O_183,N_29884,N_28353);
nor UO_184 (O_184,N_27939,N_29840);
nor UO_185 (O_185,N_29460,N_27337);
and UO_186 (O_186,N_27999,N_29718);
or UO_187 (O_187,N_27640,N_29000);
or UO_188 (O_188,N_28105,N_28135);
xnor UO_189 (O_189,N_27796,N_29775);
and UO_190 (O_190,N_27630,N_28251);
and UO_191 (O_191,N_27361,N_28765);
nor UO_192 (O_192,N_28063,N_27231);
or UO_193 (O_193,N_28647,N_29962);
xnor UO_194 (O_194,N_28910,N_27298);
and UO_195 (O_195,N_27136,N_29410);
nand UO_196 (O_196,N_28632,N_27513);
and UO_197 (O_197,N_29858,N_27909);
and UO_198 (O_198,N_29280,N_27502);
nand UO_199 (O_199,N_28222,N_27691);
nor UO_200 (O_200,N_28708,N_29009);
or UO_201 (O_201,N_27788,N_28090);
xor UO_202 (O_202,N_28686,N_29329);
and UO_203 (O_203,N_28552,N_29627);
xor UO_204 (O_204,N_27148,N_29532);
and UO_205 (O_205,N_29893,N_29844);
nor UO_206 (O_206,N_29207,N_29496);
nand UO_207 (O_207,N_28837,N_28287);
xnor UO_208 (O_208,N_28424,N_29476);
or UO_209 (O_209,N_27899,N_27905);
nand UO_210 (O_210,N_27944,N_27922);
xnor UO_211 (O_211,N_27779,N_28603);
xnor UO_212 (O_212,N_29871,N_29151);
nor UO_213 (O_213,N_27500,N_29356);
or UO_214 (O_214,N_27591,N_29230);
xor UO_215 (O_215,N_29639,N_27634);
and UO_216 (O_216,N_28083,N_29533);
and UO_217 (O_217,N_29891,N_28117);
nor UO_218 (O_218,N_28346,N_27151);
nand UO_219 (O_219,N_29857,N_27212);
nand UO_220 (O_220,N_27933,N_29104);
or UO_221 (O_221,N_28069,N_28769);
nand UO_222 (O_222,N_28940,N_28200);
or UO_223 (O_223,N_27044,N_28408);
and UO_224 (O_224,N_28032,N_29423);
nand UO_225 (O_225,N_27257,N_28378);
and UO_226 (O_226,N_27917,N_29972);
or UO_227 (O_227,N_28590,N_29591);
nand UO_228 (O_228,N_29187,N_29518);
and UO_229 (O_229,N_28358,N_28080);
xnor UO_230 (O_230,N_27921,N_28967);
xnor UO_231 (O_231,N_27628,N_27340);
or UO_232 (O_232,N_27875,N_27495);
or UO_233 (O_233,N_27641,N_28376);
nor UO_234 (O_234,N_27432,N_27472);
or UO_235 (O_235,N_27374,N_28570);
nor UO_236 (O_236,N_27664,N_29429);
nor UO_237 (O_237,N_29536,N_28812);
xor UO_238 (O_238,N_29935,N_27059);
xnor UO_239 (O_239,N_27836,N_28809);
nand UO_240 (O_240,N_29092,N_29479);
nor UO_241 (O_241,N_29059,N_28440);
and UO_242 (O_242,N_29576,N_29906);
xnor UO_243 (O_243,N_28512,N_28776);
or UO_244 (O_244,N_28921,N_27569);
nand UO_245 (O_245,N_27614,N_27428);
or UO_246 (O_246,N_29724,N_29345);
or UO_247 (O_247,N_27620,N_27831);
and UO_248 (O_248,N_27400,N_28961);
nor UO_249 (O_249,N_27419,N_27031);
xor UO_250 (O_250,N_28322,N_28459);
nor UO_251 (O_251,N_29541,N_29197);
and UO_252 (O_252,N_28033,N_28308);
and UO_253 (O_253,N_28825,N_28010);
nor UO_254 (O_254,N_29354,N_27283);
nand UO_255 (O_255,N_27558,N_28923);
or UO_256 (O_256,N_28021,N_28595);
and UO_257 (O_257,N_27734,N_29636);
nand UO_258 (O_258,N_29279,N_27588);
and UO_259 (O_259,N_28944,N_27416);
or UO_260 (O_260,N_29594,N_29176);
nand UO_261 (O_261,N_29562,N_29244);
and UO_262 (O_262,N_27138,N_27751);
and UO_263 (O_263,N_28336,N_29760);
and UO_264 (O_264,N_27656,N_28620);
and UO_265 (O_265,N_28323,N_29668);
xnor UO_266 (O_266,N_27280,N_27727);
nor UO_267 (O_267,N_28735,N_28003);
and UO_268 (O_268,N_29717,N_28816);
or UO_269 (O_269,N_29141,N_29990);
xor UO_270 (O_270,N_27011,N_29886);
nor UO_271 (O_271,N_28930,N_28299);
xor UO_272 (O_272,N_29172,N_29638);
and UO_273 (O_273,N_27721,N_28511);
nand UO_274 (O_274,N_27880,N_29768);
nand UO_275 (O_275,N_29338,N_28168);
nor UO_276 (O_276,N_28127,N_27360);
and UO_277 (O_277,N_29852,N_27801);
and UO_278 (O_278,N_29676,N_28536);
nor UO_279 (O_279,N_29430,N_29621);
and UO_280 (O_280,N_28344,N_27203);
nand UO_281 (O_281,N_28549,N_28861);
xnor UO_282 (O_282,N_29043,N_28298);
and UO_283 (O_283,N_28661,N_27335);
nand UO_284 (O_284,N_29229,N_29419);
nor UO_285 (O_285,N_27692,N_29409);
nor UO_286 (O_286,N_27985,N_28139);
xor UO_287 (O_287,N_27443,N_27205);
nor UO_288 (O_288,N_27870,N_28030);
nand UO_289 (O_289,N_28140,N_27809);
xor UO_290 (O_290,N_28518,N_27499);
nand UO_291 (O_291,N_27810,N_29249);
and UO_292 (O_292,N_28876,N_27271);
or UO_293 (O_293,N_29659,N_29177);
nand UO_294 (O_294,N_29205,N_29667);
and UO_295 (O_295,N_28501,N_27907);
xnor UO_296 (O_296,N_27889,N_28742);
and UO_297 (O_297,N_28901,N_28680);
xnor UO_298 (O_298,N_27494,N_29267);
nor UO_299 (O_299,N_28622,N_27372);
nor UO_300 (O_300,N_29396,N_28277);
or UO_301 (O_301,N_28681,N_29275);
xor UO_302 (O_302,N_27078,N_29027);
or UO_303 (O_303,N_27871,N_27051);
and UO_304 (O_304,N_29139,N_27339);
or UO_305 (O_305,N_27133,N_28793);
nand UO_306 (O_306,N_28304,N_27988);
xor UO_307 (O_307,N_29660,N_28480);
nor UO_308 (O_308,N_28648,N_28410);
nand UO_309 (O_309,N_27869,N_27086);
nor UO_310 (O_310,N_28250,N_29808);
nor UO_311 (O_311,N_27771,N_29568);
nand UO_312 (O_312,N_28301,N_27552);
xnor UO_313 (O_313,N_29957,N_29344);
nor UO_314 (O_314,N_29883,N_28414);
nor UO_315 (O_315,N_27976,N_28556);
and UO_316 (O_316,N_29922,N_27392);
or UO_317 (O_317,N_28284,N_27282);
and UO_318 (O_318,N_27610,N_28569);
xor UO_319 (O_319,N_28949,N_28659);
nor UO_320 (O_320,N_29795,N_29710);
xor UO_321 (O_321,N_28922,N_28292);
and UO_322 (O_322,N_29622,N_27979);
nor UO_323 (O_323,N_29401,N_27549);
nor UO_324 (O_324,N_29235,N_27010);
xor UO_325 (O_325,N_28332,N_28843);
xnor UO_326 (O_326,N_29865,N_27746);
and UO_327 (O_327,N_27015,N_27936);
or UO_328 (O_328,N_28011,N_27793);
or UO_329 (O_329,N_28384,N_29697);
nand UO_330 (O_330,N_29358,N_27550);
and UO_331 (O_331,N_27227,N_27341);
and UO_332 (O_332,N_29493,N_29264);
nand UO_333 (O_333,N_27693,N_28502);
and UO_334 (O_334,N_28929,N_29892);
nor UO_335 (O_335,N_28819,N_29640);
xor UO_336 (O_336,N_28070,N_27597);
or UO_337 (O_337,N_28491,N_27450);
or UO_338 (O_338,N_29513,N_27862);
xnor UO_339 (O_339,N_27932,N_28300);
or UO_340 (O_340,N_29519,N_28252);
and UO_341 (O_341,N_29528,N_29557);
or UO_342 (O_342,N_29976,N_28205);
nand UO_343 (O_343,N_29882,N_28143);
nor UO_344 (O_344,N_27546,N_29073);
and UO_345 (O_345,N_27696,N_28586);
nand UO_346 (O_346,N_29696,N_27961);
nor UO_347 (O_347,N_28048,N_29067);
nor UO_348 (O_348,N_28677,N_27168);
nor UO_349 (O_349,N_27249,N_29209);
nand UO_350 (O_350,N_28159,N_27192);
or UO_351 (O_351,N_27448,N_27876);
nand UO_352 (O_352,N_27651,N_27049);
xor UO_353 (O_353,N_28594,N_27420);
nor UO_354 (O_354,N_27789,N_28879);
or UO_355 (O_355,N_27866,N_29975);
or UO_356 (O_356,N_28014,N_28903);
nor UO_357 (O_357,N_29566,N_29744);
and UO_358 (O_358,N_27633,N_28229);
nand UO_359 (O_359,N_29310,N_29547);
xnor UO_360 (O_360,N_28400,N_27848);
and UO_361 (O_361,N_27322,N_28412);
nor UO_362 (O_362,N_27050,N_27206);
nand UO_363 (O_363,N_29543,N_29628);
or UO_364 (O_364,N_29619,N_29577);
nor UO_365 (O_365,N_28870,N_27808);
or UO_366 (O_366,N_29321,N_28206);
and UO_367 (O_367,N_27397,N_29234);
nor UO_368 (O_368,N_28892,N_28398);
nand UO_369 (O_369,N_27578,N_29992);
nand UO_370 (O_370,N_27966,N_27667);
nand UO_371 (O_371,N_29658,N_29414);
nand UO_372 (O_372,N_28433,N_27385);
nand UO_373 (O_373,N_28360,N_27514);
xnor UO_374 (O_374,N_29996,N_27737);
or UO_375 (O_375,N_29811,N_28618);
nor UO_376 (O_376,N_28704,N_29826);
and UO_377 (O_377,N_28395,N_28309);
nor UO_378 (O_378,N_27216,N_29383);
or UO_379 (O_379,N_29997,N_29567);
or UO_380 (O_380,N_29644,N_27171);
and UO_381 (O_381,N_27021,N_29880);
or UO_382 (O_382,N_29223,N_28289);
and UO_383 (O_383,N_29099,N_28666);
nand UO_384 (O_384,N_27854,N_27992);
nand UO_385 (O_385,N_29115,N_28977);
and UO_386 (O_386,N_27201,N_27371);
xor UO_387 (O_387,N_27561,N_29281);
nand UO_388 (O_388,N_29486,N_28668);
xnor UO_389 (O_389,N_28976,N_29799);
xnor UO_390 (O_390,N_29774,N_27806);
or UO_391 (O_391,N_29938,N_27193);
and UO_392 (O_392,N_29360,N_28789);
nand UO_393 (O_393,N_29825,N_27037);
nor UO_394 (O_394,N_29965,N_28148);
nor UO_395 (O_395,N_28467,N_29110);
or UO_396 (O_396,N_29539,N_29182);
nor UO_397 (O_397,N_29846,N_28665);
or UO_398 (O_398,N_29542,N_27557);
or UO_399 (O_399,N_28185,N_27660);
xor UO_400 (O_400,N_27699,N_29391);
xnor UO_401 (O_401,N_28951,N_27710);
or UO_402 (O_402,N_29304,N_27612);
nor UO_403 (O_403,N_28510,N_28952);
xor UO_404 (O_404,N_29860,N_29137);
nand UO_405 (O_405,N_29100,N_29390);
nand UO_406 (O_406,N_28259,N_29185);
or UO_407 (O_407,N_27518,N_29426);
xor UO_408 (O_408,N_28046,N_27884);
nand UO_409 (O_409,N_29489,N_27481);
and UO_410 (O_410,N_28780,N_28350);
nand UO_411 (O_411,N_27782,N_27729);
or UO_412 (O_412,N_28226,N_29450);
and UO_413 (O_413,N_28797,N_27849);
or UO_414 (O_414,N_29274,N_29483);
and UO_415 (O_415,N_29436,N_27485);
nand UO_416 (O_416,N_29245,N_28994);
nand UO_417 (O_417,N_28027,N_28389);
and UO_418 (O_418,N_29520,N_29924);
or UO_419 (O_419,N_28374,N_29854);
or UO_420 (O_420,N_27176,N_27344);
nand UO_421 (O_421,N_29218,N_28072);
xor UO_422 (O_422,N_28544,N_27731);
nor UO_423 (O_423,N_27356,N_29984);
or UO_424 (O_424,N_27376,N_27214);
nand UO_425 (O_425,N_27947,N_27066);
xor UO_426 (O_426,N_28411,N_28194);
and UO_427 (O_427,N_29895,N_27263);
or UO_428 (O_428,N_28263,N_28236);
or UO_429 (O_429,N_27145,N_27538);
and UO_430 (O_430,N_28238,N_27388);
nor UO_431 (O_431,N_27471,N_28490);
nor UO_432 (O_432,N_29866,N_29986);
and UO_433 (O_433,N_27742,N_28181);
or UO_434 (O_434,N_27726,N_27383);
xor UO_435 (O_435,N_28877,N_28736);
nand UO_436 (O_436,N_28560,N_27616);
and UO_437 (O_437,N_27841,N_27490);
and UO_438 (O_438,N_28887,N_29449);
xor UO_439 (O_439,N_29637,N_29745);
and UO_440 (O_440,N_27129,N_28878);
and UO_441 (O_441,N_28956,N_27056);
or UO_442 (O_442,N_27296,N_27937);
xnor UO_443 (O_443,N_28208,N_29406);
nand UO_444 (O_444,N_28652,N_27034);
or UO_445 (O_445,N_28792,N_28203);
nand UO_446 (O_446,N_29323,N_29664);
xor UO_447 (O_447,N_29404,N_28094);
nor UO_448 (O_448,N_27587,N_27814);
or UO_449 (O_449,N_27366,N_27260);
or UO_450 (O_450,N_28995,N_29875);
or UO_451 (O_451,N_27526,N_29969);
or UO_452 (O_452,N_29477,N_29191);
nor UO_453 (O_453,N_27713,N_29173);
or UO_454 (O_454,N_29020,N_28757);
nor UO_455 (O_455,N_28953,N_29085);
nand UO_456 (O_456,N_27241,N_29242);
nor UO_457 (O_457,N_27047,N_29060);
nor UO_458 (O_458,N_27079,N_29333);
or UO_459 (O_459,N_28192,N_28363);
nor UO_460 (O_460,N_27276,N_27097);
nor UO_461 (O_461,N_28423,N_28481);
xnor UO_462 (O_462,N_27528,N_28897);
and UO_463 (O_463,N_28709,N_29038);
and UO_464 (O_464,N_27347,N_29879);
nor UO_465 (O_465,N_28814,N_28649);
nor UO_466 (O_466,N_29427,N_29733);
and UO_467 (O_467,N_28746,N_29171);
or UO_468 (O_468,N_29017,N_28577);
nand UO_469 (O_469,N_28416,N_28602);
nand UO_470 (O_470,N_28065,N_27901);
or UO_471 (O_471,N_27874,N_29788);
nand UO_472 (O_472,N_28147,N_27955);
xor UO_473 (O_473,N_28124,N_28240);
nor UO_474 (O_474,N_27568,N_28478);
and UO_475 (O_475,N_27188,N_27245);
and UO_476 (O_476,N_27020,N_28914);
and UO_477 (O_477,N_29432,N_29079);
xor UO_478 (O_478,N_28019,N_27748);
nand UO_479 (O_479,N_29910,N_27509);
or UO_480 (O_480,N_27084,N_29090);
or UO_481 (O_481,N_27477,N_28732);
xor UO_482 (O_482,N_28617,N_27386);
or UO_483 (O_483,N_27261,N_29442);
and UO_484 (O_484,N_28778,N_28281);
or UO_485 (O_485,N_29045,N_27223);
or UO_486 (O_486,N_28744,N_27912);
xor UO_487 (O_487,N_27629,N_28172);
and UO_488 (O_488,N_27517,N_29780);
xor UO_489 (O_489,N_29929,N_29573);
and UO_490 (O_490,N_27334,N_28001);
nor UO_491 (O_491,N_29272,N_28096);
and UO_492 (O_492,N_29210,N_28642);
and UO_493 (O_493,N_27843,N_29312);
or UO_494 (O_494,N_28349,N_28904);
or UO_495 (O_495,N_27716,N_28873);
nor UO_496 (O_496,N_28115,N_29683);
or UO_497 (O_497,N_28268,N_29262);
nand UO_498 (O_498,N_27914,N_28915);
or UO_499 (O_499,N_29934,N_29352);
xnor UO_500 (O_500,N_27475,N_28161);
xor UO_501 (O_501,N_28368,N_29325);
and UO_502 (O_502,N_28209,N_29296);
and UO_503 (O_503,N_28434,N_28074);
nand UO_504 (O_504,N_29007,N_27934);
or UO_505 (O_505,N_27717,N_28762);
nand UO_506 (O_506,N_28087,N_29021);
xnor UO_507 (O_507,N_29388,N_28043);
xor UO_508 (O_508,N_29184,N_29736);
and UO_509 (O_509,N_29954,N_28554);
nor UO_510 (O_510,N_27968,N_28557);
xor UO_511 (O_511,N_28402,N_28724);
or UO_512 (O_512,N_28306,N_29677);
nor UO_513 (O_513,N_28770,N_28420);
nor UO_514 (O_514,N_27458,N_28026);
and UO_515 (O_515,N_27233,N_28959);
and UO_516 (O_516,N_27929,N_27650);
xor UO_517 (O_517,N_29482,N_27928);
or UO_518 (O_518,N_29615,N_28563);
nor UO_519 (O_519,N_27761,N_27626);
xor UO_520 (O_520,N_27155,N_27109);
or UO_521 (O_521,N_27962,N_27179);
nand UO_522 (O_522,N_28795,N_29196);
xor UO_523 (O_523,N_27785,N_27389);
nor UO_524 (O_524,N_29819,N_28320);
nor UO_525 (O_525,N_29689,N_27358);
nor UO_526 (O_526,N_28371,N_28509);
xor UO_527 (O_527,N_27680,N_29646);
nor UO_528 (O_528,N_27426,N_29631);
nor UO_529 (O_529,N_27902,N_29937);
or UO_530 (O_530,N_29387,N_27449);
or UO_531 (O_531,N_29926,N_27842);
and UO_532 (O_532,N_28838,N_28946);
xor UO_533 (O_533,N_27330,N_27314);
and UO_534 (O_534,N_29444,N_29878);
nor UO_535 (O_535,N_27211,N_28614);
nor UO_536 (O_536,N_28387,N_28484);
nor UO_537 (O_537,N_27113,N_29868);
nor UO_538 (O_538,N_27867,N_28849);
and UO_539 (O_539,N_28351,N_27225);
or UO_540 (O_540,N_28129,N_27963);
and UO_541 (O_541,N_28261,N_29600);
nand UO_542 (O_542,N_28710,N_28969);
nand UO_543 (O_543,N_29257,N_27492);
nand UO_544 (O_544,N_27462,N_28215);
or UO_545 (O_545,N_27182,N_27857);
nand UO_546 (O_546,N_29164,N_29771);
or UO_547 (O_547,N_27281,N_28815);
or UO_548 (O_548,N_29616,N_29909);
xor UO_549 (O_549,N_27355,N_29373);
nand UO_550 (O_550,N_29331,N_29226);
or UO_551 (O_551,N_28199,N_27774);
nor UO_552 (O_552,N_27491,N_27548);
and UO_553 (O_553,N_28439,N_27807);
xor UO_554 (O_554,N_29407,N_27977);
nand UO_555 (O_555,N_27199,N_28755);
and UO_556 (O_556,N_29824,N_28326);
or UO_557 (O_557,N_28198,N_29502);
nand UO_558 (O_558,N_28134,N_27743);
xor UO_559 (O_559,N_27722,N_27007);
xnor UO_560 (O_560,N_29499,N_29798);
or UO_561 (O_561,N_27275,N_29899);
nor UO_562 (O_562,N_28727,N_27756);
xor UO_563 (O_563,N_27749,N_29597);
and UO_564 (O_564,N_29923,N_27161);
xor UO_565 (O_565,N_29578,N_29468);
and UO_566 (O_566,N_29379,N_28330);
xor UO_567 (O_567,N_29132,N_28657);
xor UO_568 (O_568,N_29240,N_28885);
or UO_569 (O_569,N_28574,N_28171);
and UO_570 (O_570,N_29741,N_28548);
or UO_571 (O_571,N_29298,N_28821);
and UO_572 (O_572,N_28103,N_29967);
xor UO_573 (O_573,N_28047,N_27606);
nor UO_574 (O_574,N_29361,N_28157);
xor UO_575 (O_575,N_29606,N_28216);
xnor UO_576 (O_576,N_27094,N_27042);
and UO_577 (O_577,N_27707,N_27405);
or UO_578 (O_578,N_28919,N_29385);
or UO_579 (O_579,N_29516,N_28997);
nor UO_580 (O_580,N_28610,N_29292);
xnor UO_581 (O_581,N_29887,N_27653);
nand UO_582 (O_582,N_29447,N_27695);
xor UO_583 (O_583,N_29332,N_27980);
and UO_584 (O_584,N_29495,N_28884);
xor UO_585 (O_585,N_29114,N_28627);
xnor UO_586 (O_586,N_27351,N_27002);
and UO_587 (O_587,N_28280,N_29575);
nor UO_588 (O_588,N_27882,N_28315);
xor UO_589 (O_589,N_28868,N_27270);
xor UO_590 (O_590,N_29154,N_27230);
xor UO_591 (O_591,N_27357,N_28820);
or UO_592 (O_592,N_29106,N_28283);
or UO_593 (O_593,N_29146,N_29925);
xor UO_594 (O_594,N_29554,N_28111);
and UO_595 (O_595,N_27126,N_28369);
nor UO_596 (O_596,N_28609,N_29813);
or UO_597 (O_597,N_28045,N_29941);
or UO_598 (O_598,N_27068,N_27478);
or UO_599 (O_599,N_27169,N_27762);
nor UO_600 (O_600,N_29453,N_28968);
nor UO_601 (O_601,N_28865,N_27954);
and UO_602 (O_602,N_28012,N_28894);
nor UO_603 (O_603,N_29734,N_29605);
nand UO_604 (O_604,N_29096,N_27745);
nand UO_605 (O_605,N_29698,N_27278);
xor UO_606 (O_606,N_28380,N_27256);
xor UO_607 (O_607,N_28255,N_29351);
nor UO_608 (O_608,N_27433,N_29376);
and UO_609 (O_609,N_29920,N_28334);
xnor UO_610 (O_610,N_27081,N_27338);
nand UO_611 (O_611,N_29180,N_28007);
nor UO_612 (O_612,N_28791,N_28356);
and UO_613 (O_613,N_29582,N_27114);
or UO_614 (O_614,N_29136,N_28623);
nand UO_615 (O_615,N_27045,N_27493);
nand UO_616 (O_616,N_29770,N_27209);
and UO_617 (O_617,N_28751,N_28782);
or UO_618 (O_618,N_28370,N_27252);
nand UO_619 (O_619,N_29960,N_28102);
or UO_620 (O_620,N_27301,N_29781);
xor UO_621 (O_621,N_28406,N_27391);
and UO_622 (O_622,N_29704,N_27036);
nand UO_623 (O_623,N_27140,N_28730);
and UO_624 (O_624,N_28392,N_29551);
or UO_625 (O_625,N_27159,N_29324);
nand UO_626 (O_626,N_29349,N_27439);
or UO_627 (O_627,N_28278,N_29309);
xnor UO_628 (O_628,N_28965,N_28880);
or UO_629 (O_629,N_28886,N_29732);
or UO_630 (O_630,N_29652,N_29968);
nand UO_631 (O_631,N_29629,N_28095);
or UO_632 (O_632,N_29834,N_28813);
and UO_633 (O_633,N_27971,N_27817);
xnor UO_634 (O_634,N_29179,N_28225);
xnor UO_635 (O_635,N_28587,N_27191);
xor UO_636 (O_636,N_28177,N_27567);
and UO_637 (O_637,N_29448,N_29762);
nand UO_638 (O_638,N_29328,N_29074);
or UO_639 (O_639,N_27009,N_27319);
nand UO_640 (O_640,N_29250,N_28945);
and UO_641 (O_641,N_28670,N_28779);
nor UO_642 (O_642,N_29859,N_28415);
or UO_643 (O_643,N_29111,N_29870);
nand UO_644 (O_644,N_27313,N_29974);
nand UO_645 (O_645,N_27262,N_29951);
and UO_646 (O_646,N_27062,N_27014);
or UO_647 (O_647,N_27986,N_28364);
nor UO_648 (O_648,N_29511,N_27328);
nand UO_649 (O_649,N_29749,N_28715);
nand UO_650 (O_650,N_28840,N_27898);
nor UO_651 (O_651,N_27410,N_27354);
nor UO_652 (O_652,N_27320,N_28827);
and UO_653 (O_653,N_28219,N_28040);
nand UO_654 (O_654,N_27700,N_29307);
nand UO_655 (O_655,N_29814,N_29709);
nand UO_656 (O_656,N_27711,N_29955);
and UO_657 (O_657,N_29341,N_28864);
and UO_658 (O_658,N_27661,N_27346);
nor UO_659 (O_659,N_29585,N_29945);
or UO_660 (O_660,N_27408,N_28274);
and UO_661 (O_661,N_27637,N_27098);
xor UO_662 (O_662,N_27092,N_29527);
and UO_663 (O_663,N_29481,N_29124);
nor UO_664 (O_664,N_29855,N_27764);
or UO_665 (O_665,N_29268,N_28066);
nor UO_666 (O_666,N_28078,N_29746);
or UO_667 (O_667,N_27046,N_29441);
nand UO_668 (O_668,N_28311,N_28758);
xnor UO_669 (O_669,N_29801,N_28678);
xor UO_670 (O_670,N_28120,N_28036);
or UO_671 (O_671,N_29105,N_29003);
nor UO_672 (O_672,N_28015,N_29916);
or UO_673 (O_673,N_28173,N_28691);
nand UO_674 (O_674,N_29149,N_28195);
nand UO_675 (O_675,N_28488,N_27859);
and UO_676 (O_676,N_28149,N_29626);
nor UO_677 (O_677,N_29897,N_28888);
nor UO_678 (O_678,N_28749,N_27736);
or UO_679 (O_679,N_28393,N_28585);
nor UO_680 (O_680,N_29867,N_29049);
or UO_681 (O_681,N_29248,N_27863);
nor UO_682 (O_682,N_27750,N_28381);
xnor UO_683 (O_683,N_29613,N_27571);
nor UO_684 (O_684,N_29420,N_29491);
xnor UO_685 (O_685,N_27615,N_29320);
nand UO_686 (O_686,N_27041,N_27675);
or UO_687 (O_687,N_29408,N_27106);
nor UO_688 (O_688,N_27364,N_28009);
or UO_689 (O_689,N_28516,N_29624);
or UO_690 (O_690,N_28428,N_27226);
nand UO_691 (O_691,N_28470,N_27460);
nand UO_692 (O_692,N_28058,N_27649);
or UO_693 (O_693,N_27741,N_29222);
nand UO_694 (O_694,N_27234,N_29787);
and UO_695 (O_695,N_29050,N_27429);
nor UO_696 (O_696,N_29789,N_27287);
nand UO_697 (O_697,N_27643,N_29374);
xnor UO_698 (O_698,N_27519,N_27167);
or UO_699 (O_699,N_27728,N_29485);
xnor UO_700 (O_700,N_27890,N_29612);
xnor UO_701 (O_701,N_28637,N_28750);
nand UO_702 (O_702,N_28561,N_27124);
xnor UO_703 (O_703,N_27712,N_28465);
nor UO_704 (O_704,N_29494,N_29662);
nand UO_705 (O_705,N_29166,N_29548);
nor UO_706 (O_706,N_29537,N_29400);
or UO_707 (O_707,N_27265,N_28057);
xnor UO_708 (O_708,N_29167,N_27679);
and UO_709 (O_709,N_27953,N_29549);
nand UO_710 (O_710,N_27026,N_29699);
or UO_711 (O_711,N_27515,N_27832);
or UO_712 (O_712,N_28059,N_28477);
or UO_713 (O_713,N_27005,N_27594);
xnor UO_714 (O_714,N_28355,N_28772);
nand UO_715 (O_715,N_28175,N_28361);
nand UO_716 (O_716,N_29233,N_28089);
and UO_717 (O_717,N_29237,N_28906);
or UO_718 (O_718,N_27146,N_29695);
or UO_719 (O_719,N_28733,N_29028);
nor UO_720 (O_720,N_27894,N_27277);
nand UO_721 (O_721,N_29192,N_29721);
xnor UO_722 (O_722,N_29285,N_29731);
xor UO_723 (O_723,N_27989,N_29823);
nor UO_724 (O_724,N_28529,N_28839);
nand UO_725 (O_725,N_27022,N_29181);
nand UO_726 (O_726,N_29918,N_28365);
nor UO_727 (O_727,N_29224,N_28513);
nor UO_728 (O_728,N_29251,N_27676);
nand UO_729 (O_729,N_28017,N_29589);
or UO_730 (O_730,N_27162,N_29143);
and UO_731 (O_731,N_27959,N_28786);
or UO_732 (O_732,N_27343,N_29322);
or UO_733 (O_733,N_29221,N_28286);
xor UO_734 (O_734,N_27105,N_29134);
xor UO_735 (O_735,N_27723,N_28655);
xnor UO_736 (O_736,N_28042,N_29128);
nand UO_737 (O_737,N_27791,N_27174);
or UO_738 (O_738,N_28341,N_28186);
xnor UO_739 (O_739,N_27215,N_28731);
or UO_740 (O_740,N_29018,N_28726);
nand UO_741 (O_741,N_29308,N_27794);
and UO_742 (O_742,N_27556,N_27382);
xnor UO_743 (O_743,N_29487,N_28373);
and UO_744 (O_744,N_28798,N_28249);
or UO_745 (O_745,N_27744,N_29635);
nor UO_746 (O_746,N_28272,N_27436);
and UO_747 (O_747,N_27267,N_28482);
nor UO_748 (O_748,N_29195,N_28535);
nand UO_749 (O_749,N_27951,N_27248);
nand UO_750 (O_750,N_27003,N_28462);
xor UO_751 (O_751,N_27777,N_29842);
xor UO_752 (O_752,N_28162,N_27668);
xnor UO_753 (O_753,N_28562,N_29036);
and UO_754 (O_754,N_27773,N_29888);
or UO_755 (O_755,N_27618,N_28785);
and UO_756 (O_756,N_29165,N_28862);
or UO_757 (O_757,N_27969,N_29013);
nor UO_758 (O_758,N_27447,N_28417);
nand UO_759 (O_759,N_28531,N_27943);
nor UO_760 (O_760,N_27855,N_28004);
nor UO_761 (O_761,N_29123,N_29282);
xor UO_762 (O_762,N_28984,N_29654);
nor UO_763 (O_763,N_29540,N_28189);
nor UO_764 (O_764,N_28575,N_29121);
nor UO_765 (O_765,N_29270,N_27013);
xnor UO_766 (O_766,N_29327,N_28911);
nor UO_767 (O_767,N_29625,N_28082);
and UO_768 (O_768,N_28964,N_27850);
or UO_769 (O_769,N_27865,N_29212);
xnor UO_770 (O_770,N_27861,N_28279);
nand UO_771 (O_771,N_27434,N_27071);
or UO_772 (O_772,N_28270,N_27072);
xnor UO_773 (O_773,N_28907,N_29080);
xnor UO_774 (O_774,N_28317,N_29587);
and UO_775 (O_775,N_29581,N_27435);
nand UO_776 (O_776,N_28131,N_27960);
xnor UO_777 (O_777,N_29609,N_29550);
or UO_778 (O_778,N_27483,N_27465);
and UO_779 (O_779,N_29574,N_28737);
nand UO_780 (O_780,N_29898,N_29647);
nand UO_781 (O_781,N_28925,N_28489);
xor UO_782 (O_782,N_27603,N_29817);
and UO_783 (O_783,N_28243,N_29189);
nand UO_784 (O_784,N_28698,N_27190);
nor UO_785 (O_785,N_29831,N_28788);
and UO_786 (O_786,N_29023,N_27318);
nor UO_787 (O_787,N_27327,N_28947);
nor UO_788 (O_788,N_28418,N_28974);
xor UO_789 (O_789,N_28138,N_29063);
nor UO_790 (O_790,N_29607,N_28533);
or UO_791 (O_791,N_28612,N_27008);
xnor UO_792 (O_792,N_29186,N_28448);
or UO_793 (O_793,N_28151,N_27024);
and UO_794 (O_794,N_29681,N_27833);
or UO_795 (O_795,N_29939,N_27331);
and UO_796 (O_796,N_27560,N_28499);
nand UO_797 (O_797,N_28899,N_29919);
or UO_798 (O_798,N_29220,N_27422);
nor UO_799 (O_799,N_27573,N_29160);
xor UO_800 (O_800,N_27978,N_27120);
or UO_801 (O_801,N_29973,N_29936);
and UO_802 (O_802,N_27815,N_27139);
nand UO_803 (O_803,N_29474,N_29014);
or UO_804 (O_804,N_27284,N_27998);
xor UO_805 (O_805,N_28628,N_27345);
nand UO_806 (O_806,N_27237,N_28213);
and UO_807 (O_807,N_27821,N_29464);
or UO_808 (O_808,N_29005,N_27935);
nor UO_809 (O_809,N_27141,N_29821);
or UO_810 (O_810,N_27308,N_27646);
xnor UO_811 (O_811,N_29521,N_29498);
xnor UO_812 (O_812,N_29130,N_28580);
and UO_813 (O_813,N_29069,N_29193);
nor UO_814 (O_814,N_27829,N_27027);
nor UO_815 (O_815,N_28519,N_27165);
or UO_816 (O_816,N_29340,N_27387);
xnor UO_817 (O_817,N_28253,N_29674);
xor UO_818 (O_818,N_29425,N_29679);
nor UO_819 (O_819,N_28121,N_28589);
or UO_820 (O_820,N_27407,N_27512);
or UO_821 (O_821,N_27134,N_28928);
nand UO_822 (O_822,N_27530,N_28542);
nor UO_823 (O_823,N_29175,N_27541);
nand UO_824 (O_824,N_27040,N_28872);
xor UO_825 (O_825,N_28244,N_29411);
nor UO_826 (O_826,N_29977,N_28608);
and UO_827 (O_827,N_28056,N_27425);
xnor UO_828 (O_828,N_28830,N_28752);
xor UO_829 (O_829,N_28146,N_27299);
and UO_830 (O_830,N_28883,N_28645);
nand UO_831 (O_831,N_27533,N_27705);
xor UO_832 (O_832,N_28076,N_27342);
and UO_833 (O_833,N_28844,N_29999);
nor UO_834 (O_834,N_27642,N_29155);
and UO_835 (O_835,N_27891,N_27104);
nor UO_836 (O_836,N_27150,N_27018);
and UO_837 (O_837,N_27325,N_28613);
or UO_838 (O_838,N_28282,N_27423);
and UO_839 (O_839,N_29294,N_29048);
nor UO_840 (O_840,N_28475,N_27685);
or UO_841 (O_841,N_28294,N_27752);
and UO_842 (O_842,N_28130,N_27143);
xor UO_843 (O_843,N_27666,N_27254);
or UO_844 (O_844,N_29546,N_29118);
and UO_845 (O_845,N_28983,N_27786);
xor UO_846 (O_846,N_29228,N_29303);
xnor UO_847 (O_847,N_29712,N_29783);
or UO_848 (O_848,N_27412,N_29688);
nand UO_849 (O_849,N_28293,N_29708);
nor UO_850 (O_850,N_27763,N_27455);
nand UO_851 (O_851,N_29767,N_28771);
nand UO_852 (O_852,N_27017,N_28674);
nor UO_853 (O_853,N_28386,N_27274);
xor UO_854 (O_854,N_29236,N_28379);
xor UO_855 (O_855,N_27823,N_29422);
xor UO_856 (O_856,N_28438,N_29372);
and UO_857 (O_857,N_27677,N_29748);
nand UO_858 (O_858,N_29398,N_29084);
and UO_859 (O_859,N_27802,N_29755);
nor UO_860 (O_860,N_27730,N_27856);
or UO_861 (O_861,N_28112,N_27135);
nand UO_862 (O_862,N_29265,N_28634);
nand UO_863 (O_863,N_29336,N_27577);
and UO_864 (O_864,N_27437,N_29276);
xor UO_865 (O_865,N_28741,N_29466);
nor UO_866 (O_866,N_27735,N_27973);
or UO_867 (O_867,N_28184,N_27445);
or UO_868 (O_868,N_28239,N_28537);
or UO_869 (O_869,N_29685,N_27724);
and UO_870 (O_870,N_28970,N_29357);
xor UO_871 (O_871,N_27940,N_29794);
nor UO_872 (O_872,N_29673,N_27589);
nand UO_873 (O_873,N_29044,N_27770);
xnor UO_874 (O_874,N_28178,N_29661);
nor UO_875 (O_875,N_29653,N_27279);
nor UO_876 (O_876,N_28496,N_27131);
xnor UO_877 (O_877,N_28164,N_27479);
nand UO_878 (O_878,N_29592,N_28008);
nor UO_879 (O_879,N_29663,N_28842);
nand UO_880 (O_880,N_28307,N_29525);
and UO_881 (O_881,N_29641,N_28136);
xor UO_882 (O_882,N_29987,N_29072);
and UO_883 (O_883,N_29393,N_27438);
nand UO_884 (O_884,N_29657,N_28654);
or UO_885 (O_885,N_27194,N_27087);
and UO_886 (O_886,N_28023,N_28366);
xor UO_887 (O_887,N_28530,N_28917);
nand UO_888 (O_888,N_27091,N_27401);
and UO_889 (O_889,N_28763,N_28706);
xor UO_890 (O_890,N_27232,N_28399);
or UO_891 (O_891,N_27531,N_29047);
or UO_892 (O_892,N_27938,N_28469);
nand UO_893 (O_893,N_28022,N_27897);
or UO_894 (O_894,N_28060,N_28663);
nor UO_895 (O_895,N_28401,N_29395);
and UO_896 (O_896,N_29927,N_27409);
and UO_897 (O_897,N_29672,N_29791);
and UO_898 (O_898,N_29851,N_29053);
nand UO_899 (O_899,N_28125,N_27166);
or UO_900 (O_900,N_27456,N_29617);
and UO_901 (O_901,N_27377,N_27424);
or UO_902 (O_902,N_29706,N_27394);
nor UO_903 (O_903,N_29876,N_27349);
and UO_904 (O_904,N_29174,N_27605);
nand UO_905 (O_905,N_28443,N_29885);
xnor UO_906 (O_906,N_27183,N_28804);
nor UO_907 (O_907,N_28347,N_28611);
xnor UO_908 (O_908,N_27075,N_29590);
xor UO_909 (O_909,N_28505,N_27123);
xnor UO_910 (O_910,N_29530,N_28085);
and UO_911 (O_911,N_27063,N_28831);
nor UO_912 (O_912,N_29459,N_28803);
and UO_913 (O_913,N_27378,N_27238);
or UO_914 (O_914,N_29065,N_28362);
nand UO_915 (O_915,N_28673,N_28006);
xnor UO_916 (O_916,N_27559,N_27163);
xor UO_917 (O_917,N_28506,N_29075);
nand UO_918 (O_918,N_27454,N_29421);
or UO_919 (O_919,N_27099,N_28455);
or UO_920 (O_920,N_28859,N_29793);
nor UO_921 (O_921,N_29330,N_27684);
and UO_922 (O_922,N_29156,N_28932);
and UO_923 (O_923,N_28781,N_28975);
nor UO_924 (O_924,N_27738,N_27073);
nand UO_925 (O_925,N_28264,N_29912);
and UO_926 (O_926,N_29928,N_27369);
nor UO_927 (O_927,N_28896,N_27776);
nor UO_928 (O_928,N_27235,N_27846);
nor UO_929 (O_929,N_28237,N_27983);
and UO_930 (O_930,N_29792,N_27207);
or UO_931 (O_931,N_29515,N_27772);
xnor UO_932 (O_932,N_27228,N_29199);
and UO_933 (O_933,N_29599,N_27142);
nand UO_934 (O_934,N_27792,N_28738);
and UO_935 (O_935,N_28568,N_28672);
and UO_936 (O_936,N_28413,N_28153);
nor UO_937 (O_937,N_29126,N_29465);
nand UO_938 (O_938,N_28464,N_29461);
xor UO_939 (O_939,N_28761,N_28220);
nor UO_940 (O_940,N_27886,N_28881);
and UO_941 (O_941,N_29553,N_27799);
or UO_942 (O_942,N_29107,N_27468);
xor UO_943 (O_943,N_27294,N_27032);
nor UO_944 (O_944,N_27701,N_29786);
xnor UO_945 (O_945,N_27586,N_27180);
nor UO_946 (O_946,N_27196,N_28383);
and UO_947 (O_947,N_27828,N_29208);
or UO_948 (O_948,N_28936,N_29055);
or UO_949 (O_949,N_27775,N_27783);
nor UO_950 (O_950,N_29424,N_29415);
nand UO_951 (O_951,N_28524,N_29915);
nor UO_952 (O_952,N_29669,N_29556);
and UO_953 (O_953,N_29438,N_27547);
and UO_954 (O_954,N_28388,N_28597);
nor UO_955 (O_955,N_28920,N_28436);
xor UO_956 (O_956,N_29369,N_28232);
or UO_957 (O_957,N_27925,N_27553);
nor UO_958 (O_958,N_27627,N_29178);
nor UO_959 (O_959,N_29723,N_29287);
nand UO_960 (O_960,N_28913,N_28525);
and UO_961 (O_961,N_27473,N_28329);
and UO_962 (O_962,N_27255,N_28328);
or UO_963 (O_963,N_27268,N_29538);
or UO_964 (O_964,N_28179,N_28257);
nand UO_965 (O_965,N_27689,N_27186);
or UO_966 (O_966,N_27795,N_27484);
nand UO_967 (O_967,N_27090,N_28912);
xnor UO_968 (O_968,N_27665,N_27306);
nor UO_969 (O_969,N_28775,N_28514);
nand UO_970 (O_970,N_29517,N_27671);
and UO_971 (O_971,N_28271,N_28777);
xnor UO_972 (O_972,N_29252,N_28716);
xnor UO_973 (O_973,N_27830,N_28431);
xor UO_974 (O_974,N_29064,N_27582);
and UO_975 (O_975,N_29359,N_29719);
and UO_976 (O_976,N_27599,N_27076);
nor UO_977 (O_977,N_27754,N_27466);
or UO_978 (O_978,N_27906,N_29601);
or UO_979 (O_979,N_28133,N_27703);
nor UO_980 (O_980,N_29470,N_28266);
nor UO_981 (O_981,N_28986,N_29445);
nor UO_982 (O_982,N_28450,N_29904);
xnor UO_983 (O_983,N_28254,N_28385);
nand UO_984 (O_984,N_28288,N_28662);
nand UO_985 (O_985,N_29872,N_28053);
xor UO_986 (O_986,N_29943,N_28934);
nor UO_987 (O_987,N_27181,N_27185);
or UO_988 (O_988,N_29761,N_29750);
nor UO_989 (O_989,N_29850,N_29535);
nand UO_990 (O_990,N_27625,N_28606);
or UO_991 (O_991,N_27981,N_28555);
nor UO_992 (O_992,N_27100,N_28631);
and UO_993 (O_993,N_27516,N_28572);
nand UO_994 (O_994,N_29650,N_28823);
and UO_995 (O_995,N_29239,N_28340);
xnor UO_996 (O_996,N_28854,N_28029);
or UO_997 (O_997,N_28787,N_29116);
and UO_998 (O_998,N_28972,N_28992);
xnor UO_999 (O_999,N_28695,N_29475);
or UO_1000 (O_1000,N_28427,N_28390);
nand UO_1001 (O_1001,N_27096,N_29243);
nand UO_1002 (O_1002,N_27654,N_27994);
xor UO_1003 (O_1003,N_28829,N_27638);
nand UO_1004 (O_1004,N_29488,N_28296);
xnor UO_1005 (O_1005,N_27872,N_29246);
xor UO_1006 (O_1006,N_29025,N_27250);
or UO_1007 (O_1007,N_29894,N_28500);
and UO_1008 (O_1008,N_29822,N_27826);
nand UO_1009 (O_1009,N_29337,N_28801);
xor UO_1010 (O_1010,N_29015,N_27563);
nor UO_1011 (O_1011,N_28202,N_27060);
nor UO_1012 (O_1012,N_29261,N_28596);
or UO_1013 (O_1013,N_29727,N_28312);
or UO_1014 (O_1014,N_28545,N_27706);
xor UO_1015 (O_1015,N_28717,N_28493);
and UO_1016 (O_1016,N_27200,N_27083);
or UO_1017 (O_1017,N_29827,N_27384);
or UO_1018 (O_1018,N_27177,N_28495);
or UO_1019 (O_1019,N_27946,N_27269);
xnor UO_1020 (O_1020,N_28739,N_28578);
and UO_1021 (O_1021,N_27006,N_29877);
nor UO_1022 (O_1022,N_29259,N_27975);
nor UO_1023 (O_1023,N_28690,N_29602);
nor UO_1024 (O_1024,N_29932,N_28759);
and UO_1025 (O_1025,N_29288,N_29066);
and UO_1026 (O_1026,N_29682,N_28689);
and UO_1027 (O_1027,N_28723,N_29737);
xor UO_1028 (O_1028,N_27326,N_29201);
xor UO_1029 (O_1029,N_28486,N_28764);
nor UO_1030 (O_1030,N_27584,N_27118);
nor UO_1031 (O_1031,N_29200,N_27451);
or UO_1032 (O_1032,N_27678,N_27413);
and UO_1033 (O_1033,N_28671,N_29094);
nor UO_1034 (O_1034,N_29800,N_28333);
nor UO_1035 (O_1035,N_28895,N_29098);
nor UO_1036 (O_1036,N_28957,N_29988);
nor UO_1037 (O_1037,N_27604,N_27892);
xnor UO_1038 (O_1038,N_28588,N_29145);
xnor UO_1039 (O_1039,N_27532,N_27030);
xor UO_1040 (O_1040,N_28565,N_28960);
and UO_1041 (O_1041,N_29816,N_28855);
nand UO_1042 (O_1042,N_28382,N_28122);
nor UO_1043 (O_1043,N_27725,N_29901);
nand UO_1044 (O_1044,N_29135,N_28437);
xor UO_1045 (O_1045,N_29534,N_27645);
nor UO_1046 (O_1046,N_27246,N_27427);
and UO_1047 (O_1047,N_29054,N_28256);
or UO_1048 (O_1048,N_27623,N_27543);
nand UO_1049 (O_1049,N_29524,N_28660);
xor UO_1050 (O_1050,N_27787,N_29980);
xor UO_1051 (O_1051,N_27885,N_29862);
and UO_1052 (O_1052,N_29052,N_28591);
nor UO_1053 (O_1053,N_28093,N_29455);
or UO_1054 (O_1054,N_29529,N_27521);
xnor UO_1055 (O_1055,N_28626,N_29183);
nor UO_1056 (O_1056,N_28794,N_29443);
xor UO_1057 (O_1057,N_27715,N_29452);
nand UO_1058 (O_1058,N_28097,N_29514);
nor UO_1059 (O_1059,N_29190,N_27101);
and UO_1060 (O_1060,N_28020,N_29355);
and UO_1061 (O_1061,N_29291,N_29317);
xnor UO_1062 (O_1062,N_29979,N_27600);
xnor UO_1063 (O_1063,N_27545,N_28037);
or UO_1064 (O_1064,N_27908,N_29204);
and UO_1065 (O_1065,N_28128,N_28419);
or UO_1066 (O_1066,N_28601,N_28667);
nor UO_1067 (O_1067,N_27048,N_29754);
nor UO_1068 (O_1068,N_28988,N_29214);
nand UO_1069 (O_1069,N_27952,N_29983);
nor UO_1070 (O_1070,N_29720,N_29560);
nor UO_1071 (O_1071,N_27644,N_27272);
nand UO_1072 (O_1072,N_28234,N_28067);
xnor UO_1073 (O_1073,N_29133,N_29804);
xor UO_1074 (O_1074,N_29839,N_27990);
nor UO_1075 (O_1075,N_27510,N_28391);
and UO_1076 (O_1076,N_28479,N_28445);
nor UO_1077 (O_1077,N_29386,N_28664);
nand UO_1078 (O_1078,N_29971,N_29215);
and UO_1079 (O_1079,N_28592,N_27619);
xor UO_1080 (O_1080,N_27497,N_28224);
or UO_1081 (O_1081,N_29845,N_29835);
and UO_1082 (O_1082,N_28604,N_29752);
xnor UO_1083 (O_1083,N_29122,N_27373);
nand UO_1084 (O_1084,N_29403,N_27769);
or UO_1085 (O_1085,N_27987,N_27911);
nand UO_1086 (O_1086,N_29046,N_27804);
nand UO_1087 (O_1087,N_29701,N_29738);
and UO_1088 (O_1088,N_29260,N_28319);
and UO_1089 (O_1089,N_29034,N_27527);
nor UO_1090 (O_1090,N_29561,N_28210);
or UO_1091 (O_1091,N_28463,N_27868);
xnor UO_1092 (O_1092,N_29350,N_28916);
nor UO_1093 (O_1093,N_27074,N_29206);
or UO_1094 (O_1094,N_27805,N_29348);
nand UO_1095 (O_1095,N_27811,N_28808);
or UO_1096 (O_1096,N_28165,N_29318);
xor UO_1097 (O_1097,N_29948,N_27837);
nor UO_1098 (O_1098,N_29820,N_29417);
or UO_1099 (O_1099,N_28643,N_29559);
xnor UO_1100 (O_1100,N_29451,N_29062);
xnor UO_1101 (O_1101,N_29147,N_28728);
or UO_1102 (O_1102,N_29071,N_27157);
and UO_1103 (O_1103,N_27380,N_28452);
xor UO_1104 (O_1104,N_29437,N_29740);
nor UO_1105 (O_1105,N_28468,N_28086);
xnor UO_1106 (O_1106,N_27900,N_27350);
nand UO_1107 (O_1107,N_27709,N_28991);
xor UO_1108 (O_1108,N_29790,N_27945);
nand UO_1109 (O_1109,N_28372,N_27430);
nor UO_1110 (O_1110,N_27158,N_28354);
or UO_1111 (O_1111,N_28193,N_27580);
and UO_1112 (O_1112,N_29271,N_27112);
nand UO_1113 (O_1113,N_29763,N_29070);
nand UO_1114 (O_1114,N_27095,N_28407);
nor UO_1115 (O_1115,N_27910,N_27609);
nand UO_1116 (O_1116,N_28756,N_27598);
nand UO_1117 (O_1117,N_27414,N_29715);
nand UO_1118 (O_1118,N_28722,N_27688);
nor UO_1119 (O_1119,N_29848,N_27964);
nand UO_1120 (O_1120,N_27390,N_28028);
nor UO_1121 (O_1121,N_29900,N_27307);
nand UO_1122 (O_1122,N_27972,N_28600);
nor UO_1123 (O_1123,N_28422,N_27996);
nand UO_1124 (O_1124,N_29313,N_28273);
nor UO_1125 (O_1125,N_28106,N_27659);
nand UO_1126 (O_1126,N_27285,N_27315);
nor UO_1127 (O_1127,N_27474,N_28543);
and UO_1128 (O_1128,N_28152,N_28571);
xnor UO_1129 (O_1129,N_29334,N_27001);
nand UO_1130 (O_1130,N_29255,N_28806);
and UO_1131 (O_1131,N_29802,N_28000);
or UO_1132 (O_1132,N_28230,N_29722);
nand UO_1133 (O_1133,N_27674,N_27029);
nand UO_1134 (O_1134,N_29326,N_29434);
xnor UO_1135 (O_1135,N_28943,N_29253);
and UO_1136 (O_1136,N_29381,N_27767);
nor UO_1137 (O_1137,N_28031,N_27926);
nor UO_1138 (O_1138,N_29809,N_28630);
nor UO_1139 (O_1139,N_28989,N_28646);
or UO_1140 (O_1140,N_29853,N_29946);
and UO_1141 (O_1141,N_27302,N_28753);
and UO_1142 (O_1142,N_29095,N_29966);
nor UO_1143 (O_1143,N_28619,N_29849);
nor UO_1144 (O_1144,N_28050,N_27845);
or UO_1145 (O_1145,N_29019,N_28847);
xnor UO_1146 (O_1146,N_27881,N_28218);
nand UO_1147 (O_1147,N_28100,N_28748);
nand UO_1148 (O_1148,N_27895,N_29873);
xnor UO_1149 (O_1149,N_27942,N_27683);
xor UO_1150 (O_1150,N_29998,N_29457);
nand UO_1151 (O_1151,N_28343,N_28981);
and UO_1152 (O_1152,N_27310,N_28696);
nand UO_1153 (O_1153,N_29394,N_29523);
and UO_1154 (O_1154,N_28697,N_29508);
xor UO_1155 (O_1155,N_28743,N_27967);
nand UO_1156 (O_1156,N_29779,N_29580);
nand UO_1157 (O_1157,N_29439,N_29002);
nor UO_1158 (O_1158,N_29188,N_29109);
nor UO_1159 (O_1159,N_28693,N_29596);
or UO_1160 (O_1160,N_28621,N_29202);
xor UO_1161 (O_1161,N_29890,N_27418);
xnor UO_1162 (O_1162,N_27835,N_29828);
nand UO_1163 (O_1163,N_28073,N_29405);
nor UO_1164 (O_1164,N_27153,N_29035);
nor UO_1165 (O_1165,N_29743,N_28747);
nor UO_1166 (O_1166,N_27647,N_29364);
and UO_1167 (O_1167,N_29776,N_27000);
or UO_1168 (O_1168,N_28848,N_28725);
nor UO_1169 (O_1169,N_27381,N_28503);
nor UO_1170 (O_1170,N_27624,N_29994);
xor UO_1171 (O_1171,N_28035,N_27292);
xor UO_1172 (O_1172,N_29907,N_28766);
and UO_1173 (O_1173,N_29203,N_28700);
or UO_1174 (O_1174,N_28169,N_27739);
xor UO_1175 (O_1175,N_27572,N_28857);
xor UO_1176 (O_1176,N_29375,N_27708);
xor UO_1177 (O_1177,N_29526,N_28534);
xor UO_1178 (O_1178,N_28918,N_27336);
and UO_1179 (O_1179,N_28824,N_29756);
or UO_1180 (O_1180,N_27069,N_29500);
xnor UO_1181 (O_1181,N_27127,N_27982);
and UO_1182 (O_1182,N_29113,N_29680);
or UO_1183 (O_1183,N_27949,N_27417);
or UO_1184 (O_1184,N_28113,N_27411);
and UO_1185 (O_1185,N_28853,N_27720);
xnor UO_1186 (O_1186,N_28071,N_28327);
xnor UO_1187 (O_1187,N_29363,N_28521);
and UO_1188 (O_1188,N_27187,N_29645);
xor UO_1189 (O_1189,N_28939,N_29286);
xor UO_1190 (O_1190,N_28116,N_28302);
nand UO_1191 (O_1191,N_27016,N_27740);
nor UO_1192 (O_1192,N_27916,N_27368);
nor UO_1193 (O_1193,N_29402,N_27251);
and UO_1194 (O_1194,N_29642,N_28476);
nor UO_1195 (O_1195,N_29917,N_28441);
nand UO_1196 (O_1196,N_28182,N_28039);
nand UO_1197 (O_1197,N_27847,N_29714);
xor UO_1198 (O_1198,N_27217,N_28108);
or UO_1199 (O_1199,N_29769,N_27797);
nand UO_1200 (O_1200,N_29504,N_29366);
or UO_1201 (O_1201,N_28817,N_27229);
xnor UO_1202 (O_1202,N_29283,N_29319);
xnor UO_1203 (O_1203,N_27482,N_29138);
nand UO_1204 (O_1204,N_29273,N_27080);
and UO_1205 (O_1205,N_29728,N_27919);
xnor UO_1206 (O_1206,N_27824,N_28405);
nor UO_1207 (O_1207,N_27924,N_29902);
nor UO_1208 (O_1208,N_27353,N_28869);
or UO_1209 (O_1209,N_27534,N_28016);
nor UO_1210 (O_1210,N_29651,N_29150);
and UO_1211 (O_1211,N_27733,N_29412);
nand UO_1212 (O_1212,N_28836,N_29472);
nand UO_1213 (O_1213,N_28052,N_28528);
xor UO_1214 (O_1214,N_29042,N_28492);
nand UO_1215 (O_1215,N_28483,N_29956);
xor UO_1216 (O_1216,N_28091,N_27544);
xor UO_1217 (O_1217,N_29598,N_27300);
nand UO_1218 (O_1218,N_27879,N_28579);
nor UO_1219 (O_1219,N_27082,N_28729);
or UO_1220 (O_1220,N_29339,N_29531);
nor UO_1221 (O_1221,N_28375,N_27613);
and UO_1222 (O_1222,N_28713,N_29159);
and UO_1223 (O_1223,N_27399,N_27611);
or UO_1224 (O_1224,N_28054,N_28174);
and UO_1225 (O_1225,N_28241,N_27529);
xnor UO_1226 (O_1226,N_27259,N_28305);
nand UO_1227 (O_1227,N_27137,N_29315);
nand UO_1228 (O_1228,N_29463,N_28581);
or UO_1229 (O_1229,N_27208,N_29258);
and UO_1230 (O_1230,N_29782,N_27601);
xor UO_1231 (O_1231,N_29841,N_29247);
xor UO_1232 (O_1232,N_27593,N_27873);
nand UO_1233 (O_1233,N_27107,N_29751);
nand UO_1234 (O_1234,N_28954,N_29501);
or UO_1235 (O_1235,N_28158,N_28092);
xor UO_1236 (O_1236,N_28576,N_28985);
nor UO_1237 (O_1237,N_29254,N_29227);
nor UO_1238 (O_1238,N_29620,N_29964);
xnor UO_1239 (O_1239,N_27240,N_28246);
nor UO_1240 (O_1240,N_29656,N_29469);
or UO_1241 (O_1241,N_28055,N_28641);
nand UO_1242 (O_1242,N_29933,N_28176);
and UO_1243 (O_1243,N_28504,N_27077);
or UO_1244 (O_1244,N_29077,N_29148);
nand UO_1245 (O_1245,N_27931,N_27055);
nor UO_1246 (O_1246,N_27244,N_28227);
nand UO_1247 (O_1247,N_27913,N_28275);
nand UO_1248 (O_1248,N_29564,N_29480);
nor UO_1249 (O_1249,N_28331,N_27303);
or UO_1250 (O_1250,N_29033,N_28835);
nor UO_1251 (O_1251,N_28625,N_29950);
xnor UO_1252 (O_1252,N_28998,N_28242);
nor UO_1253 (O_1253,N_27195,N_27570);
and UO_1254 (O_1254,N_28963,N_28188);
nand UO_1255 (O_1255,N_27596,N_29803);
xor UO_1256 (O_1256,N_29368,N_28430);
nand UO_1257 (O_1257,N_29311,N_29869);
nor UO_1258 (O_1258,N_28211,N_28941);
or UO_1259 (O_1259,N_29305,N_27965);
or UO_1260 (O_1260,N_29471,N_27464);
xor UO_1261 (O_1261,N_29633,N_29671);
xnor UO_1262 (O_1262,N_28507,N_28233);
or UO_1263 (O_1263,N_28150,N_29168);
nand UO_1264 (O_1264,N_27052,N_28318);
xor UO_1265 (O_1265,N_27461,N_27457);
or UO_1266 (O_1266,N_28971,N_28321);
nand UO_1267 (O_1267,N_28948,N_27551);
or UO_1268 (O_1268,N_28688,N_29284);
nand UO_1269 (O_1269,N_28714,N_27522);
xor UO_1270 (O_1270,N_28041,N_27818);
nand UO_1271 (O_1271,N_28653,N_27766);
nor UO_1272 (O_1272,N_27053,N_29759);
xnor UO_1273 (O_1273,N_28675,N_27607);
xnor UO_1274 (O_1274,N_27441,N_29583);
nor UO_1275 (O_1275,N_28719,N_28068);
and UO_1276 (O_1276,N_28359,N_29040);
or UO_1277 (O_1277,N_29078,N_29117);
xor UO_1278 (O_1278,N_28221,N_27367);
or UO_1279 (O_1279,N_29604,N_28993);
and UO_1280 (O_1280,N_29306,N_27039);
nor UO_1281 (O_1281,N_28546,N_28828);
xor UO_1282 (O_1282,N_29726,N_27930);
xnor UO_1283 (O_1283,N_27440,N_29162);
and UO_1284 (O_1284,N_29389,N_28160);
or UO_1285 (O_1285,N_28064,N_27110);
and UO_1286 (O_1286,N_28962,N_28605);
or UO_1287 (O_1287,N_28269,N_29213);
or UO_1288 (O_1288,N_29490,N_28799);
xnor UO_1289 (O_1289,N_27883,N_28196);
and UO_1290 (O_1290,N_27431,N_28517);
and UO_1291 (O_1291,N_28999,N_28013);
xnor UO_1292 (O_1292,N_29572,N_29836);
and UO_1293 (O_1293,N_29970,N_29068);
nor UO_1294 (O_1294,N_28109,N_29586);
nand UO_1295 (O_1295,N_27329,N_28228);
nand UO_1296 (O_1296,N_27687,N_29454);
or UO_1297 (O_1297,N_29030,N_27536);
or UO_1298 (O_1298,N_27312,N_27957);
and UO_1299 (O_1299,N_27583,N_28685);
or UO_1300 (O_1300,N_29127,N_28875);
xor UO_1301 (O_1301,N_27184,N_27147);
nor UO_1302 (O_1302,N_28247,N_28498);
nor UO_1303 (O_1303,N_28005,N_27956);
nand UO_1304 (O_1304,N_27686,N_29316);
xnor UO_1305 (O_1305,N_28811,N_27501);
nor UO_1306 (O_1306,N_27375,N_27592);
xnor UO_1307 (O_1307,N_28933,N_29634);
or UO_1308 (O_1308,N_29579,N_27539);
xor UO_1309 (O_1309,N_29942,N_29593);
or UO_1310 (O_1310,N_28890,N_29484);
nand UO_1311 (O_1311,N_27877,N_27219);
nor UO_1312 (O_1312,N_29505,N_27119);
nand UO_1313 (O_1313,N_28276,N_29290);
xor UO_1314 (O_1314,N_29510,N_28342);
xnor UO_1315 (O_1315,N_29478,N_29995);
or UO_1316 (O_1316,N_28909,N_27498);
nor UO_1317 (O_1317,N_27812,N_28676);
and UO_1318 (O_1318,N_27359,N_29293);
xor UO_1319 (O_1319,N_27028,N_29001);
xnor UO_1320 (O_1320,N_28712,N_28882);
nand UO_1321 (O_1321,N_28990,N_27760);
xnor UO_1322 (O_1322,N_29678,N_28204);
nand UO_1323 (O_1323,N_27920,N_27064);
or UO_1324 (O_1324,N_29093,N_28871);
nand UO_1325 (O_1325,N_29610,N_27581);
or UO_1326 (O_1326,N_27503,N_28682);
nand UO_1327 (O_1327,N_29144,N_27253);
or UO_1328 (O_1328,N_29362,N_29120);
xnor UO_1329 (O_1329,N_28485,N_29266);
nor UO_1330 (O_1330,N_29558,N_29157);
xor UO_1331 (O_1331,N_28474,N_29753);
and UO_1332 (O_1332,N_29807,N_29497);
xor UO_1333 (O_1333,N_28867,N_29666);
and UO_1334 (O_1334,N_27415,N_27111);
xnor UO_1335 (O_1335,N_28515,N_29705);
or UO_1336 (O_1336,N_29216,N_27321);
or UO_1337 (O_1337,N_27061,N_29905);
and UO_1338 (O_1338,N_27755,N_27406);
xor UO_1339 (O_1339,N_27853,N_29061);
nand UO_1340 (O_1340,N_27555,N_29773);
nand UO_1341 (O_1341,N_28699,N_28170);
xor UO_1342 (O_1342,N_27149,N_27732);
xnor UO_1343 (O_1343,N_27210,N_29088);
nand UO_1344 (O_1344,N_27103,N_27670);
and UO_1345 (O_1345,N_29089,N_27542);
or UO_1346 (O_1346,N_27941,N_27043);
nand UO_1347 (O_1347,N_27220,N_28760);
or UO_1348 (O_1348,N_27511,N_28472);
or UO_1349 (O_1349,N_28449,N_29081);
and UO_1350 (O_1350,N_28980,N_29810);
nor UO_1351 (O_1351,N_27266,N_29632);
and UO_1352 (O_1352,N_29433,N_27264);
nor UO_1353 (O_1353,N_28166,N_29370);
or UO_1354 (O_1354,N_27974,N_28466);
nor UO_1355 (O_1355,N_28335,N_27682);
and UO_1356 (O_1356,N_27452,N_27834);
or UO_1357 (O_1357,N_27293,N_27160);
xor UO_1358 (O_1358,N_28180,N_29861);
and UO_1359 (O_1359,N_28141,N_28573);
xor UO_1360 (O_1360,N_27825,N_29940);
xor UO_1361 (O_1361,N_27370,N_27860);
and UO_1362 (O_1362,N_28201,N_28973);
nor UO_1363 (O_1363,N_28669,N_29684);
nor UO_1364 (O_1364,N_29037,N_27033);
and UO_1365 (O_1365,N_29277,N_27652);
or UO_1366 (O_1366,N_29911,N_28456);
and UO_1367 (O_1367,N_28532,N_29772);
xor UO_1368 (O_1368,N_29914,N_28701);
nor UO_1369 (O_1369,N_27480,N_28889);
xor UO_1370 (O_1370,N_27463,N_29687);
xnor UO_1371 (O_1371,N_27398,N_29806);
or UO_1372 (O_1372,N_28471,N_29777);
nor UO_1373 (O_1373,N_28644,N_27997);
nor UO_1374 (O_1374,N_27576,N_27757);
nand UO_1375 (O_1375,N_29757,N_28338);
and UO_1376 (O_1376,N_27038,N_28183);
or UO_1377 (O_1377,N_29993,N_28636);
xnor UO_1378 (O_1378,N_27247,N_29056);
nor UO_1379 (O_1379,N_27470,N_29397);
nand UO_1380 (O_1380,N_28540,N_27554);
and UO_1381 (O_1381,N_29856,N_28245);
and UO_1382 (O_1382,N_29509,N_29958);
xor UO_1383 (O_1383,N_28805,N_29608);
xor UO_1384 (O_1384,N_27421,N_29039);
and UO_1385 (O_1385,N_29231,N_29269);
and UO_1386 (O_1386,N_27204,N_29545);
nor UO_1387 (O_1387,N_29087,N_29611);
and UO_1388 (O_1388,N_27991,N_29864);
or UO_1389 (O_1389,N_29241,N_28453);
nand UO_1390 (O_1390,N_27403,N_27564);
nand UO_1391 (O_1391,N_28081,N_27323);
or UO_1392 (O_1392,N_27507,N_29832);
and UO_1393 (O_1393,N_27125,N_29838);
and UO_1394 (O_1394,N_27304,N_28212);
or UO_1395 (O_1395,N_27820,N_29353);
or UO_1396 (O_1396,N_28451,N_29153);
nand UO_1397 (O_1397,N_27803,N_29097);
and UO_1398 (O_1398,N_27719,N_28767);
nand UO_1399 (O_1399,N_29725,N_27672);
xor UO_1400 (O_1400,N_29458,N_29766);
nand UO_1401 (O_1401,N_28639,N_28421);
nor UO_1402 (O_1402,N_28190,N_28061);
or UO_1403 (O_1403,N_28104,N_28290);
or UO_1404 (O_1404,N_29032,N_27154);
and UO_1405 (O_1405,N_29703,N_28295);
xor UO_1406 (O_1406,N_28846,N_27718);
and UO_1407 (O_1407,N_29690,N_27488);
or UO_1408 (O_1408,N_27669,N_29456);
nor UO_1409 (O_1409,N_29758,N_27295);
nor UO_1410 (O_1410,N_29263,N_27562);
nor UO_1411 (O_1411,N_28860,N_27893);
nand UO_1412 (O_1412,N_28062,N_29169);
or UO_1413 (O_1413,N_27065,N_28810);
and UO_1414 (O_1414,N_28898,N_28357);
or UO_1415 (O_1415,N_27023,N_27524);
or UO_1416 (O_1416,N_29108,N_28099);
nand UO_1417 (O_1417,N_29522,N_27636);
nand UO_1418 (O_1418,N_29008,N_28650);
xnor UO_1419 (O_1419,N_29011,N_28539);
xnor UO_1420 (O_1420,N_29588,N_28740);
nand UO_1421 (O_1421,N_27459,N_29142);
and UO_1422 (O_1422,N_29462,N_27585);
nor UO_1423 (O_1423,N_28593,N_27085);
or UO_1424 (O_1424,N_27993,N_29131);
nand UO_1425 (O_1425,N_29784,N_28987);
nand UO_1426 (O_1426,N_29507,N_28396);
or UO_1427 (O_1427,N_29492,N_27057);
nor UO_1428 (O_1428,N_28841,N_27144);
xor UO_1429 (O_1429,N_28145,N_27858);
nor UO_1430 (O_1430,N_28156,N_29829);
nand UO_1431 (O_1431,N_29963,N_28551);
or UO_1432 (O_1432,N_29944,N_27221);
nand UO_1433 (O_1433,N_27504,N_27839);
nor UO_1434 (O_1434,N_29399,N_29930);
or UO_1435 (O_1435,N_28154,N_28711);
nor UO_1436 (O_1436,N_29648,N_27758);
xor UO_1437 (O_1437,N_29384,N_28926);
or UO_1438 (O_1438,N_29623,N_28567);
nor UO_1439 (O_1439,N_29219,N_27317);
and UO_1440 (O_1440,N_28858,N_29163);
or UO_1441 (O_1441,N_27690,N_29765);
or UO_1442 (O_1442,N_28314,N_27446);
and UO_1443 (O_1443,N_27467,N_27130);
nor UO_1444 (O_1444,N_27198,N_27054);
nand UO_1445 (O_1445,N_28394,N_29082);
and UO_1446 (O_1446,N_28703,N_29947);
and UO_1447 (O_1447,N_29377,N_29428);
and UO_1448 (O_1448,N_27156,N_28707);
nor UO_1449 (O_1449,N_28123,N_27927);
nand UO_1450 (O_1450,N_28845,N_27224);
nand UO_1451 (O_1451,N_27444,N_29830);
nand UO_1452 (O_1452,N_28523,N_27178);
xnor UO_1453 (O_1453,N_27590,N_29686);
and UO_1454 (O_1454,N_28979,N_28461);
and UO_1455 (O_1455,N_28267,N_28966);
xor UO_1456 (O_1456,N_29778,N_29961);
xor UO_1457 (O_1457,N_29908,N_29584);
nor UO_1458 (O_1458,N_28101,N_27442);
or UO_1459 (O_1459,N_28426,N_29010);
or UO_1460 (O_1460,N_29365,N_29785);
nand UO_1461 (O_1461,N_28520,N_29342);
xnor UO_1462 (O_1462,N_27236,N_28651);
nand UO_1463 (O_1463,N_28553,N_29194);
nor UO_1464 (O_1464,N_27851,N_27896);
nand UO_1465 (O_1465,N_27152,N_27520);
nor UO_1466 (O_1466,N_27242,N_28583);
nand UO_1467 (O_1467,N_29874,N_28745);
nand UO_1468 (O_1468,N_27681,N_27297);
and UO_1469 (O_1469,N_27784,N_28905);
and UO_1470 (O_1470,N_28893,N_29022);
nor UO_1471 (O_1471,N_28902,N_28826);
xnor UO_1472 (O_1472,N_28191,N_27918);
xor UO_1473 (O_1473,N_29863,N_29198);
or UO_1474 (O_1474,N_29431,N_27535);
or UO_1475 (O_1475,N_28079,N_27395);
xnor UO_1476 (O_1476,N_28297,N_28550);
xor UO_1477 (O_1477,N_29016,N_27396);
nor UO_1478 (O_1478,N_27070,N_27759);
and UO_1479 (O_1479,N_28044,N_28599);
nor UO_1480 (O_1480,N_29978,N_28447);
and UO_1481 (O_1481,N_27838,N_29675);
nand UO_1482 (O_1482,N_29051,N_28303);
or UO_1483 (O_1483,N_28457,N_29440);
or UO_1484 (O_1484,N_27662,N_27093);
xnor UO_1485 (O_1485,N_29739,N_29571);
or UO_1486 (O_1486,N_27175,N_28034);
nor UO_1487 (O_1487,N_27012,N_27202);
or UO_1488 (O_1488,N_28607,N_29416);
and UO_1489 (O_1489,N_29569,N_27058);
nor UO_1490 (O_1490,N_28705,N_28187);
nor UO_1491 (O_1491,N_29029,N_29603);
nor UO_1492 (O_1492,N_28197,N_28084);
nand UO_1493 (O_1493,N_28702,N_27197);
xnor UO_1494 (O_1494,N_28049,N_29413);
nor UO_1495 (O_1495,N_27575,N_28508);
and UO_1496 (O_1496,N_28262,N_29952);
and UO_1497 (O_1497,N_28624,N_28403);
nor UO_1498 (O_1498,N_29565,N_29655);
or UO_1499 (O_1499,N_29057,N_27218);
xnor UO_1500 (O_1500,N_29514,N_28233);
and UO_1501 (O_1501,N_27469,N_28732);
and UO_1502 (O_1502,N_28616,N_29889);
and UO_1503 (O_1503,N_28186,N_27516);
and UO_1504 (O_1504,N_28019,N_28815);
nor UO_1505 (O_1505,N_29565,N_29335);
and UO_1506 (O_1506,N_29618,N_28230);
and UO_1507 (O_1507,N_27542,N_28697);
or UO_1508 (O_1508,N_27596,N_29554);
nor UO_1509 (O_1509,N_28917,N_29710);
nand UO_1510 (O_1510,N_29194,N_27561);
or UO_1511 (O_1511,N_27357,N_27542);
or UO_1512 (O_1512,N_29477,N_29272);
nand UO_1513 (O_1513,N_28617,N_28879);
and UO_1514 (O_1514,N_29449,N_29193);
xor UO_1515 (O_1515,N_27734,N_27934);
and UO_1516 (O_1516,N_28184,N_28227);
or UO_1517 (O_1517,N_28524,N_27875);
or UO_1518 (O_1518,N_29693,N_27791);
nor UO_1519 (O_1519,N_27300,N_27196);
or UO_1520 (O_1520,N_28759,N_28341);
or UO_1521 (O_1521,N_28373,N_27767);
or UO_1522 (O_1522,N_27452,N_27659);
nand UO_1523 (O_1523,N_27925,N_28776);
or UO_1524 (O_1524,N_28735,N_28857);
nor UO_1525 (O_1525,N_29160,N_28433);
or UO_1526 (O_1526,N_28140,N_27061);
nor UO_1527 (O_1527,N_28144,N_27749);
xor UO_1528 (O_1528,N_28523,N_28863);
nor UO_1529 (O_1529,N_28106,N_29934);
xor UO_1530 (O_1530,N_28942,N_28938);
nand UO_1531 (O_1531,N_29088,N_28145);
nor UO_1532 (O_1532,N_29631,N_28719);
and UO_1533 (O_1533,N_27815,N_27179);
and UO_1534 (O_1534,N_27931,N_28587);
nor UO_1535 (O_1535,N_27199,N_27706);
nor UO_1536 (O_1536,N_28669,N_29372);
or UO_1537 (O_1537,N_29277,N_29805);
or UO_1538 (O_1538,N_27382,N_27225);
xnor UO_1539 (O_1539,N_27856,N_27065);
and UO_1540 (O_1540,N_29476,N_29032);
nand UO_1541 (O_1541,N_27185,N_29498);
and UO_1542 (O_1542,N_28800,N_29047);
nand UO_1543 (O_1543,N_27631,N_27322);
nor UO_1544 (O_1544,N_28023,N_27857);
nand UO_1545 (O_1545,N_28603,N_29769);
and UO_1546 (O_1546,N_29452,N_29924);
or UO_1547 (O_1547,N_28680,N_29255);
and UO_1548 (O_1548,N_29446,N_28217);
nor UO_1549 (O_1549,N_27913,N_27745);
nand UO_1550 (O_1550,N_27846,N_28013);
xor UO_1551 (O_1551,N_29073,N_28346);
or UO_1552 (O_1552,N_27592,N_29334);
xnor UO_1553 (O_1553,N_27529,N_27508);
xor UO_1554 (O_1554,N_27107,N_28394);
nor UO_1555 (O_1555,N_29914,N_28497);
nand UO_1556 (O_1556,N_28256,N_27858);
nor UO_1557 (O_1557,N_29024,N_27930);
nand UO_1558 (O_1558,N_28420,N_27959);
nand UO_1559 (O_1559,N_29366,N_27393);
or UO_1560 (O_1560,N_29151,N_29384);
nand UO_1561 (O_1561,N_28866,N_29367);
and UO_1562 (O_1562,N_29735,N_28494);
nor UO_1563 (O_1563,N_27365,N_29680);
and UO_1564 (O_1564,N_27110,N_28507);
or UO_1565 (O_1565,N_29293,N_29308);
nor UO_1566 (O_1566,N_27722,N_27681);
or UO_1567 (O_1567,N_28923,N_28598);
or UO_1568 (O_1568,N_27945,N_27896);
and UO_1569 (O_1569,N_29206,N_29642);
nor UO_1570 (O_1570,N_28231,N_29601);
or UO_1571 (O_1571,N_29776,N_29857);
or UO_1572 (O_1572,N_27103,N_27821);
or UO_1573 (O_1573,N_29953,N_27748);
or UO_1574 (O_1574,N_29861,N_28829);
nor UO_1575 (O_1575,N_29354,N_28019);
nor UO_1576 (O_1576,N_27502,N_29179);
nor UO_1577 (O_1577,N_28172,N_28250);
nand UO_1578 (O_1578,N_27598,N_29404);
xnor UO_1579 (O_1579,N_29529,N_29995);
or UO_1580 (O_1580,N_27463,N_28723);
nor UO_1581 (O_1581,N_28489,N_28096);
nor UO_1582 (O_1582,N_27241,N_28792);
nor UO_1583 (O_1583,N_29589,N_29394);
nand UO_1584 (O_1584,N_28584,N_29441);
nor UO_1585 (O_1585,N_29986,N_27660);
nor UO_1586 (O_1586,N_27906,N_27698);
or UO_1587 (O_1587,N_27342,N_27703);
xor UO_1588 (O_1588,N_28410,N_28734);
or UO_1589 (O_1589,N_28462,N_29505);
nand UO_1590 (O_1590,N_27264,N_28331);
xnor UO_1591 (O_1591,N_28934,N_29330);
xnor UO_1592 (O_1592,N_29370,N_27951);
and UO_1593 (O_1593,N_28773,N_28919);
xnor UO_1594 (O_1594,N_27811,N_27522);
xnor UO_1595 (O_1595,N_28223,N_28740);
or UO_1596 (O_1596,N_29436,N_29265);
xor UO_1597 (O_1597,N_27928,N_27149);
and UO_1598 (O_1598,N_28132,N_27824);
nor UO_1599 (O_1599,N_29065,N_27540);
or UO_1600 (O_1600,N_28606,N_29923);
or UO_1601 (O_1601,N_28183,N_27309);
or UO_1602 (O_1602,N_27114,N_28033);
nand UO_1603 (O_1603,N_28401,N_29563);
or UO_1604 (O_1604,N_28521,N_28186);
nand UO_1605 (O_1605,N_29030,N_27750);
xnor UO_1606 (O_1606,N_28282,N_28311);
and UO_1607 (O_1607,N_27889,N_29595);
or UO_1608 (O_1608,N_29967,N_29750);
and UO_1609 (O_1609,N_28541,N_27902);
and UO_1610 (O_1610,N_28807,N_29640);
or UO_1611 (O_1611,N_29073,N_27464);
and UO_1612 (O_1612,N_28433,N_28755);
nand UO_1613 (O_1613,N_27499,N_29462);
and UO_1614 (O_1614,N_28145,N_28603);
xor UO_1615 (O_1615,N_28741,N_29988);
or UO_1616 (O_1616,N_29048,N_27354);
nand UO_1617 (O_1617,N_27117,N_29818);
xor UO_1618 (O_1618,N_28934,N_27759);
and UO_1619 (O_1619,N_28476,N_29998);
xor UO_1620 (O_1620,N_29424,N_29345);
xnor UO_1621 (O_1621,N_27526,N_27731);
or UO_1622 (O_1622,N_27556,N_28613);
and UO_1623 (O_1623,N_27149,N_29954);
nor UO_1624 (O_1624,N_28225,N_28724);
xor UO_1625 (O_1625,N_27597,N_27790);
or UO_1626 (O_1626,N_28542,N_29436);
nand UO_1627 (O_1627,N_28780,N_28439);
or UO_1628 (O_1628,N_29493,N_28246);
or UO_1629 (O_1629,N_27489,N_27493);
nand UO_1630 (O_1630,N_27786,N_29730);
nor UO_1631 (O_1631,N_29631,N_27175);
nand UO_1632 (O_1632,N_29698,N_27219);
or UO_1633 (O_1633,N_27092,N_27040);
or UO_1634 (O_1634,N_29906,N_27192);
and UO_1635 (O_1635,N_27896,N_29424);
xnor UO_1636 (O_1636,N_29510,N_27353);
or UO_1637 (O_1637,N_27985,N_28413);
xor UO_1638 (O_1638,N_27376,N_29033);
nand UO_1639 (O_1639,N_29112,N_29381);
nor UO_1640 (O_1640,N_29716,N_28483);
or UO_1641 (O_1641,N_27416,N_29330);
nand UO_1642 (O_1642,N_27561,N_27592);
xnor UO_1643 (O_1643,N_28426,N_27804);
nor UO_1644 (O_1644,N_27006,N_27011);
and UO_1645 (O_1645,N_29101,N_27351);
or UO_1646 (O_1646,N_28900,N_27937);
nand UO_1647 (O_1647,N_27069,N_29670);
nand UO_1648 (O_1648,N_29382,N_27816);
nor UO_1649 (O_1649,N_29267,N_29383);
nor UO_1650 (O_1650,N_29295,N_28537);
and UO_1651 (O_1651,N_28800,N_29285);
and UO_1652 (O_1652,N_27400,N_28476);
xnor UO_1653 (O_1653,N_28800,N_27064);
or UO_1654 (O_1654,N_27213,N_27948);
and UO_1655 (O_1655,N_27520,N_28938);
nor UO_1656 (O_1656,N_28552,N_29147);
and UO_1657 (O_1657,N_29613,N_28020);
xnor UO_1658 (O_1658,N_28135,N_29813);
nand UO_1659 (O_1659,N_27485,N_27552);
xnor UO_1660 (O_1660,N_29214,N_28255);
or UO_1661 (O_1661,N_29452,N_28618);
and UO_1662 (O_1662,N_27256,N_28143);
or UO_1663 (O_1663,N_28081,N_27000);
xnor UO_1664 (O_1664,N_27666,N_29912);
nand UO_1665 (O_1665,N_29119,N_27434);
xor UO_1666 (O_1666,N_28825,N_28750);
nand UO_1667 (O_1667,N_28438,N_27024);
xor UO_1668 (O_1668,N_29450,N_28710);
and UO_1669 (O_1669,N_27311,N_27920);
or UO_1670 (O_1670,N_28773,N_29508);
and UO_1671 (O_1671,N_28337,N_29414);
xnor UO_1672 (O_1672,N_29331,N_28543);
nand UO_1673 (O_1673,N_28018,N_27675);
nor UO_1674 (O_1674,N_28830,N_28180);
nor UO_1675 (O_1675,N_29586,N_29758);
and UO_1676 (O_1676,N_28054,N_29914);
nor UO_1677 (O_1677,N_28924,N_27884);
or UO_1678 (O_1678,N_28692,N_29860);
or UO_1679 (O_1679,N_27073,N_28915);
nor UO_1680 (O_1680,N_27095,N_28655);
xor UO_1681 (O_1681,N_27238,N_27892);
nor UO_1682 (O_1682,N_28522,N_29203);
nor UO_1683 (O_1683,N_27798,N_29950);
or UO_1684 (O_1684,N_27048,N_29538);
nor UO_1685 (O_1685,N_29452,N_28487);
nor UO_1686 (O_1686,N_27078,N_27043);
or UO_1687 (O_1687,N_27379,N_29467);
nand UO_1688 (O_1688,N_27996,N_28594);
nand UO_1689 (O_1689,N_29721,N_27295);
nor UO_1690 (O_1690,N_29343,N_29941);
nand UO_1691 (O_1691,N_27273,N_27234);
and UO_1692 (O_1692,N_29240,N_27019);
or UO_1693 (O_1693,N_27411,N_27180);
nor UO_1694 (O_1694,N_29197,N_29148);
xor UO_1695 (O_1695,N_27453,N_27752);
or UO_1696 (O_1696,N_28089,N_27215);
xor UO_1697 (O_1697,N_28165,N_29195);
or UO_1698 (O_1698,N_28280,N_28427);
nand UO_1699 (O_1699,N_28436,N_29236);
or UO_1700 (O_1700,N_29904,N_28664);
or UO_1701 (O_1701,N_28814,N_29964);
and UO_1702 (O_1702,N_29883,N_27258);
xor UO_1703 (O_1703,N_28552,N_27329);
or UO_1704 (O_1704,N_28319,N_28609);
nand UO_1705 (O_1705,N_28879,N_28813);
nand UO_1706 (O_1706,N_29067,N_27956);
and UO_1707 (O_1707,N_28681,N_28293);
and UO_1708 (O_1708,N_28139,N_28105);
xnor UO_1709 (O_1709,N_28852,N_27768);
or UO_1710 (O_1710,N_29776,N_29261);
or UO_1711 (O_1711,N_27069,N_27200);
and UO_1712 (O_1712,N_29940,N_29385);
nand UO_1713 (O_1713,N_29340,N_28538);
or UO_1714 (O_1714,N_28812,N_29091);
or UO_1715 (O_1715,N_28019,N_28632);
nand UO_1716 (O_1716,N_27053,N_28087);
and UO_1717 (O_1717,N_27128,N_29561);
nor UO_1718 (O_1718,N_27677,N_29894);
nand UO_1719 (O_1719,N_29616,N_28944);
nand UO_1720 (O_1720,N_28341,N_27724);
nor UO_1721 (O_1721,N_29267,N_27868);
and UO_1722 (O_1722,N_28024,N_27687);
xnor UO_1723 (O_1723,N_28942,N_29571);
xor UO_1724 (O_1724,N_28847,N_28962);
xor UO_1725 (O_1725,N_29338,N_28999);
and UO_1726 (O_1726,N_27371,N_27474);
xor UO_1727 (O_1727,N_28767,N_29357);
and UO_1728 (O_1728,N_28535,N_27774);
xnor UO_1729 (O_1729,N_28148,N_29739);
xnor UO_1730 (O_1730,N_27000,N_28697);
and UO_1731 (O_1731,N_28678,N_29806);
xnor UO_1732 (O_1732,N_28115,N_27265);
xnor UO_1733 (O_1733,N_27581,N_29067);
nor UO_1734 (O_1734,N_29149,N_28725);
nor UO_1735 (O_1735,N_29468,N_28967);
xnor UO_1736 (O_1736,N_29313,N_27748);
xor UO_1737 (O_1737,N_27927,N_29396);
nor UO_1738 (O_1738,N_27748,N_28701);
or UO_1739 (O_1739,N_27587,N_29375);
and UO_1740 (O_1740,N_29452,N_28149);
xnor UO_1741 (O_1741,N_29546,N_28856);
nor UO_1742 (O_1742,N_29552,N_27208);
nor UO_1743 (O_1743,N_27265,N_29043);
nor UO_1744 (O_1744,N_29143,N_27913);
nand UO_1745 (O_1745,N_28008,N_28773);
or UO_1746 (O_1746,N_29933,N_27562);
or UO_1747 (O_1747,N_29221,N_28521);
xnor UO_1748 (O_1748,N_29670,N_29840);
nand UO_1749 (O_1749,N_28693,N_27446);
nand UO_1750 (O_1750,N_27314,N_28555);
nand UO_1751 (O_1751,N_28023,N_29473);
and UO_1752 (O_1752,N_27564,N_28448);
or UO_1753 (O_1753,N_29166,N_29436);
and UO_1754 (O_1754,N_28537,N_28393);
nor UO_1755 (O_1755,N_29031,N_28790);
or UO_1756 (O_1756,N_29719,N_29620);
or UO_1757 (O_1757,N_28026,N_28529);
xnor UO_1758 (O_1758,N_28730,N_29201);
or UO_1759 (O_1759,N_29239,N_29812);
xor UO_1760 (O_1760,N_27716,N_29434);
nor UO_1761 (O_1761,N_27874,N_28990);
and UO_1762 (O_1762,N_28294,N_29550);
nand UO_1763 (O_1763,N_27300,N_27380);
or UO_1764 (O_1764,N_28886,N_29682);
nor UO_1765 (O_1765,N_29835,N_28572);
or UO_1766 (O_1766,N_29091,N_29698);
xor UO_1767 (O_1767,N_27869,N_28281);
nor UO_1768 (O_1768,N_29535,N_27041);
or UO_1769 (O_1769,N_27409,N_27033);
and UO_1770 (O_1770,N_28603,N_27978);
nor UO_1771 (O_1771,N_29808,N_27200);
and UO_1772 (O_1772,N_29901,N_29599);
and UO_1773 (O_1773,N_28674,N_29999);
xnor UO_1774 (O_1774,N_29740,N_28580);
xor UO_1775 (O_1775,N_28537,N_28332);
or UO_1776 (O_1776,N_28756,N_27752);
xnor UO_1777 (O_1777,N_29127,N_29200);
and UO_1778 (O_1778,N_29433,N_29884);
or UO_1779 (O_1779,N_29402,N_27248);
nand UO_1780 (O_1780,N_28590,N_29243);
nand UO_1781 (O_1781,N_27871,N_29792);
xor UO_1782 (O_1782,N_29818,N_27787);
and UO_1783 (O_1783,N_27807,N_29598);
and UO_1784 (O_1784,N_28993,N_29509);
xor UO_1785 (O_1785,N_29024,N_28489);
or UO_1786 (O_1786,N_29417,N_28963);
xor UO_1787 (O_1787,N_29907,N_27321);
xor UO_1788 (O_1788,N_29749,N_28113);
and UO_1789 (O_1789,N_29383,N_27176);
xor UO_1790 (O_1790,N_27468,N_27828);
xor UO_1791 (O_1791,N_27045,N_29906);
or UO_1792 (O_1792,N_28439,N_27203);
nor UO_1793 (O_1793,N_28131,N_27283);
nor UO_1794 (O_1794,N_29736,N_27698);
or UO_1795 (O_1795,N_29118,N_27910);
or UO_1796 (O_1796,N_29525,N_29717);
nand UO_1797 (O_1797,N_29247,N_27529);
and UO_1798 (O_1798,N_28038,N_27616);
nor UO_1799 (O_1799,N_28659,N_29322);
or UO_1800 (O_1800,N_27583,N_29582);
and UO_1801 (O_1801,N_27935,N_27247);
or UO_1802 (O_1802,N_29370,N_28212);
nor UO_1803 (O_1803,N_27235,N_27584);
xnor UO_1804 (O_1804,N_28054,N_28394);
nor UO_1805 (O_1805,N_27367,N_29813);
nand UO_1806 (O_1806,N_27352,N_27533);
xnor UO_1807 (O_1807,N_29527,N_28426);
and UO_1808 (O_1808,N_28219,N_28252);
nor UO_1809 (O_1809,N_28458,N_29317);
or UO_1810 (O_1810,N_29893,N_28238);
nand UO_1811 (O_1811,N_28845,N_27259);
and UO_1812 (O_1812,N_29103,N_29521);
nor UO_1813 (O_1813,N_28819,N_28973);
xor UO_1814 (O_1814,N_27950,N_28383);
and UO_1815 (O_1815,N_29311,N_27000);
and UO_1816 (O_1816,N_28271,N_29050);
or UO_1817 (O_1817,N_27054,N_27630);
or UO_1818 (O_1818,N_29815,N_27192);
xor UO_1819 (O_1819,N_28607,N_28432);
nand UO_1820 (O_1820,N_28379,N_29504);
nand UO_1821 (O_1821,N_27901,N_27194);
nand UO_1822 (O_1822,N_28409,N_29288);
xnor UO_1823 (O_1823,N_27528,N_29540);
or UO_1824 (O_1824,N_29810,N_29353);
nor UO_1825 (O_1825,N_29067,N_27146);
or UO_1826 (O_1826,N_29628,N_29196);
nand UO_1827 (O_1827,N_27284,N_28643);
nor UO_1828 (O_1828,N_27314,N_27923);
and UO_1829 (O_1829,N_29572,N_28673);
nor UO_1830 (O_1830,N_27564,N_29492);
xnor UO_1831 (O_1831,N_29059,N_28669);
or UO_1832 (O_1832,N_27500,N_29037);
nor UO_1833 (O_1833,N_29441,N_29410);
xor UO_1834 (O_1834,N_27290,N_28640);
nor UO_1835 (O_1835,N_27492,N_29649);
xnor UO_1836 (O_1836,N_29498,N_27774);
xor UO_1837 (O_1837,N_28952,N_28645);
nand UO_1838 (O_1838,N_28574,N_27186);
or UO_1839 (O_1839,N_27823,N_28945);
xnor UO_1840 (O_1840,N_28486,N_29710);
nand UO_1841 (O_1841,N_27013,N_27101);
and UO_1842 (O_1842,N_28498,N_29017);
xnor UO_1843 (O_1843,N_27253,N_27798);
and UO_1844 (O_1844,N_29083,N_28166);
and UO_1845 (O_1845,N_27203,N_27236);
xor UO_1846 (O_1846,N_28643,N_28192);
nand UO_1847 (O_1847,N_29237,N_29812);
xnor UO_1848 (O_1848,N_27528,N_27992);
and UO_1849 (O_1849,N_28712,N_27363);
xnor UO_1850 (O_1850,N_27739,N_29789);
nand UO_1851 (O_1851,N_28873,N_29978);
xnor UO_1852 (O_1852,N_28722,N_28254);
nand UO_1853 (O_1853,N_27911,N_29590);
and UO_1854 (O_1854,N_27648,N_27611);
nand UO_1855 (O_1855,N_29277,N_28687);
nor UO_1856 (O_1856,N_28377,N_29157);
or UO_1857 (O_1857,N_28252,N_27255);
and UO_1858 (O_1858,N_27903,N_27824);
xnor UO_1859 (O_1859,N_29699,N_28356);
nor UO_1860 (O_1860,N_29287,N_28196);
nor UO_1861 (O_1861,N_27128,N_27648);
xnor UO_1862 (O_1862,N_29480,N_29847);
nor UO_1863 (O_1863,N_28669,N_27655);
and UO_1864 (O_1864,N_27831,N_29041);
xnor UO_1865 (O_1865,N_29042,N_29484);
or UO_1866 (O_1866,N_28871,N_28138);
xnor UO_1867 (O_1867,N_28535,N_28678);
and UO_1868 (O_1868,N_28323,N_29457);
nor UO_1869 (O_1869,N_27964,N_28222);
or UO_1870 (O_1870,N_28422,N_27091);
nand UO_1871 (O_1871,N_27205,N_28307);
nand UO_1872 (O_1872,N_29430,N_27310);
and UO_1873 (O_1873,N_29692,N_29003);
and UO_1874 (O_1874,N_29352,N_28127);
xnor UO_1875 (O_1875,N_27284,N_28314);
xnor UO_1876 (O_1876,N_27594,N_28691);
or UO_1877 (O_1877,N_28854,N_29196);
and UO_1878 (O_1878,N_28514,N_27785);
xor UO_1879 (O_1879,N_28723,N_28485);
or UO_1880 (O_1880,N_28009,N_28401);
nand UO_1881 (O_1881,N_29052,N_29810);
nor UO_1882 (O_1882,N_29149,N_29218);
xnor UO_1883 (O_1883,N_28281,N_27180);
nand UO_1884 (O_1884,N_29123,N_27218);
or UO_1885 (O_1885,N_27264,N_28148);
xnor UO_1886 (O_1886,N_27949,N_28467);
and UO_1887 (O_1887,N_29236,N_28441);
nand UO_1888 (O_1888,N_28583,N_29977);
or UO_1889 (O_1889,N_28819,N_28647);
nand UO_1890 (O_1890,N_27986,N_28313);
nand UO_1891 (O_1891,N_27942,N_28944);
and UO_1892 (O_1892,N_27823,N_28211);
nor UO_1893 (O_1893,N_29559,N_29655);
nand UO_1894 (O_1894,N_28173,N_27019);
nand UO_1895 (O_1895,N_29672,N_27675);
nand UO_1896 (O_1896,N_28235,N_29789);
nand UO_1897 (O_1897,N_27017,N_28177);
xor UO_1898 (O_1898,N_29067,N_28465);
and UO_1899 (O_1899,N_27247,N_27774);
and UO_1900 (O_1900,N_29741,N_28954);
xnor UO_1901 (O_1901,N_29017,N_28708);
and UO_1902 (O_1902,N_27944,N_28241);
nand UO_1903 (O_1903,N_28044,N_28916);
xor UO_1904 (O_1904,N_28230,N_27589);
xor UO_1905 (O_1905,N_29317,N_28254);
nor UO_1906 (O_1906,N_27430,N_27733);
nor UO_1907 (O_1907,N_27687,N_28039);
or UO_1908 (O_1908,N_27914,N_27052);
nand UO_1909 (O_1909,N_29816,N_28706);
nor UO_1910 (O_1910,N_27567,N_29129);
or UO_1911 (O_1911,N_27657,N_27081);
and UO_1912 (O_1912,N_27235,N_29905);
or UO_1913 (O_1913,N_28236,N_29970);
or UO_1914 (O_1914,N_29679,N_28347);
xor UO_1915 (O_1915,N_28355,N_29654);
nor UO_1916 (O_1916,N_28090,N_29778);
and UO_1917 (O_1917,N_28268,N_27809);
nor UO_1918 (O_1918,N_27574,N_28120);
nor UO_1919 (O_1919,N_29735,N_27814);
or UO_1920 (O_1920,N_27590,N_29647);
xor UO_1921 (O_1921,N_28428,N_29700);
xnor UO_1922 (O_1922,N_27958,N_27703);
nor UO_1923 (O_1923,N_28711,N_28352);
and UO_1924 (O_1924,N_28982,N_28077);
nand UO_1925 (O_1925,N_28280,N_29061);
xnor UO_1926 (O_1926,N_27526,N_28612);
nand UO_1927 (O_1927,N_28629,N_29716);
xnor UO_1928 (O_1928,N_29202,N_29609);
xnor UO_1929 (O_1929,N_27522,N_27325);
and UO_1930 (O_1930,N_28570,N_29903);
nor UO_1931 (O_1931,N_28612,N_27888);
and UO_1932 (O_1932,N_28932,N_28323);
nand UO_1933 (O_1933,N_28639,N_28562);
and UO_1934 (O_1934,N_28486,N_29583);
nor UO_1935 (O_1935,N_29909,N_29862);
nand UO_1936 (O_1936,N_27832,N_28873);
xnor UO_1937 (O_1937,N_27341,N_28934);
and UO_1938 (O_1938,N_28764,N_27317);
nand UO_1939 (O_1939,N_29665,N_29802);
nand UO_1940 (O_1940,N_28034,N_27638);
xor UO_1941 (O_1941,N_27819,N_28657);
nand UO_1942 (O_1942,N_27661,N_29369);
and UO_1943 (O_1943,N_29691,N_27376);
nor UO_1944 (O_1944,N_29967,N_29116);
nand UO_1945 (O_1945,N_29716,N_27892);
and UO_1946 (O_1946,N_29960,N_29174);
nor UO_1947 (O_1947,N_28413,N_28277);
nand UO_1948 (O_1948,N_28203,N_27203);
and UO_1949 (O_1949,N_29125,N_27376);
nor UO_1950 (O_1950,N_29242,N_27642);
and UO_1951 (O_1951,N_29712,N_28090);
and UO_1952 (O_1952,N_28147,N_29251);
nand UO_1953 (O_1953,N_27720,N_27678);
or UO_1954 (O_1954,N_28440,N_27664);
nand UO_1955 (O_1955,N_28034,N_29756);
or UO_1956 (O_1956,N_28516,N_29106);
xnor UO_1957 (O_1957,N_29619,N_27987);
nand UO_1958 (O_1958,N_28992,N_27558);
nand UO_1959 (O_1959,N_28649,N_27091);
nand UO_1960 (O_1960,N_28417,N_28250);
nand UO_1961 (O_1961,N_29929,N_27588);
xor UO_1962 (O_1962,N_29211,N_27371);
xor UO_1963 (O_1963,N_28109,N_28614);
nor UO_1964 (O_1964,N_27731,N_29267);
nor UO_1965 (O_1965,N_29576,N_29189);
and UO_1966 (O_1966,N_28025,N_27576);
and UO_1967 (O_1967,N_28976,N_29509);
and UO_1968 (O_1968,N_27227,N_27524);
xor UO_1969 (O_1969,N_27986,N_29271);
or UO_1970 (O_1970,N_28873,N_28785);
and UO_1971 (O_1971,N_28087,N_28606);
nand UO_1972 (O_1972,N_27115,N_27383);
nand UO_1973 (O_1973,N_28160,N_29256);
and UO_1974 (O_1974,N_28470,N_29043);
xnor UO_1975 (O_1975,N_29648,N_29906);
nand UO_1976 (O_1976,N_28999,N_29516);
and UO_1977 (O_1977,N_29439,N_28748);
nand UO_1978 (O_1978,N_29819,N_29369);
xnor UO_1979 (O_1979,N_28456,N_29890);
or UO_1980 (O_1980,N_27618,N_29361);
nand UO_1981 (O_1981,N_29651,N_27476);
and UO_1982 (O_1982,N_27639,N_27152);
nor UO_1983 (O_1983,N_29848,N_27458);
nor UO_1984 (O_1984,N_27106,N_28862);
and UO_1985 (O_1985,N_29119,N_27273);
xnor UO_1986 (O_1986,N_27303,N_27361);
xnor UO_1987 (O_1987,N_29662,N_27001);
nor UO_1988 (O_1988,N_29267,N_27271);
nor UO_1989 (O_1989,N_28647,N_27545);
xnor UO_1990 (O_1990,N_28618,N_29696);
nand UO_1991 (O_1991,N_27674,N_27031);
or UO_1992 (O_1992,N_27926,N_28449);
and UO_1993 (O_1993,N_28465,N_29824);
nand UO_1994 (O_1994,N_28168,N_29884);
nor UO_1995 (O_1995,N_27848,N_27923);
xnor UO_1996 (O_1996,N_27228,N_27163);
and UO_1997 (O_1997,N_27662,N_27364);
or UO_1998 (O_1998,N_29862,N_29172);
and UO_1999 (O_1999,N_28067,N_27393);
nor UO_2000 (O_2000,N_27973,N_29827);
nor UO_2001 (O_2001,N_27735,N_27499);
nand UO_2002 (O_2002,N_29304,N_29423);
nand UO_2003 (O_2003,N_27873,N_28567);
nor UO_2004 (O_2004,N_29148,N_29600);
nor UO_2005 (O_2005,N_29980,N_27005);
and UO_2006 (O_2006,N_27908,N_29161);
and UO_2007 (O_2007,N_28793,N_29112);
or UO_2008 (O_2008,N_27798,N_27508);
nor UO_2009 (O_2009,N_27919,N_27897);
and UO_2010 (O_2010,N_27506,N_29893);
nand UO_2011 (O_2011,N_29085,N_28008);
nor UO_2012 (O_2012,N_28784,N_29280);
nand UO_2013 (O_2013,N_29109,N_28447);
xor UO_2014 (O_2014,N_28450,N_27151);
and UO_2015 (O_2015,N_29611,N_28021);
or UO_2016 (O_2016,N_29912,N_29936);
nand UO_2017 (O_2017,N_27959,N_29929);
xor UO_2018 (O_2018,N_29307,N_28687);
nor UO_2019 (O_2019,N_28310,N_29089);
or UO_2020 (O_2020,N_28371,N_27013);
and UO_2021 (O_2021,N_28231,N_27484);
nand UO_2022 (O_2022,N_29617,N_27208);
xnor UO_2023 (O_2023,N_29563,N_27055);
nand UO_2024 (O_2024,N_28857,N_28475);
and UO_2025 (O_2025,N_29252,N_28694);
and UO_2026 (O_2026,N_27163,N_29044);
nor UO_2027 (O_2027,N_27319,N_29647);
nor UO_2028 (O_2028,N_28697,N_29008);
xnor UO_2029 (O_2029,N_28418,N_27534);
and UO_2030 (O_2030,N_28760,N_28533);
nor UO_2031 (O_2031,N_28560,N_27982);
xor UO_2032 (O_2032,N_27427,N_29378);
nand UO_2033 (O_2033,N_27167,N_28154);
xor UO_2034 (O_2034,N_28002,N_27674);
nor UO_2035 (O_2035,N_27447,N_28895);
xor UO_2036 (O_2036,N_27193,N_29239);
nand UO_2037 (O_2037,N_29253,N_28660);
xor UO_2038 (O_2038,N_28561,N_28317);
nand UO_2039 (O_2039,N_27256,N_29967);
xnor UO_2040 (O_2040,N_27274,N_29101);
or UO_2041 (O_2041,N_27653,N_28616);
or UO_2042 (O_2042,N_27307,N_29765);
nand UO_2043 (O_2043,N_27305,N_28500);
nand UO_2044 (O_2044,N_28301,N_29740);
xor UO_2045 (O_2045,N_28922,N_28050);
xnor UO_2046 (O_2046,N_27643,N_27135);
or UO_2047 (O_2047,N_27733,N_27183);
xnor UO_2048 (O_2048,N_27901,N_28946);
xnor UO_2049 (O_2049,N_29794,N_29357);
xor UO_2050 (O_2050,N_28425,N_29276);
and UO_2051 (O_2051,N_27318,N_29195);
or UO_2052 (O_2052,N_29303,N_27348);
and UO_2053 (O_2053,N_29736,N_28744);
or UO_2054 (O_2054,N_27662,N_28334);
xnor UO_2055 (O_2055,N_29447,N_29880);
and UO_2056 (O_2056,N_27678,N_27893);
and UO_2057 (O_2057,N_28696,N_27231);
or UO_2058 (O_2058,N_28049,N_27796);
nor UO_2059 (O_2059,N_28659,N_28143);
or UO_2060 (O_2060,N_29759,N_29853);
or UO_2061 (O_2061,N_28266,N_28215);
or UO_2062 (O_2062,N_28495,N_28548);
and UO_2063 (O_2063,N_29351,N_29598);
xnor UO_2064 (O_2064,N_29645,N_28766);
or UO_2065 (O_2065,N_27258,N_27893);
and UO_2066 (O_2066,N_28187,N_28428);
nor UO_2067 (O_2067,N_27380,N_28075);
and UO_2068 (O_2068,N_27097,N_29891);
or UO_2069 (O_2069,N_28263,N_28034);
nor UO_2070 (O_2070,N_27571,N_29432);
xor UO_2071 (O_2071,N_27329,N_29327);
and UO_2072 (O_2072,N_29155,N_29506);
nor UO_2073 (O_2073,N_28789,N_28950);
xnor UO_2074 (O_2074,N_29001,N_27351);
xor UO_2075 (O_2075,N_28121,N_28950);
nand UO_2076 (O_2076,N_28440,N_28074);
and UO_2077 (O_2077,N_29744,N_27911);
and UO_2078 (O_2078,N_28576,N_28717);
or UO_2079 (O_2079,N_27714,N_28283);
nand UO_2080 (O_2080,N_27204,N_28958);
or UO_2081 (O_2081,N_27947,N_29242);
or UO_2082 (O_2082,N_28226,N_27892);
or UO_2083 (O_2083,N_28527,N_27531);
and UO_2084 (O_2084,N_27186,N_27753);
nand UO_2085 (O_2085,N_29466,N_27340);
or UO_2086 (O_2086,N_29404,N_28558);
nand UO_2087 (O_2087,N_29884,N_29197);
nand UO_2088 (O_2088,N_28147,N_29494);
nor UO_2089 (O_2089,N_29647,N_28758);
nand UO_2090 (O_2090,N_29408,N_27114);
nand UO_2091 (O_2091,N_27411,N_28681);
nor UO_2092 (O_2092,N_27417,N_29410);
nor UO_2093 (O_2093,N_28882,N_29921);
xnor UO_2094 (O_2094,N_27007,N_29551);
nand UO_2095 (O_2095,N_28215,N_29128);
nand UO_2096 (O_2096,N_29537,N_28752);
xor UO_2097 (O_2097,N_28172,N_29919);
nor UO_2098 (O_2098,N_28447,N_29772);
nor UO_2099 (O_2099,N_27376,N_28458);
xnor UO_2100 (O_2100,N_28201,N_28992);
or UO_2101 (O_2101,N_29018,N_29863);
or UO_2102 (O_2102,N_29831,N_29153);
nor UO_2103 (O_2103,N_29019,N_27176);
xor UO_2104 (O_2104,N_29858,N_29832);
and UO_2105 (O_2105,N_28004,N_28526);
xor UO_2106 (O_2106,N_27261,N_29822);
or UO_2107 (O_2107,N_28893,N_29282);
or UO_2108 (O_2108,N_28428,N_28350);
and UO_2109 (O_2109,N_27973,N_28504);
nor UO_2110 (O_2110,N_27746,N_27204);
nor UO_2111 (O_2111,N_27925,N_28977);
nand UO_2112 (O_2112,N_27811,N_27912);
or UO_2113 (O_2113,N_28378,N_27158);
xor UO_2114 (O_2114,N_28733,N_29036);
and UO_2115 (O_2115,N_29133,N_27053);
xnor UO_2116 (O_2116,N_27915,N_28528);
or UO_2117 (O_2117,N_29119,N_29425);
or UO_2118 (O_2118,N_27624,N_28974);
nor UO_2119 (O_2119,N_28394,N_27063);
nor UO_2120 (O_2120,N_29928,N_27289);
nor UO_2121 (O_2121,N_27223,N_27853);
and UO_2122 (O_2122,N_28011,N_29901);
nor UO_2123 (O_2123,N_28520,N_28847);
or UO_2124 (O_2124,N_29831,N_27321);
nor UO_2125 (O_2125,N_27009,N_28453);
xnor UO_2126 (O_2126,N_27168,N_29330);
nor UO_2127 (O_2127,N_28103,N_27055);
or UO_2128 (O_2128,N_28095,N_28888);
or UO_2129 (O_2129,N_28122,N_28484);
and UO_2130 (O_2130,N_28683,N_27639);
nor UO_2131 (O_2131,N_28871,N_29764);
xor UO_2132 (O_2132,N_27407,N_29566);
nor UO_2133 (O_2133,N_29946,N_29968);
or UO_2134 (O_2134,N_29042,N_27087);
nand UO_2135 (O_2135,N_29728,N_27027);
nand UO_2136 (O_2136,N_29960,N_27815);
nor UO_2137 (O_2137,N_29072,N_27389);
or UO_2138 (O_2138,N_29658,N_27906);
or UO_2139 (O_2139,N_28957,N_27813);
nor UO_2140 (O_2140,N_29731,N_29250);
nor UO_2141 (O_2141,N_27862,N_29858);
nand UO_2142 (O_2142,N_28093,N_27741);
nor UO_2143 (O_2143,N_28282,N_28765);
nand UO_2144 (O_2144,N_28056,N_27917);
nand UO_2145 (O_2145,N_29998,N_28202);
and UO_2146 (O_2146,N_28933,N_29533);
nand UO_2147 (O_2147,N_29412,N_28239);
nor UO_2148 (O_2148,N_29861,N_29735);
nand UO_2149 (O_2149,N_27099,N_28843);
xor UO_2150 (O_2150,N_28500,N_29298);
xor UO_2151 (O_2151,N_29565,N_29524);
nor UO_2152 (O_2152,N_29810,N_28136);
nand UO_2153 (O_2153,N_29081,N_27069);
or UO_2154 (O_2154,N_28936,N_29407);
and UO_2155 (O_2155,N_27512,N_28714);
or UO_2156 (O_2156,N_29061,N_27218);
xor UO_2157 (O_2157,N_27767,N_28226);
xor UO_2158 (O_2158,N_27355,N_29154);
or UO_2159 (O_2159,N_29492,N_27083);
and UO_2160 (O_2160,N_27778,N_27691);
xnor UO_2161 (O_2161,N_27399,N_28876);
nand UO_2162 (O_2162,N_29201,N_29382);
or UO_2163 (O_2163,N_29493,N_29139);
nor UO_2164 (O_2164,N_27210,N_28126);
and UO_2165 (O_2165,N_29121,N_28774);
xnor UO_2166 (O_2166,N_28133,N_29349);
nand UO_2167 (O_2167,N_28320,N_28480);
nor UO_2168 (O_2168,N_29018,N_28560);
xor UO_2169 (O_2169,N_27749,N_28290);
or UO_2170 (O_2170,N_29778,N_27346);
or UO_2171 (O_2171,N_28925,N_27684);
nor UO_2172 (O_2172,N_29121,N_28915);
nand UO_2173 (O_2173,N_27865,N_29389);
xor UO_2174 (O_2174,N_28408,N_29413);
xnor UO_2175 (O_2175,N_28785,N_28110);
nor UO_2176 (O_2176,N_28866,N_29539);
nor UO_2177 (O_2177,N_28331,N_28448);
xor UO_2178 (O_2178,N_27514,N_29736);
or UO_2179 (O_2179,N_29312,N_29726);
nand UO_2180 (O_2180,N_27216,N_29184);
and UO_2181 (O_2181,N_27935,N_27310);
nor UO_2182 (O_2182,N_29472,N_27070);
xnor UO_2183 (O_2183,N_27467,N_27794);
nand UO_2184 (O_2184,N_27097,N_28138);
xnor UO_2185 (O_2185,N_28786,N_29997);
xor UO_2186 (O_2186,N_27096,N_28979);
and UO_2187 (O_2187,N_29238,N_28601);
and UO_2188 (O_2188,N_28056,N_28015);
and UO_2189 (O_2189,N_29743,N_28445);
nand UO_2190 (O_2190,N_28331,N_28549);
xnor UO_2191 (O_2191,N_27831,N_27080);
and UO_2192 (O_2192,N_27421,N_27829);
or UO_2193 (O_2193,N_29076,N_29308);
nand UO_2194 (O_2194,N_29187,N_27146);
or UO_2195 (O_2195,N_29301,N_28275);
and UO_2196 (O_2196,N_27008,N_29049);
and UO_2197 (O_2197,N_29583,N_27481);
or UO_2198 (O_2198,N_27764,N_27891);
nor UO_2199 (O_2199,N_27971,N_29033);
or UO_2200 (O_2200,N_28671,N_27050);
and UO_2201 (O_2201,N_28524,N_27668);
or UO_2202 (O_2202,N_28868,N_27091);
xor UO_2203 (O_2203,N_29520,N_28486);
nor UO_2204 (O_2204,N_27510,N_28635);
nand UO_2205 (O_2205,N_27485,N_27016);
nand UO_2206 (O_2206,N_27202,N_27019);
xor UO_2207 (O_2207,N_29439,N_28162);
xor UO_2208 (O_2208,N_27820,N_29369);
nand UO_2209 (O_2209,N_28620,N_27071);
or UO_2210 (O_2210,N_28778,N_29647);
or UO_2211 (O_2211,N_28699,N_28575);
xor UO_2212 (O_2212,N_28193,N_29781);
xor UO_2213 (O_2213,N_27214,N_28126);
or UO_2214 (O_2214,N_27668,N_27587);
or UO_2215 (O_2215,N_29431,N_29129);
and UO_2216 (O_2216,N_28776,N_29105);
nand UO_2217 (O_2217,N_27115,N_27450);
nor UO_2218 (O_2218,N_29356,N_27664);
nand UO_2219 (O_2219,N_28567,N_27276);
xnor UO_2220 (O_2220,N_29151,N_28885);
nor UO_2221 (O_2221,N_28339,N_27699);
and UO_2222 (O_2222,N_28764,N_29299);
or UO_2223 (O_2223,N_28081,N_27203);
and UO_2224 (O_2224,N_29086,N_27283);
nand UO_2225 (O_2225,N_29060,N_27316);
and UO_2226 (O_2226,N_28664,N_27469);
nand UO_2227 (O_2227,N_29647,N_29536);
nand UO_2228 (O_2228,N_27681,N_28731);
nand UO_2229 (O_2229,N_27194,N_28446);
nand UO_2230 (O_2230,N_29226,N_28516);
xnor UO_2231 (O_2231,N_29066,N_28793);
nor UO_2232 (O_2232,N_27794,N_27844);
and UO_2233 (O_2233,N_29525,N_27885);
nand UO_2234 (O_2234,N_29906,N_27495);
xnor UO_2235 (O_2235,N_27506,N_28077);
xnor UO_2236 (O_2236,N_27283,N_29652);
nor UO_2237 (O_2237,N_27181,N_27568);
and UO_2238 (O_2238,N_28627,N_29769);
or UO_2239 (O_2239,N_29382,N_27421);
or UO_2240 (O_2240,N_27896,N_27589);
and UO_2241 (O_2241,N_27523,N_27755);
xor UO_2242 (O_2242,N_29100,N_27533);
and UO_2243 (O_2243,N_27371,N_27137);
and UO_2244 (O_2244,N_28980,N_28645);
nor UO_2245 (O_2245,N_27101,N_29572);
nand UO_2246 (O_2246,N_27734,N_27554);
xor UO_2247 (O_2247,N_29451,N_27192);
and UO_2248 (O_2248,N_27058,N_29049);
and UO_2249 (O_2249,N_29274,N_27684);
and UO_2250 (O_2250,N_28546,N_29660);
or UO_2251 (O_2251,N_27033,N_27752);
or UO_2252 (O_2252,N_29742,N_27330);
or UO_2253 (O_2253,N_29106,N_27699);
and UO_2254 (O_2254,N_28523,N_28379);
nor UO_2255 (O_2255,N_27338,N_28728);
or UO_2256 (O_2256,N_27883,N_27602);
or UO_2257 (O_2257,N_27397,N_29592);
and UO_2258 (O_2258,N_28172,N_27931);
xnor UO_2259 (O_2259,N_29809,N_29545);
nor UO_2260 (O_2260,N_27317,N_27492);
nand UO_2261 (O_2261,N_29199,N_27607);
nor UO_2262 (O_2262,N_27448,N_27716);
nor UO_2263 (O_2263,N_28618,N_28884);
and UO_2264 (O_2264,N_28788,N_28331);
and UO_2265 (O_2265,N_27088,N_29057);
and UO_2266 (O_2266,N_28219,N_28044);
and UO_2267 (O_2267,N_29453,N_27546);
nand UO_2268 (O_2268,N_27912,N_28573);
nor UO_2269 (O_2269,N_29477,N_27569);
nor UO_2270 (O_2270,N_29054,N_29205);
and UO_2271 (O_2271,N_27552,N_27120);
nor UO_2272 (O_2272,N_28403,N_29353);
or UO_2273 (O_2273,N_29742,N_29635);
nor UO_2274 (O_2274,N_28384,N_29475);
nor UO_2275 (O_2275,N_28865,N_28784);
nor UO_2276 (O_2276,N_27212,N_28411);
nand UO_2277 (O_2277,N_27293,N_28729);
or UO_2278 (O_2278,N_29963,N_28744);
nor UO_2279 (O_2279,N_27450,N_27833);
nor UO_2280 (O_2280,N_29535,N_28731);
and UO_2281 (O_2281,N_29845,N_27417);
nor UO_2282 (O_2282,N_27955,N_27174);
nor UO_2283 (O_2283,N_27490,N_27464);
nor UO_2284 (O_2284,N_27406,N_29315);
xor UO_2285 (O_2285,N_28566,N_28242);
nor UO_2286 (O_2286,N_28937,N_27074);
and UO_2287 (O_2287,N_29597,N_28069);
and UO_2288 (O_2288,N_27920,N_27660);
nor UO_2289 (O_2289,N_27577,N_28878);
xor UO_2290 (O_2290,N_27279,N_29996);
and UO_2291 (O_2291,N_27649,N_27447);
nor UO_2292 (O_2292,N_28987,N_27745);
or UO_2293 (O_2293,N_29781,N_27841);
nor UO_2294 (O_2294,N_27393,N_29932);
nor UO_2295 (O_2295,N_29213,N_28917);
and UO_2296 (O_2296,N_28647,N_28095);
nand UO_2297 (O_2297,N_28225,N_29828);
nand UO_2298 (O_2298,N_28697,N_29892);
xor UO_2299 (O_2299,N_28445,N_27740);
nand UO_2300 (O_2300,N_29429,N_29722);
and UO_2301 (O_2301,N_29746,N_27279);
or UO_2302 (O_2302,N_28904,N_28387);
and UO_2303 (O_2303,N_28741,N_28715);
and UO_2304 (O_2304,N_27418,N_28403);
nand UO_2305 (O_2305,N_29507,N_27466);
nand UO_2306 (O_2306,N_28185,N_28761);
and UO_2307 (O_2307,N_28535,N_27084);
xor UO_2308 (O_2308,N_27779,N_29930);
and UO_2309 (O_2309,N_27548,N_28659);
xor UO_2310 (O_2310,N_28168,N_29538);
nand UO_2311 (O_2311,N_29794,N_27039);
or UO_2312 (O_2312,N_27237,N_28397);
nand UO_2313 (O_2313,N_27436,N_27489);
xor UO_2314 (O_2314,N_27809,N_29928);
or UO_2315 (O_2315,N_29899,N_29191);
nand UO_2316 (O_2316,N_29881,N_28236);
and UO_2317 (O_2317,N_27414,N_27494);
or UO_2318 (O_2318,N_27194,N_27935);
nand UO_2319 (O_2319,N_29899,N_29151);
nand UO_2320 (O_2320,N_28054,N_27671);
or UO_2321 (O_2321,N_29739,N_29903);
nor UO_2322 (O_2322,N_28704,N_27265);
and UO_2323 (O_2323,N_29925,N_29462);
nand UO_2324 (O_2324,N_28767,N_29194);
or UO_2325 (O_2325,N_28179,N_28901);
xor UO_2326 (O_2326,N_28530,N_28116);
xnor UO_2327 (O_2327,N_27508,N_27127);
and UO_2328 (O_2328,N_28498,N_29574);
or UO_2329 (O_2329,N_29124,N_28527);
or UO_2330 (O_2330,N_29799,N_28119);
nand UO_2331 (O_2331,N_29118,N_27609);
xor UO_2332 (O_2332,N_29482,N_28402);
xor UO_2333 (O_2333,N_27113,N_29611);
nand UO_2334 (O_2334,N_28205,N_29005);
nand UO_2335 (O_2335,N_27718,N_28397);
or UO_2336 (O_2336,N_28769,N_28435);
or UO_2337 (O_2337,N_29303,N_28564);
nand UO_2338 (O_2338,N_29672,N_28819);
or UO_2339 (O_2339,N_28249,N_29882);
nor UO_2340 (O_2340,N_29325,N_29283);
and UO_2341 (O_2341,N_29361,N_28552);
and UO_2342 (O_2342,N_29668,N_29297);
nor UO_2343 (O_2343,N_28343,N_27034);
xnor UO_2344 (O_2344,N_28167,N_27084);
nand UO_2345 (O_2345,N_28236,N_27772);
nor UO_2346 (O_2346,N_29439,N_28644);
xor UO_2347 (O_2347,N_29339,N_28894);
or UO_2348 (O_2348,N_29052,N_27767);
or UO_2349 (O_2349,N_27797,N_29250);
nor UO_2350 (O_2350,N_27408,N_28996);
and UO_2351 (O_2351,N_29383,N_28075);
nor UO_2352 (O_2352,N_29642,N_29765);
nor UO_2353 (O_2353,N_28251,N_28571);
xor UO_2354 (O_2354,N_29021,N_27426);
and UO_2355 (O_2355,N_29102,N_27976);
xnor UO_2356 (O_2356,N_28002,N_29958);
xnor UO_2357 (O_2357,N_28363,N_29746);
and UO_2358 (O_2358,N_28760,N_28174);
or UO_2359 (O_2359,N_28800,N_28624);
or UO_2360 (O_2360,N_28410,N_29711);
and UO_2361 (O_2361,N_27413,N_29326);
and UO_2362 (O_2362,N_29827,N_28266);
xnor UO_2363 (O_2363,N_27347,N_29944);
nor UO_2364 (O_2364,N_29771,N_29641);
and UO_2365 (O_2365,N_28531,N_29030);
xor UO_2366 (O_2366,N_29821,N_28139);
nand UO_2367 (O_2367,N_28459,N_27138);
or UO_2368 (O_2368,N_29088,N_29023);
nor UO_2369 (O_2369,N_29838,N_28324);
xnor UO_2370 (O_2370,N_29784,N_29961);
nor UO_2371 (O_2371,N_27558,N_29244);
nand UO_2372 (O_2372,N_28355,N_28530);
nor UO_2373 (O_2373,N_27335,N_29313);
nor UO_2374 (O_2374,N_28738,N_28256);
xnor UO_2375 (O_2375,N_28781,N_29323);
nand UO_2376 (O_2376,N_29042,N_28301);
xnor UO_2377 (O_2377,N_28284,N_28752);
xnor UO_2378 (O_2378,N_29010,N_28648);
xnor UO_2379 (O_2379,N_28125,N_29248);
and UO_2380 (O_2380,N_29024,N_29964);
and UO_2381 (O_2381,N_27956,N_28155);
nand UO_2382 (O_2382,N_28083,N_27831);
xnor UO_2383 (O_2383,N_28325,N_29527);
nand UO_2384 (O_2384,N_29201,N_28132);
nor UO_2385 (O_2385,N_28338,N_27727);
nand UO_2386 (O_2386,N_29032,N_28038);
or UO_2387 (O_2387,N_27645,N_27673);
nand UO_2388 (O_2388,N_29711,N_29887);
nand UO_2389 (O_2389,N_29368,N_27460);
nor UO_2390 (O_2390,N_28374,N_29988);
nor UO_2391 (O_2391,N_29645,N_28565);
and UO_2392 (O_2392,N_29157,N_27192);
nand UO_2393 (O_2393,N_28843,N_29356);
xnor UO_2394 (O_2394,N_29728,N_28919);
or UO_2395 (O_2395,N_29958,N_27908);
nand UO_2396 (O_2396,N_29659,N_28180);
and UO_2397 (O_2397,N_29370,N_27935);
and UO_2398 (O_2398,N_28604,N_28700);
nor UO_2399 (O_2399,N_29377,N_29506);
or UO_2400 (O_2400,N_28263,N_27321);
xnor UO_2401 (O_2401,N_28924,N_29789);
nand UO_2402 (O_2402,N_28852,N_27833);
or UO_2403 (O_2403,N_27013,N_29432);
nor UO_2404 (O_2404,N_28404,N_28675);
or UO_2405 (O_2405,N_27271,N_28249);
nor UO_2406 (O_2406,N_28259,N_28058);
xnor UO_2407 (O_2407,N_28989,N_28371);
xor UO_2408 (O_2408,N_28953,N_29948);
or UO_2409 (O_2409,N_28460,N_28155);
xor UO_2410 (O_2410,N_29294,N_27934);
nand UO_2411 (O_2411,N_28059,N_29576);
and UO_2412 (O_2412,N_27738,N_29526);
or UO_2413 (O_2413,N_29135,N_28633);
or UO_2414 (O_2414,N_28579,N_29286);
nor UO_2415 (O_2415,N_29855,N_29768);
nor UO_2416 (O_2416,N_28755,N_28298);
nand UO_2417 (O_2417,N_27646,N_27972);
and UO_2418 (O_2418,N_29911,N_27833);
and UO_2419 (O_2419,N_27844,N_28796);
nand UO_2420 (O_2420,N_27876,N_28469);
and UO_2421 (O_2421,N_28023,N_27904);
nor UO_2422 (O_2422,N_29590,N_29989);
or UO_2423 (O_2423,N_29708,N_28904);
nand UO_2424 (O_2424,N_29673,N_28729);
nor UO_2425 (O_2425,N_29202,N_29991);
nor UO_2426 (O_2426,N_29912,N_29283);
and UO_2427 (O_2427,N_28459,N_29990);
and UO_2428 (O_2428,N_28917,N_29611);
nor UO_2429 (O_2429,N_29308,N_28946);
nand UO_2430 (O_2430,N_28171,N_29552);
or UO_2431 (O_2431,N_29642,N_28100);
nand UO_2432 (O_2432,N_29329,N_27804);
and UO_2433 (O_2433,N_27957,N_27584);
nor UO_2434 (O_2434,N_29919,N_27585);
or UO_2435 (O_2435,N_28402,N_27927);
nor UO_2436 (O_2436,N_27272,N_27633);
and UO_2437 (O_2437,N_27460,N_27969);
xnor UO_2438 (O_2438,N_27714,N_28942);
nor UO_2439 (O_2439,N_28645,N_28926);
nand UO_2440 (O_2440,N_28390,N_29280);
xor UO_2441 (O_2441,N_29339,N_29252);
or UO_2442 (O_2442,N_27455,N_27607);
and UO_2443 (O_2443,N_28088,N_27338);
nand UO_2444 (O_2444,N_28941,N_29213);
nor UO_2445 (O_2445,N_29877,N_27379);
and UO_2446 (O_2446,N_29797,N_29118);
xor UO_2447 (O_2447,N_28173,N_27114);
nand UO_2448 (O_2448,N_27442,N_27206);
nor UO_2449 (O_2449,N_27817,N_28362);
and UO_2450 (O_2450,N_27199,N_27406);
nand UO_2451 (O_2451,N_27779,N_29319);
and UO_2452 (O_2452,N_29948,N_29050);
nand UO_2453 (O_2453,N_27580,N_27736);
or UO_2454 (O_2454,N_27312,N_27954);
and UO_2455 (O_2455,N_27401,N_27687);
or UO_2456 (O_2456,N_27629,N_29694);
nor UO_2457 (O_2457,N_29226,N_29815);
or UO_2458 (O_2458,N_27326,N_27821);
nand UO_2459 (O_2459,N_29142,N_28039);
and UO_2460 (O_2460,N_29544,N_28863);
xnor UO_2461 (O_2461,N_27494,N_27470);
xnor UO_2462 (O_2462,N_29243,N_29567);
nor UO_2463 (O_2463,N_27248,N_28384);
nor UO_2464 (O_2464,N_28660,N_29152);
nand UO_2465 (O_2465,N_29354,N_28477);
nand UO_2466 (O_2466,N_29851,N_28749);
and UO_2467 (O_2467,N_29378,N_29356);
xor UO_2468 (O_2468,N_27245,N_29601);
or UO_2469 (O_2469,N_28753,N_27125);
and UO_2470 (O_2470,N_29353,N_27781);
nand UO_2471 (O_2471,N_29997,N_27092);
nand UO_2472 (O_2472,N_27928,N_28713);
nand UO_2473 (O_2473,N_27089,N_29937);
nor UO_2474 (O_2474,N_27775,N_27063);
and UO_2475 (O_2475,N_28386,N_27572);
or UO_2476 (O_2476,N_27982,N_29913);
nand UO_2477 (O_2477,N_29454,N_29104);
and UO_2478 (O_2478,N_27542,N_27343);
or UO_2479 (O_2479,N_28275,N_28739);
nand UO_2480 (O_2480,N_27416,N_27544);
xnor UO_2481 (O_2481,N_28092,N_28187);
and UO_2482 (O_2482,N_28900,N_29895);
xnor UO_2483 (O_2483,N_28340,N_27236);
nor UO_2484 (O_2484,N_29741,N_29744);
nor UO_2485 (O_2485,N_28839,N_29505);
nor UO_2486 (O_2486,N_28441,N_28312);
nor UO_2487 (O_2487,N_28676,N_27431);
and UO_2488 (O_2488,N_29227,N_27846);
nand UO_2489 (O_2489,N_28536,N_28924);
nand UO_2490 (O_2490,N_28170,N_27494);
or UO_2491 (O_2491,N_28898,N_28075);
nand UO_2492 (O_2492,N_29565,N_28357);
nor UO_2493 (O_2493,N_28059,N_29746);
or UO_2494 (O_2494,N_27987,N_27723);
or UO_2495 (O_2495,N_27159,N_27500);
or UO_2496 (O_2496,N_29039,N_28990);
and UO_2497 (O_2497,N_27669,N_27250);
xor UO_2498 (O_2498,N_28184,N_27812);
and UO_2499 (O_2499,N_28059,N_29629);
xor UO_2500 (O_2500,N_29105,N_29972);
or UO_2501 (O_2501,N_28882,N_29229);
and UO_2502 (O_2502,N_28942,N_29372);
nor UO_2503 (O_2503,N_28702,N_27354);
xor UO_2504 (O_2504,N_28483,N_28247);
and UO_2505 (O_2505,N_29238,N_29465);
and UO_2506 (O_2506,N_27444,N_29004);
nand UO_2507 (O_2507,N_29767,N_27835);
xor UO_2508 (O_2508,N_28017,N_27255);
and UO_2509 (O_2509,N_28895,N_28037);
nor UO_2510 (O_2510,N_27559,N_27705);
or UO_2511 (O_2511,N_27603,N_27352);
nand UO_2512 (O_2512,N_28650,N_29937);
nand UO_2513 (O_2513,N_27609,N_29858);
nand UO_2514 (O_2514,N_28012,N_27558);
nor UO_2515 (O_2515,N_29293,N_29337);
nor UO_2516 (O_2516,N_28604,N_29506);
and UO_2517 (O_2517,N_27077,N_29496);
nand UO_2518 (O_2518,N_27139,N_28180);
or UO_2519 (O_2519,N_29441,N_27118);
or UO_2520 (O_2520,N_27610,N_27539);
and UO_2521 (O_2521,N_27360,N_29612);
nor UO_2522 (O_2522,N_29661,N_28033);
xor UO_2523 (O_2523,N_29321,N_29140);
or UO_2524 (O_2524,N_28795,N_29672);
xnor UO_2525 (O_2525,N_28543,N_29691);
xor UO_2526 (O_2526,N_29515,N_28478);
xor UO_2527 (O_2527,N_29071,N_29826);
nor UO_2528 (O_2528,N_27345,N_29918);
nand UO_2529 (O_2529,N_28716,N_27083);
nand UO_2530 (O_2530,N_28474,N_28534);
or UO_2531 (O_2531,N_28696,N_28623);
and UO_2532 (O_2532,N_27883,N_27003);
and UO_2533 (O_2533,N_29094,N_29680);
xnor UO_2534 (O_2534,N_29264,N_28998);
nor UO_2535 (O_2535,N_27984,N_28492);
and UO_2536 (O_2536,N_28308,N_27715);
xor UO_2537 (O_2537,N_29040,N_27515);
nand UO_2538 (O_2538,N_28568,N_28170);
and UO_2539 (O_2539,N_28265,N_28449);
nand UO_2540 (O_2540,N_28744,N_28123);
and UO_2541 (O_2541,N_28641,N_27326);
or UO_2542 (O_2542,N_28180,N_28527);
xnor UO_2543 (O_2543,N_27241,N_28940);
or UO_2544 (O_2544,N_29421,N_29321);
nand UO_2545 (O_2545,N_27281,N_28620);
nand UO_2546 (O_2546,N_27633,N_27434);
or UO_2547 (O_2547,N_27754,N_27006);
or UO_2548 (O_2548,N_28952,N_29866);
or UO_2549 (O_2549,N_28672,N_28822);
nand UO_2550 (O_2550,N_29557,N_29783);
xor UO_2551 (O_2551,N_27637,N_29632);
or UO_2552 (O_2552,N_28531,N_29127);
nand UO_2553 (O_2553,N_28715,N_27474);
nand UO_2554 (O_2554,N_29287,N_29568);
nand UO_2555 (O_2555,N_29020,N_29992);
or UO_2556 (O_2556,N_28786,N_29031);
nand UO_2557 (O_2557,N_27594,N_29048);
or UO_2558 (O_2558,N_28992,N_29779);
or UO_2559 (O_2559,N_27752,N_29136);
nor UO_2560 (O_2560,N_29402,N_27727);
xor UO_2561 (O_2561,N_27099,N_28197);
nor UO_2562 (O_2562,N_28348,N_28914);
and UO_2563 (O_2563,N_29016,N_29392);
xnor UO_2564 (O_2564,N_29979,N_28191);
nand UO_2565 (O_2565,N_27840,N_29402);
or UO_2566 (O_2566,N_27232,N_29556);
and UO_2567 (O_2567,N_27143,N_29211);
and UO_2568 (O_2568,N_29324,N_28010);
and UO_2569 (O_2569,N_28830,N_27986);
nand UO_2570 (O_2570,N_27992,N_29956);
xnor UO_2571 (O_2571,N_27245,N_28556);
nor UO_2572 (O_2572,N_27007,N_29757);
or UO_2573 (O_2573,N_28929,N_27497);
nor UO_2574 (O_2574,N_28212,N_29257);
xnor UO_2575 (O_2575,N_29896,N_28040);
or UO_2576 (O_2576,N_29684,N_28045);
nand UO_2577 (O_2577,N_29037,N_29378);
or UO_2578 (O_2578,N_28845,N_27213);
nor UO_2579 (O_2579,N_28962,N_28393);
nor UO_2580 (O_2580,N_27592,N_28409);
nor UO_2581 (O_2581,N_29479,N_29444);
or UO_2582 (O_2582,N_28301,N_27220);
nor UO_2583 (O_2583,N_27240,N_28028);
or UO_2584 (O_2584,N_29633,N_27983);
and UO_2585 (O_2585,N_28478,N_28230);
and UO_2586 (O_2586,N_28316,N_28533);
xor UO_2587 (O_2587,N_29770,N_29472);
and UO_2588 (O_2588,N_28336,N_28700);
nand UO_2589 (O_2589,N_28063,N_27909);
nor UO_2590 (O_2590,N_29479,N_27485);
xnor UO_2591 (O_2591,N_29854,N_27251);
or UO_2592 (O_2592,N_29486,N_29308);
nand UO_2593 (O_2593,N_29175,N_29085);
nor UO_2594 (O_2594,N_28963,N_27336);
or UO_2595 (O_2595,N_28783,N_27290);
and UO_2596 (O_2596,N_29137,N_28965);
and UO_2597 (O_2597,N_28504,N_29844);
or UO_2598 (O_2598,N_27880,N_29200);
xor UO_2599 (O_2599,N_28263,N_28861);
and UO_2600 (O_2600,N_29856,N_27171);
or UO_2601 (O_2601,N_27114,N_29521);
or UO_2602 (O_2602,N_29340,N_28774);
xor UO_2603 (O_2603,N_29224,N_28450);
nor UO_2604 (O_2604,N_28354,N_27234);
and UO_2605 (O_2605,N_27967,N_27102);
or UO_2606 (O_2606,N_27073,N_27830);
nor UO_2607 (O_2607,N_27361,N_29635);
nand UO_2608 (O_2608,N_28297,N_29974);
or UO_2609 (O_2609,N_29914,N_28634);
xnor UO_2610 (O_2610,N_28117,N_28918);
xnor UO_2611 (O_2611,N_27995,N_29232);
or UO_2612 (O_2612,N_29571,N_29546);
or UO_2613 (O_2613,N_28079,N_29685);
xor UO_2614 (O_2614,N_27631,N_29553);
nor UO_2615 (O_2615,N_27492,N_29380);
nor UO_2616 (O_2616,N_29868,N_27390);
nor UO_2617 (O_2617,N_29158,N_28802);
and UO_2618 (O_2618,N_29414,N_29704);
nand UO_2619 (O_2619,N_29105,N_29014);
nand UO_2620 (O_2620,N_27224,N_27565);
xnor UO_2621 (O_2621,N_28799,N_27233);
nand UO_2622 (O_2622,N_29658,N_27436);
or UO_2623 (O_2623,N_27431,N_29084);
and UO_2624 (O_2624,N_27410,N_29838);
or UO_2625 (O_2625,N_28366,N_29945);
nand UO_2626 (O_2626,N_28150,N_28580);
nand UO_2627 (O_2627,N_28284,N_29366);
nor UO_2628 (O_2628,N_28267,N_29143);
or UO_2629 (O_2629,N_29141,N_28433);
nor UO_2630 (O_2630,N_29683,N_27588);
nor UO_2631 (O_2631,N_27829,N_29719);
or UO_2632 (O_2632,N_29846,N_29953);
nor UO_2633 (O_2633,N_29387,N_27893);
nor UO_2634 (O_2634,N_29119,N_29570);
nand UO_2635 (O_2635,N_28258,N_27617);
nor UO_2636 (O_2636,N_29574,N_27877);
nor UO_2637 (O_2637,N_29827,N_29077);
and UO_2638 (O_2638,N_29441,N_28780);
or UO_2639 (O_2639,N_28874,N_28257);
nand UO_2640 (O_2640,N_28900,N_28112);
nand UO_2641 (O_2641,N_27923,N_27702);
nor UO_2642 (O_2642,N_28984,N_28432);
xor UO_2643 (O_2643,N_28936,N_29710);
and UO_2644 (O_2644,N_27572,N_28620);
and UO_2645 (O_2645,N_28590,N_28277);
nand UO_2646 (O_2646,N_27586,N_28795);
xnor UO_2647 (O_2647,N_29853,N_28192);
and UO_2648 (O_2648,N_29524,N_29548);
nand UO_2649 (O_2649,N_29243,N_27134);
xor UO_2650 (O_2650,N_28593,N_27348);
and UO_2651 (O_2651,N_28449,N_29652);
nor UO_2652 (O_2652,N_28963,N_27641);
and UO_2653 (O_2653,N_29305,N_27612);
xnor UO_2654 (O_2654,N_28366,N_29944);
or UO_2655 (O_2655,N_28260,N_28855);
nor UO_2656 (O_2656,N_29123,N_28014);
or UO_2657 (O_2657,N_29900,N_29572);
nand UO_2658 (O_2658,N_27880,N_27311);
nand UO_2659 (O_2659,N_27180,N_29349);
and UO_2660 (O_2660,N_28425,N_27300);
nor UO_2661 (O_2661,N_29598,N_28035);
nor UO_2662 (O_2662,N_27499,N_27556);
or UO_2663 (O_2663,N_28067,N_29282);
xor UO_2664 (O_2664,N_27525,N_27874);
nor UO_2665 (O_2665,N_27336,N_28048);
or UO_2666 (O_2666,N_28998,N_28682);
nand UO_2667 (O_2667,N_29729,N_28358);
and UO_2668 (O_2668,N_29939,N_28877);
xnor UO_2669 (O_2669,N_29101,N_28473);
xnor UO_2670 (O_2670,N_27623,N_27013);
and UO_2671 (O_2671,N_29511,N_27540);
xor UO_2672 (O_2672,N_27555,N_29356);
or UO_2673 (O_2673,N_29134,N_27474);
and UO_2674 (O_2674,N_29164,N_27030);
and UO_2675 (O_2675,N_27561,N_27193);
or UO_2676 (O_2676,N_28435,N_28254);
and UO_2677 (O_2677,N_28613,N_29903);
xnor UO_2678 (O_2678,N_29377,N_29770);
and UO_2679 (O_2679,N_28626,N_29069);
or UO_2680 (O_2680,N_28833,N_29564);
nand UO_2681 (O_2681,N_27108,N_29335);
nor UO_2682 (O_2682,N_29460,N_27809);
nand UO_2683 (O_2683,N_28936,N_28237);
and UO_2684 (O_2684,N_28541,N_27219);
or UO_2685 (O_2685,N_29921,N_29385);
and UO_2686 (O_2686,N_29559,N_27047);
nor UO_2687 (O_2687,N_29505,N_29665);
and UO_2688 (O_2688,N_28193,N_29584);
xor UO_2689 (O_2689,N_27000,N_29278);
xor UO_2690 (O_2690,N_28841,N_28345);
nand UO_2691 (O_2691,N_28175,N_27306);
and UO_2692 (O_2692,N_29527,N_29004);
xor UO_2693 (O_2693,N_29095,N_28783);
xor UO_2694 (O_2694,N_29821,N_29581);
nor UO_2695 (O_2695,N_29276,N_28738);
nor UO_2696 (O_2696,N_29307,N_27302);
xor UO_2697 (O_2697,N_28175,N_29978);
or UO_2698 (O_2698,N_29124,N_27304);
or UO_2699 (O_2699,N_28820,N_29844);
nand UO_2700 (O_2700,N_29916,N_29036);
or UO_2701 (O_2701,N_28479,N_29993);
nor UO_2702 (O_2702,N_29374,N_29503);
and UO_2703 (O_2703,N_28153,N_27073);
xnor UO_2704 (O_2704,N_28990,N_28697);
nor UO_2705 (O_2705,N_27081,N_28588);
and UO_2706 (O_2706,N_28368,N_29392);
nor UO_2707 (O_2707,N_27544,N_29107);
or UO_2708 (O_2708,N_27086,N_29757);
xor UO_2709 (O_2709,N_29696,N_29599);
nand UO_2710 (O_2710,N_27507,N_28065);
or UO_2711 (O_2711,N_29754,N_29240);
nand UO_2712 (O_2712,N_29988,N_29581);
nor UO_2713 (O_2713,N_29156,N_27123);
and UO_2714 (O_2714,N_29671,N_27966);
nor UO_2715 (O_2715,N_28277,N_28281);
or UO_2716 (O_2716,N_28135,N_29328);
and UO_2717 (O_2717,N_29968,N_27810);
and UO_2718 (O_2718,N_27372,N_27052);
xnor UO_2719 (O_2719,N_29472,N_28453);
nor UO_2720 (O_2720,N_28106,N_27404);
xnor UO_2721 (O_2721,N_29057,N_27791);
nor UO_2722 (O_2722,N_29602,N_29775);
nand UO_2723 (O_2723,N_27204,N_28537);
nand UO_2724 (O_2724,N_28964,N_27902);
nand UO_2725 (O_2725,N_28398,N_27090);
xor UO_2726 (O_2726,N_29056,N_28436);
xor UO_2727 (O_2727,N_29307,N_28568);
nor UO_2728 (O_2728,N_27042,N_28657);
or UO_2729 (O_2729,N_29340,N_27379);
xnor UO_2730 (O_2730,N_28245,N_28065);
nand UO_2731 (O_2731,N_27119,N_27751);
or UO_2732 (O_2732,N_29894,N_27094);
nor UO_2733 (O_2733,N_27264,N_28609);
and UO_2734 (O_2734,N_27970,N_29909);
nor UO_2735 (O_2735,N_27529,N_27838);
or UO_2736 (O_2736,N_29804,N_28238);
xor UO_2737 (O_2737,N_28625,N_28407);
nor UO_2738 (O_2738,N_29990,N_29146);
nor UO_2739 (O_2739,N_29485,N_27350);
nor UO_2740 (O_2740,N_29055,N_27245);
or UO_2741 (O_2741,N_29810,N_28996);
xor UO_2742 (O_2742,N_28603,N_29478);
nand UO_2743 (O_2743,N_29334,N_28942);
nand UO_2744 (O_2744,N_27407,N_29131);
nand UO_2745 (O_2745,N_29332,N_28554);
nor UO_2746 (O_2746,N_29315,N_27418);
and UO_2747 (O_2747,N_27332,N_28779);
or UO_2748 (O_2748,N_29956,N_29973);
nand UO_2749 (O_2749,N_29421,N_29502);
or UO_2750 (O_2750,N_27577,N_27288);
xor UO_2751 (O_2751,N_28949,N_27407);
nor UO_2752 (O_2752,N_27397,N_29969);
nand UO_2753 (O_2753,N_29246,N_28375);
or UO_2754 (O_2754,N_27717,N_29929);
nand UO_2755 (O_2755,N_29737,N_28634);
xnor UO_2756 (O_2756,N_29118,N_27096);
or UO_2757 (O_2757,N_27719,N_28517);
nor UO_2758 (O_2758,N_29023,N_28790);
and UO_2759 (O_2759,N_27021,N_28564);
or UO_2760 (O_2760,N_27147,N_29471);
and UO_2761 (O_2761,N_27173,N_29624);
or UO_2762 (O_2762,N_29129,N_29791);
or UO_2763 (O_2763,N_27016,N_27479);
and UO_2764 (O_2764,N_29998,N_28336);
nor UO_2765 (O_2765,N_28498,N_27840);
xnor UO_2766 (O_2766,N_28757,N_27724);
nor UO_2767 (O_2767,N_28385,N_28731);
and UO_2768 (O_2768,N_27345,N_29365);
xor UO_2769 (O_2769,N_28527,N_27305);
nand UO_2770 (O_2770,N_28288,N_27842);
xnor UO_2771 (O_2771,N_27910,N_29809);
nor UO_2772 (O_2772,N_28268,N_27927);
or UO_2773 (O_2773,N_27355,N_29814);
nor UO_2774 (O_2774,N_29747,N_29318);
nand UO_2775 (O_2775,N_29937,N_27027);
nand UO_2776 (O_2776,N_29165,N_29738);
and UO_2777 (O_2777,N_27412,N_27687);
nand UO_2778 (O_2778,N_28214,N_27020);
nor UO_2779 (O_2779,N_29526,N_28836);
or UO_2780 (O_2780,N_27371,N_27541);
xnor UO_2781 (O_2781,N_27090,N_29228);
nand UO_2782 (O_2782,N_27155,N_28180);
or UO_2783 (O_2783,N_29747,N_29972);
nor UO_2784 (O_2784,N_27434,N_27885);
nand UO_2785 (O_2785,N_29692,N_29081);
nand UO_2786 (O_2786,N_29333,N_27349);
or UO_2787 (O_2787,N_29526,N_29158);
nor UO_2788 (O_2788,N_28608,N_28462);
or UO_2789 (O_2789,N_29010,N_27065);
xor UO_2790 (O_2790,N_28481,N_28556);
or UO_2791 (O_2791,N_27370,N_28479);
xor UO_2792 (O_2792,N_29265,N_27000);
nor UO_2793 (O_2793,N_27109,N_29180);
or UO_2794 (O_2794,N_27669,N_28508);
nand UO_2795 (O_2795,N_28834,N_27522);
nand UO_2796 (O_2796,N_28396,N_29795);
and UO_2797 (O_2797,N_28874,N_28509);
or UO_2798 (O_2798,N_29476,N_27736);
or UO_2799 (O_2799,N_29427,N_29342);
xor UO_2800 (O_2800,N_28097,N_29216);
xor UO_2801 (O_2801,N_29997,N_28875);
and UO_2802 (O_2802,N_28464,N_28666);
nand UO_2803 (O_2803,N_29133,N_27081);
and UO_2804 (O_2804,N_28110,N_27015);
nand UO_2805 (O_2805,N_28929,N_27057);
or UO_2806 (O_2806,N_29911,N_29583);
xnor UO_2807 (O_2807,N_28611,N_27217);
nand UO_2808 (O_2808,N_27025,N_28823);
nor UO_2809 (O_2809,N_29773,N_28069);
and UO_2810 (O_2810,N_28192,N_27722);
nand UO_2811 (O_2811,N_28134,N_27368);
nand UO_2812 (O_2812,N_27033,N_28597);
xnor UO_2813 (O_2813,N_27859,N_29059);
and UO_2814 (O_2814,N_28918,N_27551);
xnor UO_2815 (O_2815,N_28990,N_27084);
nor UO_2816 (O_2816,N_27470,N_28869);
nor UO_2817 (O_2817,N_27477,N_27796);
xor UO_2818 (O_2818,N_29571,N_27814);
or UO_2819 (O_2819,N_27262,N_27648);
nor UO_2820 (O_2820,N_29495,N_28239);
nand UO_2821 (O_2821,N_27938,N_27160);
xnor UO_2822 (O_2822,N_27636,N_29015);
nor UO_2823 (O_2823,N_29376,N_28865);
nor UO_2824 (O_2824,N_29945,N_29280);
nor UO_2825 (O_2825,N_28208,N_27456);
nand UO_2826 (O_2826,N_27931,N_29180);
nand UO_2827 (O_2827,N_29619,N_28267);
or UO_2828 (O_2828,N_28468,N_28138);
xnor UO_2829 (O_2829,N_28042,N_29335);
or UO_2830 (O_2830,N_28052,N_29242);
nand UO_2831 (O_2831,N_27522,N_27532);
or UO_2832 (O_2832,N_28125,N_29343);
and UO_2833 (O_2833,N_29380,N_29884);
and UO_2834 (O_2834,N_28184,N_29075);
xnor UO_2835 (O_2835,N_28068,N_27604);
and UO_2836 (O_2836,N_27485,N_27749);
nor UO_2837 (O_2837,N_29884,N_27001);
xnor UO_2838 (O_2838,N_27569,N_29472);
or UO_2839 (O_2839,N_27010,N_29420);
nor UO_2840 (O_2840,N_28369,N_29324);
xnor UO_2841 (O_2841,N_29556,N_28858);
nand UO_2842 (O_2842,N_27819,N_27334);
xnor UO_2843 (O_2843,N_28934,N_28433);
or UO_2844 (O_2844,N_29909,N_28144);
or UO_2845 (O_2845,N_28328,N_28800);
xnor UO_2846 (O_2846,N_29050,N_27671);
nand UO_2847 (O_2847,N_27275,N_29114);
xor UO_2848 (O_2848,N_27815,N_27435);
and UO_2849 (O_2849,N_27644,N_29742);
nand UO_2850 (O_2850,N_27265,N_28090);
nor UO_2851 (O_2851,N_27272,N_29430);
nand UO_2852 (O_2852,N_28000,N_29099);
xor UO_2853 (O_2853,N_29966,N_29702);
or UO_2854 (O_2854,N_27727,N_27006);
or UO_2855 (O_2855,N_27505,N_27655);
nor UO_2856 (O_2856,N_27620,N_27371);
xnor UO_2857 (O_2857,N_29492,N_27965);
xor UO_2858 (O_2858,N_28939,N_29285);
nor UO_2859 (O_2859,N_29395,N_28032);
xnor UO_2860 (O_2860,N_28281,N_28056);
xnor UO_2861 (O_2861,N_28838,N_27040);
and UO_2862 (O_2862,N_27268,N_27393);
or UO_2863 (O_2863,N_27370,N_29569);
xnor UO_2864 (O_2864,N_27406,N_27151);
xor UO_2865 (O_2865,N_28870,N_28913);
or UO_2866 (O_2866,N_27110,N_28925);
nor UO_2867 (O_2867,N_27235,N_29546);
xnor UO_2868 (O_2868,N_27362,N_29728);
xnor UO_2869 (O_2869,N_27766,N_29562);
nand UO_2870 (O_2870,N_28608,N_28509);
nand UO_2871 (O_2871,N_29582,N_27899);
or UO_2872 (O_2872,N_29002,N_27604);
nor UO_2873 (O_2873,N_28665,N_29110);
nor UO_2874 (O_2874,N_28407,N_28813);
or UO_2875 (O_2875,N_28205,N_28833);
and UO_2876 (O_2876,N_28175,N_29427);
nand UO_2877 (O_2877,N_28017,N_27116);
nand UO_2878 (O_2878,N_29600,N_27138);
nor UO_2879 (O_2879,N_29344,N_28261);
and UO_2880 (O_2880,N_28943,N_29802);
nor UO_2881 (O_2881,N_27194,N_29070);
xnor UO_2882 (O_2882,N_28464,N_28177);
or UO_2883 (O_2883,N_28097,N_29239);
nand UO_2884 (O_2884,N_29466,N_27445);
xnor UO_2885 (O_2885,N_29178,N_27422);
nor UO_2886 (O_2886,N_28593,N_29566);
or UO_2887 (O_2887,N_28426,N_29612);
and UO_2888 (O_2888,N_28402,N_28188);
nor UO_2889 (O_2889,N_28255,N_27765);
and UO_2890 (O_2890,N_27689,N_28264);
or UO_2891 (O_2891,N_27379,N_29224);
xnor UO_2892 (O_2892,N_27586,N_28945);
nor UO_2893 (O_2893,N_29901,N_28943);
and UO_2894 (O_2894,N_29010,N_29764);
nor UO_2895 (O_2895,N_28224,N_29933);
or UO_2896 (O_2896,N_27522,N_27901);
nor UO_2897 (O_2897,N_29096,N_29069);
xor UO_2898 (O_2898,N_27103,N_27381);
nand UO_2899 (O_2899,N_29274,N_29899);
xnor UO_2900 (O_2900,N_29149,N_29527);
nand UO_2901 (O_2901,N_28035,N_27918);
nor UO_2902 (O_2902,N_27469,N_28291);
xor UO_2903 (O_2903,N_27632,N_28695);
nand UO_2904 (O_2904,N_29286,N_29534);
and UO_2905 (O_2905,N_27218,N_29691);
nor UO_2906 (O_2906,N_27897,N_29792);
nor UO_2907 (O_2907,N_28873,N_27416);
or UO_2908 (O_2908,N_28424,N_29371);
or UO_2909 (O_2909,N_27860,N_29710);
and UO_2910 (O_2910,N_27047,N_28460);
or UO_2911 (O_2911,N_29041,N_29822);
and UO_2912 (O_2912,N_27721,N_27554);
nand UO_2913 (O_2913,N_29113,N_27227);
or UO_2914 (O_2914,N_27022,N_27377);
or UO_2915 (O_2915,N_27578,N_28568);
nor UO_2916 (O_2916,N_29663,N_27965);
nand UO_2917 (O_2917,N_28465,N_27742);
xor UO_2918 (O_2918,N_28738,N_29000);
nand UO_2919 (O_2919,N_28243,N_27076);
xnor UO_2920 (O_2920,N_28919,N_28465);
and UO_2921 (O_2921,N_29926,N_28453);
or UO_2922 (O_2922,N_27425,N_28591);
nand UO_2923 (O_2923,N_27749,N_29194);
nand UO_2924 (O_2924,N_29385,N_27301);
or UO_2925 (O_2925,N_29904,N_28260);
and UO_2926 (O_2926,N_28471,N_27770);
nand UO_2927 (O_2927,N_28654,N_29245);
nor UO_2928 (O_2928,N_28539,N_27879);
and UO_2929 (O_2929,N_27584,N_29151);
and UO_2930 (O_2930,N_28731,N_28168);
and UO_2931 (O_2931,N_29214,N_29051);
and UO_2932 (O_2932,N_29681,N_29190);
or UO_2933 (O_2933,N_28820,N_27937);
xnor UO_2934 (O_2934,N_28458,N_29305);
xor UO_2935 (O_2935,N_27280,N_28422);
nor UO_2936 (O_2936,N_29676,N_28719);
nand UO_2937 (O_2937,N_28681,N_27160);
or UO_2938 (O_2938,N_27502,N_27370);
nor UO_2939 (O_2939,N_27580,N_27843);
xnor UO_2940 (O_2940,N_28223,N_28430);
xor UO_2941 (O_2941,N_27686,N_28087);
xnor UO_2942 (O_2942,N_27192,N_28718);
xor UO_2943 (O_2943,N_27412,N_29977);
nor UO_2944 (O_2944,N_28418,N_28869);
or UO_2945 (O_2945,N_29986,N_28671);
nor UO_2946 (O_2946,N_28934,N_27252);
nor UO_2947 (O_2947,N_27700,N_27763);
xor UO_2948 (O_2948,N_27768,N_29600);
xor UO_2949 (O_2949,N_29453,N_27532);
xnor UO_2950 (O_2950,N_29677,N_29464);
and UO_2951 (O_2951,N_29897,N_28413);
or UO_2952 (O_2952,N_29570,N_28996);
nand UO_2953 (O_2953,N_29249,N_29688);
or UO_2954 (O_2954,N_28607,N_27518);
and UO_2955 (O_2955,N_27418,N_29220);
xnor UO_2956 (O_2956,N_27808,N_29991);
nand UO_2957 (O_2957,N_27769,N_28607);
nor UO_2958 (O_2958,N_27901,N_27075);
xnor UO_2959 (O_2959,N_27510,N_29232);
nor UO_2960 (O_2960,N_28470,N_28695);
nand UO_2961 (O_2961,N_27011,N_27077);
and UO_2962 (O_2962,N_27134,N_27017);
xor UO_2963 (O_2963,N_27294,N_28958);
nand UO_2964 (O_2964,N_27885,N_28315);
and UO_2965 (O_2965,N_27361,N_27675);
nand UO_2966 (O_2966,N_29747,N_28688);
xor UO_2967 (O_2967,N_29468,N_28542);
or UO_2968 (O_2968,N_29303,N_29198);
nor UO_2969 (O_2969,N_29369,N_28481);
and UO_2970 (O_2970,N_28244,N_28295);
xor UO_2971 (O_2971,N_28318,N_28047);
or UO_2972 (O_2972,N_28313,N_29204);
nand UO_2973 (O_2973,N_28771,N_27845);
xnor UO_2974 (O_2974,N_29305,N_28137);
or UO_2975 (O_2975,N_29681,N_29766);
or UO_2976 (O_2976,N_29605,N_28886);
and UO_2977 (O_2977,N_27794,N_29038);
and UO_2978 (O_2978,N_29493,N_27766);
and UO_2979 (O_2979,N_28752,N_27506);
xor UO_2980 (O_2980,N_28215,N_27244);
nor UO_2981 (O_2981,N_28968,N_27800);
nand UO_2982 (O_2982,N_27252,N_27296);
nand UO_2983 (O_2983,N_29590,N_28782);
or UO_2984 (O_2984,N_27523,N_27889);
nand UO_2985 (O_2985,N_27340,N_29589);
or UO_2986 (O_2986,N_28793,N_28761);
nand UO_2987 (O_2987,N_28881,N_29462);
or UO_2988 (O_2988,N_27570,N_27479);
xnor UO_2989 (O_2989,N_27883,N_27681);
and UO_2990 (O_2990,N_29756,N_29317);
nand UO_2991 (O_2991,N_27781,N_29354);
or UO_2992 (O_2992,N_29040,N_29824);
or UO_2993 (O_2993,N_29650,N_29352);
xnor UO_2994 (O_2994,N_28391,N_27586);
or UO_2995 (O_2995,N_28952,N_27085);
xnor UO_2996 (O_2996,N_28976,N_27399);
nand UO_2997 (O_2997,N_29582,N_28469);
nor UO_2998 (O_2998,N_28854,N_28306);
xnor UO_2999 (O_2999,N_27915,N_27041);
and UO_3000 (O_3000,N_29552,N_29254);
nor UO_3001 (O_3001,N_29441,N_29155);
nor UO_3002 (O_3002,N_27001,N_27922);
xnor UO_3003 (O_3003,N_27415,N_28464);
nand UO_3004 (O_3004,N_27295,N_28934);
xnor UO_3005 (O_3005,N_29256,N_28113);
xnor UO_3006 (O_3006,N_28140,N_27952);
xor UO_3007 (O_3007,N_27157,N_29333);
nor UO_3008 (O_3008,N_28354,N_27803);
nor UO_3009 (O_3009,N_29175,N_29240);
and UO_3010 (O_3010,N_29448,N_27185);
and UO_3011 (O_3011,N_27631,N_27543);
xor UO_3012 (O_3012,N_29961,N_27579);
nand UO_3013 (O_3013,N_28133,N_28005);
and UO_3014 (O_3014,N_29997,N_29728);
xor UO_3015 (O_3015,N_29656,N_28563);
or UO_3016 (O_3016,N_28966,N_27391);
and UO_3017 (O_3017,N_29111,N_28829);
and UO_3018 (O_3018,N_28142,N_29123);
nor UO_3019 (O_3019,N_27102,N_29141);
xor UO_3020 (O_3020,N_27810,N_27521);
xor UO_3021 (O_3021,N_28534,N_29167);
xnor UO_3022 (O_3022,N_29452,N_28596);
or UO_3023 (O_3023,N_29188,N_29973);
or UO_3024 (O_3024,N_28098,N_27552);
and UO_3025 (O_3025,N_27174,N_27486);
nor UO_3026 (O_3026,N_29823,N_28955);
or UO_3027 (O_3027,N_28223,N_28816);
or UO_3028 (O_3028,N_28539,N_27473);
and UO_3029 (O_3029,N_27164,N_27668);
nor UO_3030 (O_3030,N_28893,N_28509);
xnor UO_3031 (O_3031,N_29952,N_29309);
nor UO_3032 (O_3032,N_29448,N_27213);
xor UO_3033 (O_3033,N_29879,N_29842);
xor UO_3034 (O_3034,N_29283,N_27641);
and UO_3035 (O_3035,N_29048,N_28062);
or UO_3036 (O_3036,N_28890,N_28531);
and UO_3037 (O_3037,N_28736,N_28878);
xor UO_3038 (O_3038,N_27245,N_28811);
nand UO_3039 (O_3039,N_28862,N_29845);
and UO_3040 (O_3040,N_29004,N_27460);
nor UO_3041 (O_3041,N_29277,N_29748);
or UO_3042 (O_3042,N_29628,N_28876);
and UO_3043 (O_3043,N_27044,N_27754);
or UO_3044 (O_3044,N_28447,N_28047);
nand UO_3045 (O_3045,N_29635,N_28612);
or UO_3046 (O_3046,N_27676,N_29200);
or UO_3047 (O_3047,N_27852,N_27351);
and UO_3048 (O_3048,N_27667,N_27427);
xor UO_3049 (O_3049,N_27714,N_28957);
or UO_3050 (O_3050,N_29344,N_28430);
or UO_3051 (O_3051,N_27771,N_29466);
and UO_3052 (O_3052,N_29236,N_27906);
xnor UO_3053 (O_3053,N_29183,N_27095);
and UO_3054 (O_3054,N_29136,N_28588);
and UO_3055 (O_3055,N_29223,N_28661);
nand UO_3056 (O_3056,N_29261,N_27523);
and UO_3057 (O_3057,N_28256,N_27536);
nor UO_3058 (O_3058,N_29318,N_29545);
nand UO_3059 (O_3059,N_29923,N_27464);
nor UO_3060 (O_3060,N_27350,N_28846);
nor UO_3061 (O_3061,N_27300,N_29734);
xnor UO_3062 (O_3062,N_28852,N_29475);
nor UO_3063 (O_3063,N_27811,N_27594);
and UO_3064 (O_3064,N_28642,N_29460);
xnor UO_3065 (O_3065,N_28812,N_29290);
and UO_3066 (O_3066,N_28377,N_28757);
or UO_3067 (O_3067,N_29667,N_29725);
nand UO_3068 (O_3068,N_28672,N_29416);
nand UO_3069 (O_3069,N_29341,N_28407);
nand UO_3070 (O_3070,N_27293,N_28637);
and UO_3071 (O_3071,N_28010,N_28507);
nor UO_3072 (O_3072,N_29889,N_29384);
nand UO_3073 (O_3073,N_28920,N_28349);
nor UO_3074 (O_3074,N_27555,N_29883);
nand UO_3075 (O_3075,N_29920,N_28697);
nor UO_3076 (O_3076,N_29970,N_29230);
or UO_3077 (O_3077,N_28916,N_29106);
nand UO_3078 (O_3078,N_28081,N_27177);
and UO_3079 (O_3079,N_29085,N_27004);
xnor UO_3080 (O_3080,N_27546,N_28554);
nor UO_3081 (O_3081,N_27937,N_27572);
and UO_3082 (O_3082,N_27059,N_27840);
nand UO_3083 (O_3083,N_29391,N_29512);
nor UO_3084 (O_3084,N_29180,N_27625);
and UO_3085 (O_3085,N_28130,N_28451);
xor UO_3086 (O_3086,N_27336,N_29993);
and UO_3087 (O_3087,N_28406,N_27769);
xnor UO_3088 (O_3088,N_28183,N_27019);
nand UO_3089 (O_3089,N_27672,N_28491);
nor UO_3090 (O_3090,N_28423,N_29800);
or UO_3091 (O_3091,N_27871,N_28895);
xor UO_3092 (O_3092,N_28254,N_28725);
nor UO_3093 (O_3093,N_29665,N_27563);
nand UO_3094 (O_3094,N_28793,N_29427);
nor UO_3095 (O_3095,N_29833,N_29970);
or UO_3096 (O_3096,N_29777,N_29197);
and UO_3097 (O_3097,N_29428,N_29751);
nor UO_3098 (O_3098,N_28215,N_29401);
nand UO_3099 (O_3099,N_27210,N_29554);
or UO_3100 (O_3100,N_29512,N_29038);
nor UO_3101 (O_3101,N_27723,N_29221);
and UO_3102 (O_3102,N_28414,N_27910);
nor UO_3103 (O_3103,N_29146,N_28868);
nand UO_3104 (O_3104,N_27597,N_29603);
nor UO_3105 (O_3105,N_28464,N_28410);
nor UO_3106 (O_3106,N_28595,N_28352);
and UO_3107 (O_3107,N_27822,N_29042);
or UO_3108 (O_3108,N_27240,N_28540);
or UO_3109 (O_3109,N_28497,N_29147);
xor UO_3110 (O_3110,N_27127,N_29207);
and UO_3111 (O_3111,N_27756,N_28311);
nand UO_3112 (O_3112,N_29628,N_28795);
or UO_3113 (O_3113,N_27746,N_28545);
or UO_3114 (O_3114,N_28797,N_29463);
nor UO_3115 (O_3115,N_28498,N_28237);
or UO_3116 (O_3116,N_27623,N_29859);
xnor UO_3117 (O_3117,N_27569,N_29425);
and UO_3118 (O_3118,N_27235,N_28631);
xor UO_3119 (O_3119,N_28893,N_28951);
or UO_3120 (O_3120,N_28312,N_28608);
xnor UO_3121 (O_3121,N_29551,N_29791);
nand UO_3122 (O_3122,N_27480,N_27964);
and UO_3123 (O_3123,N_29388,N_27868);
and UO_3124 (O_3124,N_27826,N_27948);
or UO_3125 (O_3125,N_29303,N_28806);
and UO_3126 (O_3126,N_28700,N_27776);
or UO_3127 (O_3127,N_29336,N_28160);
and UO_3128 (O_3128,N_29258,N_28106);
and UO_3129 (O_3129,N_28877,N_29068);
nand UO_3130 (O_3130,N_29754,N_28915);
nor UO_3131 (O_3131,N_27679,N_29625);
xor UO_3132 (O_3132,N_29563,N_28256);
nor UO_3133 (O_3133,N_29995,N_29100);
nor UO_3134 (O_3134,N_29463,N_29633);
or UO_3135 (O_3135,N_28529,N_29482);
nand UO_3136 (O_3136,N_27124,N_28280);
and UO_3137 (O_3137,N_29139,N_27621);
nor UO_3138 (O_3138,N_28074,N_29273);
or UO_3139 (O_3139,N_29428,N_29734);
xor UO_3140 (O_3140,N_27392,N_27322);
nand UO_3141 (O_3141,N_27983,N_29743);
or UO_3142 (O_3142,N_27667,N_28871);
or UO_3143 (O_3143,N_27319,N_29615);
nand UO_3144 (O_3144,N_29391,N_29534);
xor UO_3145 (O_3145,N_27733,N_27861);
xnor UO_3146 (O_3146,N_27296,N_28736);
or UO_3147 (O_3147,N_27589,N_28500);
or UO_3148 (O_3148,N_29714,N_29737);
nand UO_3149 (O_3149,N_29357,N_28825);
or UO_3150 (O_3150,N_29225,N_29316);
nor UO_3151 (O_3151,N_29763,N_29638);
nor UO_3152 (O_3152,N_27341,N_27373);
xor UO_3153 (O_3153,N_29760,N_28836);
xnor UO_3154 (O_3154,N_28451,N_29044);
nor UO_3155 (O_3155,N_29972,N_27173);
nor UO_3156 (O_3156,N_28921,N_28102);
or UO_3157 (O_3157,N_28176,N_28092);
or UO_3158 (O_3158,N_29881,N_27102);
and UO_3159 (O_3159,N_28169,N_27036);
and UO_3160 (O_3160,N_28423,N_28428);
nand UO_3161 (O_3161,N_27533,N_27422);
nand UO_3162 (O_3162,N_28699,N_29715);
xnor UO_3163 (O_3163,N_27143,N_27387);
xnor UO_3164 (O_3164,N_29249,N_27217);
and UO_3165 (O_3165,N_27416,N_27519);
nor UO_3166 (O_3166,N_27160,N_28868);
and UO_3167 (O_3167,N_28709,N_28189);
and UO_3168 (O_3168,N_28791,N_29891);
xor UO_3169 (O_3169,N_27265,N_29557);
and UO_3170 (O_3170,N_28068,N_29553);
or UO_3171 (O_3171,N_29717,N_28741);
nand UO_3172 (O_3172,N_29727,N_28564);
nor UO_3173 (O_3173,N_29145,N_27857);
xor UO_3174 (O_3174,N_27622,N_29125);
or UO_3175 (O_3175,N_29674,N_29859);
or UO_3176 (O_3176,N_28789,N_27828);
nor UO_3177 (O_3177,N_28885,N_27047);
nor UO_3178 (O_3178,N_29128,N_27307);
and UO_3179 (O_3179,N_29662,N_28507);
or UO_3180 (O_3180,N_27420,N_29910);
nand UO_3181 (O_3181,N_28590,N_29133);
or UO_3182 (O_3182,N_28666,N_29955);
or UO_3183 (O_3183,N_28122,N_29818);
and UO_3184 (O_3184,N_27592,N_27259);
and UO_3185 (O_3185,N_29201,N_27764);
or UO_3186 (O_3186,N_29791,N_27929);
and UO_3187 (O_3187,N_28517,N_29425);
nor UO_3188 (O_3188,N_29242,N_27061);
and UO_3189 (O_3189,N_29864,N_27285);
xor UO_3190 (O_3190,N_27953,N_29308);
nand UO_3191 (O_3191,N_29765,N_29997);
or UO_3192 (O_3192,N_29446,N_29198);
and UO_3193 (O_3193,N_28411,N_27051);
nor UO_3194 (O_3194,N_27011,N_28389);
or UO_3195 (O_3195,N_28831,N_27889);
nand UO_3196 (O_3196,N_28966,N_29164);
xnor UO_3197 (O_3197,N_28746,N_27639);
and UO_3198 (O_3198,N_29576,N_28376);
xnor UO_3199 (O_3199,N_28789,N_28158);
nor UO_3200 (O_3200,N_27693,N_29779);
or UO_3201 (O_3201,N_27992,N_29321);
nand UO_3202 (O_3202,N_27660,N_29413);
nor UO_3203 (O_3203,N_29244,N_28206);
and UO_3204 (O_3204,N_27679,N_28907);
or UO_3205 (O_3205,N_29227,N_29986);
or UO_3206 (O_3206,N_29664,N_29060);
and UO_3207 (O_3207,N_28170,N_27055);
xor UO_3208 (O_3208,N_27435,N_27884);
or UO_3209 (O_3209,N_27099,N_28664);
and UO_3210 (O_3210,N_29702,N_27444);
nand UO_3211 (O_3211,N_27087,N_27332);
or UO_3212 (O_3212,N_27639,N_27941);
and UO_3213 (O_3213,N_27461,N_28387);
nor UO_3214 (O_3214,N_27421,N_27419);
or UO_3215 (O_3215,N_27888,N_28275);
and UO_3216 (O_3216,N_27554,N_27976);
nand UO_3217 (O_3217,N_28822,N_28310);
or UO_3218 (O_3218,N_27968,N_28171);
nor UO_3219 (O_3219,N_27347,N_27505);
and UO_3220 (O_3220,N_29607,N_28909);
or UO_3221 (O_3221,N_29944,N_27292);
nor UO_3222 (O_3222,N_29842,N_29890);
xor UO_3223 (O_3223,N_29370,N_29477);
or UO_3224 (O_3224,N_29397,N_29957);
or UO_3225 (O_3225,N_27151,N_27351);
nand UO_3226 (O_3226,N_29314,N_27394);
and UO_3227 (O_3227,N_29525,N_27935);
nand UO_3228 (O_3228,N_28350,N_27844);
xnor UO_3229 (O_3229,N_27752,N_29893);
xor UO_3230 (O_3230,N_29373,N_27773);
xor UO_3231 (O_3231,N_29402,N_29846);
nand UO_3232 (O_3232,N_27990,N_29889);
and UO_3233 (O_3233,N_28147,N_27049);
and UO_3234 (O_3234,N_29648,N_28017);
xnor UO_3235 (O_3235,N_28900,N_29846);
xor UO_3236 (O_3236,N_28765,N_27576);
and UO_3237 (O_3237,N_27791,N_27492);
nand UO_3238 (O_3238,N_27899,N_29283);
xnor UO_3239 (O_3239,N_28551,N_29344);
and UO_3240 (O_3240,N_27346,N_28541);
nor UO_3241 (O_3241,N_27550,N_29641);
and UO_3242 (O_3242,N_28609,N_29382);
xor UO_3243 (O_3243,N_27380,N_27240);
nand UO_3244 (O_3244,N_27694,N_27416);
xor UO_3245 (O_3245,N_28458,N_29128);
nor UO_3246 (O_3246,N_28165,N_29168);
xor UO_3247 (O_3247,N_27986,N_27928);
nor UO_3248 (O_3248,N_27386,N_27342);
and UO_3249 (O_3249,N_27832,N_29727);
nor UO_3250 (O_3250,N_28878,N_28714);
nand UO_3251 (O_3251,N_29400,N_29363);
nor UO_3252 (O_3252,N_27652,N_28919);
xor UO_3253 (O_3253,N_27850,N_28091);
or UO_3254 (O_3254,N_29009,N_29368);
nand UO_3255 (O_3255,N_28839,N_28043);
nand UO_3256 (O_3256,N_28364,N_29468);
nor UO_3257 (O_3257,N_29995,N_29831);
xor UO_3258 (O_3258,N_29310,N_29601);
nor UO_3259 (O_3259,N_28115,N_27539);
nor UO_3260 (O_3260,N_28282,N_28458);
nand UO_3261 (O_3261,N_27089,N_28040);
nor UO_3262 (O_3262,N_28742,N_29604);
or UO_3263 (O_3263,N_29204,N_28084);
or UO_3264 (O_3264,N_28268,N_28420);
nand UO_3265 (O_3265,N_28680,N_28752);
and UO_3266 (O_3266,N_27737,N_29600);
nor UO_3267 (O_3267,N_28725,N_29658);
or UO_3268 (O_3268,N_27968,N_29300);
and UO_3269 (O_3269,N_29186,N_28420);
nor UO_3270 (O_3270,N_29459,N_28078);
nand UO_3271 (O_3271,N_27981,N_27283);
or UO_3272 (O_3272,N_29927,N_28764);
nor UO_3273 (O_3273,N_28033,N_27346);
nand UO_3274 (O_3274,N_27752,N_27723);
nand UO_3275 (O_3275,N_27116,N_28979);
xnor UO_3276 (O_3276,N_27374,N_29411);
xnor UO_3277 (O_3277,N_29624,N_28807);
or UO_3278 (O_3278,N_29756,N_29464);
nor UO_3279 (O_3279,N_27215,N_28441);
nand UO_3280 (O_3280,N_27558,N_28171);
xor UO_3281 (O_3281,N_28002,N_29442);
xor UO_3282 (O_3282,N_29266,N_27765);
nand UO_3283 (O_3283,N_29597,N_29230);
xor UO_3284 (O_3284,N_27637,N_29563);
and UO_3285 (O_3285,N_28958,N_28428);
nand UO_3286 (O_3286,N_28030,N_27488);
nor UO_3287 (O_3287,N_28103,N_27202);
and UO_3288 (O_3288,N_27717,N_28954);
nor UO_3289 (O_3289,N_28477,N_28792);
nor UO_3290 (O_3290,N_29081,N_27803);
or UO_3291 (O_3291,N_29979,N_27249);
or UO_3292 (O_3292,N_27786,N_29145);
or UO_3293 (O_3293,N_27499,N_27305);
nand UO_3294 (O_3294,N_27307,N_28445);
and UO_3295 (O_3295,N_28593,N_28821);
nor UO_3296 (O_3296,N_27271,N_27758);
nand UO_3297 (O_3297,N_28082,N_28737);
and UO_3298 (O_3298,N_29801,N_27889);
xor UO_3299 (O_3299,N_29189,N_29112);
nand UO_3300 (O_3300,N_29460,N_29451);
or UO_3301 (O_3301,N_27169,N_29875);
nor UO_3302 (O_3302,N_29409,N_27526);
nor UO_3303 (O_3303,N_28626,N_29421);
nand UO_3304 (O_3304,N_29653,N_27647);
nand UO_3305 (O_3305,N_29132,N_28503);
xor UO_3306 (O_3306,N_27276,N_28513);
xnor UO_3307 (O_3307,N_27017,N_28250);
or UO_3308 (O_3308,N_27831,N_27046);
nor UO_3309 (O_3309,N_29398,N_29094);
xor UO_3310 (O_3310,N_27298,N_27359);
or UO_3311 (O_3311,N_27628,N_28209);
or UO_3312 (O_3312,N_27862,N_28520);
nand UO_3313 (O_3313,N_29358,N_29446);
or UO_3314 (O_3314,N_27633,N_27295);
or UO_3315 (O_3315,N_28572,N_28411);
xnor UO_3316 (O_3316,N_28165,N_29400);
nor UO_3317 (O_3317,N_27563,N_28708);
and UO_3318 (O_3318,N_29130,N_28797);
and UO_3319 (O_3319,N_29560,N_29745);
xor UO_3320 (O_3320,N_27582,N_27346);
nand UO_3321 (O_3321,N_27622,N_29917);
nor UO_3322 (O_3322,N_28199,N_28206);
and UO_3323 (O_3323,N_27554,N_27394);
or UO_3324 (O_3324,N_27548,N_27865);
or UO_3325 (O_3325,N_29016,N_28004);
nor UO_3326 (O_3326,N_29046,N_29570);
or UO_3327 (O_3327,N_27484,N_27913);
or UO_3328 (O_3328,N_28443,N_28536);
and UO_3329 (O_3329,N_29739,N_29889);
xnor UO_3330 (O_3330,N_27182,N_29927);
xnor UO_3331 (O_3331,N_28303,N_29675);
or UO_3332 (O_3332,N_27898,N_28219);
or UO_3333 (O_3333,N_28925,N_28843);
nand UO_3334 (O_3334,N_28512,N_27596);
and UO_3335 (O_3335,N_28395,N_28383);
or UO_3336 (O_3336,N_27476,N_29948);
nand UO_3337 (O_3337,N_28965,N_28100);
and UO_3338 (O_3338,N_28941,N_28930);
xor UO_3339 (O_3339,N_29960,N_27417);
and UO_3340 (O_3340,N_29701,N_29982);
nand UO_3341 (O_3341,N_28482,N_29414);
nor UO_3342 (O_3342,N_28151,N_28876);
or UO_3343 (O_3343,N_29667,N_28595);
or UO_3344 (O_3344,N_27161,N_28933);
nand UO_3345 (O_3345,N_28406,N_29889);
nand UO_3346 (O_3346,N_28175,N_27609);
and UO_3347 (O_3347,N_28327,N_27344);
nor UO_3348 (O_3348,N_27008,N_27049);
and UO_3349 (O_3349,N_27958,N_29638);
xor UO_3350 (O_3350,N_27277,N_28083);
xor UO_3351 (O_3351,N_27389,N_28769);
or UO_3352 (O_3352,N_27781,N_27703);
xor UO_3353 (O_3353,N_29028,N_28704);
nor UO_3354 (O_3354,N_28161,N_28180);
or UO_3355 (O_3355,N_29416,N_27289);
and UO_3356 (O_3356,N_27800,N_28397);
or UO_3357 (O_3357,N_28718,N_27959);
nor UO_3358 (O_3358,N_28938,N_27562);
nor UO_3359 (O_3359,N_28902,N_27974);
and UO_3360 (O_3360,N_27621,N_27007);
and UO_3361 (O_3361,N_27195,N_27640);
nand UO_3362 (O_3362,N_28152,N_29252);
xor UO_3363 (O_3363,N_28628,N_29189);
or UO_3364 (O_3364,N_27183,N_29473);
and UO_3365 (O_3365,N_28232,N_29141);
nand UO_3366 (O_3366,N_29190,N_27423);
nor UO_3367 (O_3367,N_27940,N_29838);
or UO_3368 (O_3368,N_27511,N_28339);
nand UO_3369 (O_3369,N_29058,N_27258);
xor UO_3370 (O_3370,N_28192,N_29861);
xnor UO_3371 (O_3371,N_27741,N_27885);
and UO_3372 (O_3372,N_27121,N_27093);
nor UO_3373 (O_3373,N_28340,N_29489);
or UO_3374 (O_3374,N_28642,N_27179);
nor UO_3375 (O_3375,N_29596,N_27701);
nand UO_3376 (O_3376,N_29854,N_28155);
xor UO_3377 (O_3377,N_28874,N_28522);
nand UO_3378 (O_3378,N_29848,N_29525);
nor UO_3379 (O_3379,N_29968,N_28156);
or UO_3380 (O_3380,N_28359,N_28844);
or UO_3381 (O_3381,N_27792,N_29615);
nor UO_3382 (O_3382,N_27454,N_28895);
nand UO_3383 (O_3383,N_29511,N_28072);
nand UO_3384 (O_3384,N_29081,N_29504);
or UO_3385 (O_3385,N_27026,N_29318);
nor UO_3386 (O_3386,N_28284,N_27148);
nor UO_3387 (O_3387,N_28655,N_27395);
or UO_3388 (O_3388,N_29514,N_28399);
nor UO_3389 (O_3389,N_29148,N_29950);
nor UO_3390 (O_3390,N_28619,N_28519);
nor UO_3391 (O_3391,N_28185,N_27628);
nand UO_3392 (O_3392,N_29893,N_29034);
or UO_3393 (O_3393,N_27767,N_27041);
xor UO_3394 (O_3394,N_29312,N_29088);
and UO_3395 (O_3395,N_29252,N_28996);
and UO_3396 (O_3396,N_27933,N_27458);
and UO_3397 (O_3397,N_28064,N_27036);
xnor UO_3398 (O_3398,N_27757,N_29452);
and UO_3399 (O_3399,N_29837,N_28527);
and UO_3400 (O_3400,N_28197,N_27310);
and UO_3401 (O_3401,N_27678,N_29930);
or UO_3402 (O_3402,N_27389,N_29477);
nor UO_3403 (O_3403,N_27675,N_29610);
or UO_3404 (O_3404,N_27815,N_28379);
or UO_3405 (O_3405,N_28738,N_27490);
nor UO_3406 (O_3406,N_28561,N_27021);
nand UO_3407 (O_3407,N_29870,N_27511);
nand UO_3408 (O_3408,N_28718,N_27495);
nand UO_3409 (O_3409,N_27322,N_28625);
and UO_3410 (O_3410,N_28154,N_27251);
nor UO_3411 (O_3411,N_29378,N_29198);
nand UO_3412 (O_3412,N_27327,N_28486);
nor UO_3413 (O_3413,N_27360,N_28861);
xnor UO_3414 (O_3414,N_27517,N_27972);
xnor UO_3415 (O_3415,N_27750,N_28236);
nand UO_3416 (O_3416,N_29780,N_27599);
or UO_3417 (O_3417,N_29303,N_28635);
and UO_3418 (O_3418,N_27693,N_27484);
or UO_3419 (O_3419,N_27221,N_27910);
or UO_3420 (O_3420,N_29983,N_29564);
xnor UO_3421 (O_3421,N_29515,N_28301);
nor UO_3422 (O_3422,N_28521,N_29227);
or UO_3423 (O_3423,N_29263,N_28287);
and UO_3424 (O_3424,N_29429,N_27453);
and UO_3425 (O_3425,N_27473,N_29983);
or UO_3426 (O_3426,N_29175,N_28643);
nand UO_3427 (O_3427,N_29123,N_28186);
and UO_3428 (O_3428,N_28684,N_27129);
xor UO_3429 (O_3429,N_27723,N_28682);
nand UO_3430 (O_3430,N_29881,N_29490);
or UO_3431 (O_3431,N_29067,N_27795);
or UO_3432 (O_3432,N_27365,N_27807);
and UO_3433 (O_3433,N_28467,N_28963);
nand UO_3434 (O_3434,N_27680,N_27765);
xnor UO_3435 (O_3435,N_29255,N_28885);
xnor UO_3436 (O_3436,N_28619,N_28852);
or UO_3437 (O_3437,N_27027,N_28659);
nor UO_3438 (O_3438,N_27336,N_27051);
nor UO_3439 (O_3439,N_27209,N_27527);
and UO_3440 (O_3440,N_27343,N_27902);
and UO_3441 (O_3441,N_29598,N_27297);
nor UO_3442 (O_3442,N_28435,N_28470);
and UO_3443 (O_3443,N_28898,N_28387);
nand UO_3444 (O_3444,N_28416,N_29900);
nand UO_3445 (O_3445,N_27908,N_27924);
xor UO_3446 (O_3446,N_27451,N_29444);
xnor UO_3447 (O_3447,N_29237,N_27483);
xor UO_3448 (O_3448,N_27315,N_27043);
xnor UO_3449 (O_3449,N_29925,N_27697);
xor UO_3450 (O_3450,N_27676,N_28899);
xnor UO_3451 (O_3451,N_29704,N_27569);
nand UO_3452 (O_3452,N_29392,N_29866);
nor UO_3453 (O_3453,N_27437,N_29085);
nor UO_3454 (O_3454,N_28726,N_28819);
xor UO_3455 (O_3455,N_29514,N_28681);
nand UO_3456 (O_3456,N_28233,N_29881);
or UO_3457 (O_3457,N_28232,N_27513);
nor UO_3458 (O_3458,N_29116,N_27018);
or UO_3459 (O_3459,N_27018,N_28836);
nand UO_3460 (O_3460,N_29048,N_27819);
nor UO_3461 (O_3461,N_29668,N_29486);
and UO_3462 (O_3462,N_28734,N_27343);
xnor UO_3463 (O_3463,N_27640,N_28970);
nand UO_3464 (O_3464,N_27158,N_27559);
nand UO_3465 (O_3465,N_29909,N_29863);
or UO_3466 (O_3466,N_27601,N_27091);
nor UO_3467 (O_3467,N_28180,N_29027);
xnor UO_3468 (O_3468,N_29129,N_28102);
and UO_3469 (O_3469,N_27558,N_28776);
nor UO_3470 (O_3470,N_27978,N_29375);
nor UO_3471 (O_3471,N_29475,N_27194);
xor UO_3472 (O_3472,N_27458,N_28518);
or UO_3473 (O_3473,N_29321,N_28004);
xnor UO_3474 (O_3474,N_27892,N_28720);
xor UO_3475 (O_3475,N_29362,N_28151);
nand UO_3476 (O_3476,N_29904,N_29086);
or UO_3477 (O_3477,N_27879,N_28938);
xor UO_3478 (O_3478,N_27556,N_27414);
nor UO_3479 (O_3479,N_28697,N_28848);
nand UO_3480 (O_3480,N_28636,N_27766);
nand UO_3481 (O_3481,N_27245,N_27668);
nor UO_3482 (O_3482,N_28217,N_27739);
nand UO_3483 (O_3483,N_27292,N_28504);
nand UO_3484 (O_3484,N_27019,N_28092);
nand UO_3485 (O_3485,N_28015,N_29444);
and UO_3486 (O_3486,N_27679,N_28787);
xor UO_3487 (O_3487,N_29690,N_28897);
nor UO_3488 (O_3488,N_27416,N_28091);
or UO_3489 (O_3489,N_29044,N_27610);
and UO_3490 (O_3490,N_28618,N_28688);
xnor UO_3491 (O_3491,N_27382,N_28306);
xor UO_3492 (O_3492,N_27955,N_29233);
xnor UO_3493 (O_3493,N_29842,N_27268);
nor UO_3494 (O_3494,N_29196,N_28486);
and UO_3495 (O_3495,N_28219,N_29299);
nand UO_3496 (O_3496,N_27259,N_29580);
nand UO_3497 (O_3497,N_28348,N_27021);
nand UO_3498 (O_3498,N_27951,N_27545);
nand UO_3499 (O_3499,N_29926,N_28856);
endmodule