module basic_1000_10000_1500_20_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_645,In_570);
nor U1 (N_1,In_956,In_963);
or U2 (N_2,In_143,In_420);
nor U3 (N_3,In_798,In_607);
and U4 (N_4,In_466,In_816);
nor U5 (N_5,In_111,In_532);
and U6 (N_6,In_692,In_26);
nand U7 (N_7,In_36,In_697);
nor U8 (N_8,In_272,In_819);
nor U9 (N_9,In_855,In_809);
xnor U10 (N_10,In_455,In_558);
nor U11 (N_11,In_635,In_28);
and U12 (N_12,In_857,In_306);
and U13 (N_13,In_503,In_741);
or U14 (N_14,In_142,In_467);
nor U15 (N_15,In_8,In_890);
xor U16 (N_16,In_648,In_281);
xor U17 (N_17,In_96,In_61);
and U18 (N_18,In_110,In_826);
nand U19 (N_19,In_266,In_247);
xnor U20 (N_20,In_109,In_719);
nand U21 (N_21,In_204,In_943);
nor U22 (N_22,In_847,In_858);
and U23 (N_23,In_773,In_497);
and U24 (N_24,In_267,In_854);
nand U25 (N_25,In_241,In_401);
nand U26 (N_26,In_338,In_477);
and U27 (N_27,In_377,In_438);
and U28 (N_28,In_829,In_3);
xor U29 (N_29,In_929,In_418);
nor U30 (N_30,In_67,In_407);
and U31 (N_31,In_223,In_846);
and U32 (N_32,In_45,In_25);
nand U33 (N_33,In_140,In_557);
nor U34 (N_34,In_485,In_865);
nand U35 (N_35,In_150,In_804);
xnor U36 (N_36,In_52,In_629);
nand U37 (N_37,In_810,In_969);
xnor U38 (N_38,In_293,In_90);
or U39 (N_39,In_422,In_275);
and U40 (N_40,In_434,In_270);
or U41 (N_41,In_585,In_440);
xnor U42 (N_42,In_118,In_861);
or U43 (N_43,In_235,In_173);
xor U44 (N_44,In_144,In_791);
and U45 (N_45,In_850,In_313);
or U46 (N_46,In_742,In_716);
xor U47 (N_47,In_533,In_482);
or U48 (N_48,In_748,In_547);
and U49 (N_49,In_868,In_788);
xnor U50 (N_50,In_638,In_172);
xnor U51 (N_51,In_454,In_577);
nand U52 (N_52,In_331,In_531);
nand U53 (N_53,In_789,In_179);
and U54 (N_54,In_326,In_470);
nand U55 (N_55,In_351,In_588);
or U56 (N_56,In_794,In_991);
and U57 (N_57,In_189,In_350);
or U58 (N_58,In_589,In_955);
or U59 (N_59,In_93,In_34);
or U60 (N_60,In_750,In_537);
or U61 (N_61,In_184,In_764);
xor U62 (N_62,In_199,In_888);
xnor U63 (N_63,In_807,In_982);
xor U64 (N_64,In_453,In_727);
or U65 (N_65,In_170,In_708);
xnor U66 (N_66,In_433,In_0);
and U67 (N_67,In_29,In_898);
nand U68 (N_68,In_516,In_641);
xor U69 (N_69,In_812,In_30);
and U70 (N_70,In_835,In_479);
or U71 (N_71,In_785,In_971);
or U72 (N_72,In_555,In_592);
and U73 (N_73,In_112,In_990);
nand U74 (N_74,In_928,In_302);
or U75 (N_75,In_177,In_817);
nand U76 (N_76,In_691,In_653);
nor U77 (N_77,In_540,In_889);
nor U78 (N_78,In_800,In_566);
nand U79 (N_79,In_584,In_445);
or U80 (N_80,In_435,In_511);
nand U81 (N_81,In_625,In_209);
nand U82 (N_82,In_538,In_125);
nor U83 (N_83,In_852,In_21);
xnor U84 (N_84,In_354,In_450);
nand U85 (N_85,In_859,In_745);
and U86 (N_86,In_2,In_891);
xor U87 (N_87,In_755,In_392);
and U88 (N_88,In_406,In_149);
nor U89 (N_89,In_40,In_178);
nor U90 (N_90,In_233,In_280);
or U91 (N_91,In_341,In_636);
nor U92 (N_92,In_135,In_662);
or U93 (N_93,In_722,In_752);
xnor U94 (N_94,In_552,In_926);
xor U95 (N_95,In_290,In_307);
and U96 (N_96,In_333,In_160);
or U97 (N_97,In_996,In_604);
and U98 (N_98,In_480,In_318);
nand U99 (N_99,In_133,In_843);
xor U100 (N_100,In_549,In_188);
nand U101 (N_101,In_740,In_167);
xnor U102 (N_102,In_907,In_66);
nand U103 (N_103,In_805,In_811);
xor U104 (N_104,In_53,In_766);
xnor U105 (N_105,In_521,In_565);
and U106 (N_106,In_681,In_217);
xnor U107 (N_107,In_893,In_360);
nand U108 (N_108,In_660,In_601);
nor U109 (N_109,In_289,In_141);
nor U110 (N_110,In_298,In_175);
and U111 (N_111,In_371,In_376);
or U112 (N_112,In_504,In_905);
nor U113 (N_113,In_803,In_491);
xnor U114 (N_114,In_612,In_201);
nor U115 (N_115,In_978,In_117);
nand U116 (N_116,In_337,In_763);
and U117 (N_117,In_542,In_787);
xnor U118 (N_118,In_922,In_654);
nor U119 (N_119,In_702,In_862);
nand U120 (N_120,In_352,In_760);
or U121 (N_121,In_502,In_632);
xor U122 (N_122,In_572,In_389);
or U123 (N_123,In_359,In_863);
and U124 (N_124,In_610,In_821);
or U125 (N_125,In_122,In_545);
or U126 (N_126,In_658,In_953);
nand U127 (N_127,In_238,In_820);
nor U128 (N_128,In_134,In_769);
nor U129 (N_129,In_487,In_501);
xnor U130 (N_130,In_683,In_739);
or U131 (N_131,In_698,In_119);
nand U132 (N_132,In_291,In_274);
and U133 (N_133,In_630,In_33);
or U134 (N_134,In_534,In_260);
and U135 (N_135,In_14,In_417);
nand U136 (N_136,In_792,In_108);
and U137 (N_137,In_77,In_931);
xnor U138 (N_138,In_573,In_265);
and U139 (N_139,In_263,In_101);
or U140 (N_140,In_496,In_967);
nor U141 (N_141,In_513,In_159);
nor U142 (N_142,In_357,In_365);
xor U143 (N_143,In_631,In_308);
and U144 (N_144,In_17,In_469);
nand U145 (N_145,In_675,In_367);
and U146 (N_146,In_616,In_330);
and U147 (N_147,In_876,In_378);
and U148 (N_148,In_368,In_79);
nor U149 (N_149,In_590,In_320);
nand U150 (N_150,In_124,In_403);
xor U151 (N_151,In_309,In_214);
and U152 (N_152,In_700,In_47);
xor U153 (N_153,In_448,In_102);
nor U154 (N_154,In_32,In_414);
nor U155 (N_155,In_806,In_346);
nor U156 (N_156,In_15,In_598);
nor U157 (N_157,In_129,In_743);
nand U158 (N_158,In_737,In_814);
nor U159 (N_159,In_866,In_24);
and U160 (N_160,In_193,In_622);
nand U161 (N_161,In_459,In_85);
nor U162 (N_162,In_163,In_429);
or U163 (N_163,In_801,In_959);
or U164 (N_164,In_576,In_99);
and U165 (N_165,In_57,In_373);
nor U166 (N_166,In_180,In_7);
xnor U167 (N_167,In_297,In_424);
and U168 (N_168,In_222,In_947);
xor U169 (N_169,In_451,In_278);
or U170 (N_170,In_884,In_878);
xnor U171 (N_171,In_825,In_156);
or U172 (N_172,In_239,In_923);
and U173 (N_173,In_851,In_896);
nor U174 (N_174,In_419,In_619);
and U175 (N_175,In_594,In_568);
or U176 (N_176,In_65,In_439);
and U177 (N_177,In_164,In_191);
and U178 (N_178,In_918,In_190);
nand U179 (N_179,In_628,In_674);
and U180 (N_180,In_603,In_867);
nor U181 (N_181,In_121,In_582);
xor U182 (N_182,In_657,In_892);
xnor U183 (N_183,In_725,In_345);
and U184 (N_184,In_215,In_839);
xor U185 (N_185,In_31,In_949);
xor U186 (N_186,In_325,In_687);
nand U187 (N_187,In_751,In_207);
and U188 (N_188,In_95,In_966);
or U189 (N_189,In_633,In_883);
nor U190 (N_190,In_200,In_994);
nand U191 (N_191,In_961,In_767);
and U192 (N_192,In_525,In_828);
xnor U193 (N_193,In_372,In_489);
or U194 (N_194,In_508,In_818);
and U195 (N_195,In_369,In_637);
nor U196 (N_196,In_962,In_518);
xnor U197 (N_197,In_837,In_211);
nand U198 (N_198,In_317,In_836);
and U199 (N_199,In_483,In_759);
nor U200 (N_200,In_347,In_988);
nor U201 (N_201,In_758,In_913);
and U202 (N_202,In_286,In_600);
or U203 (N_203,In_87,In_490);
xor U204 (N_204,In_714,In_19);
xnor U205 (N_205,In_877,In_186);
and U206 (N_206,In_264,In_208);
and U207 (N_207,In_986,In_909);
or U208 (N_208,In_205,In_639);
nand U209 (N_209,In_860,In_546);
nand U210 (N_210,In_493,In_35);
and U211 (N_211,In_395,In_526);
and U212 (N_212,In_492,In_20);
nand U213 (N_213,In_405,In_409);
and U214 (N_214,In_279,In_746);
nand U215 (N_215,In_228,In_663);
nor U216 (N_216,In_599,In_756);
nor U217 (N_217,In_37,In_224);
and U218 (N_218,In_246,In_106);
and U219 (N_219,In_778,In_509);
xnor U220 (N_220,In_244,In_145);
or U221 (N_221,In_390,In_919);
or U222 (N_222,In_981,In_822);
nand U223 (N_223,In_22,In_784);
nor U224 (N_224,In_428,In_216);
xor U225 (N_225,In_212,In_56);
or U226 (N_226,In_734,In_523);
and U227 (N_227,In_54,In_271);
xnor U228 (N_228,In_934,In_673);
or U229 (N_229,In_296,In_132);
nor U230 (N_230,In_171,In_647);
xnor U231 (N_231,In_69,In_382);
and U232 (N_232,In_495,In_668);
nand U233 (N_233,In_431,In_882);
and U234 (N_234,In_586,In_176);
xnor U235 (N_235,In_795,In_258);
nor U236 (N_236,In_569,In_203);
xnor U237 (N_237,In_997,In_255);
or U238 (N_238,In_738,In_355);
and U239 (N_239,In_220,In_664);
or U240 (N_240,In_519,In_358);
nor U241 (N_241,In_301,In_973);
nand U242 (N_242,In_476,In_617);
or U243 (N_243,In_925,In_42);
or U244 (N_244,In_362,In_813);
and U245 (N_245,In_575,In_234);
and U246 (N_246,In_294,In_624);
xor U247 (N_247,In_833,In_951);
nor U248 (N_248,In_609,In_520);
and U249 (N_249,In_977,In_253);
xnor U250 (N_250,In_940,In_946);
nand U251 (N_251,In_456,In_452);
and U252 (N_252,In_960,In_396);
xnor U253 (N_253,In_731,In_128);
and U254 (N_254,In_213,In_786);
or U255 (N_255,In_535,In_507);
and U256 (N_256,In_46,In_62);
nand U257 (N_257,In_443,In_917);
nand U258 (N_258,In_985,In_989);
nand U259 (N_259,In_304,In_374);
nand U260 (N_260,In_793,In_524);
nor U261 (N_261,In_38,In_334);
xnor U262 (N_262,In_364,In_688);
nor U263 (N_263,In_621,In_70);
nand U264 (N_264,In_416,In_561);
xor U265 (N_265,In_656,In_104);
or U266 (N_266,In_9,In_644);
nand U267 (N_267,In_464,In_18);
or U268 (N_268,In_75,In_623);
or U269 (N_269,In_375,In_174);
or U270 (N_270,In_285,In_669);
nor U271 (N_271,In_83,In_232);
xnor U272 (N_272,In_721,In_505);
nor U273 (N_273,In_754,In_328);
or U274 (N_274,In_157,In_383);
and U275 (N_275,In_718,In_486);
nor U276 (N_276,In_897,In_463);
nor U277 (N_277,In_185,In_126);
and U278 (N_278,In_845,In_356);
xor U279 (N_279,In_903,In_181);
xor U280 (N_280,In_541,In_659);
and U281 (N_281,In_939,In_147);
or U282 (N_282,In_136,In_689);
and U283 (N_283,In_72,In_321);
nand U284 (N_284,In_765,In_120);
and U285 (N_285,In_51,In_363);
nor U286 (N_286,In_370,In_55);
and U287 (N_287,In_197,In_643);
xnor U288 (N_288,In_980,In_71);
nor U289 (N_289,In_640,In_595);
and U290 (N_290,In_735,In_472);
xnor U291 (N_291,In_299,In_89);
or U292 (N_292,In_684,In_642);
or U293 (N_293,In_723,In_465);
and U294 (N_294,In_76,In_550);
and U295 (N_295,In_578,In_544);
and U296 (N_296,In_522,In_536);
nand U297 (N_297,In_701,In_914);
xnor U298 (N_298,In_169,In_327);
nand U299 (N_299,In_999,In_696);
nor U300 (N_300,In_484,In_975);
nand U301 (N_301,In_710,In_153);
nand U302 (N_302,In_968,In_548);
nor U303 (N_303,In_895,In_444);
xor U304 (N_304,In_393,In_225);
nor U305 (N_305,In_100,In_500);
or U306 (N_306,In_394,In_693);
or U307 (N_307,In_924,In_732);
nor U308 (N_308,In_336,In_59);
xor U309 (N_309,In_768,In_43);
and U310 (N_310,In_243,In_98);
nand U311 (N_311,In_802,In_945);
or U312 (N_312,In_256,In_904);
nand U313 (N_313,In_626,In_387);
xor U314 (N_314,In_605,In_938);
nand U315 (N_315,In_676,In_881);
nand U316 (N_316,In_580,In_342);
or U317 (N_317,In_4,In_815);
and U318 (N_318,In_781,In_952);
or U319 (N_319,In_724,In_761);
nor U320 (N_320,In_316,In_747);
or U321 (N_321,In_48,In_397);
xor U322 (N_322,In_499,In_155);
and U323 (N_323,In_348,In_388);
nand U324 (N_324,In_615,In_166);
and U325 (N_325,In_699,In_944);
nand U326 (N_326,In_161,In_554);
xor U327 (N_327,In_97,In_183);
xor U328 (N_328,In_221,In_12);
xnor U329 (N_329,In_950,In_887);
nor U330 (N_330,In_844,In_86);
and U331 (N_331,In_634,In_425);
nand U332 (N_332,In_332,In_709);
and U333 (N_333,In_983,In_249);
nand U334 (N_334,In_283,In_335);
xor U335 (N_335,In_105,In_620);
and U336 (N_336,In_958,In_252);
nand U337 (N_337,In_974,In_921);
and U338 (N_338,In_475,In_842);
or U339 (N_339,In_678,In_206);
or U340 (N_340,In_81,In_230);
or U341 (N_341,In_563,In_10);
nand U342 (N_342,In_310,In_799);
nand U343 (N_343,In_712,In_685);
xor U344 (N_344,In_560,In_339);
nand U345 (N_345,In_972,In_257);
or U346 (N_346,In_941,In_899);
and U347 (N_347,In_58,In_717);
nand U348 (N_348,In_840,In_80);
xor U349 (N_349,In_268,In_273);
nor U350 (N_350,In_82,In_408);
or U351 (N_351,In_1,In_384);
or U352 (N_352,In_911,In_611);
xor U353 (N_353,In_462,In_984);
or U354 (N_354,In_666,In_529);
or U355 (N_355,In_386,In_195);
nor U356 (N_356,In_192,In_131);
xnor U357 (N_357,In_449,In_282);
nand U358 (N_358,In_562,In_736);
nand U359 (N_359,In_261,In_303);
or U360 (N_360,In_421,In_458);
xnor U361 (N_361,In_970,In_682);
nor U362 (N_362,In_694,In_730);
nand U363 (N_363,In_777,In_312);
nand U364 (N_364,In_830,In_571);
nor U365 (N_365,In_194,In_661);
or U366 (N_366,In_385,In_63);
xnor U367 (N_367,In_680,In_726);
and U368 (N_368,In_391,In_775);
xnor U369 (N_369,In_436,In_979);
or U370 (N_370,In_665,In_579);
or U371 (N_371,In_468,In_652);
nand U372 (N_372,In_749,In_530);
xor U373 (N_373,In_906,In_872);
nand U374 (N_374,In_103,In_292);
or U375 (N_375,In_114,In_935);
nand U376 (N_376,In_942,In_885);
and U377 (N_377,In_993,In_441);
xnor U378 (N_378,In_300,In_932);
or U379 (N_379,In_92,In_413);
xor U380 (N_380,In_430,In_559);
xnor U381 (N_381,In_227,In_553);
nand U382 (N_382,In_510,In_670);
or U383 (N_383,In_690,In_276);
or U384 (N_384,In_324,In_410);
or U385 (N_385,In_123,In_728);
or U386 (N_386,In_231,In_488);
nand U387 (N_387,In_139,In_138);
or U388 (N_388,In_782,In_920);
xnor U389 (N_389,In_936,In_720);
or U390 (N_390,In_853,In_457);
and U391 (N_391,In_762,In_528);
xor U392 (N_392,In_707,In_50);
nand U393 (N_393,In_277,In_729);
nor U394 (N_394,In_912,In_672);
nor U395 (N_395,In_987,In_380);
xor U396 (N_396,In_832,In_770);
nor U397 (N_397,In_733,In_11);
xor U398 (N_398,In_992,In_415);
nand U399 (N_399,In_74,In_242);
or U400 (N_400,In_886,In_606);
or U401 (N_401,In_695,In_262);
nand U402 (N_402,In_27,In_116);
or U403 (N_403,In_824,In_871);
nand U404 (N_404,In_73,In_827);
nand U405 (N_405,In_165,In_158);
xor U406 (N_406,In_776,In_869);
nor U407 (N_407,In_796,In_649);
nor U408 (N_408,In_219,In_514);
nand U409 (N_409,In_329,In_442);
and U410 (N_410,In_667,In_686);
or U411 (N_411,In_948,In_976);
xor U412 (N_412,In_774,In_915);
nor U413 (N_413,In_259,In_130);
nor U414 (N_414,In_91,In_583);
nand U415 (N_415,In_127,In_398);
nor U416 (N_416,In_711,In_790);
and U417 (N_417,In_902,In_597);
or U418 (N_418,In_848,In_864);
or U419 (N_419,In_284,In_596);
nand U420 (N_420,In_427,In_437);
nor U421 (N_421,In_68,In_44);
xor U422 (N_422,In_248,In_875);
nand U423 (N_423,In_744,In_6);
nand U424 (N_424,In_927,In_152);
nor U425 (N_425,In_808,In_295);
and U426 (N_426,In_361,In_340);
nand U427 (N_427,In_527,In_198);
xor U428 (N_428,In_957,In_107);
and U429 (N_429,In_411,In_512);
xor U430 (N_430,In_581,In_366);
xnor U431 (N_431,In_646,In_49);
nand U432 (N_432,In_677,In_353);
xor U433 (N_433,In_551,In_315);
or U434 (N_434,In_94,In_323);
nand U435 (N_435,In_461,In_753);
nor U436 (N_436,In_13,In_506);
xnor U437 (N_437,In_608,In_471);
xnor U438 (N_438,In_314,In_930);
nor U439 (N_439,In_704,In_446);
nor U440 (N_440,In_916,In_515);
nand U441 (N_441,In_494,In_182);
or U442 (N_442,In_287,In_757);
xnor U443 (N_443,In_910,In_154);
and U444 (N_444,In_771,In_556);
and U445 (N_445,In_933,In_478);
xor U446 (N_446,In_474,In_226);
or U447 (N_447,In_162,In_779);
or U448 (N_448,In_113,In_894);
xnor U449 (N_449,In_78,In_870);
or U450 (N_450,In_627,In_237);
or U451 (N_451,In_856,In_146);
nand U452 (N_452,In_473,In_254);
nand U453 (N_453,In_481,In_564);
xnor U454 (N_454,In_16,In_196);
or U455 (N_455,In_849,In_995);
xor U456 (N_456,In_879,In_671);
nand U457 (N_457,In_60,In_236);
nand U458 (N_458,In_618,In_715);
nor U459 (N_459,In_202,In_432);
or U460 (N_460,In_5,In_210);
nand U461 (N_461,In_498,In_901);
and U462 (N_462,In_651,In_965);
and U463 (N_463,In_954,In_305);
or U464 (N_464,In_288,In_650);
nand U465 (N_465,In_831,In_88);
nor U466 (N_466,In_269,In_311);
and U467 (N_467,In_187,In_229);
and U468 (N_468,In_381,In_998);
and U469 (N_469,In_322,In_613);
nor U470 (N_470,In_343,In_41);
or U471 (N_471,In_614,In_703);
xor U472 (N_472,In_655,In_908);
xor U473 (N_473,In_148,In_151);
nor U474 (N_474,In_834,In_64);
and U475 (N_475,In_602,In_245);
or U476 (N_476,In_460,In_823);
or U477 (N_477,In_783,In_402);
nor U478 (N_478,In_517,In_873);
xnor U479 (N_479,In_344,In_39);
nor U480 (N_480,In_880,In_349);
xor U481 (N_481,In_23,In_567);
and U482 (N_482,In_964,In_772);
or U483 (N_483,In_713,In_838);
or U484 (N_484,In_780,In_115);
nand U485 (N_485,In_218,In_447);
nand U486 (N_486,In_539,In_250);
and U487 (N_487,In_423,In_137);
or U488 (N_488,In_543,In_168);
or U489 (N_489,In_574,In_84);
or U490 (N_490,In_706,In_412);
or U491 (N_491,In_797,In_591);
and U492 (N_492,In_679,In_593);
nand U493 (N_493,In_251,In_240);
nor U494 (N_494,In_937,In_900);
nor U495 (N_495,In_705,In_426);
nor U496 (N_496,In_319,In_399);
xor U497 (N_497,In_404,In_400);
nand U498 (N_498,In_874,In_379);
xnor U499 (N_499,In_841,In_587);
nor U500 (N_500,N_54,N_10);
xnor U501 (N_501,N_232,N_304);
nor U502 (N_502,N_270,N_447);
nand U503 (N_503,N_34,N_95);
xor U504 (N_504,N_303,N_285);
or U505 (N_505,N_231,N_222);
xnor U506 (N_506,N_496,N_56);
or U507 (N_507,N_280,N_476);
nand U508 (N_508,N_217,N_373);
and U509 (N_509,N_173,N_300);
nor U510 (N_510,N_174,N_269);
nor U511 (N_511,N_310,N_256);
xnor U512 (N_512,N_37,N_474);
or U513 (N_513,N_203,N_435);
xnor U514 (N_514,N_359,N_378);
nand U515 (N_515,N_151,N_130);
and U516 (N_516,N_277,N_339);
xnor U517 (N_517,N_49,N_175);
nor U518 (N_518,N_164,N_387);
or U519 (N_519,N_40,N_115);
or U520 (N_520,N_448,N_273);
nand U521 (N_521,N_463,N_478);
nor U522 (N_522,N_464,N_453);
nor U523 (N_523,N_267,N_0);
xor U524 (N_524,N_262,N_155);
or U525 (N_525,N_237,N_185);
and U526 (N_526,N_168,N_230);
or U527 (N_527,N_132,N_67);
nor U528 (N_528,N_128,N_441);
and U529 (N_529,N_176,N_398);
and U530 (N_530,N_278,N_64);
xor U531 (N_531,N_197,N_473);
xnor U532 (N_532,N_77,N_47);
nand U533 (N_533,N_187,N_61);
or U534 (N_534,N_485,N_499);
nand U535 (N_535,N_106,N_451);
and U536 (N_536,N_389,N_434);
and U537 (N_537,N_253,N_201);
xor U538 (N_538,N_309,N_32);
or U539 (N_539,N_320,N_140);
or U540 (N_540,N_318,N_268);
or U541 (N_541,N_419,N_177);
xnor U542 (N_542,N_78,N_317);
or U543 (N_543,N_383,N_439);
nand U544 (N_544,N_401,N_257);
xor U545 (N_545,N_417,N_13);
or U546 (N_546,N_274,N_471);
nand U547 (N_547,N_199,N_143);
xor U548 (N_548,N_433,N_316);
nor U549 (N_549,N_314,N_420);
nand U550 (N_550,N_481,N_497);
and U551 (N_551,N_251,N_18);
nor U552 (N_552,N_369,N_412);
and U553 (N_553,N_319,N_264);
and U554 (N_554,N_206,N_361);
nor U555 (N_555,N_281,N_357);
nand U556 (N_556,N_221,N_353);
or U557 (N_557,N_109,N_223);
nor U558 (N_558,N_313,N_9);
and U559 (N_559,N_252,N_89);
or U560 (N_560,N_301,N_290);
and U561 (N_561,N_427,N_272);
nand U562 (N_562,N_355,N_395);
nor U563 (N_563,N_408,N_430);
nor U564 (N_564,N_422,N_402);
nor U565 (N_565,N_102,N_79);
or U566 (N_566,N_114,N_338);
and U567 (N_567,N_17,N_487);
and U568 (N_568,N_495,N_41);
nor U569 (N_569,N_216,N_215);
xor U570 (N_570,N_350,N_432);
nor U571 (N_571,N_135,N_124);
and U572 (N_572,N_169,N_324);
nor U573 (N_573,N_162,N_120);
nor U574 (N_574,N_195,N_72);
or U575 (N_575,N_43,N_352);
or U576 (N_576,N_295,N_263);
or U577 (N_577,N_287,N_38);
xor U578 (N_578,N_351,N_92);
nand U579 (N_579,N_336,N_327);
nand U580 (N_580,N_15,N_85);
nand U581 (N_581,N_192,N_414);
nor U582 (N_582,N_400,N_189);
xnor U583 (N_583,N_12,N_259);
xnor U584 (N_584,N_91,N_181);
nor U585 (N_585,N_191,N_161);
nand U586 (N_586,N_328,N_71);
xnor U587 (N_587,N_340,N_292);
nor U588 (N_588,N_362,N_19);
nor U589 (N_589,N_103,N_406);
nor U590 (N_590,N_153,N_8);
and U591 (N_591,N_90,N_243);
xnor U592 (N_592,N_229,N_475);
xnor U593 (N_593,N_51,N_358);
nor U594 (N_594,N_394,N_105);
nor U595 (N_595,N_171,N_219);
and U596 (N_596,N_126,N_299);
nor U597 (N_597,N_421,N_341);
nand U598 (N_598,N_489,N_65);
or U599 (N_599,N_266,N_202);
and U600 (N_600,N_163,N_225);
and U601 (N_601,N_138,N_329);
xor U602 (N_602,N_183,N_84);
or U603 (N_603,N_344,N_214);
nor U604 (N_604,N_70,N_3);
and U605 (N_605,N_184,N_97);
or U606 (N_606,N_288,N_148);
nand U607 (N_607,N_226,N_388);
and U608 (N_608,N_375,N_110);
xnor U609 (N_609,N_438,N_348);
or U610 (N_610,N_261,N_27);
or U611 (N_611,N_112,N_470);
or U612 (N_612,N_127,N_330);
nand U613 (N_613,N_467,N_296);
xnor U614 (N_614,N_454,N_59);
xnor U615 (N_615,N_254,N_25);
and U616 (N_616,N_260,N_53);
xor U617 (N_617,N_149,N_384);
or U618 (N_618,N_74,N_460);
and U619 (N_619,N_456,N_436);
and U620 (N_620,N_240,N_431);
xnor U621 (N_621,N_6,N_407);
nand U622 (N_622,N_486,N_233);
nor U623 (N_623,N_179,N_276);
nor U624 (N_624,N_68,N_147);
or U625 (N_625,N_386,N_356);
xor U626 (N_626,N_322,N_404);
and U627 (N_627,N_425,N_14);
xor U628 (N_628,N_469,N_413);
nand U629 (N_629,N_354,N_134);
xnor U630 (N_630,N_492,N_1);
and U631 (N_631,N_24,N_363);
xnor U632 (N_632,N_465,N_190);
xor U633 (N_633,N_411,N_33);
nor U634 (N_634,N_241,N_152);
nor U635 (N_635,N_144,N_298);
xnor U636 (N_636,N_154,N_5);
nor U637 (N_637,N_236,N_283);
nand U638 (N_638,N_380,N_347);
xnor U639 (N_639,N_325,N_100);
nand U640 (N_640,N_426,N_212);
or U641 (N_641,N_58,N_36);
and U642 (N_642,N_117,N_409);
or U643 (N_643,N_391,N_377);
nand U644 (N_644,N_160,N_121);
nor U645 (N_645,N_20,N_31);
xor U646 (N_646,N_477,N_484);
and U647 (N_647,N_326,N_423);
or U648 (N_648,N_119,N_480);
and U649 (N_649,N_131,N_87);
nor U650 (N_650,N_246,N_382);
and U651 (N_651,N_157,N_452);
xor U652 (N_652,N_145,N_86);
or U653 (N_653,N_76,N_113);
or U654 (N_654,N_118,N_200);
nand U655 (N_655,N_4,N_186);
and U656 (N_656,N_99,N_392);
nand U657 (N_657,N_188,N_137);
nor U658 (N_658,N_218,N_7);
or U659 (N_659,N_493,N_374);
and U660 (N_660,N_337,N_286);
and U661 (N_661,N_293,N_123);
or U662 (N_662,N_156,N_282);
nor U663 (N_663,N_42,N_482);
nor U664 (N_664,N_224,N_372);
xnor U665 (N_665,N_444,N_104);
xnor U666 (N_666,N_133,N_258);
or U667 (N_667,N_416,N_129);
nand U668 (N_668,N_122,N_141);
nand U669 (N_669,N_498,N_365);
nand U670 (N_670,N_483,N_405);
or U671 (N_671,N_111,N_196);
and U672 (N_672,N_159,N_468);
or U673 (N_673,N_52,N_440);
xnor U674 (N_674,N_312,N_88);
xor U675 (N_675,N_331,N_307);
or U676 (N_676,N_250,N_393);
nand U677 (N_677,N_349,N_210);
xor U678 (N_678,N_445,N_239);
and U679 (N_679,N_23,N_442);
nand U680 (N_680,N_472,N_379);
nand U681 (N_681,N_93,N_30);
nand U682 (N_682,N_390,N_205);
nand U683 (N_683,N_82,N_165);
nor U684 (N_684,N_342,N_302);
nand U685 (N_685,N_207,N_234);
or U686 (N_686,N_69,N_385);
or U687 (N_687,N_443,N_167);
or U688 (N_688,N_248,N_98);
or U689 (N_689,N_194,N_305);
or U690 (N_690,N_466,N_242);
nand U691 (N_691,N_166,N_2);
or U692 (N_692,N_308,N_381);
nand U693 (N_693,N_494,N_94);
or U694 (N_694,N_22,N_360);
or U695 (N_695,N_415,N_345);
or U696 (N_696,N_57,N_29);
nand U697 (N_697,N_139,N_399);
nand U698 (N_698,N_335,N_458);
xnor U699 (N_699,N_368,N_450);
xnor U700 (N_700,N_315,N_321);
nand U701 (N_701,N_170,N_291);
and U702 (N_702,N_367,N_289);
and U703 (N_703,N_107,N_45);
and U704 (N_704,N_172,N_81);
nand U705 (N_705,N_193,N_249);
xor U706 (N_706,N_429,N_455);
and U707 (N_707,N_284,N_424);
nor U708 (N_708,N_150,N_457);
or U709 (N_709,N_410,N_75);
nor U710 (N_710,N_479,N_26);
or U711 (N_711,N_63,N_396);
nand U712 (N_712,N_247,N_461);
nand U713 (N_713,N_271,N_490);
xor U714 (N_714,N_428,N_50);
or U715 (N_715,N_255,N_83);
and U716 (N_716,N_44,N_204);
nand U717 (N_717,N_403,N_80);
nor U718 (N_718,N_459,N_108);
nand U719 (N_719,N_306,N_275);
and U720 (N_720,N_366,N_208);
nor U721 (N_721,N_245,N_449);
or U722 (N_722,N_397,N_28);
xnor U723 (N_723,N_437,N_238);
and U724 (N_724,N_11,N_343);
and U725 (N_725,N_227,N_209);
xor U726 (N_726,N_297,N_116);
xnor U727 (N_727,N_142,N_182);
nor U728 (N_728,N_46,N_364);
or U729 (N_729,N_16,N_265);
nand U730 (N_730,N_21,N_101);
xnor U731 (N_731,N_35,N_371);
xor U732 (N_732,N_311,N_294);
nor U733 (N_733,N_211,N_323);
xnor U734 (N_734,N_235,N_66);
nand U735 (N_735,N_491,N_244);
or U736 (N_736,N_462,N_370);
nand U737 (N_737,N_62,N_332);
nor U738 (N_738,N_376,N_55);
and U739 (N_739,N_178,N_48);
nand U740 (N_740,N_96,N_158);
nor U741 (N_741,N_346,N_136);
nor U742 (N_742,N_73,N_125);
or U743 (N_743,N_333,N_488);
or U744 (N_744,N_198,N_334);
xor U745 (N_745,N_60,N_220);
xor U746 (N_746,N_446,N_146);
nand U747 (N_747,N_279,N_228);
or U748 (N_748,N_213,N_39);
or U749 (N_749,N_418,N_180);
and U750 (N_750,N_312,N_381);
or U751 (N_751,N_164,N_372);
nor U752 (N_752,N_445,N_17);
nand U753 (N_753,N_305,N_352);
or U754 (N_754,N_447,N_239);
or U755 (N_755,N_380,N_240);
nand U756 (N_756,N_21,N_418);
or U757 (N_757,N_78,N_400);
nor U758 (N_758,N_232,N_245);
xor U759 (N_759,N_389,N_211);
nor U760 (N_760,N_14,N_230);
or U761 (N_761,N_116,N_304);
nor U762 (N_762,N_73,N_370);
nand U763 (N_763,N_246,N_387);
and U764 (N_764,N_465,N_499);
xor U765 (N_765,N_330,N_350);
or U766 (N_766,N_405,N_409);
nor U767 (N_767,N_367,N_424);
xor U768 (N_768,N_479,N_147);
nor U769 (N_769,N_5,N_21);
nand U770 (N_770,N_238,N_183);
xnor U771 (N_771,N_491,N_94);
xnor U772 (N_772,N_298,N_418);
nand U773 (N_773,N_71,N_390);
or U774 (N_774,N_167,N_264);
and U775 (N_775,N_287,N_346);
nand U776 (N_776,N_89,N_441);
xnor U777 (N_777,N_259,N_122);
xor U778 (N_778,N_422,N_287);
xor U779 (N_779,N_276,N_309);
or U780 (N_780,N_238,N_143);
xnor U781 (N_781,N_234,N_302);
nor U782 (N_782,N_282,N_11);
and U783 (N_783,N_113,N_5);
or U784 (N_784,N_332,N_278);
or U785 (N_785,N_353,N_436);
or U786 (N_786,N_279,N_293);
and U787 (N_787,N_83,N_214);
or U788 (N_788,N_272,N_38);
xnor U789 (N_789,N_429,N_208);
nor U790 (N_790,N_350,N_491);
or U791 (N_791,N_261,N_18);
or U792 (N_792,N_420,N_441);
or U793 (N_793,N_69,N_83);
nand U794 (N_794,N_4,N_442);
xnor U795 (N_795,N_397,N_57);
xor U796 (N_796,N_159,N_199);
nand U797 (N_797,N_224,N_481);
nand U798 (N_798,N_23,N_89);
and U799 (N_799,N_287,N_251);
and U800 (N_800,N_265,N_175);
or U801 (N_801,N_163,N_238);
and U802 (N_802,N_212,N_290);
xnor U803 (N_803,N_40,N_28);
xor U804 (N_804,N_131,N_264);
nand U805 (N_805,N_406,N_157);
nor U806 (N_806,N_440,N_267);
nor U807 (N_807,N_449,N_93);
nor U808 (N_808,N_390,N_228);
and U809 (N_809,N_170,N_361);
nand U810 (N_810,N_297,N_275);
or U811 (N_811,N_360,N_411);
nor U812 (N_812,N_56,N_299);
or U813 (N_813,N_173,N_388);
or U814 (N_814,N_149,N_447);
and U815 (N_815,N_396,N_392);
nand U816 (N_816,N_353,N_243);
and U817 (N_817,N_83,N_161);
and U818 (N_818,N_391,N_134);
nand U819 (N_819,N_191,N_390);
xor U820 (N_820,N_62,N_40);
xnor U821 (N_821,N_239,N_401);
or U822 (N_822,N_259,N_287);
nor U823 (N_823,N_494,N_100);
nand U824 (N_824,N_447,N_39);
and U825 (N_825,N_275,N_351);
and U826 (N_826,N_345,N_253);
xor U827 (N_827,N_474,N_466);
nand U828 (N_828,N_485,N_18);
or U829 (N_829,N_23,N_68);
nor U830 (N_830,N_122,N_167);
and U831 (N_831,N_6,N_331);
and U832 (N_832,N_295,N_404);
xor U833 (N_833,N_344,N_258);
or U834 (N_834,N_498,N_346);
and U835 (N_835,N_205,N_18);
or U836 (N_836,N_155,N_358);
nor U837 (N_837,N_40,N_9);
nand U838 (N_838,N_242,N_491);
or U839 (N_839,N_159,N_457);
nand U840 (N_840,N_256,N_115);
nand U841 (N_841,N_413,N_28);
and U842 (N_842,N_273,N_287);
nor U843 (N_843,N_265,N_85);
nand U844 (N_844,N_174,N_261);
and U845 (N_845,N_91,N_27);
xor U846 (N_846,N_166,N_476);
nand U847 (N_847,N_480,N_447);
nand U848 (N_848,N_337,N_482);
or U849 (N_849,N_154,N_379);
xor U850 (N_850,N_469,N_302);
and U851 (N_851,N_98,N_217);
xnor U852 (N_852,N_489,N_376);
or U853 (N_853,N_395,N_407);
xor U854 (N_854,N_201,N_473);
nor U855 (N_855,N_146,N_313);
nor U856 (N_856,N_429,N_355);
nand U857 (N_857,N_147,N_335);
nor U858 (N_858,N_378,N_206);
nand U859 (N_859,N_219,N_266);
and U860 (N_860,N_238,N_201);
nor U861 (N_861,N_390,N_249);
nand U862 (N_862,N_236,N_435);
or U863 (N_863,N_442,N_450);
nand U864 (N_864,N_102,N_434);
nor U865 (N_865,N_126,N_409);
or U866 (N_866,N_420,N_194);
xor U867 (N_867,N_105,N_294);
xnor U868 (N_868,N_449,N_461);
and U869 (N_869,N_263,N_222);
or U870 (N_870,N_147,N_194);
nand U871 (N_871,N_231,N_399);
nor U872 (N_872,N_344,N_270);
and U873 (N_873,N_383,N_295);
nor U874 (N_874,N_237,N_253);
nand U875 (N_875,N_467,N_230);
nor U876 (N_876,N_108,N_17);
or U877 (N_877,N_89,N_141);
nor U878 (N_878,N_349,N_110);
and U879 (N_879,N_320,N_101);
xnor U880 (N_880,N_189,N_389);
nor U881 (N_881,N_150,N_492);
or U882 (N_882,N_255,N_70);
or U883 (N_883,N_326,N_201);
xnor U884 (N_884,N_497,N_486);
or U885 (N_885,N_441,N_403);
nand U886 (N_886,N_7,N_171);
and U887 (N_887,N_36,N_415);
or U888 (N_888,N_132,N_485);
or U889 (N_889,N_381,N_365);
or U890 (N_890,N_79,N_338);
or U891 (N_891,N_189,N_404);
xor U892 (N_892,N_0,N_180);
xnor U893 (N_893,N_183,N_88);
and U894 (N_894,N_308,N_405);
or U895 (N_895,N_443,N_291);
xnor U896 (N_896,N_312,N_146);
or U897 (N_897,N_123,N_264);
nor U898 (N_898,N_350,N_297);
and U899 (N_899,N_172,N_93);
xor U900 (N_900,N_185,N_467);
and U901 (N_901,N_66,N_126);
nand U902 (N_902,N_18,N_134);
and U903 (N_903,N_129,N_81);
nand U904 (N_904,N_397,N_88);
nand U905 (N_905,N_332,N_43);
xnor U906 (N_906,N_307,N_446);
or U907 (N_907,N_132,N_361);
and U908 (N_908,N_473,N_288);
nor U909 (N_909,N_189,N_244);
or U910 (N_910,N_291,N_177);
or U911 (N_911,N_453,N_391);
and U912 (N_912,N_62,N_421);
nor U913 (N_913,N_57,N_317);
nor U914 (N_914,N_387,N_470);
nand U915 (N_915,N_184,N_398);
or U916 (N_916,N_103,N_279);
nand U917 (N_917,N_246,N_350);
xor U918 (N_918,N_353,N_9);
nor U919 (N_919,N_211,N_418);
nand U920 (N_920,N_307,N_430);
and U921 (N_921,N_238,N_395);
xnor U922 (N_922,N_46,N_174);
or U923 (N_923,N_137,N_294);
nor U924 (N_924,N_242,N_109);
nor U925 (N_925,N_457,N_8);
or U926 (N_926,N_243,N_412);
nand U927 (N_927,N_150,N_289);
or U928 (N_928,N_417,N_450);
and U929 (N_929,N_206,N_68);
nand U930 (N_930,N_443,N_445);
or U931 (N_931,N_418,N_463);
nand U932 (N_932,N_391,N_407);
nand U933 (N_933,N_57,N_142);
nand U934 (N_934,N_244,N_226);
xnor U935 (N_935,N_491,N_169);
xor U936 (N_936,N_481,N_292);
nand U937 (N_937,N_350,N_316);
nand U938 (N_938,N_108,N_321);
or U939 (N_939,N_410,N_183);
or U940 (N_940,N_136,N_156);
xor U941 (N_941,N_199,N_454);
or U942 (N_942,N_94,N_498);
nor U943 (N_943,N_13,N_227);
or U944 (N_944,N_358,N_90);
or U945 (N_945,N_83,N_205);
nor U946 (N_946,N_492,N_82);
and U947 (N_947,N_6,N_302);
and U948 (N_948,N_191,N_230);
nor U949 (N_949,N_27,N_323);
or U950 (N_950,N_66,N_333);
nor U951 (N_951,N_57,N_421);
nand U952 (N_952,N_250,N_169);
nor U953 (N_953,N_281,N_128);
and U954 (N_954,N_441,N_59);
xor U955 (N_955,N_92,N_229);
or U956 (N_956,N_75,N_195);
nor U957 (N_957,N_272,N_287);
xor U958 (N_958,N_288,N_401);
nand U959 (N_959,N_120,N_45);
xnor U960 (N_960,N_139,N_134);
and U961 (N_961,N_351,N_74);
nor U962 (N_962,N_68,N_493);
or U963 (N_963,N_495,N_247);
and U964 (N_964,N_224,N_17);
nand U965 (N_965,N_284,N_72);
and U966 (N_966,N_296,N_431);
xnor U967 (N_967,N_396,N_365);
or U968 (N_968,N_13,N_118);
nor U969 (N_969,N_308,N_423);
and U970 (N_970,N_384,N_331);
xor U971 (N_971,N_366,N_398);
nor U972 (N_972,N_490,N_278);
xor U973 (N_973,N_151,N_174);
xor U974 (N_974,N_107,N_459);
nor U975 (N_975,N_195,N_340);
nor U976 (N_976,N_73,N_262);
and U977 (N_977,N_430,N_42);
xnor U978 (N_978,N_267,N_468);
nor U979 (N_979,N_469,N_32);
nor U980 (N_980,N_173,N_108);
xor U981 (N_981,N_379,N_225);
xnor U982 (N_982,N_20,N_5);
nor U983 (N_983,N_238,N_455);
nand U984 (N_984,N_290,N_106);
xnor U985 (N_985,N_381,N_275);
xor U986 (N_986,N_48,N_163);
or U987 (N_987,N_457,N_297);
and U988 (N_988,N_40,N_83);
and U989 (N_989,N_466,N_333);
or U990 (N_990,N_281,N_211);
or U991 (N_991,N_415,N_490);
and U992 (N_992,N_419,N_373);
or U993 (N_993,N_188,N_349);
and U994 (N_994,N_214,N_419);
and U995 (N_995,N_198,N_349);
and U996 (N_996,N_444,N_323);
nand U997 (N_997,N_358,N_310);
and U998 (N_998,N_443,N_497);
nor U999 (N_999,N_146,N_126);
and U1000 (N_1000,N_726,N_998);
and U1001 (N_1001,N_632,N_549);
xnor U1002 (N_1002,N_780,N_671);
xor U1003 (N_1003,N_870,N_679);
nand U1004 (N_1004,N_557,N_837);
nand U1005 (N_1005,N_638,N_530);
nor U1006 (N_1006,N_527,N_743);
nand U1007 (N_1007,N_667,N_613);
xor U1008 (N_1008,N_740,N_832);
nand U1009 (N_1009,N_920,N_827);
and U1010 (N_1010,N_548,N_725);
nand U1011 (N_1011,N_787,N_934);
nand U1012 (N_1012,N_744,N_552);
and U1013 (N_1013,N_994,N_755);
and U1014 (N_1014,N_952,N_907);
nor U1015 (N_1015,N_881,N_719);
nand U1016 (N_1016,N_500,N_783);
or U1017 (N_1017,N_721,N_931);
and U1018 (N_1018,N_945,N_944);
nand U1019 (N_1019,N_504,N_596);
and U1020 (N_1020,N_689,N_588);
xnor U1021 (N_1021,N_751,N_915);
or U1022 (N_1022,N_851,N_752);
xor U1023 (N_1023,N_763,N_695);
nand U1024 (N_1024,N_977,N_899);
nor U1025 (N_1025,N_987,N_676);
nand U1026 (N_1026,N_649,N_554);
and U1027 (N_1027,N_611,N_879);
nand U1028 (N_1028,N_801,N_760);
nand U1029 (N_1029,N_909,N_798);
nand U1030 (N_1030,N_634,N_956);
xnor U1031 (N_1031,N_631,N_584);
xor U1032 (N_1032,N_651,N_652);
xor U1033 (N_1033,N_785,N_908);
or U1034 (N_1034,N_943,N_550);
xor U1035 (N_1035,N_647,N_856);
xor U1036 (N_1036,N_947,N_960);
and U1037 (N_1037,N_929,N_581);
and U1038 (N_1038,N_720,N_556);
xor U1039 (N_1039,N_761,N_547);
nand U1040 (N_1040,N_742,N_996);
and U1041 (N_1041,N_767,N_949);
nand U1042 (N_1042,N_735,N_904);
or U1043 (N_1043,N_703,N_619);
or U1044 (N_1044,N_746,N_590);
xor U1045 (N_1045,N_933,N_655);
nand U1046 (N_1046,N_520,N_993);
xnor U1047 (N_1047,N_800,N_535);
nor U1048 (N_1048,N_525,N_635);
nor U1049 (N_1049,N_587,N_958);
xor U1050 (N_1050,N_858,N_511);
and U1051 (N_1051,N_989,N_970);
nor U1052 (N_1052,N_999,N_797);
nand U1053 (N_1053,N_646,N_670);
or U1054 (N_1054,N_806,N_985);
nand U1055 (N_1055,N_821,N_967);
xor U1056 (N_1056,N_810,N_968);
xor U1057 (N_1057,N_690,N_561);
and U1058 (N_1058,N_862,N_733);
nand U1059 (N_1059,N_809,N_568);
nor U1060 (N_1060,N_974,N_641);
xnor U1061 (N_1061,N_616,N_937);
nand U1062 (N_1062,N_653,N_512);
and U1063 (N_1063,N_747,N_845);
xor U1064 (N_1064,N_766,N_551);
xor U1065 (N_1065,N_939,N_792);
nand U1066 (N_1066,N_555,N_532);
or U1067 (N_1067,N_776,N_694);
nand U1068 (N_1068,N_836,N_546);
and U1069 (N_1069,N_519,N_893);
nor U1070 (N_1070,N_846,N_591);
xnor U1071 (N_1071,N_608,N_748);
xor U1072 (N_1072,N_901,N_618);
or U1073 (N_1073,N_749,N_501);
nor U1074 (N_1074,N_738,N_623);
or U1075 (N_1075,N_764,N_681);
or U1076 (N_1076,N_964,N_637);
xor U1077 (N_1077,N_951,N_839);
nor U1078 (N_1078,N_636,N_536);
or U1079 (N_1079,N_718,N_678);
nand U1080 (N_1080,N_789,N_788);
nand U1081 (N_1081,N_734,N_669);
nand U1082 (N_1082,N_991,N_713);
and U1083 (N_1083,N_835,N_779);
nand U1084 (N_1084,N_715,N_603);
nand U1085 (N_1085,N_615,N_852);
and U1086 (N_1086,N_875,N_658);
and U1087 (N_1087,N_804,N_697);
xnor U1088 (N_1088,N_514,N_538);
and U1089 (N_1089,N_888,N_969);
or U1090 (N_1090,N_957,N_874);
nand U1091 (N_1091,N_825,N_579);
and U1092 (N_1092,N_932,N_540);
or U1093 (N_1093,N_553,N_771);
or U1094 (N_1094,N_795,N_811);
xnor U1095 (N_1095,N_539,N_572);
or U1096 (N_1096,N_844,N_592);
or U1097 (N_1097,N_574,N_762);
nand U1098 (N_1098,N_843,N_633);
xor U1099 (N_1099,N_656,N_923);
nand U1100 (N_1100,N_600,N_509);
nor U1101 (N_1101,N_973,N_775);
and U1102 (N_1102,N_558,N_781);
or U1103 (N_1103,N_707,N_942);
xnor U1104 (N_1104,N_793,N_502);
nand U1105 (N_1105,N_891,N_950);
and U1106 (N_1106,N_817,N_883);
nand U1107 (N_1107,N_796,N_823);
xnor U1108 (N_1108,N_867,N_864);
nand U1109 (N_1109,N_685,N_575);
or U1110 (N_1110,N_595,N_505);
nor U1111 (N_1111,N_978,N_814);
xor U1112 (N_1112,N_666,N_599);
xnor U1113 (N_1113,N_571,N_570);
nor U1114 (N_1114,N_765,N_544);
and U1115 (N_1115,N_869,N_754);
xor U1116 (N_1116,N_963,N_882);
nand U1117 (N_1117,N_770,N_808);
nor U1118 (N_1118,N_887,N_576);
nor U1119 (N_1119,N_531,N_569);
and U1120 (N_1120,N_868,N_622);
xnor U1121 (N_1121,N_739,N_753);
xnor U1122 (N_1122,N_699,N_803);
nand U1123 (N_1123,N_605,N_946);
xor U1124 (N_1124,N_717,N_861);
and U1125 (N_1125,N_782,N_833);
nor U1126 (N_1126,N_626,N_979);
or U1127 (N_1127,N_838,N_709);
or U1128 (N_1128,N_683,N_773);
xor U1129 (N_1129,N_992,N_598);
and U1130 (N_1130,N_854,N_645);
or U1131 (N_1131,N_863,N_995);
or U1132 (N_1132,N_898,N_729);
or U1133 (N_1133,N_961,N_857);
or U1134 (N_1134,N_938,N_872);
xor U1135 (N_1135,N_900,N_819);
nand U1136 (N_1136,N_545,N_693);
and U1137 (N_1137,N_614,N_503);
xnor U1138 (N_1138,N_971,N_559);
nand U1139 (N_1139,N_628,N_842);
and U1140 (N_1140,N_829,N_704);
or U1141 (N_1141,N_563,N_745);
nor U1142 (N_1142,N_830,N_736);
or U1143 (N_1143,N_688,N_962);
nor U1144 (N_1144,N_702,N_813);
nand U1145 (N_1145,N_711,N_533);
xor U1146 (N_1146,N_648,N_507);
nor U1147 (N_1147,N_659,N_573);
xnor U1148 (N_1148,N_912,N_822);
and U1149 (N_1149,N_597,N_928);
or U1150 (N_1150,N_654,N_625);
and U1151 (N_1151,N_786,N_680);
xor U1152 (N_1152,N_741,N_586);
nand U1153 (N_1153,N_542,N_802);
xnor U1154 (N_1154,N_620,N_642);
or U1155 (N_1155,N_650,N_828);
xor U1156 (N_1156,N_727,N_609);
nor U1157 (N_1157,N_566,N_955);
or U1158 (N_1158,N_884,N_757);
nor U1159 (N_1159,N_853,N_737);
and U1160 (N_1160,N_583,N_914);
xor U1161 (N_1161,N_878,N_807);
nor U1162 (N_1162,N_948,N_799);
xnor U1163 (N_1163,N_758,N_664);
xor U1164 (N_1164,N_723,N_630);
nor U1165 (N_1165,N_759,N_521);
nand U1166 (N_1166,N_921,N_522);
xnor U1167 (N_1167,N_750,N_988);
nor U1168 (N_1168,N_919,N_940);
xor U1169 (N_1169,N_784,N_812);
and U1170 (N_1170,N_567,N_660);
nor U1171 (N_1171,N_663,N_824);
nor U1172 (N_1172,N_578,N_529);
nand U1173 (N_1173,N_980,N_692);
nor U1174 (N_1174,N_935,N_816);
or U1175 (N_1175,N_722,N_976);
or U1176 (N_1176,N_643,N_959);
nor U1177 (N_1177,N_585,N_589);
xnor U1178 (N_1178,N_984,N_714);
nand U1179 (N_1179,N_537,N_768);
and U1180 (N_1180,N_541,N_708);
nand U1181 (N_1181,N_665,N_716);
and U1182 (N_1182,N_657,N_865);
and U1183 (N_1183,N_691,N_954);
nor U1184 (N_1184,N_880,N_774);
nor U1185 (N_1185,N_661,N_906);
nand U1186 (N_1186,N_617,N_917);
and U1187 (N_1187,N_674,N_841);
nor U1188 (N_1188,N_518,N_885);
and U1189 (N_1189,N_602,N_965);
or U1190 (N_1190,N_582,N_925);
xor U1191 (N_1191,N_922,N_728);
and U1192 (N_1192,N_860,N_517);
nor U1193 (N_1193,N_902,N_769);
and U1194 (N_1194,N_700,N_639);
and U1195 (N_1195,N_516,N_560);
xor U1196 (N_1196,N_930,N_896);
nand U1197 (N_1197,N_818,N_778);
or U1198 (N_1198,N_668,N_756);
nor U1199 (N_1199,N_953,N_990);
or U1200 (N_1200,N_684,N_840);
xnor U1201 (N_1201,N_831,N_936);
nor U1202 (N_1202,N_580,N_903);
or U1203 (N_1203,N_918,N_565);
and U1204 (N_1204,N_866,N_966);
and U1205 (N_1205,N_847,N_859);
nor U1206 (N_1206,N_834,N_673);
nand U1207 (N_1207,N_850,N_941);
and U1208 (N_1208,N_927,N_562);
nand U1209 (N_1209,N_815,N_772);
and U1210 (N_1210,N_604,N_820);
nand U1211 (N_1211,N_916,N_601);
and U1212 (N_1212,N_805,N_577);
xnor U1213 (N_1213,N_731,N_712);
nand U1214 (N_1214,N_886,N_594);
or U1215 (N_1215,N_730,N_975);
nand U1216 (N_1216,N_911,N_826);
xor U1217 (N_1217,N_791,N_972);
nor U1218 (N_1218,N_892,N_777);
xor U1219 (N_1219,N_686,N_706);
and U1220 (N_1220,N_705,N_528);
and U1221 (N_1221,N_640,N_675);
or U1222 (N_1222,N_513,N_894);
nand U1223 (N_1223,N_794,N_593);
or U1224 (N_1224,N_523,N_644);
or U1225 (N_1225,N_997,N_629);
xnor U1226 (N_1226,N_926,N_889);
and U1227 (N_1227,N_687,N_895);
nand U1228 (N_1228,N_986,N_871);
nor U1229 (N_1229,N_607,N_515);
nor U1230 (N_1230,N_982,N_877);
and U1231 (N_1231,N_682,N_610);
xor U1232 (N_1232,N_873,N_983);
or U1233 (N_1233,N_543,N_698);
or U1234 (N_1234,N_621,N_696);
or U1235 (N_1235,N_855,N_913);
xnor U1236 (N_1236,N_510,N_724);
or U1237 (N_1237,N_677,N_981);
or U1238 (N_1238,N_564,N_662);
nand U1239 (N_1239,N_672,N_710);
nand U1240 (N_1240,N_506,N_890);
xor U1241 (N_1241,N_897,N_624);
xnor U1242 (N_1242,N_905,N_910);
or U1243 (N_1243,N_701,N_627);
nor U1244 (N_1244,N_526,N_924);
nor U1245 (N_1245,N_534,N_849);
or U1246 (N_1246,N_612,N_524);
nand U1247 (N_1247,N_848,N_606);
nand U1248 (N_1248,N_876,N_790);
nor U1249 (N_1249,N_732,N_508);
or U1250 (N_1250,N_835,N_908);
or U1251 (N_1251,N_954,N_814);
nor U1252 (N_1252,N_957,N_784);
xnor U1253 (N_1253,N_661,N_837);
nand U1254 (N_1254,N_669,N_905);
nor U1255 (N_1255,N_518,N_800);
or U1256 (N_1256,N_917,N_802);
nor U1257 (N_1257,N_624,N_885);
xnor U1258 (N_1258,N_721,N_651);
nand U1259 (N_1259,N_774,N_501);
nor U1260 (N_1260,N_955,N_517);
and U1261 (N_1261,N_963,N_745);
or U1262 (N_1262,N_903,N_820);
nand U1263 (N_1263,N_845,N_978);
or U1264 (N_1264,N_527,N_959);
xnor U1265 (N_1265,N_927,N_571);
nor U1266 (N_1266,N_653,N_831);
xor U1267 (N_1267,N_744,N_580);
nand U1268 (N_1268,N_844,N_674);
xnor U1269 (N_1269,N_552,N_967);
nand U1270 (N_1270,N_785,N_731);
or U1271 (N_1271,N_932,N_997);
nor U1272 (N_1272,N_987,N_757);
or U1273 (N_1273,N_611,N_739);
nor U1274 (N_1274,N_793,N_898);
or U1275 (N_1275,N_894,N_880);
or U1276 (N_1276,N_760,N_542);
and U1277 (N_1277,N_680,N_871);
nor U1278 (N_1278,N_824,N_936);
or U1279 (N_1279,N_959,N_677);
and U1280 (N_1280,N_803,N_733);
and U1281 (N_1281,N_817,N_926);
xnor U1282 (N_1282,N_730,N_721);
nand U1283 (N_1283,N_658,N_500);
or U1284 (N_1284,N_962,N_758);
nor U1285 (N_1285,N_695,N_571);
nand U1286 (N_1286,N_619,N_740);
xnor U1287 (N_1287,N_502,N_831);
and U1288 (N_1288,N_673,N_570);
and U1289 (N_1289,N_910,N_880);
nor U1290 (N_1290,N_933,N_974);
or U1291 (N_1291,N_760,N_563);
or U1292 (N_1292,N_534,N_787);
nor U1293 (N_1293,N_994,N_806);
or U1294 (N_1294,N_973,N_938);
and U1295 (N_1295,N_523,N_826);
and U1296 (N_1296,N_618,N_993);
nor U1297 (N_1297,N_809,N_675);
nor U1298 (N_1298,N_542,N_509);
and U1299 (N_1299,N_568,N_694);
nor U1300 (N_1300,N_852,N_715);
xnor U1301 (N_1301,N_757,N_612);
or U1302 (N_1302,N_656,N_648);
nand U1303 (N_1303,N_684,N_857);
nand U1304 (N_1304,N_932,N_732);
and U1305 (N_1305,N_817,N_557);
xnor U1306 (N_1306,N_513,N_575);
nand U1307 (N_1307,N_642,N_617);
or U1308 (N_1308,N_778,N_834);
or U1309 (N_1309,N_994,N_674);
nand U1310 (N_1310,N_616,N_677);
nand U1311 (N_1311,N_673,N_771);
or U1312 (N_1312,N_669,N_612);
or U1313 (N_1313,N_538,N_523);
or U1314 (N_1314,N_608,N_538);
nor U1315 (N_1315,N_752,N_547);
and U1316 (N_1316,N_975,N_537);
xor U1317 (N_1317,N_916,N_741);
xnor U1318 (N_1318,N_691,N_839);
nor U1319 (N_1319,N_981,N_630);
nand U1320 (N_1320,N_859,N_963);
and U1321 (N_1321,N_617,N_976);
or U1322 (N_1322,N_814,N_580);
or U1323 (N_1323,N_919,N_911);
and U1324 (N_1324,N_698,N_683);
nor U1325 (N_1325,N_784,N_937);
nor U1326 (N_1326,N_574,N_934);
or U1327 (N_1327,N_922,N_704);
nand U1328 (N_1328,N_962,N_567);
nand U1329 (N_1329,N_512,N_908);
or U1330 (N_1330,N_618,N_911);
xnor U1331 (N_1331,N_544,N_739);
nand U1332 (N_1332,N_704,N_635);
nor U1333 (N_1333,N_718,N_994);
xnor U1334 (N_1334,N_562,N_893);
and U1335 (N_1335,N_622,N_586);
nand U1336 (N_1336,N_806,N_580);
and U1337 (N_1337,N_794,N_550);
or U1338 (N_1338,N_887,N_666);
and U1339 (N_1339,N_974,N_762);
xor U1340 (N_1340,N_554,N_847);
and U1341 (N_1341,N_970,N_765);
nand U1342 (N_1342,N_962,N_862);
and U1343 (N_1343,N_809,N_657);
or U1344 (N_1344,N_710,N_856);
and U1345 (N_1345,N_938,N_569);
nand U1346 (N_1346,N_760,N_847);
or U1347 (N_1347,N_828,N_647);
nand U1348 (N_1348,N_928,N_997);
nand U1349 (N_1349,N_809,N_621);
and U1350 (N_1350,N_674,N_978);
and U1351 (N_1351,N_782,N_921);
xnor U1352 (N_1352,N_840,N_581);
xnor U1353 (N_1353,N_503,N_934);
and U1354 (N_1354,N_522,N_534);
nor U1355 (N_1355,N_588,N_811);
and U1356 (N_1356,N_885,N_830);
nor U1357 (N_1357,N_996,N_797);
nor U1358 (N_1358,N_806,N_693);
nand U1359 (N_1359,N_757,N_790);
xor U1360 (N_1360,N_948,N_612);
or U1361 (N_1361,N_662,N_856);
and U1362 (N_1362,N_817,N_637);
and U1363 (N_1363,N_877,N_671);
nor U1364 (N_1364,N_690,N_983);
or U1365 (N_1365,N_977,N_755);
xnor U1366 (N_1366,N_678,N_644);
nand U1367 (N_1367,N_960,N_950);
nand U1368 (N_1368,N_712,N_799);
nand U1369 (N_1369,N_900,N_615);
or U1370 (N_1370,N_606,N_686);
or U1371 (N_1371,N_670,N_888);
nand U1372 (N_1372,N_925,N_910);
nand U1373 (N_1373,N_620,N_930);
nand U1374 (N_1374,N_812,N_877);
nand U1375 (N_1375,N_608,N_820);
nand U1376 (N_1376,N_726,N_550);
nor U1377 (N_1377,N_543,N_851);
nor U1378 (N_1378,N_611,N_900);
xnor U1379 (N_1379,N_977,N_595);
nand U1380 (N_1380,N_621,N_681);
xnor U1381 (N_1381,N_911,N_934);
nand U1382 (N_1382,N_737,N_857);
and U1383 (N_1383,N_521,N_998);
nand U1384 (N_1384,N_824,N_666);
or U1385 (N_1385,N_598,N_537);
nor U1386 (N_1386,N_520,N_685);
nor U1387 (N_1387,N_755,N_966);
nor U1388 (N_1388,N_983,N_776);
nor U1389 (N_1389,N_988,N_688);
nor U1390 (N_1390,N_887,N_725);
and U1391 (N_1391,N_783,N_635);
and U1392 (N_1392,N_986,N_678);
nand U1393 (N_1393,N_836,N_651);
or U1394 (N_1394,N_988,N_839);
nor U1395 (N_1395,N_860,N_969);
xor U1396 (N_1396,N_810,N_773);
or U1397 (N_1397,N_684,N_961);
xnor U1398 (N_1398,N_720,N_565);
nor U1399 (N_1399,N_515,N_559);
and U1400 (N_1400,N_576,N_885);
xnor U1401 (N_1401,N_510,N_727);
and U1402 (N_1402,N_675,N_734);
and U1403 (N_1403,N_504,N_878);
and U1404 (N_1404,N_706,N_646);
nand U1405 (N_1405,N_697,N_780);
or U1406 (N_1406,N_702,N_715);
xor U1407 (N_1407,N_939,N_521);
nand U1408 (N_1408,N_801,N_583);
nor U1409 (N_1409,N_800,N_594);
or U1410 (N_1410,N_867,N_592);
and U1411 (N_1411,N_557,N_537);
or U1412 (N_1412,N_532,N_583);
nor U1413 (N_1413,N_761,N_791);
xnor U1414 (N_1414,N_910,N_746);
nor U1415 (N_1415,N_741,N_552);
nor U1416 (N_1416,N_685,N_880);
xor U1417 (N_1417,N_911,N_877);
xor U1418 (N_1418,N_604,N_731);
nor U1419 (N_1419,N_789,N_956);
nor U1420 (N_1420,N_546,N_750);
or U1421 (N_1421,N_911,N_921);
and U1422 (N_1422,N_821,N_909);
and U1423 (N_1423,N_671,N_993);
and U1424 (N_1424,N_799,N_553);
xor U1425 (N_1425,N_698,N_727);
nor U1426 (N_1426,N_730,N_958);
nor U1427 (N_1427,N_764,N_953);
nand U1428 (N_1428,N_603,N_833);
or U1429 (N_1429,N_593,N_998);
or U1430 (N_1430,N_855,N_695);
nor U1431 (N_1431,N_589,N_694);
and U1432 (N_1432,N_542,N_826);
xnor U1433 (N_1433,N_653,N_901);
or U1434 (N_1434,N_713,N_957);
or U1435 (N_1435,N_625,N_977);
nor U1436 (N_1436,N_724,N_899);
and U1437 (N_1437,N_626,N_947);
nor U1438 (N_1438,N_906,N_791);
nor U1439 (N_1439,N_510,N_625);
and U1440 (N_1440,N_599,N_562);
and U1441 (N_1441,N_560,N_832);
or U1442 (N_1442,N_873,N_813);
and U1443 (N_1443,N_619,N_771);
xnor U1444 (N_1444,N_838,N_805);
xnor U1445 (N_1445,N_848,N_882);
or U1446 (N_1446,N_707,N_592);
nand U1447 (N_1447,N_667,N_747);
nand U1448 (N_1448,N_888,N_610);
nand U1449 (N_1449,N_698,N_531);
or U1450 (N_1450,N_895,N_850);
xnor U1451 (N_1451,N_851,N_807);
nand U1452 (N_1452,N_727,N_563);
xnor U1453 (N_1453,N_951,N_701);
nand U1454 (N_1454,N_838,N_901);
or U1455 (N_1455,N_714,N_892);
nor U1456 (N_1456,N_947,N_807);
or U1457 (N_1457,N_992,N_778);
or U1458 (N_1458,N_599,N_581);
xnor U1459 (N_1459,N_521,N_660);
xnor U1460 (N_1460,N_909,N_644);
nand U1461 (N_1461,N_976,N_598);
xor U1462 (N_1462,N_643,N_866);
xnor U1463 (N_1463,N_676,N_980);
nand U1464 (N_1464,N_643,N_838);
nor U1465 (N_1465,N_990,N_757);
nor U1466 (N_1466,N_773,N_515);
or U1467 (N_1467,N_566,N_770);
or U1468 (N_1468,N_658,N_601);
or U1469 (N_1469,N_679,N_524);
and U1470 (N_1470,N_920,N_580);
nor U1471 (N_1471,N_547,N_670);
and U1472 (N_1472,N_512,N_655);
nand U1473 (N_1473,N_714,N_669);
nor U1474 (N_1474,N_611,N_811);
and U1475 (N_1475,N_723,N_957);
nor U1476 (N_1476,N_825,N_558);
nor U1477 (N_1477,N_765,N_717);
xor U1478 (N_1478,N_878,N_925);
nand U1479 (N_1479,N_725,N_866);
and U1480 (N_1480,N_849,N_519);
nand U1481 (N_1481,N_941,N_753);
and U1482 (N_1482,N_578,N_827);
nor U1483 (N_1483,N_641,N_935);
or U1484 (N_1484,N_926,N_561);
xnor U1485 (N_1485,N_805,N_913);
and U1486 (N_1486,N_798,N_729);
and U1487 (N_1487,N_614,N_799);
nor U1488 (N_1488,N_965,N_869);
and U1489 (N_1489,N_622,N_580);
nand U1490 (N_1490,N_578,N_838);
or U1491 (N_1491,N_941,N_719);
nor U1492 (N_1492,N_654,N_641);
nor U1493 (N_1493,N_827,N_812);
or U1494 (N_1494,N_778,N_655);
xor U1495 (N_1495,N_878,N_536);
xnor U1496 (N_1496,N_935,N_574);
or U1497 (N_1497,N_648,N_609);
and U1498 (N_1498,N_558,N_819);
nand U1499 (N_1499,N_847,N_550);
or U1500 (N_1500,N_1499,N_1142);
xor U1501 (N_1501,N_1040,N_1353);
and U1502 (N_1502,N_1166,N_1216);
xnor U1503 (N_1503,N_1099,N_1363);
nor U1504 (N_1504,N_1392,N_1404);
and U1505 (N_1505,N_1069,N_1478);
nor U1506 (N_1506,N_1461,N_1447);
nand U1507 (N_1507,N_1211,N_1085);
nand U1508 (N_1508,N_1480,N_1124);
nand U1509 (N_1509,N_1373,N_1222);
and U1510 (N_1510,N_1395,N_1377);
xor U1511 (N_1511,N_1173,N_1036);
and U1512 (N_1512,N_1427,N_1109);
nor U1513 (N_1513,N_1138,N_1150);
and U1514 (N_1514,N_1274,N_1000);
nor U1515 (N_1515,N_1424,N_1141);
or U1516 (N_1516,N_1301,N_1198);
nand U1517 (N_1517,N_1453,N_1001);
or U1518 (N_1518,N_1045,N_1105);
nor U1519 (N_1519,N_1039,N_1027);
nor U1520 (N_1520,N_1237,N_1153);
xnor U1521 (N_1521,N_1350,N_1359);
or U1522 (N_1522,N_1052,N_1050);
or U1523 (N_1523,N_1414,N_1464);
nand U1524 (N_1524,N_1056,N_1181);
nand U1525 (N_1525,N_1362,N_1435);
or U1526 (N_1526,N_1005,N_1335);
xor U1527 (N_1527,N_1061,N_1397);
and U1528 (N_1528,N_1175,N_1345);
xnor U1529 (N_1529,N_1187,N_1016);
and U1530 (N_1530,N_1133,N_1254);
xnor U1531 (N_1531,N_1313,N_1342);
and U1532 (N_1532,N_1223,N_1070);
or U1533 (N_1533,N_1438,N_1382);
nand U1534 (N_1534,N_1215,N_1264);
nand U1535 (N_1535,N_1148,N_1433);
nor U1536 (N_1536,N_1126,N_1064);
xnor U1537 (N_1537,N_1421,N_1008);
xnor U1538 (N_1538,N_1170,N_1365);
and U1539 (N_1539,N_1472,N_1408);
or U1540 (N_1540,N_1488,N_1169);
nand U1541 (N_1541,N_1010,N_1006);
xor U1542 (N_1542,N_1409,N_1367);
and U1543 (N_1543,N_1068,N_1086);
nor U1544 (N_1544,N_1381,N_1243);
xnor U1545 (N_1545,N_1317,N_1053);
xnor U1546 (N_1546,N_1004,N_1405);
nand U1547 (N_1547,N_1284,N_1327);
nand U1548 (N_1548,N_1297,N_1213);
nor U1549 (N_1549,N_1320,N_1432);
nand U1550 (N_1550,N_1374,N_1116);
xnor U1551 (N_1551,N_1048,N_1410);
nand U1552 (N_1552,N_1390,N_1339);
nand U1553 (N_1553,N_1046,N_1009);
or U1554 (N_1554,N_1154,N_1298);
and U1555 (N_1555,N_1292,N_1497);
nand U1556 (N_1556,N_1236,N_1445);
nand U1557 (N_1557,N_1143,N_1330);
nor U1558 (N_1558,N_1411,N_1283);
and U1559 (N_1559,N_1087,N_1097);
or U1560 (N_1560,N_1426,N_1442);
or U1561 (N_1561,N_1220,N_1078);
or U1562 (N_1562,N_1398,N_1029);
and U1563 (N_1563,N_1119,N_1376);
xor U1564 (N_1564,N_1380,N_1067);
and U1565 (N_1565,N_1309,N_1366);
nor U1566 (N_1566,N_1307,N_1192);
or U1567 (N_1567,N_1174,N_1475);
or U1568 (N_1568,N_1389,N_1384);
or U1569 (N_1569,N_1108,N_1295);
nor U1570 (N_1570,N_1144,N_1028);
or U1571 (N_1571,N_1195,N_1204);
nor U1572 (N_1572,N_1130,N_1071);
or U1573 (N_1573,N_1123,N_1232);
and U1574 (N_1574,N_1022,N_1399);
or U1575 (N_1575,N_1100,N_1332);
nor U1576 (N_1576,N_1163,N_1455);
nand U1577 (N_1577,N_1172,N_1302);
or U1578 (N_1578,N_1158,N_1055);
or U1579 (N_1579,N_1226,N_1114);
or U1580 (N_1580,N_1337,N_1280);
nor U1581 (N_1581,N_1089,N_1407);
nor U1582 (N_1582,N_1458,N_1104);
nor U1583 (N_1583,N_1315,N_1203);
nor U1584 (N_1584,N_1401,N_1075);
nand U1585 (N_1585,N_1420,N_1454);
and U1586 (N_1586,N_1128,N_1122);
xnor U1587 (N_1587,N_1155,N_1498);
and U1588 (N_1588,N_1391,N_1278);
and U1589 (N_1589,N_1256,N_1487);
nor U1590 (N_1590,N_1316,N_1031);
nor U1591 (N_1591,N_1121,N_1451);
or U1592 (N_1592,N_1357,N_1265);
nor U1593 (N_1593,N_1025,N_1033);
or U1594 (N_1594,N_1466,N_1344);
nor U1595 (N_1595,N_1465,N_1267);
or U1596 (N_1596,N_1347,N_1090);
nand U1597 (N_1597,N_1214,N_1444);
nor U1598 (N_1598,N_1191,N_1462);
xor U1599 (N_1599,N_1251,N_1245);
xor U1600 (N_1600,N_1221,N_1477);
nand U1601 (N_1601,N_1197,N_1188);
and U1602 (N_1602,N_1494,N_1452);
xnor U1603 (N_1603,N_1250,N_1208);
and U1604 (N_1604,N_1088,N_1471);
nor U1605 (N_1605,N_1176,N_1279);
xnor U1606 (N_1606,N_1467,N_1486);
and U1607 (N_1607,N_1282,N_1247);
and U1608 (N_1608,N_1019,N_1135);
xnor U1609 (N_1609,N_1288,N_1259);
xor U1610 (N_1610,N_1246,N_1326);
and U1611 (N_1611,N_1034,N_1349);
nor U1612 (N_1612,N_1129,N_1300);
nand U1613 (N_1613,N_1371,N_1358);
xor U1614 (N_1614,N_1098,N_1079);
nand U1615 (N_1615,N_1449,N_1348);
or U1616 (N_1616,N_1151,N_1492);
and U1617 (N_1617,N_1217,N_1043);
nor U1618 (N_1618,N_1329,N_1253);
nand U1619 (N_1619,N_1383,N_1396);
nand U1620 (N_1620,N_1355,N_1402);
xor U1621 (N_1621,N_1096,N_1375);
xor U1622 (N_1622,N_1092,N_1418);
nor U1623 (N_1623,N_1140,N_1314);
nand U1624 (N_1624,N_1023,N_1269);
xor U1625 (N_1625,N_1131,N_1196);
or U1626 (N_1626,N_1485,N_1352);
and U1627 (N_1627,N_1030,N_1094);
and U1628 (N_1628,N_1037,N_1060);
nand U1629 (N_1629,N_1341,N_1115);
nand U1630 (N_1630,N_1406,N_1102);
nand U1631 (N_1631,N_1178,N_1035);
and U1632 (N_1632,N_1311,N_1281);
nor U1633 (N_1633,N_1177,N_1106);
xnor U1634 (N_1634,N_1272,N_1428);
or U1635 (N_1635,N_1412,N_1066);
and U1636 (N_1636,N_1002,N_1038);
xnor U1637 (N_1637,N_1275,N_1419);
and U1638 (N_1638,N_1051,N_1474);
nor U1639 (N_1639,N_1183,N_1057);
nor U1640 (N_1640,N_1026,N_1047);
nor U1641 (N_1641,N_1145,N_1261);
nor U1642 (N_1642,N_1185,N_1491);
or U1643 (N_1643,N_1241,N_1457);
or U1644 (N_1644,N_1334,N_1328);
nor U1645 (N_1645,N_1325,N_1448);
nor U1646 (N_1646,N_1294,N_1331);
xnor U1647 (N_1647,N_1137,N_1270);
or U1648 (N_1648,N_1413,N_1062);
and U1649 (N_1649,N_1014,N_1082);
nor U1650 (N_1650,N_1430,N_1200);
xor U1651 (N_1651,N_1291,N_1489);
nand U1652 (N_1652,N_1361,N_1290);
or U1653 (N_1653,N_1120,N_1400);
xnor U1654 (N_1654,N_1072,N_1423);
xor U1655 (N_1655,N_1012,N_1224);
nor U1656 (N_1656,N_1091,N_1289);
or U1657 (N_1657,N_1493,N_1323);
xnor U1658 (N_1658,N_1230,N_1483);
nor U1659 (N_1659,N_1463,N_1205);
nor U1660 (N_1660,N_1266,N_1496);
nor U1661 (N_1661,N_1343,N_1388);
and U1662 (N_1662,N_1482,N_1425);
nor U1663 (N_1663,N_1356,N_1258);
xor U1664 (N_1664,N_1189,N_1249);
xor U1665 (N_1665,N_1268,N_1190);
nand U1666 (N_1666,N_1103,N_1385);
nand U1667 (N_1667,N_1422,N_1194);
xor U1668 (N_1668,N_1255,N_1473);
xor U1669 (N_1669,N_1257,N_1490);
xor U1670 (N_1670,N_1429,N_1437);
nand U1671 (N_1671,N_1139,N_1147);
xnor U1672 (N_1672,N_1336,N_1179);
xor U1673 (N_1673,N_1225,N_1227);
nand U1674 (N_1674,N_1273,N_1076);
nor U1675 (N_1675,N_1049,N_1322);
nand U1676 (N_1676,N_1209,N_1440);
xor U1677 (N_1677,N_1303,N_1110);
xnor U1678 (N_1678,N_1202,N_1271);
nor U1679 (N_1679,N_1495,N_1364);
or U1680 (N_1680,N_1231,N_1379);
nor U1681 (N_1681,N_1186,N_1484);
nand U1682 (N_1682,N_1113,N_1441);
and U1683 (N_1683,N_1206,N_1136);
xnor U1684 (N_1684,N_1065,N_1077);
xnor U1685 (N_1685,N_1134,N_1234);
or U1686 (N_1686,N_1238,N_1318);
and U1687 (N_1687,N_1260,N_1165);
nor U1688 (N_1688,N_1416,N_1059);
xor U1689 (N_1689,N_1007,N_1468);
or U1690 (N_1690,N_1132,N_1164);
nor U1691 (N_1691,N_1321,N_1446);
and U1692 (N_1692,N_1340,N_1058);
or U1693 (N_1693,N_1193,N_1218);
nand U1694 (N_1694,N_1011,N_1481);
nand U1695 (N_1695,N_1287,N_1476);
or U1696 (N_1696,N_1156,N_1021);
xor U1697 (N_1697,N_1394,N_1044);
nand U1698 (N_1698,N_1180,N_1277);
or U1699 (N_1699,N_1015,N_1450);
and U1700 (N_1700,N_1171,N_1470);
nor U1701 (N_1701,N_1201,N_1233);
nand U1702 (N_1702,N_1415,N_1080);
nand U1703 (N_1703,N_1370,N_1054);
nand U1704 (N_1704,N_1286,N_1013);
xnor U1705 (N_1705,N_1403,N_1378);
or U1706 (N_1706,N_1263,N_1219);
nand U1707 (N_1707,N_1112,N_1293);
xnor U1708 (N_1708,N_1101,N_1117);
xnor U1709 (N_1709,N_1393,N_1443);
nor U1710 (N_1710,N_1235,N_1386);
nand U1711 (N_1711,N_1436,N_1207);
or U1712 (N_1712,N_1387,N_1239);
and U1713 (N_1713,N_1360,N_1479);
nand U1714 (N_1714,N_1354,N_1439);
and U1715 (N_1715,N_1333,N_1240);
or U1716 (N_1716,N_1372,N_1063);
or U1717 (N_1717,N_1431,N_1084);
or U1718 (N_1718,N_1162,N_1338);
xor U1719 (N_1719,N_1024,N_1167);
xor U1720 (N_1720,N_1125,N_1262);
nor U1721 (N_1721,N_1324,N_1149);
xor U1722 (N_1722,N_1041,N_1319);
xor U1723 (N_1723,N_1159,N_1346);
xor U1724 (N_1724,N_1146,N_1460);
or U1725 (N_1725,N_1081,N_1107);
nor U1726 (N_1726,N_1093,N_1161);
and U1727 (N_1727,N_1434,N_1244);
or U1728 (N_1728,N_1212,N_1073);
xnor U1729 (N_1729,N_1312,N_1276);
nand U1730 (N_1730,N_1308,N_1229);
or U1731 (N_1731,N_1252,N_1469);
or U1732 (N_1732,N_1095,N_1118);
nor U1733 (N_1733,N_1296,N_1304);
nand U1734 (N_1734,N_1306,N_1168);
nor U1735 (N_1735,N_1248,N_1018);
nand U1736 (N_1736,N_1417,N_1042);
nor U1737 (N_1737,N_1160,N_1228);
and U1738 (N_1738,N_1157,N_1242);
xnor U1739 (N_1739,N_1182,N_1017);
nor U1740 (N_1740,N_1305,N_1456);
xnor U1741 (N_1741,N_1111,N_1351);
or U1742 (N_1742,N_1003,N_1199);
xor U1743 (N_1743,N_1020,N_1083);
nand U1744 (N_1744,N_1310,N_1285);
xor U1745 (N_1745,N_1299,N_1368);
xor U1746 (N_1746,N_1369,N_1184);
nor U1747 (N_1747,N_1032,N_1074);
xor U1748 (N_1748,N_1459,N_1152);
or U1749 (N_1749,N_1127,N_1210);
or U1750 (N_1750,N_1048,N_1449);
xnor U1751 (N_1751,N_1211,N_1099);
or U1752 (N_1752,N_1462,N_1040);
nor U1753 (N_1753,N_1423,N_1203);
or U1754 (N_1754,N_1448,N_1455);
and U1755 (N_1755,N_1442,N_1441);
or U1756 (N_1756,N_1456,N_1242);
xnor U1757 (N_1757,N_1106,N_1439);
nor U1758 (N_1758,N_1435,N_1253);
nand U1759 (N_1759,N_1322,N_1005);
or U1760 (N_1760,N_1332,N_1259);
nand U1761 (N_1761,N_1319,N_1385);
nand U1762 (N_1762,N_1118,N_1247);
and U1763 (N_1763,N_1008,N_1190);
xor U1764 (N_1764,N_1192,N_1126);
nand U1765 (N_1765,N_1026,N_1269);
and U1766 (N_1766,N_1482,N_1018);
xnor U1767 (N_1767,N_1488,N_1448);
and U1768 (N_1768,N_1489,N_1389);
nor U1769 (N_1769,N_1244,N_1287);
and U1770 (N_1770,N_1453,N_1096);
nor U1771 (N_1771,N_1143,N_1342);
nand U1772 (N_1772,N_1052,N_1464);
nor U1773 (N_1773,N_1274,N_1462);
nor U1774 (N_1774,N_1400,N_1392);
xnor U1775 (N_1775,N_1362,N_1120);
and U1776 (N_1776,N_1353,N_1073);
or U1777 (N_1777,N_1119,N_1419);
and U1778 (N_1778,N_1095,N_1316);
xnor U1779 (N_1779,N_1159,N_1428);
and U1780 (N_1780,N_1043,N_1446);
nand U1781 (N_1781,N_1093,N_1309);
nor U1782 (N_1782,N_1016,N_1346);
and U1783 (N_1783,N_1172,N_1299);
or U1784 (N_1784,N_1033,N_1499);
or U1785 (N_1785,N_1366,N_1022);
and U1786 (N_1786,N_1064,N_1492);
and U1787 (N_1787,N_1420,N_1220);
nand U1788 (N_1788,N_1380,N_1387);
nor U1789 (N_1789,N_1353,N_1345);
nor U1790 (N_1790,N_1352,N_1220);
and U1791 (N_1791,N_1217,N_1122);
xnor U1792 (N_1792,N_1403,N_1274);
and U1793 (N_1793,N_1245,N_1480);
xor U1794 (N_1794,N_1027,N_1013);
xor U1795 (N_1795,N_1006,N_1098);
nand U1796 (N_1796,N_1356,N_1465);
or U1797 (N_1797,N_1240,N_1303);
and U1798 (N_1798,N_1112,N_1189);
nor U1799 (N_1799,N_1058,N_1345);
xor U1800 (N_1800,N_1166,N_1382);
nor U1801 (N_1801,N_1432,N_1136);
and U1802 (N_1802,N_1281,N_1387);
nand U1803 (N_1803,N_1363,N_1047);
and U1804 (N_1804,N_1237,N_1021);
nor U1805 (N_1805,N_1269,N_1186);
or U1806 (N_1806,N_1272,N_1418);
xnor U1807 (N_1807,N_1306,N_1130);
or U1808 (N_1808,N_1064,N_1149);
or U1809 (N_1809,N_1210,N_1163);
xnor U1810 (N_1810,N_1151,N_1000);
nand U1811 (N_1811,N_1268,N_1160);
nor U1812 (N_1812,N_1041,N_1358);
nor U1813 (N_1813,N_1349,N_1308);
nand U1814 (N_1814,N_1056,N_1010);
nand U1815 (N_1815,N_1133,N_1441);
and U1816 (N_1816,N_1302,N_1115);
and U1817 (N_1817,N_1345,N_1303);
and U1818 (N_1818,N_1435,N_1088);
nor U1819 (N_1819,N_1309,N_1072);
or U1820 (N_1820,N_1482,N_1476);
nor U1821 (N_1821,N_1227,N_1212);
or U1822 (N_1822,N_1207,N_1021);
and U1823 (N_1823,N_1209,N_1462);
and U1824 (N_1824,N_1085,N_1123);
and U1825 (N_1825,N_1045,N_1403);
nand U1826 (N_1826,N_1407,N_1298);
xnor U1827 (N_1827,N_1318,N_1050);
nor U1828 (N_1828,N_1159,N_1239);
nor U1829 (N_1829,N_1378,N_1155);
nand U1830 (N_1830,N_1372,N_1446);
xnor U1831 (N_1831,N_1401,N_1489);
xor U1832 (N_1832,N_1385,N_1099);
nand U1833 (N_1833,N_1423,N_1432);
nand U1834 (N_1834,N_1353,N_1282);
xor U1835 (N_1835,N_1371,N_1447);
and U1836 (N_1836,N_1308,N_1224);
or U1837 (N_1837,N_1273,N_1326);
or U1838 (N_1838,N_1469,N_1273);
nand U1839 (N_1839,N_1113,N_1170);
xnor U1840 (N_1840,N_1499,N_1089);
nor U1841 (N_1841,N_1266,N_1078);
xor U1842 (N_1842,N_1032,N_1439);
or U1843 (N_1843,N_1372,N_1433);
and U1844 (N_1844,N_1391,N_1246);
or U1845 (N_1845,N_1250,N_1295);
or U1846 (N_1846,N_1199,N_1095);
nand U1847 (N_1847,N_1386,N_1186);
xnor U1848 (N_1848,N_1122,N_1114);
or U1849 (N_1849,N_1006,N_1309);
nor U1850 (N_1850,N_1051,N_1480);
nor U1851 (N_1851,N_1354,N_1436);
and U1852 (N_1852,N_1037,N_1389);
nor U1853 (N_1853,N_1223,N_1450);
nand U1854 (N_1854,N_1188,N_1443);
nor U1855 (N_1855,N_1017,N_1103);
or U1856 (N_1856,N_1394,N_1123);
xnor U1857 (N_1857,N_1391,N_1008);
nor U1858 (N_1858,N_1381,N_1298);
or U1859 (N_1859,N_1327,N_1436);
nor U1860 (N_1860,N_1339,N_1267);
and U1861 (N_1861,N_1262,N_1110);
and U1862 (N_1862,N_1302,N_1483);
xnor U1863 (N_1863,N_1331,N_1221);
xor U1864 (N_1864,N_1437,N_1185);
nor U1865 (N_1865,N_1378,N_1094);
xnor U1866 (N_1866,N_1384,N_1036);
nand U1867 (N_1867,N_1099,N_1220);
xnor U1868 (N_1868,N_1293,N_1130);
nor U1869 (N_1869,N_1222,N_1253);
xnor U1870 (N_1870,N_1009,N_1440);
xnor U1871 (N_1871,N_1214,N_1386);
nor U1872 (N_1872,N_1430,N_1266);
or U1873 (N_1873,N_1412,N_1013);
and U1874 (N_1874,N_1375,N_1451);
nor U1875 (N_1875,N_1084,N_1372);
or U1876 (N_1876,N_1074,N_1300);
nor U1877 (N_1877,N_1251,N_1123);
nand U1878 (N_1878,N_1365,N_1267);
or U1879 (N_1879,N_1028,N_1424);
or U1880 (N_1880,N_1000,N_1232);
or U1881 (N_1881,N_1352,N_1347);
xor U1882 (N_1882,N_1128,N_1251);
or U1883 (N_1883,N_1351,N_1459);
or U1884 (N_1884,N_1449,N_1235);
xnor U1885 (N_1885,N_1309,N_1389);
xnor U1886 (N_1886,N_1047,N_1155);
nand U1887 (N_1887,N_1286,N_1447);
xor U1888 (N_1888,N_1453,N_1482);
nor U1889 (N_1889,N_1143,N_1364);
and U1890 (N_1890,N_1359,N_1238);
and U1891 (N_1891,N_1257,N_1187);
nand U1892 (N_1892,N_1000,N_1174);
or U1893 (N_1893,N_1174,N_1215);
and U1894 (N_1894,N_1312,N_1105);
nor U1895 (N_1895,N_1179,N_1499);
nand U1896 (N_1896,N_1233,N_1239);
nand U1897 (N_1897,N_1234,N_1055);
or U1898 (N_1898,N_1207,N_1294);
and U1899 (N_1899,N_1480,N_1304);
or U1900 (N_1900,N_1239,N_1083);
and U1901 (N_1901,N_1048,N_1010);
nand U1902 (N_1902,N_1382,N_1296);
and U1903 (N_1903,N_1159,N_1453);
and U1904 (N_1904,N_1327,N_1263);
nand U1905 (N_1905,N_1070,N_1324);
or U1906 (N_1906,N_1421,N_1218);
or U1907 (N_1907,N_1348,N_1357);
nand U1908 (N_1908,N_1248,N_1229);
nand U1909 (N_1909,N_1174,N_1071);
nor U1910 (N_1910,N_1277,N_1407);
nor U1911 (N_1911,N_1482,N_1286);
nor U1912 (N_1912,N_1108,N_1358);
xor U1913 (N_1913,N_1059,N_1141);
nor U1914 (N_1914,N_1465,N_1194);
and U1915 (N_1915,N_1064,N_1281);
and U1916 (N_1916,N_1026,N_1159);
or U1917 (N_1917,N_1284,N_1173);
nor U1918 (N_1918,N_1309,N_1376);
or U1919 (N_1919,N_1420,N_1124);
or U1920 (N_1920,N_1402,N_1093);
and U1921 (N_1921,N_1380,N_1039);
xnor U1922 (N_1922,N_1481,N_1092);
xnor U1923 (N_1923,N_1305,N_1333);
nand U1924 (N_1924,N_1155,N_1112);
and U1925 (N_1925,N_1153,N_1028);
or U1926 (N_1926,N_1381,N_1492);
nor U1927 (N_1927,N_1267,N_1476);
nor U1928 (N_1928,N_1148,N_1141);
nand U1929 (N_1929,N_1488,N_1383);
xnor U1930 (N_1930,N_1358,N_1091);
and U1931 (N_1931,N_1385,N_1175);
or U1932 (N_1932,N_1258,N_1048);
nand U1933 (N_1933,N_1004,N_1093);
and U1934 (N_1934,N_1224,N_1067);
nand U1935 (N_1935,N_1357,N_1453);
xnor U1936 (N_1936,N_1173,N_1456);
xnor U1937 (N_1937,N_1032,N_1169);
xor U1938 (N_1938,N_1314,N_1375);
nor U1939 (N_1939,N_1468,N_1427);
nand U1940 (N_1940,N_1460,N_1289);
and U1941 (N_1941,N_1384,N_1119);
xor U1942 (N_1942,N_1203,N_1373);
xor U1943 (N_1943,N_1157,N_1159);
xor U1944 (N_1944,N_1099,N_1484);
or U1945 (N_1945,N_1081,N_1466);
nor U1946 (N_1946,N_1114,N_1382);
nor U1947 (N_1947,N_1307,N_1349);
and U1948 (N_1948,N_1251,N_1146);
nand U1949 (N_1949,N_1418,N_1385);
and U1950 (N_1950,N_1427,N_1083);
nand U1951 (N_1951,N_1391,N_1245);
nand U1952 (N_1952,N_1085,N_1178);
nor U1953 (N_1953,N_1188,N_1147);
nand U1954 (N_1954,N_1495,N_1422);
xnor U1955 (N_1955,N_1141,N_1137);
nand U1956 (N_1956,N_1196,N_1193);
nor U1957 (N_1957,N_1391,N_1077);
and U1958 (N_1958,N_1116,N_1046);
and U1959 (N_1959,N_1309,N_1065);
xnor U1960 (N_1960,N_1482,N_1185);
xnor U1961 (N_1961,N_1198,N_1106);
or U1962 (N_1962,N_1357,N_1067);
nand U1963 (N_1963,N_1218,N_1220);
nand U1964 (N_1964,N_1320,N_1405);
nand U1965 (N_1965,N_1356,N_1246);
nor U1966 (N_1966,N_1481,N_1396);
and U1967 (N_1967,N_1389,N_1163);
nand U1968 (N_1968,N_1262,N_1374);
or U1969 (N_1969,N_1318,N_1495);
nor U1970 (N_1970,N_1221,N_1499);
nand U1971 (N_1971,N_1445,N_1164);
nor U1972 (N_1972,N_1064,N_1396);
or U1973 (N_1973,N_1299,N_1220);
xnor U1974 (N_1974,N_1229,N_1483);
xnor U1975 (N_1975,N_1277,N_1274);
xnor U1976 (N_1976,N_1036,N_1046);
xor U1977 (N_1977,N_1427,N_1002);
nand U1978 (N_1978,N_1009,N_1256);
xor U1979 (N_1979,N_1241,N_1038);
and U1980 (N_1980,N_1262,N_1360);
nand U1981 (N_1981,N_1079,N_1052);
or U1982 (N_1982,N_1070,N_1338);
or U1983 (N_1983,N_1290,N_1236);
nand U1984 (N_1984,N_1022,N_1176);
and U1985 (N_1985,N_1175,N_1215);
nand U1986 (N_1986,N_1182,N_1245);
xnor U1987 (N_1987,N_1094,N_1388);
nand U1988 (N_1988,N_1079,N_1473);
xor U1989 (N_1989,N_1403,N_1019);
nor U1990 (N_1990,N_1221,N_1281);
and U1991 (N_1991,N_1258,N_1016);
and U1992 (N_1992,N_1140,N_1028);
and U1993 (N_1993,N_1326,N_1442);
xor U1994 (N_1994,N_1036,N_1070);
or U1995 (N_1995,N_1230,N_1257);
and U1996 (N_1996,N_1377,N_1030);
or U1997 (N_1997,N_1356,N_1034);
nor U1998 (N_1998,N_1268,N_1263);
xnor U1999 (N_1999,N_1471,N_1336);
and U2000 (N_2000,N_1908,N_1988);
nor U2001 (N_2001,N_1858,N_1731);
and U2002 (N_2002,N_1693,N_1957);
xor U2003 (N_2003,N_1742,N_1572);
or U2004 (N_2004,N_1932,N_1897);
nand U2005 (N_2005,N_1788,N_1822);
nor U2006 (N_2006,N_1717,N_1582);
nor U2007 (N_2007,N_1749,N_1698);
nor U2008 (N_2008,N_1782,N_1548);
or U2009 (N_2009,N_1661,N_1672);
nor U2010 (N_2010,N_1707,N_1701);
nor U2011 (N_2011,N_1947,N_1839);
nand U2012 (N_2012,N_1571,N_1600);
and U2013 (N_2013,N_1654,N_1724);
and U2014 (N_2014,N_1870,N_1502);
nor U2015 (N_2015,N_1627,N_1781);
nor U2016 (N_2016,N_1877,N_1635);
nor U2017 (N_2017,N_1694,N_1990);
nor U2018 (N_2018,N_1629,N_1823);
and U2019 (N_2019,N_1562,N_1676);
or U2020 (N_2020,N_1843,N_1609);
and U2021 (N_2021,N_1765,N_1856);
nand U2022 (N_2022,N_1678,N_1533);
and U2023 (N_2023,N_1814,N_1682);
nand U2024 (N_2024,N_1828,N_1993);
nand U2025 (N_2025,N_1518,N_1515);
nor U2026 (N_2026,N_1683,N_1720);
and U2027 (N_2027,N_1784,N_1697);
and U2028 (N_2028,N_1962,N_1913);
nand U2029 (N_2029,N_1702,N_1555);
and U2030 (N_2030,N_1653,N_1973);
nand U2031 (N_2031,N_1815,N_1535);
or U2032 (N_2032,N_1968,N_1700);
and U2033 (N_2033,N_1925,N_1873);
nor U2034 (N_2034,N_1736,N_1779);
and U2035 (N_2035,N_1588,N_1774);
and U2036 (N_2036,N_1639,N_1912);
xnor U2037 (N_2037,N_1622,N_1597);
xnor U2038 (N_2038,N_1705,N_1921);
xnor U2039 (N_2039,N_1744,N_1785);
and U2040 (N_2040,N_1824,N_1794);
nor U2041 (N_2041,N_1630,N_1687);
or U2042 (N_2042,N_1837,N_1586);
nand U2043 (N_2043,N_1941,N_1906);
xnor U2044 (N_2044,N_1650,N_1699);
and U2045 (N_2045,N_1849,N_1671);
nand U2046 (N_2046,N_1505,N_1916);
and U2047 (N_2047,N_1902,N_1714);
or U2048 (N_2048,N_1624,N_1611);
or U2049 (N_2049,N_1727,N_1884);
xnor U2050 (N_2050,N_1734,N_1549);
and U2051 (N_2051,N_1748,N_1959);
xor U2052 (N_2052,N_1660,N_1580);
nand U2053 (N_2053,N_1532,N_1751);
or U2054 (N_2054,N_1547,N_1799);
and U2055 (N_2055,N_1704,N_1722);
xnor U2056 (N_2056,N_1918,N_1716);
nor U2057 (N_2057,N_1718,N_1613);
or U2058 (N_2058,N_1934,N_1960);
xnor U2059 (N_2059,N_1541,N_1768);
and U2060 (N_2060,N_1787,N_1521);
nand U2061 (N_2061,N_1556,N_1667);
nand U2062 (N_2062,N_1776,N_1589);
xor U2063 (N_2063,N_1816,N_1999);
xnor U2064 (N_2064,N_1989,N_1735);
xnor U2065 (N_2065,N_1965,N_1692);
or U2066 (N_2066,N_1543,N_1685);
xor U2067 (N_2067,N_1967,N_1775);
nand U2068 (N_2068,N_1830,N_1504);
nand U2069 (N_2069,N_1848,N_1576);
and U2070 (N_2070,N_1590,N_1542);
nand U2071 (N_2071,N_1806,N_1778);
nor U2072 (N_2072,N_1938,N_1651);
xnor U2073 (N_2073,N_1979,N_1537);
nor U2074 (N_2074,N_1844,N_1710);
and U2075 (N_2075,N_1869,N_1767);
and U2076 (N_2076,N_1757,N_1804);
and U2077 (N_2077,N_1610,N_1991);
nor U2078 (N_2078,N_1866,N_1706);
or U2079 (N_2079,N_1636,N_1675);
xor U2080 (N_2080,N_1620,N_1560);
xor U2081 (N_2081,N_1838,N_1516);
or U2082 (N_2082,N_1669,N_1577);
nand U2083 (N_2083,N_1551,N_1644);
xor U2084 (N_2084,N_1926,N_1570);
nand U2085 (N_2085,N_1893,N_1786);
nand U2086 (N_2086,N_1500,N_1587);
xnor U2087 (N_2087,N_1688,N_1859);
nor U2088 (N_2088,N_1553,N_1833);
nor U2089 (N_2089,N_1637,N_1602);
and U2090 (N_2090,N_1910,N_1796);
and U2091 (N_2091,N_1840,N_1759);
and U2092 (N_2092,N_1743,N_1691);
nor U2093 (N_2093,N_1545,N_1561);
xor U2094 (N_2094,N_1880,N_1845);
or U2095 (N_2095,N_1964,N_1997);
nor U2096 (N_2096,N_1819,N_1566);
or U2097 (N_2097,N_1987,N_1770);
xor U2098 (N_2098,N_1857,N_1758);
nor U2099 (N_2099,N_1747,N_1812);
nand U2100 (N_2100,N_1657,N_1821);
nand U2101 (N_2101,N_1971,N_1604);
nor U2102 (N_2102,N_1852,N_1829);
nand U2103 (N_2103,N_1865,N_1656);
or U2104 (N_2104,N_1998,N_1511);
xor U2105 (N_2105,N_1876,N_1595);
nand U2106 (N_2106,N_1575,N_1649);
nor U2107 (N_2107,N_1746,N_1861);
nor U2108 (N_2108,N_1867,N_1536);
or U2109 (N_2109,N_1899,N_1510);
xor U2110 (N_2110,N_1646,N_1801);
nand U2111 (N_2111,N_1820,N_1726);
xor U2112 (N_2112,N_1593,N_1922);
and U2113 (N_2113,N_1777,N_1733);
xnor U2114 (N_2114,N_1937,N_1623);
and U2115 (N_2115,N_1970,N_1855);
nor U2116 (N_2116,N_1780,N_1573);
nor U2117 (N_2117,N_1550,N_1728);
nor U2118 (N_2118,N_1607,N_1984);
xnor U2119 (N_2119,N_1567,N_1557);
nand U2120 (N_2120,N_1591,N_1860);
nand U2121 (N_2121,N_1885,N_1565);
and U2122 (N_2122,N_1889,N_1836);
nand U2123 (N_2123,N_1948,N_1863);
nand U2124 (N_2124,N_1883,N_1868);
nand U2125 (N_2125,N_1696,N_1841);
nand U2126 (N_2126,N_1642,N_1558);
and U2127 (N_2127,N_1513,N_1723);
xor U2128 (N_2128,N_1559,N_1983);
and U2129 (N_2129,N_1544,N_1955);
xor U2130 (N_2130,N_1772,N_1529);
nand U2131 (N_2131,N_1752,N_1679);
xor U2132 (N_2132,N_1626,N_1802);
or U2133 (N_2133,N_1929,N_1940);
xnor U2134 (N_2134,N_1753,N_1755);
xor U2135 (N_2135,N_1882,N_1892);
nand U2136 (N_2136,N_1583,N_1891);
and U2137 (N_2137,N_1878,N_1632);
nor U2138 (N_2138,N_1517,N_1879);
nor U2139 (N_2139,N_1818,N_1638);
and U2140 (N_2140,N_1578,N_1931);
or U2141 (N_2141,N_1564,N_1825);
xnor U2142 (N_2142,N_1581,N_1608);
and U2143 (N_2143,N_1975,N_1506);
xnor U2144 (N_2144,N_1648,N_1729);
xor U2145 (N_2145,N_1905,N_1792);
nor U2146 (N_2146,N_1956,N_1641);
or U2147 (N_2147,N_1862,N_1842);
and U2148 (N_2148,N_1834,N_1605);
nand U2149 (N_2149,N_1616,N_1982);
nor U2150 (N_2150,N_1614,N_1503);
nor U2151 (N_2151,N_1871,N_1737);
xnor U2152 (N_2152,N_1526,N_1509);
or U2153 (N_2153,N_1994,N_1663);
or U2154 (N_2154,N_1942,N_1766);
nor U2155 (N_2155,N_1914,N_1986);
or U2156 (N_2156,N_1810,N_1527);
and U2157 (N_2157,N_1946,N_1789);
or U2158 (N_2158,N_1647,N_1917);
xor U2159 (N_2159,N_1612,N_1514);
nor U2160 (N_2160,N_1945,N_1674);
nor U2161 (N_2161,N_1813,N_1793);
or U2162 (N_2162,N_1992,N_1708);
nor U2163 (N_2163,N_1525,N_1546);
and U2164 (N_2164,N_1936,N_1769);
and U2165 (N_2165,N_1596,N_1520);
nand U2166 (N_2166,N_1668,N_1740);
nor U2167 (N_2167,N_1713,N_1930);
nand U2168 (N_2168,N_1904,N_1978);
and U2169 (N_2169,N_1935,N_1750);
nand U2170 (N_2170,N_1985,N_1763);
and U2171 (N_2171,N_1976,N_1501);
and U2172 (N_2172,N_1850,N_1530);
and U2173 (N_2173,N_1640,N_1915);
or U2174 (N_2174,N_1958,N_1835);
nor U2175 (N_2175,N_1584,N_1592);
and U2176 (N_2176,N_1508,N_1771);
nand U2177 (N_2177,N_1563,N_1528);
nand U2178 (N_2178,N_1911,N_1606);
and U2179 (N_2179,N_1795,N_1791);
and U2180 (N_2180,N_1898,N_1888);
xnor U2181 (N_2181,N_1534,N_1619);
and U2182 (N_2182,N_1895,N_1598);
nand U2183 (N_2183,N_1659,N_1631);
or U2184 (N_2184,N_1670,N_1618);
nand U2185 (N_2185,N_1512,N_1761);
nand U2186 (N_2186,N_1800,N_1864);
xnor U2187 (N_2187,N_1754,N_1603);
or U2188 (N_2188,N_1625,N_1980);
nor U2189 (N_2189,N_1797,N_1943);
or U2190 (N_2190,N_1643,N_1507);
or U2191 (N_2191,N_1522,N_1540);
nand U2192 (N_2192,N_1617,N_1949);
xnor U2193 (N_2193,N_1923,N_1805);
or U2194 (N_2194,N_1809,N_1851);
nand U2195 (N_2195,N_1712,N_1756);
nor U2196 (N_2196,N_1519,N_1826);
nand U2197 (N_2197,N_1677,N_1933);
and U2198 (N_2198,N_1939,N_1601);
nand U2199 (N_2199,N_1741,N_1539);
nand U2200 (N_2200,N_1621,N_1554);
and U2201 (N_2201,N_1599,N_1924);
nand U2202 (N_2202,N_1531,N_1961);
xor U2203 (N_2203,N_1974,N_1645);
xnor U2204 (N_2204,N_1725,N_1886);
xor U2205 (N_2205,N_1711,N_1523);
or U2206 (N_2206,N_1538,N_1881);
nor U2207 (N_2207,N_1690,N_1745);
or U2208 (N_2208,N_1944,N_1954);
or U2209 (N_2209,N_1633,N_1890);
nor U2210 (N_2210,N_1739,N_1783);
xor U2211 (N_2211,N_1634,N_1903);
or U2212 (N_2212,N_1807,N_1664);
xnor U2213 (N_2213,N_1853,N_1875);
and U2214 (N_2214,N_1798,N_1615);
and U2215 (N_2215,N_1966,N_1662);
and U2216 (N_2216,N_1673,N_1680);
and U2217 (N_2217,N_1977,N_1665);
or U2218 (N_2218,N_1569,N_1574);
nor U2219 (N_2219,N_1817,N_1831);
or U2220 (N_2220,N_1658,N_1928);
nand U2221 (N_2221,N_1764,N_1951);
or U2222 (N_2222,N_1773,N_1684);
nor U2223 (N_2223,N_1681,N_1594);
or U2224 (N_2224,N_1666,N_1950);
and U2225 (N_2225,N_1832,N_1920);
xnor U2226 (N_2226,N_1995,N_1900);
nand U2227 (N_2227,N_1887,N_1568);
and U2228 (N_2228,N_1703,N_1732);
xnor U2229 (N_2229,N_1846,N_1709);
xnor U2230 (N_2230,N_1803,N_1715);
nor U2231 (N_2231,N_1969,N_1827);
nor U2232 (N_2232,N_1909,N_1963);
xnor U2233 (N_2233,N_1907,N_1730);
xor U2234 (N_2234,N_1972,N_1981);
or U2235 (N_2235,N_1952,N_1896);
nand U2236 (N_2236,N_1790,N_1872);
xnor U2237 (N_2237,N_1689,N_1524);
or U2238 (N_2238,N_1953,N_1579);
nor U2239 (N_2239,N_1552,N_1854);
nor U2240 (N_2240,N_1927,N_1894);
or U2241 (N_2241,N_1808,N_1721);
xor U2242 (N_2242,N_1760,N_1686);
nand U2243 (N_2243,N_1652,N_1655);
and U2244 (N_2244,N_1919,N_1762);
nor U2245 (N_2245,N_1847,N_1738);
and U2246 (N_2246,N_1901,N_1695);
nand U2247 (N_2247,N_1628,N_1874);
and U2248 (N_2248,N_1719,N_1996);
nor U2249 (N_2249,N_1585,N_1811);
or U2250 (N_2250,N_1610,N_1611);
nand U2251 (N_2251,N_1581,N_1573);
xnor U2252 (N_2252,N_1762,N_1837);
xnor U2253 (N_2253,N_1861,N_1988);
xor U2254 (N_2254,N_1868,N_1673);
nand U2255 (N_2255,N_1906,N_1618);
or U2256 (N_2256,N_1915,N_1655);
nor U2257 (N_2257,N_1542,N_1963);
nand U2258 (N_2258,N_1758,N_1739);
or U2259 (N_2259,N_1643,N_1773);
and U2260 (N_2260,N_1998,N_1938);
nor U2261 (N_2261,N_1900,N_1991);
nor U2262 (N_2262,N_1558,N_1532);
or U2263 (N_2263,N_1780,N_1713);
and U2264 (N_2264,N_1872,N_1697);
xor U2265 (N_2265,N_1790,N_1674);
nor U2266 (N_2266,N_1623,N_1943);
and U2267 (N_2267,N_1599,N_1995);
and U2268 (N_2268,N_1502,N_1721);
nand U2269 (N_2269,N_1905,N_1778);
nor U2270 (N_2270,N_1991,N_1683);
xnor U2271 (N_2271,N_1646,N_1766);
xnor U2272 (N_2272,N_1525,N_1855);
nand U2273 (N_2273,N_1956,N_1795);
and U2274 (N_2274,N_1860,N_1611);
or U2275 (N_2275,N_1983,N_1696);
and U2276 (N_2276,N_1945,N_1931);
nor U2277 (N_2277,N_1758,N_1801);
nand U2278 (N_2278,N_1914,N_1623);
and U2279 (N_2279,N_1842,N_1942);
nand U2280 (N_2280,N_1760,N_1511);
nor U2281 (N_2281,N_1510,N_1784);
nor U2282 (N_2282,N_1898,N_1974);
or U2283 (N_2283,N_1871,N_1785);
xor U2284 (N_2284,N_1870,N_1624);
and U2285 (N_2285,N_1531,N_1515);
and U2286 (N_2286,N_1855,N_1725);
and U2287 (N_2287,N_1531,N_1633);
xor U2288 (N_2288,N_1895,N_1968);
and U2289 (N_2289,N_1814,N_1846);
or U2290 (N_2290,N_1832,N_1511);
nand U2291 (N_2291,N_1961,N_1850);
xnor U2292 (N_2292,N_1725,N_1787);
and U2293 (N_2293,N_1586,N_1928);
and U2294 (N_2294,N_1550,N_1750);
and U2295 (N_2295,N_1747,N_1867);
or U2296 (N_2296,N_1858,N_1617);
xnor U2297 (N_2297,N_1877,N_1805);
and U2298 (N_2298,N_1766,N_1909);
nor U2299 (N_2299,N_1538,N_1895);
and U2300 (N_2300,N_1535,N_1921);
nand U2301 (N_2301,N_1950,N_1686);
nand U2302 (N_2302,N_1799,N_1809);
or U2303 (N_2303,N_1548,N_1681);
and U2304 (N_2304,N_1930,N_1521);
xnor U2305 (N_2305,N_1936,N_1964);
nand U2306 (N_2306,N_1995,N_1606);
nand U2307 (N_2307,N_1718,N_1668);
nor U2308 (N_2308,N_1840,N_1658);
and U2309 (N_2309,N_1998,N_1508);
nand U2310 (N_2310,N_1655,N_1697);
nand U2311 (N_2311,N_1540,N_1754);
and U2312 (N_2312,N_1921,N_1910);
nand U2313 (N_2313,N_1917,N_1757);
nand U2314 (N_2314,N_1818,N_1786);
xnor U2315 (N_2315,N_1590,N_1743);
and U2316 (N_2316,N_1619,N_1790);
and U2317 (N_2317,N_1795,N_1675);
or U2318 (N_2318,N_1658,N_1918);
xor U2319 (N_2319,N_1918,N_1730);
xor U2320 (N_2320,N_1830,N_1578);
nor U2321 (N_2321,N_1888,N_1846);
and U2322 (N_2322,N_1522,N_1609);
and U2323 (N_2323,N_1549,N_1724);
xnor U2324 (N_2324,N_1588,N_1931);
xnor U2325 (N_2325,N_1583,N_1995);
nand U2326 (N_2326,N_1667,N_1649);
and U2327 (N_2327,N_1806,N_1545);
and U2328 (N_2328,N_1886,N_1608);
nor U2329 (N_2329,N_1955,N_1761);
xor U2330 (N_2330,N_1901,N_1606);
nor U2331 (N_2331,N_1679,N_1758);
and U2332 (N_2332,N_1507,N_1575);
xor U2333 (N_2333,N_1769,N_1684);
xor U2334 (N_2334,N_1952,N_1631);
nor U2335 (N_2335,N_1986,N_1558);
or U2336 (N_2336,N_1858,N_1862);
nand U2337 (N_2337,N_1627,N_1795);
and U2338 (N_2338,N_1936,N_1801);
xor U2339 (N_2339,N_1902,N_1992);
nand U2340 (N_2340,N_1965,N_1925);
nor U2341 (N_2341,N_1938,N_1747);
xnor U2342 (N_2342,N_1874,N_1797);
xnor U2343 (N_2343,N_1731,N_1541);
or U2344 (N_2344,N_1568,N_1861);
or U2345 (N_2345,N_1689,N_1751);
or U2346 (N_2346,N_1789,N_1636);
and U2347 (N_2347,N_1624,N_1538);
and U2348 (N_2348,N_1707,N_1991);
nor U2349 (N_2349,N_1835,N_1853);
and U2350 (N_2350,N_1780,N_1567);
or U2351 (N_2351,N_1543,N_1863);
and U2352 (N_2352,N_1552,N_1991);
or U2353 (N_2353,N_1631,N_1988);
nand U2354 (N_2354,N_1761,N_1827);
nor U2355 (N_2355,N_1590,N_1551);
nor U2356 (N_2356,N_1784,N_1563);
or U2357 (N_2357,N_1659,N_1892);
or U2358 (N_2358,N_1752,N_1503);
and U2359 (N_2359,N_1671,N_1638);
nand U2360 (N_2360,N_1650,N_1705);
nand U2361 (N_2361,N_1979,N_1843);
or U2362 (N_2362,N_1502,N_1557);
xor U2363 (N_2363,N_1979,N_1828);
nor U2364 (N_2364,N_1797,N_1635);
nand U2365 (N_2365,N_1715,N_1750);
or U2366 (N_2366,N_1822,N_1979);
and U2367 (N_2367,N_1557,N_1602);
xor U2368 (N_2368,N_1786,N_1505);
xor U2369 (N_2369,N_1668,N_1633);
or U2370 (N_2370,N_1580,N_1865);
and U2371 (N_2371,N_1510,N_1922);
xor U2372 (N_2372,N_1666,N_1725);
nor U2373 (N_2373,N_1675,N_1729);
or U2374 (N_2374,N_1605,N_1789);
or U2375 (N_2375,N_1717,N_1536);
nand U2376 (N_2376,N_1725,N_1844);
nand U2377 (N_2377,N_1677,N_1895);
or U2378 (N_2378,N_1763,N_1731);
and U2379 (N_2379,N_1917,N_1889);
or U2380 (N_2380,N_1629,N_1670);
or U2381 (N_2381,N_1502,N_1712);
xnor U2382 (N_2382,N_1631,N_1814);
or U2383 (N_2383,N_1540,N_1531);
and U2384 (N_2384,N_1857,N_1702);
and U2385 (N_2385,N_1737,N_1675);
xnor U2386 (N_2386,N_1513,N_1632);
nor U2387 (N_2387,N_1722,N_1742);
nor U2388 (N_2388,N_1996,N_1635);
nor U2389 (N_2389,N_1805,N_1958);
nand U2390 (N_2390,N_1842,N_1876);
xnor U2391 (N_2391,N_1877,N_1532);
or U2392 (N_2392,N_1582,N_1644);
nor U2393 (N_2393,N_1972,N_1642);
nor U2394 (N_2394,N_1834,N_1742);
xnor U2395 (N_2395,N_1731,N_1971);
nor U2396 (N_2396,N_1714,N_1875);
or U2397 (N_2397,N_1829,N_1758);
or U2398 (N_2398,N_1895,N_1565);
and U2399 (N_2399,N_1630,N_1740);
and U2400 (N_2400,N_1886,N_1876);
or U2401 (N_2401,N_1815,N_1657);
xnor U2402 (N_2402,N_1988,N_1724);
and U2403 (N_2403,N_1622,N_1731);
and U2404 (N_2404,N_1877,N_1615);
and U2405 (N_2405,N_1852,N_1813);
nor U2406 (N_2406,N_1923,N_1999);
nand U2407 (N_2407,N_1710,N_1741);
xnor U2408 (N_2408,N_1797,N_1815);
and U2409 (N_2409,N_1803,N_1526);
nand U2410 (N_2410,N_1605,N_1568);
nand U2411 (N_2411,N_1528,N_1920);
or U2412 (N_2412,N_1676,N_1882);
and U2413 (N_2413,N_1926,N_1537);
or U2414 (N_2414,N_1514,N_1565);
and U2415 (N_2415,N_1830,N_1827);
and U2416 (N_2416,N_1787,N_1567);
nand U2417 (N_2417,N_1964,N_1959);
and U2418 (N_2418,N_1689,N_1564);
xor U2419 (N_2419,N_1963,N_1510);
nor U2420 (N_2420,N_1786,N_1673);
nand U2421 (N_2421,N_1506,N_1687);
xor U2422 (N_2422,N_1932,N_1589);
or U2423 (N_2423,N_1656,N_1591);
xnor U2424 (N_2424,N_1786,N_1564);
and U2425 (N_2425,N_1946,N_1525);
or U2426 (N_2426,N_1979,N_1819);
nand U2427 (N_2427,N_1573,N_1880);
or U2428 (N_2428,N_1869,N_1979);
and U2429 (N_2429,N_1741,N_1706);
and U2430 (N_2430,N_1559,N_1890);
or U2431 (N_2431,N_1873,N_1780);
nor U2432 (N_2432,N_1732,N_1531);
and U2433 (N_2433,N_1969,N_1953);
nor U2434 (N_2434,N_1995,N_1700);
xor U2435 (N_2435,N_1603,N_1901);
nor U2436 (N_2436,N_1682,N_1741);
nand U2437 (N_2437,N_1837,N_1729);
nand U2438 (N_2438,N_1541,N_1992);
or U2439 (N_2439,N_1601,N_1850);
xnor U2440 (N_2440,N_1516,N_1836);
nand U2441 (N_2441,N_1696,N_1962);
xnor U2442 (N_2442,N_1677,N_1710);
or U2443 (N_2443,N_1579,N_1652);
and U2444 (N_2444,N_1831,N_1736);
and U2445 (N_2445,N_1919,N_1711);
and U2446 (N_2446,N_1867,N_1941);
nor U2447 (N_2447,N_1722,N_1525);
xnor U2448 (N_2448,N_1740,N_1601);
and U2449 (N_2449,N_1702,N_1799);
and U2450 (N_2450,N_1775,N_1764);
or U2451 (N_2451,N_1803,N_1930);
and U2452 (N_2452,N_1714,N_1513);
nor U2453 (N_2453,N_1663,N_1824);
or U2454 (N_2454,N_1883,N_1854);
and U2455 (N_2455,N_1897,N_1631);
and U2456 (N_2456,N_1657,N_1818);
or U2457 (N_2457,N_1736,N_1985);
nand U2458 (N_2458,N_1528,N_1968);
and U2459 (N_2459,N_1887,N_1873);
or U2460 (N_2460,N_1691,N_1617);
nor U2461 (N_2461,N_1678,N_1600);
or U2462 (N_2462,N_1506,N_1832);
or U2463 (N_2463,N_1953,N_1518);
nand U2464 (N_2464,N_1808,N_1922);
nand U2465 (N_2465,N_1552,N_1749);
and U2466 (N_2466,N_1893,N_1711);
and U2467 (N_2467,N_1859,N_1734);
nand U2468 (N_2468,N_1886,N_1541);
nor U2469 (N_2469,N_1819,N_1906);
nand U2470 (N_2470,N_1718,N_1645);
or U2471 (N_2471,N_1721,N_1857);
and U2472 (N_2472,N_1542,N_1652);
nand U2473 (N_2473,N_1870,N_1769);
or U2474 (N_2474,N_1552,N_1595);
nand U2475 (N_2475,N_1752,N_1912);
nand U2476 (N_2476,N_1653,N_1725);
nand U2477 (N_2477,N_1805,N_1663);
nand U2478 (N_2478,N_1931,N_1841);
nor U2479 (N_2479,N_1809,N_1733);
xor U2480 (N_2480,N_1517,N_1613);
or U2481 (N_2481,N_1861,N_1654);
nor U2482 (N_2482,N_1974,N_1697);
xor U2483 (N_2483,N_1986,N_1836);
nor U2484 (N_2484,N_1543,N_1551);
and U2485 (N_2485,N_1987,N_1646);
and U2486 (N_2486,N_1918,N_1826);
nor U2487 (N_2487,N_1621,N_1660);
or U2488 (N_2488,N_1500,N_1732);
or U2489 (N_2489,N_1751,N_1836);
or U2490 (N_2490,N_1692,N_1880);
or U2491 (N_2491,N_1733,N_1820);
xor U2492 (N_2492,N_1591,N_1527);
or U2493 (N_2493,N_1873,N_1541);
nand U2494 (N_2494,N_1716,N_1571);
nand U2495 (N_2495,N_1736,N_1581);
nand U2496 (N_2496,N_1573,N_1911);
and U2497 (N_2497,N_1985,N_1815);
nand U2498 (N_2498,N_1898,N_1749);
nand U2499 (N_2499,N_1899,N_1669);
and U2500 (N_2500,N_2417,N_2342);
and U2501 (N_2501,N_2421,N_2491);
or U2502 (N_2502,N_2096,N_2123);
xnor U2503 (N_2503,N_2095,N_2168);
xor U2504 (N_2504,N_2405,N_2035);
xor U2505 (N_2505,N_2238,N_2171);
or U2506 (N_2506,N_2235,N_2314);
xnor U2507 (N_2507,N_2222,N_2190);
or U2508 (N_2508,N_2220,N_2376);
or U2509 (N_2509,N_2056,N_2034);
or U2510 (N_2510,N_2079,N_2495);
or U2511 (N_2511,N_2151,N_2447);
xnor U2512 (N_2512,N_2204,N_2023);
and U2513 (N_2513,N_2442,N_2305);
xnor U2514 (N_2514,N_2464,N_2289);
xnor U2515 (N_2515,N_2488,N_2354);
nor U2516 (N_2516,N_2191,N_2101);
xor U2517 (N_2517,N_2025,N_2106);
and U2518 (N_2518,N_2043,N_2318);
nor U2519 (N_2519,N_2154,N_2327);
nor U2520 (N_2520,N_2391,N_2005);
or U2521 (N_2521,N_2343,N_2384);
xor U2522 (N_2522,N_2073,N_2399);
and U2523 (N_2523,N_2155,N_2382);
and U2524 (N_2524,N_2487,N_2370);
nand U2525 (N_2525,N_2250,N_2387);
nand U2526 (N_2526,N_2490,N_2273);
or U2527 (N_2527,N_2226,N_2252);
nor U2528 (N_2528,N_2437,N_2419);
nand U2529 (N_2529,N_2335,N_2129);
or U2530 (N_2530,N_2030,N_2348);
nor U2531 (N_2531,N_2429,N_2361);
nand U2532 (N_2532,N_2020,N_2069);
xnor U2533 (N_2533,N_2051,N_2213);
or U2534 (N_2534,N_2446,N_2149);
nor U2535 (N_2535,N_2140,N_2219);
xnor U2536 (N_2536,N_2356,N_2368);
or U2537 (N_2537,N_2074,N_2479);
or U2538 (N_2538,N_2138,N_2424);
xor U2539 (N_2539,N_2481,N_2156);
or U2540 (N_2540,N_2227,N_2320);
nand U2541 (N_2541,N_2071,N_2440);
nand U2542 (N_2542,N_2077,N_2102);
and U2543 (N_2543,N_2249,N_2054);
nor U2544 (N_2544,N_2459,N_2346);
and U2545 (N_2545,N_2359,N_2298);
nand U2546 (N_2546,N_2482,N_2211);
nor U2547 (N_2547,N_2414,N_2409);
and U2548 (N_2548,N_2205,N_2325);
or U2549 (N_2549,N_2053,N_2261);
nand U2550 (N_2550,N_2278,N_2036);
nand U2551 (N_2551,N_2108,N_2013);
xnor U2552 (N_2552,N_2124,N_2306);
nor U2553 (N_2553,N_2258,N_2009);
xnor U2554 (N_2554,N_2286,N_2264);
nand U2555 (N_2555,N_2497,N_2199);
xnor U2556 (N_2556,N_2097,N_2247);
nor U2557 (N_2557,N_2435,N_2060);
and U2558 (N_2558,N_2089,N_2179);
nand U2559 (N_2559,N_2494,N_2100);
or U2560 (N_2560,N_2115,N_2443);
nor U2561 (N_2561,N_2357,N_2350);
and U2562 (N_2562,N_2290,N_2111);
xor U2563 (N_2563,N_2090,N_2347);
and U2564 (N_2564,N_2087,N_2420);
nor U2565 (N_2565,N_2283,N_2113);
or U2566 (N_2566,N_2416,N_2112);
nor U2567 (N_2567,N_2334,N_2478);
xnor U2568 (N_2568,N_2277,N_2485);
and U2569 (N_2569,N_2031,N_2126);
and U2570 (N_2570,N_2322,N_2326);
or U2571 (N_2571,N_2048,N_2208);
nand U2572 (N_2572,N_2017,N_2174);
and U2573 (N_2573,N_2344,N_2144);
nand U2574 (N_2574,N_2225,N_2122);
xnor U2575 (N_2575,N_2324,N_2366);
nor U2576 (N_2576,N_2145,N_2426);
xor U2577 (N_2577,N_2055,N_2469);
nand U2578 (N_2578,N_2489,N_2180);
or U2579 (N_2579,N_2265,N_2068);
nor U2580 (N_2580,N_2128,N_2312);
or U2581 (N_2581,N_2170,N_2331);
or U2582 (N_2582,N_2449,N_2007);
or U2583 (N_2583,N_2285,N_2223);
nor U2584 (N_2584,N_2224,N_2460);
xor U2585 (N_2585,N_2098,N_2455);
xor U2586 (N_2586,N_2300,N_2181);
nand U2587 (N_2587,N_2232,N_2175);
nand U2588 (N_2588,N_2125,N_2270);
nor U2589 (N_2589,N_2423,N_2038);
xnor U2590 (N_2590,N_2483,N_2019);
nor U2591 (N_2591,N_2160,N_2292);
xor U2592 (N_2592,N_2130,N_2461);
xnor U2593 (N_2593,N_2301,N_2014);
nor U2594 (N_2594,N_2133,N_2498);
or U2595 (N_2595,N_2063,N_2099);
xor U2596 (N_2596,N_2291,N_2203);
nand U2597 (N_2597,N_2165,N_2003);
xor U2598 (N_2598,N_2159,N_2064);
and U2599 (N_2599,N_2315,N_2243);
and U2600 (N_2600,N_2187,N_2373);
xor U2601 (N_2601,N_2109,N_2476);
nor U2602 (N_2602,N_2212,N_2454);
nand U2603 (N_2603,N_2215,N_2287);
xnor U2604 (N_2604,N_2137,N_2418);
and U2605 (N_2605,N_2255,N_2297);
and U2606 (N_2606,N_2338,N_2193);
and U2607 (N_2607,N_2282,N_2186);
nor U2608 (N_2608,N_2016,N_2379);
nor U2609 (N_2609,N_2177,N_2148);
and U2610 (N_2610,N_2022,N_2351);
nand U2611 (N_2611,N_2248,N_2294);
xor U2612 (N_2612,N_2406,N_2234);
nor U2613 (N_2613,N_2217,N_2393);
xnor U2614 (N_2614,N_2448,N_2037);
and U2615 (N_2615,N_2044,N_2396);
nor U2616 (N_2616,N_2355,N_2345);
and U2617 (N_2617,N_2385,N_2093);
and U2618 (N_2618,N_2052,N_2018);
nor U2619 (N_2619,N_2092,N_2364);
and U2620 (N_2620,N_2404,N_2002);
xor U2621 (N_2621,N_2242,N_2229);
nor U2622 (N_2622,N_2336,N_2067);
nor U2623 (N_2623,N_2245,N_2163);
nand U2624 (N_2624,N_2083,N_2371);
or U2625 (N_2625,N_2272,N_2164);
nor U2626 (N_2626,N_2280,N_2457);
nor U2627 (N_2627,N_2015,N_2425);
or U2628 (N_2628,N_2178,N_2057);
nand U2629 (N_2629,N_2288,N_2275);
nor U2630 (N_2630,N_2276,N_2375);
and U2631 (N_2631,N_2441,N_2267);
nor U2632 (N_2632,N_2323,N_2062);
nand U2633 (N_2633,N_2358,N_2374);
nor U2634 (N_2634,N_2076,N_2380);
and U2635 (N_2635,N_2408,N_2228);
xor U2636 (N_2636,N_2263,N_2281);
xnor U2637 (N_2637,N_2474,N_2117);
or U2638 (N_2638,N_2244,N_2192);
nor U2639 (N_2639,N_2104,N_2430);
or U2640 (N_2640,N_2162,N_2422);
or U2641 (N_2641,N_2296,N_2352);
or U2642 (N_2642,N_2195,N_2050);
or U2643 (N_2643,N_2237,N_2450);
nor U2644 (N_2644,N_2365,N_2021);
and U2645 (N_2645,N_2086,N_2372);
nor U2646 (N_2646,N_2059,N_2012);
and U2647 (N_2647,N_2339,N_2011);
nand U2648 (N_2648,N_2027,N_2172);
and U2649 (N_2649,N_2214,N_2363);
xor U2650 (N_2650,N_2153,N_2400);
nor U2651 (N_2651,N_2369,N_2198);
nand U2652 (N_2652,N_2332,N_2231);
nand U2653 (N_2653,N_2236,N_2189);
xor U2654 (N_2654,N_2209,N_2394);
xor U2655 (N_2655,N_2493,N_2029);
xnor U2656 (N_2656,N_2284,N_2197);
xor U2657 (N_2657,N_2496,N_2088);
xor U2658 (N_2658,N_2360,N_2196);
xor U2659 (N_2659,N_2202,N_2028);
nor U2660 (N_2660,N_2321,N_2184);
xor U2661 (N_2661,N_2456,N_2047);
or U2662 (N_2662,N_2049,N_2246);
nor U2663 (N_2663,N_2407,N_2377);
xnor U2664 (N_2664,N_2006,N_2157);
or U2665 (N_2665,N_2110,N_2010);
nand U2666 (N_2666,N_2472,N_2026);
and U2667 (N_2667,N_2042,N_2000);
nor U2668 (N_2668,N_2254,N_2433);
nand U2669 (N_2669,N_2158,N_2239);
xor U2670 (N_2670,N_2432,N_2438);
nor U2671 (N_2671,N_2230,N_2072);
nand U2672 (N_2672,N_2458,N_2081);
and U2673 (N_2673,N_2210,N_2462);
xor U2674 (N_2674,N_2107,N_2136);
nor U2675 (N_2675,N_2453,N_2094);
and U2676 (N_2676,N_2152,N_2166);
nand U2677 (N_2677,N_2127,N_2415);
nor U2678 (N_2678,N_2032,N_2135);
xor U2679 (N_2679,N_2182,N_2311);
nand U2680 (N_2680,N_2295,N_2431);
or U2681 (N_2681,N_2139,N_2467);
or U2682 (N_2682,N_2259,N_2183);
nand U2683 (N_2683,N_2266,N_2388);
nand U2684 (N_2684,N_2241,N_2045);
xnor U2685 (N_2685,N_2221,N_2468);
xnor U2686 (N_2686,N_2046,N_2389);
and U2687 (N_2687,N_2120,N_2480);
nor U2688 (N_2688,N_2121,N_2040);
nor U2689 (N_2689,N_2176,N_2084);
nand U2690 (N_2690,N_2328,N_2341);
and U2691 (N_2691,N_2173,N_2367);
xnor U2692 (N_2692,N_2240,N_2085);
xor U2693 (N_2693,N_2378,N_2251);
nand U2694 (N_2694,N_2233,N_2317);
nor U2695 (N_2695,N_2473,N_2041);
nor U2696 (N_2696,N_2309,N_2340);
nor U2697 (N_2697,N_2492,N_2066);
nand U2698 (N_2698,N_2024,N_2119);
nor U2699 (N_2699,N_2116,N_2253);
nor U2700 (N_2700,N_2411,N_2161);
xor U2701 (N_2701,N_2398,N_2033);
and U2702 (N_2702,N_2392,N_2465);
nor U2703 (N_2703,N_2444,N_2381);
nor U2704 (N_2704,N_2188,N_2452);
and U2705 (N_2705,N_2004,N_2439);
nor U2706 (N_2706,N_2362,N_2065);
or U2707 (N_2707,N_2397,N_2082);
nor U2708 (N_2708,N_2477,N_2436);
xnor U2709 (N_2709,N_2262,N_2413);
nand U2710 (N_2710,N_2299,N_2080);
xor U2711 (N_2711,N_2268,N_2279);
or U2712 (N_2712,N_2169,N_2134);
or U2713 (N_2713,N_2070,N_2383);
and U2714 (N_2714,N_2206,N_2390);
nand U2715 (N_2715,N_2218,N_2260);
nor U2716 (N_2716,N_2185,N_2131);
nor U2717 (N_2717,N_2142,N_2132);
or U2718 (N_2718,N_2147,N_2316);
xor U2719 (N_2719,N_2271,N_2091);
nand U2720 (N_2720,N_2463,N_2058);
xnor U2721 (N_2721,N_2201,N_2403);
nor U2722 (N_2722,N_2207,N_2269);
nand U2723 (N_2723,N_2216,N_2307);
and U2724 (N_2724,N_2410,N_2471);
or U2725 (N_2725,N_2333,N_2308);
nand U2726 (N_2726,N_2313,N_2499);
nor U2727 (N_2727,N_2475,N_2075);
nor U2728 (N_2728,N_2310,N_2401);
and U2729 (N_2729,N_2402,N_2486);
nand U2730 (N_2730,N_2143,N_2293);
and U2731 (N_2731,N_2078,N_2146);
xor U2732 (N_2732,N_2330,N_2114);
nor U2733 (N_2733,N_2319,N_2008);
nand U2734 (N_2734,N_2039,N_2412);
nand U2735 (N_2735,N_2337,N_2103);
or U2736 (N_2736,N_2118,N_2001);
or U2737 (N_2737,N_2303,N_2274);
nor U2738 (N_2738,N_2445,N_2466);
or U2739 (N_2739,N_2451,N_2105);
nor U2740 (N_2740,N_2141,N_2302);
xor U2741 (N_2741,N_2257,N_2353);
nor U2742 (N_2742,N_2434,N_2484);
or U2743 (N_2743,N_2167,N_2349);
and U2744 (N_2744,N_2194,N_2386);
nand U2745 (N_2745,N_2150,N_2061);
nor U2746 (N_2746,N_2470,N_2200);
nor U2747 (N_2747,N_2395,N_2427);
xnor U2748 (N_2748,N_2256,N_2428);
or U2749 (N_2749,N_2329,N_2304);
xnor U2750 (N_2750,N_2316,N_2034);
nand U2751 (N_2751,N_2134,N_2482);
nor U2752 (N_2752,N_2331,N_2249);
nor U2753 (N_2753,N_2156,N_2106);
or U2754 (N_2754,N_2468,N_2182);
xor U2755 (N_2755,N_2217,N_2428);
and U2756 (N_2756,N_2017,N_2283);
or U2757 (N_2757,N_2427,N_2031);
or U2758 (N_2758,N_2387,N_2062);
nor U2759 (N_2759,N_2168,N_2016);
nor U2760 (N_2760,N_2296,N_2493);
nand U2761 (N_2761,N_2052,N_2377);
and U2762 (N_2762,N_2051,N_2304);
and U2763 (N_2763,N_2027,N_2277);
nor U2764 (N_2764,N_2442,N_2441);
and U2765 (N_2765,N_2199,N_2182);
nor U2766 (N_2766,N_2497,N_2024);
xor U2767 (N_2767,N_2425,N_2054);
nor U2768 (N_2768,N_2351,N_2167);
xor U2769 (N_2769,N_2207,N_2358);
and U2770 (N_2770,N_2092,N_2335);
and U2771 (N_2771,N_2451,N_2373);
xor U2772 (N_2772,N_2341,N_2093);
nor U2773 (N_2773,N_2371,N_2485);
and U2774 (N_2774,N_2169,N_2125);
or U2775 (N_2775,N_2092,N_2260);
nor U2776 (N_2776,N_2064,N_2495);
or U2777 (N_2777,N_2447,N_2155);
or U2778 (N_2778,N_2277,N_2311);
xor U2779 (N_2779,N_2464,N_2157);
xnor U2780 (N_2780,N_2044,N_2212);
or U2781 (N_2781,N_2402,N_2237);
or U2782 (N_2782,N_2476,N_2074);
nand U2783 (N_2783,N_2203,N_2127);
xor U2784 (N_2784,N_2062,N_2429);
nand U2785 (N_2785,N_2322,N_2108);
and U2786 (N_2786,N_2374,N_2382);
nor U2787 (N_2787,N_2026,N_2475);
nand U2788 (N_2788,N_2328,N_2170);
nand U2789 (N_2789,N_2359,N_2334);
nand U2790 (N_2790,N_2227,N_2222);
nor U2791 (N_2791,N_2244,N_2485);
or U2792 (N_2792,N_2455,N_2075);
and U2793 (N_2793,N_2011,N_2269);
or U2794 (N_2794,N_2123,N_2158);
xnor U2795 (N_2795,N_2409,N_2270);
and U2796 (N_2796,N_2139,N_2173);
xor U2797 (N_2797,N_2237,N_2193);
nor U2798 (N_2798,N_2476,N_2117);
nand U2799 (N_2799,N_2230,N_2088);
nand U2800 (N_2800,N_2294,N_2478);
nand U2801 (N_2801,N_2256,N_2473);
xor U2802 (N_2802,N_2453,N_2079);
and U2803 (N_2803,N_2377,N_2328);
nand U2804 (N_2804,N_2085,N_2479);
and U2805 (N_2805,N_2019,N_2243);
and U2806 (N_2806,N_2396,N_2353);
xor U2807 (N_2807,N_2326,N_2157);
and U2808 (N_2808,N_2265,N_2282);
nand U2809 (N_2809,N_2194,N_2018);
and U2810 (N_2810,N_2257,N_2024);
nand U2811 (N_2811,N_2422,N_2420);
xor U2812 (N_2812,N_2029,N_2147);
nor U2813 (N_2813,N_2040,N_2186);
nand U2814 (N_2814,N_2369,N_2235);
and U2815 (N_2815,N_2469,N_2243);
nand U2816 (N_2816,N_2473,N_2498);
or U2817 (N_2817,N_2364,N_2416);
or U2818 (N_2818,N_2299,N_2070);
and U2819 (N_2819,N_2285,N_2458);
nor U2820 (N_2820,N_2146,N_2364);
or U2821 (N_2821,N_2332,N_2268);
or U2822 (N_2822,N_2128,N_2227);
and U2823 (N_2823,N_2410,N_2291);
nand U2824 (N_2824,N_2407,N_2383);
and U2825 (N_2825,N_2025,N_2387);
xor U2826 (N_2826,N_2118,N_2013);
nand U2827 (N_2827,N_2086,N_2476);
nor U2828 (N_2828,N_2020,N_2047);
nand U2829 (N_2829,N_2118,N_2207);
or U2830 (N_2830,N_2455,N_2236);
or U2831 (N_2831,N_2110,N_2263);
or U2832 (N_2832,N_2365,N_2071);
xor U2833 (N_2833,N_2458,N_2300);
and U2834 (N_2834,N_2414,N_2125);
nand U2835 (N_2835,N_2419,N_2136);
or U2836 (N_2836,N_2393,N_2162);
xor U2837 (N_2837,N_2085,N_2097);
or U2838 (N_2838,N_2134,N_2455);
xor U2839 (N_2839,N_2065,N_2250);
or U2840 (N_2840,N_2120,N_2497);
xor U2841 (N_2841,N_2392,N_2332);
and U2842 (N_2842,N_2296,N_2478);
xnor U2843 (N_2843,N_2072,N_2290);
or U2844 (N_2844,N_2248,N_2257);
or U2845 (N_2845,N_2003,N_2028);
nand U2846 (N_2846,N_2223,N_2043);
xor U2847 (N_2847,N_2252,N_2135);
or U2848 (N_2848,N_2479,N_2317);
xnor U2849 (N_2849,N_2495,N_2487);
nand U2850 (N_2850,N_2264,N_2138);
and U2851 (N_2851,N_2139,N_2236);
or U2852 (N_2852,N_2021,N_2374);
nor U2853 (N_2853,N_2309,N_2179);
or U2854 (N_2854,N_2151,N_2261);
and U2855 (N_2855,N_2213,N_2306);
and U2856 (N_2856,N_2080,N_2470);
and U2857 (N_2857,N_2056,N_2084);
nand U2858 (N_2858,N_2149,N_2195);
nand U2859 (N_2859,N_2385,N_2282);
and U2860 (N_2860,N_2360,N_2263);
and U2861 (N_2861,N_2198,N_2227);
nand U2862 (N_2862,N_2114,N_2017);
or U2863 (N_2863,N_2446,N_2463);
nor U2864 (N_2864,N_2087,N_2432);
nand U2865 (N_2865,N_2046,N_2205);
nand U2866 (N_2866,N_2080,N_2138);
nor U2867 (N_2867,N_2017,N_2187);
nand U2868 (N_2868,N_2319,N_2382);
and U2869 (N_2869,N_2403,N_2359);
nand U2870 (N_2870,N_2442,N_2347);
or U2871 (N_2871,N_2124,N_2434);
nand U2872 (N_2872,N_2217,N_2354);
or U2873 (N_2873,N_2179,N_2169);
or U2874 (N_2874,N_2407,N_2072);
nand U2875 (N_2875,N_2230,N_2251);
nor U2876 (N_2876,N_2311,N_2323);
and U2877 (N_2877,N_2134,N_2241);
or U2878 (N_2878,N_2466,N_2224);
and U2879 (N_2879,N_2125,N_2309);
xnor U2880 (N_2880,N_2163,N_2442);
or U2881 (N_2881,N_2122,N_2352);
xor U2882 (N_2882,N_2296,N_2303);
xnor U2883 (N_2883,N_2479,N_2415);
nand U2884 (N_2884,N_2468,N_2358);
nand U2885 (N_2885,N_2089,N_2464);
nand U2886 (N_2886,N_2049,N_2487);
nor U2887 (N_2887,N_2059,N_2050);
nor U2888 (N_2888,N_2432,N_2117);
nor U2889 (N_2889,N_2238,N_2484);
and U2890 (N_2890,N_2231,N_2322);
or U2891 (N_2891,N_2386,N_2334);
and U2892 (N_2892,N_2147,N_2046);
nor U2893 (N_2893,N_2427,N_2047);
and U2894 (N_2894,N_2242,N_2497);
and U2895 (N_2895,N_2439,N_2484);
xor U2896 (N_2896,N_2260,N_2117);
or U2897 (N_2897,N_2264,N_2257);
and U2898 (N_2898,N_2091,N_2422);
or U2899 (N_2899,N_2473,N_2340);
nor U2900 (N_2900,N_2451,N_2447);
nor U2901 (N_2901,N_2473,N_2214);
nor U2902 (N_2902,N_2359,N_2251);
xnor U2903 (N_2903,N_2129,N_2287);
and U2904 (N_2904,N_2298,N_2050);
xnor U2905 (N_2905,N_2125,N_2344);
or U2906 (N_2906,N_2077,N_2011);
and U2907 (N_2907,N_2292,N_2164);
nand U2908 (N_2908,N_2413,N_2049);
xor U2909 (N_2909,N_2122,N_2384);
or U2910 (N_2910,N_2311,N_2010);
xnor U2911 (N_2911,N_2459,N_2128);
xor U2912 (N_2912,N_2410,N_2285);
and U2913 (N_2913,N_2254,N_2382);
xor U2914 (N_2914,N_2155,N_2282);
nor U2915 (N_2915,N_2249,N_2270);
and U2916 (N_2916,N_2032,N_2238);
and U2917 (N_2917,N_2197,N_2193);
nand U2918 (N_2918,N_2312,N_2390);
nor U2919 (N_2919,N_2057,N_2110);
nor U2920 (N_2920,N_2006,N_2016);
xor U2921 (N_2921,N_2381,N_2099);
nand U2922 (N_2922,N_2411,N_2032);
xor U2923 (N_2923,N_2207,N_2017);
or U2924 (N_2924,N_2243,N_2098);
nand U2925 (N_2925,N_2331,N_2089);
or U2926 (N_2926,N_2491,N_2070);
xnor U2927 (N_2927,N_2453,N_2008);
and U2928 (N_2928,N_2339,N_2069);
and U2929 (N_2929,N_2110,N_2412);
nor U2930 (N_2930,N_2264,N_2353);
and U2931 (N_2931,N_2163,N_2132);
or U2932 (N_2932,N_2053,N_2461);
nand U2933 (N_2933,N_2353,N_2208);
xor U2934 (N_2934,N_2275,N_2495);
and U2935 (N_2935,N_2292,N_2305);
xnor U2936 (N_2936,N_2006,N_2375);
or U2937 (N_2937,N_2441,N_2163);
nor U2938 (N_2938,N_2177,N_2350);
and U2939 (N_2939,N_2058,N_2198);
nor U2940 (N_2940,N_2001,N_2445);
and U2941 (N_2941,N_2348,N_2051);
nand U2942 (N_2942,N_2051,N_2303);
and U2943 (N_2943,N_2360,N_2232);
nand U2944 (N_2944,N_2392,N_2173);
and U2945 (N_2945,N_2047,N_2129);
nor U2946 (N_2946,N_2252,N_2395);
nor U2947 (N_2947,N_2174,N_2025);
xnor U2948 (N_2948,N_2488,N_2459);
nand U2949 (N_2949,N_2064,N_2023);
or U2950 (N_2950,N_2240,N_2453);
or U2951 (N_2951,N_2275,N_2191);
nand U2952 (N_2952,N_2281,N_2429);
and U2953 (N_2953,N_2245,N_2307);
nand U2954 (N_2954,N_2385,N_2163);
nand U2955 (N_2955,N_2269,N_2069);
and U2956 (N_2956,N_2076,N_2090);
or U2957 (N_2957,N_2337,N_2270);
nor U2958 (N_2958,N_2134,N_2323);
or U2959 (N_2959,N_2102,N_2353);
or U2960 (N_2960,N_2050,N_2179);
nand U2961 (N_2961,N_2365,N_2488);
nor U2962 (N_2962,N_2405,N_2487);
and U2963 (N_2963,N_2200,N_2166);
and U2964 (N_2964,N_2251,N_2300);
xor U2965 (N_2965,N_2268,N_2374);
or U2966 (N_2966,N_2061,N_2132);
xor U2967 (N_2967,N_2048,N_2356);
nor U2968 (N_2968,N_2022,N_2300);
nand U2969 (N_2969,N_2445,N_2009);
and U2970 (N_2970,N_2441,N_2224);
nor U2971 (N_2971,N_2295,N_2413);
or U2972 (N_2972,N_2181,N_2168);
or U2973 (N_2973,N_2447,N_2053);
or U2974 (N_2974,N_2494,N_2092);
nor U2975 (N_2975,N_2474,N_2373);
or U2976 (N_2976,N_2249,N_2174);
or U2977 (N_2977,N_2326,N_2084);
nor U2978 (N_2978,N_2211,N_2147);
nand U2979 (N_2979,N_2304,N_2493);
nand U2980 (N_2980,N_2013,N_2094);
nor U2981 (N_2981,N_2087,N_2479);
or U2982 (N_2982,N_2296,N_2330);
nand U2983 (N_2983,N_2188,N_2484);
nor U2984 (N_2984,N_2115,N_2447);
nor U2985 (N_2985,N_2358,N_2472);
or U2986 (N_2986,N_2073,N_2495);
nand U2987 (N_2987,N_2459,N_2314);
xnor U2988 (N_2988,N_2145,N_2054);
and U2989 (N_2989,N_2300,N_2271);
and U2990 (N_2990,N_2230,N_2415);
and U2991 (N_2991,N_2217,N_2187);
xor U2992 (N_2992,N_2054,N_2331);
xor U2993 (N_2993,N_2414,N_2420);
or U2994 (N_2994,N_2022,N_2100);
xnor U2995 (N_2995,N_2242,N_2406);
and U2996 (N_2996,N_2495,N_2233);
and U2997 (N_2997,N_2375,N_2107);
nor U2998 (N_2998,N_2038,N_2018);
nand U2999 (N_2999,N_2263,N_2354);
xnor U3000 (N_3000,N_2534,N_2897);
or U3001 (N_3001,N_2876,N_2825);
nand U3002 (N_3002,N_2948,N_2646);
nand U3003 (N_3003,N_2577,N_2996);
and U3004 (N_3004,N_2706,N_2958);
nand U3005 (N_3005,N_2853,N_2529);
nand U3006 (N_3006,N_2874,N_2630);
xor U3007 (N_3007,N_2500,N_2538);
or U3008 (N_3008,N_2769,N_2603);
nor U3009 (N_3009,N_2916,N_2802);
nand U3010 (N_3010,N_2522,N_2644);
and U3011 (N_3011,N_2528,N_2701);
nor U3012 (N_3012,N_2821,N_2896);
nor U3013 (N_3013,N_2679,N_2531);
nand U3014 (N_3014,N_2953,N_2660);
and U3015 (N_3015,N_2847,N_2928);
nand U3016 (N_3016,N_2940,N_2804);
nor U3017 (N_3017,N_2653,N_2602);
or U3018 (N_3018,N_2540,N_2517);
and U3019 (N_3019,N_2915,N_2803);
nor U3020 (N_3020,N_2886,N_2748);
nand U3021 (N_3021,N_2667,N_2725);
nand U3022 (N_3022,N_2558,N_2910);
nand U3023 (N_3023,N_2979,N_2614);
nand U3024 (N_3024,N_2519,N_2892);
xnor U3025 (N_3025,N_2641,N_2645);
nor U3026 (N_3026,N_2521,N_2741);
xor U3027 (N_3027,N_2530,N_2723);
nand U3028 (N_3028,N_2759,N_2815);
xor U3029 (N_3029,N_2911,N_2676);
or U3030 (N_3030,N_2999,N_2840);
nand U3031 (N_3031,N_2733,N_2505);
nor U3032 (N_3032,N_2728,N_2978);
xnor U3033 (N_3033,N_2939,N_2836);
nand U3034 (N_3034,N_2852,N_2581);
or U3035 (N_3035,N_2511,N_2616);
nor U3036 (N_3036,N_2729,N_2560);
and U3037 (N_3037,N_2787,N_2790);
xor U3038 (N_3038,N_2634,N_2643);
or U3039 (N_3039,N_2514,N_2833);
and U3040 (N_3040,N_2651,N_2975);
nor U3041 (N_3041,N_2649,N_2848);
nor U3042 (N_3042,N_2627,N_2745);
or U3043 (N_3043,N_2889,N_2633);
and U3044 (N_3044,N_2995,N_2887);
xnor U3045 (N_3045,N_2515,N_2970);
xor U3046 (N_3046,N_2687,N_2718);
nand U3047 (N_3047,N_2596,N_2609);
nor U3048 (N_3048,N_2772,N_2883);
and U3049 (N_3049,N_2544,N_2561);
and U3050 (N_3050,N_2582,N_2749);
or U3051 (N_3051,N_2942,N_2754);
and U3052 (N_3052,N_2684,N_2888);
and U3053 (N_3053,N_2795,N_2980);
or U3054 (N_3054,N_2762,N_2782);
nand U3055 (N_3055,N_2924,N_2512);
nor U3056 (N_3056,N_2779,N_2583);
or U3057 (N_3057,N_2721,N_2696);
nor U3058 (N_3058,N_2981,N_2568);
nand U3059 (N_3059,N_2793,N_2501);
nand U3060 (N_3060,N_2824,N_2920);
xor U3061 (N_3061,N_2699,N_2952);
or U3062 (N_3062,N_2593,N_2554);
or U3063 (N_3063,N_2600,N_2605);
nor U3064 (N_3064,N_2599,N_2771);
xor U3065 (N_3065,N_2993,N_2907);
nand U3066 (N_3066,N_2758,N_2677);
and U3067 (N_3067,N_2909,N_2800);
or U3068 (N_3068,N_2869,N_2868);
nand U3069 (N_3069,N_2757,N_2575);
nand U3070 (N_3070,N_2674,N_2751);
or U3071 (N_3071,N_2797,N_2722);
nor U3072 (N_3072,N_2893,N_2965);
and U3073 (N_3073,N_2933,N_2595);
nand U3074 (N_3074,N_2835,N_2918);
nand U3075 (N_3075,N_2564,N_2923);
or U3076 (N_3076,N_2601,N_2855);
nor U3077 (N_3077,N_2552,N_2691);
xor U3078 (N_3078,N_2610,N_2672);
or U3079 (N_3079,N_2623,N_2624);
nor U3080 (N_3080,N_2932,N_2811);
nand U3081 (N_3081,N_2826,N_2525);
nor U3082 (N_3082,N_2827,N_2982);
nand U3083 (N_3083,N_2956,N_2670);
nand U3084 (N_3084,N_2508,N_2556);
xnor U3085 (N_3085,N_2579,N_2866);
nor U3086 (N_3086,N_2550,N_2668);
nand U3087 (N_3087,N_2807,N_2744);
or U3088 (N_3088,N_2792,N_2776);
nor U3089 (N_3089,N_2551,N_2647);
and U3090 (N_3090,N_2941,N_2740);
xnor U3091 (N_3091,N_2708,N_2565);
or U3092 (N_3092,N_2929,N_2693);
nor U3093 (N_3093,N_2781,N_2526);
xor U3094 (N_3094,N_2695,N_2694);
nand U3095 (N_3095,N_2997,N_2770);
or U3096 (N_3096,N_2764,N_2871);
nand U3097 (N_3097,N_2832,N_2656);
nand U3098 (N_3098,N_2654,N_2700);
xnor U3099 (N_3099,N_2523,N_2843);
nand U3100 (N_3100,N_2655,N_2613);
or U3101 (N_3101,N_2845,N_2681);
nor U3102 (N_3102,N_2882,N_2806);
or U3103 (N_3103,N_2716,N_2503);
and U3104 (N_3104,N_2799,N_2927);
xor U3105 (N_3105,N_2894,N_2831);
nand U3106 (N_3106,N_2620,N_2714);
and U3107 (N_3107,N_2713,N_2900);
xnor U3108 (N_3108,N_2664,N_2973);
xor U3109 (N_3109,N_2865,N_2686);
nor U3110 (N_3110,N_2704,N_2798);
or U3111 (N_3111,N_2612,N_2536);
xor U3112 (N_3112,N_2917,N_2912);
and U3113 (N_3113,N_2930,N_2870);
and U3114 (N_3114,N_2625,N_2709);
xor U3115 (N_3115,N_2904,N_2559);
and U3116 (N_3116,N_2765,N_2658);
nor U3117 (N_3117,N_2990,N_2961);
xnor U3118 (N_3118,N_2678,N_2618);
xnor U3119 (N_3119,N_2985,N_2563);
or U3120 (N_3120,N_2592,N_2830);
and U3121 (N_3121,N_2922,N_2527);
or U3122 (N_3122,N_2860,N_2947);
and U3123 (N_3123,N_2663,N_2669);
xor U3124 (N_3124,N_2862,N_2705);
or U3125 (N_3125,N_2502,N_2775);
or U3126 (N_3126,N_2743,N_2629);
or U3127 (N_3127,N_2959,N_2969);
xnor U3128 (N_3128,N_2532,N_2931);
nand U3129 (N_3129,N_2584,N_2842);
nor U3130 (N_3130,N_2650,N_2546);
nand U3131 (N_3131,N_2750,N_2507);
nor U3132 (N_3132,N_2884,N_2591);
and U3133 (N_3133,N_2727,N_2573);
or U3134 (N_3134,N_2680,N_2937);
nand U3135 (N_3135,N_2574,N_2987);
and U3136 (N_3136,N_2533,N_2549);
nor U3137 (N_3137,N_2587,N_2657);
or U3138 (N_3138,N_2566,N_2976);
nand U3139 (N_3139,N_2877,N_2607);
and U3140 (N_3140,N_2838,N_2784);
nand U3141 (N_3141,N_2611,N_2992);
or U3142 (N_3142,N_2880,N_2968);
and U3143 (N_3143,N_2822,N_2829);
nand U3144 (N_3144,N_2903,N_2783);
xnor U3145 (N_3145,N_2908,N_2518);
nor U3146 (N_3146,N_2662,N_2777);
or U3147 (N_3147,N_2617,N_2682);
nor U3148 (N_3148,N_2785,N_2542);
and U3149 (N_3149,N_2801,N_2814);
nor U3150 (N_3150,N_2895,N_2755);
xor U3151 (N_3151,N_2632,N_2766);
nand U3152 (N_3152,N_2683,N_2925);
nand U3153 (N_3153,N_2638,N_2712);
nor U3154 (N_3154,N_2977,N_2513);
xor U3155 (N_3155,N_2988,N_2547);
or U3156 (N_3156,N_2626,N_2752);
xor U3157 (N_3157,N_2813,N_2690);
xor U3158 (N_3158,N_2944,N_2901);
and U3159 (N_3159,N_2703,N_2742);
nand U3160 (N_3160,N_2934,N_2585);
and U3161 (N_3161,N_2535,N_2872);
xnor U3162 (N_3162,N_2966,N_2688);
nor U3163 (N_3163,N_2994,N_2805);
xnor U3164 (N_3164,N_2606,N_2841);
xor U3165 (N_3165,N_2780,N_2639);
or U3166 (N_3166,N_2562,N_2571);
nor U3167 (N_3167,N_2586,N_2820);
and U3168 (N_3168,N_2962,N_2516);
or U3169 (N_3169,N_2671,N_2955);
or U3170 (N_3170,N_2590,N_2545);
and U3171 (N_3171,N_2850,N_2857);
and U3172 (N_3172,N_2636,N_2567);
nor U3173 (N_3173,N_2761,N_2796);
nand U3174 (N_3174,N_2726,N_2951);
xor U3175 (N_3175,N_2875,N_2823);
xor U3176 (N_3176,N_2789,N_2763);
xor U3177 (N_3177,N_2898,N_2812);
nor U3178 (N_3178,N_2753,N_2637);
nand U3179 (N_3179,N_2986,N_2778);
xor U3180 (N_3180,N_2572,N_2879);
nor U3181 (N_3181,N_2891,N_2756);
xor U3182 (N_3182,N_2859,N_2767);
or U3183 (N_3183,N_2867,N_2998);
or U3184 (N_3184,N_2984,N_2808);
xnor U3185 (N_3185,N_2537,N_2739);
nor U3186 (N_3186,N_2899,N_2863);
nor U3187 (N_3187,N_2828,N_2957);
nand U3188 (N_3188,N_2724,N_2816);
nand U3189 (N_3189,N_2746,N_2510);
xor U3190 (N_3190,N_2991,N_2858);
or U3191 (N_3191,N_2819,N_2738);
xor U3192 (N_3192,N_2856,N_2715);
xnor U3193 (N_3193,N_2989,N_2817);
nand U3194 (N_3194,N_2737,N_2692);
and U3195 (N_3195,N_2570,N_2818);
nor U3196 (N_3196,N_2971,N_2509);
nand U3197 (N_3197,N_2661,N_2949);
and U3198 (N_3198,N_2938,N_2707);
nor U3199 (N_3199,N_2926,N_2885);
nand U3200 (N_3200,N_2839,N_2648);
and U3201 (N_3201,N_2619,N_2553);
or U3202 (N_3202,N_2640,N_2675);
nor U3203 (N_3203,N_2878,N_2734);
or U3204 (N_3204,N_2697,N_2946);
and U3205 (N_3205,N_2861,N_2578);
nand U3206 (N_3206,N_2631,N_2557);
and U3207 (N_3207,N_2588,N_2936);
and U3208 (N_3208,N_2844,N_2642);
xnor U3209 (N_3209,N_2881,N_2773);
nand U3210 (N_3210,N_2873,N_2506);
and U3211 (N_3211,N_2849,N_2921);
nand U3212 (N_3212,N_2665,N_2543);
nand U3213 (N_3213,N_2589,N_2604);
and U3214 (N_3214,N_2730,N_2524);
xnor U3215 (N_3215,N_2788,N_2837);
nand U3216 (N_3216,N_2702,N_2615);
xor U3217 (N_3217,N_2666,N_2659);
nand U3218 (N_3218,N_2628,N_2580);
xnor U3219 (N_3219,N_2954,N_2791);
xor U3220 (N_3220,N_2735,N_2731);
and U3221 (N_3221,N_2539,N_2945);
or U3222 (N_3222,N_2504,N_2711);
and U3223 (N_3223,N_2594,N_2736);
nor U3224 (N_3224,N_2720,N_2794);
xor U3225 (N_3225,N_2786,N_2964);
xor U3226 (N_3226,N_2732,N_2555);
and U3227 (N_3227,N_2710,N_2621);
nand U3228 (N_3228,N_2698,N_2902);
and U3229 (N_3229,N_2905,N_2569);
nor U3230 (N_3230,N_2967,N_2809);
nand U3231 (N_3231,N_2673,N_2768);
or U3232 (N_3232,N_2689,N_2685);
nand U3233 (N_3233,N_2774,N_2598);
nand U3234 (N_3234,N_2919,N_2960);
nor U3235 (N_3235,N_2972,N_2846);
or U3236 (N_3236,N_2597,N_2548);
xor U3237 (N_3237,N_2913,N_2943);
nor U3238 (N_3238,N_2864,N_2851);
nor U3239 (N_3239,N_2717,N_2622);
xor U3240 (N_3240,N_2935,N_2760);
xnor U3241 (N_3241,N_2974,N_2520);
and U3242 (N_3242,N_2906,N_2652);
nand U3243 (N_3243,N_2635,N_2719);
xor U3244 (N_3244,N_2810,N_2963);
nand U3245 (N_3245,N_2541,N_2890);
xnor U3246 (N_3246,N_2914,N_2608);
xnor U3247 (N_3247,N_2854,N_2950);
or U3248 (N_3248,N_2576,N_2983);
nand U3249 (N_3249,N_2834,N_2747);
or U3250 (N_3250,N_2688,N_2747);
or U3251 (N_3251,N_2622,N_2658);
or U3252 (N_3252,N_2656,N_2546);
and U3253 (N_3253,N_2869,N_2827);
nand U3254 (N_3254,N_2584,N_2846);
nor U3255 (N_3255,N_2558,N_2609);
or U3256 (N_3256,N_2736,N_2922);
nand U3257 (N_3257,N_2898,N_2879);
nor U3258 (N_3258,N_2602,N_2622);
nand U3259 (N_3259,N_2696,N_2983);
nor U3260 (N_3260,N_2724,N_2611);
or U3261 (N_3261,N_2984,N_2985);
nand U3262 (N_3262,N_2915,N_2680);
xnor U3263 (N_3263,N_2588,N_2916);
nand U3264 (N_3264,N_2702,N_2551);
or U3265 (N_3265,N_2804,N_2809);
nor U3266 (N_3266,N_2921,N_2905);
nand U3267 (N_3267,N_2506,N_2685);
and U3268 (N_3268,N_2643,N_2536);
or U3269 (N_3269,N_2706,N_2735);
or U3270 (N_3270,N_2918,N_2655);
xor U3271 (N_3271,N_2712,N_2722);
xor U3272 (N_3272,N_2813,N_2507);
xnor U3273 (N_3273,N_2531,N_2764);
and U3274 (N_3274,N_2571,N_2951);
and U3275 (N_3275,N_2832,N_2591);
or U3276 (N_3276,N_2968,N_2614);
nor U3277 (N_3277,N_2696,N_2688);
nand U3278 (N_3278,N_2605,N_2764);
or U3279 (N_3279,N_2630,N_2895);
and U3280 (N_3280,N_2910,N_2567);
and U3281 (N_3281,N_2752,N_2714);
or U3282 (N_3282,N_2506,N_2823);
or U3283 (N_3283,N_2540,N_2852);
nand U3284 (N_3284,N_2647,N_2985);
nor U3285 (N_3285,N_2703,N_2558);
and U3286 (N_3286,N_2720,N_2609);
xnor U3287 (N_3287,N_2775,N_2787);
xor U3288 (N_3288,N_2672,N_2848);
nand U3289 (N_3289,N_2516,N_2894);
and U3290 (N_3290,N_2859,N_2679);
nor U3291 (N_3291,N_2991,N_2904);
xor U3292 (N_3292,N_2887,N_2649);
xor U3293 (N_3293,N_2958,N_2565);
and U3294 (N_3294,N_2993,N_2848);
and U3295 (N_3295,N_2665,N_2690);
and U3296 (N_3296,N_2870,N_2989);
and U3297 (N_3297,N_2738,N_2589);
or U3298 (N_3298,N_2739,N_2834);
and U3299 (N_3299,N_2941,N_2584);
and U3300 (N_3300,N_2770,N_2658);
or U3301 (N_3301,N_2509,N_2591);
and U3302 (N_3302,N_2886,N_2879);
xor U3303 (N_3303,N_2768,N_2956);
nand U3304 (N_3304,N_2504,N_2714);
nand U3305 (N_3305,N_2819,N_2645);
nor U3306 (N_3306,N_2929,N_2806);
nand U3307 (N_3307,N_2981,N_2824);
nor U3308 (N_3308,N_2938,N_2506);
xor U3309 (N_3309,N_2811,N_2521);
and U3310 (N_3310,N_2540,N_2752);
xnor U3311 (N_3311,N_2737,N_2983);
nor U3312 (N_3312,N_2958,N_2518);
nand U3313 (N_3313,N_2588,N_2626);
and U3314 (N_3314,N_2617,N_2643);
or U3315 (N_3315,N_2657,N_2565);
or U3316 (N_3316,N_2635,N_2836);
nor U3317 (N_3317,N_2970,N_2758);
and U3318 (N_3318,N_2709,N_2547);
and U3319 (N_3319,N_2622,N_2762);
or U3320 (N_3320,N_2876,N_2595);
and U3321 (N_3321,N_2588,N_2947);
and U3322 (N_3322,N_2572,N_2917);
or U3323 (N_3323,N_2765,N_2913);
nor U3324 (N_3324,N_2741,N_2591);
nor U3325 (N_3325,N_2984,N_2736);
and U3326 (N_3326,N_2670,N_2707);
xor U3327 (N_3327,N_2819,N_2591);
xor U3328 (N_3328,N_2515,N_2928);
xor U3329 (N_3329,N_2602,N_2978);
and U3330 (N_3330,N_2563,N_2507);
or U3331 (N_3331,N_2861,N_2855);
nand U3332 (N_3332,N_2793,N_2886);
or U3333 (N_3333,N_2557,N_2915);
nand U3334 (N_3334,N_2789,N_2570);
nand U3335 (N_3335,N_2945,N_2876);
xor U3336 (N_3336,N_2637,N_2792);
nor U3337 (N_3337,N_2919,N_2878);
nand U3338 (N_3338,N_2679,N_2741);
nand U3339 (N_3339,N_2876,N_2841);
nand U3340 (N_3340,N_2579,N_2888);
and U3341 (N_3341,N_2746,N_2823);
nor U3342 (N_3342,N_2906,N_2812);
and U3343 (N_3343,N_2620,N_2888);
xor U3344 (N_3344,N_2707,N_2545);
xnor U3345 (N_3345,N_2531,N_2632);
xor U3346 (N_3346,N_2533,N_2978);
xor U3347 (N_3347,N_2505,N_2538);
nand U3348 (N_3348,N_2621,N_2915);
nand U3349 (N_3349,N_2804,N_2557);
and U3350 (N_3350,N_2583,N_2928);
nor U3351 (N_3351,N_2994,N_2606);
xor U3352 (N_3352,N_2918,N_2906);
or U3353 (N_3353,N_2866,N_2963);
nor U3354 (N_3354,N_2832,N_2698);
nand U3355 (N_3355,N_2565,N_2937);
nand U3356 (N_3356,N_2908,N_2950);
nand U3357 (N_3357,N_2895,N_2873);
nor U3358 (N_3358,N_2861,N_2937);
nand U3359 (N_3359,N_2903,N_2509);
nand U3360 (N_3360,N_2768,N_2760);
or U3361 (N_3361,N_2819,N_2637);
nor U3362 (N_3362,N_2622,N_2819);
xor U3363 (N_3363,N_2791,N_2658);
or U3364 (N_3364,N_2731,N_2910);
nor U3365 (N_3365,N_2942,N_2910);
and U3366 (N_3366,N_2797,N_2634);
and U3367 (N_3367,N_2795,N_2892);
xor U3368 (N_3368,N_2577,N_2669);
nor U3369 (N_3369,N_2976,N_2564);
nand U3370 (N_3370,N_2622,N_2682);
nor U3371 (N_3371,N_2681,N_2743);
and U3372 (N_3372,N_2593,N_2662);
and U3373 (N_3373,N_2885,N_2633);
nor U3374 (N_3374,N_2556,N_2613);
xor U3375 (N_3375,N_2506,N_2805);
nor U3376 (N_3376,N_2867,N_2954);
nor U3377 (N_3377,N_2906,N_2917);
nand U3378 (N_3378,N_2560,N_2523);
nor U3379 (N_3379,N_2538,N_2567);
or U3380 (N_3380,N_2929,N_2999);
and U3381 (N_3381,N_2872,N_2693);
nand U3382 (N_3382,N_2734,N_2863);
nor U3383 (N_3383,N_2659,N_2533);
or U3384 (N_3384,N_2513,N_2745);
xnor U3385 (N_3385,N_2807,N_2800);
nand U3386 (N_3386,N_2942,N_2739);
xor U3387 (N_3387,N_2555,N_2743);
nor U3388 (N_3388,N_2642,N_2636);
nand U3389 (N_3389,N_2649,N_2648);
and U3390 (N_3390,N_2967,N_2762);
xor U3391 (N_3391,N_2503,N_2665);
xnor U3392 (N_3392,N_2764,N_2916);
nand U3393 (N_3393,N_2784,N_2634);
or U3394 (N_3394,N_2816,N_2672);
or U3395 (N_3395,N_2811,N_2561);
xor U3396 (N_3396,N_2994,N_2889);
or U3397 (N_3397,N_2957,N_2693);
nor U3398 (N_3398,N_2688,N_2685);
nand U3399 (N_3399,N_2962,N_2557);
xor U3400 (N_3400,N_2690,N_2520);
nand U3401 (N_3401,N_2789,N_2983);
nor U3402 (N_3402,N_2588,N_2867);
xnor U3403 (N_3403,N_2576,N_2857);
xor U3404 (N_3404,N_2776,N_2870);
xnor U3405 (N_3405,N_2707,N_2962);
and U3406 (N_3406,N_2970,N_2617);
xor U3407 (N_3407,N_2610,N_2810);
xor U3408 (N_3408,N_2623,N_2773);
nand U3409 (N_3409,N_2657,N_2540);
or U3410 (N_3410,N_2846,N_2953);
nor U3411 (N_3411,N_2867,N_2615);
xor U3412 (N_3412,N_2526,N_2925);
and U3413 (N_3413,N_2693,N_2641);
xor U3414 (N_3414,N_2710,N_2604);
nand U3415 (N_3415,N_2735,N_2589);
and U3416 (N_3416,N_2644,N_2535);
xor U3417 (N_3417,N_2841,N_2822);
or U3418 (N_3418,N_2948,N_2776);
nor U3419 (N_3419,N_2701,N_2930);
and U3420 (N_3420,N_2861,N_2565);
and U3421 (N_3421,N_2950,N_2990);
xor U3422 (N_3422,N_2756,N_2946);
nor U3423 (N_3423,N_2624,N_2984);
nor U3424 (N_3424,N_2839,N_2652);
nor U3425 (N_3425,N_2778,N_2637);
xor U3426 (N_3426,N_2607,N_2614);
xnor U3427 (N_3427,N_2512,N_2942);
and U3428 (N_3428,N_2605,N_2822);
nand U3429 (N_3429,N_2648,N_2825);
xor U3430 (N_3430,N_2568,N_2788);
and U3431 (N_3431,N_2899,N_2997);
nand U3432 (N_3432,N_2876,N_2844);
xor U3433 (N_3433,N_2610,N_2503);
nor U3434 (N_3434,N_2697,N_2578);
and U3435 (N_3435,N_2792,N_2540);
nand U3436 (N_3436,N_2861,N_2710);
nor U3437 (N_3437,N_2659,N_2782);
and U3438 (N_3438,N_2960,N_2514);
nor U3439 (N_3439,N_2539,N_2996);
nand U3440 (N_3440,N_2653,N_2785);
xor U3441 (N_3441,N_2623,N_2513);
xor U3442 (N_3442,N_2661,N_2663);
nand U3443 (N_3443,N_2578,N_2501);
or U3444 (N_3444,N_2812,N_2535);
nor U3445 (N_3445,N_2650,N_2817);
xor U3446 (N_3446,N_2505,N_2953);
and U3447 (N_3447,N_2855,N_2955);
xnor U3448 (N_3448,N_2889,N_2921);
xnor U3449 (N_3449,N_2654,N_2669);
and U3450 (N_3450,N_2772,N_2837);
and U3451 (N_3451,N_2953,N_2652);
or U3452 (N_3452,N_2789,N_2644);
and U3453 (N_3453,N_2726,N_2823);
xor U3454 (N_3454,N_2890,N_2693);
nor U3455 (N_3455,N_2779,N_2709);
xor U3456 (N_3456,N_2578,N_2824);
xor U3457 (N_3457,N_2919,N_2809);
and U3458 (N_3458,N_2789,N_2834);
and U3459 (N_3459,N_2566,N_2685);
or U3460 (N_3460,N_2885,N_2872);
or U3461 (N_3461,N_2767,N_2594);
nor U3462 (N_3462,N_2521,N_2751);
nor U3463 (N_3463,N_2700,N_2598);
and U3464 (N_3464,N_2809,N_2565);
and U3465 (N_3465,N_2608,N_2663);
and U3466 (N_3466,N_2553,N_2807);
or U3467 (N_3467,N_2565,N_2951);
xnor U3468 (N_3468,N_2901,N_2604);
nor U3469 (N_3469,N_2700,N_2816);
nand U3470 (N_3470,N_2738,N_2845);
and U3471 (N_3471,N_2899,N_2606);
and U3472 (N_3472,N_2725,N_2899);
and U3473 (N_3473,N_2599,N_2536);
and U3474 (N_3474,N_2687,N_2594);
xor U3475 (N_3475,N_2779,N_2865);
and U3476 (N_3476,N_2821,N_2723);
nor U3477 (N_3477,N_2513,N_2777);
xor U3478 (N_3478,N_2562,N_2573);
xor U3479 (N_3479,N_2959,N_2580);
xor U3480 (N_3480,N_2651,N_2508);
nor U3481 (N_3481,N_2757,N_2749);
or U3482 (N_3482,N_2532,N_2876);
nor U3483 (N_3483,N_2862,N_2515);
nor U3484 (N_3484,N_2829,N_2669);
or U3485 (N_3485,N_2993,N_2881);
and U3486 (N_3486,N_2615,N_2822);
or U3487 (N_3487,N_2867,N_2823);
xnor U3488 (N_3488,N_2521,N_2725);
nand U3489 (N_3489,N_2758,N_2967);
nand U3490 (N_3490,N_2642,N_2815);
nand U3491 (N_3491,N_2554,N_2733);
or U3492 (N_3492,N_2926,N_2846);
xor U3493 (N_3493,N_2568,N_2888);
and U3494 (N_3494,N_2616,N_2612);
nor U3495 (N_3495,N_2785,N_2850);
or U3496 (N_3496,N_2841,N_2562);
xnor U3497 (N_3497,N_2807,N_2660);
or U3498 (N_3498,N_2869,N_2558);
nand U3499 (N_3499,N_2947,N_2871);
xnor U3500 (N_3500,N_3004,N_3358);
and U3501 (N_3501,N_3496,N_3447);
or U3502 (N_3502,N_3161,N_3481);
and U3503 (N_3503,N_3178,N_3245);
nor U3504 (N_3504,N_3468,N_3127);
or U3505 (N_3505,N_3373,N_3405);
and U3506 (N_3506,N_3219,N_3132);
and U3507 (N_3507,N_3054,N_3304);
and U3508 (N_3508,N_3267,N_3163);
or U3509 (N_3509,N_3195,N_3118);
nor U3510 (N_3510,N_3317,N_3239);
and U3511 (N_3511,N_3255,N_3439);
nand U3512 (N_3512,N_3353,N_3167);
nand U3513 (N_3513,N_3395,N_3103);
nand U3514 (N_3514,N_3303,N_3284);
nand U3515 (N_3515,N_3370,N_3423);
nor U3516 (N_3516,N_3123,N_3046);
xnor U3517 (N_3517,N_3124,N_3011);
nor U3518 (N_3518,N_3386,N_3055);
or U3519 (N_3519,N_3042,N_3329);
nor U3520 (N_3520,N_3295,N_3384);
xnor U3521 (N_3521,N_3053,N_3250);
nand U3522 (N_3522,N_3360,N_3394);
nand U3523 (N_3523,N_3069,N_3309);
nand U3524 (N_3524,N_3049,N_3265);
and U3525 (N_3525,N_3473,N_3105);
or U3526 (N_3526,N_3474,N_3002);
nand U3527 (N_3527,N_3085,N_3351);
xor U3528 (N_3528,N_3216,N_3442);
nor U3529 (N_3529,N_3153,N_3312);
nand U3530 (N_3530,N_3210,N_3179);
or U3531 (N_3531,N_3410,N_3440);
or U3532 (N_3532,N_3006,N_3414);
and U3533 (N_3533,N_3258,N_3359);
or U3534 (N_3534,N_3252,N_3148);
xor U3535 (N_3535,N_3346,N_3343);
nor U3536 (N_3536,N_3413,N_3285);
or U3537 (N_3537,N_3480,N_3321);
nor U3538 (N_3538,N_3368,N_3154);
nand U3539 (N_3539,N_3288,N_3084);
nor U3540 (N_3540,N_3251,N_3450);
or U3541 (N_3541,N_3269,N_3024);
and U3542 (N_3542,N_3256,N_3398);
nor U3543 (N_3543,N_3418,N_3347);
nor U3544 (N_3544,N_3009,N_3232);
and U3545 (N_3545,N_3490,N_3170);
xnor U3546 (N_3546,N_3478,N_3025);
or U3547 (N_3547,N_3019,N_3455);
xnor U3548 (N_3548,N_3070,N_3488);
nor U3549 (N_3549,N_3198,N_3235);
and U3550 (N_3550,N_3137,N_3104);
nor U3551 (N_3551,N_3102,N_3047);
nor U3552 (N_3552,N_3451,N_3315);
nor U3553 (N_3553,N_3067,N_3086);
or U3554 (N_3554,N_3291,N_3027);
or U3555 (N_3555,N_3248,N_3402);
nand U3556 (N_3556,N_3459,N_3068);
nand U3557 (N_3557,N_3058,N_3409);
xor U3558 (N_3558,N_3445,N_3378);
and U3559 (N_3559,N_3129,N_3032);
or U3560 (N_3560,N_3408,N_3456);
xnor U3561 (N_3561,N_3231,N_3296);
and U3562 (N_3562,N_3131,N_3262);
or U3563 (N_3563,N_3015,N_3390);
xnor U3564 (N_3564,N_3172,N_3101);
nor U3565 (N_3565,N_3354,N_3246);
xor U3566 (N_3566,N_3007,N_3159);
nor U3567 (N_3567,N_3033,N_3357);
nand U3568 (N_3568,N_3164,N_3274);
nand U3569 (N_3569,N_3493,N_3376);
and U3570 (N_3570,N_3145,N_3112);
xnor U3571 (N_3571,N_3377,N_3141);
xnor U3572 (N_3572,N_3319,N_3100);
or U3573 (N_3573,N_3469,N_3362);
or U3574 (N_3574,N_3120,N_3234);
nand U3575 (N_3575,N_3115,N_3472);
nand U3576 (N_3576,N_3106,N_3109);
and U3577 (N_3577,N_3243,N_3200);
xor U3578 (N_3578,N_3114,N_3140);
nand U3579 (N_3579,N_3134,N_3371);
nand U3580 (N_3580,N_3217,N_3090);
and U3581 (N_3581,N_3444,N_3162);
nand U3582 (N_3582,N_3150,N_3318);
or U3583 (N_3583,N_3412,N_3466);
and U3584 (N_3584,N_3177,N_3282);
xor U3585 (N_3585,N_3186,N_3224);
nand U3586 (N_3586,N_3207,N_3041);
or U3587 (N_3587,N_3365,N_3043);
xnor U3588 (N_3588,N_3079,N_3397);
xor U3589 (N_3589,N_3345,N_3151);
and U3590 (N_3590,N_3066,N_3181);
or U3591 (N_3591,N_3021,N_3268);
or U3592 (N_3592,N_3077,N_3196);
and U3593 (N_3593,N_3421,N_3372);
nand U3594 (N_3594,N_3475,N_3254);
nor U3595 (N_3595,N_3333,N_3157);
and U3596 (N_3596,N_3453,N_3454);
nand U3597 (N_3597,N_3095,N_3119);
xnor U3598 (N_3598,N_3283,N_3197);
or U3599 (N_3599,N_3193,N_3272);
nand U3600 (N_3600,N_3208,N_3143);
nor U3601 (N_3601,N_3460,N_3449);
and U3602 (N_3602,N_3199,N_3188);
and U3603 (N_3603,N_3314,N_3320);
nor U3604 (N_3604,N_3223,N_3367);
and U3605 (N_3605,N_3416,N_3470);
xnor U3606 (N_3606,N_3341,N_3051);
nor U3607 (N_3607,N_3215,N_3204);
xnor U3608 (N_3608,N_3273,N_3180);
and U3609 (N_3609,N_3206,N_3281);
xor U3610 (N_3610,N_3301,N_3044);
nor U3611 (N_3611,N_3498,N_3093);
and U3612 (N_3612,N_3436,N_3429);
nor U3613 (N_3613,N_3125,N_3014);
and U3614 (N_3614,N_3494,N_3108);
nor U3615 (N_3615,N_3016,N_3146);
nor U3616 (N_3616,N_3165,N_3420);
xnor U3617 (N_3617,N_3432,N_3270);
xor U3618 (N_3618,N_3383,N_3411);
xnor U3619 (N_3619,N_3244,N_3316);
nand U3620 (N_3620,N_3363,N_3342);
and U3621 (N_3621,N_3430,N_3205);
nor U3622 (N_3622,N_3417,N_3324);
nand U3623 (N_3623,N_3415,N_3082);
nor U3624 (N_3624,N_3489,N_3184);
or U3625 (N_3625,N_3030,N_3220);
and U3626 (N_3626,N_3203,N_3361);
or U3627 (N_3627,N_3116,N_3407);
xor U3628 (N_3628,N_3052,N_3128);
or U3629 (N_3629,N_3117,N_3168);
xor U3630 (N_3630,N_3001,N_3097);
nor U3631 (N_3631,N_3308,N_3448);
xnor U3632 (N_3632,N_3374,N_3160);
xnor U3633 (N_3633,N_3158,N_3213);
xnor U3634 (N_3634,N_3393,N_3144);
nand U3635 (N_3635,N_3326,N_3352);
and U3636 (N_3636,N_3458,N_3214);
nand U3637 (N_3637,N_3406,N_3392);
xnor U3638 (N_3638,N_3031,N_3350);
nand U3639 (N_3639,N_3096,N_3428);
nor U3640 (N_3640,N_3422,N_3382);
and U3641 (N_3641,N_3380,N_3266);
xor U3642 (N_3642,N_3045,N_3107);
xnor U3643 (N_3643,N_3228,N_3280);
nand U3644 (N_3644,N_3322,N_3292);
or U3645 (N_3645,N_3388,N_3387);
xnor U3646 (N_3646,N_3483,N_3133);
nand U3647 (N_3647,N_3190,N_3189);
and U3648 (N_3648,N_3149,N_3089);
nand U3649 (N_3649,N_3065,N_3221);
nor U3650 (N_3650,N_3139,N_3340);
xor U3651 (N_3651,N_3113,N_3187);
and U3652 (N_3652,N_3048,N_3401);
nor U3653 (N_3653,N_3039,N_3355);
nand U3654 (N_3654,N_3135,N_3438);
nand U3655 (N_3655,N_3479,N_3330);
nor U3656 (N_3656,N_3003,N_3130);
xnor U3657 (N_3657,N_3344,N_3110);
and U3658 (N_3658,N_3237,N_3400);
or U3659 (N_3659,N_3297,N_3443);
xor U3660 (N_3660,N_3306,N_3183);
nand U3661 (N_3661,N_3491,N_3427);
or U3662 (N_3662,N_3328,N_3484);
xnor U3663 (N_3663,N_3062,N_3111);
nand U3664 (N_3664,N_3092,N_3476);
nand U3665 (N_3665,N_3310,N_3486);
nand U3666 (N_3666,N_3076,N_3307);
nand U3667 (N_3667,N_3034,N_3461);
nand U3668 (N_3668,N_3075,N_3121);
nand U3669 (N_3669,N_3467,N_3081);
or U3670 (N_3670,N_3294,N_3477);
nand U3671 (N_3671,N_3336,N_3389);
or U3672 (N_3672,N_3040,N_3099);
xor U3673 (N_3673,N_3169,N_3356);
nand U3674 (N_3674,N_3156,N_3492);
and U3675 (N_3675,N_3441,N_3012);
nor U3676 (N_3676,N_3375,N_3175);
xor U3677 (N_3677,N_3264,N_3211);
and U3678 (N_3678,N_3038,N_3334);
nand U3679 (N_3679,N_3259,N_3257);
nand U3680 (N_3680,N_3080,N_3457);
xor U3681 (N_3681,N_3059,N_3325);
nand U3682 (N_3682,N_3300,N_3202);
and U3683 (N_3683,N_3277,N_3072);
or U3684 (N_3684,N_3174,N_3236);
or U3685 (N_3685,N_3233,N_3299);
xnor U3686 (N_3686,N_3403,N_3385);
and U3687 (N_3687,N_3289,N_3419);
and U3688 (N_3688,N_3227,N_3173);
nand U3689 (N_3689,N_3229,N_3074);
and U3690 (N_3690,N_3017,N_3305);
xnor U3691 (N_3691,N_3396,N_3018);
or U3692 (N_3692,N_3276,N_3176);
or U3693 (N_3693,N_3242,N_3087);
and U3694 (N_3694,N_3426,N_3126);
nand U3695 (N_3695,N_3327,N_3369);
and U3696 (N_3696,N_3286,N_3253);
xor U3697 (N_3697,N_3035,N_3434);
and U3698 (N_3698,N_3263,N_3366);
and U3699 (N_3699,N_3194,N_3147);
and U3700 (N_3700,N_3379,N_3060);
xor U3701 (N_3701,N_3339,N_3391);
and U3702 (N_3702,N_3138,N_3098);
or U3703 (N_3703,N_3249,N_3349);
nor U3704 (N_3704,N_3381,N_3332);
nor U3705 (N_3705,N_3290,N_3495);
or U3706 (N_3706,N_3094,N_3485);
nor U3707 (N_3707,N_3050,N_3425);
xnor U3708 (N_3708,N_3071,N_3013);
nor U3709 (N_3709,N_3302,N_3424);
nor U3710 (N_3710,N_3008,N_3298);
nand U3711 (N_3711,N_3348,N_3287);
or U3712 (N_3712,N_3499,N_3010);
nor U3713 (N_3713,N_3240,N_3311);
xor U3714 (N_3714,N_3142,N_3061);
xor U3715 (N_3715,N_3446,N_3364);
xnor U3716 (N_3716,N_3078,N_3225);
nor U3717 (N_3717,N_3192,N_3404);
nand U3718 (N_3718,N_3023,N_3020);
xor U3719 (N_3719,N_3230,N_3260);
nor U3720 (N_3720,N_3088,N_3122);
and U3721 (N_3721,N_3191,N_3155);
nor U3722 (N_3722,N_3064,N_3029);
nand U3723 (N_3723,N_3338,N_3497);
nand U3724 (N_3724,N_3222,N_3218);
nand U3725 (N_3725,N_3331,N_3226);
nor U3726 (N_3726,N_3185,N_3293);
and U3727 (N_3727,N_3022,N_3279);
xor U3728 (N_3728,N_3136,N_3152);
nand U3729 (N_3729,N_3471,N_3431);
nor U3730 (N_3730,N_3337,N_3437);
nand U3731 (N_3731,N_3487,N_3026);
nor U3732 (N_3732,N_3212,N_3462);
nand U3733 (N_3733,N_3463,N_3166);
or U3734 (N_3734,N_3201,N_3209);
nand U3735 (N_3735,N_3482,N_3063);
and U3736 (N_3736,N_3083,N_3323);
nor U3737 (N_3737,N_3238,N_3056);
and U3738 (N_3738,N_3091,N_3452);
nor U3739 (N_3739,N_3335,N_3000);
nor U3740 (N_3740,N_3278,N_3057);
xnor U3741 (N_3741,N_3073,N_3028);
xnor U3742 (N_3742,N_3433,N_3271);
nor U3743 (N_3743,N_3465,N_3036);
and U3744 (N_3744,N_3182,N_3037);
and U3745 (N_3745,N_3313,N_3464);
and U3746 (N_3746,N_3005,N_3247);
nor U3747 (N_3747,N_3171,N_3261);
xnor U3748 (N_3748,N_3275,N_3399);
nand U3749 (N_3749,N_3435,N_3241);
and U3750 (N_3750,N_3221,N_3041);
and U3751 (N_3751,N_3434,N_3357);
nand U3752 (N_3752,N_3342,N_3008);
nand U3753 (N_3753,N_3285,N_3210);
or U3754 (N_3754,N_3279,N_3442);
or U3755 (N_3755,N_3439,N_3469);
xor U3756 (N_3756,N_3476,N_3086);
nor U3757 (N_3757,N_3250,N_3352);
and U3758 (N_3758,N_3012,N_3123);
xnor U3759 (N_3759,N_3459,N_3479);
nor U3760 (N_3760,N_3469,N_3228);
and U3761 (N_3761,N_3015,N_3181);
nor U3762 (N_3762,N_3341,N_3012);
xor U3763 (N_3763,N_3498,N_3012);
nor U3764 (N_3764,N_3330,N_3453);
or U3765 (N_3765,N_3150,N_3305);
xor U3766 (N_3766,N_3284,N_3013);
or U3767 (N_3767,N_3309,N_3253);
nand U3768 (N_3768,N_3357,N_3091);
xnor U3769 (N_3769,N_3062,N_3307);
and U3770 (N_3770,N_3250,N_3330);
and U3771 (N_3771,N_3137,N_3477);
nor U3772 (N_3772,N_3129,N_3156);
or U3773 (N_3773,N_3408,N_3227);
or U3774 (N_3774,N_3098,N_3205);
xnor U3775 (N_3775,N_3457,N_3182);
and U3776 (N_3776,N_3383,N_3486);
nor U3777 (N_3777,N_3415,N_3385);
and U3778 (N_3778,N_3367,N_3444);
nor U3779 (N_3779,N_3410,N_3064);
xor U3780 (N_3780,N_3131,N_3289);
or U3781 (N_3781,N_3255,N_3253);
xor U3782 (N_3782,N_3013,N_3464);
and U3783 (N_3783,N_3091,N_3088);
xnor U3784 (N_3784,N_3220,N_3295);
and U3785 (N_3785,N_3249,N_3373);
nor U3786 (N_3786,N_3180,N_3371);
nor U3787 (N_3787,N_3348,N_3314);
xor U3788 (N_3788,N_3219,N_3098);
nor U3789 (N_3789,N_3056,N_3062);
or U3790 (N_3790,N_3413,N_3431);
nor U3791 (N_3791,N_3497,N_3046);
nand U3792 (N_3792,N_3309,N_3163);
xor U3793 (N_3793,N_3152,N_3441);
nor U3794 (N_3794,N_3080,N_3342);
or U3795 (N_3795,N_3398,N_3074);
xnor U3796 (N_3796,N_3454,N_3270);
nor U3797 (N_3797,N_3433,N_3338);
and U3798 (N_3798,N_3334,N_3130);
xnor U3799 (N_3799,N_3270,N_3061);
or U3800 (N_3800,N_3278,N_3170);
or U3801 (N_3801,N_3474,N_3259);
xor U3802 (N_3802,N_3194,N_3120);
or U3803 (N_3803,N_3150,N_3208);
nand U3804 (N_3804,N_3394,N_3074);
nor U3805 (N_3805,N_3221,N_3222);
or U3806 (N_3806,N_3033,N_3417);
xor U3807 (N_3807,N_3012,N_3117);
nand U3808 (N_3808,N_3203,N_3305);
and U3809 (N_3809,N_3017,N_3054);
and U3810 (N_3810,N_3463,N_3068);
nor U3811 (N_3811,N_3250,N_3203);
and U3812 (N_3812,N_3241,N_3144);
nor U3813 (N_3813,N_3434,N_3094);
nor U3814 (N_3814,N_3450,N_3144);
nand U3815 (N_3815,N_3220,N_3422);
xnor U3816 (N_3816,N_3311,N_3226);
and U3817 (N_3817,N_3463,N_3491);
nor U3818 (N_3818,N_3004,N_3110);
nor U3819 (N_3819,N_3185,N_3103);
xnor U3820 (N_3820,N_3116,N_3099);
nand U3821 (N_3821,N_3256,N_3062);
xnor U3822 (N_3822,N_3016,N_3392);
nand U3823 (N_3823,N_3320,N_3274);
nor U3824 (N_3824,N_3119,N_3254);
or U3825 (N_3825,N_3250,N_3001);
nor U3826 (N_3826,N_3362,N_3393);
nand U3827 (N_3827,N_3425,N_3261);
nand U3828 (N_3828,N_3098,N_3143);
and U3829 (N_3829,N_3419,N_3425);
xnor U3830 (N_3830,N_3317,N_3006);
nand U3831 (N_3831,N_3103,N_3031);
nand U3832 (N_3832,N_3403,N_3020);
nand U3833 (N_3833,N_3304,N_3473);
nand U3834 (N_3834,N_3370,N_3457);
nand U3835 (N_3835,N_3365,N_3002);
and U3836 (N_3836,N_3182,N_3079);
or U3837 (N_3837,N_3475,N_3184);
nor U3838 (N_3838,N_3097,N_3205);
nand U3839 (N_3839,N_3297,N_3183);
or U3840 (N_3840,N_3198,N_3136);
nor U3841 (N_3841,N_3493,N_3112);
or U3842 (N_3842,N_3452,N_3023);
xor U3843 (N_3843,N_3324,N_3322);
or U3844 (N_3844,N_3108,N_3233);
nor U3845 (N_3845,N_3433,N_3258);
nand U3846 (N_3846,N_3253,N_3290);
and U3847 (N_3847,N_3264,N_3184);
nor U3848 (N_3848,N_3167,N_3256);
nor U3849 (N_3849,N_3356,N_3387);
xnor U3850 (N_3850,N_3158,N_3003);
nand U3851 (N_3851,N_3020,N_3155);
and U3852 (N_3852,N_3351,N_3277);
and U3853 (N_3853,N_3260,N_3032);
and U3854 (N_3854,N_3345,N_3260);
xor U3855 (N_3855,N_3468,N_3405);
xnor U3856 (N_3856,N_3126,N_3054);
nor U3857 (N_3857,N_3311,N_3054);
and U3858 (N_3858,N_3238,N_3033);
xor U3859 (N_3859,N_3114,N_3287);
xor U3860 (N_3860,N_3224,N_3288);
xnor U3861 (N_3861,N_3078,N_3418);
nand U3862 (N_3862,N_3300,N_3135);
nand U3863 (N_3863,N_3398,N_3494);
xor U3864 (N_3864,N_3261,N_3217);
nand U3865 (N_3865,N_3264,N_3404);
nand U3866 (N_3866,N_3400,N_3444);
nor U3867 (N_3867,N_3495,N_3307);
nor U3868 (N_3868,N_3209,N_3004);
nand U3869 (N_3869,N_3427,N_3315);
nand U3870 (N_3870,N_3027,N_3117);
and U3871 (N_3871,N_3157,N_3161);
nor U3872 (N_3872,N_3441,N_3406);
or U3873 (N_3873,N_3427,N_3286);
or U3874 (N_3874,N_3268,N_3285);
and U3875 (N_3875,N_3267,N_3479);
and U3876 (N_3876,N_3039,N_3395);
or U3877 (N_3877,N_3346,N_3153);
or U3878 (N_3878,N_3200,N_3264);
nand U3879 (N_3879,N_3161,N_3431);
or U3880 (N_3880,N_3482,N_3450);
xnor U3881 (N_3881,N_3080,N_3095);
nor U3882 (N_3882,N_3485,N_3351);
and U3883 (N_3883,N_3307,N_3366);
or U3884 (N_3884,N_3302,N_3303);
nand U3885 (N_3885,N_3085,N_3456);
or U3886 (N_3886,N_3462,N_3372);
xor U3887 (N_3887,N_3153,N_3099);
nand U3888 (N_3888,N_3028,N_3243);
nand U3889 (N_3889,N_3449,N_3261);
nand U3890 (N_3890,N_3454,N_3152);
or U3891 (N_3891,N_3055,N_3178);
nor U3892 (N_3892,N_3411,N_3227);
nor U3893 (N_3893,N_3354,N_3127);
nor U3894 (N_3894,N_3188,N_3494);
and U3895 (N_3895,N_3329,N_3277);
xor U3896 (N_3896,N_3406,N_3096);
and U3897 (N_3897,N_3226,N_3139);
or U3898 (N_3898,N_3443,N_3374);
nand U3899 (N_3899,N_3432,N_3104);
nor U3900 (N_3900,N_3256,N_3350);
and U3901 (N_3901,N_3236,N_3296);
nor U3902 (N_3902,N_3330,N_3059);
and U3903 (N_3903,N_3120,N_3213);
or U3904 (N_3904,N_3415,N_3435);
nor U3905 (N_3905,N_3344,N_3277);
nand U3906 (N_3906,N_3259,N_3080);
nor U3907 (N_3907,N_3291,N_3477);
nand U3908 (N_3908,N_3431,N_3015);
nor U3909 (N_3909,N_3492,N_3374);
or U3910 (N_3910,N_3246,N_3406);
nand U3911 (N_3911,N_3077,N_3113);
nor U3912 (N_3912,N_3245,N_3265);
nor U3913 (N_3913,N_3400,N_3378);
nand U3914 (N_3914,N_3296,N_3080);
or U3915 (N_3915,N_3270,N_3444);
xnor U3916 (N_3916,N_3167,N_3334);
or U3917 (N_3917,N_3029,N_3014);
nor U3918 (N_3918,N_3407,N_3095);
nand U3919 (N_3919,N_3043,N_3100);
and U3920 (N_3920,N_3379,N_3365);
or U3921 (N_3921,N_3091,N_3258);
nor U3922 (N_3922,N_3332,N_3459);
and U3923 (N_3923,N_3342,N_3425);
and U3924 (N_3924,N_3459,N_3225);
xor U3925 (N_3925,N_3256,N_3356);
nand U3926 (N_3926,N_3333,N_3438);
nand U3927 (N_3927,N_3202,N_3010);
and U3928 (N_3928,N_3203,N_3056);
nor U3929 (N_3929,N_3358,N_3108);
nand U3930 (N_3930,N_3341,N_3149);
xnor U3931 (N_3931,N_3301,N_3172);
nor U3932 (N_3932,N_3210,N_3206);
xor U3933 (N_3933,N_3018,N_3071);
nand U3934 (N_3934,N_3287,N_3357);
and U3935 (N_3935,N_3052,N_3155);
or U3936 (N_3936,N_3019,N_3420);
or U3937 (N_3937,N_3054,N_3241);
and U3938 (N_3938,N_3104,N_3173);
xor U3939 (N_3939,N_3105,N_3049);
xor U3940 (N_3940,N_3126,N_3176);
and U3941 (N_3941,N_3308,N_3414);
or U3942 (N_3942,N_3241,N_3114);
or U3943 (N_3943,N_3008,N_3362);
nand U3944 (N_3944,N_3309,N_3453);
or U3945 (N_3945,N_3366,N_3249);
and U3946 (N_3946,N_3427,N_3006);
or U3947 (N_3947,N_3131,N_3430);
or U3948 (N_3948,N_3390,N_3458);
nand U3949 (N_3949,N_3388,N_3164);
or U3950 (N_3950,N_3195,N_3391);
nor U3951 (N_3951,N_3381,N_3018);
xor U3952 (N_3952,N_3154,N_3214);
nand U3953 (N_3953,N_3381,N_3088);
nor U3954 (N_3954,N_3036,N_3094);
and U3955 (N_3955,N_3159,N_3073);
and U3956 (N_3956,N_3122,N_3135);
xor U3957 (N_3957,N_3483,N_3416);
or U3958 (N_3958,N_3457,N_3385);
nand U3959 (N_3959,N_3038,N_3110);
and U3960 (N_3960,N_3332,N_3366);
nand U3961 (N_3961,N_3401,N_3415);
xnor U3962 (N_3962,N_3339,N_3447);
nor U3963 (N_3963,N_3177,N_3469);
xnor U3964 (N_3964,N_3157,N_3391);
or U3965 (N_3965,N_3406,N_3130);
or U3966 (N_3966,N_3205,N_3328);
or U3967 (N_3967,N_3340,N_3367);
or U3968 (N_3968,N_3210,N_3052);
nand U3969 (N_3969,N_3335,N_3169);
nand U3970 (N_3970,N_3378,N_3184);
nor U3971 (N_3971,N_3195,N_3085);
or U3972 (N_3972,N_3079,N_3418);
nand U3973 (N_3973,N_3488,N_3395);
and U3974 (N_3974,N_3231,N_3457);
nor U3975 (N_3975,N_3281,N_3243);
xor U3976 (N_3976,N_3158,N_3437);
nand U3977 (N_3977,N_3098,N_3060);
and U3978 (N_3978,N_3314,N_3162);
or U3979 (N_3979,N_3343,N_3102);
xor U3980 (N_3980,N_3402,N_3404);
or U3981 (N_3981,N_3475,N_3403);
nand U3982 (N_3982,N_3229,N_3414);
nor U3983 (N_3983,N_3147,N_3439);
and U3984 (N_3984,N_3461,N_3106);
xor U3985 (N_3985,N_3404,N_3439);
and U3986 (N_3986,N_3139,N_3356);
or U3987 (N_3987,N_3493,N_3012);
nor U3988 (N_3988,N_3197,N_3238);
nor U3989 (N_3989,N_3031,N_3121);
xnor U3990 (N_3990,N_3417,N_3132);
nand U3991 (N_3991,N_3029,N_3004);
or U3992 (N_3992,N_3284,N_3359);
nor U3993 (N_3993,N_3444,N_3421);
or U3994 (N_3994,N_3159,N_3162);
or U3995 (N_3995,N_3231,N_3453);
and U3996 (N_3996,N_3475,N_3304);
nand U3997 (N_3997,N_3012,N_3470);
nor U3998 (N_3998,N_3203,N_3270);
or U3999 (N_3999,N_3060,N_3164);
nand U4000 (N_4000,N_3705,N_3638);
or U4001 (N_4001,N_3525,N_3701);
nor U4002 (N_4002,N_3874,N_3587);
nand U4003 (N_4003,N_3500,N_3650);
and U4004 (N_4004,N_3858,N_3846);
nand U4005 (N_4005,N_3516,N_3967);
xnor U4006 (N_4006,N_3850,N_3855);
or U4007 (N_4007,N_3821,N_3983);
and U4008 (N_4008,N_3753,N_3656);
or U4009 (N_4009,N_3907,N_3839);
xnor U4010 (N_4010,N_3621,N_3976);
nand U4011 (N_4011,N_3805,N_3767);
nor U4012 (N_4012,N_3684,N_3580);
nand U4013 (N_4013,N_3643,N_3704);
or U4014 (N_4014,N_3849,N_3848);
or U4015 (N_4015,N_3870,N_3790);
nor U4016 (N_4016,N_3997,N_3810);
and U4017 (N_4017,N_3714,N_3977);
nand U4018 (N_4018,N_3632,N_3744);
and U4019 (N_4019,N_3601,N_3694);
and U4020 (N_4020,N_3964,N_3854);
nand U4021 (N_4021,N_3519,N_3702);
nor U4022 (N_4022,N_3865,N_3573);
or U4023 (N_4023,N_3813,N_3824);
and U4024 (N_4024,N_3512,N_3737);
xnor U4025 (N_4025,N_3706,N_3970);
or U4026 (N_4026,N_3615,N_3528);
nor U4027 (N_4027,N_3623,N_3537);
xnor U4028 (N_4028,N_3642,N_3772);
xor U4029 (N_4029,N_3777,N_3722);
and U4030 (N_4030,N_3914,N_3838);
nand U4031 (N_4031,N_3734,N_3610);
or U4032 (N_4032,N_3872,N_3775);
nand U4033 (N_4033,N_3984,N_3857);
and U4034 (N_4034,N_3604,N_3646);
and U4035 (N_4035,N_3598,N_3718);
xnor U4036 (N_4036,N_3513,N_3617);
nor U4037 (N_4037,N_3585,N_3928);
xnor U4038 (N_4038,N_3531,N_3963);
or U4039 (N_4039,N_3745,N_3711);
nor U4040 (N_4040,N_3916,N_3940);
xnor U4041 (N_4041,N_3817,N_3904);
and U4042 (N_4042,N_3504,N_3524);
and U4043 (N_4043,N_3756,N_3981);
and U4044 (N_4044,N_3933,N_3719);
nand U4045 (N_4045,N_3811,N_3797);
nor U4046 (N_4046,N_3826,N_3809);
xnor U4047 (N_4047,N_3781,N_3716);
nand U4048 (N_4048,N_3842,N_3888);
nor U4049 (N_4049,N_3886,N_3629);
nor U4050 (N_4050,N_3517,N_3724);
and U4051 (N_4051,N_3686,N_3551);
or U4052 (N_4052,N_3560,N_3910);
nand U4053 (N_4053,N_3890,N_3565);
nand U4054 (N_4054,N_3644,N_3979);
and U4055 (N_4055,N_3978,N_3900);
nor U4056 (N_4056,N_3553,N_3789);
or U4057 (N_4057,N_3840,N_3721);
or U4058 (N_4058,N_3577,N_3628);
nand U4059 (N_4059,N_3815,N_3653);
nor U4060 (N_4060,N_3785,N_3699);
nand U4061 (N_4061,N_3540,N_3994);
or U4062 (N_4062,N_3582,N_3627);
and U4063 (N_4063,N_3959,N_3903);
or U4064 (N_4064,N_3796,N_3990);
or U4065 (N_4065,N_3827,N_3541);
nor U4066 (N_4066,N_3735,N_3507);
nor U4067 (N_4067,N_3556,N_3662);
nor U4068 (N_4068,N_3947,N_3901);
nor U4069 (N_4069,N_3602,N_3866);
and U4070 (N_4070,N_3639,N_3511);
nand U4071 (N_4071,N_3521,N_3503);
and U4072 (N_4072,N_3955,N_3931);
or U4073 (N_4073,N_3668,N_3989);
nand U4074 (N_4074,N_3812,N_3946);
xnor U4075 (N_4075,N_3912,N_3712);
nand U4076 (N_4076,N_3759,N_3829);
or U4077 (N_4077,N_3841,N_3885);
nand U4078 (N_4078,N_3856,N_3864);
xnor U4079 (N_4079,N_3729,N_3820);
or U4080 (N_4080,N_3895,N_3637);
nor U4081 (N_4081,N_3526,N_3697);
nand U4082 (N_4082,N_3869,N_3625);
or U4083 (N_4083,N_3852,N_3794);
nor U4084 (N_4084,N_3581,N_3835);
or U4085 (N_4085,N_3715,N_3562);
or U4086 (N_4086,N_3986,N_3793);
or U4087 (N_4087,N_3927,N_3645);
and U4088 (N_4088,N_3816,N_3879);
and U4089 (N_4089,N_3802,N_3633);
or U4090 (N_4090,N_3570,N_3666);
or U4091 (N_4091,N_3825,N_3937);
and U4092 (N_4092,N_3923,N_3619);
or U4093 (N_4093,N_3593,N_3698);
and U4094 (N_4094,N_3635,N_3607);
nor U4095 (N_4095,N_3682,N_3616);
or U4096 (N_4096,N_3762,N_3834);
nand U4097 (N_4097,N_3943,N_3634);
xnor U4098 (N_4098,N_3761,N_3655);
and U4099 (N_4099,N_3932,N_3594);
and U4100 (N_4100,N_3938,N_3542);
nand U4101 (N_4101,N_3731,N_3717);
nand U4102 (N_4102,N_3787,N_3550);
xor U4103 (N_4103,N_3768,N_3993);
and U4104 (N_4104,N_3893,N_3754);
nor U4105 (N_4105,N_3693,N_3544);
nor U4106 (N_4106,N_3514,N_3522);
and U4107 (N_4107,N_3863,N_3720);
xor U4108 (N_4108,N_3539,N_3784);
nand U4109 (N_4109,N_3620,N_3626);
and U4110 (N_4110,N_3660,N_3678);
and U4111 (N_4111,N_3742,N_3700);
nand U4112 (N_4112,N_3774,N_3867);
or U4113 (N_4113,N_3683,N_3941);
nor U4114 (N_4114,N_3748,N_3680);
xor U4115 (N_4115,N_3992,N_3944);
nand U4116 (N_4116,N_3911,N_3962);
xor U4117 (N_4117,N_3611,N_3728);
or U4118 (N_4118,N_3833,N_3592);
nand U4119 (N_4119,N_3727,N_3501);
and U4120 (N_4120,N_3956,N_3736);
and U4121 (N_4121,N_3534,N_3568);
xnor U4122 (N_4122,N_3533,N_3641);
or U4123 (N_4123,N_3915,N_3887);
xor U4124 (N_4124,N_3764,N_3597);
nand U4125 (N_4125,N_3588,N_3624);
nor U4126 (N_4126,N_3672,N_3792);
and U4127 (N_4127,N_3965,N_3859);
xnor U4128 (N_4128,N_3935,N_3703);
xor U4129 (N_4129,N_3898,N_3523);
or U4130 (N_4130,N_3822,N_3726);
or U4131 (N_4131,N_3558,N_3877);
and U4132 (N_4132,N_3750,N_3640);
nand U4133 (N_4133,N_3770,N_3707);
nor U4134 (N_4134,N_3832,N_3819);
or U4135 (N_4135,N_3599,N_3998);
or U4136 (N_4136,N_3883,N_3747);
nand U4137 (N_4137,N_3807,N_3861);
nand U4138 (N_4138,N_3584,N_3880);
or U4139 (N_4139,N_3926,N_3559);
and U4140 (N_4140,N_3548,N_3687);
nand U4141 (N_4141,N_3782,N_3681);
nor U4142 (N_4142,N_3891,N_3571);
and U4143 (N_4143,N_3689,N_3674);
nand U4144 (N_4144,N_3606,N_3739);
or U4145 (N_4145,N_3974,N_3676);
xnor U4146 (N_4146,N_3892,N_3791);
xnor U4147 (N_4147,N_3949,N_3723);
nand U4148 (N_4148,N_3969,N_3665);
or U4149 (N_4149,N_3612,N_3889);
xnor U4150 (N_4150,N_3740,N_3982);
xnor U4151 (N_4151,N_3980,N_3899);
or U4152 (N_4152,N_3876,N_3806);
and U4153 (N_4153,N_3743,N_3882);
and U4154 (N_4154,N_3613,N_3710);
nand U4155 (N_4155,N_3590,N_3661);
or U4156 (N_4156,N_3913,N_3567);
nand U4157 (N_4157,N_3988,N_3520);
nor U4158 (N_4158,N_3690,N_3506);
or U4159 (N_4159,N_3563,N_3948);
or U4160 (N_4160,N_3917,N_3905);
nand U4161 (N_4161,N_3902,N_3614);
or U4162 (N_4162,N_3667,N_3968);
and U4163 (N_4163,N_3725,N_3878);
or U4164 (N_4164,N_3830,N_3545);
nand U4165 (N_4165,N_3897,N_3778);
or U4166 (N_4166,N_3828,N_3975);
xnor U4167 (N_4167,N_3675,N_3589);
and U4168 (N_4168,N_3999,N_3884);
nand U4169 (N_4169,N_3936,N_3942);
and U4170 (N_4170,N_3713,N_3765);
xnor U4171 (N_4171,N_3804,N_3631);
nand U4172 (N_4172,N_3554,N_3773);
xor U4173 (N_4173,N_3508,N_3783);
nor U4174 (N_4174,N_3741,N_3749);
nor U4175 (N_4175,N_3738,N_3795);
nor U4176 (N_4176,N_3799,N_3755);
nor U4177 (N_4177,N_3618,N_3991);
or U4178 (N_4178,N_3871,N_3786);
nor U4179 (N_4179,N_3579,N_3502);
nand U4180 (N_4180,N_3578,N_3847);
or U4181 (N_4181,N_3746,N_3549);
xnor U4182 (N_4182,N_3798,N_3771);
or U4183 (N_4183,N_3909,N_3730);
nor U4184 (N_4184,N_3752,N_3985);
or U4185 (N_4185,N_3538,N_3657);
nor U4186 (N_4186,N_3596,N_3708);
and U4187 (N_4187,N_3875,N_3868);
nand U4188 (N_4188,N_3945,N_3732);
nor U4189 (N_4189,N_3921,N_3677);
xnor U4190 (N_4190,N_3555,N_3966);
xnor U4191 (N_4191,N_3543,N_3605);
nor U4192 (N_4192,N_3803,N_3664);
or U4193 (N_4193,N_3814,N_3801);
xnor U4194 (N_4194,N_3788,N_3961);
or U4195 (N_4195,N_3757,N_3574);
and U4196 (N_4196,N_3603,N_3929);
xnor U4197 (N_4197,N_3557,N_3939);
nor U4198 (N_4198,N_3630,N_3647);
or U4199 (N_4199,N_3987,N_3530);
nand U4200 (N_4200,N_3505,N_3954);
nor U4201 (N_4201,N_3844,N_3649);
or U4202 (N_4202,N_3922,N_3583);
or U4203 (N_4203,N_3836,N_3995);
or U4204 (N_4204,N_3779,N_3695);
nor U4205 (N_4205,N_3566,N_3873);
and U4206 (N_4206,N_3659,N_3860);
nor U4207 (N_4207,N_3532,N_3776);
or U4208 (N_4208,N_3953,N_3595);
nand U4209 (N_4209,N_3851,N_3670);
nor U4210 (N_4210,N_3509,N_3572);
xor U4211 (N_4211,N_3651,N_3823);
nand U4212 (N_4212,N_3853,N_3924);
and U4213 (N_4213,N_3569,N_3818);
nor U4214 (N_4214,N_3685,N_3679);
xnor U4215 (N_4215,N_3957,N_3654);
and U4216 (N_4216,N_3862,N_3609);
and U4217 (N_4217,N_3763,N_3663);
nor U4218 (N_4218,N_3845,N_3951);
nand U4219 (N_4219,N_3600,N_3546);
xor U4220 (N_4220,N_3586,N_3894);
xor U4221 (N_4221,N_3766,N_3510);
or U4222 (N_4222,N_3671,N_3536);
and U4223 (N_4223,N_3648,N_3881);
xnor U4224 (N_4224,N_3733,N_3691);
nand U4225 (N_4225,N_3843,N_3960);
and U4226 (N_4226,N_3971,N_3696);
nand U4227 (N_4227,N_3780,N_3652);
xnor U4228 (N_4228,N_3908,N_3958);
or U4229 (N_4229,N_3527,N_3751);
and U4230 (N_4230,N_3950,N_3658);
nor U4231 (N_4231,N_3996,N_3930);
xnor U4232 (N_4232,N_3688,N_3709);
xor U4233 (N_4233,N_3831,N_3669);
nor U4234 (N_4234,N_3760,N_3952);
or U4235 (N_4235,N_3972,N_3973);
or U4236 (N_4236,N_3515,N_3808);
xor U4237 (N_4237,N_3837,N_3529);
or U4238 (N_4238,N_3561,N_3575);
nor U4239 (N_4239,N_3906,N_3564);
nand U4240 (N_4240,N_3934,N_3800);
xnor U4241 (N_4241,N_3673,N_3591);
nor U4242 (N_4242,N_3552,N_3622);
nand U4243 (N_4243,N_3692,N_3518);
nor U4244 (N_4244,N_3608,N_3925);
or U4245 (N_4245,N_3919,N_3918);
xor U4246 (N_4246,N_3636,N_3758);
nor U4247 (N_4247,N_3535,N_3769);
or U4248 (N_4248,N_3896,N_3547);
and U4249 (N_4249,N_3920,N_3576);
xnor U4250 (N_4250,N_3832,N_3736);
nor U4251 (N_4251,N_3568,N_3918);
and U4252 (N_4252,N_3812,N_3972);
nand U4253 (N_4253,N_3938,N_3755);
and U4254 (N_4254,N_3850,N_3768);
and U4255 (N_4255,N_3611,N_3744);
nor U4256 (N_4256,N_3997,N_3878);
xor U4257 (N_4257,N_3683,N_3899);
and U4258 (N_4258,N_3661,N_3806);
nor U4259 (N_4259,N_3659,N_3585);
nand U4260 (N_4260,N_3775,N_3720);
and U4261 (N_4261,N_3834,N_3899);
or U4262 (N_4262,N_3960,N_3645);
xnor U4263 (N_4263,N_3732,N_3941);
nand U4264 (N_4264,N_3954,N_3571);
xnor U4265 (N_4265,N_3743,N_3535);
nor U4266 (N_4266,N_3755,N_3701);
xor U4267 (N_4267,N_3681,N_3909);
nor U4268 (N_4268,N_3587,N_3847);
xnor U4269 (N_4269,N_3736,N_3629);
and U4270 (N_4270,N_3527,N_3812);
nand U4271 (N_4271,N_3634,N_3864);
nand U4272 (N_4272,N_3529,N_3838);
and U4273 (N_4273,N_3662,N_3891);
or U4274 (N_4274,N_3842,N_3952);
or U4275 (N_4275,N_3714,N_3696);
nand U4276 (N_4276,N_3745,N_3706);
and U4277 (N_4277,N_3912,N_3936);
or U4278 (N_4278,N_3622,N_3947);
xor U4279 (N_4279,N_3934,N_3619);
and U4280 (N_4280,N_3623,N_3538);
nor U4281 (N_4281,N_3953,N_3740);
and U4282 (N_4282,N_3563,N_3846);
nand U4283 (N_4283,N_3681,N_3828);
nand U4284 (N_4284,N_3713,N_3562);
or U4285 (N_4285,N_3909,N_3983);
or U4286 (N_4286,N_3890,N_3789);
nand U4287 (N_4287,N_3792,N_3831);
or U4288 (N_4288,N_3856,N_3797);
nor U4289 (N_4289,N_3931,N_3803);
or U4290 (N_4290,N_3759,N_3651);
nor U4291 (N_4291,N_3764,N_3959);
nand U4292 (N_4292,N_3959,N_3612);
nand U4293 (N_4293,N_3573,N_3686);
and U4294 (N_4294,N_3517,N_3891);
nor U4295 (N_4295,N_3504,N_3675);
xor U4296 (N_4296,N_3569,N_3930);
xnor U4297 (N_4297,N_3911,N_3764);
nor U4298 (N_4298,N_3801,N_3741);
nand U4299 (N_4299,N_3957,N_3803);
xor U4300 (N_4300,N_3501,N_3720);
nand U4301 (N_4301,N_3684,N_3872);
nor U4302 (N_4302,N_3813,N_3517);
nor U4303 (N_4303,N_3682,N_3860);
nor U4304 (N_4304,N_3681,N_3766);
nand U4305 (N_4305,N_3722,N_3959);
or U4306 (N_4306,N_3953,N_3553);
or U4307 (N_4307,N_3535,N_3695);
or U4308 (N_4308,N_3999,N_3900);
nand U4309 (N_4309,N_3809,N_3548);
nor U4310 (N_4310,N_3563,N_3917);
xor U4311 (N_4311,N_3512,N_3794);
xor U4312 (N_4312,N_3942,N_3824);
nand U4313 (N_4313,N_3810,N_3837);
nor U4314 (N_4314,N_3759,N_3810);
xor U4315 (N_4315,N_3790,N_3919);
xnor U4316 (N_4316,N_3904,N_3999);
or U4317 (N_4317,N_3565,N_3888);
and U4318 (N_4318,N_3684,N_3532);
xnor U4319 (N_4319,N_3600,N_3841);
nor U4320 (N_4320,N_3642,N_3661);
nor U4321 (N_4321,N_3708,N_3865);
and U4322 (N_4322,N_3929,N_3977);
xor U4323 (N_4323,N_3541,N_3951);
nor U4324 (N_4324,N_3925,N_3533);
xnor U4325 (N_4325,N_3576,N_3936);
xor U4326 (N_4326,N_3965,N_3810);
xnor U4327 (N_4327,N_3657,N_3769);
xnor U4328 (N_4328,N_3755,N_3655);
nand U4329 (N_4329,N_3577,N_3932);
or U4330 (N_4330,N_3615,N_3671);
nor U4331 (N_4331,N_3595,N_3535);
or U4332 (N_4332,N_3581,N_3928);
nand U4333 (N_4333,N_3731,N_3862);
nor U4334 (N_4334,N_3785,N_3836);
nand U4335 (N_4335,N_3594,N_3945);
xor U4336 (N_4336,N_3897,N_3942);
or U4337 (N_4337,N_3809,N_3998);
nor U4338 (N_4338,N_3660,N_3980);
or U4339 (N_4339,N_3636,N_3919);
nor U4340 (N_4340,N_3553,N_3741);
xnor U4341 (N_4341,N_3540,N_3744);
or U4342 (N_4342,N_3508,N_3542);
and U4343 (N_4343,N_3817,N_3955);
nand U4344 (N_4344,N_3619,N_3673);
nand U4345 (N_4345,N_3979,N_3778);
nor U4346 (N_4346,N_3703,N_3873);
or U4347 (N_4347,N_3980,N_3768);
xnor U4348 (N_4348,N_3985,N_3561);
or U4349 (N_4349,N_3585,N_3632);
and U4350 (N_4350,N_3765,N_3524);
and U4351 (N_4351,N_3520,N_3967);
nor U4352 (N_4352,N_3644,N_3895);
and U4353 (N_4353,N_3944,N_3941);
nor U4354 (N_4354,N_3906,N_3646);
nor U4355 (N_4355,N_3566,N_3856);
xor U4356 (N_4356,N_3714,N_3550);
xor U4357 (N_4357,N_3857,N_3891);
and U4358 (N_4358,N_3965,N_3982);
and U4359 (N_4359,N_3695,N_3784);
nor U4360 (N_4360,N_3549,N_3765);
nor U4361 (N_4361,N_3724,N_3664);
or U4362 (N_4362,N_3656,N_3578);
and U4363 (N_4363,N_3873,N_3775);
and U4364 (N_4364,N_3540,N_3587);
and U4365 (N_4365,N_3671,N_3582);
xor U4366 (N_4366,N_3993,N_3672);
xor U4367 (N_4367,N_3783,N_3879);
xnor U4368 (N_4368,N_3963,N_3975);
nand U4369 (N_4369,N_3605,N_3773);
nand U4370 (N_4370,N_3600,N_3886);
and U4371 (N_4371,N_3678,N_3886);
nor U4372 (N_4372,N_3639,N_3704);
nand U4373 (N_4373,N_3553,N_3542);
xor U4374 (N_4374,N_3683,N_3823);
nor U4375 (N_4375,N_3793,N_3985);
or U4376 (N_4376,N_3999,N_3883);
xnor U4377 (N_4377,N_3938,N_3764);
xor U4378 (N_4378,N_3722,N_3895);
or U4379 (N_4379,N_3561,N_3622);
nor U4380 (N_4380,N_3682,N_3824);
nand U4381 (N_4381,N_3814,N_3747);
nor U4382 (N_4382,N_3908,N_3918);
nor U4383 (N_4383,N_3935,N_3919);
and U4384 (N_4384,N_3721,N_3668);
or U4385 (N_4385,N_3592,N_3684);
nor U4386 (N_4386,N_3703,N_3689);
nand U4387 (N_4387,N_3539,N_3696);
or U4388 (N_4388,N_3974,N_3584);
xnor U4389 (N_4389,N_3924,N_3739);
or U4390 (N_4390,N_3694,N_3831);
or U4391 (N_4391,N_3514,N_3659);
nand U4392 (N_4392,N_3791,N_3867);
or U4393 (N_4393,N_3635,N_3610);
nor U4394 (N_4394,N_3901,N_3736);
nor U4395 (N_4395,N_3767,N_3960);
or U4396 (N_4396,N_3835,N_3674);
or U4397 (N_4397,N_3818,N_3517);
nor U4398 (N_4398,N_3702,N_3628);
nand U4399 (N_4399,N_3560,N_3648);
xor U4400 (N_4400,N_3749,N_3775);
and U4401 (N_4401,N_3864,N_3632);
or U4402 (N_4402,N_3977,N_3659);
and U4403 (N_4403,N_3779,N_3676);
and U4404 (N_4404,N_3566,N_3851);
nand U4405 (N_4405,N_3784,N_3993);
nand U4406 (N_4406,N_3813,N_3611);
or U4407 (N_4407,N_3754,N_3777);
nand U4408 (N_4408,N_3698,N_3535);
nand U4409 (N_4409,N_3883,N_3519);
nor U4410 (N_4410,N_3647,N_3511);
or U4411 (N_4411,N_3608,N_3943);
and U4412 (N_4412,N_3610,N_3942);
and U4413 (N_4413,N_3558,N_3688);
nand U4414 (N_4414,N_3941,N_3759);
or U4415 (N_4415,N_3557,N_3825);
and U4416 (N_4416,N_3712,N_3800);
nand U4417 (N_4417,N_3500,N_3837);
nand U4418 (N_4418,N_3623,N_3687);
nor U4419 (N_4419,N_3662,N_3752);
nor U4420 (N_4420,N_3664,N_3659);
or U4421 (N_4421,N_3570,N_3671);
and U4422 (N_4422,N_3997,N_3979);
xor U4423 (N_4423,N_3501,N_3760);
nand U4424 (N_4424,N_3638,N_3513);
or U4425 (N_4425,N_3845,N_3584);
nor U4426 (N_4426,N_3800,N_3746);
nor U4427 (N_4427,N_3819,N_3601);
nand U4428 (N_4428,N_3816,N_3779);
xor U4429 (N_4429,N_3759,N_3790);
nand U4430 (N_4430,N_3562,N_3761);
xor U4431 (N_4431,N_3534,N_3817);
or U4432 (N_4432,N_3852,N_3627);
or U4433 (N_4433,N_3575,N_3644);
nor U4434 (N_4434,N_3678,N_3781);
and U4435 (N_4435,N_3513,N_3916);
nand U4436 (N_4436,N_3627,N_3725);
or U4437 (N_4437,N_3804,N_3916);
xnor U4438 (N_4438,N_3582,N_3870);
nand U4439 (N_4439,N_3787,N_3659);
nand U4440 (N_4440,N_3634,N_3512);
and U4441 (N_4441,N_3755,N_3725);
nor U4442 (N_4442,N_3974,N_3778);
nand U4443 (N_4443,N_3636,N_3650);
or U4444 (N_4444,N_3699,N_3796);
or U4445 (N_4445,N_3615,N_3685);
nand U4446 (N_4446,N_3671,N_3982);
and U4447 (N_4447,N_3860,N_3533);
nand U4448 (N_4448,N_3857,N_3552);
or U4449 (N_4449,N_3741,N_3938);
nand U4450 (N_4450,N_3971,N_3700);
nor U4451 (N_4451,N_3989,N_3769);
and U4452 (N_4452,N_3536,N_3878);
nand U4453 (N_4453,N_3516,N_3889);
and U4454 (N_4454,N_3737,N_3724);
or U4455 (N_4455,N_3674,N_3632);
and U4456 (N_4456,N_3564,N_3980);
and U4457 (N_4457,N_3527,N_3651);
xor U4458 (N_4458,N_3866,N_3977);
and U4459 (N_4459,N_3590,N_3895);
and U4460 (N_4460,N_3853,N_3860);
or U4461 (N_4461,N_3636,N_3996);
or U4462 (N_4462,N_3526,N_3525);
or U4463 (N_4463,N_3670,N_3986);
or U4464 (N_4464,N_3879,N_3997);
xor U4465 (N_4465,N_3648,N_3685);
xor U4466 (N_4466,N_3997,N_3500);
or U4467 (N_4467,N_3918,N_3698);
and U4468 (N_4468,N_3573,N_3720);
or U4469 (N_4469,N_3598,N_3979);
and U4470 (N_4470,N_3940,N_3834);
xnor U4471 (N_4471,N_3508,N_3697);
or U4472 (N_4472,N_3689,N_3933);
nand U4473 (N_4473,N_3863,N_3989);
or U4474 (N_4474,N_3936,N_3729);
nor U4475 (N_4475,N_3777,N_3942);
nand U4476 (N_4476,N_3803,N_3819);
nor U4477 (N_4477,N_3745,N_3510);
or U4478 (N_4478,N_3841,N_3606);
nand U4479 (N_4479,N_3937,N_3668);
xor U4480 (N_4480,N_3989,N_3831);
nand U4481 (N_4481,N_3957,N_3708);
or U4482 (N_4482,N_3979,N_3935);
or U4483 (N_4483,N_3534,N_3830);
nand U4484 (N_4484,N_3931,N_3981);
nor U4485 (N_4485,N_3736,N_3535);
nand U4486 (N_4486,N_3784,N_3655);
or U4487 (N_4487,N_3596,N_3762);
xnor U4488 (N_4488,N_3568,N_3761);
nand U4489 (N_4489,N_3706,N_3944);
xnor U4490 (N_4490,N_3961,N_3936);
nor U4491 (N_4491,N_3757,N_3586);
xnor U4492 (N_4492,N_3748,N_3849);
and U4493 (N_4493,N_3786,N_3730);
nor U4494 (N_4494,N_3746,N_3581);
or U4495 (N_4495,N_3798,N_3624);
xnor U4496 (N_4496,N_3527,N_3948);
or U4497 (N_4497,N_3615,N_3959);
nand U4498 (N_4498,N_3569,N_3552);
xnor U4499 (N_4499,N_3897,N_3874);
nor U4500 (N_4500,N_4003,N_4266);
and U4501 (N_4501,N_4120,N_4194);
nor U4502 (N_4502,N_4082,N_4118);
and U4503 (N_4503,N_4161,N_4019);
and U4504 (N_4504,N_4395,N_4045);
nor U4505 (N_4505,N_4034,N_4234);
nand U4506 (N_4506,N_4157,N_4098);
and U4507 (N_4507,N_4095,N_4466);
xor U4508 (N_4508,N_4491,N_4424);
xnor U4509 (N_4509,N_4027,N_4015);
nand U4510 (N_4510,N_4293,N_4298);
xnor U4511 (N_4511,N_4277,N_4427);
or U4512 (N_4512,N_4192,N_4428);
nor U4513 (N_4513,N_4220,N_4342);
xor U4514 (N_4514,N_4049,N_4106);
and U4515 (N_4515,N_4265,N_4474);
and U4516 (N_4516,N_4290,N_4442);
nor U4517 (N_4517,N_4473,N_4047);
or U4518 (N_4518,N_4068,N_4496);
nand U4519 (N_4519,N_4207,N_4330);
xnor U4520 (N_4520,N_4413,N_4262);
nor U4521 (N_4521,N_4248,N_4339);
nor U4522 (N_4522,N_4079,N_4141);
nand U4523 (N_4523,N_4421,N_4305);
and U4524 (N_4524,N_4255,N_4356);
xor U4525 (N_4525,N_4004,N_4477);
or U4526 (N_4526,N_4406,N_4016);
xnor U4527 (N_4527,N_4012,N_4401);
nand U4528 (N_4528,N_4455,N_4479);
or U4529 (N_4529,N_4076,N_4494);
nor U4530 (N_4530,N_4060,N_4375);
or U4531 (N_4531,N_4493,N_4077);
nand U4532 (N_4532,N_4202,N_4002);
nor U4533 (N_4533,N_4402,N_4454);
or U4534 (N_4534,N_4272,N_4052);
xnor U4535 (N_4535,N_4259,N_4389);
nand U4536 (N_4536,N_4008,N_4124);
nand U4537 (N_4537,N_4149,N_4351);
and U4538 (N_4538,N_4179,N_4196);
nand U4539 (N_4539,N_4245,N_4303);
xor U4540 (N_4540,N_4000,N_4185);
xnor U4541 (N_4541,N_4144,N_4097);
nand U4542 (N_4542,N_4445,N_4468);
or U4543 (N_4543,N_4464,N_4386);
nor U4544 (N_4544,N_4116,N_4180);
nand U4545 (N_4545,N_4282,N_4319);
and U4546 (N_4546,N_4136,N_4490);
xor U4547 (N_4547,N_4289,N_4457);
and U4548 (N_4548,N_4054,N_4066);
and U4549 (N_4549,N_4200,N_4013);
and U4550 (N_4550,N_4417,N_4204);
nand U4551 (N_4551,N_4415,N_4126);
and U4552 (N_4552,N_4101,N_4155);
nand U4553 (N_4553,N_4397,N_4295);
or U4554 (N_4554,N_4093,N_4300);
or U4555 (N_4555,N_4405,N_4297);
or U4556 (N_4556,N_4354,N_4355);
and U4557 (N_4557,N_4193,N_4286);
xor U4558 (N_4558,N_4326,N_4203);
xnor U4559 (N_4559,N_4432,N_4214);
and U4560 (N_4560,N_4311,N_4434);
nor U4561 (N_4561,N_4344,N_4288);
and U4562 (N_4562,N_4377,N_4380);
and U4563 (N_4563,N_4212,N_4195);
nor U4564 (N_4564,N_4021,N_4143);
nand U4565 (N_4565,N_4362,N_4190);
nand U4566 (N_4566,N_4050,N_4310);
xor U4567 (N_4567,N_4152,N_4170);
nor U4568 (N_4568,N_4285,N_4062);
nor U4569 (N_4569,N_4256,N_4283);
nor U4570 (N_4570,N_4430,N_4167);
and U4571 (N_4571,N_4217,N_4410);
or U4572 (N_4572,N_4264,N_4487);
or U4573 (N_4573,N_4110,N_4073);
nor U4574 (N_4574,N_4274,N_4348);
xnor U4575 (N_4575,N_4041,N_4221);
xnor U4576 (N_4576,N_4233,N_4419);
and U4577 (N_4577,N_4053,N_4105);
nor U4578 (N_4578,N_4206,N_4373);
or U4579 (N_4579,N_4132,N_4125);
nand U4580 (N_4580,N_4215,N_4044);
or U4581 (N_4581,N_4462,N_4173);
or U4582 (N_4582,N_4061,N_4369);
and U4583 (N_4583,N_4183,N_4322);
xor U4584 (N_4584,N_4001,N_4372);
nand U4585 (N_4585,N_4017,N_4357);
nor U4586 (N_4586,N_4318,N_4018);
and U4587 (N_4587,N_4114,N_4365);
nor U4588 (N_4588,N_4481,N_4460);
nor U4589 (N_4589,N_4242,N_4439);
and U4590 (N_4590,N_4036,N_4112);
nor U4591 (N_4591,N_4270,N_4005);
xnor U4592 (N_4592,N_4287,N_4168);
or U4593 (N_4593,N_4399,N_4440);
nand U4594 (N_4594,N_4317,N_4361);
and U4595 (N_4595,N_4228,N_4391);
and U4596 (N_4596,N_4497,N_4441);
or U4597 (N_4597,N_4463,N_4321);
or U4598 (N_4598,N_4250,N_4184);
nand U4599 (N_4599,N_4086,N_4331);
or U4600 (N_4600,N_4191,N_4235);
or U4601 (N_4601,N_4307,N_4396);
or U4602 (N_4602,N_4129,N_4345);
or U4603 (N_4603,N_4387,N_4394);
nor U4604 (N_4604,N_4058,N_4324);
nor U4605 (N_4605,N_4178,N_4325);
and U4606 (N_4606,N_4131,N_4418);
nor U4607 (N_4607,N_4032,N_4480);
nor U4608 (N_4608,N_4343,N_4230);
or U4609 (N_4609,N_4227,N_4056);
nand U4610 (N_4610,N_4469,N_4431);
nor U4611 (N_4611,N_4216,N_4156);
or U4612 (N_4612,N_4094,N_4301);
and U4613 (N_4613,N_4336,N_4091);
nor U4614 (N_4614,N_4411,N_4291);
nor U4615 (N_4615,N_4360,N_4188);
xor U4616 (N_4616,N_4224,N_4231);
xor U4617 (N_4617,N_4029,N_4009);
xor U4618 (N_4618,N_4145,N_4099);
and U4619 (N_4619,N_4456,N_4089);
or U4620 (N_4620,N_4461,N_4241);
nand U4621 (N_4621,N_4452,N_4181);
and U4622 (N_4622,N_4448,N_4346);
and U4623 (N_4623,N_4218,N_4476);
or U4624 (N_4624,N_4407,N_4025);
nand U4625 (N_4625,N_4294,N_4085);
nor U4626 (N_4626,N_4171,N_4363);
xnor U4627 (N_4627,N_4254,N_4040);
nor U4628 (N_4628,N_4371,N_4223);
nor U4629 (N_4629,N_4172,N_4482);
xor U4630 (N_4630,N_4103,N_4446);
and U4631 (N_4631,N_4467,N_4420);
nor U4632 (N_4632,N_4258,N_4051);
nor U4633 (N_4633,N_4280,N_4299);
or U4634 (N_4634,N_4088,N_4022);
nor U4635 (N_4635,N_4253,N_4353);
nor U4636 (N_4636,N_4121,N_4334);
or U4637 (N_4637,N_4292,N_4281);
nor U4638 (N_4638,N_4064,N_4388);
xnor U4639 (N_4639,N_4252,N_4123);
and U4640 (N_4640,N_4384,N_4475);
or U4641 (N_4641,N_4160,N_4453);
nor U4642 (N_4642,N_4147,N_4139);
nand U4643 (N_4643,N_4057,N_4451);
nor U4644 (N_4644,N_4409,N_4247);
or U4645 (N_4645,N_4083,N_4176);
xnor U4646 (N_4646,N_4390,N_4080);
nand U4647 (N_4647,N_4037,N_4059);
or U4648 (N_4648,N_4308,N_4314);
nand U4649 (N_4649,N_4425,N_4043);
xor U4650 (N_4650,N_4166,N_4028);
or U4651 (N_4651,N_4304,N_4443);
nand U4652 (N_4652,N_4031,N_4133);
nand U4653 (N_4653,N_4219,N_4198);
or U4654 (N_4654,N_4358,N_4393);
or U4655 (N_4655,N_4329,N_4039);
nand U4656 (N_4656,N_4333,N_4006);
nand U4657 (N_4657,N_4100,N_4422);
and U4658 (N_4658,N_4302,N_4492);
or U4659 (N_4659,N_4150,N_4134);
and U4660 (N_4660,N_4400,N_4007);
or U4661 (N_4661,N_4213,N_4385);
nor U4662 (N_4662,N_4140,N_4119);
or U4663 (N_4663,N_4090,N_4251);
nor U4664 (N_4664,N_4197,N_4323);
xnor U4665 (N_4665,N_4163,N_4164);
nand U4666 (N_4666,N_4312,N_4412);
or U4667 (N_4667,N_4313,N_4332);
or U4668 (N_4668,N_4158,N_4024);
nor U4669 (N_4669,N_4162,N_4175);
xor U4670 (N_4670,N_4065,N_4340);
nand U4671 (N_4671,N_4260,N_4046);
xnor U4672 (N_4672,N_4499,N_4261);
and U4673 (N_4673,N_4284,N_4146);
and U4674 (N_4674,N_4426,N_4240);
xor U4675 (N_4675,N_4199,N_4137);
nor U4676 (N_4676,N_4279,N_4465);
xor U4677 (N_4677,N_4169,N_4392);
or U4678 (N_4678,N_4023,N_4069);
xnor U4679 (N_4679,N_4084,N_4296);
nand U4680 (N_4680,N_4483,N_4403);
or U4681 (N_4681,N_4488,N_4055);
nor U4682 (N_4682,N_4135,N_4078);
or U4683 (N_4683,N_4225,N_4239);
and U4684 (N_4684,N_4267,N_4379);
and U4685 (N_4685,N_4165,N_4485);
nor U4686 (N_4686,N_4376,N_4367);
xor U4687 (N_4687,N_4316,N_4368);
xnor U4688 (N_4688,N_4115,N_4438);
xnor U4689 (N_4689,N_4489,N_4142);
nand U4690 (N_4690,N_4208,N_4472);
nor U4691 (N_4691,N_4177,N_4229);
nand U4692 (N_4692,N_4370,N_4237);
nor U4693 (N_4693,N_4201,N_4130);
nor U4694 (N_4694,N_4416,N_4246);
nor U4695 (N_4695,N_4398,N_4102);
xnor U4696 (N_4696,N_4092,N_4238);
nand U4697 (N_4697,N_4347,N_4249);
nand U4698 (N_4698,N_4081,N_4471);
or U4699 (N_4699,N_4182,N_4075);
nor U4700 (N_4700,N_4341,N_4486);
or U4701 (N_4701,N_4128,N_4484);
or U4702 (N_4702,N_4435,N_4122);
or U4703 (N_4703,N_4010,N_4359);
or U4704 (N_4704,N_4063,N_4408);
nand U4705 (N_4705,N_4459,N_4148);
xnor U4706 (N_4706,N_4209,N_4433);
xor U4707 (N_4707,N_4072,N_4127);
and U4708 (N_4708,N_4278,N_4187);
or U4709 (N_4709,N_4153,N_4074);
nand U4710 (N_4710,N_4275,N_4374);
nand U4711 (N_4711,N_4269,N_4273);
or U4712 (N_4712,N_4035,N_4033);
and U4713 (N_4713,N_4449,N_4236);
nor U4714 (N_4714,N_4349,N_4154);
xnor U4715 (N_4715,N_4107,N_4096);
or U4716 (N_4716,N_4450,N_4328);
xor U4717 (N_4717,N_4186,N_4067);
and U4718 (N_4718,N_4268,N_4383);
and U4719 (N_4719,N_4271,N_4087);
or U4720 (N_4720,N_4495,N_4352);
nand U4721 (N_4721,N_4404,N_4210);
and U4722 (N_4722,N_4138,N_4211);
nand U4723 (N_4723,N_4470,N_4014);
or U4724 (N_4724,N_4243,N_4020);
nor U4725 (N_4725,N_4070,N_4335);
xnor U4726 (N_4726,N_4315,N_4030);
and U4727 (N_4727,N_4263,N_4026);
or U4728 (N_4728,N_4042,N_4117);
nor U4729 (N_4729,N_4382,N_4222);
and U4730 (N_4730,N_4109,N_4437);
xnor U4731 (N_4731,N_4444,N_4381);
xor U4732 (N_4732,N_4159,N_4108);
nor U4733 (N_4733,N_4320,N_4306);
nor U4734 (N_4734,N_4337,N_4423);
or U4735 (N_4735,N_4048,N_4071);
and U4736 (N_4736,N_4232,N_4338);
and U4737 (N_4737,N_4309,N_4447);
xnor U4738 (N_4738,N_4257,N_4104);
or U4739 (N_4739,N_4478,N_4276);
nand U4740 (N_4740,N_4327,N_4111);
nor U4741 (N_4741,N_4244,N_4226);
or U4742 (N_4742,N_4189,N_4366);
nor U4743 (N_4743,N_4151,N_4113);
nor U4744 (N_4744,N_4498,N_4350);
and U4745 (N_4745,N_4174,N_4458);
nor U4746 (N_4746,N_4364,N_4436);
and U4747 (N_4747,N_4429,N_4011);
nor U4748 (N_4748,N_4378,N_4205);
nand U4749 (N_4749,N_4414,N_4038);
and U4750 (N_4750,N_4466,N_4433);
xor U4751 (N_4751,N_4309,N_4381);
and U4752 (N_4752,N_4247,N_4008);
or U4753 (N_4753,N_4040,N_4025);
and U4754 (N_4754,N_4170,N_4362);
or U4755 (N_4755,N_4225,N_4397);
xnor U4756 (N_4756,N_4124,N_4386);
nor U4757 (N_4757,N_4237,N_4234);
nand U4758 (N_4758,N_4077,N_4015);
and U4759 (N_4759,N_4181,N_4361);
nor U4760 (N_4760,N_4324,N_4152);
and U4761 (N_4761,N_4315,N_4345);
nand U4762 (N_4762,N_4183,N_4068);
or U4763 (N_4763,N_4173,N_4368);
nor U4764 (N_4764,N_4174,N_4027);
or U4765 (N_4765,N_4373,N_4232);
nor U4766 (N_4766,N_4440,N_4010);
or U4767 (N_4767,N_4482,N_4292);
nand U4768 (N_4768,N_4340,N_4313);
or U4769 (N_4769,N_4446,N_4285);
xor U4770 (N_4770,N_4455,N_4400);
or U4771 (N_4771,N_4203,N_4139);
and U4772 (N_4772,N_4039,N_4110);
and U4773 (N_4773,N_4026,N_4462);
nor U4774 (N_4774,N_4058,N_4036);
and U4775 (N_4775,N_4243,N_4412);
or U4776 (N_4776,N_4007,N_4021);
xor U4777 (N_4777,N_4239,N_4221);
and U4778 (N_4778,N_4456,N_4331);
xnor U4779 (N_4779,N_4099,N_4483);
xor U4780 (N_4780,N_4003,N_4075);
and U4781 (N_4781,N_4459,N_4129);
xor U4782 (N_4782,N_4034,N_4193);
xnor U4783 (N_4783,N_4082,N_4085);
and U4784 (N_4784,N_4371,N_4267);
or U4785 (N_4785,N_4395,N_4000);
or U4786 (N_4786,N_4089,N_4399);
and U4787 (N_4787,N_4031,N_4264);
nand U4788 (N_4788,N_4497,N_4475);
and U4789 (N_4789,N_4333,N_4419);
nand U4790 (N_4790,N_4281,N_4302);
nand U4791 (N_4791,N_4365,N_4235);
or U4792 (N_4792,N_4048,N_4407);
xor U4793 (N_4793,N_4407,N_4176);
and U4794 (N_4794,N_4215,N_4018);
xnor U4795 (N_4795,N_4086,N_4443);
nand U4796 (N_4796,N_4162,N_4443);
nor U4797 (N_4797,N_4437,N_4369);
and U4798 (N_4798,N_4004,N_4483);
nor U4799 (N_4799,N_4299,N_4424);
xnor U4800 (N_4800,N_4077,N_4111);
and U4801 (N_4801,N_4216,N_4031);
xnor U4802 (N_4802,N_4253,N_4360);
xnor U4803 (N_4803,N_4170,N_4261);
and U4804 (N_4804,N_4031,N_4293);
xnor U4805 (N_4805,N_4386,N_4390);
nor U4806 (N_4806,N_4424,N_4451);
or U4807 (N_4807,N_4360,N_4244);
and U4808 (N_4808,N_4281,N_4385);
xnor U4809 (N_4809,N_4339,N_4478);
xnor U4810 (N_4810,N_4004,N_4429);
and U4811 (N_4811,N_4455,N_4062);
nand U4812 (N_4812,N_4274,N_4091);
nor U4813 (N_4813,N_4399,N_4290);
or U4814 (N_4814,N_4247,N_4328);
xor U4815 (N_4815,N_4172,N_4428);
nor U4816 (N_4816,N_4406,N_4071);
nor U4817 (N_4817,N_4187,N_4452);
and U4818 (N_4818,N_4338,N_4310);
nand U4819 (N_4819,N_4201,N_4023);
nand U4820 (N_4820,N_4496,N_4268);
and U4821 (N_4821,N_4177,N_4463);
nor U4822 (N_4822,N_4097,N_4273);
nand U4823 (N_4823,N_4395,N_4288);
and U4824 (N_4824,N_4380,N_4102);
and U4825 (N_4825,N_4198,N_4494);
and U4826 (N_4826,N_4280,N_4088);
and U4827 (N_4827,N_4076,N_4301);
nor U4828 (N_4828,N_4490,N_4450);
xnor U4829 (N_4829,N_4207,N_4383);
xor U4830 (N_4830,N_4353,N_4102);
xor U4831 (N_4831,N_4466,N_4488);
xor U4832 (N_4832,N_4329,N_4051);
and U4833 (N_4833,N_4204,N_4157);
xnor U4834 (N_4834,N_4207,N_4306);
nand U4835 (N_4835,N_4393,N_4491);
xor U4836 (N_4836,N_4301,N_4199);
nor U4837 (N_4837,N_4329,N_4014);
xor U4838 (N_4838,N_4429,N_4102);
nand U4839 (N_4839,N_4209,N_4158);
xor U4840 (N_4840,N_4389,N_4452);
nor U4841 (N_4841,N_4388,N_4175);
or U4842 (N_4842,N_4455,N_4299);
nor U4843 (N_4843,N_4063,N_4002);
nor U4844 (N_4844,N_4326,N_4050);
nor U4845 (N_4845,N_4062,N_4057);
or U4846 (N_4846,N_4037,N_4139);
and U4847 (N_4847,N_4163,N_4187);
nor U4848 (N_4848,N_4140,N_4099);
or U4849 (N_4849,N_4132,N_4358);
and U4850 (N_4850,N_4202,N_4182);
xor U4851 (N_4851,N_4412,N_4493);
xor U4852 (N_4852,N_4388,N_4247);
xnor U4853 (N_4853,N_4452,N_4026);
or U4854 (N_4854,N_4081,N_4493);
nand U4855 (N_4855,N_4052,N_4488);
xor U4856 (N_4856,N_4324,N_4345);
or U4857 (N_4857,N_4382,N_4349);
xor U4858 (N_4858,N_4463,N_4053);
nor U4859 (N_4859,N_4277,N_4044);
or U4860 (N_4860,N_4364,N_4154);
xor U4861 (N_4861,N_4076,N_4118);
and U4862 (N_4862,N_4305,N_4163);
or U4863 (N_4863,N_4241,N_4117);
and U4864 (N_4864,N_4212,N_4364);
nand U4865 (N_4865,N_4194,N_4476);
or U4866 (N_4866,N_4057,N_4178);
nand U4867 (N_4867,N_4088,N_4219);
and U4868 (N_4868,N_4183,N_4007);
nor U4869 (N_4869,N_4161,N_4222);
or U4870 (N_4870,N_4030,N_4036);
nand U4871 (N_4871,N_4081,N_4468);
or U4872 (N_4872,N_4162,N_4167);
xnor U4873 (N_4873,N_4374,N_4000);
nand U4874 (N_4874,N_4110,N_4380);
nand U4875 (N_4875,N_4018,N_4433);
xor U4876 (N_4876,N_4024,N_4110);
xnor U4877 (N_4877,N_4413,N_4234);
or U4878 (N_4878,N_4074,N_4353);
or U4879 (N_4879,N_4311,N_4485);
and U4880 (N_4880,N_4393,N_4202);
or U4881 (N_4881,N_4291,N_4028);
and U4882 (N_4882,N_4313,N_4234);
nand U4883 (N_4883,N_4409,N_4318);
xor U4884 (N_4884,N_4014,N_4412);
or U4885 (N_4885,N_4461,N_4148);
nor U4886 (N_4886,N_4319,N_4314);
xor U4887 (N_4887,N_4282,N_4216);
or U4888 (N_4888,N_4169,N_4040);
nor U4889 (N_4889,N_4046,N_4206);
and U4890 (N_4890,N_4473,N_4376);
nand U4891 (N_4891,N_4266,N_4151);
nand U4892 (N_4892,N_4261,N_4216);
nand U4893 (N_4893,N_4279,N_4216);
nor U4894 (N_4894,N_4171,N_4217);
and U4895 (N_4895,N_4283,N_4042);
nand U4896 (N_4896,N_4242,N_4156);
nor U4897 (N_4897,N_4322,N_4129);
and U4898 (N_4898,N_4271,N_4413);
and U4899 (N_4899,N_4251,N_4379);
and U4900 (N_4900,N_4436,N_4043);
and U4901 (N_4901,N_4149,N_4203);
nor U4902 (N_4902,N_4496,N_4291);
nand U4903 (N_4903,N_4060,N_4247);
and U4904 (N_4904,N_4458,N_4366);
nand U4905 (N_4905,N_4250,N_4350);
xnor U4906 (N_4906,N_4031,N_4278);
nor U4907 (N_4907,N_4120,N_4052);
nand U4908 (N_4908,N_4052,N_4357);
nor U4909 (N_4909,N_4426,N_4191);
nand U4910 (N_4910,N_4465,N_4294);
and U4911 (N_4911,N_4160,N_4310);
xnor U4912 (N_4912,N_4305,N_4228);
or U4913 (N_4913,N_4158,N_4493);
xor U4914 (N_4914,N_4176,N_4317);
and U4915 (N_4915,N_4462,N_4070);
xor U4916 (N_4916,N_4212,N_4430);
nand U4917 (N_4917,N_4416,N_4209);
and U4918 (N_4918,N_4133,N_4310);
nand U4919 (N_4919,N_4266,N_4411);
xnor U4920 (N_4920,N_4269,N_4208);
and U4921 (N_4921,N_4408,N_4242);
nor U4922 (N_4922,N_4484,N_4478);
or U4923 (N_4923,N_4448,N_4181);
or U4924 (N_4924,N_4228,N_4426);
xor U4925 (N_4925,N_4022,N_4344);
nor U4926 (N_4926,N_4218,N_4487);
nand U4927 (N_4927,N_4310,N_4485);
xor U4928 (N_4928,N_4206,N_4461);
and U4929 (N_4929,N_4375,N_4360);
nand U4930 (N_4930,N_4203,N_4338);
or U4931 (N_4931,N_4442,N_4063);
nor U4932 (N_4932,N_4086,N_4159);
or U4933 (N_4933,N_4431,N_4405);
or U4934 (N_4934,N_4121,N_4275);
or U4935 (N_4935,N_4478,N_4050);
nor U4936 (N_4936,N_4349,N_4310);
nand U4937 (N_4937,N_4345,N_4260);
and U4938 (N_4938,N_4103,N_4094);
and U4939 (N_4939,N_4456,N_4497);
xnor U4940 (N_4940,N_4222,N_4002);
nor U4941 (N_4941,N_4010,N_4239);
nand U4942 (N_4942,N_4050,N_4244);
and U4943 (N_4943,N_4459,N_4133);
and U4944 (N_4944,N_4274,N_4231);
and U4945 (N_4945,N_4330,N_4339);
xor U4946 (N_4946,N_4170,N_4063);
nand U4947 (N_4947,N_4309,N_4431);
nand U4948 (N_4948,N_4419,N_4261);
nand U4949 (N_4949,N_4277,N_4280);
or U4950 (N_4950,N_4099,N_4176);
nand U4951 (N_4951,N_4343,N_4147);
or U4952 (N_4952,N_4379,N_4390);
xor U4953 (N_4953,N_4167,N_4440);
nor U4954 (N_4954,N_4148,N_4110);
nand U4955 (N_4955,N_4026,N_4253);
nand U4956 (N_4956,N_4108,N_4263);
or U4957 (N_4957,N_4023,N_4006);
xnor U4958 (N_4958,N_4191,N_4128);
nand U4959 (N_4959,N_4376,N_4180);
and U4960 (N_4960,N_4166,N_4470);
or U4961 (N_4961,N_4321,N_4047);
or U4962 (N_4962,N_4219,N_4007);
xnor U4963 (N_4963,N_4076,N_4110);
xor U4964 (N_4964,N_4045,N_4219);
or U4965 (N_4965,N_4085,N_4408);
or U4966 (N_4966,N_4025,N_4084);
nand U4967 (N_4967,N_4270,N_4464);
and U4968 (N_4968,N_4390,N_4040);
or U4969 (N_4969,N_4427,N_4161);
and U4970 (N_4970,N_4053,N_4298);
nor U4971 (N_4971,N_4102,N_4215);
xnor U4972 (N_4972,N_4040,N_4214);
xor U4973 (N_4973,N_4324,N_4133);
nor U4974 (N_4974,N_4048,N_4164);
nand U4975 (N_4975,N_4166,N_4095);
xnor U4976 (N_4976,N_4204,N_4385);
and U4977 (N_4977,N_4111,N_4123);
or U4978 (N_4978,N_4216,N_4440);
and U4979 (N_4979,N_4121,N_4356);
or U4980 (N_4980,N_4083,N_4339);
nor U4981 (N_4981,N_4315,N_4314);
or U4982 (N_4982,N_4033,N_4183);
and U4983 (N_4983,N_4237,N_4168);
and U4984 (N_4984,N_4089,N_4194);
xor U4985 (N_4985,N_4110,N_4302);
xnor U4986 (N_4986,N_4348,N_4156);
nor U4987 (N_4987,N_4324,N_4061);
nor U4988 (N_4988,N_4375,N_4346);
or U4989 (N_4989,N_4360,N_4018);
nor U4990 (N_4990,N_4067,N_4248);
nor U4991 (N_4991,N_4101,N_4230);
or U4992 (N_4992,N_4264,N_4332);
or U4993 (N_4993,N_4148,N_4134);
nand U4994 (N_4994,N_4413,N_4086);
and U4995 (N_4995,N_4441,N_4324);
nand U4996 (N_4996,N_4280,N_4249);
nor U4997 (N_4997,N_4226,N_4240);
nand U4998 (N_4998,N_4130,N_4221);
or U4999 (N_4999,N_4156,N_4495);
and U5000 (N_5000,N_4532,N_4911);
nor U5001 (N_5001,N_4610,N_4642);
and U5002 (N_5002,N_4530,N_4677);
xnor U5003 (N_5003,N_4947,N_4929);
nor U5004 (N_5004,N_4556,N_4658);
or U5005 (N_5005,N_4617,N_4982);
nand U5006 (N_5006,N_4662,N_4942);
and U5007 (N_5007,N_4673,N_4900);
nor U5008 (N_5008,N_4652,N_4754);
or U5009 (N_5009,N_4503,N_4772);
nand U5010 (N_5010,N_4558,N_4576);
xnor U5011 (N_5011,N_4629,N_4748);
and U5012 (N_5012,N_4737,N_4913);
and U5013 (N_5013,N_4813,N_4605);
and U5014 (N_5014,N_4705,N_4870);
nand U5015 (N_5015,N_4998,N_4835);
xor U5016 (N_5016,N_4654,N_4946);
or U5017 (N_5017,N_4923,N_4537);
and U5018 (N_5018,N_4630,N_4839);
or U5019 (N_5019,N_4843,N_4612);
or U5020 (N_5020,N_4846,N_4964);
nor U5021 (N_5021,N_4564,N_4917);
nand U5022 (N_5022,N_4738,N_4620);
and U5023 (N_5023,N_4663,N_4882);
nand U5024 (N_5024,N_4587,N_4904);
nand U5025 (N_5025,N_4722,N_4824);
xnor U5026 (N_5026,N_4603,N_4586);
xnor U5027 (N_5027,N_4571,N_4906);
and U5028 (N_5028,N_4749,N_4959);
or U5029 (N_5029,N_4800,N_4762);
nor U5030 (N_5030,N_4809,N_4599);
nor U5031 (N_5031,N_4579,N_4999);
xnor U5032 (N_5032,N_4508,N_4514);
xor U5033 (N_5033,N_4893,N_4950);
xor U5034 (N_5034,N_4624,N_4667);
nand U5035 (N_5035,N_4968,N_4692);
and U5036 (N_5036,N_4957,N_4615);
or U5037 (N_5037,N_4821,N_4674);
and U5038 (N_5038,N_4940,N_4535);
and U5039 (N_5039,N_4918,N_4907);
nor U5040 (N_5040,N_4747,N_4768);
nor U5041 (N_5041,N_4962,N_4689);
nand U5042 (N_5042,N_4729,N_4596);
or U5043 (N_5043,N_4553,N_4626);
nor U5044 (N_5044,N_4854,N_4788);
nor U5045 (N_5045,N_4698,N_4715);
or U5046 (N_5046,N_4896,N_4789);
or U5047 (N_5047,N_4770,N_4636);
or U5048 (N_5048,N_4894,N_4986);
nor U5049 (N_5049,N_4803,N_4575);
nand U5050 (N_5050,N_4811,N_4802);
xnor U5051 (N_5051,N_4822,N_4855);
nor U5052 (N_5052,N_4613,N_4841);
xor U5053 (N_5053,N_4951,N_4621);
xor U5054 (N_5054,N_4625,N_4786);
or U5055 (N_5055,N_4996,N_4676);
nand U5056 (N_5056,N_4644,N_4509);
or U5057 (N_5057,N_4505,N_4672);
and U5058 (N_5058,N_4682,N_4944);
or U5059 (N_5059,N_4700,N_4860);
nand U5060 (N_5060,N_4543,N_4932);
xnor U5061 (N_5061,N_4874,N_4512);
or U5062 (N_5062,N_4561,N_4686);
or U5063 (N_5063,N_4892,N_4725);
nor U5064 (N_5064,N_4542,N_4830);
xnor U5065 (N_5065,N_4949,N_4752);
and U5066 (N_5066,N_4814,N_4775);
or U5067 (N_5067,N_4753,N_4647);
xnor U5068 (N_5068,N_4721,N_4719);
nand U5069 (N_5069,N_4602,N_4941);
xor U5070 (N_5070,N_4559,N_4836);
nand U5071 (N_5071,N_4521,N_4659);
and U5072 (N_5072,N_4718,N_4798);
or U5073 (N_5073,N_4759,N_4655);
xnor U5074 (N_5074,N_4536,N_4981);
nand U5075 (N_5075,N_4777,N_4970);
nor U5076 (N_5076,N_4792,N_4879);
xor U5077 (N_5077,N_4651,N_4867);
nand U5078 (N_5078,N_4693,N_4616);
and U5079 (N_5079,N_4908,N_4552);
or U5080 (N_5080,N_4538,N_4588);
and U5081 (N_5081,N_4591,N_4875);
xor U5082 (N_5082,N_4608,N_4948);
xor U5083 (N_5083,N_4799,N_4953);
nor U5084 (N_5084,N_4598,N_4847);
or U5085 (N_5085,N_4745,N_4891);
and U5086 (N_5086,N_4888,N_4601);
nand U5087 (N_5087,N_4842,N_4766);
or U5088 (N_5088,N_4975,N_4736);
xor U5089 (N_5089,N_4983,N_4580);
nor U5090 (N_5090,N_4781,N_4680);
nor U5091 (N_5091,N_4681,N_4808);
xnor U5092 (N_5092,N_4660,N_4816);
nor U5093 (N_5093,N_4704,N_4921);
nand U5094 (N_5094,N_4963,N_4726);
xnor U5095 (N_5095,N_4831,N_4887);
nor U5096 (N_5096,N_4628,N_4779);
nand U5097 (N_5097,N_4684,N_4611);
or U5098 (N_5098,N_4504,N_4746);
nand U5099 (N_5099,N_4534,N_4510);
and U5100 (N_5100,N_4773,N_4861);
and U5101 (N_5101,N_4614,N_4837);
nand U5102 (N_5102,N_4685,N_4989);
xor U5103 (N_5103,N_4910,N_4528);
nor U5104 (N_5104,N_4895,N_4890);
or U5105 (N_5105,N_4812,N_4639);
nor U5106 (N_5106,N_4820,N_4665);
or U5107 (N_5107,N_4774,N_4883);
and U5108 (N_5108,N_4834,N_4683);
nand U5109 (N_5109,N_4872,N_4661);
nand U5110 (N_5110,N_4703,N_4701);
xor U5111 (N_5111,N_4666,N_4540);
and U5112 (N_5112,N_4697,N_4934);
nand U5113 (N_5113,N_4584,N_4524);
nor U5114 (N_5114,N_4868,N_4741);
nor U5115 (N_5115,N_4618,N_4997);
xnor U5116 (N_5116,N_4866,N_4585);
nand U5117 (N_5117,N_4756,N_4589);
nand U5118 (N_5118,N_4991,N_4827);
and U5119 (N_5119,N_4702,N_4516);
nor U5120 (N_5120,N_4761,N_4902);
and U5121 (N_5121,N_4936,N_4863);
and U5122 (N_5122,N_4594,N_4711);
nor U5123 (N_5123,N_4967,N_4646);
nand U5124 (N_5124,N_4547,N_4873);
nor U5125 (N_5125,N_4699,N_4577);
nand U5126 (N_5126,N_4649,N_4730);
and U5127 (N_5127,N_4995,N_4574);
xnor U5128 (N_5128,N_4664,N_4817);
and U5129 (N_5129,N_4764,N_4525);
and U5130 (N_5130,N_4551,N_4669);
nor U5131 (N_5131,N_4937,N_4832);
xnor U5132 (N_5132,N_4898,N_4671);
nor U5133 (N_5133,N_4901,N_4507);
or U5134 (N_5134,N_4688,N_4760);
nor U5135 (N_5135,N_4978,N_4815);
nand U5136 (N_5136,N_4912,N_4653);
xnor U5137 (N_5137,N_4784,N_4919);
nand U5138 (N_5138,N_4818,N_4765);
nor U5139 (N_5139,N_4573,N_4568);
and U5140 (N_5140,N_4522,N_4709);
or U5141 (N_5141,N_4876,N_4858);
and U5142 (N_5142,N_4527,N_4993);
or U5143 (N_5143,N_4994,N_4716);
xor U5144 (N_5144,N_4724,N_4903);
nand U5145 (N_5145,N_4782,N_4560);
nor U5146 (N_5146,N_4713,N_4750);
and U5147 (N_5147,N_4670,N_4511);
or U5148 (N_5148,N_4740,N_4733);
nor U5149 (N_5149,N_4570,N_4793);
nor U5150 (N_5150,N_4545,N_4501);
and U5151 (N_5151,N_4717,N_4555);
nand U5152 (N_5152,N_4889,N_4739);
xnor U5153 (N_5153,N_4541,N_4791);
nor U5154 (N_5154,N_4915,N_4776);
or U5155 (N_5155,N_4632,N_4992);
nand U5156 (N_5156,N_4925,N_4529);
nor U5157 (N_5157,N_4966,N_4960);
xnor U5158 (N_5158,N_4961,N_4563);
nor U5159 (N_5159,N_4657,N_4933);
and U5160 (N_5160,N_4848,N_4723);
and U5161 (N_5161,N_4634,N_4526);
or U5162 (N_5162,N_4857,N_4865);
or U5163 (N_5163,N_4965,N_4952);
xor U5164 (N_5164,N_4668,N_4710);
and U5165 (N_5165,N_4985,N_4707);
xor U5166 (N_5166,N_4833,N_4980);
xnor U5167 (N_5167,N_4977,N_4590);
and U5168 (N_5168,N_4886,N_4922);
nor U5169 (N_5169,N_4878,N_4548);
nor U5170 (N_5170,N_4609,N_4714);
nor U5171 (N_5171,N_4897,N_4973);
nor U5172 (N_5172,N_4955,N_4757);
or U5173 (N_5173,N_4604,N_4797);
xor U5174 (N_5174,N_4743,N_4850);
xnor U5175 (N_5175,N_4881,N_4939);
nor U5176 (N_5176,N_4862,N_4582);
nand U5177 (N_5177,N_4905,N_4708);
or U5178 (N_5178,N_4758,N_4988);
and U5179 (N_5179,N_4852,N_4627);
nor U5180 (N_5180,N_4931,N_4869);
xor U5181 (N_5181,N_4720,N_4622);
xnor U5182 (N_5182,N_4806,N_4945);
or U5183 (N_5183,N_4593,N_4924);
or U5184 (N_5184,N_4731,N_4819);
or U5185 (N_5185,N_4823,N_4938);
and U5186 (N_5186,N_4849,N_4694);
or U5187 (N_5187,N_4780,N_4927);
nor U5188 (N_5188,N_4578,N_4518);
xor U5189 (N_5189,N_4734,N_4956);
and U5190 (N_5190,N_4979,N_4597);
and U5191 (N_5191,N_4675,N_4517);
nor U5192 (N_5192,N_4728,N_4853);
nand U5193 (N_5193,N_4643,N_4928);
or U5194 (N_5194,N_4971,N_4523);
xnor U5195 (N_5195,N_4506,N_4519);
nor U5196 (N_5196,N_4755,N_4641);
nor U5197 (N_5197,N_4678,N_4549);
nand U5198 (N_5198,N_4696,N_4783);
or U5199 (N_5199,N_4744,N_4567);
nand U5200 (N_5200,N_4829,N_4899);
or U5201 (N_5201,N_4691,N_4840);
and U5202 (N_5202,N_4844,N_4990);
nand U5203 (N_5203,N_4695,N_4796);
nor U5204 (N_5204,N_4972,N_4914);
or U5205 (N_5205,N_4557,N_4801);
nor U5206 (N_5206,N_4648,N_4871);
xor U5207 (N_5207,N_4600,N_4954);
xor U5208 (N_5208,N_4502,N_4920);
or U5209 (N_5209,N_4631,N_4732);
nor U5210 (N_5210,N_4607,N_4825);
and U5211 (N_5211,N_4807,N_4909);
or U5212 (N_5212,N_4984,N_4581);
or U5213 (N_5213,N_4637,N_4785);
or U5214 (N_5214,N_4916,N_4767);
xor U5215 (N_5215,N_4763,N_4880);
and U5216 (N_5216,N_4885,N_4640);
nand U5217 (N_5217,N_4969,N_4805);
xnor U5218 (N_5218,N_4550,N_4565);
nor U5219 (N_5219,N_4804,N_4531);
xnor U5220 (N_5220,N_4515,N_4690);
xnor U5221 (N_5221,N_4751,N_4769);
and U5222 (N_5222,N_4851,N_4656);
and U5223 (N_5223,N_4884,N_4595);
and U5224 (N_5224,N_4794,N_4645);
xor U5225 (N_5225,N_4533,N_4727);
nor U5226 (N_5226,N_4566,N_4742);
or U5227 (N_5227,N_4958,N_4795);
xor U5228 (N_5228,N_4987,N_4619);
nand U5229 (N_5229,N_4864,N_4650);
and U5230 (N_5230,N_4544,N_4546);
and U5231 (N_5231,N_4569,N_4633);
nor U5232 (N_5232,N_4712,N_4562);
or U5233 (N_5233,N_4572,N_4592);
and U5234 (N_5234,N_4500,N_4838);
or U5235 (N_5235,N_4826,N_4679);
nor U5236 (N_5236,N_4943,N_4877);
nand U5237 (N_5237,N_4856,N_4606);
or U5238 (N_5238,N_4513,N_4583);
or U5239 (N_5239,N_4828,N_4976);
or U5240 (N_5240,N_4790,N_4554);
or U5241 (N_5241,N_4735,N_4623);
or U5242 (N_5242,N_4638,N_4859);
nand U5243 (N_5243,N_4935,N_4520);
xnor U5244 (N_5244,N_4771,N_4974);
and U5245 (N_5245,N_4539,N_4930);
or U5246 (N_5246,N_4778,N_4810);
nand U5247 (N_5247,N_4635,N_4706);
nand U5248 (N_5248,N_4687,N_4787);
xor U5249 (N_5249,N_4926,N_4845);
xnor U5250 (N_5250,N_4986,N_4693);
or U5251 (N_5251,N_4597,N_4691);
nand U5252 (N_5252,N_4852,N_4766);
nand U5253 (N_5253,N_4973,N_4590);
nor U5254 (N_5254,N_4683,N_4537);
nor U5255 (N_5255,N_4613,N_4780);
nor U5256 (N_5256,N_4858,N_4600);
nor U5257 (N_5257,N_4652,N_4598);
or U5258 (N_5258,N_4654,N_4966);
or U5259 (N_5259,N_4542,N_4829);
nand U5260 (N_5260,N_4876,N_4863);
or U5261 (N_5261,N_4935,N_4706);
xor U5262 (N_5262,N_4973,N_4992);
nor U5263 (N_5263,N_4598,N_4864);
and U5264 (N_5264,N_4626,N_4611);
nand U5265 (N_5265,N_4783,N_4877);
xor U5266 (N_5266,N_4731,N_4618);
and U5267 (N_5267,N_4905,N_4872);
or U5268 (N_5268,N_4720,N_4580);
nor U5269 (N_5269,N_4744,N_4509);
xor U5270 (N_5270,N_4541,N_4838);
nand U5271 (N_5271,N_4904,N_4620);
nor U5272 (N_5272,N_4564,N_4658);
nor U5273 (N_5273,N_4766,N_4554);
nor U5274 (N_5274,N_4847,N_4845);
nor U5275 (N_5275,N_4896,N_4981);
nor U5276 (N_5276,N_4906,N_4764);
or U5277 (N_5277,N_4891,N_4580);
xnor U5278 (N_5278,N_4674,N_4684);
or U5279 (N_5279,N_4782,N_4566);
or U5280 (N_5280,N_4902,N_4766);
and U5281 (N_5281,N_4821,N_4905);
and U5282 (N_5282,N_4778,N_4605);
nor U5283 (N_5283,N_4830,N_4842);
nand U5284 (N_5284,N_4546,N_4557);
and U5285 (N_5285,N_4861,N_4912);
xnor U5286 (N_5286,N_4736,N_4546);
nor U5287 (N_5287,N_4553,N_4957);
nor U5288 (N_5288,N_4979,N_4581);
xor U5289 (N_5289,N_4914,N_4750);
or U5290 (N_5290,N_4908,N_4518);
and U5291 (N_5291,N_4746,N_4861);
and U5292 (N_5292,N_4585,N_4937);
nand U5293 (N_5293,N_4828,N_4993);
nor U5294 (N_5294,N_4845,N_4633);
xnor U5295 (N_5295,N_4887,N_4739);
and U5296 (N_5296,N_4842,N_4769);
nand U5297 (N_5297,N_4748,N_4969);
or U5298 (N_5298,N_4798,N_4839);
nor U5299 (N_5299,N_4879,N_4615);
nand U5300 (N_5300,N_4526,N_4910);
xor U5301 (N_5301,N_4744,N_4801);
or U5302 (N_5302,N_4928,N_4616);
and U5303 (N_5303,N_4728,N_4933);
nand U5304 (N_5304,N_4863,N_4905);
xor U5305 (N_5305,N_4731,N_4891);
xor U5306 (N_5306,N_4722,N_4756);
xnor U5307 (N_5307,N_4835,N_4544);
nand U5308 (N_5308,N_4813,N_4748);
xnor U5309 (N_5309,N_4650,N_4660);
and U5310 (N_5310,N_4712,N_4564);
or U5311 (N_5311,N_4531,N_4932);
nor U5312 (N_5312,N_4561,N_4977);
or U5313 (N_5313,N_4629,N_4613);
nor U5314 (N_5314,N_4750,N_4688);
and U5315 (N_5315,N_4817,N_4614);
nand U5316 (N_5316,N_4831,N_4700);
nor U5317 (N_5317,N_4927,N_4665);
or U5318 (N_5318,N_4844,N_4792);
or U5319 (N_5319,N_4781,N_4804);
nor U5320 (N_5320,N_4926,N_4611);
nand U5321 (N_5321,N_4824,N_4663);
nor U5322 (N_5322,N_4987,N_4633);
and U5323 (N_5323,N_4675,N_4531);
nand U5324 (N_5324,N_4877,N_4656);
or U5325 (N_5325,N_4512,N_4567);
xor U5326 (N_5326,N_4940,N_4523);
nand U5327 (N_5327,N_4644,N_4720);
xnor U5328 (N_5328,N_4613,N_4913);
nand U5329 (N_5329,N_4889,N_4917);
xnor U5330 (N_5330,N_4978,N_4526);
nor U5331 (N_5331,N_4977,N_4608);
or U5332 (N_5332,N_4930,N_4583);
or U5333 (N_5333,N_4843,N_4854);
nand U5334 (N_5334,N_4625,N_4963);
xor U5335 (N_5335,N_4754,N_4934);
nand U5336 (N_5336,N_4937,N_4587);
nand U5337 (N_5337,N_4606,N_4870);
nand U5338 (N_5338,N_4962,N_4691);
xor U5339 (N_5339,N_4558,N_4802);
and U5340 (N_5340,N_4789,N_4821);
nand U5341 (N_5341,N_4925,N_4698);
or U5342 (N_5342,N_4888,N_4554);
nor U5343 (N_5343,N_4876,N_4926);
xor U5344 (N_5344,N_4542,N_4872);
xnor U5345 (N_5345,N_4720,N_4573);
or U5346 (N_5346,N_4921,N_4936);
nor U5347 (N_5347,N_4976,N_4630);
and U5348 (N_5348,N_4951,N_4625);
or U5349 (N_5349,N_4882,N_4731);
nor U5350 (N_5350,N_4698,N_4643);
nand U5351 (N_5351,N_4935,N_4640);
nor U5352 (N_5352,N_4835,N_4710);
nand U5353 (N_5353,N_4727,N_4620);
and U5354 (N_5354,N_4940,N_4825);
and U5355 (N_5355,N_4829,N_4824);
nor U5356 (N_5356,N_4748,N_4568);
or U5357 (N_5357,N_4540,N_4815);
nor U5358 (N_5358,N_4984,N_4964);
or U5359 (N_5359,N_4521,N_4777);
nand U5360 (N_5360,N_4502,N_4531);
xor U5361 (N_5361,N_4573,N_4638);
nand U5362 (N_5362,N_4633,N_4644);
and U5363 (N_5363,N_4707,N_4998);
nor U5364 (N_5364,N_4567,N_4546);
xor U5365 (N_5365,N_4904,N_4963);
nand U5366 (N_5366,N_4874,N_4696);
and U5367 (N_5367,N_4724,N_4760);
nand U5368 (N_5368,N_4677,N_4851);
xnor U5369 (N_5369,N_4746,N_4541);
xor U5370 (N_5370,N_4949,N_4919);
nand U5371 (N_5371,N_4708,N_4939);
nand U5372 (N_5372,N_4781,N_4885);
xnor U5373 (N_5373,N_4857,N_4550);
nor U5374 (N_5374,N_4729,N_4961);
and U5375 (N_5375,N_4529,N_4663);
xnor U5376 (N_5376,N_4837,N_4818);
nand U5377 (N_5377,N_4699,N_4823);
xor U5378 (N_5378,N_4583,N_4515);
xnor U5379 (N_5379,N_4758,N_4606);
xor U5380 (N_5380,N_4900,N_4854);
nand U5381 (N_5381,N_4531,N_4622);
nor U5382 (N_5382,N_4575,N_4756);
and U5383 (N_5383,N_4856,N_4583);
and U5384 (N_5384,N_4708,N_4825);
or U5385 (N_5385,N_4639,N_4974);
or U5386 (N_5386,N_4693,N_4870);
nor U5387 (N_5387,N_4538,N_4795);
or U5388 (N_5388,N_4740,N_4782);
or U5389 (N_5389,N_4895,N_4828);
and U5390 (N_5390,N_4512,N_4552);
xor U5391 (N_5391,N_4880,N_4670);
and U5392 (N_5392,N_4811,N_4838);
nor U5393 (N_5393,N_4841,N_4874);
xnor U5394 (N_5394,N_4754,N_4981);
xor U5395 (N_5395,N_4945,N_4579);
nor U5396 (N_5396,N_4771,N_4815);
and U5397 (N_5397,N_4775,N_4857);
and U5398 (N_5398,N_4510,N_4570);
nand U5399 (N_5399,N_4874,N_4662);
nand U5400 (N_5400,N_4761,N_4859);
xor U5401 (N_5401,N_4907,N_4953);
or U5402 (N_5402,N_4584,N_4712);
xnor U5403 (N_5403,N_4565,N_4573);
or U5404 (N_5404,N_4906,N_4941);
xor U5405 (N_5405,N_4740,N_4920);
nor U5406 (N_5406,N_4633,N_4591);
or U5407 (N_5407,N_4844,N_4793);
nand U5408 (N_5408,N_4521,N_4634);
and U5409 (N_5409,N_4700,N_4938);
and U5410 (N_5410,N_4565,N_4704);
xnor U5411 (N_5411,N_4589,N_4824);
and U5412 (N_5412,N_4822,N_4920);
or U5413 (N_5413,N_4583,N_4908);
nor U5414 (N_5414,N_4791,N_4927);
or U5415 (N_5415,N_4973,N_4615);
nor U5416 (N_5416,N_4702,N_4999);
nor U5417 (N_5417,N_4557,N_4888);
nor U5418 (N_5418,N_4670,N_4717);
and U5419 (N_5419,N_4507,N_4580);
or U5420 (N_5420,N_4559,N_4905);
or U5421 (N_5421,N_4976,N_4506);
xor U5422 (N_5422,N_4801,N_4993);
nor U5423 (N_5423,N_4845,N_4848);
and U5424 (N_5424,N_4741,N_4597);
nand U5425 (N_5425,N_4805,N_4799);
or U5426 (N_5426,N_4702,N_4781);
nand U5427 (N_5427,N_4770,N_4598);
xor U5428 (N_5428,N_4931,N_4971);
and U5429 (N_5429,N_4532,N_4759);
or U5430 (N_5430,N_4816,N_4738);
and U5431 (N_5431,N_4636,N_4995);
xor U5432 (N_5432,N_4883,N_4706);
nor U5433 (N_5433,N_4557,N_4588);
nand U5434 (N_5434,N_4554,N_4541);
and U5435 (N_5435,N_4640,N_4532);
nand U5436 (N_5436,N_4581,N_4994);
and U5437 (N_5437,N_4684,N_4866);
nand U5438 (N_5438,N_4799,N_4826);
nand U5439 (N_5439,N_4784,N_4699);
and U5440 (N_5440,N_4873,N_4612);
nand U5441 (N_5441,N_4616,N_4821);
xnor U5442 (N_5442,N_4682,N_4532);
xor U5443 (N_5443,N_4661,N_4715);
and U5444 (N_5444,N_4809,N_4807);
or U5445 (N_5445,N_4876,N_4603);
and U5446 (N_5446,N_4628,N_4797);
xnor U5447 (N_5447,N_4647,N_4775);
nand U5448 (N_5448,N_4997,N_4622);
nand U5449 (N_5449,N_4613,N_4805);
or U5450 (N_5450,N_4839,N_4736);
nand U5451 (N_5451,N_4990,N_4532);
xnor U5452 (N_5452,N_4712,N_4959);
or U5453 (N_5453,N_4738,N_4743);
nand U5454 (N_5454,N_4895,N_4686);
and U5455 (N_5455,N_4545,N_4978);
and U5456 (N_5456,N_4997,N_4540);
xnor U5457 (N_5457,N_4878,N_4500);
or U5458 (N_5458,N_4578,N_4879);
or U5459 (N_5459,N_4574,N_4909);
and U5460 (N_5460,N_4879,N_4980);
nor U5461 (N_5461,N_4643,N_4970);
xor U5462 (N_5462,N_4876,N_4867);
nor U5463 (N_5463,N_4740,N_4658);
xnor U5464 (N_5464,N_4896,N_4670);
nand U5465 (N_5465,N_4568,N_4643);
nor U5466 (N_5466,N_4992,N_4538);
or U5467 (N_5467,N_4973,N_4665);
and U5468 (N_5468,N_4819,N_4828);
xor U5469 (N_5469,N_4958,N_4538);
nor U5470 (N_5470,N_4972,N_4758);
and U5471 (N_5471,N_4500,N_4983);
or U5472 (N_5472,N_4816,N_4542);
nor U5473 (N_5473,N_4963,N_4997);
and U5474 (N_5474,N_4858,N_4844);
nand U5475 (N_5475,N_4951,N_4824);
and U5476 (N_5476,N_4922,N_4880);
nor U5477 (N_5477,N_4698,N_4748);
or U5478 (N_5478,N_4997,N_4570);
and U5479 (N_5479,N_4966,N_4550);
or U5480 (N_5480,N_4991,N_4657);
nor U5481 (N_5481,N_4726,N_4582);
xor U5482 (N_5482,N_4838,N_4681);
xnor U5483 (N_5483,N_4867,N_4894);
xnor U5484 (N_5484,N_4501,N_4713);
xnor U5485 (N_5485,N_4642,N_4946);
and U5486 (N_5486,N_4688,N_4502);
or U5487 (N_5487,N_4830,N_4677);
and U5488 (N_5488,N_4512,N_4892);
and U5489 (N_5489,N_4536,N_4790);
nor U5490 (N_5490,N_4603,N_4983);
nand U5491 (N_5491,N_4599,N_4989);
and U5492 (N_5492,N_4788,N_4908);
or U5493 (N_5493,N_4883,N_4510);
or U5494 (N_5494,N_4656,N_4763);
xor U5495 (N_5495,N_4634,N_4660);
xor U5496 (N_5496,N_4623,N_4851);
and U5497 (N_5497,N_4517,N_4658);
xnor U5498 (N_5498,N_4561,N_4549);
and U5499 (N_5499,N_4858,N_4945);
xor U5500 (N_5500,N_5130,N_5136);
nor U5501 (N_5501,N_5091,N_5341);
and U5502 (N_5502,N_5240,N_5206);
xor U5503 (N_5503,N_5405,N_5114);
and U5504 (N_5504,N_5155,N_5330);
xnor U5505 (N_5505,N_5318,N_5342);
nor U5506 (N_5506,N_5243,N_5310);
and U5507 (N_5507,N_5456,N_5477);
or U5508 (N_5508,N_5192,N_5375);
or U5509 (N_5509,N_5436,N_5270);
nand U5510 (N_5510,N_5175,N_5075);
nand U5511 (N_5511,N_5464,N_5413);
and U5512 (N_5512,N_5360,N_5095);
xor U5513 (N_5513,N_5268,N_5150);
and U5514 (N_5514,N_5218,N_5471);
and U5515 (N_5515,N_5197,N_5368);
nand U5516 (N_5516,N_5497,N_5339);
xor U5517 (N_5517,N_5242,N_5458);
xor U5518 (N_5518,N_5113,N_5427);
nand U5519 (N_5519,N_5381,N_5323);
nand U5520 (N_5520,N_5221,N_5418);
nand U5521 (N_5521,N_5306,N_5085);
or U5522 (N_5522,N_5467,N_5146);
nand U5523 (N_5523,N_5144,N_5369);
nor U5524 (N_5524,N_5217,N_5331);
or U5525 (N_5525,N_5069,N_5321);
xnor U5526 (N_5526,N_5058,N_5292);
and U5527 (N_5527,N_5042,N_5047);
nor U5528 (N_5528,N_5241,N_5393);
nand U5529 (N_5529,N_5401,N_5455);
or U5530 (N_5530,N_5134,N_5064);
nor U5531 (N_5531,N_5082,N_5067);
nor U5532 (N_5532,N_5450,N_5459);
nor U5533 (N_5533,N_5283,N_5382);
and U5534 (N_5534,N_5356,N_5475);
xor U5535 (N_5535,N_5311,N_5016);
nand U5536 (N_5536,N_5320,N_5127);
and U5537 (N_5537,N_5279,N_5380);
xor U5538 (N_5538,N_5207,N_5313);
nand U5539 (N_5539,N_5247,N_5244);
nor U5540 (N_5540,N_5271,N_5407);
nand U5541 (N_5541,N_5389,N_5005);
xnor U5542 (N_5542,N_5423,N_5481);
nor U5543 (N_5543,N_5319,N_5084);
nor U5544 (N_5544,N_5294,N_5024);
and U5545 (N_5545,N_5037,N_5433);
or U5546 (N_5546,N_5326,N_5062);
or U5547 (N_5547,N_5183,N_5489);
and U5548 (N_5548,N_5296,N_5374);
xnor U5549 (N_5549,N_5073,N_5122);
and U5550 (N_5550,N_5081,N_5088);
nand U5551 (N_5551,N_5052,N_5324);
nor U5552 (N_5552,N_5300,N_5487);
and U5553 (N_5553,N_5055,N_5430);
xnor U5554 (N_5554,N_5246,N_5226);
xor U5555 (N_5555,N_5090,N_5302);
and U5556 (N_5556,N_5277,N_5143);
nand U5557 (N_5557,N_5275,N_5280);
or U5558 (N_5558,N_5424,N_5220);
xnor U5559 (N_5559,N_5057,N_5404);
nor U5560 (N_5560,N_5013,N_5045);
and U5561 (N_5561,N_5317,N_5435);
nor U5562 (N_5562,N_5021,N_5204);
xor U5563 (N_5563,N_5256,N_5149);
and U5564 (N_5564,N_5291,N_5499);
nand U5565 (N_5565,N_5128,N_5139);
and U5566 (N_5566,N_5138,N_5030);
nand U5567 (N_5567,N_5309,N_5012);
or U5568 (N_5568,N_5232,N_5169);
nand U5569 (N_5569,N_5031,N_5225);
nand U5570 (N_5570,N_5019,N_5412);
nor U5571 (N_5571,N_5336,N_5432);
xor U5572 (N_5572,N_5308,N_5403);
nor U5573 (N_5573,N_5325,N_5262);
nand U5574 (N_5574,N_5202,N_5109);
nand U5575 (N_5575,N_5181,N_5337);
nand U5576 (N_5576,N_5008,N_5453);
nor U5577 (N_5577,N_5440,N_5495);
nand U5578 (N_5578,N_5186,N_5190);
nand U5579 (N_5579,N_5429,N_5224);
xnor U5580 (N_5580,N_5026,N_5480);
xnor U5581 (N_5581,N_5223,N_5102);
xor U5582 (N_5582,N_5040,N_5269);
xor U5583 (N_5583,N_5153,N_5361);
xor U5584 (N_5584,N_5151,N_5002);
and U5585 (N_5585,N_5120,N_5406);
and U5586 (N_5586,N_5060,N_5355);
nor U5587 (N_5587,N_5473,N_5391);
nor U5588 (N_5588,N_5235,N_5379);
xor U5589 (N_5589,N_5288,N_5438);
and U5590 (N_5590,N_5056,N_5168);
nor U5591 (N_5591,N_5101,N_5295);
nand U5592 (N_5592,N_5108,N_5080);
nand U5593 (N_5593,N_5007,N_5219);
nand U5594 (N_5594,N_5209,N_5408);
xnor U5595 (N_5595,N_5451,N_5478);
nor U5596 (N_5596,N_5216,N_5099);
xnor U5597 (N_5597,N_5327,N_5170);
and U5598 (N_5598,N_5188,N_5133);
nor U5599 (N_5599,N_5043,N_5135);
and U5600 (N_5600,N_5034,N_5329);
xor U5601 (N_5601,N_5274,N_5299);
or U5602 (N_5602,N_5365,N_5184);
and U5603 (N_5603,N_5293,N_5472);
xor U5604 (N_5604,N_5328,N_5041);
nand U5605 (N_5605,N_5431,N_5350);
xor U5606 (N_5606,N_5322,N_5098);
nand U5607 (N_5607,N_5257,N_5196);
xnor U5608 (N_5608,N_5213,N_5287);
xor U5609 (N_5609,N_5238,N_5236);
nor U5610 (N_5610,N_5035,N_5063);
nor U5611 (N_5611,N_5398,N_5419);
and U5612 (N_5612,N_5145,N_5415);
nand U5613 (N_5613,N_5033,N_5229);
nor U5614 (N_5614,N_5373,N_5001);
and U5615 (N_5615,N_5061,N_5089);
nor U5616 (N_5616,N_5364,N_5290);
or U5617 (N_5617,N_5178,N_5399);
xor U5618 (N_5618,N_5441,N_5346);
nand U5619 (N_5619,N_5140,N_5121);
and U5620 (N_5620,N_5068,N_5189);
nor U5621 (N_5621,N_5230,N_5263);
and U5622 (N_5622,N_5039,N_5316);
nand U5623 (N_5623,N_5484,N_5416);
nor U5624 (N_5624,N_5286,N_5006);
nor U5625 (N_5625,N_5023,N_5193);
or U5626 (N_5626,N_5402,N_5254);
nor U5627 (N_5627,N_5461,N_5264);
or U5628 (N_5628,N_5352,N_5173);
xnor U5629 (N_5629,N_5179,N_5417);
nand U5630 (N_5630,N_5191,N_5434);
nand U5631 (N_5631,N_5386,N_5298);
and U5632 (N_5632,N_5260,N_5180);
xor U5633 (N_5633,N_5425,N_5083);
xor U5634 (N_5634,N_5029,N_5383);
and U5635 (N_5635,N_5333,N_5428);
or U5636 (N_5636,N_5131,N_5314);
or U5637 (N_5637,N_5396,N_5200);
nand U5638 (N_5638,N_5071,N_5214);
and U5639 (N_5639,N_5048,N_5359);
xor U5640 (N_5640,N_5237,N_5493);
nor U5641 (N_5641,N_5111,N_5312);
or U5642 (N_5642,N_5259,N_5228);
and U5643 (N_5643,N_5367,N_5129);
nor U5644 (N_5644,N_5258,N_5152);
nand U5645 (N_5645,N_5172,N_5483);
and U5646 (N_5646,N_5362,N_5276);
or U5647 (N_5647,N_5304,N_5148);
nand U5648 (N_5648,N_5462,N_5249);
and U5649 (N_5649,N_5390,N_5198);
nand U5650 (N_5650,N_5465,N_5115);
nor U5651 (N_5651,N_5053,N_5201);
nor U5652 (N_5652,N_5015,N_5025);
nand U5653 (N_5653,N_5385,N_5490);
xor U5654 (N_5654,N_5491,N_5156);
xor U5655 (N_5655,N_5100,N_5273);
and U5656 (N_5656,N_5018,N_5446);
and U5657 (N_5657,N_5059,N_5301);
nand U5658 (N_5658,N_5124,N_5103);
nand U5659 (N_5659,N_5315,N_5421);
nor U5660 (N_5660,N_5051,N_5496);
or U5661 (N_5661,N_5332,N_5203);
and U5662 (N_5662,N_5261,N_5482);
xnor U5663 (N_5663,N_5439,N_5066);
and U5664 (N_5664,N_5255,N_5392);
xnor U5665 (N_5665,N_5160,N_5466);
or U5666 (N_5666,N_5376,N_5074);
and U5667 (N_5667,N_5445,N_5227);
nor U5668 (N_5668,N_5366,N_5038);
nand U5669 (N_5669,N_5278,N_5400);
xnor U5670 (N_5670,N_5253,N_5234);
nor U5671 (N_5671,N_5265,N_5094);
and U5672 (N_5672,N_5447,N_5284);
nand U5673 (N_5673,N_5022,N_5092);
or U5674 (N_5674,N_5251,N_5372);
xor U5675 (N_5675,N_5165,N_5028);
nand U5676 (N_5676,N_5289,N_5159);
nand U5677 (N_5677,N_5387,N_5104);
nor U5678 (N_5678,N_5065,N_5454);
nor U5679 (N_5679,N_5036,N_5443);
or U5680 (N_5680,N_5351,N_5394);
xnor U5681 (N_5681,N_5303,N_5378);
and U5682 (N_5682,N_5344,N_5334);
nand U5683 (N_5683,N_5017,N_5486);
xor U5684 (N_5684,N_5117,N_5046);
nand U5685 (N_5685,N_5164,N_5281);
and U5686 (N_5686,N_5370,N_5363);
and U5687 (N_5687,N_5414,N_5014);
or U5688 (N_5688,N_5116,N_5195);
nor U5689 (N_5689,N_5215,N_5498);
or U5690 (N_5690,N_5132,N_5449);
or U5691 (N_5691,N_5087,N_5347);
xnor U5692 (N_5692,N_5492,N_5272);
and U5693 (N_5693,N_5166,N_5452);
nand U5694 (N_5694,N_5476,N_5105);
xor U5695 (N_5695,N_5126,N_5070);
nand U5696 (N_5696,N_5171,N_5282);
nor U5697 (N_5697,N_5010,N_5354);
nand U5698 (N_5698,N_5032,N_5123);
and U5699 (N_5699,N_5106,N_5371);
nor U5700 (N_5700,N_5463,N_5147);
nand U5701 (N_5701,N_5410,N_5422);
nor U5702 (N_5702,N_5488,N_5470);
or U5703 (N_5703,N_5093,N_5177);
nor U5704 (N_5704,N_5485,N_5266);
xnor U5705 (N_5705,N_5076,N_5110);
or U5706 (N_5706,N_5125,N_5137);
nor U5707 (N_5707,N_5285,N_5158);
xnor U5708 (N_5708,N_5118,N_5444);
nor U5709 (N_5709,N_5112,N_5077);
nor U5710 (N_5710,N_5267,N_5163);
nor U5711 (N_5711,N_5162,N_5161);
xor U5712 (N_5712,N_5020,N_5377);
and U5713 (N_5713,N_5460,N_5468);
and U5714 (N_5714,N_5194,N_5174);
and U5715 (N_5715,N_5011,N_5009);
nand U5716 (N_5716,N_5211,N_5297);
nand U5717 (N_5717,N_5049,N_5167);
nand U5718 (N_5718,N_5054,N_5239);
and U5719 (N_5719,N_5426,N_5307);
or U5720 (N_5720,N_5479,N_5086);
xnor U5721 (N_5721,N_5335,N_5141);
and U5722 (N_5722,N_5199,N_5494);
and U5723 (N_5723,N_5409,N_5182);
and U5724 (N_5724,N_5119,N_5222);
or U5725 (N_5725,N_5044,N_5388);
and U5726 (N_5726,N_5395,N_5208);
xor U5727 (N_5727,N_5096,N_5343);
xnor U5728 (N_5728,N_5420,N_5107);
nor U5729 (N_5729,N_5340,N_5079);
nand U5730 (N_5730,N_5353,N_5384);
nand U5731 (N_5731,N_5050,N_5474);
xnor U5732 (N_5732,N_5072,N_5078);
xor U5733 (N_5733,N_5252,N_5231);
nor U5734 (N_5734,N_5176,N_5397);
and U5735 (N_5735,N_5437,N_5448);
or U5736 (N_5736,N_5411,N_5210);
xor U5737 (N_5737,N_5157,N_5305);
and U5738 (N_5738,N_5245,N_5000);
xnor U5739 (N_5739,N_5154,N_5004);
or U5740 (N_5740,N_5003,N_5349);
xor U5741 (N_5741,N_5027,N_5348);
or U5742 (N_5742,N_5250,N_5457);
or U5743 (N_5743,N_5185,N_5212);
or U5744 (N_5744,N_5248,N_5338);
nand U5745 (N_5745,N_5097,N_5358);
and U5746 (N_5746,N_5142,N_5233);
xor U5747 (N_5747,N_5442,N_5357);
and U5748 (N_5748,N_5345,N_5187);
xnor U5749 (N_5749,N_5469,N_5205);
xor U5750 (N_5750,N_5398,N_5003);
nor U5751 (N_5751,N_5083,N_5201);
nor U5752 (N_5752,N_5163,N_5358);
or U5753 (N_5753,N_5068,N_5169);
nor U5754 (N_5754,N_5354,N_5039);
nand U5755 (N_5755,N_5362,N_5056);
and U5756 (N_5756,N_5338,N_5185);
or U5757 (N_5757,N_5052,N_5282);
and U5758 (N_5758,N_5203,N_5067);
and U5759 (N_5759,N_5035,N_5199);
and U5760 (N_5760,N_5240,N_5409);
nor U5761 (N_5761,N_5294,N_5198);
nand U5762 (N_5762,N_5495,N_5273);
or U5763 (N_5763,N_5079,N_5449);
nor U5764 (N_5764,N_5237,N_5133);
nand U5765 (N_5765,N_5351,N_5249);
nand U5766 (N_5766,N_5410,N_5388);
or U5767 (N_5767,N_5105,N_5422);
nand U5768 (N_5768,N_5200,N_5177);
nor U5769 (N_5769,N_5299,N_5166);
nor U5770 (N_5770,N_5255,N_5228);
and U5771 (N_5771,N_5358,N_5029);
or U5772 (N_5772,N_5451,N_5414);
or U5773 (N_5773,N_5314,N_5032);
or U5774 (N_5774,N_5121,N_5124);
nand U5775 (N_5775,N_5112,N_5276);
or U5776 (N_5776,N_5100,N_5245);
or U5777 (N_5777,N_5021,N_5140);
xor U5778 (N_5778,N_5202,N_5251);
or U5779 (N_5779,N_5351,N_5484);
or U5780 (N_5780,N_5460,N_5060);
nand U5781 (N_5781,N_5420,N_5036);
nor U5782 (N_5782,N_5018,N_5237);
or U5783 (N_5783,N_5220,N_5006);
or U5784 (N_5784,N_5355,N_5412);
nor U5785 (N_5785,N_5182,N_5341);
and U5786 (N_5786,N_5405,N_5343);
or U5787 (N_5787,N_5227,N_5042);
nor U5788 (N_5788,N_5116,N_5425);
or U5789 (N_5789,N_5284,N_5283);
xor U5790 (N_5790,N_5294,N_5277);
or U5791 (N_5791,N_5397,N_5255);
nor U5792 (N_5792,N_5218,N_5317);
xnor U5793 (N_5793,N_5122,N_5264);
nor U5794 (N_5794,N_5436,N_5155);
xnor U5795 (N_5795,N_5054,N_5107);
and U5796 (N_5796,N_5348,N_5142);
xnor U5797 (N_5797,N_5373,N_5008);
or U5798 (N_5798,N_5410,N_5318);
nor U5799 (N_5799,N_5033,N_5030);
and U5800 (N_5800,N_5211,N_5456);
or U5801 (N_5801,N_5220,N_5299);
xor U5802 (N_5802,N_5282,N_5039);
nand U5803 (N_5803,N_5108,N_5382);
nand U5804 (N_5804,N_5447,N_5245);
or U5805 (N_5805,N_5351,N_5184);
nand U5806 (N_5806,N_5096,N_5119);
nand U5807 (N_5807,N_5381,N_5364);
or U5808 (N_5808,N_5165,N_5477);
or U5809 (N_5809,N_5323,N_5054);
nor U5810 (N_5810,N_5223,N_5246);
nor U5811 (N_5811,N_5094,N_5138);
xnor U5812 (N_5812,N_5479,N_5054);
and U5813 (N_5813,N_5451,N_5197);
xnor U5814 (N_5814,N_5023,N_5269);
nor U5815 (N_5815,N_5119,N_5297);
nand U5816 (N_5816,N_5472,N_5122);
xnor U5817 (N_5817,N_5440,N_5181);
or U5818 (N_5818,N_5167,N_5323);
nand U5819 (N_5819,N_5428,N_5026);
nand U5820 (N_5820,N_5228,N_5083);
nor U5821 (N_5821,N_5229,N_5014);
and U5822 (N_5822,N_5246,N_5477);
nor U5823 (N_5823,N_5109,N_5462);
nor U5824 (N_5824,N_5392,N_5036);
nor U5825 (N_5825,N_5052,N_5064);
and U5826 (N_5826,N_5168,N_5080);
or U5827 (N_5827,N_5120,N_5069);
nor U5828 (N_5828,N_5016,N_5088);
nor U5829 (N_5829,N_5274,N_5036);
or U5830 (N_5830,N_5410,N_5456);
nand U5831 (N_5831,N_5101,N_5418);
nor U5832 (N_5832,N_5111,N_5319);
and U5833 (N_5833,N_5240,N_5342);
nand U5834 (N_5834,N_5408,N_5442);
nand U5835 (N_5835,N_5173,N_5134);
nor U5836 (N_5836,N_5486,N_5112);
nor U5837 (N_5837,N_5471,N_5148);
nor U5838 (N_5838,N_5410,N_5257);
or U5839 (N_5839,N_5469,N_5454);
xor U5840 (N_5840,N_5471,N_5261);
or U5841 (N_5841,N_5072,N_5383);
or U5842 (N_5842,N_5169,N_5195);
and U5843 (N_5843,N_5162,N_5284);
nor U5844 (N_5844,N_5330,N_5447);
nand U5845 (N_5845,N_5053,N_5385);
nand U5846 (N_5846,N_5479,N_5285);
nor U5847 (N_5847,N_5379,N_5177);
xor U5848 (N_5848,N_5125,N_5402);
or U5849 (N_5849,N_5477,N_5070);
nor U5850 (N_5850,N_5188,N_5127);
and U5851 (N_5851,N_5454,N_5317);
or U5852 (N_5852,N_5178,N_5309);
nand U5853 (N_5853,N_5316,N_5409);
nor U5854 (N_5854,N_5094,N_5219);
nand U5855 (N_5855,N_5274,N_5145);
nor U5856 (N_5856,N_5470,N_5237);
nor U5857 (N_5857,N_5110,N_5121);
or U5858 (N_5858,N_5002,N_5177);
or U5859 (N_5859,N_5374,N_5124);
or U5860 (N_5860,N_5443,N_5453);
or U5861 (N_5861,N_5230,N_5339);
or U5862 (N_5862,N_5183,N_5330);
xnor U5863 (N_5863,N_5262,N_5393);
nor U5864 (N_5864,N_5185,N_5038);
and U5865 (N_5865,N_5309,N_5380);
or U5866 (N_5866,N_5445,N_5036);
nor U5867 (N_5867,N_5225,N_5183);
and U5868 (N_5868,N_5106,N_5133);
or U5869 (N_5869,N_5352,N_5122);
nand U5870 (N_5870,N_5406,N_5295);
nor U5871 (N_5871,N_5280,N_5353);
xor U5872 (N_5872,N_5173,N_5088);
or U5873 (N_5873,N_5079,N_5423);
xnor U5874 (N_5874,N_5236,N_5453);
or U5875 (N_5875,N_5196,N_5052);
xnor U5876 (N_5876,N_5329,N_5192);
or U5877 (N_5877,N_5082,N_5299);
or U5878 (N_5878,N_5433,N_5292);
and U5879 (N_5879,N_5286,N_5198);
nand U5880 (N_5880,N_5344,N_5330);
and U5881 (N_5881,N_5434,N_5165);
or U5882 (N_5882,N_5305,N_5219);
nand U5883 (N_5883,N_5420,N_5262);
and U5884 (N_5884,N_5167,N_5432);
nor U5885 (N_5885,N_5175,N_5104);
or U5886 (N_5886,N_5205,N_5224);
nand U5887 (N_5887,N_5270,N_5439);
and U5888 (N_5888,N_5398,N_5390);
and U5889 (N_5889,N_5218,N_5465);
nor U5890 (N_5890,N_5326,N_5116);
and U5891 (N_5891,N_5152,N_5143);
xor U5892 (N_5892,N_5272,N_5073);
xnor U5893 (N_5893,N_5345,N_5005);
nor U5894 (N_5894,N_5185,N_5010);
nand U5895 (N_5895,N_5417,N_5278);
nand U5896 (N_5896,N_5463,N_5076);
and U5897 (N_5897,N_5250,N_5355);
xnor U5898 (N_5898,N_5019,N_5419);
nand U5899 (N_5899,N_5080,N_5237);
and U5900 (N_5900,N_5298,N_5345);
nand U5901 (N_5901,N_5195,N_5092);
nand U5902 (N_5902,N_5434,N_5081);
nand U5903 (N_5903,N_5198,N_5422);
nand U5904 (N_5904,N_5417,N_5127);
and U5905 (N_5905,N_5370,N_5220);
or U5906 (N_5906,N_5485,N_5424);
and U5907 (N_5907,N_5002,N_5024);
nor U5908 (N_5908,N_5223,N_5292);
xor U5909 (N_5909,N_5212,N_5335);
nor U5910 (N_5910,N_5258,N_5486);
nand U5911 (N_5911,N_5199,N_5309);
nand U5912 (N_5912,N_5014,N_5032);
nand U5913 (N_5913,N_5153,N_5215);
and U5914 (N_5914,N_5289,N_5475);
and U5915 (N_5915,N_5109,N_5048);
or U5916 (N_5916,N_5077,N_5380);
nor U5917 (N_5917,N_5373,N_5169);
xor U5918 (N_5918,N_5466,N_5190);
nand U5919 (N_5919,N_5259,N_5374);
xnor U5920 (N_5920,N_5012,N_5133);
and U5921 (N_5921,N_5233,N_5225);
or U5922 (N_5922,N_5323,N_5428);
and U5923 (N_5923,N_5107,N_5461);
nor U5924 (N_5924,N_5099,N_5175);
or U5925 (N_5925,N_5367,N_5441);
xor U5926 (N_5926,N_5454,N_5286);
xnor U5927 (N_5927,N_5073,N_5265);
xnor U5928 (N_5928,N_5328,N_5068);
nand U5929 (N_5929,N_5179,N_5282);
nand U5930 (N_5930,N_5385,N_5446);
nand U5931 (N_5931,N_5114,N_5467);
xnor U5932 (N_5932,N_5379,N_5381);
xnor U5933 (N_5933,N_5091,N_5280);
nand U5934 (N_5934,N_5376,N_5423);
nor U5935 (N_5935,N_5416,N_5355);
and U5936 (N_5936,N_5110,N_5417);
and U5937 (N_5937,N_5051,N_5086);
nand U5938 (N_5938,N_5128,N_5248);
nand U5939 (N_5939,N_5388,N_5227);
nand U5940 (N_5940,N_5443,N_5172);
nor U5941 (N_5941,N_5035,N_5021);
nand U5942 (N_5942,N_5314,N_5293);
and U5943 (N_5943,N_5316,N_5051);
and U5944 (N_5944,N_5412,N_5342);
xnor U5945 (N_5945,N_5097,N_5489);
nand U5946 (N_5946,N_5278,N_5066);
nor U5947 (N_5947,N_5098,N_5342);
and U5948 (N_5948,N_5073,N_5362);
xnor U5949 (N_5949,N_5074,N_5437);
or U5950 (N_5950,N_5281,N_5483);
nor U5951 (N_5951,N_5434,N_5248);
and U5952 (N_5952,N_5053,N_5196);
xor U5953 (N_5953,N_5412,N_5211);
xnor U5954 (N_5954,N_5237,N_5444);
and U5955 (N_5955,N_5274,N_5128);
and U5956 (N_5956,N_5066,N_5207);
nor U5957 (N_5957,N_5169,N_5099);
nand U5958 (N_5958,N_5043,N_5033);
nor U5959 (N_5959,N_5187,N_5112);
or U5960 (N_5960,N_5301,N_5105);
and U5961 (N_5961,N_5268,N_5054);
nand U5962 (N_5962,N_5163,N_5137);
and U5963 (N_5963,N_5367,N_5048);
and U5964 (N_5964,N_5106,N_5072);
nand U5965 (N_5965,N_5457,N_5203);
xnor U5966 (N_5966,N_5049,N_5192);
nand U5967 (N_5967,N_5399,N_5235);
xnor U5968 (N_5968,N_5041,N_5238);
and U5969 (N_5969,N_5147,N_5148);
nor U5970 (N_5970,N_5107,N_5185);
xnor U5971 (N_5971,N_5490,N_5022);
nor U5972 (N_5972,N_5293,N_5161);
xnor U5973 (N_5973,N_5033,N_5481);
xor U5974 (N_5974,N_5253,N_5163);
nor U5975 (N_5975,N_5072,N_5354);
or U5976 (N_5976,N_5256,N_5329);
or U5977 (N_5977,N_5065,N_5473);
and U5978 (N_5978,N_5169,N_5338);
nor U5979 (N_5979,N_5372,N_5375);
or U5980 (N_5980,N_5423,N_5331);
nand U5981 (N_5981,N_5215,N_5073);
and U5982 (N_5982,N_5475,N_5343);
or U5983 (N_5983,N_5169,N_5035);
nor U5984 (N_5984,N_5422,N_5241);
nand U5985 (N_5985,N_5263,N_5217);
or U5986 (N_5986,N_5481,N_5059);
nor U5987 (N_5987,N_5180,N_5155);
and U5988 (N_5988,N_5131,N_5243);
or U5989 (N_5989,N_5482,N_5331);
nand U5990 (N_5990,N_5061,N_5057);
and U5991 (N_5991,N_5177,N_5040);
nand U5992 (N_5992,N_5205,N_5297);
and U5993 (N_5993,N_5485,N_5197);
and U5994 (N_5994,N_5295,N_5206);
xnor U5995 (N_5995,N_5047,N_5320);
and U5996 (N_5996,N_5324,N_5473);
or U5997 (N_5997,N_5488,N_5354);
nand U5998 (N_5998,N_5151,N_5306);
nand U5999 (N_5999,N_5078,N_5325);
or U6000 (N_6000,N_5880,N_5567);
nand U6001 (N_6001,N_5740,N_5841);
nor U6002 (N_6002,N_5758,N_5868);
or U6003 (N_6003,N_5619,N_5729);
nand U6004 (N_6004,N_5983,N_5789);
nor U6005 (N_6005,N_5562,N_5528);
or U6006 (N_6006,N_5664,N_5766);
or U6007 (N_6007,N_5920,N_5612);
or U6008 (N_6008,N_5725,N_5749);
nand U6009 (N_6009,N_5627,N_5691);
nand U6010 (N_6010,N_5713,N_5505);
nand U6011 (N_6011,N_5879,N_5600);
nand U6012 (N_6012,N_5863,N_5977);
or U6013 (N_6013,N_5836,N_5950);
xor U6014 (N_6014,N_5886,N_5685);
nand U6015 (N_6015,N_5915,N_5913);
and U6016 (N_6016,N_5774,N_5927);
nand U6017 (N_6017,N_5792,N_5830);
nor U6018 (N_6018,N_5502,N_5511);
xor U6019 (N_6019,N_5787,N_5862);
xnor U6020 (N_6020,N_5738,N_5723);
nand U6021 (N_6021,N_5904,N_5508);
nor U6022 (N_6022,N_5605,N_5721);
nor U6023 (N_6023,N_5663,N_5793);
xor U6024 (N_6024,N_5805,N_5907);
and U6025 (N_6025,N_5584,N_5959);
and U6026 (N_6026,N_5697,N_5719);
and U6027 (N_6027,N_5651,N_5641);
nand U6028 (N_6028,N_5896,N_5504);
and U6029 (N_6029,N_5763,N_5530);
and U6030 (N_6030,N_5799,N_5745);
nor U6031 (N_6031,N_5616,N_5784);
nand U6032 (N_6032,N_5773,N_5547);
or U6033 (N_6033,N_5996,N_5964);
or U6034 (N_6034,N_5992,N_5694);
xor U6035 (N_6035,N_5929,N_5515);
nor U6036 (N_6036,N_5974,N_5662);
nand U6037 (N_6037,N_5575,N_5620);
or U6038 (N_6038,N_5639,N_5644);
nand U6039 (N_6039,N_5760,N_5518);
xor U6040 (N_6040,N_5550,N_5585);
nor U6041 (N_6041,N_5642,N_5589);
xnor U6042 (N_6042,N_5901,N_5531);
nand U6043 (N_6043,N_5903,N_5768);
and U6044 (N_6044,N_5744,N_5970);
or U6045 (N_6045,N_5806,N_5791);
xor U6046 (N_6046,N_5577,N_5590);
or U6047 (N_6047,N_5971,N_5536);
or U6048 (N_6048,N_5917,N_5810);
xor U6049 (N_6049,N_5888,N_5638);
xnor U6050 (N_6050,N_5565,N_5637);
xnor U6051 (N_6051,N_5512,N_5724);
xor U6052 (N_6052,N_5846,N_5981);
or U6053 (N_6053,N_5842,N_5626);
or U6054 (N_6054,N_5849,N_5594);
nor U6055 (N_6055,N_5803,N_5614);
or U6056 (N_6056,N_5876,N_5720);
or U6057 (N_6057,N_5683,N_5670);
nor U6058 (N_6058,N_5543,N_5899);
or U6059 (N_6059,N_5608,N_5801);
nand U6060 (N_6060,N_5598,N_5742);
and U6061 (N_6061,N_5561,N_5857);
and U6062 (N_6062,N_5672,N_5759);
nor U6063 (N_6063,N_5905,N_5615);
nor U6064 (N_6064,N_5835,N_5556);
nand U6065 (N_6065,N_5624,N_5999);
xnor U6066 (N_6066,N_5889,N_5623);
or U6067 (N_6067,N_5555,N_5667);
xnor U6068 (N_6068,N_5731,N_5786);
nor U6069 (N_6069,N_5957,N_5963);
or U6070 (N_6070,N_5815,N_5647);
or U6071 (N_6071,N_5581,N_5973);
or U6072 (N_6072,N_5937,N_5859);
or U6073 (N_6073,N_5928,N_5912);
xnor U6074 (N_6074,N_5794,N_5750);
or U6075 (N_6075,N_5501,N_5798);
or U6076 (N_6076,N_5826,N_5610);
nand U6077 (N_6077,N_5533,N_5892);
xor U6078 (N_6078,N_5700,N_5780);
and U6079 (N_6079,N_5711,N_5781);
nand U6080 (N_6080,N_5761,N_5715);
nand U6081 (N_6081,N_5945,N_5884);
and U6082 (N_6082,N_5534,N_5748);
or U6083 (N_6083,N_5772,N_5571);
nand U6084 (N_6084,N_5537,N_5931);
and U6085 (N_6085,N_5676,N_5596);
nand U6086 (N_6086,N_5869,N_5628);
nand U6087 (N_6087,N_5607,N_5510);
nand U6088 (N_6088,N_5703,N_5573);
nor U6089 (N_6089,N_5795,N_5958);
xnor U6090 (N_6090,N_5506,N_5895);
nand U6091 (N_6091,N_5737,N_5542);
or U6092 (N_6092,N_5707,N_5526);
nand U6093 (N_6093,N_5513,N_5746);
nand U6094 (N_6094,N_5943,N_5881);
nand U6095 (N_6095,N_5788,N_5669);
nand U6096 (N_6096,N_5661,N_5779);
nand U6097 (N_6097,N_5591,N_5821);
xor U6098 (N_6098,N_5986,N_5960);
nor U6099 (N_6099,N_5712,N_5932);
and U6100 (N_6100,N_5710,N_5617);
xnor U6101 (N_6101,N_5674,N_5718);
nor U6102 (N_6102,N_5717,N_5618);
nand U6103 (N_6103,N_5601,N_5633);
xnor U6104 (N_6104,N_5613,N_5546);
and U6105 (N_6105,N_5563,N_5878);
nor U6106 (N_6106,N_5611,N_5539);
xor U6107 (N_6107,N_5574,N_5853);
xor U6108 (N_6108,N_5517,N_5681);
nand U6109 (N_6109,N_5656,N_5893);
xor U6110 (N_6110,N_5756,N_5762);
nor U6111 (N_6111,N_5521,N_5906);
nor U6112 (N_6112,N_5509,N_5910);
xnor U6113 (N_6113,N_5993,N_5566);
and U6114 (N_6114,N_5856,N_5606);
xnor U6115 (N_6115,N_5705,N_5765);
xnor U6116 (N_6116,N_5934,N_5666);
nor U6117 (N_6117,N_5679,N_5660);
or U6118 (N_6118,N_5771,N_5914);
and U6119 (N_6119,N_5630,N_5682);
nor U6120 (N_6120,N_5854,N_5948);
xnor U6121 (N_6121,N_5877,N_5852);
xnor U6122 (N_6122,N_5688,N_5797);
or U6123 (N_6123,N_5671,N_5597);
nand U6124 (N_6124,N_5757,N_5800);
xor U6125 (N_6125,N_5743,N_5783);
or U6126 (N_6126,N_5535,N_5726);
xnor U6127 (N_6127,N_5538,N_5752);
or U6128 (N_6128,N_5603,N_5769);
or U6129 (N_6129,N_5940,N_5695);
nand U6130 (N_6130,N_5549,N_5673);
xnor U6131 (N_6131,N_5936,N_5790);
nand U6132 (N_6132,N_5902,N_5930);
or U6133 (N_6133,N_5754,N_5827);
nor U6134 (N_6134,N_5524,N_5976);
nand U6135 (N_6135,N_5557,N_5956);
and U6136 (N_6136,N_5954,N_5753);
and U6137 (N_6137,N_5997,N_5875);
and U6138 (N_6138,N_5885,N_5552);
xor U6139 (N_6139,N_5995,N_5592);
and U6140 (N_6140,N_5916,N_5657);
or U6141 (N_6141,N_5693,N_5829);
or U6142 (N_6142,N_5775,N_5838);
and U6143 (N_6143,N_5655,N_5944);
xnor U6144 (N_6144,N_5668,N_5541);
and U6145 (N_6145,N_5558,N_5734);
nor U6146 (N_6146,N_5599,N_5870);
xor U6147 (N_6147,N_5646,N_5825);
xor U6148 (N_6148,N_5687,N_5975);
xor U6149 (N_6149,N_5861,N_5527);
nor U6150 (N_6150,N_5858,N_5570);
nor U6151 (N_6151,N_5559,N_5516);
and U6152 (N_6152,N_5621,N_5820);
nand U6153 (N_6153,N_5982,N_5522);
nand U6154 (N_6154,N_5819,N_5658);
and U6155 (N_6155,N_5947,N_5921);
xnor U6156 (N_6156,N_5716,N_5987);
and U6157 (N_6157,N_5953,N_5698);
nor U6158 (N_6158,N_5696,N_5851);
nor U6159 (N_6159,N_5702,N_5985);
nand U6160 (N_6160,N_5923,N_5529);
xor U6161 (N_6161,N_5747,N_5919);
and U6162 (N_6162,N_5949,N_5785);
xor U6163 (N_6163,N_5514,N_5812);
nand U6164 (N_6164,N_5817,N_5816);
or U6165 (N_6165,N_5837,N_5586);
nor U6166 (N_6166,N_5689,N_5978);
nand U6167 (N_6167,N_5860,N_5545);
xnor U6168 (N_6168,N_5872,N_5935);
nor U6169 (N_6169,N_5652,N_5850);
or U6170 (N_6170,N_5796,N_5519);
nand U6171 (N_6171,N_5727,N_5969);
nor U6172 (N_6172,N_5828,N_5891);
nor U6173 (N_6173,N_5728,N_5952);
nand U6174 (N_6174,N_5972,N_5887);
nor U6175 (N_6175,N_5523,N_5831);
nor U6176 (N_6176,N_5569,N_5548);
nor U6177 (N_6177,N_5554,N_5640);
nand U6178 (N_6178,N_5532,N_5938);
nand U6179 (N_6179,N_5507,N_5553);
or U6180 (N_6180,N_5649,N_5629);
nand U6181 (N_6181,N_5968,N_5701);
nor U6182 (N_6182,N_5882,N_5874);
or U6183 (N_6183,N_5708,N_5848);
nor U6184 (N_6184,N_5873,N_5777);
or U6185 (N_6185,N_5578,N_5941);
nand U6186 (N_6186,N_5933,N_5813);
and U6187 (N_6187,N_5867,N_5951);
nand U6188 (N_6188,N_5855,N_5544);
xor U6189 (N_6189,N_5736,N_5994);
or U6190 (N_6190,N_5942,N_5751);
xor U6191 (N_6191,N_5843,N_5714);
nand U6192 (N_6192,N_5909,N_5755);
or U6193 (N_6193,N_5686,N_5706);
nand U6194 (N_6194,N_5840,N_5609);
and U6195 (N_6195,N_5834,N_5908);
nor U6196 (N_6196,N_5645,N_5864);
nand U6197 (N_6197,N_5582,N_5926);
and U6198 (N_6198,N_5764,N_5823);
nand U6199 (N_6199,N_5804,N_5551);
and U6200 (N_6200,N_5654,N_5814);
xor U6201 (N_6201,N_5739,N_5730);
and U6202 (N_6202,N_5900,N_5939);
nor U6203 (N_6203,N_5722,N_5579);
and U6204 (N_6204,N_5692,N_5809);
or U6205 (N_6205,N_5989,N_5776);
and U6206 (N_6206,N_5832,N_5980);
or U6207 (N_6207,N_5650,N_5807);
nand U6208 (N_6208,N_5699,N_5818);
or U6209 (N_6209,N_5955,N_5845);
xor U6210 (N_6210,N_5967,N_5979);
nand U6211 (N_6211,N_5500,N_5733);
xor U6212 (N_6212,N_5824,N_5593);
nand U6213 (N_6213,N_5580,N_5767);
xor U6214 (N_6214,N_5677,N_5588);
nor U6215 (N_6215,N_5890,N_5897);
nor U6216 (N_6216,N_5984,N_5924);
nor U6217 (N_6217,N_5675,N_5898);
xor U6218 (N_6218,N_5811,N_5961);
and U6219 (N_6219,N_5634,N_5839);
or U6220 (N_6220,N_5587,N_5732);
nand U6221 (N_6221,N_5922,N_5966);
xnor U6222 (N_6222,N_5871,N_5680);
and U6223 (N_6223,N_5648,N_5782);
nand U6224 (N_6224,N_5802,N_5659);
and U6225 (N_6225,N_5865,N_5990);
xnor U6226 (N_6226,N_5946,N_5709);
xor U6227 (N_6227,N_5525,N_5770);
nor U6228 (N_6228,N_5735,N_5503);
nand U6229 (N_6229,N_5690,N_5991);
xnor U6230 (N_6230,N_5583,N_5741);
and U6231 (N_6231,N_5520,N_5576);
nand U6232 (N_6232,N_5918,N_5883);
or U6233 (N_6233,N_5678,N_5622);
and U6234 (N_6234,N_5998,N_5778);
or U6235 (N_6235,N_5925,N_5540);
nor U6236 (N_6236,N_5847,N_5894);
or U6237 (N_6237,N_5822,N_5965);
xnor U6238 (N_6238,N_5962,N_5568);
and U6239 (N_6239,N_5602,N_5572);
and U6240 (N_6240,N_5564,N_5604);
or U6241 (N_6241,N_5833,N_5704);
nor U6242 (N_6242,N_5653,N_5684);
nand U6243 (N_6243,N_5643,N_5636);
xnor U6244 (N_6244,N_5665,N_5632);
nand U6245 (N_6245,N_5866,N_5595);
and U6246 (N_6246,N_5988,N_5631);
xnor U6247 (N_6247,N_5808,N_5844);
and U6248 (N_6248,N_5635,N_5560);
and U6249 (N_6249,N_5625,N_5911);
and U6250 (N_6250,N_5909,N_5544);
nor U6251 (N_6251,N_5762,N_5629);
and U6252 (N_6252,N_5652,N_5758);
nand U6253 (N_6253,N_5511,N_5687);
xor U6254 (N_6254,N_5642,N_5550);
nand U6255 (N_6255,N_5857,N_5624);
nand U6256 (N_6256,N_5707,N_5627);
or U6257 (N_6257,N_5762,N_5531);
nand U6258 (N_6258,N_5886,N_5894);
nand U6259 (N_6259,N_5673,N_5826);
or U6260 (N_6260,N_5898,N_5699);
nor U6261 (N_6261,N_5965,N_5732);
nor U6262 (N_6262,N_5726,N_5709);
and U6263 (N_6263,N_5777,N_5902);
or U6264 (N_6264,N_5669,N_5907);
nand U6265 (N_6265,N_5793,N_5664);
or U6266 (N_6266,N_5785,N_5559);
nor U6267 (N_6267,N_5563,N_5706);
nor U6268 (N_6268,N_5506,N_5878);
nor U6269 (N_6269,N_5850,N_5784);
nand U6270 (N_6270,N_5920,N_5592);
xor U6271 (N_6271,N_5851,N_5825);
and U6272 (N_6272,N_5801,N_5756);
nor U6273 (N_6273,N_5694,N_5749);
nor U6274 (N_6274,N_5961,N_5526);
nor U6275 (N_6275,N_5655,N_5605);
and U6276 (N_6276,N_5786,N_5670);
nor U6277 (N_6277,N_5812,N_5594);
xnor U6278 (N_6278,N_5624,N_5926);
nand U6279 (N_6279,N_5631,N_5994);
nand U6280 (N_6280,N_5759,N_5651);
and U6281 (N_6281,N_5565,N_5978);
or U6282 (N_6282,N_5621,N_5841);
nand U6283 (N_6283,N_5556,N_5963);
xnor U6284 (N_6284,N_5706,N_5752);
nand U6285 (N_6285,N_5770,N_5533);
xor U6286 (N_6286,N_5516,N_5568);
nor U6287 (N_6287,N_5548,N_5881);
xor U6288 (N_6288,N_5736,N_5815);
nor U6289 (N_6289,N_5673,N_5927);
and U6290 (N_6290,N_5557,N_5745);
and U6291 (N_6291,N_5618,N_5755);
nand U6292 (N_6292,N_5546,N_5821);
and U6293 (N_6293,N_5659,N_5655);
nor U6294 (N_6294,N_5714,N_5848);
nor U6295 (N_6295,N_5933,N_5565);
nand U6296 (N_6296,N_5585,N_5922);
or U6297 (N_6297,N_5628,N_5796);
xnor U6298 (N_6298,N_5872,N_5885);
xor U6299 (N_6299,N_5858,N_5975);
nor U6300 (N_6300,N_5940,N_5964);
or U6301 (N_6301,N_5557,N_5650);
nor U6302 (N_6302,N_5870,N_5887);
or U6303 (N_6303,N_5862,N_5931);
nor U6304 (N_6304,N_5999,N_5914);
xnor U6305 (N_6305,N_5808,N_5573);
nand U6306 (N_6306,N_5848,N_5876);
and U6307 (N_6307,N_5916,N_5700);
nor U6308 (N_6308,N_5917,N_5977);
or U6309 (N_6309,N_5671,N_5988);
or U6310 (N_6310,N_5641,N_5675);
nor U6311 (N_6311,N_5526,N_5519);
nand U6312 (N_6312,N_5905,N_5847);
nand U6313 (N_6313,N_5834,N_5849);
nand U6314 (N_6314,N_5540,N_5793);
nand U6315 (N_6315,N_5789,N_5692);
or U6316 (N_6316,N_5870,N_5794);
or U6317 (N_6317,N_5788,N_5931);
xor U6318 (N_6318,N_5976,N_5703);
xor U6319 (N_6319,N_5866,N_5579);
xor U6320 (N_6320,N_5567,N_5657);
nor U6321 (N_6321,N_5923,N_5871);
nand U6322 (N_6322,N_5544,N_5994);
nand U6323 (N_6323,N_5829,N_5933);
and U6324 (N_6324,N_5762,N_5827);
or U6325 (N_6325,N_5974,N_5825);
nand U6326 (N_6326,N_5789,N_5517);
nor U6327 (N_6327,N_5514,N_5620);
and U6328 (N_6328,N_5969,N_5548);
or U6329 (N_6329,N_5658,N_5611);
or U6330 (N_6330,N_5887,N_5912);
and U6331 (N_6331,N_5957,N_5509);
or U6332 (N_6332,N_5870,N_5792);
nand U6333 (N_6333,N_5810,N_5627);
or U6334 (N_6334,N_5561,N_5927);
or U6335 (N_6335,N_5582,N_5843);
nand U6336 (N_6336,N_5761,N_5552);
and U6337 (N_6337,N_5518,N_5818);
or U6338 (N_6338,N_5840,N_5839);
nor U6339 (N_6339,N_5652,N_5576);
nor U6340 (N_6340,N_5772,N_5856);
and U6341 (N_6341,N_5738,N_5857);
nor U6342 (N_6342,N_5834,N_5922);
xor U6343 (N_6343,N_5672,N_5904);
nand U6344 (N_6344,N_5571,N_5683);
nand U6345 (N_6345,N_5998,N_5930);
or U6346 (N_6346,N_5990,N_5996);
nor U6347 (N_6347,N_5746,N_5972);
and U6348 (N_6348,N_5657,N_5539);
and U6349 (N_6349,N_5518,N_5719);
and U6350 (N_6350,N_5594,N_5697);
or U6351 (N_6351,N_5998,N_5909);
nand U6352 (N_6352,N_5899,N_5833);
and U6353 (N_6353,N_5819,N_5773);
or U6354 (N_6354,N_5819,N_5991);
xnor U6355 (N_6355,N_5753,N_5739);
and U6356 (N_6356,N_5552,N_5591);
xor U6357 (N_6357,N_5557,N_5895);
xor U6358 (N_6358,N_5592,N_5898);
nor U6359 (N_6359,N_5712,N_5740);
xor U6360 (N_6360,N_5772,N_5949);
nand U6361 (N_6361,N_5570,N_5766);
nor U6362 (N_6362,N_5747,N_5778);
nor U6363 (N_6363,N_5998,N_5712);
and U6364 (N_6364,N_5639,N_5587);
or U6365 (N_6365,N_5943,N_5607);
xor U6366 (N_6366,N_5654,N_5951);
or U6367 (N_6367,N_5760,N_5660);
nand U6368 (N_6368,N_5605,N_5682);
xor U6369 (N_6369,N_5621,N_5712);
or U6370 (N_6370,N_5803,N_5510);
nor U6371 (N_6371,N_5891,N_5862);
and U6372 (N_6372,N_5583,N_5917);
nor U6373 (N_6373,N_5787,N_5633);
or U6374 (N_6374,N_5641,N_5576);
or U6375 (N_6375,N_5879,N_5960);
and U6376 (N_6376,N_5828,N_5526);
or U6377 (N_6377,N_5935,N_5899);
or U6378 (N_6378,N_5967,N_5655);
nor U6379 (N_6379,N_5640,N_5536);
xnor U6380 (N_6380,N_5914,N_5717);
xnor U6381 (N_6381,N_5783,N_5941);
or U6382 (N_6382,N_5762,N_5769);
xnor U6383 (N_6383,N_5607,N_5896);
nor U6384 (N_6384,N_5701,N_5510);
nand U6385 (N_6385,N_5588,N_5500);
or U6386 (N_6386,N_5798,N_5618);
xor U6387 (N_6387,N_5581,N_5982);
nor U6388 (N_6388,N_5713,N_5712);
nand U6389 (N_6389,N_5553,N_5583);
nand U6390 (N_6390,N_5760,N_5644);
or U6391 (N_6391,N_5627,N_5701);
xnor U6392 (N_6392,N_5771,N_5701);
and U6393 (N_6393,N_5974,N_5831);
nand U6394 (N_6394,N_5552,N_5777);
nand U6395 (N_6395,N_5840,N_5629);
xor U6396 (N_6396,N_5772,N_5925);
xnor U6397 (N_6397,N_5671,N_5689);
xor U6398 (N_6398,N_5621,N_5596);
and U6399 (N_6399,N_5768,N_5504);
nand U6400 (N_6400,N_5769,N_5699);
nor U6401 (N_6401,N_5889,N_5756);
nand U6402 (N_6402,N_5987,N_5581);
xnor U6403 (N_6403,N_5621,N_5653);
or U6404 (N_6404,N_5775,N_5948);
and U6405 (N_6405,N_5806,N_5813);
xor U6406 (N_6406,N_5606,N_5812);
nor U6407 (N_6407,N_5768,N_5721);
and U6408 (N_6408,N_5967,N_5502);
and U6409 (N_6409,N_5722,N_5885);
nor U6410 (N_6410,N_5919,N_5891);
or U6411 (N_6411,N_5654,N_5624);
nor U6412 (N_6412,N_5938,N_5906);
and U6413 (N_6413,N_5955,N_5777);
nor U6414 (N_6414,N_5607,N_5863);
xnor U6415 (N_6415,N_5872,N_5990);
xor U6416 (N_6416,N_5938,N_5840);
and U6417 (N_6417,N_5621,N_5969);
nor U6418 (N_6418,N_5913,N_5778);
nand U6419 (N_6419,N_5683,N_5856);
nor U6420 (N_6420,N_5542,N_5616);
and U6421 (N_6421,N_5732,N_5920);
or U6422 (N_6422,N_5734,N_5842);
nand U6423 (N_6423,N_5797,N_5591);
nand U6424 (N_6424,N_5990,N_5873);
or U6425 (N_6425,N_5606,N_5638);
nand U6426 (N_6426,N_5579,N_5837);
nor U6427 (N_6427,N_5656,N_5787);
and U6428 (N_6428,N_5898,N_5818);
nand U6429 (N_6429,N_5757,N_5615);
xor U6430 (N_6430,N_5976,N_5749);
xnor U6431 (N_6431,N_5983,N_5972);
or U6432 (N_6432,N_5707,N_5501);
and U6433 (N_6433,N_5638,N_5825);
and U6434 (N_6434,N_5808,N_5706);
xor U6435 (N_6435,N_5580,N_5822);
and U6436 (N_6436,N_5934,N_5920);
xnor U6437 (N_6437,N_5685,N_5560);
or U6438 (N_6438,N_5698,N_5540);
nor U6439 (N_6439,N_5715,N_5746);
xnor U6440 (N_6440,N_5907,N_5896);
xnor U6441 (N_6441,N_5864,N_5641);
xor U6442 (N_6442,N_5540,N_5638);
nor U6443 (N_6443,N_5986,N_5605);
xnor U6444 (N_6444,N_5998,N_5728);
xor U6445 (N_6445,N_5559,N_5839);
xnor U6446 (N_6446,N_5763,N_5789);
nor U6447 (N_6447,N_5517,N_5827);
and U6448 (N_6448,N_5747,N_5752);
nand U6449 (N_6449,N_5648,N_5925);
or U6450 (N_6450,N_5746,N_5636);
nand U6451 (N_6451,N_5575,N_5821);
nand U6452 (N_6452,N_5791,N_5708);
or U6453 (N_6453,N_5925,N_5727);
nor U6454 (N_6454,N_5707,N_5973);
xor U6455 (N_6455,N_5898,N_5822);
and U6456 (N_6456,N_5633,N_5793);
nor U6457 (N_6457,N_5751,N_5628);
nor U6458 (N_6458,N_5998,N_5870);
xor U6459 (N_6459,N_5542,N_5569);
xnor U6460 (N_6460,N_5531,N_5609);
nor U6461 (N_6461,N_5835,N_5932);
xor U6462 (N_6462,N_5797,N_5624);
nand U6463 (N_6463,N_5830,N_5921);
nand U6464 (N_6464,N_5844,N_5571);
nor U6465 (N_6465,N_5620,N_5863);
xnor U6466 (N_6466,N_5515,N_5879);
nor U6467 (N_6467,N_5631,N_5619);
nor U6468 (N_6468,N_5674,N_5738);
and U6469 (N_6469,N_5818,N_5963);
xor U6470 (N_6470,N_5845,N_5629);
nand U6471 (N_6471,N_5688,N_5791);
nor U6472 (N_6472,N_5769,N_5759);
or U6473 (N_6473,N_5814,N_5930);
xnor U6474 (N_6474,N_5862,N_5821);
or U6475 (N_6475,N_5749,N_5981);
xor U6476 (N_6476,N_5790,N_5928);
and U6477 (N_6477,N_5971,N_5760);
nand U6478 (N_6478,N_5903,N_5996);
xor U6479 (N_6479,N_5893,N_5992);
and U6480 (N_6480,N_5543,N_5592);
or U6481 (N_6481,N_5580,N_5758);
and U6482 (N_6482,N_5616,N_5954);
and U6483 (N_6483,N_5908,N_5609);
or U6484 (N_6484,N_5529,N_5928);
or U6485 (N_6485,N_5634,N_5972);
and U6486 (N_6486,N_5917,N_5811);
or U6487 (N_6487,N_5909,N_5637);
xor U6488 (N_6488,N_5863,N_5749);
and U6489 (N_6489,N_5693,N_5767);
nor U6490 (N_6490,N_5886,N_5630);
nor U6491 (N_6491,N_5869,N_5890);
or U6492 (N_6492,N_5694,N_5542);
or U6493 (N_6493,N_5651,N_5997);
and U6494 (N_6494,N_5566,N_5750);
xor U6495 (N_6495,N_5984,N_5640);
nand U6496 (N_6496,N_5604,N_5828);
nor U6497 (N_6497,N_5898,N_5998);
nor U6498 (N_6498,N_5997,N_5619);
xnor U6499 (N_6499,N_5503,N_5886);
xnor U6500 (N_6500,N_6481,N_6022);
nor U6501 (N_6501,N_6447,N_6129);
or U6502 (N_6502,N_6315,N_6291);
nor U6503 (N_6503,N_6024,N_6175);
nand U6504 (N_6504,N_6397,N_6245);
and U6505 (N_6505,N_6444,N_6302);
and U6506 (N_6506,N_6325,N_6206);
nand U6507 (N_6507,N_6450,N_6027);
nand U6508 (N_6508,N_6280,N_6340);
or U6509 (N_6509,N_6037,N_6352);
nand U6510 (N_6510,N_6294,N_6219);
and U6511 (N_6511,N_6035,N_6462);
nand U6512 (N_6512,N_6139,N_6162);
xnor U6513 (N_6513,N_6008,N_6056);
nor U6514 (N_6514,N_6090,N_6190);
xor U6515 (N_6515,N_6395,N_6229);
or U6516 (N_6516,N_6073,N_6279);
nand U6517 (N_6517,N_6427,N_6100);
and U6518 (N_6518,N_6307,N_6230);
and U6519 (N_6519,N_6041,N_6042);
nor U6520 (N_6520,N_6211,N_6263);
nand U6521 (N_6521,N_6109,N_6240);
nor U6522 (N_6522,N_6417,N_6493);
nand U6523 (N_6523,N_6087,N_6184);
and U6524 (N_6524,N_6030,N_6265);
and U6525 (N_6525,N_6028,N_6440);
and U6526 (N_6526,N_6078,N_6418);
nand U6527 (N_6527,N_6074,N_6264);
nand U6528 (N_6528,N_6198,N_6277);
or U6529 (N_6529,N_6303,N_6257);
nor U6530 (N_6530,N_6285,N_6068);
xnor U6531 (N_6531,N_6466,N_6009);
nand U6532 (N_6532,N_6490,N_6498);
nand U6533 (N_6533,N_6351,N_6367);
xnor U6534 (N_6534,N_6083,N_6318);
and U6535 (N_6535,N_6428,N_6054);
xnor U6536 (N_6536,N_6414,N_6251);
nand U6537 (N_6537,N_6301,N_6416);
xnor U6538 (N_6538,N_6284,N_6254);
xnor U6539 (N_6539,N_6298,N_6120);
nor U6540 (N_6540,N_6225,N_6415);
and U6541 (N_6541,N_6411,N_6306);
xor U6542 (N_6542,N_6084,N_6443);
or U6543 (N_6543,N_6072,N_6448);
or U6544 (N_6544,N_6386,N_6153);
or U6545 (N_6545,N_6218,N_6259);
nor U6546 (N_6546,N_6317,N_6452);
or U6547 (N_6547,N_6193,N_6321);
and U6548 (N_6548,N_6131,N_6207);
and U6549 (N_6549,N_6112,N_6402);
and U6550 (N_6550,N_6123,N_6365);
xnor U6551 (N_6551,N_6103,N_6373);
nor U6552 (N_6552,N_6154,N_6220);
nand U6553 (N_6553,N_6043,N_6347);
nor U6554 (N_6554,N_6449,N_6314);
xnor U6555 (N_6555,N_6460,N_6216);
nand U6556 (N_6556,N_6354,N_6065);
nand U6557 (N_6557,N_6194,N_6126);
nand U6558 (N_6558,N_6172,N_6155);
nand U6559 (N_6559,N_6250,N_6375);
or U6560 (N_6560,N_6470,N_6342);
xor U6561 (N_6561,N_6274,N_6086);
or U6562 (N_6562,N_6483,N_6010);
or U6563 (N_6563,N_6262,N_6080);
nand U6564 (N_6564,N_6069,N_6442);
nand U6565 (N_6565,N_6282,N_6001);
nand U6566 (N_6566,N_6143,N_6370);
or U6567 (N_6567,N_6478,N_6094);
or U6568 (N_6568,N_6473,N_6164);
and U6569 (N_6569,N_6401,N_6376);
nor U6570 (N_6570,N_6324,N_6025);
or U6571 (N_6571,N_6379,N_6005);
and U6572 (N_6572,N_6296,N_6289);
and U6573 (N_6573,N_6276,N_6359);
or U6574 (N_6574,N_6149,N_6432);
nand U6575 (N_6575,N_6079,N_6044);
and U6576 (N_6576,N_6369,N_6075);
or U6577 (N_6577,N_6286,N_6210);
nand U6578 (N_6578,N_6145,N_6396);
and U6579 (N_6579,N_6170,N_6406);
xor U6580 (N_6580,N_6261,N_6186);
xor U6581 (N_6581,N_6290,N_6297);
nor U6582 (N_6582,N_6492,N_6016);
xor U6583 (N_6583,N_6469,N_6408);
nand U6584 (N_6584,N_6021,N_6039);
nand U6585 (N_6585,N_6144,N_6424);
and U6586 (N_6586,N_6268,N_6475);
and U6587 (N_6587,N_6082,N_6322);
or U6588 (N_6588,N_6288,N_6337);
xor U6589 (N_6589,N_6356,N_6157);
and U6590 (N_6590,N_6111,N_6439);
or U6591 (N_6591,N_6343,N_6384);
nor U6592 (N_6592,N_6203,N_6063);
or U6593 (N_6593,N_6032,N_6390);
nor U6594 (N_6594,N_6057,N_6147);
nand U6595 (N_6595,N_6105,N_6255);
or U6596 (N_6596,N_6436,N_6477);
or U6597 (N_6597,N_6004,N_6256);
nand U6598 (N_6598,N_6106,N_6361);
or U6599 (N_6599,N_6031,N_6467);
and U6600 (N_6600,N_6199,N_6388);
or U6601 (N_6601,N_6096,N_6422);
or U6602 (N_6602,N_6383,N_6161);
xnor U6603 (N_6603,N_6434,N_6104);
nand U6604 (N_6604,N_6189,N_6445);
nand U6605 (N_6605,N_6013,N_6474);
xor U6606 (N_6606,N_6341,N_6171);
xor U6607 (N_6607,N_6130,N_6468);
and U6608 (N_6608,N_6209,N_6159);
nor U6609 (N_6609,N_6231,N_6266);
nor U6610 (N_6610,N_6249,N_6348);
nand U6611 (N_6611,N_6399,N_6196);
xnor U6612 (N_6612,N_6300,N_6067);
xnor U6613 (N_6613,N_6116,N_6237);
nor U6614 (N_6614,N_6465,N_6000);
and U6615 (N_6615,N_6410,N_6260);
nand U6616 (N_6616,N_6246,N_6125);
xor U6617 (N_6617,N_6034,N_6227);
xor U6618 (N_6618,N_6364,N_6185);
xor U6619 (N_6619,N_6305,N_6456);
or U6620 (N_6620,N_6393,N_6309);
xnor U6621 (N_6621,N_6201,N_6479);
xor U6622 (N_6622,N_6350,N_6114);
nor U6623 (N_6623,N_6033,N_6187);
nand U6624 (N_6624,N_6156,N_6191);
xor U6625 (N_6625,N_6316,N_6213);
and U6626 (N_6626,N_6150,N_6311);
xnor U6627 (N_6627,N_6463,N_6328);
nor U6628 (N_6628,N_6183,N_6215);
nor U6629 (N_6629,N_6258,N_6046);
and U6630 (N_6630,N_6006,N_6205);
and U6631 (N_6631,N_6482,N_6308);
xnor U6632 (N_6632,N_6239,N_6121);
or U6633 (N_6633,N_6387,N_6148);
nand U6634 (N_6634,N_6243,N_6458);
nand U6635 (N_6635,N_6115,N_6441);
nor U6636 (N_6636,N_6292,N_6029);
xor U6637 (N_6637,N_6212,N_6461);
nor U6638 (N_6638,N_6053,N_6488);
nand U6639 (N_6639,N_6208,N_6197);
nor U6640 (N_6640,N_6494,N_6093);
nand U6641 (N_6641,N_6108,N_6007);
xor U6642 (N_6642,N_6122,N_6398);
and U6643 (N_6643,N_6329,N_6242);
xnor U6644 (N_6644,N_6140,N_6099);
or U6645 (N_6645,N_6451,N_6052);
xor U6646 (N_6646,N_6113,N_6381);
xor U6647 (N_6647,N_6182,N_6454);
nor U6648 (N_6648,N_6012,N_6232);
nand U6649 (N_6649,N_6163,N_6038);
nand U6650 (N_6650,N_6382,N_6214);
and U6651 (N_6651,N_6345,N_6374);
or U6652 (N_6652,N_6421,N_6331);
nor U6653 (N_6653,N_6177,N_6489);
or U6654 (N_6654,N_6088,N_6176);
nor U6655 (N_6655,N_6158,N_6195);
or U6656 (N_6656,N_6048,N_6433);
or U6657 (N_6657,N_6491,N_6287);
xor U6658 (N_6658,N_6378,N_6138);
or U6659 (N_6659,N_6313,N_6366);
and U6660 (N_6660,N_6050,N_6036);
xor U6661 (N_6661,N_6102,N_6179);
nor U6662 (N_6662,N_6485,N_6059);
and U6663 (N_6663,N_6327,N_6455);
or U6664 (N_6664,N_6495,N_6134);
xnor U6665 (N_6665,N_6235,N_6497);
and U6666 (N_6666,N_6055,N_6430);
and U6667 (N_6667,N_6101,N_6281);
nor U6668 (N_6668,N_6368,N_6459);
and U6669 (N_6669,N_6472,N_6045);
nor U6670 (N_6670,N_6070,N_6110);
nor U6671 (N_6671,N_6226,N_6200);
or U6672 (N_6672,N_6423,N_6233);
xnor U6673 (N_6673,N_6480,N_6336);
and U6674 (N_6674,N_6295,N_6160);
nor U6675 (N_6675,N_6496,N_6169);
nand U6676 (N_6676,N_6426,N_6064);
or U6677 (N_6677,N_6438,N_6071);
xnor U6678 (N_6678,N_6133,N_6435);
or U6679 (N_6679,N_6419,N_6174);
nand U6680 (N_6680,N_6124,N_6471);
or U6681 (N_6681,N_6453,N_6339);
xnor U6682 (N_6682,N_6061,N_6077);
or U6683 (N_6683,N_6377,N_6275);
nand U6684 (N_6684,N_6349,N_6412);
nand U6685 (N_6685,N_6446,N_6253);
xnor U6686 (N_6686,N_6023,N_6142);
and U6687 (N_6687,N_6118,N_6017);
nor U6688 (N_6688,N_6323,N_6425);
or U6689 (N_6689,N_6135,N_6484);
or U6690 (N_6690,N_6335,N_6362);
nand U6691 (N_6691,N_6404,N_6270);
xnor U6692 (N_6692,N_6132,N_6310);
nor U6693 (N_6693,N_6003,N_6181);
nand U6694 (N_6694,N_6420,N_6476);
nand U6695 (N_6695,N_6391,N_6049);
nor U6696 (N_6696,N_6092,N_6019);
and U6697 (N_6697,N_6091,N_6018);
xor U6698 (N_6698,N_6217,N_6358);
and U6699 (N_6699,N_6241,N_6269);
or U6700 (N_6700,N_6372,N_6026);
or U6701 (N_6701,N_6293,N_6167);
or U6702 (N_6702,N_6014,N_6283);
nand U6703 (N_6703,N_6338,N_6221);
xnor U6704 (N_6704,N_6299,N_6085);
nand U6705 (N_6705,N_6344,N_6141);
nor U6706 (N_6706,N_6389,N_6152);
or U6707 (N_6707,N_6178,N_6247);
xnor U6708 (N_6708,N_6151,N_6371);
nor U6709 (N_6709,N_6271,N_6180);
nand U6710 (N_6710,N_6188,N_6499);
and U6711 (N_6711,N_6400,N_6058);
nor U6712 (N_6712,N_6431,N_6204);
xor U6713 (N_6713,N_6363,N_6011);
or U6714 (N_6714,N_6236,N_6248);
xor U6715 (N_6715,N_6332,N_6403);
and U6716 (N_6716,N_6409,N_6334);
nand U6717 (N_6717,N_6128,N_6165);
nor U6718 (N_6718,N_6224,N_6238);
and U6719 (N_6719,N_6355,N_6272);
xor U6720 (N_6720,N_6346,N_6136);
xor U6721 (N_6721,N_6252,N_6486);
nand U6722 (N_6722,N_6360,N_6223);
nor U6723 (N_6723,N_6320,N_6089);
nor U6724 (N_6724,N_6312,N_6107);
or U6725 (N_6725,N_6146,N_6405);
or U6726 (N_6726,N_6040,N_6385);
nand U6727 (N_6727,N_6117,N_6051);
and U6728 (N_6728,N_6137,N_6166);
nand U6729 (N_6729,N_6394,N_6020);
and U6730 (N_6730,N_6353,N_6076);
nor U6731 (N_6731,N_6487,N_6380);
and U6732 (N_6732,N_6097,N_6330);
xnor U6733 (N_6733,N_6168,N_6407);
xor U6734 (N_6734,N_6060,N_6457);
or U6735 (N_6735,N_6062,N_6437);
nand U6736 (N_6736,N_6228,N_6304);
and U6737 (N_6737,N_6047,N_6413);
xor U6738 (N_6738,N_6357,N_6002);
or U6739 (N_6739,N_6333,N_6267);
nand U6740 (N_6740,N_6081,N_6319);
or U6741 (N_6741,N_6202,N_6015);
or U6742 (N_6742,N_6244,N_6273);
nand U6743 (N_6743,N_6326,N_6119);
and U6744 (N_6744,N_6222,N_6192);
xnor U6745 (N_6745,N_6127,N_6066);
xnor U6746 (N_6746,N_6392,N_6234);
xor U6747 (N_6747,N_6464,N_6095);
xor U6748 (N_6748,N_6173,N_6429);
nor U6749 (N_6749,N_6098,N_6278);
and U6750 (N_6750,N_6433,N_6396);
nand U6751 (N_6751,N_6046,N_6311);
xor U6752 (N_6752,N_6085,N_6231);
nor U6753 (N_6753,N_6447,N_6105);
and U6754 (N_6754,N_6418,N_6285);
xnor U6755 (N_6755,N_6384,N_6465);
xor U6756 (N_6756,N_6473,N_6097);
nor U6757 (N_6757,N_6118,N_6176);
xnor U6758 (N_6758,N_6469,N_6441);
xor U6759 (N_6759,N_6326,N_6179);
and U6760 (N_6760,N_6356,N_6203);
xor U6761 (N_6761,N_6141,N_6171);
xnor U6762 (N_6762,N_6173,N_6387);
xor U6763 (N_6763,N_6246,N_6047);
nand U6764 (N_6764,N_6247,N_6276);
nor U6765 (N_6765,N_6199,N_6092);
nor U6766 (N_6766,N_6186,N_6367);
and U6767 (N_6767,N_6471,N_6247);
and U6768 (N_6768,N_6358,N_6064);
nand U6769 (N_6769,N_6239,N_6425);
xor U6770 (N_6770,N_6091,N_6457);
nor U6771 (N_6771,N_6235,N_6450);
xnor U6772 (N_6772,N_6437,N_6360);
nor U6773 (N_6773,N_6013,N_6393);
xor U6774 (N_6774,N_6017,N_6302);
nor U6775 (N_6775,N_6341,N_6137);
and U6776 (N_6776,N_6414,N_6283);
nor U6777 (N_6777,N_6484,N_6321);
nor U6778 (N_6778,N_6189,N_6276);
xor U6779 (N_6779,N_6348,N_6407);
xnor U6780 (N_6780,N_6263,N_6410);
or U6781 (N_6781,N_6090,N_6357);
xnor U6782 (N_6782,N_6036,N_6346);
and U6783 (N_6783,N_6130,N_6234);
or U6784 (N_6784,N_6439,N_6091);
nor U6785 (N_6785,N_6430,N_6159);
nand U6786 (N_6786,N_6355,N_6070);
and U6787 (N_6787,N_6145,N_6402);
xor U6788 (N_6788,N_6448,N_6482);
or U6789 (N_6789,N_6042,N_6065);
or U6790 (N_6790,N_6167,N_6350);
xnor U6791 (N_6791,N_6138,N_6104);
nand U6792 (N_6792,N_6380,N_6400);
xnor U6793 (N_6793,N_6266,N_6211);
and U6794 (N_6794,N_6078,N_6101);
or U6795 (N_6795,N_6207,N_6046);
xnor U6796 (N_6796,N_6338,N_6294);
nand U6797 (N_6797,N_6124,N_6385);
nor U6798 (N_6798,N_6268,N_6403);
xnor U6799 (N_6799,N_6074,N_6212);
or U6800 (N_6800,N_6169,N_6446);
nand U6801 (N_6801,N_6245,N_6435);
xnor U6802 (N_6802,N_6471,N_6061);
nand U6803 (N_6803,N_6474,N_6020);
nand U6804 (N_6804,N_6291,N_6157);
or U6805 (N_6805,N_6052,N_6338);
and U6806 (N_6806,N_6496,N_6274);
nand U6807 (N_6807,N_6401,N_6175);
and U6808 (N_6808,N_6073,N_6438);
and U6809 (N_6809,N_6285,N_6190);
nand U6810 (N_6810,N_6284,N_6074);
nand U6811 (N_6811,N_6198,N_6145);
xnor U6812 (N_6812,N_6257,N_6481);
xnor U6813 (N_6813,N_6213,N_6201);
or U6814 (N_6814,N_6209,N_6119);
nand U6815 (N_6815,N_6159,N_6314);
or U6816 (N_6816,N_6201,N_6341);
nand U6817 (N_6817,N_6114,N_6437);
nand U6818 (N_6818,N_6047,N_6022);
nand U6819 (N_6819,N_6278,N_6450);
nor U6820 (N_6820,N_6478,N_6056);
nand U6821 (N_6821,N_6037,N_6460);
xor U6822 (N_6822,N_6457,N_6365);
nor U6823 (N_6823,N_6318,N_6191);
nand U6824 (N_6824,N_6069,N_6372);
or U6825 (N_6825,N_6420,N_6396);
or U6826 (N_6826,N_6358,N_6114);
and U6827 (N_6827,N_6180,N_6011);
nor U6828 (N_6828,N_6072,N_6475);
xnor U6829 (N_6829,N_6006,N_6156);
or U6830 (N_6830,N_6081,N_6393);
nand U6831 (N_6831,N_6309,N_6446);
nand U6832 (N_6832,N_6051,N_6294);
nand U6833 (N_6833,N_6489,N_6304);
nor U6834 (N_6834,N_6316,N_6403);
nor U6835 (N_6835,N_6034,N_6308);
or U6836 (N_6836,N_6465,N_6325);
and U6837 (N_6837,N_6140,N_6400);
nand U6838 (N_6838,N_6328,N_6252);
xor U6839 (N_6839,N_6035,N_6457);
nor U6840 (N_6840,N_6097,N_6303);
nor U6841 (N_6841,N_6479,N_6003);
and U6842 (N_6842,N_6484,N_6030);
nor U6843 (N_6843,N_6471,N_6015);
xor U6844 (N_6844,N_6197,N_6312);
nand U6845 (N_6845,N_6472,N_6066);
or U6846 (N_6846,N_6234,N_6384);
xnor U6847 (N_6847,N_6435,N_6466);
xnor U6848 (N_6848,N_6404,N_6127);
xnor U6849 (N_6849,N_6338,N_6106);
or U6850 (N_6850,N_6202,N_6398);
or U6851 (N_6851,N_6155,N_6270);
or U6852 (N_6852,N_6045,N_6077);
nor U6853 (N_6853,N_6080,N_6137);
xor U6854 (N_6854,N_6486,N_6400);
or U6855 (N_6855,N_6363,N_6499);
or U6856 (N_6856,N_6252,N_6082);
xnor U6857 (N_6857,N_6212,N_6442);
and U6858 (N_6858,N_6058,N_6242);
nor U6859 (N_6859,N_6177,N_6455);
nor U6860 (N_6860,N_6463,N_6379);
nand U6861 (N_6861,N_6455,N_6281);
nand U6862 (N_6862,N_6491,N_6183);
nand U6863 (N_6863,N_6375,N_6045);
nand U6864 (N_6864,N_6039,N_6343);
nor U6865 (N_6865,N_6449,N_6184);
or U6866 (N_6866,N_6235,N_6111);
nor U6867 (N_6867,N_6361,N_6412);
and U6868 (N_6868,N_6066,N_6123);
and U6869 (N_6869,N_6459,N_6059);
or U6870 (N_6870,N_6407,N_6419);
and U6871 (N_6871,N_6455,N_6318);
nor U6872 (N_6872,N_6461,N_6002);
nor U6873 (N_6873,N_6021,N_6462);
nor U6874 (N_6874,N_6283,N_6304);
xnor U6875 (N_6875,N_6109,N_6257);
xnor U6876 (N_6876,N_6311,N_6168);
xor U6877 (N_6877,N_6144,N_6126);
or U6878 (N_6878,N_6250,N_6153);
and U6879 (N_6879,N_6250,N_6351);
and U6880 (N_6880,N_6203,N_6372);
nand U6881 (N_6881,N_6441,N_6206);
nand U6882 (N_6882,N_6104,N_6287);
nor U6883 (N_6883,N_6028,N_6293);
nor U6884 (N_6884,N_6475,N_6371);
nand U6885 (N_6885,N_6363,N_6260);
nor U6886 (N_6886,N_6489,N_6383);
nand U6887 (N_6887,N_6160,N_6102);
and U6888 (N_6888,N_6459,N_6043);
nor U6889 (N_6889,N_6252,N_6231);
nand U6890 (N_6890,N_6087,N_6136);
nand U6891 (N_6891,N_6476,N_6472);
xor U6892 (N_6892,N_6424,N_6302);
or U6893 (N_6893,N_6110,N_6378);
nor U6894 (N_6894,N_6012,N_6403);
or U6895 (N_6895,N_6441,N_6240);
and U6896 (N_6896,N_6272,N_6196);
or U6897 (N_6897,N_6348,N_6144);
nor U6898 (N_6898,N_6465,N_6048);
or U6899 (N_6899,N_6363,N_6299);
xor U6900 (N_6900,N_6185,N_6444);
nand U6901 (N_6901,N_6236,N_6225);
xor U6902 (N_6902,N_6470,N_6482);
nand U6903 (N_6903,N_6228,N_6439);
nor U6904 (N_6904,N_6142,N_6258);
xor U6905 (N_6905,N_6076,N_6305);
nand U6906 (N_6906,N_6294,N_6046);
nor U6907 (N_6907,N_6148,N_6466);
nand U6908 (N_6908,N_6300,N_6164);
xnor U6909 (N_6909,N_6099,N_6338);
and U6910 (N_6910,N_6012,N_6089);
xnor U6911 (N_6911,N_6044,N_6187);
nor U6912 (N_6912,N_6003,N_6016);
nand U6913 (N_6913,N_6240,N_6406);
or U6914 (N_6914,N_6128,N_6223);
and U6915 (N_6915,N_6065,N_6348);
nand U6916 (N_6916,N_6407,N_6268);
nor U6917 (N_6917,N_6195,N_6456);
or U6918 (N_6918,N_6360,N_6034);
nor U6919 (N_6919,N_6269,N_6476);
and U6920 (N_6920,N_6395,N_6252);
or U6921 (N_6921,N_6221,N_6446);
xnor U6922 (N_6922,N_6468,N_6470);
or U6923 (N_6923,N_6434,N_6111);
xnor U6924 (N_6924,N_6252,N_6124);
and U6925 (N_6925,N_6218,N_6327);
xor U6926 (N_6926,N_6421,N_6197);
xor U6927 (N_6927,N_6201,N_6158);
xnor U6928 (N_6928,N_6154,N_6047);
nor U6929 (N_6929,N_6115,N_6474);
xnor U6930 (N_6930,N_6302,N_6383);
nand U6931 (N_6931,N_6116,N_6194);
and U6932 (N_6932,N_6146,N_6329);
or U6933 (N_6933,N_6451,N_6148);
and U6934 (N_6934,N_6232,N_6024);
nand U6935 (N_6935,N_6302,N_6021);
nand U6936 (N_6936,N_6156,N_6209);
and U6937 (N_6937,N_6481,N_6287);
nor U6938 (N_6938,N_6097,N_6140);
nor U6939 (N_6939,N_6380,N_6368);
xor U6940 (N_6940,N_6313,N_6265);
nor U6941 (N_6941,N_6329,N_6454);
or U6942 (N_6942,N_6383,N_6320);
nor U6943 (N_6943,N_6458,N_6004);
nor U6944 (N_6944,N_6056,N_6229);
nand U6945 (N_6945,N_6385,N_6208);
and U6946 (N_6946,N_6489,N_6361);
nor U6947 (N_6947,N_6008,N_6137);
nand U6948 (N_6948,N_6087,N_6231);
and U6949 (N_6949,N_6324,N_6033);
nand U6950 (N_6950,N_6156,N_6405);
nor U6951 (N_6951,N_6093,N_6318);
and U6952 (N_6952,N_6250,N_6437);
xnor U6953 (N_6953,N_6271,N_6119);
nor U6954 (N_6954,N_6087,N_6203);
or U6955 (N_6955,N_6332,N_6033);
nor U6956 (N_6956,N_6400,N_6454);
nor U6957 (N_6957,N_6205,N_6304);
or U6958 (N_6958,N_6417,N_6445);
and U6959 (N_6959,N_6139,N_6187);
xor U6960 (N_6960,N_6438,N_6007);
nor U6961 (N_6961,N_6104,N_6368);
and U6962 (N_6962,N_6126,N_6470);
xnor U6963 (N_6963,N_6068,N_6096);
and U6964 (N_6964,N_6123,N_6038);
nand U6965 (N_6965,N_6054,N_6490);
nor U6966 (N_6966,N_6362,N_6075);
or U6967 (N_6967,N_6498,N_6313);
nand U6968 (N_6968,N_6463,N_6397);
nor U6969 (N_6969,N_6372,N_6303);
nor U6970 (N_6970,N_6364,N_6245);
nor U6971 (N_6971,N_6476,N_6455);
or U6972 (N_6972,N_6045,N_6455);
and U6973 (N_6973,N_6210,N_6120);
nor U6974 (N_6974,N_6190,N_6097);
xnor U6975 (N_6975,N_6205,N_6452);
or U6976 (N_6976,N_6277,N_6302);
and U6977 (N_6977,N_6201,N_6069);
and U6978 (N_6978,N_6370,N_6248);
and U6979 (N_6979,N_6398,N_6334);
and U6980 (N_6980,N_6444,N_6167);
xnor U6981 (N_6981,N_6466,N_6499);
and U6982 (N_6982,N_6381,N_6168);
xor U6983 (N_6983,N_6440,N_6383);
xor U6984 (N_6984,N_6355,N_6482);
nor U6985 (N_6985,N_6013,N_6001);
and U6986 (N_6986,N_6255,N_6186);
xor U6987 (N_6987,N_6019,N_6455);
or U6988 (N_6988,N_6071,N_6440);
or U6989 (N_6989,N_6373,N_6324);
nor U6990 (N_6990,N_6436,N_6023);
nand U6991 (N_6991,N_6126,N_6036);
nor U6992 (N_6992,N_6487,N_6307);
nand U6993 (N_6993,N_6429,N_6367);
xnor U6994 (N_6994,N_6049,N_6310);
and U6995 (N_6995,N_6245,N_6484);
xnor U6996 (N_6996,N_6312,N_6313);
and U6997 (N_6997,N_6035,N_6175);
xnor U6998 (N_6998,N_6241,N_6155);
nand U6999 (N_6999,N_6359,N_6123);
or U7000 (N_7000,N_6575,N_6656);
xnor U7001 (N_7001,N_6636,N_6865);
xnor U7002 (N_7002,N_6517,N_6763);
nand U7003 (N_7003,N_6782,N_6707);
nor U7004 (N_7004,N_6728,N_6740);
or U7005 (N_7005,N_6722,N_6886);
xnor U7006 (N_7006,N_6847,N_6798);
nand U7007 (N_7007,N_6818,N_6824);
or U7008 (N_7008,N_6972,N_6982);
nand U7009 (N_7009,N_6553,N_6927);
nand U7010 (N_7010,N_6540,N_6905);
and U7011 (N_7011,N_6993,N_6966);
xor U7012 (N_7012,N_6866,N_6817);
xnor U7013 (N_7013,N_6959,N_6533);
nor U7014 (N_7014,N_6608,N_6796);
xnor U7015 (N_7015,N_6916,N_6692);
xnor U7016 (N_7016,N_6820,N_6879);
nor U7017 (N_7017,N_6730,N_6781);
or U7018 (N_7018,N_6565,N_6822);
nand U7019 (N_7019,N_6543,N_6750);
xnor U7020 (N_7020,N_6881,N_6634);
nand U7021 (N_7021,N_6925,N_6623);
or U7022 (N_7022,N_6601,N_6518);
or U7023 (N_7023,N_6621,N_6978);
nand U7024 (N_7024,N_6742,N_6594);
nand U7025 (N_7025,N_6778,N_6811);
xnor U7026 (N_7026,N_6584,N_6838);
or U7027 (N_7027,N_6840,N_6851);
nor U7028 (N_7028,N_6668,N_6785);
and U7029 (N_7029,N_6902,N_6526);
nor U7030 (N_7030,N_6985,N_6967);
nor U7031 (N_7031,N_6821,N_6706);
nor U7032 (N_7032,N_6749,N_6952);
nor U7033 (N_7033,N_6609,N_6637);
nor U7034 (N_7034,N_6615,N_6994);
nor U7035 (N_7035,N_6729,N_6748);
and U7036 (N_7036,N_6950,N_6557);
and U7037 (N_7037,N_6956,N_6743);
nand U7038 (N_7038,N_6981,N_6772);
or U7039 (N_7039,N_6585,N_6857);
or U7040 (N_7040,N_6829,N_6936);
and U7041 (N_7041,N_6542,N_6566);
and U7042 (N_7042,N_6712,N_6669);
or U7043 (N_7043,N_6622,N_6509);
nor U7044 (N_7044,N_6777,N_6568);
nand U7045 (N_7045,N_6655,N_6776);
nand U7046 (N_7046,N_6976,N_6853);
xnor U7047 (N_7047,N_6702,N_6854);
nand U7048 (N_7048,N_6843,N_6582);
and U7049 (N_7049,N_6697,N_6979);
xor U7050 (N_7050,N_6567,N_6823);
nor U7051 (N_7051,N_6834,N_6643);
or U7052 (N_7052,N_6805,N_6904);
or U7053 (N_7053,N_6774,N_6974);
or U7054 (N_7054,N_6793,N_6635);
nor U7055 (N_7055,N_6684,N_6769);
nor U7056 (N_7056,N_6718,N_6593);
and U7057 (N_7057,N_6989,N_6650);
nor U7058 (N_7058,N_6986,N_6765);
and U7059 (N_7059,N_6987,N_6733);
xor U7060 (N_7060,N_6665,N_6912);
nand U7061 (N_7061,N_6771,N_6929);
nand U7062 (N_7062,N_6984,N_6558);
xor U7063 (N_7063,N_6563,N_6619);
nor U7064 (N_7064,N_6875,N_6794);
or U7065 (N_7065,N_6600,N_6858);
xor U7066 (N_7066,N_6973,N_6832);
nor U7067 (N_7067,N_6897,N_6835);
xor U7068 (N_7068,N_6685,N_6536);
xor U7069 (N_7069,N_6795,N_6638);
nand U7070 (N_7070,N_6999,N_6644);
nand U7071 (N_7071,N_6528,N_6519);
xnor U7072 (N_7072,N_6842,N_6539);
and U7073 (N_7073,N_6719,N_6696);
xor U7074 (N_7074,N_6887,N_6760);
and U7075 (N_7075,N_6864,N_6955);
nand U7076 (N_7076,N_6928,N_6764);
nor U7077 (N_7077,N_6627,N_6524);
nand U7078 (N_7078,N_6647,N_6918);
or U7079 (N_7079,N_6694,N_6991);
or U7080 (N_7080,N_6554,N_6537);
and U7081 (N_7081,N_6852,N_6888);
or U7082 (N_7082,N_6738,N_6522);
and U7083 (N_7083,N_6573,N_6525);
or U7084 (N_7084,N_6671,N_6680);
nor U7085 (N_7085,N_6597,N_6751);
and U7086 (N_7086,N_6731,N_6732);
and U7087 (N_7087,N_6812,N_6693);
and U7088 (N_7088,N_6552,N_6755);
nand U7089 (N_7089,N_6964,N_6859);
nand U7090 (N_7090,N_6534,N_6971);
xnor U7091 (N_7091,N_6523,N_6954);
or U7092 (N_7092,N_6577,N_6930);
nand U7093 (N_7093,N_6734,N_6583);
nor U7094 (N_7094,N_6633,N_6931);
and U7095 (N_7095,N_6687,N_6848);
xor U7096 (N_7096,N_6899,N_6963);
and U7097 (N_7097,N_6616,N_6695);
or U7098 (N_7098,N_6983,N_6675);
xor U7099 (N_7099,N_6937,N_6690);
xnor U7100 (N_7100,N_6970,N_6556);
nand U7101 (N_7101,N_6646,N_6890);
and U7102 (N_7102,N_6502,N_6574);
nor U7103 (N_7103,N_6758,N_6784);
xnor U7104 (N_7104,N_6614,N_6773);
xor U7105 (N_7105,N_6704,N_6658);
and U7106 (N_7106,N_6957,N_6513);
nand U7107 (N_7107,N_6648,N_6739);
nand U7108 (N_7108,N_6910,N_6882);
nand U7109 (N_7109,N_6746,N_6741);
xor U7110 (N_7110,N_6711,N_6977);
xnor U7111 (N_7111,N_6663,N_6560);
nor U7112 (N_7112,N_6913,N_6681);
nand U7113 (N_7113,N_6767,N_6571);
and U7114 (N_7114,N_6700,N_6612);
xnor U7115 (N_7115,N_6884,N_6603);
xnor U7116 (N_7116,N_6761,N_6724);
nand U7117 (N_7117,N_6723,N_6998);
or U7118 (N_7118,N_6786,N_6703);
xor U7119 (N_7119,N_6894,N_6649);
or U7120 (N_7120,N_6862,N_6896);
nand U7121 (N_7121,N_6673,N_6641);
xnor U7122 (N_7122,N_6968,N_6555);
xnor U7123 (N_7123,N_6944,N_6815);
xnor U7124 (N_7124,N_6576,N_6801);
nand U7125 (N_7125,N_6903,N_6992);
and U7126 (N_7126,N_6855,N_6961);
and U7127 (N_7127,N_6507,N_6578);
and U7128 (N_7128,N_6878,N_6744);
nand U7129 (N_7129,N_6779,N_6876);
or U7130 (N_7130,N_6503,N_6988);
and U7131 (N_7131,N_6531,N_6506);
or U7132 (N_7132,N_6813,N_6908);
nand U7133 (N_7133,N_6947,N_6591);
nor U7134 (N_7134,N_6893,N_6868);
nor U7135 (N_7135,N_6996,N_6883);
and U7136 (N_7136,N_6709,N_6735);
and U7137 (N_7137,N_6725,N_6624);
and U7138 (N_7138,N_6980,N_6892);
nand U7139 (N_7139,N_6901,N_6791);
or U7140 (N_7140,N_6639,N_6827);
and U7141 (N_7141,N_6550,N_6629);
and U7142 (N_7142,N_6599,N_6628);
nand U7143 (N_7143,N_6588,N_6547);
and U7144 (N_7144,N_6521,N_6872);
or U7145 (N_7145,N_6666,N_6686);
nand U7146 (N_7146,N_6911,N_6631);
or U7147 (N_7147,N_6877,N_6688);
nor U7148 (N_7148,N_6962,N_6787);
nand U7149 (N_7149,N_6714,N_6651);
and U7150 (N_7150,N_6825,N_6907);
and U7151 (N_7151,N_6505,N_6652);
and U7152 (N_7152,N_6933,N_6662);
xnor U7153 (N_7153,N_6932,N_6721);
or U7154 (N_7154,N_6800,N_6610);
or U7155 (N_7155,N_6831,N_6799);
and U7156 (N_7156,N_6653,N_6790);
or U7157 (N_7157,N_6898,N_6544);
nand U7158 (N_7158,N_6803,N_6500);
xor U7159 (N_7159,N_6511,N_6562);
nand U7160 (N_7160,N_6891,N_6846);
xnor U7161 (N_7161,N_6920,N_6736);
or U7162 (N_7162,N_6672,N_6532);
xnor U7163 (N_7163,N_6589,N_6924);
and U7164 (N_7164,N_6630,N_6515);
nand U7165 (N_7165,N_6661,N_6869);
nor U7166 (N_7166,N_6586,N_6807);
or U7167 (N_7167,N_6863,N_6889);
nand U7168 (N_7168,N_6770,N_6926);
xor U7169 (N_7169,N_6757,N_6683);
nor U7170 (N_7170,N_6581,N_6870);
nor U7171 (N_7171,N_6551,N_6860);
nand U7172 (N_7172,N_6995,N_6545);
nor U7173 (N_7173,N_6965,N_6530);
nor U7174 (N_7174,N_6788,N_6538);
nor U7175 (N_7175,N_6969,N_6900);
and U7176 (N_7176,N_6921,N_6516);
nand U7177 (N_7177,N_6762,N_6766);
xnor U7178 (N_7178,N_6605,N_6759);
nand U7179 (N_7179,N_6940,N_6579);
or U7180 (N_7180,N_6942,N_6837);
or U7181 (N_7181,N_6654,N_6512);
nor U7182 (N_7182,N_6935,N_6943);
and U7183 (N_7183,N_6645,N_6720);
xnor U7184 (N_7184,N_6915,N_6792);
and U7185 (N_7185,N_6607,N_6845);
nand U7186 (N_7186,N_6569,N_6660);
or U7187 (N_7187,N_6828,N_6885);
xnor U7188 (N_7188,N_6844,N_6780);
nand U7189 (N_7189,N_6914,N_6919);
xnor U7190 (N_7190,N_6753,N_6997);
xnor U7191 (N_7191,N_6691,N_6939);
and U7192 (N_7192,N_6747,N_6768);
and U7193 (N_7193,N_6708,N_6836);
nand U7194 (N_7194,N_6559,N_6873);
xnor U7195 (N_7195,N_6867,N_6611);
nand U7196 (N_7196,N_6951,N_6529);
xnor U7197 (N_7197,N_6737,N_6923);
and U7198 (N_7198,N_6679,N_6689);
and U7199 (N_7199,N_6948,N_6841);
nor U7200 (N_7200,N_6640,N_6839);
xnor U7201 (N_7201,N_6667,N_6826);
xnor U7202 (N_7202,N_6726,N_6909);
and U7203 (N_7203,N_6657,N_6632);
xor U7204 (N_7204,N_6564,N_6713);
nor U7205 (N_7205,N_6922,N_6783);
or U7206 (N_7206,N_6561,N_6514);
xor U7207 (N_7207,N_6789,N_6596);
xor U7208 (N_7208,N_6587,N_6941);
or U7209 (N_7209,N_6880,N_6945);
nand U7210 (N_7210,N_6674,N_6810);
nor U7211 (N_7211,N_6804,N_6809);
xnor U7212 (N_7212,N_6625,N_6990);
nand U7213 (N_7213,N_6850,N_6745);
or U7214 (N_7214,N_6549,N_6659);
nor U7215 (N_7215,N_6819,N_6682);
or U7216 (N_7216,N_6670,N_6874);
xor U7217 (N_7217,N_6806,N_6756);
xor U7218 (N_7218,N_6572,N_6606);
and U7219 (N_7219,N_6527,N_6595);
xnor U7220 (N_7220,N_6678,N_6946);
or U7221 (N_7221,N_6958,N_6613);
nand U7222 (N_7222,N_6501,N_6580);
or U7223 (N_7223,N_6833,N_6535);
or U7224 (N_7224,N_6802,N_6510);
nor U7225 (N_7225,N_6830,N_6504);
nor U7226 (N_7226,N_6677,N_6960);
or U7227 (N_7227,N_6775,N_6727);
nand U7228 (N_7228,N_6705,N_6676);
and U7229 (N_7229,N_6541,N_6715);
nand U7230 (N_7230,N_6620,N_6592);
nand U7231 (N_7231,N_6849,N_6710);
nor U7232 (N_7232,N_6949,N_6934);
xor U7233 (N_7233,N_6520,N_6856);
or U7234 (N_7234,N_6508,N_6938);
nor U7235 (N_7235,N_6797,N_6754);
nor U7236 (N_7236,N_6642,N_6717);
nand U7237 (N_7237,N_6975,N_6602);
xnor U7238 (N_7238,N_6752,N_6816);
or U7239 (N_7239,N_6548,N_6814);
nor U7240 (N_7240,N_6617,N_6618);
nand U7241 (N_7241,N_6808,N_6861);
or U7242 (N_7242,N_6895,N_6570);
xor U7243 (N_7243,N_6906,N_6917);
and U7244 (N_7244,N_6699,N_6716);
or U7245 (N_7245,N_6698,N_6626);
nor U7246 (N_7246,N_6590,N_6953);
and U7247 (N_7247,N_6546,N_6604);
nand U7248 (N_7248,N_6598,N_6664);
and U7249 (N_7249,N_6871,N_6701);
nor U7250 (N_7250,N_6843,N_6927);
xnor U7251 (N_7251,N_6944,N_6922);
or U7252 (N_7252,N_6504,N_6697);
xnor U7253 (N_7253,N_6501,N_6958);
nor U7254 (N_7254,N_6789,N_6866);
or U7255 (N_7255,N_6951,N_6874);
and U7256 (N_7256,N_6726,N_6917);
xor U7257 (N_7257,N_6899,N_6508);
nor U7258 (N_7258,N_6829,N_6833);
nand U7259 (N_7259,N_6572,N_6845);
nand U7260 (N_7260,N_6915,N_6688);
or U7261 (N_7261,N_6947,N_6783);
or U7262 (N_7262,N_6771,N_6689);
nor U7263 (N_7263,N_6558,N_6525);
nor U7264 (N_7264,N_6871,N_6818);
nand U7265 (N_7265,N_6687,N_6918);
and U7266 (N_7266,N_6953,N_6988);
xor U7267 (N_7267,N_6737,N_6696);
and U7268 (N_7268,N_6678,N_6991);
xor U7269 (N_7269,N_6923,N_6664);
nor U7270 (N_7270,N_6671,N_6670);
and U7271 (N_7271,N_6614,N_6932);
xnor U7272 (N_7272,N_6702,N_6792);
nor U7273 (N_7273,N_6896,N_6742);
nor U7274 (N_7274,N_6962,N_6918);
nor U7275 (N_7275,N_6600,N_6501);
nand U7276 (N_7276,N_6942,N_6943);
or U7277 (N_7277,N_6952,N_6971);
and U7278 (N_7278,N_6863,N_6829);
nor U7279 (N_7279,N_6695,N_6710);
nand U7280 (N_7280,N_6582,N_6534);
and U7281 (N_7281,N_6605,N_6607);
xor U7282 (N_7282,N_6788,N_6689);
and U7283 (N_7283,N_6903,N_6953);
or U7284 (N_7284,N_6618,N_6749);
nand U7285 (N_7285,N_6861,N_6659);
xnor U7286 (N_7286,N_6866,N_6874);
nor U7287 (N_7287,N_6703,N_6927);
nor U7288 (N_7288,N_6587,N_6658);
or U7289 (N_7289,N_6954,N_6845);
nand U7290 (N_7290,N_6794,N_6720);
nand U7291 (N_7291,N_6590,N_6920);
nand U7292 (N_7292,N_6882,N_6871);
xnor U7293 (N_7293,N_6582,N_6518);
and U7294 (N_7294,N_6570,N_6515);
xnor U7295 (N_7295,N_6665,N_6835);
nor U7296 (N_7296,N_6958,N_6893);
xnor U7297 (N_7297,N_6820,N_6552);
or U7298 (N_7298,N_6999,N_6834);
and U7299 (N_7299,N_6674,N_6962);
nor U7300 (N_7300,N_6509,N_6748);
xor U7301 (N_7301,N_6649,N_6814);
and U7302 (N_7302,N_6514,N_6625);
and U7303 (N_7303,N_6740,N_6611);
nor U7304 (N_7304,N_6682,N_6538);
and U7305 (N_7305,N_6677,N_6622);
xor U7306 (N_7306,N_6703,N_6609);
nor U7307 (N_7307,N_6765,N_6568);
or U7308 (N_7308,N_6821,N_6871);
or U7309 (N_7309,N_6777,N_6666);
nand U7310 (N_7310,N_6899,N_6755);
or U7311 (N_7311,N_6667,N_6820);
nand U7312 (N_7312,N_6864,N_6663);
or U7313 (N_7313,N_6974,N_6550);
nand U7314 (N_7314,N_6576,N_6696);
nor U7315 (N_7315,N_6639,N_6747);
nand U7316 (N_7316,N_6635,N_6824);
nor U7317 (N_7317,N_6775,N_6840);
nand U7318 (N_7318,N_6920,N_6869);
nand U7319 (N_7319,N_6834,N_6837);
and U7320 (N_7320,N_6563,N_6892);
and U7321 (N_7321,N_6883,N_6871);
or U7322 (N_7322,N_6639,N_6718);
or U7323 (N_7323,N_6654,N_6881);
or U7324 (N_7324,N_6605,N_6877);
nor U7325 (N_7325,N_6943,N_6972);
or U7326 (N_7326,N_6617,N_6611);
nor U7327 (N_7327,N_6752,N_6566);
and U7328 (N_7328,N_6854,N_6987);
or U7329 (N_7329,N_6856,N_6708);
and U7330 (N_7330,N_6799,N_6616);
nor U7331 (N_7331,N_6568,N_6660);
and U7332 (N_7332,N_6712,N_6808);
nand U7333 (N_7333,N_6984,N_6994);
xor U7334 (N_7334,N_6774,N_6835);
xor U7335 (N_7335,N_6582,N_6653);
and U7336 (N_7336,N_6872,N_6743);
nor U7337 (N_7337,N_6856,N_6871);
nand U7338 (N_7338,N_6683,N_6532);
xnor U7339 (N_7339,N_6657,N_6952);
nor U7340 (N_7340,N_6705,N_6567);
nand U7341 (N_7341,N_6588,N_6805);
or U7342 (N_7342,N_6795,N_6744);
xor U7343 (N_7343,N_6847,N_6957);
and U7344 (N_7344,N_6788,N_6553);
and U7345 (N_7345,N_6751,N_6723);
xnor U7346 (N_7346,N_6878,N_6760);
nand U7347 (N_7347,N_6887,N_6538);
and U7348 (N_7348,N_6951,N_6894);
nand U7349 (N_7349,N_6500,N_6758);
nand U7350 (N_7350,N_6725,N_6776);
nor U7351 (N_7351,N_6992,N_6785);
and U7352 (N_7352,N_6738,N_6840);
and U7353 (N_7353,N_6766,N_6925);
nor U7354 (N_7354,N_6829,N_6800);
and U7355 (N_7355,N_6733,N_6822);
nor U7356 (N_7356,N_6657,N_6836);
nand U7357 (N_7357,N_6712,N_6909);
xor U7358 (N_7358,N_6580,N_6683);
and U7359 (N_7359,N_6542,N_6952);
xnor U7360 (N_7360,N_6928,N_6745);
nand U7361 (N_7361,N_6852,N_6573);
nand U7362 (N_7362,N_6792,N_6764);
xnor U7363 (N_7363,N_6823,N_6921);
or U7364 (N_7364,N_6723,N_6585);
and U7365 (N_7365,N_6746,N_6551);
nor U7366 (N_7366,N_6869,N_6804);
or U7367 (N_7367,N_6557,N_6711);
and U7368 (N_7368,N_6543,N_6549);
or U7369 (N_7369,N_6571,N_6784);
and U7370 (N_7370,N_6722,N_6922);
and U7371 (N_7371,N_6888,N_6850);
nor U7372 (N_7372,N_6726,N_6775);
nand U7373 (N_7373,N_6813,N_6680);
or U7374 (N_7374,N_6977,N_6661);
and U7375 (N_7375,N_6630,N_6609);
and U7376 (N_7376,N_6763,N_6738);
or U7377 (N_7377,N_6642,N_6526);
nand U7378 (N_7378,N_6815,N_6852);
and U7379 (N_7379,N_6503,N_6973);
xor U7380 (N_7380,N_6754,N_6956);
xor U7381 (N_7381,N_6895,N_6751);
nor U7382 (N_7382,N_6812,N_6919);
xor U7383 (N_7383,N_6806,N_6921);
nor U7384 (N_7384,N_6985,N_6976);
and U7385 (N_7385,N_6643,N_6614);
xor U7386 (N_7386,N_6894,N_6561);
xor U7387 (N_7387,N_6582,N_6975);
and U7388 (N_7388,N_6885,N_6887);
nand U7389 (N_7389,N_6805,N_6636);
and U7390 (N_7390,N_6532,N_6637);
nor U7391 (N_7391,N_6911,N_6605);
or U7392 (N_7392,N_6842,N_6939);
or U7393 (N_7393,N_6677,N_6733);
xor U7394 (N_7394,N_6925,N_6534);
xnor U7395 (N_7395,N_6633,N_6748);
nand U7396 (N_7396,N_6901,N_6833);
nand U7397 (N_7397,N_6831,N_6728);
or U7398 (N_7398,N_6894,N_6943);
xnor U7399 (N_7399,N_6596,N_6649);
or U7400 (N_7400,N_6646,N_6786);
nor U7401 (N_7401,N_6589,N_6635);
or U7402 (N_7402,N_6693,N_6715);
nor U7403 (N_7403,N_6729,N_6774);
and U7404 (N_7404,N_6506,N_6733);
nand U7405 (N_7405,N_6912,N_6776);
and U7406 (N_7406,N_6784,N_6996);
nand U7407 (N_7407,N_6848,N_6991);
or U7408 (N_7408,N_6693,N_6647);
nor U7409 (N_7409,N_6741,N_6780);
and U7410 (N_7410,N_6677,N_6986);
xor U7411 (N_7411,N_6746,N_6988);
and U7412 (N_7412,N_6781,N_6680);
nand U7413 (N_7413,N_6654,N_6511);
nor U7414 (N_7414,N_6501,N_6630);
xor U7415 (N_7415,N_6591,N_6715);
nand U7416 (N_7416,N_6647,N_6817);
xnor U7417 (N_7417,N_6761,N_6728);
nor U7418 (N_7418,N_6803,N_6513);
nand U7419 (N_7419,N_6714,N_6971);
or U7420 (N_7420,N_6877,N_6730);
and U7421 (N_7421,N_6809,N_6640);
xor U7422 (N_7422,N_6534,N_6623);
and U7423 (N_7423,N_6902,N_6897);
nand U7424 (N_7424,N_6600,N_6656);
and U7425 (N_7425,N_6565,N_6692);
nand U7426 (N_7426,N_6614,N_6597);
xnor U7427 (N_7427,N_6744,N_6528);
or U7428 (N_7428,N_6758,N_6771);
nand U7429 (N_7429,N_6672,N_6769);
nor U7430 (N_7430,N_6557,N_6975);
xnor U7431 (N_7431,N_6747,N_6591);
or U7432 (N_7432,N_6991,N_6638);
or U7433 (N_7433,N_6675,N_6593);
nand U7434 (N_7434,N_6961,N_6617);
nor U7435 (N_7435,N_6849,N_6751);
nand U7436 (N_7436,N_6985,N_6970);
xor U7437 (N_7437,N_6742,N_6920);
and U7438 (N_7438,N_6566,N_6647);
nand U7439 (N_7439,N_6786,N_6833);
and U7440 (N_7440,N_6742,N_6986);
or U7441 (N_7441,N_6627,N_6567);
or U7442 (N_7442,N_6680,N_6688);
and U7443 (N_7443,N_6962,N_6994);
nand U7444 (N_7444,N_6519,N_6835);
or U7445 (N_7445,N_6703,N_6908);
nand U7446 (N_7446,N_6705,N_6725);
xnor U7447 (N_7447,N_6670,N_6833);
nand U7448 (N_7448,N_6787,N_6665);
nand U7449 (N_7449,N_6950,N_6971);
xnor U7450 (N_7450,N_6720,N_6760);
xnor U7451 (N_7451,N_6745,N_6886);
nor U7452 (N_7452,N_6845,N_6543);
or U7453 (N_7453,N_6592,N_6673);
nor U7454 (N_7454,N_6687,N_6779);
xnor U7455 (N_7455,N_6841,N_6740);
or U7456 (N_7456,N_6612,N_6815);
nand U7457 (N_7457,N_6528,N_6549);
and U7458 (N_7458,N_6996,N_6816);
or U7459 (N_7459,N_6926,N_6641);
nand U7460 (N_7460,N_6632,N_6672);
nor U7461 (N_7461,N_6604,N_6867);
and U7462 (N_7462,N_6953,N_6760);
nor U7463 (N_7463,N_6612,N_6973);
or U7464 (N_7464,N_6859,N_6661);
nor U7465 (N_7465,N_6930,N_6607);
and U7466 (N_7466,N_6981,N_6949);
nor U7467 (N_7467,N_6651,N_6834);
nor U7468 (N_7468,N_6940,N_6913);
nor U7469 (N_7469,N_6693,N_6933);
xnor U7470 (N_7470,N_6665,N_6695);
and U7471 (N_7471,N_6900,N_6940);
nand U7472 (N_7472,N_6942,N_6624);
nand U7473 (N_7473,N_6878,N_6712);
xnor U7474 (N_7474,N_6819,N_6800);
or U7475 (N_7475,N_6732,N_6850);
nand U7476 (N_7476,N_6583,N_6810);
xnor U7477 (N_7477,N_6727,N_6645);
nand U7478 (N_7478,N_6794,N_6978);
nand U7479 (N_7479,N_6625,N_6787);
nand U7480 (N_7480,N_6743,N_6739);
and U7481 (N_7481,N_6957,N_6628);
and U7482 (N_7482,N_6817,N_6829);
nand U7483 (N_7483,N_6863,N_6665);
nand U7484 (N_7484,N_6850,N_6744);
nor U7485 (N_7485,N_6569,N_6703);
xor U7486 (N_7486,N_6593,N_6587);
nor U7487 (N_7487,N_6923,N_6873);
or U7488 (N_7488,N_6852,N_6595);
xor U7489 (N_7489,N_6550,N_6827);
or U7490 (N_7490,N_6986,N_6626);
or U7491 (N_7491,N_6554,N_6661);
xor U7492 (N_7492,N_6917,N_6618);
xor U7493 (N_7493,N_6674,N_6890);
nor U7494 (N_7494,N_6969,N_6828);
nand U7495 (N_7495,N_6754,N_6999);
xnor U7496 (N_7496,N_6891,N_6771);
xnor U7497 (N_7497,N_6703,N_6760);
and U7498 (N_7498,N_6766,N_6986);
xnor U7499 (N_7499,N_6869,N_6757);
nand U7500 (N_7500,N_7474,N_7195);
nor U7501 (N_7501,N_7233,N_7316);
and U7502 (N_7502,N_7134,N_7018);
and U7503 (N_7503,N_7486,N_7380);
xor U7504 (N_7504,N_7061,N_7019);
and U7505 (N_7505,N_7057,N_7127);
or U7506 (N_7506,N_7494,N_7144);
and U7507 (N_7507,N_7475,N_7011);
nand U7508 (N_7508,N_7010,N_7361);
nor U7509 (N_7509,N_7014,N_7277);
nand U7510 (N_7510,N_7304,N_7098);
nand U7511 (N_7511,N_7420,N_7188);
or U7512 (N_7512,N_7143,N_7293);
nand U7513 (N_7513,N_7251,N_7250);
xnor U7514 (N_7514,N_7036,N_7200);
or U7515 (N_7515,N_7184,N_7303);
or U7516 (N_7516,N_7295,N_7084);
nand U7517 (N_7517,N_7301,N_7159);
and U7518 (N_7518,N_7059,N_7377);
and U7519 (N_7519,N_7360,N_7418);
and U7520 (N_7520,N_7024,N_7083);
nand U7521 (N_7521,N_7442,N_7214);
nand U7522 (N_7522,N_7222,N_7359);
and U7523 (N_7523,N_7165,N_7462);
or U7524 (N_7524,N_7283,N_7108);
nand U7525 (N_7525,N_7070,N_7311);
or U7526 (N_7526,N_7048,N_7458);
xnor U7527 (N_7527,N_7490,N_7022);
nand U7528 (N_7528,N_7315,N_7308);
or U7529 (N_7529,N_7110,N_7479);
xnor U7530 (N_7530,N_7260,N_7470);
xnor U7531 (N_7531,N_7421,N_7082);
nor U7532 (N_7532,N_7254,N_7473);
or U7533 (N_7533,N_7234,N_7065);
or U7534 (N_7534,N_7428,N_7149);
nand U7535 (N_7535,N_7419,N_7258);
or U7536 (N_7536,N_7148,N_7236);
and U7537 (N_7537,N_7317,N_7069);
or U7538 (N_7538,N_7116,N_7383);
xor U7539 (N_7539,N_7128,N_7118);
or U7540 (N_7540,N_7422,N_7286);
and U7541 (N_7541,N_7297,N_7152);
nand U7542 (N_7542,N_7080,N_7169);
and U7543 (N_7543,N_7412,N_7459);
xor U7544 (N_7544,N_7212,N_7272);
or U7545 (N_7545,N_7203,N_7163);
xnor U7546 (N_7546,N_7046,N_7464);
and U7547 (N_7547,N_7215,N_7298);
xnor U7548 (N_7548,N_7241,N_7100);
and U7549 (N_7549,N_7035,N_7211);
nand U7550 (N_7550,N_7404,N_7399);
xor U7551 (N_7551,N_7284,N_7114);
or U7552 (N_7552,N_7385,N_7274);
or U7553 (N_7553,N_7410,N_7440);
nand U7554 (N_7554,N_7288,N_7193);
xor U7555 (N_7555,N_7405,N_7294);
nor U7556 (N_7556,N_7463,N_7223);
xor U7557 (N_7557,N_7173,N_7088);
xor U7558 (N_7558,N_7471,N_7480);
xnor U7559 (N_7559,N_7497,N_7492);
and U7560 (N_7560,N_7239,N_7041);
xor U7561 (N_7561,N_7091,N_7278);
nor U7562 (N_7562,N_7495,N_7244);
nor U7563 (N_7563,N_7089,N_7006);
nor U7564 (N_7564,N_7056,N_7264);
nand U7565 (N_7565,N_7265,N_7289);
nor U7566 (N_7566,N_7457,N_7228);
and U7567 (N_7567,N_7472,N_7003);
nor U7568 (N_7568,N_7229,N_7266);
xnor U7569 (N_7569,N_7324,N_7235);
nor U7570 (N_7570,N_7273,N_7125);
or U7571 (N_7571,N_7181,N_7431);
or U7572 (N_7572,N_7153,N_7281);
and U7573 (N_7573,N_7325,N_7269);
or U7574 (N_7574,N_7197,N_7130);
and U7575 (N_7575,N_7042,N_7077);
nand U7576 (N_7576,N_7392,N_7106);
and U7577 (N_7577,N_7452,N_7224);
and U7578 (N_7578,N_7226,N_7290);
or U7579 (N_7579,N_7007,N_7105);
or U7580 (N_7580,N_7285,N_7073);
and U7581 (N_7581,N_7104,N_7271);
xnor U7582 (N_7582,N_7496,N_7139);
nor U7583 (N_7583,N_7395,N_7300);
xor U7584 (N_7584,N_7432,N_7230);
or U7585 (N_7585,N_7085,N_7342);
and U7586 (N_7586,N_7255,N_7112);
nor U7587 (N_7587,N_7238,N_7190);
nor U7588 (N_7588,N_7199,N_7232);
and U7589 (N_7589,N_7373,N_7326);
or U7590 (N_7590,N_7086,N_7060);
nand U7591 (N_7591,N_7068,N_7033);
nand U7592 (N_7592,N_7156,N_7338);
xnor U7593 (N_7593,N_7052,N_7252);
nor U7594 (N_7594,N_7102,N_7242);
and U7595 (N_7595,N_7339,N_7292);
xnor U7596 (N_7596,N_7240,N_7146);
and U7597 (N_7597,N_7306,N_7346);
xnor U7598 (N_7598,N_7465,N_7047);
nor U7599 (N_7599,N_7245,N_7180);
nor U7600 (N_7600,N_7075,N_7142);
nand U7601 (N_7601,N_7424,N_7382);
and U7602 (N_7602,N_7225,N_7466);
nand U7603 (N_7603,N_7256,N_7078);
nand U7604 (N_7604,N_7093,N_7488);
xnor U7605 (N_7605,N_7357,N_7141);
xor U7606 (N_7606,N_7012,N_7337);
nand U7607 (N_7607,N_7013,N_7484);
and U7608 (N_7608,N_7429,N_7177);
nor U7609 (N_7609,N_7367,N_7436);
xor U7610 (N_7610,N_7220,N_7362);
or U7611 (N_7611,N_7121,N_7476);
or U7612 (N_7612,N_7498,N_7454);
nand U7613 (N_7613,N_7031,N_7145);
xor U7614 (N_7614,N_7002,N_7243);
and U7615 (N_7615,N_7341,N_7335);
xor U7616 (N_7616,N_7351,N_7167);
xnor U7617 (N_7617,N_7206,N_7123);
or U7618 (N_7618,N_7333,N_7249);
nand U7619 (N_7619,N_7210,N_7029);
nor U7620 (N_7620,N_7015,N_7231);
nand U7621 (N_7621,N_7066,N_7423);
nand U7622 (N_7622,N_7468,N_7364);
xnor U7623 (N_7623,N_7191,N_7433);
nand U7624 (N_7624,N_7170,N_7435);
or U7625 (N_7625,N_7322,N_7262);
or U7626 (N_7626,N_7328,N_7321);
or U7627 (N_7627,N_7209,N_7032);
xor U7628 (N_7628,N_7489,N_7179);
nor U7629 (N_7629,N_7296,N_7120);
and U7630 (N_7630,N_7138,N_7217);
or U7631 (N_7631,N_7336,N_7027);
and U7632 (N_7632,N_7081,N_7004);
and U7633 (N_7633,N_7379,N_7349);
nor U7634 (N_7634,N_7099,N_7332);
nor U7635 (N_7635,N_7441,N_7388);
xnor U7636 (N_7636,N_7402,N_7072);
nor U7637 (N_7637,N_7058,N_7071);
xor U7638 (N_7638,N_7017,N_7387);
xor U7639 (N_7639,N_7263,N_7166);
xnor U7640 (N_7640,N_7347,N_7168);
nand U7641 (N_7641,N_7270,N_7446);
nand U7642 (N_7642,N_7450,N_7447);
or U7643 (N_7643,N_7461,N_7136);
and U7644 (N_7644,N_7493,N_7299);
nand U7645 (N_7645,N_7135,N_7049);
nor U7646 (N_7646,N_7064,N_7430);
nor U7647 (N_7647,N_7096,N_7327);
nand U7648 (N_7648,N_7400,N_7378);
nand U7649 (N_7649,N_7095,N_7371);
xor U7650 (N_7650,N_7381,N_7318);
nand U7651 (N_7651,N_7067,N_7227);
nor U7652 (N_7652,N_7202,N_7055);
xor U7653 (N_7653,N_7097,N_7122);
or U7654 (N_7654,N_7408,N_7111);
and U7655 (N_7655,N_7449,N_7183);
nand U7656 (N_7656,N_7157,N_7023);
nor U7657 (N_7657,N_7026,N_7276);
nor U7658 (N_7658,N_7314,N_7030);
nand U7659 (N_7659,N_7375,N_7374);
nor U7660 (N_7660,N_7354,N_7054);
xor U7661 (N_7661,N_7398,N_7140);
and U7662 (N_7662,N_7219,N_7185);
and U7663 (N_7663,N_7154,N_7267);
xor U7664 (N_7664,N_7103,N_7074);
nor U7665 (N_7665,N_7365,N_7247);
nor U7666 (N_7666,N_7455,N_7482);
xnor U7667 (N_7667,N_7133,N_7391);
and U7668 (N_7668,N_7028,N_7034);
or U7669 (N_7669,N_7040,N_7370);
nor U7670 (N_7670,N_7119,N_7129);
and U7671 (N_7671,N_7350,N_7376);
and U7672 (N_7672,N_7045,N_7323);
or U7673 (N_7673,N_7407,N_7309);
nor U7674 (N_7674,N_7204,N_7147);
or U7675 (N_7675,N_7115,N_7356);
nor U7676 (N_7676,N_7389,N_7192);
xor U7677 (N_7677,N_7016,N_7481);
xor U7678 (N_7678,N_7394,N_7182);
and U7679 (N_7679,N_7396,N_7008);
nand U7680 (N_7680,N_7174,N_7038);
and U7681 (N_7681,N_7443,N_7319);
nor U7682 (N_7682,N_7094,N_7268);
or U7683 (N_7683,N_7390,N_7403);
xnor U7684 (N_7684,N_7310,N_7305);
xnor U7685 (N_7685,N_7437,N_7107);
and U7686 (N_7686,N_7216,N_7487);
or U7687 (N_7687,N_7090,N_7384);
or U7688 (N_7688,N_7434,N_7050);
nor U7689 (N_7689,N_7313,N_7280);
and U7690 (N_7690,N_7162,N_7161);
or U7691 (N_7691,N_7416,N_7330);
nand U7692 (N_7692,N_7397,N_7025);
xor U7693 (N_7693,N_7261,N_7079);
or U7694 (N_7694,N_7363,N_7287);
xnor U7695 (N_7695,N_7001,N_7248);
and U7696 (N_7696,N_7372,N_7087);
xnor U7697 (N_7697,N_7246,N_7151);
nor U7698 (N_7698,N_7453,N_7413);
and U7699 (N_7699,N_7386,N_7051);
xor U7700 (N_7700,N_7196,N_7483);
or U7701 (N_7701,N_7340,N_7158);
and U7702 (N_7702,N_7160,N_7021);
nand U7703 (N_7703,N_7417,N_7207);
xnor U7704 (N_7704,N_7150,N_7499);
nor U7705 (N_7705,N_7092,N_7155);
and U7706 (N_7706,N_7175,N_7076);
xor U7707 (N_7707,N_7329,N_7414);
nand U7708 (N_7708,N_7352,N_7164);
xnor U7709 (N_7709,N_7439,N_7198);
nand U7710 (N_7710,N_7425,N_7005);
and U7711 (N_7711,N_7109,N_7478);
or U7712 (N_7712,N_7237,N_7427);
xor U7713 (N_7713,N_7456,N_7124);
nor U7714 (N_7714,N_7320,N_7218);
or U7715 (N_7715,N_7409,N_7187);
and U7716 (N_7716,N_7291,N_7355);
nor U7717 (N_7717,N_7369,N_7132);
nor U7718 (N_7718,N_7366,N_7176);
xor U7719 (N_7719,N_7368,N_7000);
nor U7720 (N_7720,N_7172,N_7444);
or U7721 (N_7721,N_7348,N_7415);
and U7722 (N_7722,N_7137,N_7194);
or U7723 (N_7723,N_7221,N_7171);
or U7724 (N_7724,N_7101,N_7393);
and U7725 (N_7725,N_7126,N_7113);
or U7726 (N_7726,N_7253,N_7205);
nand U7727 (N_7727,N_7331,N_7020);
xnor U7728 (N_7728,N_7053,N_7279);
nor U7729 (N_7729,N_7401,N_7445);
nor U7730 (N_7730,N_7063,N_7460);
nand U7731 (N_7731,N_7302,N_7343);
nand U7732 (N_7732,N_7469,N_7039);
nand U7733 (N_7733,N_7344,N_7477);
and U7734 (N_7734,N_7037,N_7448);
xnor U7735 (N_7735,N_7353,N_7009);
nor U7736 (N_7736,N_7334,N_7208);
and U7737 (N_7737,N_7438,N_7213);
and U7738 (N_7738,N_7044,N_7117);
nand U7739 (N_7739,N_7043,N_7467);
nor U7740 (N_7740,N_7201,N_7189);
and U7741 (N_7741,N_7282,N_7491);
xnor U7742 (N_7742,N_7426,N_7345);
nor U7743 (N_7743,N_7062,N_7131);
nor U7744 (N_7744,N_7178,N_7451);
nand U7745 (N_7745,N_7358,N_7411);
or U7746 (N_7746,N_7485,N_7406);
nand U7747 (N_7747,N_7312,N_7307);
nor U7748 (N_7748,N_7257,N_7275);
nand U7749 (N_7749,N_7186,N_7259);
and U7750 (N_7750,N_7391,N_7092);
and U7751 (N_7751,N_7495,N_7057);
nor U7752 (N_7752,N_7307,N_7026);
or U7753 (N_7753,N_7248,N_7153);
or U7754 (N_7754,N_7096,N_7180);
or U7755 (N_7755,N_7208,N_7154);
xor U7756 (N_7756,N_7142,N_7111);
nor U7757 (N_7757,N_7075,N_7106);
or U7758 (N_7758,N_7060,N_7296);
nand U7759 (N_7759,N_7248,N_7112);
and U7760 (N_7760,N_7252,N_7273);
or U7761 (N_7761,N_7159,N_7216);
or U7762 (N_7762,N_7115,N_7352);
or U7763 (N_7763,N_7347,N_7179);
nor U7764 (N_7764,N_7413,N_7041);
nor U7765 (N_7765,N_7280,N_7099);
nand U7766 (N_7766,N_7128,N_7328);
or U7767 (N_7767,N_7070,N_7324);
or U7768 (N_7768,N_7054,N_7186);
or U7769 (N_7769,N_7353,N_7245);
and U7770 (N_7770,N_7033,N_7349);
or U7771 (N_7771,N_7406,N_7438);
nand U7772 (N_7772,N_7273,N_7320);
and U7773 (N_7773,N_7354,N_7344);
xor U7774 (N_7774,N_7350,N_7140);
nor U7775 (N_7775,N_7332,N_7139);
or U7776 (N_7776,N_7306,N_7058);
or U7777 (N_7777,N_7447,N_7476);
and U7778 (N_7778,N_7466,N_7219);
nor U7779 (N_7779,N_7280,N_7087);
xor U7780 (N_7780,N_7273,N_7454);
nand U7781 (N_7781,N_7060,N_7116);
nand U7782 (N_7782,N_7249,N_7391);
or U7783 (N_7783,N_7315,N_7120);
and U7784 (N_7784,N_7115,N_7043);
nand U7785 (N_7785,N_7074,N_7145);
and U7786 (N_7786,N_7297,N_7291);
xnor U7787 (N_7787,N_7312,N_7348);
nor U7788 (N_7788,N_7055,N_7113);
xor U7789 (N_7789,N_7483,N_7105);
or U7790 (N_7790,N_7412,N_7229);
nor U7791 (N_7791,N_7443,N_7025);
or U7792 (N_7792,N_7346,N_7090);
nand U7793 (N_7793,N_7366,N_7158);
nor U7794 (N_7794,N_7467,N_7307);
xor U7795 (N_7795,N_7289,N_7272);
nor U7796 (N_7796,N_7020,N_7138);
or U7797 (N_7797,N_7367,N_7198);
or U7798 (N_7798,N_7350,N_7417);
or U7799 (N_7799,N_7151,N_7133);
nor U7800 (N_7800,N_7396,N_7225);
nor U7801 (N_7801,N_7219,N_7258);
nand U7802 (N_7802,N_7148,N_7035);
or U7803 (N_7803,N_7407,N_7205);
and U7804 (N_7804,N_7353,N_7312);
nor U7805 (N_7805,N_7367,N_7304);
xor U7806 (N_7806,N_7104,N_7333);
or U7807 (N_7807,N_7071,N_7029);
or U7808 (N_7808,N_7162,N_7398);
xor U7809 (N_7809,N_7173,N_7158);
or U7810 (N_7810,N_7013,N_7095);
nand U7811 (N_7811,N_7119,N_7177);
or U7812 (N_7812,N_7085,N_7381);
nor U7813 (N_7813,N_7480,N_7436);
and U7814 (N_7814,N_7385,N_7439);
xnor U7815 (N_7815,N_7252,N_7084);
and U7816 (N_7816,N_7224,N_7409);
or U7817 (N_7817,N_7050,N_7077);
nand U7818 (N_7818,N_7141,N_7334);
xor U7819 (N_7819,N_7121,N_7410);
xor U7820 (N_7820,N_7137,N_7436);
or U7821 (N_7821,N_7047,N_7166);
or U7822 (N_7822,N_7487,N_7238);
xor U7823 (N_7823,N_7444,N_7148);
or U7824 (N_7824,N_7047,N_7215);
or U7825 (N_7825,N_7415,N_7024);
and U7826 (N_7826,N_7412,N_7246);
nand U7827 (N_7827,N_7024,N_7284);
nor U7828 (N_7828,N_7037,N_7143);
nor U7829 (N_7829,N_7282,N_7406);
nand U7830 (N_7830,N_7495,N_7126);
nor U7831 (N_7831,N_7481,N_7488);
xnor U7832 (N_7832,N_7477,N_7359);
xor U7833 (N_7833,N_7303,N_7442);
nor U7834 (N_7834,N_7379,N_7126);
nand U7835 (N_7835,N_7159,N_7494);
nor U7836 (N_7836,N_7336,N_7309);
and U7837 (N_7837,N_7278,N_7490);
xnor U7838 (N_7838,N_7137,N_7147);
nand U7839 (N_7839,N_7089,N_7495);
and U7840 (N_7840,N_7073,N_7288);
xnor U7841 (N_7841,N_7252,N_7205);
and U7842 (N_7842,N_7223,N_7094);
nor U7843 (N_7843,N_7275,N_7162);
nor U7844 (N_7844,N_7476,N_7127);
nor U7845 (N_7845,N_7251,N_7134);
and U7846 (N_7846,N_7466,N_7264);
or U7847 (N_7847,N_7479,N_7397);
or U7848 (N_7848,N_7186,N_7124);
or U7849 (N_7849,N_7360,N_7294);
and U7850 (N_7850,N_7100,N_7272);
nor U7851 (N_7851,N_7253,N_7131);
or U7852 (N_7852,N_7355,N_7127);
and U7853 (N_7853,N_7435,N_7012);
nand U7854 (N_7854,N_7003,N_7066);
nand U7855 (N_7855,N_7186,N_7120);
xor U7856 (N_7856,N_7286,N_7125);
nand U7857 (N_7857,N_7194,N_7007);
nand U7858 (N_7858,N_7106,N_7031);
nor U7859 (N_7859,N_7233,N_7292);
xor U7860 (N_7860,N_7006,N_7248);
and U7861 (N_7861,N_7085,N_7048);
or U7862 (N_7862,N_7162,N_7465);
nor U7863 (N_7863,N_7410,N_7016);
or U7864 (N_7864,N_7417,N_7013);
and U7865 (N_7865,N_7433,N_7294);
or U7866 (N_7866,N_7442,N_7253);
and U7867 (N_7867,N_7107,N_7300);
nor U7868 (N_7868,N_7379,N_7442);
nand U7869 (N_7869,N_7063,N_7213);
and U7870 (N_7870,N_7136,N_7308);
xor U7871 (N_7871,N_7242,N_7464);
or U7872 (N_7872,N_7386,N_7219);
nand U7873 (N_7873,N_7332,N_7419);
or U7874 (N_7874,N_7012,N_7097);
nor U7875 (N_7875,N_7170,N_7202);
nand U7876 (N_7876,N_7071,N_7085);
nand U7877 (N_7877,N_7288,N_7058);
nor U7878 (N_7878,N_7326,N_7101);
and U7879 (N_7879,N_7345,N_7262);
xnor U7880 (N_7880,N_7239,N_7371);
nor U7881 (N_7881,N_7391,N_7461);
and U7882 (N_7882,N_7467,N_7151);
xor U7883 (N_7883,N_7141,N_7142);
xnor U7884 (N_7884,N_7464,N_7327);
nand U7885 (N_7885,N_7457,N_7341);
nor U7886 (N_7886,N_7184,N_7459);
and U7887 (N_7887,N_7134,N_7204);
nand U7888 (N_7888,N_7324,N_7330);
nor U7889 (N_7889,N_7022,N_7143);
xnor U7890 (N_7890,N_7293,N_7415);
and U7891 (N_7891,N_7114,N_7192);
nand U7892 (N_7892,N_7032,N_7172);
nand U7893 (N_7893,N_7114,N_7151);
nand U7894 (N_7894,N_7399,N_7156);
nand U7895 (N_7895,N_7377,N_7088);
nor U7896 (N_7896,N_7414,N_7106);
or U7897 (N_7897,N_7225,N_7227);
nor U7898 (N_7898,N_7384,N_7058);
xnor U7899 (N_7899,N_7402,N_7238);
and U7900 (N_7900,N_7430,N_7345);
nand U7901 (N_7901,N_7149,N_7153);
nor U7902 (N_7902,N_7126,N_7375);
and U7903 (N_7903,N_7457,N_7452);
nand U7904 (N_7904,N_7080,N_7260);
nand U7905 (N_7905,N_7343,N_7433);
and U7906 (N_7906,N_7272,N_7327);
nor U7907 (N_7907,N_7085,N_7088);
nand U7908 (N_7908,N_7341,N_7348);
xor U7909 (N_7909,N_7134,N_7043);
and U7910 (N_7910,N_7063,N_7157);
xor U7911 (N_7911,N_7276,N_7193);
nand U7912 (N_7912,N_7279,N_7246);
and U7913 (N_7913,N_7289,N_7263);
xor U7914 (N_7914,N_7099,N_7466);
nand U7915 (N_7915,N_7082,N_7233);
xnor U7916 (N_7916,N_7369,N_7027);
nand U7917 (N_7917,N_7259,N_7224);
and U7918 (N_7918,N_7227,N_7379);
nand U7919 (N_7919,N_7129,N_7105);
xnor U7920 (N_7920,N_7271,N_7138);
nor U7921 (N_7921,N_7255,N_7302);
nand U7922 (N_7922,N_7338,N_7236);
nor U7923 (N_7923,N_7088,N_7067);
xnor U7924 (N_7924,N_7061,N_7418);
xor U7925 (N_7925,N_7476,N_7489);
or U7926 (N_7926,N_7279,N_7346);
nand U7927 (N_7927,N_7240,N_7366);
or U7928 (N_7928,N_7370,N_7066);
or U7929 (N_7929,N_7310,N_7007);
and U7930 (N_7930,N_7211,N_7293);
and U7931 (N_7931,N_7453,N_7086);
nor U7932 (N_7932,N_7402,N_7360);
or U7933 (N_7933,N_7383,N_7039);
xor U7934 (N_7934,N_7420,N_7415);
nand U7935 (N_7935,N_7173,N_7278);
nand U7936 (N_7936,N_7136,N_7071);
or U7937 (N_7937,N_7372,N_7262);
nand U7938 (N_7938,N_7167,N_7312);
and U7939 (N_7939,N_7141,N_7127);
xnor U7940 (N_7940,N_7263,N_7152);
nand U7941 (N_7941,N_7306,N_7211);
nand U7942 (N_7942,N_7076,N_7449);
or U7943 (N_7943,N_7432,N_7179);
nor U7944 (N_7944,N_7036,N_7498);
nor U7945 (N_7945,N_7016,N_7464);
nand U7946 (N_7946,N_7067,N_7222);
nand U7947 (N_7947,N_7309,N_7408);
and U7948 (N_7948,N_7017,N_7424);
nand U7949 (N_7949,N_7353,N_7003);
and U7950 (N_7950,N_7352,N_7343);
or U7951 (N_7951,N_7395,N_7490);
or U7952 (N_7952,N_7353,N_7123);
nor U7953 (N_7953,N_7169,N_7125);
nor U7954 (N_7954,N_7282,N_7064);
nor U7955 (N_7955,N_7064,N_7193);
and U7956 (N_7956,N_7269,N_7046);
xor U7957 (N_7957,N_7416,N_7207);
and U7958 (N_7958,N_7170,N_7347);
and U7959 (N_7959,N_7254,N_7436);
and U7960 (N_7960,N_7385,N_7167);
or U7961 (N_7961,N_7161,N_7061);
nor U7962 (N_7962,N_7068,N_7477);
or U7963 (N_7963,N_7144,N_7230);
xnor U7964 (N_7964,N_7313,N_7466);
and U7965 (N_7965,N_7035,N_7381);
xor U7966 (N_7966,N_7127,N_7402);
or U7967 (N_7967,N_7460,N_7370);
nand U7968 (N_7968,N_7345,N_7215);
or U7969 (N_7969,N_7407,N_7166);
xor U7970 (N_7970,N_7009,N_7266);
or U7971 (N_7971,N_7391,N_7105);
and U7972 (N_7972,N_7205,N_7399);
nand U7973 (N_7973,N_7248,N_7119);
or U7974 (N_7974,N_7014,N_7067);
or U7975 (N_7975,N_7371,N_7481);
nor U7976 (N_7976,N_7266,N_7023);
xnor U7977 (N_7977,N_7023,N_7231);
nor U7978 (N_7978,N_7278,N_7211);
xor U7979 (N_7979,N_7185,N_7241);
nor U7980 (N_7980,N_7011,N_7482);
nor U7981 (N_7981,N_7124,N_7424);
or U7982 (N_7982,N_7396,N_7335);
and U7983 (N_7983,N_7487,N_7323);
nor U7984 (N_7984,N_7210,N_7401);
or U7985 (N_7985,N_7080,N_7347);
and U7986 (N_7986,N_7290,N_7208);
nor U7987 (N_7987,N_7393,N_7147);
nor U7988 (N_7988,N_7268,N_7278);
or U7989 (N_7989,N_7381,N_7068);
and U7990 (N_7990,N_7087,N_7290);
nand U7991 (N_7991,N_7168,N_7014);
nand U7992 (N_7992,N_7288,N_7228);
and U7993 (N_7993,N_7014,N_7412);
and U7994 (N_7994,N_7416,N_7229);
xor U7995 (N_7995,N_7027,N_7002);
xor U7996 (N_7996,N_7324,N_7301);
nor U7997 (N_7997,N_7253,N_7356);
and U7998 (N_7998,N_7249,N_7198);
xor U7999 (N_7999,N_7370,N_7061);
nand U8000 (N_8000,N_7616,N_7711);
and U8001 (N_8001,N_7821,N_7947);
and U8002 (N_8002,N_7690,N_7559);
nand U8003 (N_8003,N_7517,N_7659);
xnor U8004 (N_8004,N_7533,N_7555);
nand U8005 (N_8005,N_7924,N_7814);
nand U8006 (N_8006,N_7512,N_7648);
and U8007 (N_8007,N_7591,N_7743);
or U8008 (N_8008,N_7799,N_7791);
or U8009 (N_8009,N_7553,N_7828);
nand U8010 (N_8010,N_7674,N_7696);
xnor U8011 (N_8011,N_7515,N_7573);
nand U8012 (N_8012,N_7632,N_7557);
nor U8013 (N_8013,N_7840,N_7992);
nand U8014 (N_8014,N_7815,N_7704);
or U8015 (N_8015,N_7646,N_7508);
or U8016 (N_8016,N_7778,N_7755);
nor U8017 (N_8017,N_7671,N_7505);
nor U8018 (N_8018,N_7619,N_7862);
nand U8019 (N_8019,N_7570,N_7919);
and U8020 (N_8020,N_7695,N_7590);
xor U8021 (N_8021,N_7945,N_7863);
and U8022 (N_8022,N_7528,N_7628);
nor U8023 (N_8023,N_7750,N_7621);
nor U8024 (N_8024,N_7857,N_7661);
and U8025 (N_8025,N_7527,N_7685);
nand U8026 (N_8026,N_7982,N_7891);
nand U8027 (N_8027,N_7532,N_7904);
and U8028 (N_8028,N_7804,N_7538);
or U8029 (N_8029,N_7562,N_7941);
or U8030 (N_8030,N_7903,N_7726);
xor U8031 (N_8031,N_7795,N_7595);
nor U8032 (N_8032,N_7762,N_7680);
nor U8033 (N_8033,N_7763,N_7751);
nor U8034 (N_8034,N_7725,N_7733);
nand U8035 (N_8035,N_7567,N_7594);
or U8036 (N_8036,N_7723,N_7965);
nand U8037 (N_8037,N_7636,N_7881);
xor U8038 (N_8038,N_7883,N_7705);
xnor U8039 (N_8039,N_7768,N_7842);
and U8040 (N_8040,N_7806,N_7601);
and U8041 (N_8041,N_7959,N_7753);
nand U8042 (N_8042,N_7727,N_7805);
nor U8043 (N_8043,N_7776,N_7735);
nor U8044 (N_8044,N_7874,N_7906);
and U8045 (N_8045,N_7630,N_7608);
nor U8046 (N_8046,N_7544,N_7740);
nor U8047 (N_8047,N_7966,N_7820);
nand U8048 (N_8048,N_7866,N_7558);
nor U8049 (N_8049,N_7757,N_7638);
or U8050 (N_8050,N_7599,N_7925);
nor U8051 (N_8051,N_7810,N_7689);
xnor U8052 (N_8052,N_7998,N_7789);
xnor U8053 (N_8053,N_7730,N_7737);
or U8054 (N_8054,N_7949,N_7961);
nand U8055 (N_8055,N_7835,N_7930);
nand U8056 (N_8056,N_7698,N_7653);
and U8057 (N_8057,N_7975,N_7641);
nor U8058 (N_8058,N_7932,N_7770);
or U8059 (N_8059,N_7662,N_7644);
and U8060 (N_8060,N_7513,N_7584);
nand U8061 (N_8061,N_7660,N_7542);
and U8062 (N_8062,N_7909,N_7536);
xor U8063 (N_8063,N_7817,N_7780);
and U8064 (N_8064,N_7784,N_7859);
and U8065 (N_8065,N_7718,N_7502);
xnor U8066 (N_8066,N_7772,N_7860);
or U8067 (N_8067,N_7955,N_7715);
nand U8068 (N_8068,N_7869,N_7957);
and U8069 (N_8069,N_7877,N_7731);
nor U8070 (N_8070,N_7938,N_7978);
or U8071 (N_8071,N_7501,N_7734);
or U8072 (N_8072,N_7958,N_7574);
or U8073 (N_8073,N_7652,N_7886);
and U8074 (N_8074,N_7972,N_7971);
nor U8075 (N_8075,N_7892,N_7525);
or U8076 (N_8076,N_7803,N_7645);
nand U8077 (N_8077,N_7767,N_7822);
xnor U8078 (N_8078,N_7576,N_7546);
or U8079 (N_8079,N_7607,N_7639);
nor U8080 (N_8080,N_7537,N_7995);
nor U8081 (N_8081,N_7769,N_7758);
xor U8082 (N_8082,N_7667,N_7716);
and U8083 (N_8083,N_7597,N_7624);
nor U8084 (N_8084,N_7854,N_7953);
or U8085 (N_8085,N_7617,N_7896);
or U8086 (N_8086,N_7708,N_7600);
or U8087 (N_8087,N_7897,N_7974);
nor U8088 (N_8088,N_7640,N_7592);
nor U8089 (N_8089,N_7848,N_7876);
xnor U8090 (N_8090,N_7765,N_7677);
or U8091 (N_8091,N_7986,N_7732);
nor U8092 (N_8092,N_7623,N_7937);
and U8093 (N_8093,N_7752,N_7818);
nand U8094 (N_8094,N_7686,N_7707);
xor U8095 (N_8095,N_7681,N_7787);
nor U8096 (N_8096,N_7613,N_7626);
nand U8097 (N_8097,N_7720,N_7916);
and U8098 (N_8098,N_7552,N_7606);
nor U8099 (N_8099,N_7976,N_7988);
nor U8100 (N_8100,N_7847,N_7846);
nand U8101 (N_8101,N_7913,N_7530);
or U8102 (N_8102,N_7738,N_7794);
xnor U8103 (N_8103,N_7921,N_7614);
or U8104 (N_8104,N_7907,N_7990);
and U8105 (N_8105,N_7816,N_7654);
xnor U8106 (N_8106,N_7663,N_7510);
or U8107 (N_8107,N_7657,N_7692);
xor U8108 (N_8108,N_7593,N_7699);
xnor U8109 (N_8109,N_7811,N_7887);
nand U8110 (N_8110,N_7761,N_7518);
nor U8111 (N_8111,N_7843,N_7893);
xor U8112 (N_8112,N_7741,N_7809);
or U8113 (N_8113,N_7724,N_7878);
xnor U8114 (N_8114,N_7968,N_7611);
nor U8115 (N_8115,N_7861,N_7849);
nand U8116 (N_8116,N_7951,N_7545);
nand U8117 (N_8117,N_7523,N_7929);
or U8118 (N_8118,N_7952,N_7580);
or U8119 (N_8119,N_7845,N_7808);
xnor U8120 (N_8120,N_7717,N_7826);
and U8121 (N_8121,N_7571,N_7651);
nand U8122 (N_8122,N_7844,N_7813);
and U8123 (N_8123,N_7775,N_7801);
nand U8124 (N_8124,N_7588,N_7710);
xor U8125 (N_8125,N_7979,N_7867);
nand U8126 (N_8126,N_7500,N_7864);
xnor U8127 (N_8127,N_7694,N_7933);
xor U8128 (N_8128,N_7931,N_7839);
or U8129 (N_8129,N_7868,N_7964);
nand U8130 (N_8130,N_7910,N_7792);
or U8131 (N_8131,N_7785,N_7850);
nor U8132 (N_8132,N_7788,N_7550);
nor U8133 (N_8133,N_7855,N_7798);
xor U8134 (N_8134,N_7678,N_7920);
or U8135 (N_8135,N_7977,N_7534);
and U8136 (N_8136,N_7577,N_7911);
nand U8137 (N_8137,N_7889,N_7650);
xor U8138 (N_8138,N_7985,N_7541);
nor U8139 (N_8139,N_7946,N_7746);
xor U8140 (N_8140,N_7983,N_7719);
xor U8141 (N_8141,N_7669,N_7970);
xor U8142 (N_8142,N_7918,N_7915);
xor U8143 (N_8143,N_7980,N_7962);
nand U8144 (N_8144,N_7637,N_7880);
nor U8145 (N_8145,N_7908,N_7566);
or U8146 (N_8146,N_7547,N_7543);
or U8147 (N_8147,N_7631,N_7668);
nand U8148 (N_8148,N_7742,N_7928);
or U8149 (N_8149,N_7782,N_7647);
nor U8150 (N_8150,N_7643,N_7526);
nor U8151 (N_8151,N_7994,N_7879);
xnor U8152 (N_8152,N_7587,N_7954);
and U8153 (N_8153,N_7996,N_7511);
nand U8154 (N_8154,N_7745,N_7923);
or U8155 (N_8155,N_7830,N_7598);
or U8156 (N_8156,N_7771,N_7605);
xnor U8157 (N_8157,N_7756,N_7882);
or U8158 (N_8158,N_7890,N_7898);
nand U8159 (N_8159,N_7781,N_7516);
or U8160 (N_8160,N_7684,N_7540);
and U8161 (N_8161,N_7569,N_7712);
xor U8162 (N_8162,N_7841,N_7926);
nor U8163 (N_8163,N_7520,N_7833);
and U8164 (N_8164,N_7675,N_7539);
nor U8165 (N_8165,N_7851,N_7853);
or U8166 (N_8166,N_7509,N_7714);
nand U8167 (N_8167,N_7852,N_7575);
or U8168 (N_8168,N_7672,N_7514);
xnor U8169 (N_8169,N_7506,N_7936);
nand U8170 (N_8170,N_7800,N_7917);
or U8171 (N_8171,N_7825,N_7635);
or U8172 (N_8172,N_7560,N_7549);
nor U8173 (N_8173,N_7610,N_7629);
or U8174 (N_8174,N_7688,N_7589);
or U8175 (N_8175,N_7942,N_7940);
nand U8176 (N_8176,N_7529,N_7670);
nand U8177 (N_8177,N_7673,N_7873);
nor U8178 (N_8178,N_7535,N_7999);
and U8179 (N_8179,N_7665,N_7615);
and U8180 (N_8180,N_7894,N_7895);
nor U8181 (N_8181,N_7691,N_7902);
nor U8182 (N_8182,N_7701,N_7900);
nor U8183 (N_8183,N_7749,N_7697);
nor U8184 (N_8184,N_7683,N_7578);
or U8185 (N_8185,N_7922,N_7656);
xor U8186 (N_8186,N_7649,N_7831);
nor U8187 (N_8187,N_7747,N_7875);
xnor U8188 (N_8188,N_7989,N_7948);
and U8189 (N_8189,N_7905,N_7790);
and U8190 (N_8190,N_7759,N_7773);
or U8191 (N_8191,N_7779,N_7797);
nor U8192 (N_8192,N_7604,N_7524);
or U8193 (N_8193,N_7997,N_7884);
nor U8194 (N_8194,N_7618,N_7682);
and U8195 (N_8195,N_7981,N_7991);
nor U8196 (N_8196,N_7872,N_7812);
nor U8197 (N_8197,N_7522,N_7777);
and U8198 (N_8198,N_7693,N_7581);
xor U8199 (N_8199,N_7658,N_7993);
xnor U8200 (N_8200,N_7967,N_7796);
xor U8201 (N_8201,N_7585,N_7807);
nor U8202 (N_8202,N_7634,N_7565);
nand U8203 (N_8203,N_7579,N_7960);
or U8204 (N_8204,N_7944,N_7721);
nor U8205 (N_8205,N_7582,N_7824);
or U8206 (N_8206,N_7563,N_7722);
nor U8207 (N_8207,N_7973,N_7620);
xnor U8208 (N_8208,N_7766,N_7950);
nor U8209 (N_8209,N_7503,N_7865);
and U8210 (N_8210,N_7802,N_7956);
nand U8211 (N_8211,N_7834,N_7561);
nor U8212 (N_8212,N_7736,N_7912);
and U8213 (N_8213,N_7519,N_7642);
or U8214 (N_8214,N_7838,N_7786);
nand U8215 (N_8215,N_7703,N_7856);
nor U8216 (N_8216,N_7551,N_7939);
nor U8217 (N_8217,N_7748,N_7633);
or U8218 (N_8218,N_7603,N_7793);
xor U8219 (N_8219,N_7664,N_7602);
nor U8220 (N_8220,N_7564,N_7548);
nand U8221 (N_8221,N_7702,N_7679);
nor U8222 (N_8222,N_7521,N_7531);
or U8223 (N_8223,N_7687,N_7625);
nand U8224 (N_8224,N_7709,N_7969);
xnor U8225 (N_8225,N_7819,N_7764);
xor U8226 (N_8226,N_7612,N_7568);
xor U8227 (N_8227,N_7774,N_7823);
nand U8228 (N_8228,N_7556,N_7899);
xor U8229 (N_8229,N_7836,N_7934);
and U8230 (N_8230,N_7984,N_7622);
nand U8231 (N_8231,N_7507,N_7885);
xnor U8232 (N_8232,N_7739,N_7700);
nor U8233 (N_8233,N_7706,N_7914);
and U8234 (N_8234,N_7888,N_7871);
nand U8235 (N_8235,N_7870,N_7943);
or U8236 (N_8236,N_7858,N_7729);
or U8237 (N_8237,N_7832,N_7554);
and U8238 (N_8238,N_7713,N_7666);
xor U8239 (N_8239,N_7728,N_7609);
nand U8240 (N_8240,N_7760,N_7583);
nand U8241 (N_8241,N_7935,N_7837);
nand U8242 (N_8242,N_7596,N_7655);
xnor U8243 (N_8243,N_7987,N_7504);
nor U8244 (N_8244,N_7783,N_7676);
xor U8245 (N_8245,N_7744,N_7827);
xor U8246 (N_8246,N_7754,N_7586);
nor U8247 (N_8247,N_7963,N_7627);
or U8248 (N_8248,N_7572,N_7829);
xnor U8249 (N_8249,N_7901,N_7927);
xor U8250 (N_8250,N_7738,N_7764);
and U8251 (N_8251,N_7814,N_7836);
and U8252 (N_8252,N_7803,N_7871);
nand U8253 (N_8253,N_7610,N_7978);
or U8254 (N_8254,N_7816,N_7884);
and U8255 (N_8255,N_7760,N_7818);
and U8256 (N_8256,N_7957,N_7847);
or U8257 (N_8257,N_7635,N_7676);
xnor U8258 (N_8258,N_7598,N_7716);
nand U8259 (N_8259,N_7794,N_7693);
xnor U8260 (N_8260,N_7560,N_7936);
nor U8261 (N_8261,N_7738,N_7670);
nor U8262 (N_8262,N_7583,N_7811);
or U8263 (N_8263,N_7701,N_7652);
nand U8264 (N_8264,N_7934,N_7559);
or U8265 (N_8265,N_7502,N_7710);
or U8266 (N_8266,N_7904,N_7794);
nor U8267 (N_8267,N_7644,N_7948);
or U8268 (N_8268,N_7682,N_7957);
nand U8269 (N_8269,N_7752,N_7595);
nor U8270 (N_8270,N_7925,N_7717);
or U8271 (N_8271,N_7978,N_7602);
or U8272 (N_8272,N_7823,N_7779);
and U8273 (N_8273,N_7910,N_7944);
or U8274 (N_8274,N_7796,N_7984);
and U8275 (N_8275,N_7611,N_7804);
xor U8276 (N_8276,N_7835,N_7560);
nor U8277 (N_8277,N_7506,N_7926);
or U8278 (N_8278,N_7969,N_7834);
or U8279 (N_8279,N_7631,N_7922);
xor U8280 (N_8280,N_7658,N_7619);
nand U8281 (N_8281,N_7958,N_7572);
or U8282 (N_8282,N_7620,N_7573);
or U8283 (N_8283,N_7746,N_7962);
nand U8284 (N_8284,N_7501,N_7544);
nor U8285 (N_8285,N_7515,N_7617);
xnor U8286 (N_8286,N_7621,N_7788);
and U8287 (N_8287,N_7897,N_7608);
and U8288 (N_8288,N_7649,N_7705);
nor U8289 (N_8289,N_7770,N_7705);
or U8290 (N_8290,N_7569,N_7760);
xnor U8291 (N_8291,N_7966,N_7882);
nand U8292 (N_8292,N_7636,N_7907);
nor U8293 (N_8293,N_7513,N_7916);
xnor U8294 (N_8294,N_7968,N_7847);
and U8295 (N_8295,N_7757,N_7972);
xnor U8296 (N_8296,N_7945,N_7565);
or U8297 (N_8297,N_7670,N_7768);
nand U8298 (N_8298,N_7609,N_7848);
or U8299 (N_8299,N_7791,N_7539);
nand U8300 (N_8300,N_7929,N_7808);
nand U8301 (N_8301,N_7927,N_7856);
nor U8302 (N_8302,N_7512,N_7620);
xnor U8303 (N_8303,N_7930,N_7823);
and U8304 (N_8304,N_7933,N_7966);
and U8305 (N_8305,N_7948,N_7517);
and U8306 (N_8306,N_7755,N_7589);
nand U8307 (N_8307,N_7892,N_7942);
nor U8308 (N_8308,N_7707,N_7850);
nor U8309 (N_8309,N_7867,N_7724);
and U8310 (N_8310,N_7543,N_7634);
or U8311 (N_8311,N_7712,N_7948);
or U8312 (N_8312,N_7527,N_7845);
and U8313 (N_8313,N_7609,N_7672);
nor U8314 (N_8314,N_7721,N_7653);
and U8315 (N_8315,N_7965,N_7589);
nor U8316 (N_8316,N_7563,N_7695);
or U8317 (N_8317,N_7633,N_7870);
and U8318 (N_8318,N_7538,N_7894);
xor U8319 (N_8319,N_7700,N_7903);
nand U8320 (N_8320,N_7775,N_7888);
and U8321 (N_8321,N_7922,N_7589);
or U8322 (N_8322,N_7617,N_7890);
nand U8323 (N_8323,N_7574,N_7511);
nor U8324 (N_8324,N_7939,N_7512);
xnor U8325 (N_8325,N_7687,N_7517);
and U8326 (N_8326,N_7559,N_7891);
xor U8327 (N_8327,N_7850,N_7692);
xor U8328 (N_8328,N_7681,N_7902);
or U8329 (N_8329,N_7673,N_7747);
nand U8330 (N_8330,N_7763,N_7756);
nor U8331 (N_8331,N_7989,N_7733);
and U8332 (N_8332,N_7868,N_7995);
xnor U8333 (N_8333,N_7568,N_7531);
and U8334 (N_8334,N_7778,N_7657);
nor U8335 (N_8335,N_7919,N_7507);
nor U8336 (N_8336,N_7632,N_7556);
or U8337 (N_8337,N_7783,N_7825);
nand U8338 (N_8338,N_7521,N_7582);
and U8339 (N_8339,N_7738,N_7537);
and U8340 (N_8340,N_7528,N_7870);
or U8341 (N_8341,N_7967,N_7646);
xor U8342 (N_8342,N_7985,N_7946);
nand U8343 (N_8343,N_7779,N_7703);
and U8344 (N_8344,N_7544,N_7840);
nor U8345 (N_8345,N_7555,N_7709);
xor U8346 (N_8346,N_7612,N_7942);
nor U8347 (N_8347,N_7830,N_7629);
xnor U8348 (N_8348,N_7887,N_7944);
xor U8349 (N_8349,N_7664,N_7508);
nand U8350 (N_8350,N_7836,N_7548);
nor U8351 (N_8351,N_7853,N_7944);
and U8352 (N_8352,N_7965,N_7576);
nand U8353 (N_8353,N_7977,N_7965);
nor U8354 (N_8354,N_7502,N_7509);
and U8355 (N_8355,N_7970,N_7772);
nor U8356 (N_8356,N_7792,N_7997);
or U8357 (N_8357,N_7677,N_7999);
nor U8358 (N_8358,N_7792,N_7794);
nand U8359 (N_8359,N_7899,N_7993);
nor U8360 (N_8360,N_7967,N_7580);
and U8361 (N_8361,N_7934,N_7871);
or U8362 (N_8362,N_7564,N_7678);
xor U8363 (N_8363,N_7608,N_7800);
nand U8364 (N_8364,N_7647,N_7619);
or U8365 (N_8365,N_7630,N_7992);
or U8366 (N_8366,N_7929,N_7569);
nor U8367 (N_8367,N_7735,N_7852);
xnor U8368 (N_8368,N_7928,N_7802);
xnor U8369 (N_8369,N_7816,N_7651);
nor U8370 (N_8370,N_7578,N_7894);
and U8371 (N_8371,N_7928,N_7926);
nor U8372 (N_8372,N_7762,N_7998);
xor U8373 (N_8373,N_7734,N_7617);
and U8374 (N_8374,N_7630,N_7575);
and U8375 (N_8375,N_7961,N_7811);
xor U8376 (N_8376,N_7804,N_7976);
or U8377 (N_8377,N_7953,N_7755);
or U8378 (N_8378,N_7987,N_7975);
or U8379 (N_8379,N_7740,N_7634);
xor U8380 (N_8380,N_7989,N_7919);
and U8381 (N_8381,N_7514,N_7948);
and U8382 (N_8382,N_7785,N_7570);
and U8383 (N_8383,N_7953,N_7800);
xor U8384 (N_8384,N_7942,N_7768);
or U8385 (N_8385,N_7596,N_7764);
nand U8386 (N_8386,N_7574,N_7784);
xnor U8387 (N_8387,N_7960,N_7747);
nor U8388 (N_8388,N_7571,N_7945);
and U8389 (N_8389,N_7596,N_7551);
or U8390 (N_8390,N_7794,N_7533);
nand U8391 (N_8391,N_7515,N_7971);
nor U8392 (N_8392,N_7866,N_7983);
nand U8393 (N_8393,N_7794,N_7556);
and U8394 (N_8394,N_7553,N_7551);
xnor U8395 (N_8395,N_7708,N_7777);
nand U8396 (N_8396,N_7552,N_7627);
nand U8397 (N_8397,N_7511,N_7542);
nor U8398 (N_8398,N_7665,N_7635);
and U8399 (N_8399,N_7651,N_7990);
nor U8400 (N_8400,N_7688,N_7948);
or U8401 (N_8401,N_7582,N_7545);
xor U8402 (N_8402,N_7658,N_7698);
or U8403 (N_8403,N_7630,N_7545);
and U8404 (N_8404,N_7609,N_7888);
and U8405 (N_8405,N_7603,N_7914);
xnor U8406 (N_8406,N_7676,N_7970);
and U8407 (N_8407,N_7792,N_7772);
xnor U8408 (N_8408,N_7509,N_7912);
nand U8409 (N_8409,N_7610,N_7965);
or U8410 (N_8410,N_7676,N_7723);
nor U8411 (N_8411,N_7834,N_7868);
xnor U8412 (N_8412,N_7662,N_7837);
and U8413 (N_8413,N_7884,N_7956);
xnor U8414 (N_8414,N_7805,N_7523);
xor U8415 (N_8415,N_7925,N_7602);
and U8416 (N_8416,N_7755,N_7974);
and U8417 (N_8417,N_7861,N_7815);
or U8418 (N_8418,N_7698,N_7504);
and U8419 (N_8419,N_7747,N_7566);
xnor U8420 (N_8420,N_7609,N_7857);
nor U8421 (N_8421,N_7506,N_7970);
nand U8422 (N_8422,N_7563,N_7509);
nand U8423 (N_8423,N_7556,N_7722);
nor U8424 (N_8424,N_7864,N_7878);
or U8425 (N_8425,N_7860,N_7929);
xor U8426 (N_8426,N_7804,N_7951);
and U8427 (N_8427,N_7951,N_7966);
or U8428 (N_8428,N_7886,N_7989);
nand U8429 (N_8429,N_7779,N_7563);
nor U8430 (N_8430,N_7570,N_7660);
nor U8431 (N_8431,N_7784,N_7829);
or U8432 (N_8432,N_7530,N_7982);
nor U8433 (N_8433,N_7914,N_7885);
and U8434 (N_8434,N_7995,N_7807);
nand U8435 (N_8435,N_7684,N_7972);
and U8436 (N_8436,N_7751,N_7961);
nand U8437 (N_8437,N_7582,N_7718);
nor U8438 (N_8438,N_7733,N_7909);
nor U8439 (N_8439,N_7863,N_7549);
nor U8440 (N_8440,N_7821,N_7971);
or U8441 (N_8441,N_7883,N_7816);
or U8442 (N_8442,N_7887,N_7517);
xnor U8443 (N_8443,N_7722,N_7566);
nor U8444 (N_8444,N_7595,N_7538);
nand U8445 (N_8445,N_7807,N_7611);
or U8446 (N_8446,N_7940,N_7875);
nand U8447 (N_8447,N_7552,N_7840);
and U8448 (N_8448,N_7573,N_7731);
xnor U8449 (N_8449,N_7732,N_7886);
nand U8450 (N_8450,N_7729,N_7645);
and U8451 (N_8451,N_7529,N_7576);
nor U8452 (N_8452,N_7937,N_7946);
or U8453 (N_8453,N_7941,N_7707);
xnor U8454 (N_8454,N_7868,N_7773);
xor U8455 (N_8455,N_7649,N_7909);
or U8456 (N_8456,N_7514,N_7614);
xnor U8457 (N_8457,N_7782,N_7541);
or U8458 (N_8458,N_7665,N_7767);
nor U8459 (N_8459,N_7569,N_7627);
xor U8460 (N_8460,N_7672,N_7998);
or U8461 (N_8461,N_7786,N_7884);
nand U8462 (N_8462,N_7607,N_7625);
or U8463 (N_8463,N_7572,N_7824);
xnor U8464 (N_8464,N_7858,N_7931);
nand U8465 (N_8465,N_7896,N_7624);
or U8466 (N_8466,N_7657,N_7590);
xor U8467 (N_8467,N_7635,N_7948);
or U8468 (N_8468,N_7946,N_7641);
xnor U8469 (N_8469,N_7874,N_7501);
xor U8470 (N_8470,N_7856,N_7992);
nand U8471 (N_8471,N_7603,N_7685);
and U8472 (N_8472,N_7915,N_7954);
nand U8473 (N_8473,N_7664,N_7944);
nor U8474 (N_8474,N_7995,N_7840);
xor U8475 (N_8475,N_7900,N_7936);
nand U8476 (N_8476,N_7622,N_7822);
nand U8477 (N_8477,N_7993,N_7579);
and U8478 (N_8478,N_7606,N_7958);
nor U8479 (N_8479,N_7786,N_7803);
or U8480 (N_8480,N_7507,N_7901);
nor U8481 (N_8481,N_7904,N_7568);
nand U8482 (N_8482,N_7729,N_7673);
nor U8483 (N_8483,N_7523,N_7637);
nand U8484 (N_8484,N_7777,N_7798);
or U8485 (N_8485,N_7837,N_7772);
or U8486 (N_8486,N_7621,N_7774);
xnor U8487 (N_8487,N_7512,N_7793);
xnor U8488 (N_8488,N_7660,N_7910);
nand U8489 (N_8489,N_7650,N_7981);
nand U8490 (N_8490,N_7787,N_7812);
or U8491 (N_8491,N_7913,N_7748);
or U8492 (N_8492,N_7510,N_7542);
or U8493 (N_8493,N_7993,N_7759);
nor U8494 (N_8494,N_7610,N_7979);
or U8495 (N_8495,N_7771,N_7641);
nand U8496 (N_8496,N_7636,N_7694);
nand U8497 (N_8497,N_7832,N_7962);
nand U8498 (N_8498,N_7593,N_7927);
nand U8499 (N_8499,N_7533,N_7973);
xnor U8500 (N_8500,N_8183,N_8370);
and U8501 (N_8501,N_8019,N_8084);
nor U8502 (N_8502,N_8016,N_8240);
nand U8503 (N_8503,N_8280,N_8160);
and U8504 (N_8504,N_8281,N_8158);
nor U8505 (N_8505,N_8277,N_8461);
xor U8506 (N_8506,N_8422,N_8418);
nand U8507 (N_8507,N_8327,N_8341);
xor U8508 (N_8508,N_8361,N_8390);
and U8509 (N_8509,N_8484,N_8115);
or U8510 (N_8510,N_8425,N_8362);
xnor U8511 (N_8511,N_8163,N_8437);
or U8512 (N_8512,N_8384,N_8079);
or U8513 (N_8513,N_8460,N_8048);
nor U8514 (N_8514,N_8325,N_8412);
nor U8515 (N_8515,N_8143,N_8347);
or U8516 (N_8516,N_8131,N_8416);
or U8517 (N_8517,N_8231,N_8103);
nor U8518 (N_8518,N_8287,N_8176);
nor U8519 (N_8519,N_8093,N_8100);
and U8520 (N_8520,N_8272,N_8442);
or U8521 (N_8521,N_8132,N_8088);
or U8522 (N_8522,N_8137,N_8085);
nand U8523 (N_8523,N_8128,N_8112);
nor U8524 (N_8524,N_8333,N_8237);
xnor U8525 (N_8525,N_8266,N_8138);
xor U8526 (N_8526,N_8031,N_8056);
nor U8527 (N_8527,N_8166,N_8273);
or U8528 (N_8528,N_8123,N_8499);
or U8529 (N_8529,N_8342,N_8090);
nand U8530 (N_8530,N_8331,N_8365);
or U8531 (N_8531,N_8097,N_8459);
or U8532 (N_8532,N_8409,N_8028);
nor U8533 (N_8533,N_8201,N_8414);
nand U8534 (N_8534,N_8136,N_8044);
xnor U8535 (N_8535,N_8379,N_8117);
and U8536 (N_8536,N_8014,N_8025);
and U8537 (N_8537,N_8336,N_8236);
nor U8538 (N_8538,N_8239,N_8456);
nor U8539 (N_8539,N_8279,N_8076);
and U8540 (N_8540,N_8184,N_8058);
nand U8541 (N_8541,N_8440,N_8434);
xor U8542 (N_8542,N_8039,N_8289);
nand U8543 (N_8543,N_8064,N_8351);
nor U8544 (N_8544,N_8488,N_8151);
nor U8545 (N_8545,N_8145,N_8017);
and U8546 (N_8546,N_8452,N_8400);
nor U8547 (N_8547,N_8135,N_8029);
or U8548 (N_8548,N_8448,N_8062);
and U8549 (N_8549,N_8455,N_8008);
and U8550 (N_8550,N_8405,N_8344);
nor U8551 (N_8551,N_8155,N_8490);
nand U8552 (N_8552,N_8478,N_8492);
or U8553 (N_8553,N_8156,N_8439);
and U8554 (N_8554,N_8330,N_8108);
nor U8555 (N_8555,N_8173,N_8080);
and U8556 (N_8556,N_8253,N_8348);
and U8557 (N_8557,N_8431,N_8116);
or U8558 (N_8558,N_8329,N_8209);
nor U8559 (N_8559,N_8152,N_8495);
or U8560 (N_8560,N_8038,N_8269);
nand U8561 (N_8561,N_8380,N_8335);
nand U8562 (N_8562,N_8377,N_8120);
nor U8563 (N_8563,N_8323,N_8047);
nor U8564 (N_8564,N_8469,N_8319);
nand U8565 (N_8565,N_8105,N_8350);
nand U8566 (N_8566,N_8052,N_8227);
nand U8567 (N_8567,N_8334,N_8352);
nor U8568 (N_8568,N_8095,N_8216);
nand U8569 (N_8569,N_8197,N_8321);
xnor U8570 (N_8570,N_8118,N_8213);
or U8571 (N_8571,N_8394,N_8114);
xnor U8572 (N_8572,N_8177,N_8193);
nand U8573 (N_8573,N_8001,N_8161);
and U8574 (N_8574,N_8376,N_8026);
nand U8575 (N_8575,N_8398,N_8186);
and U8576 (N_8576,N_8003,N_8206);
nor U8577 (N_8577,N_8192,N_8243);
xor U8578 (N_8578,N_8435,N_8067);
and U8579 (N_8579,N_8489,N_8157);
xor U8580 (N_8580,N_8200,N_8312);
and U8581 (N_8581,N_8389,N_8358);
nand U8582 (N_8582,N_8401,N_8444);
nand U8583 (N_8583,N_8104,N_8252);
and U8584 (N_8584,N_8445,N_8109);
nand U8585 (N_8585,N_8170,N_8254);
nand U8586 (N_8586,N_8072,N_8450);
xor U8587 (N_8587,N_8133,N_8018);
and U8588 (N_8588,N_8451,N_8270);
or U8589 (N_8589,N_8395,N_8241);
nand U8590 (N_8590,N_8308,N_8476);
xnor U8591 (N_8591,N_8413,N_8168);
nor U8592 (N_8592,N_8102,N_8147);
or U8593 (N_8593,N_8233,N_8221);
nor U8594 (N_8594,N_8196,N_8436);
nand U8595 (N_8595,N_8260,N_8311);
and U8596 (N_8596,N_8180,N_8055);
or U8597 (N_8597,N_8073,N_8217);
nor U8598 (N_8598,N_8081,N_8144);
nand U8599 (N_8599,N_8122,N_8096);
nor U8600 (N_8600,N_8282,N_8402);
and U8601 (N_8601,N_8393,N_8214);
xnor U8602 (N_8602,N_8089,N_8406);
nand U8603 (N_8603,N_8391,N_8315);
or U8604 (N_8604,N_8367,N_8199);
nor U8605 (N_8605,N_8276,N_8392);
nand U8606 (N_8606,N_8234,N_8245);
and U8607 (N_8607,N_8467,N_8020);
xor U8608 (N_8608,N_8374,N_8487);
nor U8609 (N_8609,N_8433,N_8417);
nand U8610 (N_8610,N_8092,N_8007);
and U8611 (N_8611,N_8320,N_8288);
and U8612 (N_8612,N_8203,N_8043);
xor U8613 (N_8613,N_8346,N_8458);
and U8614 (N_8614,N_8408,N_8332);
nand U8615 (N_8615,N_8212,N_8068);
and U8616 (N_8616,N_8202,N_8054);
or U8617 (N_8617,N_8378,N_8383);
xnor U8618 (N_8618,N_8162,N_8002);
or U8619 (N_8619,N_8283,N_8153);
and U8620 (N_8620,N_8050,N_8441);
or U8621 (N_8621,N_8286,N_8472);
or U8622 (N_8622,N_8185,N_8388);
nor U8623 (N_8623,N_8188,N_8305);
nand U8624 (N_8624,N_8191,N_8264);
or U8625 (N_8625,N_8360,N_8078);
and U8626 (N_8626,N_8204,N_8470);
nand U8627 (N_8627,N_8187,N_8368);
nor U8628 (N_8628,N_8235,N_8310);
nand U8629 (N_8629,N_8284,N_8005);
or U8630 (N_8630,N_8298,N_8317);
and U8631 (N_8631,N_8110,N_8337);
xor U8632 (N_8632,N_8167,N_8290);
xnor U8633 (N_8633,N_8042,N_8396);
or U8634 (N_8634,N_8232,N_8359);
nand U8635 (N_8635,N_8053,N_8485);
nor U8636 (N_8636,N_8000,N_8430);
and U8637 (N_8637,N_8263,N_8009);
nand U8638 (N_8638,N_8195,N_8140);
nor U8639 (N_8639,N_8306,N_8465);
xnor U8640 (N_8640,N_8292,N_8285);
xnor U8641 (N_8641,N_8242,N_8149);
nor U8642 (N_8642,N_8248,N_8424);
or U8643 (N_8643,N_8297,N_8419);
nand U8644 (N_8644,N_8494,N_8210);
or U8645 (N_8645,N_8271,N_8075);
or U8646 (N_8646,N_8011,N_8371);
nand U8647 (N_8647,N_8256,N_8070);
nor U8648 (N_8648,N_8012,N_8190);
nor U8649 (N_8649,N_8318,N_8074);
nand U8650 (N_8650,N_8491,N_8101);
or U8651 (N_8651,N_8345,N_8295);
nor U8652 (N_8652,N_8473,N_8219);
nor U8653 (N_8653,N_8126,N_8246);
or U8654 (N_8654,N_8326,N_8077);
nand U8655 (N_8655,N_8071,N_8420);
nand U8656 (N_8656,N_8322,N_8274);
xor U8657 (N_8657,N_8134,N_8404);
or U8658 (N_8658,N_8159,N_8127);
xnor U8659 (N_8659,N_8015,N_8215);
nor U8660 (N_8660,N_8482,N_8139);
and U8661 (N_8661,N_8293,N_8174);
and U8662 (N_8662,N_8049,N_8010);
or U8663 (N_8663,N_8069,N_8303);
nand U8664 (N_8664,N_8004,N_8498);
or U8665 (N_8665,N_8375,N_8205);
xor U8666 (N_8666,N_8238,N_8294);
nand U8667 (N_8667,N_8033,N_8497);
and U8668 (N_8668,N_8356,N_8363);
and U8669 (N_8669,N_8399,N_8141);
nor U8670 (N_8670,N_8211,N_8429);
nand U8671 (N_8671,N_8182,N_8432);
or U8672 (N_8672,N_8154,N_8421);
nand U8673 (N_8673,N_8449,N_8369);
and U8674 (N_8674,N_8302,N_8423);
nor U8675 (N_8675,N_8453,N_8194);
and U8676 (N_8676,N_8259,N_8354);
and U8677 (N_8677,N_8454,N_8407);
and U8678 (N_8678,N_8148,N_8475);
xor U8679 (N_8679,N_8107,N_8051);
xor U8680 (N_8680,N_8468,N_8258);
nor U8681 (N_8681,N_8098,N_8403);
or U8682 (N_8682,N_8249,N_8471);
nor U8683 (N_8683,N_8316,N_8106);
nor U8684 (N_8684,N_8121,N_8063);
nand U8685 (N_8685,N_8324,N_8113);
or U8686 (N_8686,N_8275,N_8046);
xor U8687 (N_8687,N_8343,N_8129);
nor U8688 (N_8688,N_8481,N_8457);
or U8689 (N_8689,N_8427,N_8304);
or U8690 (N_8690,N_8372,N_8082);
or U8691 (N_8691,N_8385,N_8111);
nor U8692 (N_8692,N_8169,N_8223);
xnor U8693 (N_8693,N_8065,N_8268);
xnor U8694 (N_8694,N_8447,N_8387);
or U8695 (N_8695,N_8066,N_8023);
nor U8696 (N_8696,N_8036,N_8030);
xor U8697 (N_8697,N_8314,N_8338);
and U8698 (N_8698,N_8386,N_8222);
nor U8699 (N_8699,N_8091,N_8267);
and U8700 (N_8700,N_8446,N_8483);
nand U8701 (N_8701,N_8355,N_8037);
nand U8702 (N_8702,N_8045,N_8251);
and U8703 (N_8703,N_8099,N_8124);
nor U8704 (N_8704,N_8443,N_8059);
and U8705 (N_8705,N_8462,N_8299);
nor U8706 (N_8706,N_8171,N_8119);
nor U8707 (N_8707,N_8250,N_8463);
and U8708 (N_8708,N_8340,N_8309);
nand U8709 (N_8709,N_8179,N_8150);
nand U8710 (N_8710,N_8301,N_8230);
or U8711 (N_8711,N_8493,N_8060);
xnor U8712 (N_8712,N_8040,N_8226);
and U8713 (N_8713,N_8130,N_8278);
xnor U8714 (N_8714,N_8415,N_8480);
and U8715 (N_8715,N_8032,N_8428);
xnor U8716 (N_8716,N_8057,N_8027);
and U8717 (N_8717,N_8164,N_8021);
and U8718 (N_8718,N_8041,N_8291);
or U8719 (N_8719,N_8165,N_8486);
or U8720 (N_8720,N_8218,N_8353);
xor U8721 (N_8721,N_8464,N_8208);
nor U8722 (N_8722,N_8366,N_8172);
and U8723 (N_8723,N_8313,N_8328);
and U8724 (N_8724,N_8474,N_8479);
xnor U8725 (N_8725,N_8125,N_8034);
nor U8726 (N_8726,N_8142,N_8296);
nand U8727 (N_8727,N_8220,N_8426);
xor U8728 (N_8728,N_8261,N_8438);
nor U8729 (N_8729,N_8262,N_8265);
or U8730 (N_8730,N_8247,N_8086);
nor U8731 (N_8731,N_8357,N_8229);
nand U8732 (N_8732,N_8224,N_8189);
and U8733 (N_8733,N_8178,N_8207);
nor U8734 (N_8734,N_8339,N_8146);
or U8735 (N_8735,N_8382,N_8255);
nand U8736 (N_8736,N_8300,N_8373);
or U8737 (N_8737,N_8225,N_8198);
nor U8738 (N_8738,N_8410,N_8381);
xnor U8739 (N_8739,N_8228,N_8083);
nand U8740 (N_8740,N_8024,N_8181);
nor U8741 (N_8741,N_8364,N_8477);
or U8742 (N_8742,N_8307,N_8006);
nand U8743 (N_8743,N_8087,N_8061);
nor U8744 (N_8744,N_8244,N_8094);
and U8745 (N_8745,N_8257,N_8349);
xor U8746 (N_8746,N_8035,N_8466);
nor U8747 (N_8747,N_8397,N_8411);
nand U8748 (N_8748,N_8175,N_8022);
nand U8749 (N_8749,N_8496,N_8013);
nor U8750 (N_8750,N_8283,N_8001);
nor U8751 (N_8751,N_8153,N_8009);
and U8752 (N_8752,N_8302,N_8341);
xor U8753 (N_8753,N_8160,N_8017);
nand U8754 (N_8754,N_8267,N_8052);
nor U8755 (N_8755,N_8124,N_8424);
nand U8756 (N_8756,N_8333,N_8425);
nand U8757 (N_8757,N_8487,N_8457);
and U8758 (N_8758,N_8328,N_8017);
nor U8759 (N_8759,N_8230,N_8270);
nor U8760 (N_8760,N_8169,N_8106);
or U8761 (N_8761,N_8050,N_8467);
nor U8762 (N_8762,N_8035,N_8471);
xnor U8763 (N_8763,N_8351,N_8335);
nor U8764 (N_8764,N_8070,N_8254);
xor U8765 (N_8765,N_8230,N_8434);
nand U8766 (N_8766,N_8186,N_8239);
and U8767 (N_8767,N_8167,N_8111);
or U8768 (N_8768,N_8277,N_8294);
nand U8769 (N_8769,N_8354,N_8283);
or U8770 (N_8770,N_8252,N_8256);
or U8771 (N_8771,N_8139,N_8420);
nor U8772 (N_8772,N_8147,N_8136);
or U8773 (N_8773,N_8173,N_8268);
nand U8774 (N_8774,N_8064,N_8156);
and U8775 (N_8775,N_8382,N_8102);
and U8776 (N_8776,N_8431,N_8290);
and U8777 (N_8777,N_8271,N_8360);
or U8778 (N_8778,N_8210,N_8451);
or U8779 (N_8779,N_8181,N_8306);
nand U8780 (N_8780,N_8095,N_8249);
or U8781 (N_8781,N_8161,N_8137);
nand U8782 (N_8782,N_8285,N_8073);
nand U8783 (N_8783,N_8484,N_8240);
and U8784 (N_8784,N_8463,N_8262);
or U8785 (N_8785,N_8455,N_8146);
nor U8786 (N_8786,N_8336,N_8118);
and U8787 (N_8787,N_8306,N_8498);
xnor U8788 (N_8788,N_8155,N_8277);
nor U8789 (N_8789,N_8286,N_8186);
or U8790 (N_8790,N_8347,N_8454);
nand U8791 (N_8791,N_8196,N_8240);
or U8792 (N_8792,N_8006,N_8270);
nand U8793 (N_8793,N_8195,N_8079);
xor U8794 (N_8794,N_8145,N_8438);
or U8795 (N_8795,N_8209,N_8249);
xnor U8796 (N_8796,N_8187,N_8149);
or U8797 (N_8797,N_8153,N_8106);
and U8798 (N_8798,N_8321,N_8490);
and U8799 (N_8799,N_8440,N_8484);
and U8800 (N_8800,N_8396,N_8364);
nand U8801 (N_8801,N_8489,N_8220);
xor U8802 (N_8802,N_8367,N_8413);
and U8803 (N_8803,N_8283,N_8180);
nand U8804 (N_8804,N_8417,N_8333);
nor U8805 (N_8805,N_8060,N_8007);
xor U8806 (N_8806,N_8154,N_8422);
nand U8807 (N_8807,N_8126,N_8444);
and U8808 (N_8808,N_8467,N_8234);
nand U8809 (N_8809,N_8043,N_8318);
nor U8810 (N_8810,N_8310,N_8427);
nor U8811 (N_8811,N_8235,N_8473);
nand U8812 (N_8812,N_8140,N_8158);
nor U8813 (N_8813,N_8486,N_8281);
or U8814 (N_8814,N_8375,N_8301);
nand U8815 (N_8815,N_8259,N_8322);
xor U8816 (N_8816,N_8459,N_8465);
and U8817 (N_8817,N_8228,N_8423);
nor U8818 (N_8818,N_8306,N_8180);
nor U8819 (N_8819,N_8367,N_8118);
nand U8820 (N_8820,N_8132,N_8033);
nor U8821 (N_8821,N_8021,N_8117);
or U8822 (N_8822,N_8090,N_8002);
and U8823 (N_8823,N_8166,N_8463);
and U8824 (N_8824,N_8078,N_8328);
or U8825 (N_8825,N_8165,N_8094);
or U8826 (N_8826,N_8479,N_8068);
and U8827 (N_8827,N_8403,N_8226);
nand U8828 (N_8828,N_8312,N_8005);
or U8829 (N_8829,N_8091,N_8436);
nor U8830 (N_8830,N_8257,N_8348);
nand U8831 (N_8831,N_8261,N_8322);
and U8832 (N_8832,N_8460,N_8058);
and U8833 (N_8833,N_8141,N_8077);
or U8834 (N_8834,N_8248,N_8267);
xnor U8835 (N_8835,N_8365,N_8013);
xnor U8836 (N_8836,N_8417,N_8350);
nor U8837 (N_8837,N_8307,N_8348);
or U8838 (N_8838,N_8426,N_8427);
and U8839 (N_8839,N_8445,N_8288);
nor U8840 (N_8840,N_8382,N_8433);
nor U8841 (N_8841,N_8350,N_8377);
nor U8842 (N_8842,N_8137,N_8017);
or U8843 (N_8843,N_8211,N_8103);
nand U8844 (N_8844,N_8458,N_8135);
nor U8845 (N_8845,N_8316,N_8197);
and U8846 (N_8846,N_8210,N_8215);
nor U8847 (N_8847,N_8496,N_8371);
and U8848 (N_8848,N_8409,N_8287);
or U8849 (N_8849,N_8263,N_8316);
or U8850 (N_8850,N_8005,N_8376);
nor U8851 (N_8851,N_8255,N_8309);
and U8852 (N_8852,N_8441,N_8103);
or U8853 (N_8853,N_8427,N_8476);
and U8854 (N_8854,N_8243,N_8139);
xnor U8855 (N_8855,N_8132,N_8438);
or U8856 (N_8856,N_8455,N_8151);
xnor U8857 (N_8857,N_8164,N_8377);
xor U8858 (N_8858,N_8045,N_8212);
nor U8859 (N_8859,N_8255,N_8139);
xnor U8860 (N_8860,N_8312,N_8125);
xor U8861 (N_8861,N_8100,N_8027);
or U8862 (N_8862,N_8320,N_8469);
nand U8863 (N_8863,N_8293,N_8455);
and U8864 (N_8864,N_8477,N_8376);
nor U8865 (N_8865,N_8271,N_8349);
and U8866 (N_8866,N_8326,N_8293);
or U8867 (N_8867,N_8485,N_8288);
and U8868 (N_8868,N_8258,N_8094);
nand U8869 (N_8869,N_8160,N_8103);
and U8870 (N_8870,N_8434,N_8346);
xnor U8871 (N_8871,N_8479,N_8173);
or U8872 (N_8872,N_8284,N_8387);
nand U8873 (N_8873,N_8029,N_8272);
nand U8874 (N_8874,N_8478,N_8112);
xor U8875 (N_8875,N_8250,N_8148);
nor U8876 (N_8876,N_8048,N_8118);
nor U8877 (N_8877,N_8326,N_8069);
xnor U8878 (N_8878,N_8307,N_8075);
xor U8879 (N_8879,N_8200,N_8252);
and U8880 (N_8880,N_8218,N_8298);
nand U8881 (N_8881,N_8340,N_8431);
and U8882 (N_8882,N_8151,N_8436);
nand U8883 (N_8883,N_8374,N_8207);
xnor U8884 (N_8884,N_8388,N_8068);
nor U8885 (N_8885,N_8292,N_8052);
and U8886 (N_8886,N_8161,N_8099);
or U8887 (N_8887,N_8067,N_8068);
or U8888 (N_8888,N_8157,N_8178);
nor U8889 (N_8889,N_8335,N_8127);
nand U8890 (N_8890,N_8323,N_8383);
nand U8891 (N_8891,N_8279,N_8278);
and U8892 (N_8892,N_8007,N_8067);
and U8893 (N_8893,N_8135,N_8339);
xnor U8894 (N_8894,N_8106,N_8107);
or U8895 (N_8895,N_8397,N_8359);
xor U8896 (N_8896,N_8110,N_8340);
nor U8897 (N_8897,N_8005,N_8222);
and U8898 (N_8898,N_8131,N_8087);
xor U8899 (N_8899,N_8037,N_8201);
or U8900 (N_8900,N_8156,N_8412);
and U8901 (N_8901,N_8156,N_8079);
nor U8902 (N_8902,N_8024,N_8084);
or U8903 (N_8903,N_8020,N_8147);
and U8904 (N_8904,N_8243,N_8461);
nand U8905 (N_8905,N_8452,N_8448);
nor U8906 (N_8906,N_8464,N_8395);
nand U8907 (N_8907,N_8327,N_8063);
nand U8908 (N_8908,N_8362,N_8013);
nor U8909 (N_8909,N_8410,N_8267);
nor U8910 (N_8910,N_8332,N_8229);
or U8911 (N_8911,N_8173,N_8017);
and U8912 (N_8912,N_8167,N_8068);
nor U8913 (N_8913,N_8243,N_8208);
and U8914 (N_8914,N_8030,N_8022);
nand U8915 (N_8915,N_8051,N_8433);
xor U8916 (N_8916,N_8288,N_8167);
xnor U8917 (N_8917,N_8128,N_8333);
or U8918 (N_8918,N_8099,N_8356);
nor U8919 (N_8919,N_8390,N_8220);
nand U8920 (N_8920,N_8077,N_8404);
and U8921 (N_8921,N_8135,N_8315);
nor U8922 (N_8922,N_8237,N_8345);
xnor U8923 (N_8923,N_8078,N_8226);
or U8924 (N_8924,N_8168,N_8126);
nand U8925 (N_8925,N_8342,N_8367);
or U8926 (N_8926,N_8021,N_8082);
nand U8927 (N_8927,N_8301,N_8132);
xnor U8928 (N_8928,N_8355,N_8017);
nand U8929 (N_8929,N_8449,N_8119);
nor U8930 (N_8930,N_8150,N_8277);
xnor U8931 (N_8931,N_8363,N_8033);
xnor U8932 (N_8932,N_8255,N_8200);
nor U8933 (N_8933,N_8045,N_8345);
nor U8934 (N_8934,N_8373,N_8377);
nor U8935 (N_8935,N_8214,N_8043);
nand U8936 (N_8936,N_8028,N_8233);
nor U8937 (N_8937,N_8476,N_8411);
xor U8938 (N_8938,N_8032,N_8415);
and U8939 (N_8939,N_8007,N_8075);
or U8940 (N_8940,N_8374,N_8110);
or U8941 (N_8941,N_8051,N_8461);
nor U8942 (N_8942,N_8413,N_8462);
nand U8943 (N_8943,N_8404,N_8186);
or U8944 (N_8944,N_8225,N_8141);
nand U8945 (N_8945,N_8125,N_8196);
xnor U8946 (N_8946,N_8141,N_8307);
nand U8947 (N_8947,N_8378,N_8314);
nor U8948 (N_8948,N_8404,N_8046);
nand U8949 (N_8949,N_8163,N_8182);
xnor U8950 (N_8950,N_8294,N_8115);
or U8951 (N_8951,N_8419,N_8030);
nand U8952 (N_8952,N_8173,N_8420);
and U8953 (N_8953,N_8050,N_8279);
nand U8954 (N_8954,N_8381,N_8175);
nor U8955 (N_8955,N_8031,N_8210);
xor U8956 (N_8956,N_8129,N_8153);
and U8957 (N_8957,N_8162,N_8132);
or U8958 (N_8958,N_8066,N_8239);
nand U8959 (N_8959,N_8499,N_8188);
nor U8960 (N_8960,N_8431,N_8346);
or U8961 (N_8961,N_8370,N_8347);
xnor U8962 (N_8962,N_8005,N_8341);
and U8963 (N_8963,N_8244,N_8089);
and U8964 (N_8964,N_8210,N_8200);
and U8965 (N_8965,N_8263,N_8254);
nand U8966 (N_8966,N_8187,N_8225);
and U8967 (N_8967,N_8043,N_8339);
nand U8968 (N_8968,N_8392,N_8376);
nand U8969 (N_8969,N_8115,N_8106);
nand U8970 (N_8970,N_8009,N_8092);
xor U8971 (N_8971,N_8334,N_8128);
nand U8972 (N_8972,N_8148,N_8017);
xnor U8973 (N_8973,N_8198,N_8181);
nand U8974 (N_8974,N_8288,N_8137);
or U8975 (N_8975,N_8238,N_8227);
xnor U8976 (N_8976,N_8486,N_8102);
nor U8977 (N_8977,N_8002,N_8246);
nor U8978 (N_8978,N_8132,N_8418);
nor U8979 (N_8979,N_8299,N_8309);
or U8980 (N_8980,N_8070,N_8152);
or U8981 (N_8981,N_8028,N_8323);
and U8982 (N_8982,N_8166,N_8070);
or U8983 (N_8983,N_8090,N_8134);
xnor U8984 (N_8984,N_8080,N_8018);
nor U8985 (N_8985,N_8318,N_8258);
and U8986 (N_8986,N_8122,N_8172);
or U8987 (N_8987,N_8047,N_8199);
nor U8988 (N_8988,N_8039,N_8228);
or U8989 (N_8989,N_8229,N_8237);
or U8990 (N_8990,N_8364,N_8043);
or U8991 (N_8991,N_8011,N_8490);
and U8992 (N_8992,N_8339,N_8057);
and U8993 (N_8993,N_8487,N_8123);
nor U8994 (N_8994,N_8359,N_8054);
or U8995 (N_8995,N_8016,N_8001);
and U8996 (N_8996,N_8198,N_8032);
or U8997 (N_8997,N_8235,N_8248);
and U8998 (N_8998,N_8387,N_8193);
xor U8999 (N_8999,N_8051,N_8392);
and U9000 (N_9000,N_8806,N_8925);
nand U9001 (N_9001,N_8669,N_8729);
nor U9002 (N_9002,N_8767,N_8510);
xnor U9003 (N_9003,N_8962,N_8550);
or U9004 (N_9004,N_8682,N_8737);
xnor U9005 (N_9005,N_8952,N_8526);
or U9006 (N_9006,N_8829,N_8919);
nand U9007 (N_9007,N_8522,N_8882);
and U9008 (N_9008,N_8553,N_8556);
nand U9009 (N_9009,N_8921,N_8643);
xnor U9010 (N_9010,N_8817,N_8613);
nand U9011 (N_9011,N_8527,N_8726);
and U9012 (N_9012,N_8579,N_8740);
and U9013 (N_9013,N_8695,N_8838);
nor U9014 (N_9014,N_8834,N_8936);
or U9015 (N_9015,N_8886,N_8532);
nand U9016 (N_9016,N_8575,N_8990);
nand U9017 (N_9017,N_8754,N_8803);
and U9018 (N_9018,N_8753,N_8612);
nor U9019 (N_9019,N_8694,N_8582);
or U9020 (N_9020,N_8800,N_8667);
xor U9021 (N_9021,N_8988,N_8614);
and U9022 (N_9022,N_8734,N_8622);
nand U9023 (N_9023,N_8965,N_8585);
or U9024 (N_9024,N_8616,N_8648);
xor U9025 (N_9025,N_8996,N_8552);
or U9026 (N_9026,N_8787,N_8948);
nand U9027 (N_9027,N_8647,N_8914);
nor U9028 (N_9028,N_8673,N_8619);
or U9029 (N_9029,N_8814,N_8644);
and U9030 (N_9030,N_8594,N_8651);
nor U9031 (N_9031,N_8560,N_8650);
and U9032 (N_9032,N_8720,N_8781);
xor U9033 (N_9033,N_8958,N_8696);
nand U9034 (N_9034,N_8758,N_8777);
xnor U9035 (N_9035,N_8653,N_8601);
and U9036 (N_9036,N_8769,N_8828);
and U9037 (N_9037,N_8702,N_8946);
xor U9038 (N_9038,N_8706,N_8540);
nand U9039 (N_9039,N_8855,N_8507);
nand U9040 (N_9040,N_8813,N_8779);
xor U9041 (N_9041,N_8799,N_8693);
nand U9042 (N_9042,N_8700,N_8699);
or U9043 (N_9043,N_8608,N_8891);
and U9044 (N_9044,N_8609,N_8991);
nand U9045 (N_9045,N_8606,N_8785);
xor U9046 (N_9046,N_8853,N_8519);
nor U9047 (N_9047,N_8501,N_8536);
and U9048 (N_9048,N_8557,N_8618);
nand U9049 (N_9049,N_8620,N_8827);
or U9050 (N_9050,N_8697,N_8820);
or U9051 (N_9051,N_8658,N_8857);
and U9052 (N_9052,N_8610,N_8636);
and U9053 (N_9053,N_8561,N_8551);
nand U9054 (N_9054,N_8583,N_8851);
xor U9055 (N_9055,N_8905,N_8535);
or U9056 (N_9056,N_8595,N_8832);
and U9057 (N_9057,N_8778,N_8796);
xor U9058 (N_9058,N_8877,N_8733);
nand U9059 (N_9059,N_8854,N_8816);
and U9060 (N_9060,N_8562,N_8591);
nor U9061 (N_9061,N_8587,N_8748);
and U9062 (N_9062,N_8548,N_8961);
nor U9063 (N_9063,N_8727,N_8752);
or U9064 (N_9064,N_8791,N_8933);
xor U9065 (N_9065,N_8987,N_8892);
or U9066 (N_9066,N_8964,N_8843);
or U9067 (N_9067,N_8626,N_8711);
nand U9068 (N_9068,N_8995,N_8874);
or U9069 (N_9069,N_8760,N_8804);
nor U9070 (N_9070,N_8588,N_8980);
and U9071 (N_9071,N_8528,N_8631);
and U9072 (N_9072,N_8633,N_8662);
or U9073 (N_9073,N_8652,N_8683);
nand U9074 (N_9074,N_8848,N_8703);
and U9075 (N_9075,N_8978,N_8634);
nor U9076 (N_9076,N_8539,N_8504);
or U9077 (N_9077,N_8993,N_8811);
xnor U9078 (N_9078,N_8934,N_8768);
nand U9079 (N_9079,N_8704,N_8598);
nor U9080 (N_9080,N_8688,N_8516);
nand U9081 (N_9081,N_8765,N_8661);
xnor U9082 (N_9082,N_8833,N_8543);
nand U9083 (N_9083,N_8564,N_8969);
or U9084 (N_9084,N_8782,N_8932);
or U9085 (N_9085,N_8549,N_8523);
nor U9086 (N_9086,N_8982,N_8736);
xnor U9087 (N_9087,N_8893,N_8937);
nor U9088 (N_9088,N_8502,N_8907);
nand U9089 (N_9089,N_8596,N_8705);
nor U9090 (N_9090,N_8685,N_8773);
xnor U9091 (N_9091,N_8847,N_8865);
xor U9092 (N_9092,N_8590,N_8567);
and U9093 (N_9093,N_8617,N_8698);
or U9094 (N_9094,N_8917,N_8846);
and U9095 (N_9095,N_8898,N_8538);
nor U9096 (N_9096,N_8565,N_8772);
nor U9097 (N_9097,N_8534,N_8895);
and U9098 (N_9098,N_8568,N_8750);
nor U9099 (N_9099,N_8862,N_8655);
nor U9100 (N_9100,N_8708,N_8666);
and U9101 (N_9101,N_8623,N_8544);
or U9102 (N_9102,N_8597,N_8656);
and U9103 (N_9103,N_8860,N_8569);
or U9104 (N_9104,N_8629,N_8878);
nor U9105 (N_9105,N_8639,N_8805);
xnor U9106 (N_9106,N_8976,N_8869);
xor U9107 (N_9107,N_8784,N_8716);
nor U9108 (N_9108,N_8863,N_8979);
and U9109 (N_9109,N_8665,N_8554);
nor U9110 (N_9110,N_8624,N_8795);
or U9111 (N_9111,N_8837,N_8889);
or U9112 (N_9112,N_8566,N_8867);
nor U9113 (N_9113,N_8722,N_8581);
xnor U9114 (N_9114,N_8941,N_8732);
or U9115 (N_9115,N_8676,N_8763);
xor U9116 (N_9116,N_8728,N_8984);
and U9117 (N_9117,N_8738,N_8635);
xor U9118 (N_9118,N_8992,N_8592);
and U9119 (N_9119,N_8967,N_8576);
nand U9120 (N_9120,N_8894,N_8972);
or U9121 (N_9121,N_8999,N_8808);
nor U9122 (N_9122,N_8928,N_8835);
nand U9123 (N_9123,N_8850,N_8640);
xor U9124 (N_9124,N_8599,N_8500);
nor U9125 (N_9125,N_8951,N_8807);
and U9126 (N_9126,N_8646,N_8884);
nor U9127 (N_9127,N_8718,N_8953);
nand U9128 (N_9128,N_8517,N_8775);
nor U9129 (N_9129,N_8824,N_8801);
or U9130 (N_9130,N_8896,N_8836);
or U9131 (N_9131,N_8637,N_8723);
and U9132 (N_9132,N_8611,N_8783);
or U9133 (N_9133,N_8710,N_8989);
nand U9134 (N_9134,N_8881,N_8657);
and U9135 (N_9135,N_8915,N_8920);
nor U9136 (N_9136,N_8842,N_8521);
xor U9137 (N_9137,N_8981,N_8947);
and U9138 (N_9138,N_8998,N_8674);
xnor U9139 (N_9139,N_8849,N_8844);
and U9140 (N_9140,N_8687,N_8959);
or U9141 (N_9141,N_8861,N_8963);
and U9142 (N_9142,N_8840,N_8970);
nor U9143 (N_9143,N_8714,N_8912);
and U9144 (N_9144,N_8715,N_8717);
nand U9145 (N_9145,N_8883,N_8830);
and U9146 (N_9146,N_8759,N_8638);
nor U9147 (N_9147,N_8515,N_8997);
nor U9148 (N_9148,N_8600,N_8770);
or U9149 (N_9149,N_8913,N_8764);
xor U9150 (N_9150,N_8577,N_8712);
and U9151 (N_9151,N_8621,N_8537);
nor U9152 (N_9152,N_8572,N_8871);
nand U9153 (N_9153,N_8880,N_8529);
and U9154 (N_9154,N_8985,N_8627);
nor U9155 (N_9155,N_8918,N_8812);
xnor U9156 (N_9156,N_8823,N_8939);
nand U9157 (N_9157,N_8686,N_8745);
xor U9158 (N_9158,N_8931,N_8776);
xnor U9159 (N_9159,N_8868,N_8821);
xnor U9160 (N_9160,N_8902,N_8659);
nand U9161 (N_9161,N_8520,N_8794);
nor U9162 (N_9162,N_8604,N_8671);
xnor U9163 (N_9163,N_8731,N_8692);
nand U9164 (N_9164,N_8899,N_8940);
and U9165 (N_9165,N_8825,N_8739);
nor U9166 (N_9166,N_8873,N_8766);
and U9167 (N_9167,N_8761,N_8815);
or U9168 (N_9168,N_8690,N_8910);
xnor U9169 (N_9169,N_8788,N_8802);
or U9170 (N_9170,N_8573,N_8742);
xnor U9171 (N_9171,N_8872,N_8542);
nor U9172 (N_9172,N_8906,N_8904);
or U9173 (N_9173,N_8818,N_8831);
nor U9174 (N_9174,N_8935,N_8689);
nor U9175 (N_9175,N_8945,N_8663);
xor U9176 (N_9176,N_8681,N_8555);
xor U9177 (N_9177,N_8649,N_8675);
xnor U9178 (N_9178,N_8743,N_8508);
nand U9179 (N_9179,N_8615,N_8533);
or U9180 (N_9180,N_8839,N_8879);
nor U9181 (N_9181,N_8509,N_8645);
and U9182 (N_9182,N_8810,N_8747);
xor U9183 (N_9183,N_8589,N_8870);
xor U9184 (N_9184,N_8574,N_8943);
nand U9185 (N_9185,N_8672,N_8630);
xnor U9186 (N_9186,N_8744,N_8927);
xnor U9187 (N_9187,N_8680,N_8797);
or U9188 (N_9188,N_8709,N_8664);
xnor U9189 (N_9189,N_8513,N_8809);
and U9190 (N_9190,N_8570,N_8930);
xnor U9191 (N_9191,N_8563,N_8875);
nand U9192 (N_9192,N_8819,N_8684);
or U9193 (N_9193,N_8789,N_8793);
nor U9194 (N_9194,N_8841,N_8559);
and U9195 (N_9195,N_8571,N_8713);
or U9196 (N_9196,N_8580,N_8960);
xor U9197 (N_9197,N_8909,N_8746);
or U9198 (N_9198,N_8603,N_8944);
or U9199 (N_9199,N_8955,N_8957);
and U9200 (N_9200,N_8668,N_8774);
or U9201 (N_9201,N_8890,N_8950);
xnor U9202 (N_9202,N_8654,N_8798);
nor U9203 (N_9203,N_8701,N_8975);
xor U9204 (N_9204,N_8751,N_8670);
nand U9205 (N_9205,N_8558,N_8923);
and U9206 (N_9206,N_8911,N_8924);
and U9207 (N_9207,N_8605,N_8628);
nor U9208 (N_9208,N_8792,N_8983);
xor U9209 (N_9209,N_8578,N_8586);
or U9210 (N_9210,N_8531,N_8505);
and U9211 (N_9211,N_8771,N_8790);
xnor U9212 (N_9212,N_8584,N_8786);
and U9213 (N_9213,N_8660,N_8942);
or U9214 (N_9214,N_8625,N_8900);
nor U9215 (N_9215,N_8922,N_8547);
xnor U9216 (N_9216,N_8721,N_8954);
nor U9217 (N_9217,N_8929,N_8525);
and U9218 (N_9218,N_8977,N_8741);
and U9219 (N_9219,N_8506,N_8887);
and U9220 (N_9220,N_8719,N_8524);
nand U9221 (N_9221,N_8677,N_8897);
or U9222 (N_9222,N_8749,N_8546);
and U9223 (N_9223,N_8974,N_8757);
and U9224 (N_9224,N_8949,N_8724);
or U9225 (N_9225,N_8762,N_8916);
nand U9226 (N_9226,N_8971,N_8885);
and U9227 (N_9227,N_8530,N_8903);
nand U9228 (N_9228,N_8514,N_8780);
nand U9229 (N_9229,N_8901,N_8966);
nand U9230 (N_9230,N_8956,N_8973);
or U9231 (N_9231,N_8679,N_8691);
nand U9232 (N_9232,N_8642,N_8826);
xnor U9233 (N_9233,N_8876,N_8756);
xor U9234 (N_9234,N_8908,N_8602);
or U9235 (N_9235,N_8730,N_8503);
nor U9236 (N_9236,N_8822,N_8607);
or U9237 (N_9237,N_8545,N_8968);
or U9238 (N_9238,N_8845,N_8866);
nor U9239 (N_9239,N_8541,N_8707);
and U9240 (N_9240,N_8678,N_8725);
or U9241 (N_9241,N_8994,N_8859);
nand U9242 (N_9242,N_8852,N_8938);
nand U9243 (N_9243,N_8593,N_8518);
or U9244 (N_9244,N_8632,N_8986);
nor U9245 (N_9245,N_8858,N_8641);
or U9246 (N_9246,N_8888,N_8511);
nor U9247 (N_9247,N_8856,N_8512);
xnor U9248 (N_9248,N_8926,N_8755);
and U9249 (N_9249,N_8864,N_8735);
or U9250 (N_9250,N_8623,N_8860);
nand U9251 (N_9251,N_8859,N_8610);
nand U9252 (N_9252,N_8970,N_8697);
and U9253 (N_9253,N_8699,N_8867);
or U9254 (N_9254,N_8958,N_8806);
xnor U9255 (N_9255,N_8744,N_8930);
nor U9256 (N_9256,N_8678,N_8943);
xor U9257 (N_9257,N_8841,N_8962);
xnor U9258 (N_9258,N_8526,N_8620);
and U9259 (N_9259,N_8875,N_8853);
or U9260 (N_9260,N_8645,N_8836);
nand U9261 (N_9261,N_8787,N_8500);
or U9262 (N_9262,N_8686,N_8878);
nor U9263 (N_9263,N_8829,N_8931);
nor U9264 (N_9264,N_8804,N_8797);
nand U9265 (N_9265,N_8580,N_8875);
and U9266 (N_9266,N_8912,N_8553);
or U9267 (N_9267,N_8688,N_8832);
and U9268 (N_9268,N_8797,N_8627);
and U9269 (N_9269,N_8998,N_8578);
xnor U9270 (N_9270,N_8838,N_8983);
xor U9271 (N_9271,N_8884,N_8986);
or U9272 (N_9272,N_8584,N_8620);
nor U9273 (N_9273,N_8885,N_8528);
and U9274 (N_9274,N_8826,N_8991);
nand U9275 (N_9275,N_8935,N_8546);
nand U9276 (N_9276,N_8538,N_8722);
or U9277 (N_9277,N_8686,N_8940);
or U9278 (N_9278,N_8938,N_8755);
xnor U9279 (N_9279,N_8823,N_8866);
xnor U9280 (N_9280,N_8643,N_8967);
or U9281 (N_9281,N_8711,N_8927);
xor U9282 (N_9282,N_8880,N_8686);
nand U9283 (N_9283,N_8797,N_8559);
nand U9284 (N_9284,N_8846,N_8797);
nor U9285 (N_9285,N_8591,N_8821);
nor U9286 (N_9286,N_8547,N_8726);
or U9287 (N_9287,N_8588,N_8841);
nand U9288 (N_9288,N_8886,N_8598);
and U9289 (N_9289,N_8513,N_8998);
nand U9290 (N_9290,N_8667,N_8611);
xor U9291 (N_9291,N_8876,N_8755);
nor U9292 (N_9292,N_8662,N_8880);
or U9293 (N_9293,N_8642,N_8853);
nor U9294 (N_9294,N_8581,N_8735);
nand U9295 (N_9295,N_8875,N_8543);
nor U9296 (N_9296,N_8778,N_8934);
nor U9297 (N_9297,N_8980,N_8705);
nor U9298 (N_9298,N_8548,N_8594);
or U9299 (N_9299,N_8801,N_8853);
and U9300 (N_9300,N_8912,N_8781);
nor U9301 (N_9301,N_8596,N_8773);
or U9302 (N_9302,N_8737,N_8824);
or U9303 (N_9303,N_8601,N_8702);
xor U9304 (N_9304,N_8787,N_8946);
nor U9305 (N_9305,N_8956,N_8627);
xnor U9306 (N_9306,N_8677,N_8575);
nor U9307 (N_9307,N_8806,N_8599);
nor U9308 (N_9308,N_8917,N_8630);
or U9309 (N_9309,N_8981,N_8938);
or U9310 (N_9310,N_8650,N_8776);
or U9311 (N_9311,N_8528,N_8923);
nor U9312 (N_9312,N_8719,N_8699);
xor U9313 (N_9313,N_8556,N_8604);
nand U9314 (N_9314,N_8560,N_8641);
nor U9315 (N_9315,N_8819,N_8573);
or U9316 (N_9316,N_8862,N_8734);
nand U9317 (N_9317,N_8529,N_8543);
or U9318 (N_9318,N_8844,N_8583);
or U9319 (N_9319,N_8952,N_8741);
and U9320 (N_9320,N_8539,N_8895);
xor U9321 (N_9321,N_8889,N_8815);
or U9322 (N_9322,N_8791,N_8780);
xor U9323 (N_9323,N_8966,N_8505);
xor U9324 (N_9324,N_8509,N_8834);
nor U9325 (N_9325,N_8747,N_8886);
and U9326 (N_9326,N_8680,N_8735);
or U9327 (N_9327,N_8749,N_8658);
nand U9328 (N_9328,N_8992,N_8524);
or U9329 (N_9329,N_8735,N_8628);
and U9330 (N_9330,N_8617,N_8857);
or U9331 (N_9331,N_8922,N_8821);
nand U9332 (N_9332,N_8974,N_8580);
or U9333 (N_9333,N_8955,N_8842);
or U9334 (N_9334,N_8849,N_8720);
xor U9335 (N_9335,N_8516,N_8693);
nor U9336 (N_9336,N_8862,N_8972);
xor U9337 (N_9337,N_8862,N_8855);
nand U9338 (N_9338,N_8529,N_8995);
xnor U9339 (N_9339,N_8534,N_8762);
or U9340 (N_9340,N_8930,N_8786);
xor U9341 (N_9341,N_8929,N_8753);
nor U9342 (N_9342,N_8847,N_8551);
nand U9343 (N_9343,N_8637,N_8737);
nor U9344 (N_9344,N_8665,N_8817);
and U9345 (N_9345,N_8938,N_8614);
or U9346 (N_9346,N_8916,N_8744);
nor U9347 (N_9347,N_8841,N_8783);
xnor U9348 (N_9348,N_8666,N_8514);
nand U9349 (N_9349,N_8550,N_8872);
xor U9350 (N_9350,N_8906,N_8741);
or U9351 (N_9351,N_8692,N_8591);
and U9352 (N_9352,N_8838,N_8675);
xor U9353 (N_9353,N_8588,N_8883);
and U9354 (N_9354,N_8536,N_8649);
xor U9355 (N_9355,N_8592,N_8713);
xnor U9356 (N_9356,N_8959,N_8520);
and U9357 (N_9357,N_8994,N_8739);
nor U9358 (N_9358,N_8887,N_8564);
and U9359 (N_9359,N_8744,N_8685);
xnor U9360 (N_9360,N_8823,N_8736);
and U9361 (N_9361,N_8535,N_8599);
nand U9362 (N_9362,N_8546,N_8900);
nand U9363 (N_9363,N_8519,N_8788);
or U9364 (N_9364,N_8689,N_8616);
and U9365 (N_9365,N_8542,N_8771);
nand U9366 (N_9366,N_8600,N_8604);
nand U9367 (N_9367,N_8791,N_8915);
and U9368 (N_9368,N_8770,N_8740);
nor U9369 (N_9369,N_8629,N_8660);
nor U9370 (N_9370,N_8839,N_8608);
and U9371 (N_9371,N_8964,N_8986);
or U9372 (N_9372,N_8679,N_8641);
and U9373 (N_9373,N_8776,N_8535);
nor U9374 (N_9374,N_8792,N_8752);
or U9375 (N_9375,N_8768,N_8908);
and U9376 (N_9376,N_8565,N_8931);
nor U9377 (N_9377,N_8659,N_8737);
nand U9378 (N_9378,N_8787,N_8589);
nor U9379 (N_9379,N_8678,N_8669);
or U9380 (N_9380,N_8876,N_8618);
nand U9381 (N_9381,N_8719,N_8662);
or U9382 (N_9382,N_8886,N_8722);
and U9383 (N_9383,N_8569,N_8570);
xnor U9384 (N_9384,N_8574,N_8511);
or U9385 (N_9385,N_8512,N_8511);
and U9386 (N_9386,N_8975,N_8681);
or U9387 (N_9387,N_8645,N_8681);
nand U9388 (N_9388,N_8779,N_8661);
and U9389 (N_9389,N_8627,N_8503);
and U9390 (N_9390,N_8544,N_8509);
nor U9391 (N_9391,N_8638,N_8552);
nor U9392 (N_9392,N_8530,N_8815);
nand U9393 (N_9393,N_8678,N_8506);
or U9394 (N_9394,N_8747,N_8799);
nor U9395 (N_9395,N_8642,N_8726);
or U9396 (N_9396,N_8955,N_8696);
and U9397 (N_9397,N_8972,N_8728);
nor U9398 (N_9398,N_8712,N_8878);
or U9399 (N_9399,N_8771,N_8663);
nand U9400 (N_9400,N_8505,N_8638);
nand U9401 (N_9401,N_8537,N_8743);
nand U9402 (N_9402,N_8701,N_8628);
and U9403 (N_9403,N_8798,N_8529);
nand U9404 (N_9404,N_8767,N_8630);
and U9405 (N_9405,N_8824,N_8790);
and U9406 (N_9406,N_8516,N_8966);
and U9407 (N_9407,N_8527,N_8522);
xnor U9408 (N_9408,N_8777,N_8988);
nand U9409 (N_9409,N_8998,N_8801);
nand U9410 (N_9410,N_8500,N_8604);
or U9411 (N_9411,N_8825,N_8569);
and U9412 (N_9412,N_8620,N_8735);
and U9413 (N_9413,N_8526,N_8728);
nand U9414 (N_9414,N_8511,N_8626);
and U9415 (N_9415,N_8658,N_8747);
or U9416 (N_9416,N_8903,N_8836);
xor U9417 (N_9417,N_8751,N_8867);
xnor U9418 (N_9418,N_8712,N_8524);
and U9419 (N_9419,N_8925,N_8792);
nand U9420 (N_9420,N_8848,N_8680);
or U9421 (N_9421,N_8570,N_8929);
xnor U9422 (N_9422,N_8936,N_8984);
or U9423 (N_9423,N_8651,N_8654);
nor U9424 (N_9424,N_8848,N_8810);
and U9425 (N_9425,N_8552,N_8728);
xnor U9426 (N_9426,N_8994,N_8646);
and U9427 (N_9427,N_8722,N_8655);
nor U9428 (N_9428,N_8549,N_8799);
and U9429 (N_9429,N_8986,N_8984);
nand U9430 (N_9430,N_8883,N_8628);
and U9431 (N_9431,N_8633,N_8723);
nor U9432 (N_9432,N_8611,N_8727);
xnor U9433 (N_9433,N_8942,N_8914);
or U9434 (N_9434,N_8732,N_8897);
xor U9435 (N_9435,N_8957,N_8936);
and U9436 (N_9436,N_8815,N_8744);
and U9437 (N_9437,N_8796,N_8840);
and U9438 (N_9438,N_8892,N_8715);
nor U9439 (N_9439,N_8879,N_8882);
nor U9440 (N_9440,N_8637,N_8641);
and U9441 (N_9441,N_8585,N_8895);
and U9442 (N_9442,N_8733,N_8644);
nand U9443 (N_9443,N_8776,N_8563);
xnor U9444 (N_9444,N_8634,N_8635);
xnor U9445 (N_9445,N_8866,N_8882);
and U9446 (N_9446,N_8526,N_8817);
xor U9447 (N_9447,N_8755,N_8567);
nand U9448 (N_9448,N_8571,N_8532);
xor U9449 (N_9449,N_8573,N_8931);
and U9450 (N_9450,N_8601,N_8925);
nand U9451 (N_9451,N_8893,N_8628);
or U9452 (N_9452,N_8918,N_8743);
nor U9453 (N_9453,N_8778,N_8523);
nor U9454 (N_9454,N_8511,N_8561);
or U9455 (N_9455,N_8940,N_8715);
xor U9456 (N_9456,N_8772,N_8779);
or U9457 (N_9457,N_8920,N_8991);
and U9458 (N_9458,N_8812,N_8639);
nor U9459 (N_9459,N_8853,N_8752);
or U9460 (N_9460,N_8591,N_8723);
and U9461 (N_9461,N_8793,N_8764);
xnor U9462 (N_9462,N_8895,N_8565);
xor U9463 (N_9463,N_8712,N_8582);
nor U9464 (N_9464,N_8774,N_8676);
xor U9465 (N_9465,N_8996,N_8951);
and U9466 (N_9466,N_8586,N_8639);
and U9467 (N_9467,N_8960,N_8952);
nand U9468 (N_9468,N_8811,N_8523);
xnor U9469 (N_9469,N_8820,N_8622);
nand U9470 (N_9470,N_8992,N_8856);
nand U9471 (N_9471,N_8729,N_8589);
nand U9472 (N_9472,N_8946,N_8919);
and U9473 (N_9473,N_8505,N_8827);
or U9474 (N_9474,N_8726,N_8543);
nor U9475 (N_9475,N_8646,N_8526);
xnor U9476 (N_9476,N_8787,N_8820);
and U9477 (N_9477,N_8780,N_8762);
and U9478 (N_9478,N_8700,N_8835);
xnor U9479 (N_9479,N_8513,N_8837);
or U9480 (N_9480,N_8607,N_8908);
nor U9481 (N_9481,N_8893,N_8522);
nand U9482 (N_9482,N_8921,N_8803);
nand U9483 (N_9483,N_8881,N_8896);
xnor U9484 (N_9484,N_8608,N_8701);
nor U9485 (N_9485,N_8997,N_8762);
and U9486 (N_9486,N_8612,N_8616);
and U9487 (N_9487,N_8642,N_8500);
xnor U9488 (N_9488,N_8607,N_8739);
nand U9489 (N_9489,N_8796,N_8771);
and U9490 (N_9490,N_8638,N_8985);
and U9491 (N_9491,N_8638,N_8870);
nor U9492 (N_9492,N_8672,N_8656);
nor U9493 (N_9493,N_8639,N_8834);
xor U9494 (N_9494,N_8589,N_8646);
and U9495 (N_9495,N_8770,N_8854);
and U9496 (N_9496,N_8543,N_8920);
or U9497 (N_9497,N_8684,N_8869);
or U9498 (N_9498,N_8605,N_8576);
nand U9499 (N_9499,N_8986,N_8752);
xnor U9500 (N_9500,N_9048,N_9338);
nor U9501 (N_9501,N_9109,N_9020);
nand U9502 (N_9502,N_9251,N_9231);
or U9503 (N_9503,N_9267,N_9101);
and U9504 (N_9504,N_9221,N_9033);
or U9505 (N_9505,N_9166,N_9117);
xor U9506 (N_9506,N_9055,N_9031);
or U9507 (N_9507,N_9167,N_9461);
or U9508 (N_9508,N_9256,N_9200);
and U9509 (N_9509,N_9034,N_9174);
and U9510 (N_9510,N_9410,N_9337);
nand U9511 (N_9511,N_9148,N_9437);
and U9512 (N_9512,N_9196,N_9252);
nand U9513 (N_9513,N_9136,N_9211);
nor U9514 (N_9514,N_9001,N_9038);
xor U9515 (N_9515,N_9406,N_9115);
nand U9516 (N_9516,N_9016,N_9495);
or U9517 (N_9517,N_9325,N_9287);
nand U9518 (N_9518,N_9216,N_9318);
nor U9519 (N_9519,N_9379,N_9364);
xor U9520 (N_9520,N_9181,N_9201);
nor U9521 (N_9521,N_9343,N_9341);
nand U9522 (N_9522,N_9208,N_9183);
or U9523 (N_9523,N_9250,N_9476);
nand U9524 (N_9524,N_9039,N_9254);
or U9525 (N_9525,N_9123,N_9004);
nor U9526 (N_9526,N_9145,N_9046);
and U9527 (N_9527,N_9085,N_9035);
or U9528 (N_9528,N_9297,N_9207);
nand U9529 (N_9529,N_9296,N_9422);
or U9530 (N_9530,N_9356,N_9053);
nand U9531 (N_9531,N_9172,N_9150);
nor U9532 (N_9532,N_9059,N_9402);
or U9533 (N_9533,N_9158,N_9224);
or U9534 (N_9534,N_9336,N_9306);
nor U9535 (N_9535,N_9449,N_9490);
nor U9536 (N_9536,N_9178,N_9245);
xnor U9537 (N_9537,N_9486,N_9271);
xor U9538 (N_9538,N_9481,N_9458);
or U9539 (N_9539,N_9403,N_9023);
nand U9540 (N_9540,N_9442,N_9353);
nand U9541 (N_9541,N_9180,N_9433);
nand U9542 (N_9542,N_9303,N_9078);
nand U9543 (N_9543,N_9460,N_9041);
nor U9544 (N_9544,N_9420,N_9463);
or U9545 (N_9545,N_9195,N_9096);
or U9546 (N_9546,N_9143,N_9161);
xor U9547 (N_9547,N_9242,N_9398);
nand U9548 (N_9548,N_9329,N_9083);
xnor U9549 (N_9549,N_9198,N_9236);
nand U9550 (N_9550,N_9484,N_9488);
or U9551 (N_9551,N_9399,N_9134);
and U9552 (N_9552,N_9247,N_9194);
xor U9553 (N_9553,N_9400,N_9452);
nor U9554 (N_9554,N_9068,N_9259);
xor U9555 (N_9555,N_9446,N_9372);
or U9556 (N_9556,N_9319,N_9385);
or U9557 (N_9557,N_9210,N_9137);
or U9558 (N_9558,N_9025,N_9071);
and U9559 (N_9559,N_9238,N_9474);
nand U9560 (N_9560,N_9139,N_9080);
and U9561 (N_9561,N_9088,N_9368);
and U9562 (N_9562,N_9072,N_9431);
nand U9563 (N_9563,N_9010,N_9413);
and U9564 (N_9564,N_9185,N_9387);
and U9565 (N_9565,N_9301,N_9441);
or U9566 (N_9566,N_9465,N_9171);
nor U9567 (N_9567,N_9454,N_9040);
and U9568 (N_9568,N_9013,N_9322);
or U9569 (N_9569,N_9065,N_9307);
or U9570 (N_9570,N_9005,N_9237);
nand U9571 (N_9571,N_9036,N_9469);
nand U9572 (N_9572,N_9478,N_9348);
nand U9573 (N_9573,N_9386,N_9113);
nand U9574 (N_9574,N_9027,N_9396);
nor U9575 (N_9575,N_9324,N_9104);
nand U9576 (N_9576,N_9135,N_9186);
or U9577 (N_9577,N_9054,N_9388);
and U9578 (N_9578,N_9008,N_9483);
and U9579 (N_9579,N_9350,N_9017);
nor U9580 (N_9580,N_9073,N_9373);
nor U9581 (N_9581,N_9280,N_9149);
and U9582 (N_9582,N_9007,N_9082);
or U9583 (N_9583,N_9173,N_9432);
nand U9584 (N_9584,N_9276,N_9089);
nor U9585 (N_9585,N_9380,N_9006);
nand U9586 (N_9586,N_9225,N_9220);
nand U9587 (N_9587,N_9191,N_9384);
or U9588 (N_9588,N_9187,N_9009);
xnor U9589 (N_9589,N_9428,N_9057);
or U9590 (N_9590,N_9435,N_9327);
nand U9591 (N_9591,N_9351,N_9299);
xnor U9592 (N_9592,N_9045,N_9049);
or U9593 (N_9593,N_9443,N_9480);
and U9594 (N_9594,N_9206,N_9241);
xnor U9595 (N_9595,N_9367,N_9393);
and U9596 (N_9596,N_9290,N_9357);
or U9597 (N_9597,N_9391,N_9074);
xnor U9598 (N_9598,N_9118,N_9315);
xor U9599 (N_9599,N_9000,N_9121);
and U9600 (N_9600,N_9248,N_9347);
xor U9601 (N_9601,N_9122,N_9240);
nor U9602 (N_9602,N_9365,N_9294);
or U9603 (N_9603,N_9244,N_9044);
nand U9604 (N_9604,N_9266,N_9439);
nand U9605 (N_9605,N_9392,N_9147);
and U9606 (N_9606,N_9098,N_9093);
and U9607 (N_9607,N_9494,N_9272);
xnor U9608 (N_9608,N_9157,N_9485);
or U9609 (N_9609,N_9355,N_9103);
or U9610 (N_9610,N_9475,N_9190);
xor U9611 (N_9611,N_9014,N_9361);
and U9612 (N_9612,N_9119,N_9345);
nand U9613 (N_9613,N_9346,N_9226);
or U9614 (N_9614,N_9340,N_9164);
nor U9615 (N_9615,N_9366,N_9026);
nand U9616 (N_9616,N_9107,N_9378);
xor U9617 (N_9617,N_9138,N_9492);
xor U9618 (N_9618,N_9470,N_9414);
or U9619 (N_9619,N_9199,N_9275);
xor U9620 (N_9620,N_9155,N_9423);
or U9621 (N_9621,N_9270,N_9067);
xnor U9622 (N_9622,N_9412,N_9144);
nand U9623 (N_9623,N_9335,N_9124);
or U9624 (N_9624,N_9202,N_9168);
nand U9625 (N_9625,N_9419,N_9305);
xor U9626 (N_9626,N_9300,N_9451);
or U9627 (N_9627,N_9030,N_9298);
nand U9628 (N_9628,N_9142,N_9462);
xnor U9629 (N_9629,N_9170,N_9427);
or U9630 (N_9630,N_9448,N_9456);
or U9631 (N_9631,N_9283,N_9421);
xnor U9632 (N_9632,N_9383,N_9028);
or U9633 (N_9633,N_9112,N_9471);
or U9634 (N_9634,N_9349,N_9232);
nor U9635 (N_9635,N_9024,N_9105);
or U9636 (N_9636,N_9404,N_9152);
and U9637 (N_9637,N_9424,N_9243);
and U9638 (N_9638,N_9309,N_9050);
nand U9639 (N_9639,N_9311,N_9192);
xor U9640 (N_9640,N_9417,N_9457);
xnor U9641 (N_9641,N_9116,N_9175);
and U9642 (N_9642,N_9111,N_9496);
or U9643 (N_9643,N_9019,N_9091);
xnor U9644 (N_9644,N_9429,N_9012);
nand U9645 (N_9645,N_9255,N_9092);
xnor U9646 (N_9646,N_9162,N_9097);
or U9647 (N_9647,N_9289,N_9288);
xor U9648 (N_9648,N_9022,N_9015);
or U9649 (N_9649,N_9189,N_9331);
nand U9650 (N_9650,N_9131,N_9263);
xor U9651 (N_9651,N_9360,N_9376);
nor U9652 (N_9652,N_9405,N_9308);
nor U9653 (N_9653,N_9156,N_9169);
or U9654 (N_9654,N_9265,N_9100);
and U9655 (N_9655,N_9440,N_9472);
nand U9656 (N_9656,N_9227,N_9438);
or U9657 (N_9657,N_9094,N_9077);
and U9658 (N_9658,N_9102,N_9295);
xor U9659 (N_9659,N_9377,N_9127);
and U9660 (N_9660,N_9051,N_9323);
and U9661 (N_9661,N_9214,N_9179);
nor U9662 (N_9662,N_9467,N_9262);
nor U9663 (N_9663,N_9268,N_9445);
and U9664 (N_9664,N_9160,N_9370);
nor U9665 (N_9665,N_9277,N_9018);
nand U9666 (N_9666,N_9302,N_9493);
and U9667 (N_9667,N_9430,N_9163);
nor U9668 (N_9668,N_9217,N_9132);
or U9669 (N_9669,N_9062,N_9293);
and U9670 (N_9670,N_9408,N_9409);
nand U9671 (N_9671,N_9076,N_9159);
and U9672 (N_9672,N_9459,N_9052);
nand U9673 (N_9673,N_9099,N_9213);
nor U9674 (N_9674,N_9333,N_9334);
or U9675 (N_9675,N_9029,N_9032);
xor U9676 (N_9676,N_9130,N_9269);
xnor U9677 (N_9677,N_9182,N_9284);
nand U9678 (N_9678,N_9063,N_9090);
or U9679 (N_9679,N_9278,N_9426);
nand U9680 (N_9680,N_9497,N_9416);
or U9681 (N_9681,N_9235,N_9193);
nand U9682 (N_9682,N_9390,N_9291);
xnor U9683 (N_9683,N_9253,N_9258);
or U9684 (N_9684,N_9316,N_9285);
and U9685 (N_9685,N_9095,N_9418);
nor U9686 (N_9686,N_9060,N_9079);
or U9687 (N_9687,N_9128,N_9371);
and U9688 (N_9688,N_9129,N_9395);
xnor U9689 (N_9689,N_9218,N_9184);
nand U9690 (N_9690,N_9140,N_9491);
xor U9691 (N_9691,N_9363,N_9215);
nor U9692 (N_9692,N_9344,N_9205);
xnor U9693 (N_9693,N_9197,N_9279);
nor U9694 (N_9694,N_9106,N_9487);
or U9695 (N_9695,N_9042,N_9229);
nand U9696 (N_9696,N_9146,N_9075);
nand U9697 (N_9697,N_9069,N_9056);
nor U9698 (N_9698,N_9282,N_9321);
or U9699 (N_9699,N_9153,N_9081);
nor U9700 (N_9700,N_9257,N_9249);
and U9701 (N_9701,N_9310,N_9087);
xnor U9702 (N_9702,N_9133,N_9264);
and U9703 (N_9703,N_9394,N_9228);
or U9704 (N_9704,N_9342,N_9482);
nor U9705 (N_9705,N_9219,N_9209);
nor U9706 (N_9706,N_9313,N_9468);
nor U9707 (N_9707,N_9234,N_9314);
xnor U9708 (N_9708,N_9369,N_9382);
nand U9709 (N_9709,N_9108,N_9401);
nand U9710 (N_9710,N_9233,N_9498);
nor U9711 (N_9711,N_9320,N_9479);
xor U9712 (N_9712,N_9260,N_9415);
xor U9713 (N_9713,N_9434,N_9274);
nor U9714 (N_9714,N_9188,N_9436);
nand U9715 (N_9715,N_9246,N_9312);
or U9716 (N_9716,N_9058,N_9281);
nor U9717 (N_9717,N_9086,N_9477);
nand U9718 (N_9718,N_9002,N_9411);
or U9719 (N_9719,N_9154,N_9444);
and U9720 (N_9720,N_9466,N_9273);
xor U9721 (N_9721,N_9397,N_9359);
xnor U9722 (N_9722,N_9204,N_9230);
nand U9723 (N_9723,N_9381,N_9212);
or U9724 (N_9724,N_9021,N_9114);
xor U9725 (N_9725,N_9455,N_9354);
or U9726 (N_9726,N_9165,N_9177);
nand U9727 (N_9727,N_9499,N_9043);
and U9728 (N_9728,N_9326,N_9066);
xnor U9729 (N_9729,N_9037,N_9450);
nand U9730 (N_9730,N_9261,N_9239);
nand U9731 (N_9731,N_9352,N_9304);
and U9732 (N_9732,N_9203,N_9064);
or U9733 (N_9733,N_9011,N_9407);
and U9734 (N_9734,N_9317,N_9222);
or U9735 (N_9735,N_9425,N_9126);
nand U9736 (N_9736,N_9473,N_9489);
xnor U9737 (N_9737,N_9375,N_9223);
nand U9738 (N_9738,N_9120,N_9141);
nand U9739 (N_9739,N_9151,N_9125);
and U9740 (N_9740,N_9374,N_9362);
or U9741 (N_9741,N_9330,N_9464);
or U9742 (N_9742,N_9061,N_9176);
nand U9743 (N_9743,N_9070,N_9328);
and U9744 (N_9744,N_9332,N_9358);
xor U9745 (N_9745,N_9084,N_9389);
or U9746 (N_9746,N_9447,N_9286);
or U9747 (N_9747,N_9292,N_9110);
nor U9748 (N_9748,N_9047,N_9453);
xor U9749 (N_9749,N_9339,N_9003);
nor U9750 (N_9750,N_9031,N_9429);
xor U9751 (N_9751,N_9422,N_9130);
nor U9752 (N_9752,N_9494,N_9315);
nand U9753 (N_9753,N_9092,N_9334);
nor U9754 (N_9754,N_9416,N_9007);
and U9755 (N_9755,N_9022,N_9101);
xor U9756 (N_9756,N_9346,N_9338);
or U9757 (N_9757,N_9389,N_9253);
nor U9758 (N_9758,N_9028,N_9254);
and U9759 (N_9759,N_9442,N_9009);
and U9760 (N_9760,N_9320,N_9166);
nor U9761 (N_9761,N_9402,N_9363);
xnor U9762 (N_9762,N_9390,N_9190);
and U9763 (N_9763,N_9332,N_9388);
nand U9764 (N_9764,N_9377,N_9093);
and U9765 (N_9765,N_9067,N_9334);
or U9766 (N_9766,N_9135,N_9480);
nand U9767 (N_9767,N_9059,N_9123);
or U9768 (N_9768,N_9244,N_9163);
or U9769 (N_9769,N_9312,N_9089);
nand U9770 (N_9770,N_9296,N_9178);
and U9771 (N_9771,N_9195,N_9002);
nand U9772 (N_9772,N_9389,N_9434);
or U9773 (N_9773,N_9178,N_9342);
or U9774 (N_9774,N_9400,N_9053);
or U9775 (N_9775,N_9024,N_9449);
nor U9776 (N_9776,N_9210,N_9410);
xnor U9777 (N_9777,N_9164,N_9444);
xnor U9778 (N_9778,N_9022,N_9389);
xor U9779 (N_9779,N_9180,N_9131);
nand U9780 (N_9780,N_9197,N_9206);
nor U9781 (N_9781,N_9391,N_9428);
and U9782 (N_9782,N_9002,N_9404);
xnor U9783 (N_9783,N_9314,N_9324);
or U9784 (N_9784,N_9469,N_9280);
and U9785 (N_9785,N_9366,N_9133);
nand U9786 (N_9786,N_9380,N_9323);
nor U9787 (N_9787,N_9171,N_9036);
nand U9788 (N_9788,N_9051,N_9183);
nor U9789 (N_9789,N_9362,N_9418);
nand U9790 (N_9790,N_9282,N_9249);
nand U9791 (N_9791,N_9458,N_9207);
or U9792 (N_9792,N_9390,N_9146);
xor U9793 (N_9793,N_9187,N_9297);
xor U9794 (N_9794,N_9092,N_9451);
nand U9795 (N_9795,N_9344,N_9463);
xnor U9796 (N_9796,N_9414,N_9169);
xnor U9797 (N_9797,N_9408,N_9487);
and U9798 (N_9798,N_9025,N_9044);
or U9799 (N_9799,N_9333,N_9172);
nand U9800 (N_9800,N_9455,N_9293);
xor U9801 (N_9801,N_9180,N_9152);
nand U9802 (N_9802,N_9006,N_9376);
nor U9803 (N_9803,N_9000,N_9277);
or U9804 (N_9804,N_9275,N_9484);
nand U9805 (N_9805,N_9365,N_9114);
nand U9806 (N_9806,N_9443,N_9065);
xor U9807 (N_9807,N_9120,N_9098);
or U9808 (N_9808,N_9265,N_9173);
xnor U9809 (N_9809,N_9426,N_9020);
xor U9810 (N_9810,N_9084,N_9313);
nand U9811 (N_9811,N_9106,N_9451);
nand U9812 (N_9812,N_9323,N_9024);
and U9813 (N_9813,N_9390,N_9100);
and U9814 (N_9814,N_9355,N_9420);
xor U9815 (N_9815,N_9326,N_9259);
and U9816 (N_9816,N_9067,N_9407);
nand U9817 (N_9817,N_9224,N_9096);
or U9818 (N_9818,N_9062,N_9436);
or U9819 (N_9819,N_9498,N_9416);
xnor U9820 (N_9820,N_9455,N_9460);
nor U9821 (N_9821,N_9310,N_9291);
nand U9822 (N_9822,N_9217,N_9478);
xnor U9823 (N_9823,N_9451,N_9207);
and U9824 (N_9824,N_9109,N_9301);
nor U9825 (N_9825,N_9299,N_9175);
and U9826 (N_9826,N_9455,N_9320);
nor U9827 (N_9827,N_9371,N_9247);
nor U9828 (N_9828,N_9117,N_9126);
or U9829 (N_9829,N_9460,N_9493);
nor U9830 (N_9830,N_9333,N_9312);
nand U9831 (N_9831,N_9261,N_9348);
nand U9832 (N_9832,N_9152,N_9247);
xnor U9833 (N_9833,N_9007,N_9284);
nand U9834 (N_9834,N_9499,N_9109);
or U9835 (N_9835,N_9285,N_9287);
or U9836 (N_9836,N_9439,N_9275);
nor U9837 (N_9837,N_9015,N_9180);
or U9838 (N_9838,N_9366,N_9286);
xor U9839 (N_9839,N_9476,N_9275);
nor U9840 (N_9840,N_9131,N_9433);
nor U9841 (N_9841,N_9317,N_9225);
or U9842 (N_9842,N_9160,N_9123);
xor U9843 (N_9843,N_9373,N_9196);
nand U9844 (N_9844,N_9170,N_9333);
nand U9845 (N_9845,N_9024,N_9162);
or U9846 (N_9846,N_9478,N_9407);
nor U9847 (N_9847,N_9441,N_9197);
or U9848 (N_9848,N_9273,N_9004);
nand U9849 (N_9849,N_9455,N_9145);
and U9850 (N_9850,N_9111,N_9181);
nand U9851 (N_9851,N_9437,N_9035);
or U9852 (N_9852,N_9003,N_9196);
nor U9853 (N_9853,N_9177,N_9435);
nor U9854 (N_9854,N_9123,N_9212);
or U9855 (N_9855,N_9351,N_9287);
or U9856 (N_9856,N_9476,N_9194);
and U9857 (N_9857,N_9092,N_9407);
and U9858 (N_9858,N_9325,N_9477);
xor U9859 (N_9859,N_9047,N_9256);
xor U9860 (N_9860,N_9147,N_9362);
xnor U9861 (N_9861,N_9341,N_9161);
nand U9862 (N_9862,N_9425,N_9222);
nand U9863 (N_9863,N_9000,N_9225);
or U9864 (N_9864,N_9305,N_9295);
nand U9865 (N_9865,N_9132,N_9199);
or U9866 (N_9866,N_9110,N_9418);
nand U9867 (N_9867,N_9103,N_9061);
nand U9868 (N_9868,N_9282,N_9028);
nor U9869 (N_9869,N_9190,N_9300);
nor U9870 (N_9870,N_9340,N_9035);
nand U9871 (N_9871,N_9242,N_9323);
or U9872 (N_9872,N_9403,N_9281);
xor U9873 (N_9873,N_9262,N_9013);
nand U9874 (N_9874,N_9068,N_9112);
nor U9875 (N_9875,N_9313,N_9018);
or U9876 (N_9876,N_9336,N_9466);
or U9877 (N_9877,N_9403,N_9385);
xnor U9878 (N_9878,N_9160,N_9254);
nand U9879 (N_9879,N_9233,N_9384);
or U9880 (N_9880,N_9380,N_9385);
and U9881 (N_9881,N_9455,N_9205);
and U9882 (N_9882,N_9416,N_9453);
nor U9883 (N_9883,N_9107,N_9395);
or U9884 (N_9884,N_9329,N_9027);
and U9885 (N_9885,N_9322,N_9038);
and U9886 (N_9886,N_9302,N_9452);
xor U9887 (N_9887,N_9373,N_9379);
or U9888 (N_9888,N_9467,N_9310);
xnor U9889 (N_9889,N_9025,N_9407);
or U9890 (N_9890,N_9411,N_9359);
xnor U9891 (N_9891,N_9486,N_9176);
xor U9892 (N_9892,N_9372,N_9214);
nor U9893 (N_9893,N_9285,N_9175);
nand U9894 (N_9894,N_9276,N_9039);
nor U9895 (N_9895,N_9492,N_9185);
xor U9896 (N_9896,N_9476,N_9146);
or U9897 (N_9897,N_9358,N_9015);
nor U9898 (N_9898,N_9081,N_9326);
and U9899 (N_9899,N_9012,N_9017);
and U9900 (N_9900,N_9247,N_9478);
nand U9901 (N_9901,N_9030,N_9436);
and U9902 (N_9902,N_9271,N_9254);
nor U9903 (N_9903,N_9180,N_9200);
xnor U9904 (N_9904,N_9205,N_9479);
nand U9905 (N_9905,N_9119,N_9164);
or U9906 (N_9906,N_9328,N_9238);
or U9907 (N_9907,N_9082,N_9300);
and U9908 (N_9908,N_9054,N_9008);
xnor U9909 (N_9909,N_9209,N_9333);
nor U9910 (N_9910,N_9241,N_9378);
nor U9911 (N_9911,N_9408,N_9363);
nor U9912 (N_9912,N_9122,N_9297);
nor U9913 (N_9913,N_9135,N_9091);
nor U9914 (N_9914,N_9122,N_9039);
nand U9915 (N_9915,N_9291,N_9003);
and U9916 (N_9916,N_9425,N_9427);
nor U9917 (N_9917,N_9404,N_9274);
nor U9918 (N_9918,N_9333,N_9108);
and U9919 (N_9919,N_9156,N_9202);
nor U9920 (N_9920,N_9107,N_9418);
or U9921 (N_9921,N_9399,N_9224);
and U9922 (N_9922,N_9115,N_9496);
nor U9923 (N_9923,N_9351,N_9424);
nand U9924 (N_9924,N_9117,N_9194);
xnor U9925 (N_9925,N_9253,N_9478);
nor U9926 (N_9926,N_9014,N_9264);
and U9927 (N_9927,N_9344,N_9206);
and U9928 (N_9928,N_9334,N_9036);
or U9929 (N_9929,N_9055,N_9157);
and U9930 (N_9930,N_9210,N_9318);
and U9931 (N_9931,N_9384,N_9310);
nand U9932 (N_9932,N_9145,N_9123);
and U9933 (N_9933,N_9198,N_9424);
nor U9934 (N_9934,N_9119,N_9343);
or U9935 (N_9935,N_9002,N_9095);
and U9936 (N_9936,N_9377,N_9231);
or U9937 (N_9937,N_9070,N_9233);
nor U9938 (N_9938,N_9416,N_9200);
or U9939 (N_9939,N_9440,N_9297);
and U9940 (N_9940,N_9332,N_9404);
xor U9941 (N_9941,N_9488,N_9048);
xnor U9942 (N_9942,N_9092,N_9382);
xnor U9943 (N_9943,N_9094,N_9153);
and U9944 (N_9944,N_9271,N_9068);
nor U9945 (N_9945,N_9216,N_9310);
and U9946 (N_9946,N_9421,N_9474);
or U9947 (N_9947,N_9324,N_9041);
xnor U9948 (N_9948,N_9021,N_9136);
or U9949 (N_9949,N_9256,N_9316);
xnor U9950 (N_9950,N_9424,N_9241);
nand U9951 (N_9951,N_9150,N_9108);
xnor U9952 (N_9952,N_9085,N_9204);
and U9953 (N_9953,N_9462,N_9293);
xnor U9954 (N_9954,N_9148,N_9083);
nor U9955 (N_9955,N_9279,N_9122);
and U9956 (N_9956,N_9459,N_9154);
nand U9957 (N_9957,N_9324,N_9031);
xnor U9958 (N_9958,N_9260,N_9448);
and U9959 (N_9959,N_9217,N_9379);
xor U9960 (N_9960,N_9486,N_9170);
xnor U9961 (N_9961,N_9458,N_9146);
or U9962 (N_9962,N_9456,N_9413);
or U9963 (N_9963,N_9415,N_9417);
nand U9964 (N_9964,N_9367,N_9429);
nor U9965 (N_9965,N_9051,N_9037);
nor U9966 (N_9966,N_9203,N_9146);
nand U9967 (N_9967,N_9175,N_9226);
xor U9968 (N_9968,N_9175,N_9247);
xnor U9969 (N_9969,N_9389,N_9258);
nor U9970 (N_9970,N_9321,N_9266);
or U9971 (N_9971,N_9272,N_9368);
and U9972 (N_9972,N_9425,N_9224);
or U9973 (N_9973,N_9477,N_9359);
nor U9974 (N_9974,N_9319,N_9413);
or U9975 (N_9975,N_9180,N_9379);
nand U9976 (N_9976,N_9348,N_9184);
and U9977 (N_9977,N_9199,N_9305);
nand U9978 (N_9978,N_9495,N_9419);
and U9979 (N_9979,N_9368,N_9085);
nor U9980 (N_9980,N_9108,N_9138);
or U9981 (N_9981,N_9473,N_9010);
nor U9982 (N_9982,N_9362,N_9177);
or U9983 (N_9983,N_9135,N_9120);
nand U9984 (N_9984,N_9387,N_9315);
nand U9985 (N_9985,N_9466,N_9186);
and U9986 (N_9986,N_9234,N_9167);
or U9987 (N_9987,N_9425,N_9432);
xnor U9988 (N_9988,N_9398,N_9454);
nand U9989 (N_9989,N_9054,N_9057);
or U9990 (N_9990,N_9188,N_9326);
nor U9991 (N_9991,N_9369,N_9177);
or U9992 (N_9992,N_9029,N_9277);
nand U9993 (N_9993,N_9378,N_9089);
nor U9994 (N_9994,N_9329,N_9141);
nand U9995 (N_9995,N_9010,N_9083);
nand U9996 (N_9996,N_9145,N_9131);
and U9997 (N_9997,N_9069,N_9150);
xor U9998 (N_9998,N_9178,N_9120);
or U9999 (N_9999,N_9245,N_9081);
nor UO_0 (O_0,N_9925,N_9766);
xor UO_1 (O_1,N_9971,N_9592);
nor UO_2 (O_2,N_9929,N_9693);
nand UO_3 (O_3,N_9579,N_9876);
and UO_4 (O_4,N_9632,N_9783);
nand UO_5 (O_5,N_9906,N_9989);
xor UO_6 (O_6,N_9904,N_9558);
or UO_7 (O_7,N_9886,N_9712);
nand UO_8 (O_8,N_9577,N_9718);
nor UO_9 (O_9,N_9782,N_9556);
nand UO_10 (O_10,N_9798,N_9963);
or UO_11 (O_11,N_9566,N_9986);
or UO_12 (O_12,N_9542,N_9832);
xor UO_13 (O_13,N_9786,N_9868);
xnor UO_14 (O_14,N_9842,N_9979);
nor UO_15 (O_15,N_9760,N_9841);
and UO_16 (O_16,N_9994,N_9801);
xnor UO_17 (O_17,N_9500,N_9649);
or UO_18 (O_18,N_9888,N_9526);
and UO_19 (O_19,N_9624,N_9763);
and UO_20 (O_20,N_9557,N_9825);
nor UO_21 (O_21,N_9992,N_9941);
nand UO_22 (O_22,N_9799,N_9748);
nand UO_23 (O_23,N_9590,N_9501);
xor UO_24 (O_24,N_9513,N_9749);
and UO_25 (O_25,N_9974,N_9978);
and UO_26 (O_26,N_9584,N_9713);
nor UO_27 (O_27,N_9741,N_9933);
nor UO_28 (O_28,N_9787,N_9525);
and UO_29 (O_29,N_9602,N_9678);
nand UO_30 (O_30,N_9761,N_9729);
xnor UO_31 (O_31,N_9769,N_9725);
nor UO_32 (O_32,N_9637,N_9685);
nor UO_33 (O_33,N_9747,N_9613);
nand UO_34 (O_34,N_9908,N_9936);
or UO_35 (O_35,N_9569,N_9515);
and UO_36 (O_36,N_9957,N_9744);
or UO_37 (O_37,N_9879,N_9669);
or UO_38 (O_38,N_9504,N_9607);
xnor UO_39 (O_39,N_9830,N_9991);
xnor UO_40 (O_40,N_9634,N_9924);
and UO_41 (O_41,N_9671,N_9968);
nand UO_42 (O_42,N_9919,N_9719);
and UO_43 (O_43,N_9511,N_9596);
xnor UO_44 (O_44,N_9785,N_9739);
or UO_45 (O_45,N_9883,N_9606);
nor UO_46 (O_46,N_9840,N_9716);
or UO_47 (O_47,N_9539,N_9853);
nand UO_48 (O_48,N_9625,N_9582);
and UO_49 (O_49,N_9930,N_9772);
and UO_50 (O_50,N_9647,N_9848);
nor UO_51 (O_51,N_9820,N_9838);
and UO_52 (O_52,N_9640,N_9949);
or UO_53 (O_53,N_9554,N_9823);
nor UO_54 (O_54,N_9854,N_9656);
nand UO_55 (O_55,N_9921,N_9628);
xor UO_56 (O_56,N_9984,N_9960);
or UO_57 (O_57,N_9997,N_9752);
nor UO_58 (O_58,N_9561,N_9808);
xnor UO_59 (O_59,N_9896,N_9604);
and UO_60 (O_60,N_9911,N_9845);
and UO_61 (O_61,N_9977,N_9810);
and UO_62 (O_62,N_9870,N_9524);
nand UO_63 (O_63,N_9814,N_9586);
nor UO_64 (O_64,N_9740,N_9675);
and UO_65 (O_65,N_9812,N_9616);
xor UO_66 (O_66,N_9573,N_9605);
and UO_67 (O_67,N_9756,N_9527);
or UO_68 (O_68,N_9519,N_9973);
xnor UO_69 (O_69,N_9630,N_9891);
or UO_70 (O_70,N_9563,N_9934);
nand UO_71 (O_71,N_9548,N_9790);
and UO_72 (O_72,N_9967,N_9806);
and UO_73 (O_73,N_9884,N_9950);
xor UO_74 (O_74,N_9633,N_9535);
or UO_75 (O_75,N_9560,N_9784);
xor UO_76 (O_76,N_9843,N_9619);
xnor UO_77 (O_77,N_9754,N_9775);
or UO_78 (O_78,N_9518,N_9594);
or UO_79 (O_79,N_9551,N_9947);
and UO_80 (O_80,N_9597,N_9581);
nor UO_81 (O_81,N_9550,N_9796);
xnor UO_82 (O_82,N_9909,N_9878);
xnor UO_83 (O_83,N_9762,N_9797);
xor UO_84 (O_84,N_9861,N_9564);
nor UO_85 (O_85,N_9965,N_9610);
nor UO_86 (O_86,N_9738,N_9734);
xnor UO_87 (O_87,N_9807,N_9774);
nor UO_88 (O_88,N_9863,N_9612);
nand UO_89 (O_89,N_9534,N_9860);
and UO_90 (O_90,N_9530,N_9636);
nor UO_91 (O_91,N_9804,N_9826);
and UO_92 (O_92,N_9710,N_9966);
xor UO_93 (O_93,N_9684,N_9846);
nor UO_94 (O_94,N_9847,N_9707);
nor UO_95 (O_95,N_9767,N_9578);
xnor UO_96 (O_96,N_9601,N_9758);
and UO_97 (O_97,N_9850,N_9621);
and UO_98 (O_98,N_9920,N_9750);
or UO_99 (O_99,N_9720,N_9828);
nor UO_100 (O_100,N_9559,N_9692);
or UO_101 (O_101,N_9708,N_9727);
xor UO_102 (O_102,N_9755,N_9664);
nand UO_103 (O_103,N_9673,N_9733);
nand UO_104 (O_104,N_9654,N_9976);
and UO_105 (O_105,N_9536,N_9617);
xor UO_106 (O_106,N_9588,N_9682);
nand UO_107 (O_107,N_9877,N_9901);
and UO_108 (O_108,N_9817,N_9824);
or UO_109 (O_109,N_9611,N_9507);
nor UO_110 (O_110,N_9653,N_9737);
xnor UO_111 (O_111,N_9913,N_9887);
or UO_112 (O_112,N_9657,N_9988);
xor UO_113 (O_113,N_9764,N_9618);
nand UO_114 (O_114,N_9598,N_9779);
or UO_115 (O_115,N_9773,N_9655);
or UO_116 (O_116,N_9969,N_9918);
xor UO_117 (O_117,N_9662,N_9958);
xnor UO_118 (O_118,N_9732,N_9943);
nor UO_119 (O_119,N_9627,N_9572);
xor UO_120 (O_120,N_9852,N_9609);
nor UO_121 (O_121,N_9857,N_9659);
or UO_122 (O_122,N_9660,N_9996);
and UO_123 (O_123,N_9895,N_9593);
and UO_124 (O_124,N_9856,N_9952);
or UO_125 (O_125,N_9910,N_9809);
xnor UO_126 (O_126,N_9698,N_9690);
and UO_127 (O_127,N_9699,N_9874);
and UO_128 (O_128,N_9702,N_9757);
nor UO_129 (O_129,N_9506,N_9704);
or UO_130 (O_130,N_9873,N_9917);
nand UO_131 (O_131,N_9570,N_9851);
nor UO_132 (O_132,N_9509,N_9905);
nand UO_133 (O_133,N_9945,N_9665);
and UO_134 (O_134,N_9962,N_9736);
nor UO_135 (O_135,N_9975,N_9717);
or UO_136 (O_136,N_9781,N_9789);
nand UO_137 (O_137,N_9803,N_9948);
or UO_138 (O_138,N_9663,N_9765);
or UO_139 (O_139,N_9651,N_9946);
and UO_140 (O_140,N_9916,N_9776);
nor UO_141 (O_141,N_9589,N_9932);
nand UO_142 (O_142,N_9714,N_9990);
or UO_143 (O_143,N_9768,N_9700);
nor UO_144 (O_144,N_9638,N_9697);
nand UO_145 (O_145,N_9677,N_9922);
nand UO_146 (O_146,N_9872,N_9742);
and UO_147 (O_147,N_9686,N_9746);
nor UO_148 (O_148,N_9529,N_9818);
nand UO_149 (O_149,N_9722,N_9844);
nand UO_150 (O_150,N_9939,N_9726);
nand UO_151 (O_151,N_9753,N_9687);
xnor UO_152 (O_152,N_9964,N_9993);
and UO_153 (O_153,N_9658,N_9800);
nor UO_154 (O_154,N_9689,N_9795);
nor UO_155 (O_155,N_9585,N_9829);
xnor UO_156 (O_156,N_9580,N_9695);
or UO_157 (O_157,N_9696,N_9982);
nand UO_158 (O_158,N_9902,N_9538);
nand UO_159 (O_159,N_9938,N_9721);
nand UO_160 (O_160,N_9959,N_9892);
and UO_161 (O_161,N_9547,N_9953);
nor UO_162 (O_162,N_9517,N_9723);
nor UO_163 (O_163,N_9885,N_9981);
xnor UO_164 (O_164,N_9935,N_9701);
nor UO_165 (O_165,N_9599,N_9780);
or UO_166 (O_166,N_9552,N_9859);
and UO_167 (O_167,N_9571,N_9691);
or UO_168 (O_168,N_9839,N_9822);
nand UO_169 (O_169,N_9703,N_9562);
nand UO_170 (O_170,N_9837,N_9866);
nand UO_171 (O_171,N_9543,N_9635);
and UO_172 (O_172,N_9648,N_9546);
nand UO_173 (O_173,N_9999,N_9813);
xnor UO_174 (O_174,N_9899,N_9890);
xor UO_175 (O_175,N_9942,N_9553);
nor UO_176 (O_176,N_9864,N_9680);
or UO_177 (O_177,N_9759,N_9591);
and UO_178 (O_178,N_9912,N_9502);
and UO_179 (O_179,N_9620,N_9623);
xnor UO_180 (O_180,N_9537,N_9565);
nor UO_181 (O_181,N_9792,N_9514);
and UO_182 (O_182,N_9642,N_9641);
or UO_183 (O_183,N_9724,N_9834);
xor UO_184 (O_184,N_9770,N_9907);
or UO_185 (O_185,N_9816,N_9927);
xor UO_186 (O_186,N_9652,N_9743);
or UO_187 (O_187,N_9614,N_9631);
or UO_188 (O_188,N_9626,N_9893);
xnor UO_189 (O_189,N_9674,N_9555);
or UO_190 (O_190,N_9954,N_9831);
xor UO_191 (O_191,N_9666,N_9728);
or UO_192 (O_192,N_9815,N_9849);
nor UO_193 (O_193,N_9972,N_9615);
nand UO_194 (O_194,N_9676,N_9833);
or UO_195 (O_195,N_9670,N_9882);
or UO_196 (O_196,N_9867,N_9510);
and UO_197 (O_197,N_9528,N_9875);
or UO_198 (O_198,N_9576,N_9894);
nand UO_199 (O_199,N_9928,N_9587);
and UO_200 (O_200,N_9520,N_9865);
nor UO_201 (O_201,N_9681,N_9532);
nor UO_202 (O_202,N_9523,N_9923);
xnor UO_203 (O_203,N_9937,N_9745);
xnor UO_204 (O_204,N_9567,N_9944);
nor UO_205 (O_205,N_9603,N_9650);
nand UO_206 (O_206,N_9987,N_9771);
nor UO_207 (O_207,N_9705,N_9512);
and UO_208 (O_208,N_9940,N_9955);
nand UO_209 (O_209,N_9531,N_9836);
nand UO_210 (O_210,N_9855,N_9583);
and UO_211 (O_211,N_9545,N_9898);
or UO_212 (O_212,N_9516,N_9629);
or UO_213 (O_213,N_9931,N_9998);
xor UO_214 (O_214,N_9679,N_9926);
and UO_215 (O_215,N_9788,N_9794);
and UO_216 (O_216,N_9683,N_9541);
nor UO_217 (O_217,N_9793,N_9903);
or UO_218 (O_218,N_9731,N_9672);
or UO_219 (O_219,N_9730,N_9951);
nor UO_220 (O_220,N_9821,N_9661);
and UO_221 (O_221,N_9915,N_9622);
or UO_222 (O_222,N_9715,N_9897);
nand UO_223 (O_223,N_9595,N_9871);
or UO_224 (O_224,N_9667,N_9711);
nand UO_225 (O_225,N_9533,N_9869);
nor UO_226 (O_226,N_9646,N_9503);
nor UO_227 (O_227,N_9961,N_9709);
and UO_228 (O_228,N_9880,N_9549);
or UO_229 (O_229,N_9778,N_9574);
nor UO_230 (O_230,N_9694,N_9568);
nand UO_231 (O_231,N_9575,N_9688);
nand UO_232 (O_232,N_9544,N_9835);
nand UO_233 (O_233,N_9881,N_9644);
and UO_234 (O_234,N_9858,N_9505);
xnor UO_235 (O_235,N_9827,N_9639);
nor UO_236 (O_236,N_9914,N_9956);
nand UO_237 (O_237,N_9805,N_9735);
nand UO_238 (O_238,N_9791,N_9777);
and UO_239 (O_239,N_9521,N_9522);
and UO_240 (O_240,N_9751,N_9706);
nor UO_241 (O_241,N_9508,N_9980);
and UO_242 (O_242,N_9608,N_9600);
nand UO_243 (O_243,N_9540,N_9889);
nand UO_244 (O_244,N_9811,N_9983);
and UO_245 (O_245,N_9819,N_9668);
and UO_246 (O_246,N_9862,N_9985);
nand UO_247 (O_247,N_9995,N_9900);
nor UO_248 (O_248,N_9643,N_9802);
or UO_249 (O_249,N_9645,N_9970);
nand UO_250 (O_250,N_9650,N_9633);
nor UO_251 (O_251,N_9829,N_9999);
nand UO_252 (O_252,N_9705,N_9969);
and UO_253 (O_253,N_9983,N_9886);
or UO_254 (O_254,N_9972,N_9631);
and UO_255 (O_255,N_9535,N_9597);
xor UO_256 (O_256,N_9821,N_9851);
xor UO_257 (O_257,N_9667,N_9863);
xnor UO_258 (O_258,N_9585,N_9763);
or UO_259 (O_259,N_9703,N_9578);
nand UO_260 (O_260,N_9846,N_9679);
nor UO_261 (O_261,N_9977,N_9647);
or UO_262 (O_262,N_9533,N_9837);
and UO_263 (O_263,N_9674,N_9857);
nand UO_264 (O_264,N_9870,N_9912);
xor UO_265 (O_265,N_9945,N_9921);
xor UO_266 (O_266,N_9947,N_9973);
xnor UO_267 (O_267,N_9757,N_9816);
xor UO_268 (O_268,N_9721,N_9692);
nand UO_269 (O_269,N_9696,N_9857);
nor UO_270 (O_270,N_9803,N_9583);
xor UO_271 (O_271,N_9701,N_9622);
xor UO_272 (O_272,N_9771,N_9719);
nand UO_273 (O_273,N_9965,N_9672);
or UO_274 (O_274,N_9548,N_9546);
nor UO_275 (O_275,N_9988,N_9729);
nor UO_276 (O_276,N_9974,N_9553);
nor UO_277 (O_277,N_9871,N_9813);
nor UO_278 (O_278,N_9797,N_9655);
xnor UO_279 (O_279,N_9845,N_9970);
and UO_280 (O_280,N_9726,N_9584);
and UO_281 (O_281,N_9922,N_9595);
nor UO_282 (O_282,N_9583,N_9973);
nor UO_283 (O_283,N_9539,N_9802);
and UO_284 (O_284,N_9924,N_9668);
nand UO_285 (O_285,N_9688,N_9803);
or UO_286 (O_286,N_9664,N_9732);
nor UO_287 (O_287,N_9758,N_9652);
xnor UO_288 (O_288,N_9634,N_9581);
and UO_289 (O_289,N_9842,N_9646);
nor UO_290 (O_290,N_9619,N_9639);
nand UO_291 (O_291,N_9846,N_9515);
xor UO_292 (O_292,N_9558,N_9567);
xor UO_293 (O_293,N_9558,N_9645);
xnor UO_294 (O_294,N_9546,N_9999);
or UO_295 (O_295,N_9541,N_9957);
xnor UO_296 (O_296,N_9969,N_9772);
nand UO_297 (O_297,N_9549,N_9672);
nor UO_298 (O_298,N_9644,N_9612);
nor UO_299 (O_299,N_9840,N_9927);
nand UO_300 (O_300,N_9559,N_9741);
and UO_301 (O_301,N_9710,N_9511);
and UO_302 (O_302,N_9750,N_9890);
nand UO_303 (O_303,N_9944,N_9885);
nand UO_304 (O_304,N_9814,N_9989);
xor UO_305 (O_305,N_9820,N_9742);
nor UO_306 (O_306,N_9692,N_9751);
or UO_307 (O_307,N_9828,N_9760);
nor UO_308 (O_308,N_9906,N_9733);
xnor UO_309 (O_309,N_9571,N_9849);
and UO_310 (O_310,N_9571,N_9778);
nand UO_311 (O_311,N_9906,N_9763);
nor UO_312 (O_312,N_9850,N_9506);
nor UO_313 (O_313,N_9656,N_9909);
or UO_314 (O_314,N_9709,N_9846);
and UO_315 (O_315,N_9895,N_9551);
and UO_316 (O_316,N_9977,N_9851);
nand UO_317 (O_317,N_9873,N_9688);
nor UO_318 (O_318,N_9764,N_9910);
or UO_319 (O_319,N_9866,N_9502);
nand UO_320 (O_320,N_9914,N_9737);
xnor UO_321 (O_321,N_9724,N_9785);
nand UO_322 (O_322,N_9650,N_9691);
or UO_323 (O_323,N_9538,N_9719);
nor UO_324 (O_324,N_9553,N_9656);
or UO_325 (O_325,N_9775,N_9860);
or UO_326 (O_326,N_9909,N_9581);
and UO_327 (O_327,N_9979,N_9540);
and UO_328 (O_328,N_9782,N_9578);
nand UO_329 (O_329,N_9795,N_9647);
nand UO_330 (O_330,N_9938,N_9580);
and UO_331 (O_331,N_9610,N_9995);
and UO_332 (O_332,N_9957,N_9930);
xnor UO_333 (O_333,N_9702,N_9706);
or UO_334 (O_334,N_9566,N_9596);
xnor UO_335 (O_335,N_9830,N_9864);
and UO_336 (O_336,N_9774,N_9536);
and UO_337 (O_337,N_9752,N_9871);
xor UO_338 (O_338,N_9735,N_9609);
xnor UO_339 (O_339,N_9904,N_9913);
or UO_340 (O_340,N_9979,N_9765);
or UO_341 (O_341,N_9688,N_9792);
nor UO_342 (O_342,N_9702,N_9715);
and UO_343 (O_343,N_9664,N_9610);
nor UO_344 (O_344,N_9583,N_9846);
nor UO_345 (O_345,N_9732,N_9637);
and UO_346 (O_346,N_9716,N_9645);
nor UO_347 (O_347,N_9549,N_9648);
and UO_348 (O_348,N_9750,N_9546);
xnor UO_349 (O_349,N_9831,N_9904);
or UO_350 (O_350,N_9824,N_9607);
xnor UO_351 (O_351,N_9861,N_9797);
nand UO_352 (O_352,N_9521,N_9642);
nor UO_353 (O_353,N_9580,N_9585);
or UO_354 (O_354,N_9770,N_9552);
or UO_355 (O_355,N_9621,N_9879);
and UO_356 (O_356,N_9937,N_9654);
xnor UO_357 (O_357,N_9538,N_9817);
and UO_358 (O_358,N_9676,N_9677);
nor UO_359 (O_359,N_9970,N_9836);
or UO_360 (O_360,N_9806,N_9525);
nor UO_361 (O_361,N_9690,N_9648);
and UO_362 (O_362,N_9960,N_9593);
xnor UO_363 (O_363,N_9885,N_9861);
xor UO_364 (O_364,N_9859,N_9936);
nor UO_365 (O_365,N_9994,N_9646);
nor UO_366 (O_366,N_9568,N_9758);
nor UO_367 (O_367,N_9891,N_9611);
nor UO_368 (O_368,N_9844,N_9731);
and UO_369 (O_369,N_9776,N_9561);
xnor UO_370 (O_370,N_9612,N_9999);
or UO_371 (O_371,N_9829,N_9825);
or UO_372 (O_372,N_9769,N_9858);
and UO_373 (O_373,N_9503,N_9713);
or UO_374 (O_374,N_9992,N_9743);
nor UO_375 (O_375,N_9608,N_9525);
nand UO_376 (O_376,N_9819,N_9584);
or UO_377 (O_377,N_9900,N_9788);
or UO_378 (O_378,N_9752,N_9783);
nor UO_379 (O_379,N_9873,N_9672);
or UO_380 (O_380,N_9935,N_9910);
xor UO_381 (O_381,N_9514,N_9896);
or UO_382 (O_382,N_9542,N_9892);
nor UO_383 (O_383,N_9925,N_9581);
xor UO_384 (O_384,N_9831,N_9661);
xor UO_385 (O_385,N_9732,N_9760);
xor UO_386 (O_386,N_9815,N_9875);
nor UO_387 (O_387,N_9776,N_9703);
xor UO_388 (O_388,N_9715,N_9692);
and UO_389 (O_389,N_9711,N_9502);
nand UO_390 (O_390,N_9904,N_9778);
nand UO_391 (O_391,N_9659,N_9641);
nor UO_392 (O_392,N_9777,N_9612);
and UO_393 (O_393,N_9966,N_9986);
or UO_394 (O_394,N_9693,N_9519);
xnor UO_395 (O_395,N_9808,N_9706);
or UO_396 (O_396,N_9710,N_9859);
nand UO_397 (O_397,N_9771,N_9991);
and UO_398 (O_398,N_9812,N_9914);
nor UO_399 (O_399,N_9541,N_9609);
nor UO_400 (O_400,N_9870,N_9700);
or UO_401 (O_401,N_9857,N_9710);
nor UO_402 (O_402,N_9565,N_9841);
and UO_403 (O_403,N_9950,N_9974);
and UO_404 (O_404,N_9719,N_9619);
and UO_405 (O_405,N_9924,N_9944);
nand UO_406 (O_406,N_9647,N_9583);
or UO_407 (O_407,N_9889,N_9597);
and UO_408 (O_408,N_9684,N_9515);
or UO_409 (O_409,N_9507,N_9742);
and UO_410 (O_410,N_9618,N_9669);
nand UO_411 (O_411,N_9913,N_9749);
nand UO_412 (O_412,N_9500,N_9949);
and UO_413 (O_413,N_9626,N_9788);
nor UO_414 (O_414,N_9829,N_9720);
and UO_415 (O_415,N_9909,N_9838);
nand UO_416 (O_416,N_9606,N_9696);
nand UO_417 (O_417,N_9997,N_9781);
xnor UO_418 (O_418,N_9915,N_9653);
or UO_419 (O_419,N_9885,N_9998);
nand UO_420 (O_420,N_9884,N_9555);
nor UO_421 (O_421,N_9706,N_9531);
nor UO_422 (O_422,N_9976,N_9931);
and UO_423 (O_423,N_9529,N_9558);
nor UO_424 (O_424,N_9725,N_9510);
and UO_425 (O_425,N_9736,N_9608);
nor UO_426 (O_426,N_9861,N_9532);
nor UO_427 (O_427,N_9980,N_9628);
or UO_428 (O_428,N_9686,N_9736);
or UO_429 (O_429,N_9996,N_9719);
xor UO_430 (O_430,N_9798,N_9720);
xnor UO_431 (O_431,N_9598,N_9865);
and UO_432 (O_432,N_9603,N_9774);
nand UO_433 (O_433,N_9595,N_9980);
and UO_434 (O_434,N_9598,N_9925);
or UO_435 (O_435,N_9715,N_9884);
nor UO_436 (O_436,N_9608,N_9999);
or UO_437 (O_437,N_9534,N_9588);
or UO_438 (O_438,N_9817,N_9588);
xor UO_439 (O_439,N_9887,N_9685);
and UO_440 (O_440,N_9787,N_9553);
nand UO_441 (O_441,N_9786,N_9862);
nor UO_442 (O_442,N_9717,N_9695);
and UO_443 (O_443,N_9726,N_9900);
nand UO_444 (O_444,N_9822,N_9589);
xor UO_445 (O_445,N_9938,N_9525);
nand UO_446 (O_446,N_9625,N_9534);
xnor UO_447 (O_447,N_9686,N_9622);
or UO_448 (O_448,N_9855,N_9641);
or UO_449 (O_449,N_9631,N_9966);
or UO_450 (O_450,N_9522,N_9793);
xor UO_451 (O_451,N_9708,N_9804);
nand UO_452 (O_452,N_9644,N_9717);
or UO_453 (O_453,N_9823,N_9632);
or UO_454 (O_454,N_9613,N_9930);
xnor UO_455 (O_455,N_9786,N_9553);
nand UO_456 (O_456,N_9548,N_9775);
xor UO_457 (O_457,N_9502,N_9967);
or UO_458 (O_458,N_9571,N_9645);
or UO_459 (O_459,N_9783,N_9751);
xor UO_460 (O_460,N_9768,N_9835);
nand UO_461 (O_461,N_9856,N_9595);
and UO_462 (O_462,N_9917,N_9838);
nor UO_463 (O_463,N_9769,N_9755);
or UO_464 (O_464,N_9585,N_9899);
xor UO_465 (O_465,N_9687,N_9782);
and UO_466 (O_466,N_9803,N_9660);
and UO_467 (O_467,N_9878,N_9916);
and UO_468 (O_468,N_9981,N_9902);
nor UO_469 (O_469,N_9625,N_9786);
or UO_470 (O_470,N_9966,N_9640);
xnor UO_471 (O_471,N_9551,N_9547);
nor UO_472 (O_472,N_9949,N_9875);
xor UO_473 (O_473,N_9545,N_9616);
xnor UO_474 (O_474,N_9658,N_9625);
nor UO_475 (O_475,N_9555,N_9604);
nand UO_476 (O_476,N_9738,N_9977);
nor UO_477 (O_477,N_9634,N_9967);
xnor UO_478 (O_478,N_9559,N_9654);
nand UO_479 (O_479,N_9950,N_9534);
nand UO_480 (O_480,N_9775,N_9982);
nand UO_481 (O_481,N_9903,N_9503);
xor UO_482 (O_482,N_9781,N_9778);
nor UO_483 (O_483,N_9607,N_9886);
xor UO_484 (O_484,N_9814,N_9798);
nand UO_485 (O_485,N_9730,N_9984);
and UO_486 (O_486,N_9706,N_9719);
xnor UO_487 (O_487,N_9713,N_9695);
xnor UO_488 (O_488,N_9961,N_9941);
nand UO_489 (O_489,N_9868,N_9942);
nor UO_490 (O_490,N_9810,N_9918);
nand UO_491 (O_491,N_9928,N_9788);
or UO_492 (O_492,N_9516,N_9562);
nor UO_493 (O_493,N_9681,N_9998);
and UO_494 (O_494,N_9985,N_9824);
or UO_495 (O_495,N_9986,N_9699);
or UO_496 (O_496,N_9912,N_9949);
and UO_497 (O_497,N_9937,N_9915);
and UO_498 (O_498,N_9644,N_9804);
or UO_499 (O_499,N_9592,N_9951);
or UO_500 (O_500,N_9865,N_9876);
nand UO_501 (O_501,N_9906,N_9917);
nand UO_502 (O_502,N_9615,N_9577);
or UO_503 (O_503,N_9534,N_9500);
nor UO_504 (O_504,N_9679,N_9950);
nand UO_505 (O_505,N_9821,N_9992);
and UO_506 (O_506,N_9719,N_9854);
xnor UO_507 (O_507,N_9867,N_9811);
xnor UO_508 (O_508,N_9960,N_9997);
nor UO_509 (O_509,N_9897,N_9976);
nand UO_510 (O_510,N_9903,N_9713);
or UO_511 (O_511,N_9792,N_9672);
nor UO_512 (O_512,N_9753,N_9708);
and UO_513 (O_513,N_9924,N_9701);
nor UO_514 (O_514,N_9752,N_9556);
and UO_515 (O_515,N_9779,N_9626);
nand UO_516 (O_516,N_9761,N_9664);
xor UO_517 (O_517,N_9512,N_9669);
nor UO_518 (O_518,N_9622,N_9921);
xnor UO_519 (O_519,N_9888,N_9933);
and UO_520 (O_520,N_9504,N_9923);
or UO_521 (O_521,N_9504,N_9644);
and UO_522 (O_522,N_9648,N_9668);
or UO_523 (O_523,N_9723,N_9964);
nand UO_524 (O_524,N_9948,N_9563);
xor UO_525 (O_525,N_9781,N_9700);
nor UO_526 (O_526,N_9541,N_9945);
xnor UO_527 (O_527,N_9868,N_9508);
or UO_528 (O_528,N_9519,N_9556);
nor UO_529 (O_529,N_9810,N_9967);
nand UO_530 (O_530,N_9557,N_9506);
nor UO_531 (O_531,N_9830,N_9731);
nor UO_532 (O_532,N_9907,N_9661);
xor UO_533 (O_533,N_9775,N_9854);
or UO_534 (O_534,N_9914,N_9597);
and UO_535 (O_535,N_9975,N_9761);
xnor UO_536 (O_536,N_9988,N_9725);
xor UO_537 (O_537,N_9540,N_9541);
or UO_538 (O_538,N_9667,N_9698);
nand UO_539 (O_539,N_9974,N_9618);
nor UO_540 (O_540,N_9587,N_9604);
and UO_541 (O_541,N_9859,N_9783);
nand UO_542 (O_542,N_9818,N_9609);
or UO_543 (O_543,N_9909,N_9957);
nor UO_544 (O_544,N_9609,N_9660);
and UO_545 (O_545,N_9730,N_9788);
or UO_546 (O_546,N_9947,N_9563);
and UO_547 (O_547,N_9830,N_9882);
or UO_548 (O_548,N_9867,N_9935);
and UO_549 (O_549,N_9724,N_9556);
and UO_550 (O_550,N_9662,N_9913);
nand UO_551 (O_551,N_9742,N_9727);
or UO_552 (O_552,N_9743,N_9500);
nor UO_553 (O_553,N_9577,N_9831);
xnor UO_554 (O_554,N_9862,N_9522);
xor UO_555 (O_555,N_9913,N_9521);
nor UO_556 (O_556,N_9554,N_9720);
nor UO_557 (O_557,N_9905,N_9734);
nor UO_558 (O_558,N_9728,N_9941);
nand UO_559 (O_559,N_9831,N_9738);
xor UO_560 (O_560,N_9704,N_9805);
and UO_561 (O_561,N_9912,N_9574);
xor UO_562 (O_562,N_9604,N_9705);
nor UO_563 (O_563,N_9857,N_9515);
and UO_564 (O_564,N_9596,N_9890);
and UO_565 (O_565,N_9701,N_9630);
xor UO_566 (O_566,N_9959,N_9816);
nor UO_567 (O_567,N_9862,N_9934);
nand UO_568 (O_568,N_9570,N_9687);
nor UO_569 (O_569,N_9809,N_9927);
nor UO_570 (O_570,N_9876,N_9910);
and UO_571 (O_571,N_9981,N_9623);
xnor UO_572 (O_572,N_9918,N_9690);
nand UO_573 (O_573,N_9854,N_9831);
and UO_574 (O_574,N_9606,N_9536);
or UO_575 (O_575,N_9743,N_9889);
and UO_576 (O_576,N_9746,N_9867);
nor UO_577 (O_577,N_9871,N_9756);
nand UO_578 (O_578,N_9575,N_9958);
and UO_579 (O_579,N_9950,N_9762);
nor UO_580 (O_580,N_9992,N_9757);
xor UO_581 (O_581,N_9545,N_9981);
or UO_582 (O_582,N_9793,N_9535);
xor UO_583 (O_583,N_9643,N_9640);
nand UO_584 (O_584,N_9513,N_9936);
and UO_585 (O_585,N_9545,N_9982);
nor UO_586 (O_586,N_9586,N_9661);
xor UO_587 (O_587,N_9716,N_9521);
nand UO_588 (O_588,N_9561,N_9800);
xor UO_589 (O_589,N_9602,N_9753);
xor UO_590 (O_590,N_9853,N_9538);
nand UO_591 (O_591,N_9987,N_9741);
and UO_592 (O_592,N_9812,N_9816);
nor UO_593 (O_593,N_9733,N_9737);
and UO_594 (O_594,N_9622,N_9873);
nand UO_595 (O_595,N_9683,N_9928);
or UO_596 (O_596,N_9759,N_9800);
nand UO_597 (O_597,N_9531,N_9878);
or UO_598 (O_598,N_9799,N_9637);
and UO_599 (O_599,N_9832,N_9865);
or UO_600 (O_600,N_9560,N_9924);
and UO_601 (O_601,N_9955,N_9574);
nor UO_602 (O_602,N_9751,N_9943);
nand UO_603 (O_603,N_9779,N_9547);
nor UO_604 (O_604,N_9841,N_9735);
and UO_605 (O_605,N_9789,N_9941);
nand UO_606 (O_606,N_9669,N_9754);
xnor UO_607 (O_607,N_9776,N_9661);
nand UO_608 (O_608,N_9680,N_9618);
and UO_609 (O_609,N_9957,N_9890);
and UO_610 (O_610,N_9503,N_9812);
and UO_611 (O_611,N_9698,N_9629);
and UO_612 (O_612,N_9605,N_9579);
or UO_613 (O_613,N_9676,N_9776);
or UO_614 (O_614,N_9529,N_9644);
or UO_615 (O_615,N_9923,N_9516);
nor UO_616 (O_616,N_9874,N_9968);
xnor UO_617 (O_617,N_9837,N_9976);
nand UO_618 (O_618,N_9593,N_9501);
or UO_619 (O_619,N_9967,N_9508);
nand UO_620 (O_620,N_9887,N_9878);
nand UO_621 (O_621,N_9882,N_9707);
and UO_622 (O_622,N_9648,N_9991);
nand UO_623 (O_623,N_9974,N_9656);
nor UO_624 (O_624,N_9765,N_9772);
and UO_625 (O_625,N_9799,N_9872);
xor UO_626 (O_626,N_9869,N_9515);
nor UO_627 (O_627,N_9523,N_9565);
nor UO_628 (O_628,N_9567,N_9641);
xnor UO_629 (O_629,N_9873,N_9807);
xnor UO_630 (O_630,N_9608,N_9897);
nor UO_631 (O_631,N_9698,N_9763);
nand UO_632 (O_632,N_9639,N_9505);
and UO_633 (O_633,N_9872,N_9923);
or UO_634 (O_634,N_9602,N_9906);
nand UO_635 (O_635,N_9937,N_9562);
nand UO_636 (O_636,N_9663,N_9993);
nor UO_637 (O_637,N_9890,N_9997);
or UO_638 (O_638,N_9964,N_9861);
or UO_639 (O_639,N_9874,N_9528);
nor UO_640 (O_640,N_9980,N_9600);
xnor UO_641 (O_641,N_9648,N_9885);
xnor UO_642 (O_642,N_9589,N_9685);
nand UO_643 (O_643,N_9960,N_9993);
nor UO_644 (O_644,N_9653,N_9820);
nand UO_645 (O_645,N_9684,N_9809);
or UO_646 (O_646,N_9582,N_9818);
and UO_647 (O_647,N_9872,N_9734);
or UO_648 (O_648,N_9527,N_9535);
nor UO_649 (O_649,N_9706,N_9982);
or UO_650 (O_650,N_9855,N_9831);
and UO_651 (O_651,N_9959,N_9568);
xor UO_652 (O_652,N_9744,N_9971);
xnor UO_653 (O_653,N_9781,N_9595);
or UO_654 (O_654,N_9677,N_9740);
xnor UO_655 (O_655,N_9596,N_9510);
and UO_656 (O_656,N_9754,N_9890);
or UO_657 (O_657,N_9622,N_9699);
nand UO_658 (O_658,N_9713,N_9799);
and UO_659 (O_659,N_9765,N_9676);
nor UO_660 (O_660,N_9740,N_9500);
or UO_661 (O_661,N_9810,N_9671);
nor UO_662 (O_662,N_9852,N_9858);
and UO_663 (O_663,N_9960,N_9687);
and UO_664 (O_664,N_9564,N_9703);
and UO_665 (O_665,N_9512,N_9697);
nand UO_666 (O_666,N_9566,N_9662);
and UO_667 (O_667,N_9777,N_9983);
and UO_668 (O_668,N_9866,N_9743);
or UO_669 (O_669,N_9566,N_9754);
nand UO_670 (O_670,N_9990,N_9997);
xor UO_671 (O_671,N_9749,N_9547);
xnor UO_672 (O_672,N_9711,N_9601);
nand UO_673 (O_673,N_9851,N_9553);
or UO_674 (O_674,N_9832,N_9625);
or UO_675 (O_675,N_9959,N_9646);
and UO_676 (O_676,N_9935,N_9663);
nand UO_677 (O_677,N_9695,N_9602);
nand UO_678 (O_678,N_9993,N_9711);
and UO_679 (O_679,N_9864,N_9862);
xnor UO_680 (O_680,N_9572,N_9503);
xnor UO_681 (O_681,N_9542,N_9969);
nand UO_682 (O_682,N_9840,N_9778);
or UO_683 (O_683,N_9509,N_9723);
nand UO_684 (O_684,N_9888,N_9669);
or UO_685 (O_685,N_9984,N_9637);
xnor UO_686 (O_686,N_9580,N_9618);
or UO_687 (O_687,N_9695,N_9987);
and UO_688 (O_688,N_9967,N_9847);
nor UO_689 (O_689,N_9514,N_9539);
or UO_690 (O_690,N_9748,N_9687);
or UO_691 (O_691,N_9637,N_9942);
xnor UO_692 (O_692,N_9940,N_9598);
or UO_693 (O_693,N_9871,N_9833);
nor UO_694 (O_694,N_9811,N_9871);
nand UO_695 (O_695,N_9967,N_9933);
and UO_696 (O_696,N_9868,N_9672);
and UO_697 (O_697,N_9727,N_9534);
nand UO_698 (O_698,N_9799,N_9527);
or UO_699 (O_699,N_9908,N_9648);
or UO_700 (O_700,N_9866,N_9848);
or UO_701 (O_701,N_9718,N_9782);
and UO_702 (O_702,N_9826,N_9829);
nor UO_703 (O_703,N_9636,N_9563);
xor UO_704 (O_704,N_9793,N_9824);
nand UO_705 (O_705,N_9874,N_9784);
xnor UO_706 (O_706,N_9962,N_9653);
nor UO_707 (O_707,N_9542,N_9634);
nor UO_708 (O_708,N_9684,N_9975);
xnor UO_709 (O_709,N_9985,N_9792);
xor UO_710 (O_710,N_9935,N_9808);
or UO_711 (O_711,N_9897,N_9657);
nor UO_712 (O_712,N_9943,N_9771);
xnor UO_713 (O_713,N_9945,N_9535);
nand UO_714 (O_714,N_9940,N_9587);
and UO_715 (O_715,N_9985,N_9977);
nand UO_716 (O_716,N_9976,N_9832);
nor UO_717 (O_717,N_9553,N_9753);
nand UO_718 (O_718,N_9675,N_9910);
and UO_719 (O_719,N_9944,N_9648);
nand UO_720 (O_720,N_9708,N_9916);
nor UO_721 (O_721,N_9673,N_9591);
nor UO_722 (O_722,N_9958,N_9939);
or UO_723 (O_723,N_9879,N_9575);
xor UO_724 (O_724,N_9597,N_9966);
or UO_725 (O_725,N_9971,N_9590);
xnor UO_726 (O_726,N_9519,N_9543);
and UO_727 (O_727,N_9571,N_9827);
nor UO_728 (O_728,N_9519,N_9655);
nand UO_729 (O_729,N_9732,N_9906);
xnor UO_730 (O_730,N_9560,N_9725);
nor UO_731 (O_731,N_9645,N_9533);
nor UO_732 (O_732,N_9891,N_9665);
nand UO_733 (O_733,N_9989,N_9794);
and UO_734 (O_734,N_9697,N_9967);
nand UO_735 (O_735,N_9618,N_9563);
and UO_736 (O_736,N_9588,N_9587);
nand UO_737 (O_737,N_9694,N_9994);
xnor UO_738 (O_738,N_9934,N_9673);
nor UO_739 (O_739,N_9877,N_9945);
xnor UO_740 (O_740,N_9786,N_9722);
nand UO_741 (O_741,N_9698,N_9916);
and UO_742 (O_742,N_9584,N_9994);
xor UO_743 (O_743,N_9751,N_9750);
and UO_744 (O_744,N_9786,N_9692);
nand UO_745 (O_745,N_9873,N_9969);
xor UO_746 (O_746,N_9519,N_9970);
or UO_747 (O_747,N_9910,N_9791);
nand UO_748 (O_748,N_9508,N_9772);
or UO_749 (O_749,N_9927,N_9964);
and UO_750 (O_750,N_9695,N_9508);
or UO_751 (O_751,N_9663,N_9697);
xor UO_752 (O_752,N_9913,N_9947);
xor UO_753 (O_753,N_9594,N_9536);
nor UO_754 (O_754,N_9776,N_9748);
nor UO_755 (O_755,N_9735,N_9909);
xnor UO_756 (O_756,N_9603,N_9907);
or UO_757 (O_757,N_9808,N_9516);
xnor UO_758 (O_758,N_9529,N_9787);
and UO_759 (O_759,N_9746,N_9661);
or UO_760 (O_760,N_9716,N_9776);
nand UO_761 (O_761,N_9523,N_9596);
xnor UO_762 (O_762,N_9871,N_9740);
and UO_763 (O_763,N_9544,N_9811);
and UO_764 (O_764,N_9957,N_9619);
nand UO_765 (O_765,N_9655,N_9960);
xor UO_766 (O_766,N_9845,N_9736);
xnor UO_767 (O_767,N_9694,N_9697);
and UO_768 (O_768,N_9580,N_9648);
xor UO_769 (O_769,N_9520,N_9585);
or UO_770 (O_770,N_9652,N_9903);
xor UO_771 (O_771,N_9668,N_9623);
nor UO_772 (O_772,N_9584,N_9778);
or UO_773 (O_773,N_9841,N_9753);
xnor UO_774 (O_774,N_9857,N_9614);
and UO_775 (O_775,N_9536,N_9951);
or UO_776 (O_776,N_9689,N_9605);
nand UO_777 (O_777,N_9745,N_9855);
nor UO_778 (O_778,N_9629,N_9589);
nand UO_779 (O_779,N_9762,N_9559);
or UO_780 (O_780,N_9937,N_9732);
and UO_781 (O_781,N_9820,N_9908);
nand UO_782 (O_782,N_9821,N_9606);
nand UO_783 (O_783,N_9682,N_9689);
or UO_784 (O_784,N_9665,N_9599);
and UO_785 (O_785,N_9684,N_9766);
nor UO_786 (O_786,N_9635,N_9633);
xor UO_787 (O_787,N_9708,N_9874);
and UO_788 (O_788,N_9754,N_9707);
or UO_789 (O_789,N_9512,N_9840);
nand UO_790 (O_790,N_9917,N_9986);
xnor UO_791 (O_791,N_9571,N_9815);
xnor UO_792 (O_792,N_9760,N_9863);
or UO_793 (O_793,N_9840,N_9634);
or UO_794 (O_794,N_9987,N_9888);
nand UO_795 (O_795,N_9930,N_9605);
nor UO_796 (O_796,N_9937,N_9647);
nor UO_797 (O_797,N_9502,N_9896);
and UO_798 (O_798,N_9966,N_9574);
xor UO_799 (O_799,N_9523,N_9549);
nand UO_800 (O_800,N_9633,N_9775);
nor UO_801 (O_801,N_9985,N_9514);
nor UO_802 (O_802,N_9997,N_9929);
xor UO_803 (O_803,N_9833,N_9860);
and UO_804 (O_804,N_9600,N_9874);
xor UO_805 (O_805,N_9749,N_9757);
or UO_806 (O_806,N_9856,N_9591);
nor UO_807 (O_807,N_9882,N_9846);
or UO_808 (O_808,N_9811,N_9573);
xnor UO_809 (O_809,N_9559,N_9936);
or UO_810 (O_810,N_9784,N_9782);
nor UO_811 (O_811,N_9932,N_9970);
nor UO_812 (O_812,N_9861,N_9643);
nand UO_813 (O_813,N_9686,N_9884);
or UO_814 (O_814,N_9689,N_9817);
xnor UO_815 (O_815,N_9967,N_9630);
and UO_816 (O_816,N_9549,N_9997);
nand UO_817 (O_817,N_9543,N_9937);
xor UO_818 (O_818,N_9642,N_9658);
nand UO_819 (O_819,N_9651,N_9701);
or UO_820 (O_820,N_9592,N_9778);
or UO_821 (O_821,N_9717,N_9584);
xor UO_822 (O_822,N_9853,N_9950);
nor UO_823 (O_823,N_9831,N_9745);
and UO_824 (O_824,N_9754,N_9815);
and UO_825 (O_825,N_9914,N_9603);
nand UO_826 (O_826,N_9890,N_9952);
nor UO_827 (O_827,N_9524,N_9817);
nand UO_828 (O_828,N_9733,N_9990);
nor UO_829 (O_829,N_9803,N_9695);
nor UO_830 (O_830,N_9943,N_9795);
xor UO_831 (O_831,N_9668,N_9734);
xor UO_832 (O_832,N_9962,N_9701);
or UO_833 (O_833,N_9517,N_9789);
and UO_834 (O_834,N_9923,N_9806);
and UO_835 (O_835,N_9799,N_9928);
xnor UO_836 (O_836,N_9875,N_9684);
xnor UO_837 (O_837,N_9816,N_9516);
xor UO_838 (O_838,N_9974,N_9972);
and UO_839 (O_839,N_9813,N_9537);
or UO_840 (O_840,N_9910,N_9726);
nand UO_841 (O_841,N_9590,N_9596);
xnor UO_842 (O_842,N_9577,N_9755);
nand UO_843 (O_843,N_9726,N_9733);
xor UO_844 (O_844,N_9856,N_9980);
nand UO_845 (O_845,N_9677,N_9817);
nor UO_846 (O_846,N_9658,N_9871);
or UO_847 (O_847,N_9842,N_9734);
or UO_848 (O_848,N_9602,N_9611);
and UO_849 (O_849,N_9995,N_9618);
or UO_850 (O_850,N_9944,N_9925);
xnor UO_851 (O_851,N_9843,N_9892);
nand UO_852 (O_852,N_9830,N_9892);
or UO_853 (O_853,N_9760,N_9897);
or UO_854 (O_854,N_9604,N_9670);
xor UO_855 (O_855,N_9922,N_9749);
or UO_856 (O_856,N_9997,N_9523);
or UO_857 (O_857,N_9780,N_9600);
nor UO_858 (O_858,N_9869,N_9681);
and UO_859 (O_859,N_9504,N_9962);
nand UO_860 (O_860,N_9820,N_9806);
nand UO_861 (O_861,N_9585,N_9892);
and UO_862 (O_862,N_9718,N_9575);
xor UO_863 (O_863,N_9806,N_9659);
nand UO_864 (O_864,N_9898,N_9586);
xnor UO_865 (O_865,N_9808,N_9809);
nand UO_866 (O_866,N_9534,N_9993);
nand UO_867 (O_867,N_9589,N_9659);
xor UO_868 (O_868,N_9703,N_9800);
and UO_869 (O_869,N_9593,N_9799);
xor UO_870 (O_870,N_9859,N_9738);
and UO_871 (O_871,N_9646,N_9644);
xor UO_872 (O_872,N_9776,N_9580);
or UO_873 (O_873,N_9958,N_9790);
and UO_874 (O_874,N_9786,N_9579);
or UO_875 (O_875,N_9882,N_9685);
xor UO_876 (O_876,N_9859,N_9838);
xor UO_877 (O_877,N_9582,N_9580);
xnor UO_878 (O_878,N_9937,N_9713);
or UO_879 (O_879,N_9582,N_9754);
or UO_880 (O_880,N_9795,N_9636);
nor UO_881 (O_881,N_9656,N_9756);
nor UO_882 (O_882,N_9674,N_9530);
and UO_883 (O_883,N_9555,N_9881);
xnor UO_884 (O_884,N_9826,N_9628);
and UO_885 (O_885,N_9823,N_9839);
nor UO_886 (O_886,N_9716,N_9884);
and UO_887 (O_887,N_9779,N_9688);
and UO_888 (O_888,N_9913,N_9844);
nand UO_889 (O_889,N_9601,N_9991);
or UO_890 (O_890,N_9671,N_9543);
and UO_891 (O_891,N_9736,N_9668);
nand UO_892 (O_892,N_9791,N_9772);
and UO_893 (O_893,N_9844,N_9867);
and UO_894 (O_894,N_9731,N_9935);
nor UO_895 (O_895,N_9576,N_9844);
nor UO_896 (O_896,N_9993,N_9580);
xor UO_897 (O_897,N_9773,N_9744);
xnor UO_898 (O_898,N_9770,N_9780);
or UO_899 (O_899,N_9849,N_9974);
and UO_900 (O_900,N_9793,N_9907);
nor UO_901 (O_901,N_9653,N_9655);
or UO_902 (O_902,N_9598,N_9700);
xor UO_903 (O_903,N_9620,N_9587);
nand UO_904 (O_904,N_9626,N_9930);
or UO_905 (O_905,N_9981,N_9583);
or UO_906 (O_906,N_9812,N_9839);
xor UO_907 (O_907,N_9666,N_9766);
and UO_908 (O_908,N_9884,N_9653);
nor UO_909 (O_909,N_9956,N_9863);
and UO_910 (O_910,N_9886,N_9626);
or UO_911 (O_911,N_9706,N_9760);
xnor UO_912 (O_912,N_9803,N_9919);
and UO_913 (O_913,N_9596,N_9945);
nor UO_914 (O_914,N_9833,N_9576);
nand UO_915 (O_915,N_9935,N_9933);
or UO_916 (O_916,N_9567,N_9698);
xor UO_917 (O_917,N_9990,N_9686);
or UO_918 (O_918,N_9514,N_9880);
or UO_919 (O_919,N_9961,N_9882);
and UO_920 (O_920,N_9723,N_9962);
nand UO_921 (O_921,N_9727,N_9794);
or UO_922 (O_922,N_9525,N_9764);
nand UO_923 (O_923,N_9675,N_9819);
nor UO_924 (O_924,N_9744,N_9912);
or UO_925 (O_925,N_9924,N_9950);
and UO_926 (O_926,N_9785,N_9940);
xnor UO_927 (O_927,N_9812,N_9668);
nand UO_928 (O_928,N_9843,N_9937);
and UO_929 (O_929,N_9950,N_9609);
xor UO_930 (O_930,N_9521,N_9731);
xnor UO_931 (O_931,N_9976,N_9972);
nor UO_932 (O_932,N_9860,N_9817);
nand UO_933 (O_933,N_9819,N_9542);
and UO_934 (O_934,N_9816,N_9712);
xor UO_935 (O_935,N_9646,N_9657);
or UO_936 (O_936,N_9792,N_9622);
or UO_937 (O_937,N_9742,N_9745);
nand UO_938 (O_938,N_9857,N_9940);
xnor UO_939 (O_939,N_9933,N_9837);
nand UO_940 (O_940,N_9606,N_9907);
nand UO_941 (O_941,N_9609,N_9883);
and UO_942 (O_942,N_9690,N_9672);
nor UO_943 (O_943,N_9815,N_9817);
nor UO_944 (O_944,N_9851,N_9833);
or UO_945 (O_945,N_9981,N_9953);
or UO_946 (O_946,N_9508,N_9786);
nand UO_947 (O_947,N_9737,N_9603);
xnor UO_948 (O_948,N_9719,N_9807);
xor UO_949 (O_949,N_9783,N_9830);
nor UO_950 (O_950,N_9743,N_9566);
or UO_951 (O_951,N_9930,N_9843);
nand UO_952 (O_952,N_9543,N_9649);
nand UO_953 (O_953,N_9679,N_9561);
and UO_954 (O_954,N_9840,N_9758);
or UO_955 (O_955,N_9506,N_9678);
or UO_956 (O_956,N_9959,N_9715);
xor UO_957 (O_957,N_9605,N_9794);
xnor UO_958 (O_958,N_9862,N_9855);
nand UO_959 (O_959,N_9882,N_9576);
nand UO_960 (O_960,N_9944,N_9503);
nand UO_961 (O_961,N_9719,N_9986);
xnor UO_962 (O_962,N_9674,N_9738);
and UO_963 (O_963,N_9718,N_9744);
and UO_964 (O_964,N_9712,N_9965);
nor UO_965 (O_965,N_9524,N_9716);
nor UO_966 (O_966,N_9617,N_9597);
or UO_967 (O_967,N_9642,N_9722);
nand UO_968 (O_968,N_9857,N_9891);
and UO_969 (O_969,N_9758,N_9993);
nand UO_970 (O_970,N_9704,N_9991);
xor UO_971 (O_971,N_9732,N_9920);
nor UO_972 (O_972,N_9674,N_9824);
and UO_973 (O_973,N_9522,N_9531);
and UO_974 (O_974,N_9884,N_9604);
nor UO_975 (O_975,N_9606,N_9889);
xnor UO_976 (O_976,N_9820,N_9744);
xnor UO_977 (O_977,N_9672,N_9962);
or UO_978 (O_978,N_9794,N_9830);
and UO_979 (O_979,N_9801,N_9673);
or UO_980 (O_980,N_9761,N_9869);
and UO_981 (O_981,N_9611,N_9900);
nand UO_982 (O_982,N_9629,N_9713);
nor UO_983 (O_983,N_9977,N_9942);
or UO_984 (O_984,N_9614,N_9647);
or UO_985 (O_985,N_9908,N_9534);
nor UO_986 (O_986,N_9893,N_9629);
nand UO_987 (O_987,N_9752,N_9874);
or UO_988 (O_988,N_9623,N_9539);
nand UO_989 (O_989,N_9738,N_9603);
and UO_990 (O_990,N_9972,N_9853);
nand UO_991 (O_991,N_9627,N_9548);
nor UO_992 (O_992,N_9632,N_9946);
nand UO_993 (O_993,N_9869,N_9822);
nor UO_994 (O_994,N_9609,N_9911);
nor UO_995 (O_995,N_9980,N_9692);
and UO_996 (O_996,N_9923,N_9665);
xor UO_997 (O_997,N_9634,N_9637);
xor UO_998 (O_998,N_9544,N_9913);
xor UO_999 (O_999,N_9923,N_9796);
and UO_1000 (O_1000,N_9560,N_9513);
and UO_1001 (O_1001,N_9889,N_9977);
xor UO_1002 (O_1002,N_9575,N_9750);
or UO_1003 (O_1003,N_9703,N_9736);
nand UO_1004 (O_1004,N_9857,N_9643);
and UO_1005 (O_1005,N_9797,N_9956);
xnor UO_1006 (O_1006,N_9840,N_9781);
or UO_1007 (O_1007,N_9691,N_9960);
xnor UO_1008 (O_1008,N_9898,N_9977);
or UO_1009 (O_1009,N_9910,N_9546);
nor UO_1010 (O_1010,N_9951,N_9919);
xor UO_1011 (O_1011,N_9751,N_9947);
nor UO_1012 (O_1012,N_9674,N_9596);
or UO_1013 (O_1013,N_9557,N_9606);
and UO_1014 (O_1014,N_9930,N_9822);
nor UO_1015 (O_1015,N_9770,N_9602);
and UO_1016 (O_1016,N_9923,N_9873);
xnor UO_1017 (O_1017,N_9602,N_9797);
and UO_1018 (O_1018,N_9845,N_9501);
nand UO_1019 (O_1019,N_9620,N_9901);
or UO_1020 (O_1020,N_9638,N_9783);
nand UO_1021 (O_1021,N_9700,N_9922);
or UO_1022 (O_1022,N_9760,N_9620);
and UO_1023 (O_1023,N_9937,N_9750);
or UO_1024 (O_1024,N_9651,N_9542);
or UO_1025 (O_1025,N_9550,N_9583);
or UO_1026 (O_1026,N_9801,N_9990);
nor UO_1027 (O_1027,N_9956,N_9624);
or UO_1028 (O_1028,N_9607,N_9817);
nand UO_1029 (O_1029,N_9712,N_9544);
nand UO_1030 (O_1030,N_9732,N_9718);
xor UO_1031 (O_1031,N_9544,N_9526);
nand UO_1032 (O_1032,N_9847,N_9713);
nand UO_1033 (O_1033,N_9985,N_9856);
and UO_1034 (O_1034,N_9645,N_9588);
or UO_1035 (O_1035,N_9686,N_9701);
nand UO_1036 (O_1036,N_9792,N_9903);
nand UO_1037 (O_1037,N_9505,N_9605);
xor UO_1038 (O_1038,N_9585,N_9774);
nor UO_1039 (O_1039,N_9676,N_9970);
nor UO_1040 (O_1040,N_9723,N_9969);
nand UO_1041 (O_1041,N_9552,N_9667);
nand UO_1042 (O_1042,N_9760,N_9912);
or UO_1043 (O_1043,N_9877,N_9740);
nand UO_1044 (O_1044,N_9738,N_9755);
nand UO_1045 (O_1045,N_9887,N_9642);
nand UO_1046 (O_1046,N_9669,N_9563);
and UO_1047 (O_1047,N_9951,N_9644);
nand UO_1048 (O_1048,N_9647,N_9934);
nand UO_1049 (O_1049,N_9726,N_9723);
xnor UO_1050 (O_1050,N_9560,N_9834);
nor UO_1051 (O_1051,N_9680,N_9858);
and UO_1052 (O_1052,N_9886,N_9919);
nand UO_1053 (O_1053,N_9844,N_9649);
nor UO_1054 (O_1054,N_9778,N_9753);
xor UO_1055 (O_1055,N_9896,N_9849);
xnor UO_1056 (O_1056,N_9512,N_9936);
and UO_1057 (O_1057,N_9996,N_9544);
xor UO_1058 (O_1058,N_9773,N_9686);
or UO_1059 (O_1059,N_9503,N_9967);
or UO_1060 (O_1060,N_9771,N_9674);
and UO_1061 (O_1061,N_9967,N_9765);
nand UO_1062 (O_1062,N_9896,N_9735);
nor UO_1063 (O_1063,N_9983,N_9897);
nand UO_1064 (O_1064,N_9643,N_9581);
nor UO_1065 (O_1065,N_9816,N_9738);
and UO_1066 (O_1066,N_9551,N_9596);
or UO_1067 (O_1067,N_9875,N_9868);
nor UO_1068 (O_1068,N_9876,N_9516);
nor UO_1069 (O_1069,N_9523,N_9656);
or UO_1070 (O_1070,N_9505,N_9851);
xnor UO_1071 (O_1071,N_9825,N_9582);
nand UO_1072 (O_1072,N_9783,N_9604);
and UO_1073 (O_1073,N_9735,N_9852);
xor UO_1074 (O_1074,N_9860,N_9856);
xor UO_1075 (O_1075,N_9856,N_9909);
nand UO_1076 (O_1076,N_9642,N_9790);
nand UO_1077 (O_1077,N_9719,N_9965);
xor UO_1078 (O_1078,N_9666,N_9784);
xnor UO_1079 (O_1079,N_9841,N_9636);
nor UO_1080 (O_1080,N_9647,N_9626);
and UO_1081 (O_1081,N_9696,N_9658);
nand UO_1082 (O_1082,N_9622,N_9641);
nand UO_1083 (O_1083,N_9725,N_9642);
nor UO_1084 (O_1084,N_9688,N_9804);
and UO_1085 (O_1085,N_9808,N_9858);
or UO_1086 (O_1086,N_9750,N_9648);
and UO_1087 (O_1087,N_9732,N_9504);
and UO_1088 (O_1088,N_9654,N_9552);
or UO_1089 (O_1089,N_9643,N_9651);
nor UO_1090 (O_1090,N_9597,N_9669);
xor UO_1091 (O_1091,N_9888,N_9591);
xor UO_1092 (O_1092,N_9626,N_9688);
and UO_1093 (O_1093,N_9873,N_9583);
nand UO_1094 (O_1094,N_9653,N_9558);
and UO_1095 (O_1095,N_9870,N_9977);
or UO_1096 (O_1096,N_9942,N_9716);
xnor UO_1097 (O_1097,N_9946,N_9888);
nand UO_1098 (O_1098,N_9979,N_9562);
nand UO_1099 (O_1099,N_9707,N_9538);
nor UO_1100 (O_1100,N_9955,N_9626);
nor UO_1101 (O_1101,N_9829,N_9995);
or UO_1102 (O_1102,N_9509,N_9953);
xor UO_1103 (O_1103,N_9635,N_9517);
nand UO_1104 (O_1104,N_9893,N_9777);
nand UO_1105 (O_1105,N_9910,N_9542);
nand UO_1106 (O_1106,N_9751,N_9739);
and UO_1107 (O_1107,N_9660,N_9944);
or UO_1108 (O_1108,N_9615,N_9721);
and UO_1109 (O_1109,N_9954,N_9512);
nand UO_1110 (O_1110,N_9950,N_9688);
nand UO_1111 (O_1111,N_9596,N_9895);
or UO_1112 (O_1112,N_9864,N_9914);
and UO_1113 (O_1113,N_9927,N_9658);
nor UO_1114 (O_1114,N_9715,N_9784);
xor UO_1115 (O_1115,N_9866,N_9832);
nand UO_1116 (O_1116,N_9943,N_9817);
xnor UO_1117 (O_1117,N_9567,N_9722);
and UO_1118 (O_1118,N_9888,N_9755);
or UO_1119 (O_1119,N_9538,N_9747);
nand UO_1120 (O_1120,N_9762,N_9673);
or UO_1121 (O_1121,N_9807,N_9724);
xnor UO_1122 (O_1122,N_9825,N_9556);
nand UO_1123 (O_1123,N_9766,N_9621);
and UO_1124 (O_1124,N_9881,N_9896);
nor UO_1125 (O_1125,N_9899,N_9706);
and UO_1126 (O_1126,N_9750,N_9563);
nor UO_1127 (O_1127,N_9832,N_9951);
nor UO_1128 (O_1128,N_9706,N_9756);
or UO_1129 (O_1129,N_9551,N_9892);
and UO_1130 (O_1130,N_9894,N_9709);
nor UO_1131 (O_1131,N_9983,N_9793);
xor UO_1132 (O_1132,N_9567,N_9715);
nor UO_1133 (O_1133,N_9939,N_9926);
xor UO_1134 (O_1134,N_9890,N_9981);
and UO_1135 (O_1135,N_9975,N_9648);
xor UO_1136 (O_1136,N_9804,N_9640);
nand UO_1137 (O_1137,N_9908,N_9984);
or UO_1138 (O_1138,N_9955,N_9935);
nor UO_1139 (O_1139,N_9791,N_9749);
nand UO_1140 (O_1140,N_9886,N_9746);
xor UO_1141 (O_1141,N_9929,N_9539);
and UO_1142 (O_1142,N_9702,N_9676);
nand UO_1143 (O_1143,N_9513,N_9821);
nor UO_1144 (O_1144,N_9688,N_9658);
and UO_1145 (O_1145,N_9596,N_9604);
or UO_1146 (O_1146,N_9592,N_9583);
xnor UO_1147 (O_1147,N_9509,N_9990);
and UO_1148 (O_1148,N_9773,N_9865);
nor UO_1149 (O_1149,N_9959,N_9519);
nor UO_1150 (O_1150,N_9567,N_9703);
or UO_1151 (O_1151,N_9656,N_9847);
or UO_1152 (O_1152,N_9722,N_9619);
or UO_1153 (O_1153,N_9641,N_9529);
nor UO_1154 (O_1154,N_9736,N_9901);
and UO_1155 (O_1155,N_9672,N_9666);
or UO_1156 (O_1156,N_9744,N_9575);
xnor UO_1157 (O_1157,N_9982,N_9509);
and UO_1158 (O_1158,N_9818,N_9825);
nand UO_1159 (O_1159,N_9547,N_9902);
nand UO_1160 (O_1160,N_9788,N_9664);
nand UO_1161 (O_1161,N_9638,N_9660);
nand UO_1162 (O_1162,N_9878,N_9703);
or UO_1163 (O_1163,N_9902,N_9747);
nand UO_1164 (O_1164,N_9535,N_9770);
xnor UO_1165 (O_1165,N_9611,N_9669);
or UO_1166 (O_1166,N_9510,N_9931);
nand UO_1167 (O_1167,N_9815,N_9723);
or UO_1168 (O_1168,N_9502,N_9693);
xor UO_1169 (O_1169,N_9731,N_9863);
nand UO_1170 (O_1170,N_9563,N_9640);
or UO_1171 (O_1171,N_9826,N_9739);
xor UO_1172 (O_1172,N_9776,N_9972);
nor UO_1173 (O_1173,N_9779,N_9724);
or UO_1174 (O_1174,N_9851,N_9504);
or UO_1175 (O_1175,N_9682,N_9862);
and UO_1176 (O_1176,N_9690,N_9513);
xor UO_1177 (O_1177,N_9559,N_9715);
or UO_1178 (O_1178,N_9801,N_9963);
and UO_1179 (O_1179,N_9509,N_9976);
xor UO_1180 (O_1180,N_9624,N_9796);
and UO_1181 (O_1181,N_9547,N_9712);
nor UO_1182 (O_1182,N_9838,N_9701);
nor UO_1183 (O_1183,N_9679,N_9731);
and UO_1184 (O_1184,N_9839,N_9519);
nor UO_1185 (O_1185,N_9982,N_9836);
nor UO_1186 (O_1186,N_9678,N_9531);
nand UO_1187 (O_1187,N_9694,N_9602);
and UO_1188 (O_1188,N_9922,N_9509);
nand UO_1189 (O_1189,N_9757,N_9714);
xnor UO_1190 (O_1190,N_9816,N_9837);
xnor UO_1191 (O_1191,N_9886,N_9682);
or UO_1192 (O_1192,N_9601,N_9930);
nand UO_1193 (O_1193,N_9679,N_9570);
nand UO_1194 (O_1194,N_9967,N_9908);
or UO_1195 (O_1195,N_9615,N_9826);
and UO_1196 (O_1196,N_9944,N_9709);
xor UO_1197 (O_1197,N_9823,N_9518);
xnor UO_1198 (O_1198,N_9672,N_9602);
and UO_1199 (O_1199,N_9642,N_9788);
nor UO_1200 (O_1200,N_9634,N_9730);
nand UO_1201 (O_1201,N_9810,N_9939);
xnor UO_1202 (O_1202,N_9572,N_9927);
nand UO_1203 (O_1203,N_9506,N_9653);
or UO_1204 (O_1204,N_9605,N_9957);
xnor UO_1205 (O_1205,N_9544,N_9536);
and UO_1206 (O_1206,N_9949,N_9940);
nand UO_1207 (O_1207,N_9603,N_9677);
nor UO_1208 (O_1208,N_9786,N_9990);
and UO_1209 (O_1209,N_9547,N_9612);
nor UO_1210 (O_1210,N_9553,N_9860);
nor UO_1211 (O_1211,N_9721,N_9747);
or UO_1212 (O_1212,N_9941,N_9761);
or UO_1213 (O_1213,N_9882,N_9644);
nor UO_1214 (O_1214,N_9689,N_9766);
or UO_1215 (O_1215,N_9714,N_9512);
xor UO_1216 (O_1216,N_9546,N_9744);
xnor UO_1217 (O_1217,N_9603,N_9661);
nand UO_1218 (O_1218,N_9937,N_9679);
xor UO_1219 (O_1219,N_9857,N_9955);
nand UO_1220 (O_1220,N_9999,N_9788);
nor UO_1221 (O_1221,N_9754,N_9967);
xnor UO_1222 (O_1222,N_9941,N_9653);
nand UO_1223 (O_1223,N_9588,N_9843);
xor UO_1224 (O_1224,N_9642,N_9617);
xnor UO_1225 (O_1225,N_9909,N_9770);
nor UO_1226 (O_1226,N_9522,N_9920);
or UO_1227 (O_1227,N_9539,N_9728);
and UO_1228 (O_1228,N_9844,N_9971);
nand UO_1229 (O_1229,N_9649,N_9666);
xnor UO_1230 (O_1230,N_9567,N_9628);
xnor UO_1231 (O_1231,N_9839,N_9724);
nand UO_1232 (O_1232,N_9775,N_9688);
nand UO_1233 (O_1233,N_9567,N_9889);
xor UO_1234 (O_1234,N_9976,N_9581);
nand UO_1235 (O_1235,N_9628,N_9914);
xor UO_1236 (O_1236,N_9837,N_9877);
nand UO_1237 (O_1237,N_9770,N_9751);
and UO_1238 (O_1238,N_9797,N_9898);
or UO_1239 (O_1239,N_9767,N_9788);
and UO_1240 (O_1240,N_9625,N_9632);
and UO_1241 (O_1241,N_9735,N_9729);
or UO_1242 (O_1242,N_9760,N_9837);
or UO_1243 (O_1243,N_9973,N_9626);
or UO_1244 (O_1244,N_9756,N_9847);
nor UO_1245 (O_1245,N_9979,N_9691);
nor UO_1246 (O_1246,N_9632,N_9837);
xor UO_1247 (O_1247,N_9893,N_9543);
nor UO_1248 (O_1248,N_9641,N_9873);
nand UO_1249 (O_1249,N_9854,N_9707);
and UO_1250 (O_1250,N_9728,N_9598);
or UO_1251 (O_1251,N_9948,N_9534);
nand UO_1252 (O_1252,N_9636,N_9923);
xor UO_1253 (O_1253,N_9612,N_9969);
and UO_1254 (O_1254,N_9942,N_9839);
nand UO_1255 (O_1255,N_9688,N_9600);
or UO_1256 (O_1256,N_9935,N_9516);
xnor UO_1257 (O_1257,N_9831,N_9646);
nor UO_1258 (O_1258,N_9854,N_9694);
and UO_1259 (O_1259,N_9919,N_9907);
and UO_1260 (O_1260,N_9700,N_9690);
nor UO_1261 (O_1261,N_9724,N_9928);
or UO_1262 (O_1262,N_9801,N_9727);
nor UO_1263 (O_1263,N_9897,N_9831);
and UO_1264 (O_1264,N_9942,N_9929);
nand UO_1265 (O_1265,N_9720,N_9807);
nor UO_1266 (O_1266,N_9824,N_9894);
nor UO_1267 (O_1267,N_9742,N_9911);
nand UO_1268 (O_1268,N_9694,N_9729);
and UO_1269 (O_1269,N_9558,N_9985);
xnor UO_1270 (O_1270,N_9961,N_9756);
nand UO_1271 (O_1271,N_9972,N_9702);
nor UO_1272 (O_1272,N_9882,N_9767);
nand UO_1273 (O_1273,N_9861,N_9990);
nor UO_1274 (O_1274,N_9972,N_9818);
xnor UO_1275 (O_1275,N_9687,N_9595);
and UO_1276 (O_1276,N_9874,N_9936);
nand UO_1277 (O_1277,N_9787,N_9923);
nand UO_1278 (O_1278,N_9541,N_9978);
and UO_1279 (O_1279,N_9997,N_9953);
and UO_1280 (O_1280,N_9948,N_9569);
and UO_1281 (O_1281,N_9585,N_9929);
and UO_1282 (O_1282,N_9885,N_9654);
nor UO_1283 (O_1283,N_9781,N_9986);
nand UO_1284 (O_1284,N_9634,N_9694);
and UO_1285 (O_1285,N_9509,N_9802);
or UO_1286 (O_1286,N_9975,N_9698);
xnor UO_1287 (O_1287,N_9612,N_9718);
or UO_1288 (O_1288,N_9886,N_9847);
xnor UO_1289 (O_1289,N_9762,N_9956);
or UO_1290 (O_1290,N_9833,N_9913);
and UO_1291 (O_1291,N_9878,N_9985);
nor UO_1292 (O_1292,N_9699,N_9927);
nand UO_1293 (O_1293,N_9694,N_9646);
xor UO_1294 (O_1294,N_9880,N_9990);
xnor UO_1295 (O_1295,N_9714,N_9607);
nor UO_1296 (O_1296,N_9582,N_9891);
nand UO_1297 (O_1297,N_9776,N_9890);
nor UO_1298 (O_1298,N_9639,N_9787);
nand UO_1299 (O_1299,N_9574,N_9546);
nor UO_1300 (O_1300,N_9682,N_9993);
xor UO_1301 (O_1301,N_9505,N_9938);
and UO_1302 (O_1302,N_9876,N_9617);
nand UO_1303 (O_1303,N_9778,N_9670);
or UO_1304 (O_1304,N_9719,N_9959);
and UO_1305 (O_1305,N_9839,N_9628);
nor UO_1306 (O_1306,N_9923,N_9592);
and UO_1307 (O_1307,N_9624,N_9677);
or UO_1308 (O_1308,N_9564,N_9975);
nand UO_1309 (O_1309,N_9716,N_9929);
and UO_1310 (O_1310,N_9581,N_9702);
xor UO_1311 (O_1311,N_9899,N_9653);
and UO_1312 (O_1312,N_9616,N_9558);
nor UO_1313 (O_1313,N_9905,N_9896);
nor UO_1314 (O_1314,N_9643,N_9979);
nand UO_1315 (O_1315,N_9873,N_9944);
nand UO_1316 (O_1316,N_9667,N_9823);
or UO_1317 (O_1317,N_9705,N_9567);
or UO_1318 (O_1318,N_9750,N_9772);
nand UO_1319 (O_1319,N_9730,N_9605);
nand UO_1320 (O_1320,N_9801,N_9500);
nand UO_1321 (O_1321,N_9801,N_9785);
and UO_1322 (O_1322,N_9873,N_9564);
nand UO_1323 (O_1323,N_9831,N_9696);
and UO_1324 (O_1324,N_9785,N_9858);
nand UO_1325 (O_1325,N_9582,N_9539);
or UO_1326 (O_1326,N_9760,N_9832);
and UO_1327 (O_1327,N_9815,N_9519);
nor UO_1328 (O_1328,N_9535,N_9968);
nand UO_1329 (O_1329,N_9731,N_9873);
and UO_1330 (O_1330,N_9685,N_9697);
nor UO_1331 (O_1331,N_9959,N_9777);
and UO_1332 (O_1332,N_9754,N_9837);
xor UO_1333 (O_1333,N_9686,N_9942);
nor UO_1334 (O_1334,N_9735,N_9586);
nand UO_1335 (O_1335,N_9639,N_9847);
nand UO_1336 (O_1336,N_9873,N_9862);
xnor UO_1337 (O_1337,N_9715,N_9876);
and UO_1338 (O_1338,N_9556,N_9911);
nor UO_1339 (O_1339,N_9964,N_9863);
nor UO_1340 (O_1340,N_9534,N_9697);
nand UO_1341 (O_1341,N_9887,N_9832);
or UO_1342 (O_1342,N_9729,N_9891);
and UO_1343 (O_1343,N_9762,N_9657);
or UO_1344 (O_1344,N_9716,N_9867);
and UO_1345 (O_1345,N_9815,N_9888);
and UO_1346 (O_1346,N_9973,N_9822);
or UO_1347 (O_1347,N_9826,N_9979);
xor UO_1348 (O_1348,N_9662,N_9895);
nor UO_1349 (O_1349,N_9652,N_9800);
or UO_1350 (O_1350,N_9789,N_9980);
and UO_1351 (O_1351,N_9842,N_9833);
nor UO_1352 (O_1352,N_9576,N_9768);
nand UO_1353 (O_1353,N_9994,N_9701);
nand UO_1354 (O_1354,N_9523,N_9900);
xnor UO_1355 (O_1355,N_9628,N_9686);
or UO_1356 (O_1356,N_9709,N_9659);
or UO_1357 (O_1357,N_9544,N_9823);
nor UO_1358 (O_1358,N_9612,N_9887);
nand UO_1359 (O_1359,N_9875,N_9819);
nand UO_1360 (O_1360,N_9882,N_9819);
nand UO_1361 (O_1361,N_9606,N_9574);
nand UO_1362 (O_1362,N_9999,N_9594);
nand UO_1363 (O_1363,N_9646,N_9531);
and UO_1364 (O_1364,N_9590,N_9766);
xor UO_1365 (O_1365,N_9541,N_9600);
xnor UO_1366 (O_1366,N_9979,N_9820);
nand UO_1367 (O_1367,N_9572,N_9713);
or UO_1368 (O_1368,N_9842,N_9777);
nand UO_1369 (O_1369,N_9623,N_9959);
or UO_1370 (O_1370,N_9783,N_9969);
xnor UO_1371 (O_1371,N_9955,N_9689);
or UO_1372 (O_1372,N_9871,N_9545);
nand UO_1373 (O_1373,N_9948,N_9612);
xor UO_1374 (O_1374,N_9946,N_9772);
nand UO_1375 (O_1375,N_9766,N_9787);
or UO_1376 (O_1376,N_9515,N_9982);
and UO_1377 (O_1377,N_9714,N_9699);
nor UO_1378 (O_1378,N_9809,N_9876);
and UO_1379 (O_1379,N_9942,N_9905);
nand UO_1380 (O_1380,N_9552,N_9633);
or UO_1381 (O_1381,N_9729,N_9522);
and UO_1382 (O_1382,N_9926,N_9603);
nor UO_1383 (O_1383,N_9527,N_9798);
and UO_1384 (O_1384,N_9815,N_9818);
or UO_1385 (O_1385,N_9745,N_9841);
and UO_1386 (O_1386,N_9538,N_9662);
nor UO_1387 (O_1387,N_9778,N_9980);
xnor UO_1388 (O_1388,N_9916,N_9794);
and UO_1389 (O_1389,N_9633,N_9551);
or UO_1390 (O_1390,N_9607,N_9891);
nor UO_1391 (O_1391,N_9653,N_9796);
xor UO_1392 (O_1392,N_9563,N_9776);
or UO_1393 (O_1393,N_9753,N_9945);
xnor UO_1394 (O_1394,N_9704,N_9585);
and UO_1395 (O_1395,N_9743,N_9956);
nand UO_1396 (O_1396,N_9557,N_9940);
and UO_1397 (O_1397,N_9884,N_9773);
nor UO_1398 (O_1398,N_9972,N_9515);
xor UO_1399 (O_1399,N_9919,N_9755);
xor UO_1400 (O_1400,N_9904,N_9563);
nand UO_1401 (O_1401,N_9672,N_9647);
nor UO_1402 (O_1402,N_9875,N_9717);
xor UO_1403 (O_1403,N_9691,N_9936);
xor UO_1404 (O_1404,N_9834,N_9637);
nor UO_1405 (O_1405,N_9996,N_9947);
xor UO_1406 (O_1406,N_9526,N_9861);
nor UO_1407 (O_1407,N_9798,N_9768);
and UO_1408 (O_1408,N_9927,N_9742);
and UO_1409 (O_1409,N_9917,N_9589);
and UO_1410 (O_1410,N_9777,N_9598);
nand UO_1411 (O_1411,N_9848,N_9791);
nor UO_1412 (O_1412,N_9981,N_9820);
nand UO_1413 (O_1413,N_9615,N_9624);
nor UO_1414 (O_1414,N_9837,N_9939);
or UO_1415 (O_1415,N_9829,N_9568);
or UO_1416 (O_1416,N_9655,N_9711);
or UO_1417 (O_1417,N_9827,N_9630);
xor UO_1418 (O_1418,N_9588,N_9637);
or UO_1419 (O_1419,N_9535,N_9548);
nor UO_1420 (O_1420,N_9940,N_9946);
nand UO_1421 (O_1421,N_9526,N_9853);
and UO_1422 (O_1422,N_9564,N_9842);
or UO_1423 (O_1423,N_9987,N_9561);
xor UO_1424 (O_1424,N_9846,N_9564);
nand UO_1425 (O_1425,N_9587,N_9597);
nand UO_1426 (O_1426,N_9787,N_9966);
or UO_1427 (O_1427,N_9987,N_9644);
or UO_1428 (O_1428,N_9631,N_9941);
nor UO_1429 (O_1429,N_9576,N_9977);
nand UO_1430 (O_1430,N_9926,N_9863);
and UO_1431 (O_1431,N_9747,N_9594);
nand UO_1432 (O_1432,N_9686,N_9877);
nor UO_1433 (O_1433,N_9557,N_9847);
nor UO_1434 (O_1434,N_9653,N_9782);
and UO_1435 (O_1435,N_9819,N_9985);
nor UO_1436 (O_1436,N_9594,N_9590);
nand UO_1437 (O_1437,N_9947,N_9506);
nor UO_1438 (O_1438,N_9567,N_9569);
xnor UO_1439 (O_1439,N_9719,N_9579);
or UO_1440 (O_1440,N_9968,N_9665);
nand UO_1441 (O_1441,N_9964,N_9854);
and UO_1442 (O_1442,N_9709,N_9629);
and UO_1443 (O_1443,N_9521,N_9929);
xor UO_1444 (O_1444,N_9660,N_9646);
xor UO_1445 (O_1445,N_9853,N_9981);
nand UO_1446 (O_1446,N_9547,N_9513);
and UO_1447 (O_1447,N_9900,N_9793);
nand UO_1448 (O_1448,N_9840,N_9917);
nand UO_1449 (O_1449,N_9632,N_9704);
or UO_1450 (O_1450,N_9830,N_9524);
xnor UO_1451 (O_1451,N_9510,N_9899);
or UO_1452 (O_1452,N_9660,N_9828);
xnor UO_1453 (O_1453,N_9502,N_9597);
xor UO_1454 (O_1454,N_9752,N_9625);
and UO_1455 (O_1455,N_9657,N_9743);
nand UO_1456 (O_1456,N_9525,N_9864);
xor UO_1457 (O_1457,N_9936,N_9765);
nand UO_1458 (O_1458,N_9705,N_9942);
or UO_1459 (O_1459,N_9850,N_9783);
and UO_1460 (O_1460,N_9830,N_9862);
and UO_1461 (O_1461,N_9743,N_9703);
nor UO_1462 (O_1462,N_9662,N_9816);
nor UO_1463 (O_1463,N_9527,N_9659);
or UO_1464 (O_1464,N_9880,N_9867);
or UO_1465 (O_1465,N_9842,N_9613);
nor UO_1466 (O_1466,N_9688,N_9629);
xnor UO_1467 (O_1467,N_9813,N_9680);
and UO_1468 (O_1468,N_9851,N_9778);
or UO_1469 (O_1469,N_9890,N_9974);
nor UO_1470 (O_1470,N_9678,N_9545);
and UO_1471 (O_1471,N_9630,N_9562);
xor UO_1472 (O_1472,N_9898,N_9546);
and UO_1473 (O_1473,N_9987,N_9898);
xnor UO_1474 (O_1474,N_9687,N_9673);
and UO_1475 (O_1475,N_9569,N_9902);
or UO_1476 (O_1476,N_9902,N_9857);
xor UO_1477 (O_1477,N_9635,N_9694);
or UO_1478 (O_1478,N_9685,N_9922);
xnor UO_1479 (O_1479,N_9716,N_9996);
xnor UO_1480 (O_1480,N_9535,N_9560);
xor UO_1481 (O_1481,N_9552,N_9885);
or UO_1482 (O_1482,N_9646,N_9978);
and UO_1483 (O_1483,N_9969,N_9744);
nor UO_1484 (O_1484,N_9847,N_9820);
nor UO_1485 (O_1485,N_9812,N_9656);
nand UO_1486 (O_1486,N_9607,N_9832);
nand UO_1487 (O_1487,N_9810,N_9934);
xnor UO_1488 (O_1488,N_9844,N_9533);
or UO_1489 (O_1489,N_9921,N_9653);
nor UO_1490 (O_1490,N_9849,N_9853);
nor UO_1491 (O_1491,N_9704,N_9504);
or UO_1492 (O_1492,N_9806,N_9591);
and UO_1493 (O_1493,N_9756,N_9551);
xor UO_1494 (O_1494,N_9710,N_9702);
xor UO_1495 (O_1495,N_9868,N_9617);
nor UO_1496 (O_1496,N_9835,N_9585);
xnor UO_1497 (O_1497,N_9784,N_9949);
nor UO_1498 (O_1498,N_9501,N_9968);
and UO_1499 (O_1499,N_9811,N_9724);
endmodule